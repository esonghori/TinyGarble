
module hamming ( x, y, o );
  input [1599:0] x;
  input [1599:0] y;
  output [10:0] o;
  wire   n38259, n38260, n38261, n38262, n38263, n38264, n38265, n38266,
         n38267, n38268, n38269, n38270, n38271, n38272, n38273, n38274,
         n38275, n38276, n38277, n38278, n38279, n38280, n38281, n38282,
         n38283, n38284, n38285, n38286, n38287, n38288, n38289, n38290,
         n38291, n38292, n38293, n38294, n38295, n38296, n38297, n38298,
         n38299, n38300, n38301, n38302, n38303, n38304, n38305, n38306,
         n38307, n38308, n38309, n38310, n38311, n38312, n38313, n38314,
         n38315, n38316, n38317, n38318, n38319, n38320, n38321, n38322,
         n38323, n38324, n38325, n38326, n38327, n38328, n38329, n38330,
         n38331, n38332, n38333, n38334, n38335, n38336, n38337, n38338,
         n38339, n38340, n38341, n38342, n38343, n38344, n38345, n38346,
         n38347, n38348, n38349, n38350, n38351, n38352, n38353, n38354,
         n38355, n38356, n38357, n38358, n38359, n38360, n38361, n38362,
         n38363, n38364, n38365, n38366, n38367, n38368, n38369, n38370,
         n38371, n38372, n38373, n38374, n38375, n38376, n38377, n38378,
         n38379, n38380, n38381, n38382, n38383, n38384, n38385, n38386,
         n38387, n38388, n38389, n38390, n38391, n38392, n38393, n38394,
         n38395, n38396, n38397, n38398, n38399, n38400, n38401, n38402,
         n38403, n38404, n38405, n38406, n38407, n38408, n38409, n38410,
         n38411, n38412, n38413, n38414, n38415, n38416, n38417, n38418,
         n38419, n38420, n38421, n38422, n38423, n38424, n38425, n38426,
         n38427, n38428, n38429, n38430, n38431, n38432, n38433, n38434,
         n38435, n38436, n38437, n38438, n38439, n38440, n38441, n38442,
         n38443, n38444, n38445, n38446, n38447, n38448, n38449, n38450,
         n38451, n38452, n38453, n38454, n38455, n38456, n38457, n38458,
         n38459, n38460, n38461, n38462, n38463, n38464, n38465, n38466,
         n38467, n38468, n38469, n38470, n38471, n38472, n38473, n38474,
         n38475, n38476, n38477, n38478, n38479, n38480, n38481, n38482,
         n38483, n38484, n38485, n38486, n38487, n38488, n38489, n38490,
         n38491, n38492, n38493, n38494, n38495, n38496, n38497, n38498,
         n38499, n38500, n38501, n38502, n38503, n38504, n38505, n38506,
         n38507, n38508, n38509, n38510, n38511, n38512, n38513, n38514,
         n38515, n38516, n38517, n38518, n38519, n38520, n38521, n38522,
         n38523, n38524, n38525, n38526, n38527, n38528, n38529, n38530,
         n38531, n38532, n38533, n38534, n38535, n38536, n38537, n38538,
         n38539, n38540, n38541, n38542, n38543, n38544, n38545, n38546,
         n38547, n38548, n38549, n38550, n38551, n38552, n38553, n38554,
         n38555, n38556, n38557, n38558, n38559, n38560, n38561, n38562,
         n38563, n38564, n38565, n38566, n38567, n38568, n38569, n38570,
         n38571, n38572, n38573, n38574, n38575, n38576, n38577, n38578,
         n38579, n38580, n38581, n38582, n38583, n38584, n38585, n38586,
         n38587, n38588, n38589, n38590, n38591, n38592, n38593, n38594,
         n38595, n38596, n38597, n38598, n38599, n38600, n38601, n38602,
         n38603, n38604, n38605, n38606, n38607, n38608, n38609, n38610,
         n38611, n38612, n38613, n38614, n38615, n38616, n38617, n38618,
         n38619, n38620, n38621, n38622, n38623, n38624, n38625, n38626,
         n38627, n38628, n38629, n38630, n38631, n38632, n38633, n38634,
         n38635, n38636, n38637, n38638, n38639, n38640, n38641, n38642,
         n38643, n38644, n38645, n38646, n38647, n38648, n38649, n38650,
         n38651, n38652, n38653, n38654, n38655, n38656, n38657, n38658,
         n38659, n38660, n38661, n38662, n38663, n38664, n38665, n38666,
         n38667, n38668, n38669, n38670, n38671, n38672, n38673, n38674,
         n38675, n38676, n38677, n38678, n38679, n38680, n38681, n38682,
         n38683, n38684, n38685, n38686, n38687, n38688, n38689, n38690,
         n38691, n38692, n38693, n38694, n38695, n38696, n38697, n38698,
         n38699, n38700, n38701, n38702, n38703, n38704, n38705, n38706,
         n38707, n38708, n38709, n38710, n38711, n38712, n38713, n38714,
         n38715, n38716, n38717, n38718, n38719, n38720, n38721, n38722,
         n38723, n38724, n38725, n38726, n38727, n38728, n38729, n38730,
         n38731, n38732, n38733, n38734, n38735, n38736, n38737, n38738,
         n38739, n38740, n38741, n38742, n38743, n38744, n38745, n38746,
         n38747, n38748, n38749, n38750, n38751, n38752, n38753, n38754,
         n38755, n38756, n38757, n38758, n38759, n38760, n38761, n38762,
         n38763, n38764, n38765, n38766, n38767, n38768, n38769, n38770,
         n38771, n38772, n38773, n38774, n38775, n38776, n38777, n38778,
         n38779, n38780, n38781, n38782, n38783, n38784, n38785, n38786,
         n38787, n38788, n38789, n38790, n38791, n38792, n38793, n38794,
         n38795, n38796, n38797, n38798, n38799, n38800, n38801, n38802,
         n38803, n38804, n38805, n38806, n38807, n38808, n38809, n38810,
         n38811, n38812, n38813, n38814, n38815, n38816, n38817, n38818,
         n38819, n38820, n38821, n38822, n38823, n38824, n38825, n38826,
         n38827, n38828, n38829, n38830, n38831, n38832, n38833, n38834,
         n38835, n38836, n38837, n38838, n38839, n38840, n38841, n38842,
         n38843, n38844, n38845, n38846, n38847, n38848, n38849, n38850,
         n38851, n38852, n38853, n38854, n38855, n38856, n38857, n38858,
         n38859, n38860, n38861, n38862, n38863, n38864, n38865, n38866,
         n38867, n38868, n38869, n38870, n38871, n38872, n38873, n38874,
         n38875, n38876, n38877, n38878, n38879, n38880, n38881, n38882,
         n38883, n38884, n38885, n38886, n38887, n38888, n38889, n38890,
         n38891, n38892, n38893, n38894, n38895, n38896, n38897, n38898,
         n38899, n38900, n38901, n38902, n38903, n38904, n38905, n38906,
         n38907, n38908, n38909, n38910, n38911, n38912, n38913, n38914,
         n38915, n38916, n38917, n38918, n38919, n38920, n38921, n38922,
         n38923, n38924, n38925, n38926, n38927, n38928, n38929, n38930,
         n38931, n38932, n38933, n38934, n38935, n38936, n38937, n38938,
         n38939, n38940, n38941, n38942, n38943, n38944, n38945, n38946,
         n38947, n38948, n38949, n38950, n38951, n38952, n38953, n38954,
         n38955, n38956, n38957, n38958, n38959, n38960, n38961, n38962,
         n38963, n38964, n38965, n38966, n38967, n38968, n38969, n38970,
         n38971, n38972, n38973, n38974, n38975, n38976, n38977, n38978,
         n38979, n38980, n38981, n38982, n38983, n38984, n38985, n38986,
         n38987, n38988, n38989, n38990, n38991, n38992, n38993, n38994,
         n38995, n38996, n38997, n38998, n38999, n39000, n39001, n39002,
         n39003, n39004, n39005, n39006, n39007, n39008, n39009, n39010,
         n39011, n39012, n39013, n39014, n39015, n39016, n39017, n39018,
         n39019, n39020, n39021, n39022, n39023, n39024, n39025, n39026,
         n39027, n39028, n39029, n39030, n39031, n39032, n39033, n39034,
         n39035, n39036, n39037, n39038, n39039, n39040, n39041, n39042,
         n39043, n39044, n39045, n39046, n39047, n39048, n39049, n39050,
         n39051, n39052, n39053, n39054, n39055, n39056, n39057, n39058,
         n39059, n39060, n39061, n39062, n39063, n39064, n39065, n39066,
         n39067, n39068, n39069, n39070, n39071, n39072, n39073, n39074,
         n39075, n39076, n39077, n39078, n39079, n39080, n39081, n39082,
         n39083, n39084, n39085, n39086, n39087, n39088, n39089, n39090,
         n39091, n39092, n39093, n39094, n39095, n39096, n39097, n39098,
         n39099, n39100, n39101, n39102, n39103, n39104, n39105, n39106,
         n39107, n39108, n39109, n39110, n39111, n39112, n39113, n39114,
         n39115, n39116, n39117, n39118, n39119, n39120, n39121, n39122,
         n39123, n39124, n39125, n39126, n39127, n39128, n39129, n39130,
         n39131, n39132, n39133, n39134, n39135, n39136, n39137, n39138,
         n39139, n39140, n39141, n39142, n39143, n39144, n39145, n39146,
         n39147, n39148, n39149, n39150, n39151, n39152, n39153, n39154,
         n39155, n39156, n39157, n39158, n39159, n39160, n39161, n39162,
         n39163, n39164, n39165, n39166, n39167, n39168, n39169, n39170,
         n39171, n39172, n39173, n39174, n39175, n39176, n39177, n39178,
         n39179, n39180, n39181, n39182, n39183, n39184, n39185, n39186,
         n39187, n39188, n39189, n39190, n39191, n39192, n39193, n39194,
         n39195, n39196, n39197, n39198, n39199, n39200, n39201, n39202,
         n39203, n39204, n39205, n39206, n39207, n39208, n39209, n39210,
         n39211, n39212, n39213, n39214, n39215, n39216, n39217, n39218,
         n39219, n39220, n39221, n39222, n39223, n39224, n39225, n39226,
         n39227, n39228, n39229, n39230, n39231, n39232, n39233, n39234,
         n39235, n39236, n39237, n39238, n39239, n39240, n39241, n39242,
         n39243, n39244, n39245, n39246, n39247, n39248, n39249, n39250,
         n39251, n39252, n39253, n39254, n39255, n39256, n39257, n39258,
         n39259, n39260, n39261, n39262, n39263, n39264, n39265, n39266,
         n39267, n39268, n39269, n39270, n39271, n39272, n39273, n39274,
         n39275, n39276, n39277, n39278, n39279, n39280, n39281, n39282,
         n39283, n39284, n39285, n39286, n39287, n39288, n39289, n39290,
         n39291, n39292, n39293, n39294, n39295, n39296, n39297, n39298,
         n39299, n39300, n39301, n39302, n39303, n39304, n39305, n39306,
         n39307, n39308, n39309, n39310, n39311, n39312, n39313, n39314,
         n39315, n39316, n39317, n39318, n39319, n39320, n39321, n39322,
         n39323, n39324, n39325, n39326, n39327, n39328, n39329, n39330,
         n39331, n39332, n39333, n39334, n39335, n39336, n39337, n39338,
         n39339, n39340, n39341, n39342, n39343, n39344, n39345, n39346,
         n39347, n39348, n39349, n39350, n39351, n39352, n39353, n39354,
         n39355, n39356, n39357, n39358, n39359, n39360, n39361, n39362,
         n39363, n39364, n39365, n39366, n39367, n39368, n39369, n39370,
         n39371, n39372, n39373, n39374, n39375, n39376, n39377, n39378,
         n39379, n39380, n39381, n39382, n39383, n39384, n39385, n39386,
         n39387, n39388, n39389, n39390, n39391, n39392, n39393, n39394,
         n39395, n39396, n39397, n39398, n39399, n39400, n39401, n39402,
         n39403, n39404, n39405, n39406, n39407, n39408, n39409, n39410,
         n39411, n39412, n39413, n39414, n39415, n39416, n39417, n39418,
         n39419, n39420, n39421, n39422, n39423, n39424, n39425, n39426,
         n39427, n39428, n39429, n39430, n39431, n39432, n39433, n39434,
         n39435, n39436, n39437, n39438, n39439, n39440, n39441, n39442,
         n39443, n39444, n39445, n39446, n39447, n39448, n39449, n39450,
         n39451, n39452, n39453, n39454, n39455, n39456, n39457, n39458,
         n39459, n39460, n39461, n39462, n39463, n39464, n39465, n39466,
         n39467, n39468, n39469, n39470, n39471, n39472, n39473, n39474,
         n39475, n39476, n39477, n39478, n39479, n39480, n39481, n39482,
         n39483, n39484, n39485, n39486, n39487, n39488, n39489, n39490,
         n39491, n39492, n39493, n39494, n39495, n39496, n39497, n39498,
         n39499, n39500, n39501, n39502, n39503, n39504, n39505, n39506,
         n39507, n39508, n39509, n39510, n39511, n39512, n39513, n39514,
         n39515, n39516, n39517, n39518, n39519, n39520, n39521, n39522,
         n39523, n39524, n39525, n39526, n39527, n39528, n39529, n39530,
         n39531, n39532, n39533, n39534, n39535, n39536, n39537, n39538,
         n39539, n39540, n39541, n39542, n39543, n39544, n39545, n39546,
         n39547, n39548, n39549, n39550, n39551, n39552, n39553, n39554,
         n39555, n39556, n39557, n39558, n39559, n39560, n39561, n39562,
         n39563, n39564, n39565, n39566, n39567, n39568, n39569, n39570,
         n39571, n39572, n39573, n39574, n39575, n39576, n39577, n39578,
         n39579, n39580, n39581, n39582, n39583, n39584, n39585, n39586,
         n39587, n39588, n39589, n39590, n39591, n39592, n39593, n39594,
         n39595, n39596, n39597, n39598, n39599, n39600, n39601, n39602,
         n39603, n39604, n39605, n39606, n39607, n39608, n39609, n39610,
         n39611, n39612, n39613, n39614, n39615, n39616, n39617, n39618,
         n39619, n39620, n39621, n39622, n39623, n39624, n39625, n39626,
         n39627, n39628, n39629, n39630, n39631, n39632, n39633, n39634,
         n39635, n39636, n39637, n39638, n39639, n39640, n39641, n39642,
         n39643, n39644, n39645, n39646, n39647, n39648, n39649, n39650,
         n39651, n39652, n39653, n39654, n39655, n39656, n39657, n39658,
         n39659, n39660, n39661, n39662, n39663, n39664, n39665, n39666,
         n39667, n39668, n39669, n39670, n39671, n39672, n39673, n39674,
         n39675, n39676, n39677, n39678, n39679, n39680, n39681, n39682,
         n39683, n39684, n39685, n39686, n39687, n39688, n39689, n39690,
         n39691, n39692, n39693, n39694, n39695, n39696, n39697, n39698,
         n39699, n39700, n39701, n39702, n39703, n39704, n39705, n39706,
         n39707, n39708, n39709, n39710, n39711, n39712, n39713, n39714,
         n39715, n39716, n39717, n39718, n39719, n39720, n39721, n39722,
         n39723, n39724, n39725, n39726, n39727, n39728, n39729, n39730,
         n39731, n39732, n39733, n39734, n39735, n39736, n39737, n39738,
         n39739, n39740, n39741, n39742, n39743, n39744, n39745, n39746,
         n39747, n39748, n39749, n39750, n39751, n39752, n39753, n39754,
         n39755, n39756, n39757, n39758, n39759, n39760, n39761, n39762,
         n39763, n39764, n39765, n39766, n39767, n39768, n39769, n39770,
         n39771, n39772, n39773, n39774, n39775, n39776, n39777, n39778,
         n39779, n39780, n39781, n39782, n39783, n39784, n39785, n39786,
         n39787, n39788, n39789, n39790, n39791, n39792, n39793, n39794,
         n39795, n39796, n39797, n39798, n39799, n39800, n39801, n39802,
         n39803, n39804, n39805, n39806, n39807, n39808, n39809, n39810,
         n39811, n39812, n39813, n39814, n39815, n39816, n39817, n39818,
         n39819, n39820, n39821, n39822, n39823, n39824, n39825, n39826,
         n39827, n39828, n39829, n39830, n39831, n39832, n39833, n39834,
         n39835, n39836, n39837, n39838, n39839, n39840, n39841, n39842,
         n39843, n39844, n39845, n39846, n39847, n39848, n39849, n39850,
         n39851, n39852, n39853, n39854, n39855, n39856, n39857, n39858,
         n39859, n39860, n39861, n39862, n39863, n39864, n39865, n39866,
         n39867, n39868, n39869, n39870, n39871, n39872, n39873, n39874,
         n39875, n39876, n39877, n39878, n39879, n39880, n39881, n39882,
         n39883, n39884, n39885, n39886, n39887, n39888, n39889, n39890,
         n39891, n39892, n39893, n39894, n39895, n39896, n39897, n39898,
         n39899, n39900, n39901, n39902, n39903, n39904, n39905, n39906,
         n39907, n39908, n39909, n39910, n39911, n39912, n39913, n39914,
         n39915, n39916, n39917, n39918, n39919, n39920, n39921, n39922,
         n39923, n39924, n39925, n39926, n39927, n39928, n39929, n39930,
         n39931, n39932, n39933, n39934, n39935, n39936, n39937, n39938,
         n39939, n39940, n39941, n39942, n39943, n39944, n39945, n39946,
         n39947, n39948, n39949, n39950, n39951, n39952, n39953, n39954,
         n39955, n39956, n39957, n39958, n39959, n39960, n39961, n39962,
         n39963, n39964, n39965, n39966, n39967, n39968, n39969, n39970,
         n39971, n39972, n39973, n39974, n39975, n39976, n39977, n39978,
         n39979, n39980, n39981, n39982, n39983, n39984, n39985, n39986,
         n39987, n39988, n39989, n39990, n39991, n39992, n39993, n39994,
         n39995, n39996, n39997, n39998, n39999, n40000, n40001, n40002,
         n40003, n40004, n40005, n40006, n40007, n40008, n40009, n40010,
         n40011, n40012, n40013, n40014, n40015, n40016, n40017, n40018,
         n40019, n40020, n40021, n40022, n40023, n40024, n40025, n40026,
         n40027, n40028, n40029, n40030, n40031, n40032, n40033, n40034,
         n40035, n40036, n40037, n40038, n40039, n40040, n40041, n40042,
         n40043, n40044, n40045, n40046, n40047, n40048, n40049, n40050,
         n40051, n40052, n40053, n40054, n40055, n40056, n40057, n40058,
         n40059, n40060, n40061, n40062, n40063, n40064, n40065, n40066,
         n40067, n40068, n40069, n40070, n40071, n40072, n40073, n40074,
         n40075, n40076, n40077, n40078, n40079, n40080, n40081, n40082,
         n40083, n40084, n40085, n40086, n40087, n40088, n40089, n40090,
         n40091, n40092, n40093, n40094, n40095, n40096, n40097, n40098,
         n40099, n40100, n40101, n40102, n40103, n40104, n40105, n40106,
         n40107, n40108, n40109, n40110, n40111, n40112, n40113, n40114,
         n40115, n40116, n40117, n40118, n40119, n40120, n40121, n40122,
         n40123, n40124, n40125, n40126, n40127, n40128, n40129, n40130,
         n40131, n40132, n40133, n40134, n40135, n40136, n40137, n40138,
         n40139, n40140, n40141, n40142, n40143, n40144, n40145, n40146,
         n40147, n40148, n40149, n40150, n40151, n40152, n40153, n40154,
         n40155, n40156, n40157, n40158, n40159, n40160, n40161, n40162,
         n40163, n40164, n40165, n40166, n40167, n40168, n40169, n40170,
         n40171, n40172, n40173, n40174, n40175, n40176, n40177, n40178,
         n40179, n40180, n40181, n40182, n40183, n40184, n40185, n40186,
         n40187, n40188, n40189, n40190, n40191, n40192, n40193, n40194,
         n40195, n40196, n40197, n40198, n40199, n40200, n40201, n40202,
         n40203, n40204, n40205, n40206, n40207, n40208, n40209, n40210,
         n40211, n40212, n40213, n40214, n40215, n40216, n40217, n40218,
         n40219, n40220, n40221, n40222, n40223, n40224, n40225, n40226,
         n40227, n40228, n40229, n40230, n40231, n40232, n40233, n40234,
         n40235, n40236, n40237, n40238, n40239, n40240, n40241, n40242,
         n40243, n40244, n40245, n40246, n40247, n40248, n40249, n40250,
         n40251, n40252, n40253, n40254, n40255, n40256, n40257, n40258,
         n40259, n40260, n40261, n40262, n40263, n40264, n40265, n40266,
         n40267, n40268, n40269, n40270, n40271, n40272, n40273, n40274,
         n40275, n40276, n40277, n40278, n40279, n40280, n40281, n40282,
         n40283, n40284, n40285, n40286, n40287, n40288, n40289, n40290,
         n40291, n40292, n40293, n40294, n40295, n40296, n40297, n40298,
         n40299, n40300, n40301, n40302, n40303, n40304, n40305, n40306,
         n40307, n40308, n40309, n40310, n40311, n40312, n40313, n40314,
         n40315, n40316, n40317, n40318, n40319, n40320, n40321, n40322,
         n40323, n40324, n40325, n40326, n40327, n40328, n40329, n40330,
         n40331, n40332, n40333, n40334, n40335, n40336, n40337, n40338,
         n40339, n40340, n40341, n40342, n40343, n40344, n40345, n40346,
         n40347, n40348, n40349, n40350, n40351, n40352, n40353, n40354,
         n40355, n40356, n40357, n40358, n40359, n40360, n40361, n40362,
         n40363, n40364, n40365, n40366, n40367, n40368, n40369, n40370,
         n40371, n40372, n40373, n40374, n40375, n40376, n40377, n40378,
         n40379, n40380, n40381, n40382, n40383, n40384, n40385, n40386,
         n40387, n40388, n40389, n40390, n40391, n40392, n40393, n40394,
         n40395, n40396, n40397, n40398, n40399, n40400, n40401, n40402,
         n40403, n40404, n40405, n40406, n40407, n40408, n40409, n40410,
         n40411, n40412, n40413, n40414, n40415, n40416, n40417, n40418,
         n40419, n40420, n40421, n40422, n40423, n40424, n40425, n40426,
         n40427, n40428, n40429, n40430, n40431, n40432, n40433, n40434,
         n40435, n40436, n40437, n40438, n40439, n40440, n40441, n40442,
         n40443, n40444, n40445, n40446, n40447, n40448, n40449, n40450,
         n40451, n40452, n40453, n40454, n40455, n40456, n40457, n40458,
         n40459, n40460, n40461, n40462, n40463, n40464, n40465, n40466,
         n40467, n40468, n40469, n40470, n40471, n40472, n40473, n40474,
         n40475, n40476, n40477, n40478, n40479, n40480, n40481, n40482,
         n40483, n40484, n40485, n40486, n40487, n40488, n40489, n40490,
         n40491, n40492, n40493, n40494, n40495, n40496, n40497, n40498,
         n40499, n40500, n40501, n40502, n40503, n40504, n40505, n40506,
         n40507, n40508, n40509, n40510, n40511, n40512, n40513, n40514,
         n40515, n40516, n40517, n40518, n40519, n40520, n40521, n40522,
         n40523, n40524, n40525, n40526, n40527, n40528, n40529, n40530,
         n40531, n40532, n40533, n40534, n40535, n40536, n40537, n40538,
         n40539, n40540, n40541, n40542, n40543, n40544, n40545, n40546,
         n40547, n40548, n40549, n40550, n40551, n40552, n40553, n40554,
         n40555, n40556, n40557, n40558, n40559, n40560, n40561, n40562,
         n40563, n40564, n40565, n40566, n40567, n40568, n40569, n40570,
         n40571, n40572, n40573, n40574, n40575, n40576, n40577, n40578,
         n40579, n40580, n40581, n40582, n40583, n40584, n40585, n40586,
         n40587, n40588, n40589, n40590, n40591, n40592, n40593, n40594,
         n40595, n40596, n40597, n40598, n40599, n40600, n40601, n40602,
         n40603, n40604, n40605, n40606, n40607, n40608, n40609, n40610,
         n40611, n40612, n40613, n40614, n40615, n40616, n40617, n40618,
         n40619, n40620, n40621, n40622, n40623, n40624, n40625, n40626,
         n40627, n40628, n40629, n40630, n40631, n40632, n40633, n40634,
         n40635, n40636, n40637, n40638, n40639, n40640, n40641, n40642,
         n40643, n40644, n40645, n40646, n40647, n40648, n40649, n40650,
         n40651, n40652, n40653, n40654, n40655, n40656, n40657, n40658,
         n40659, n40660, n40661, n40662, n40663, n40664, n40665, n40666,
         n40667, n40668, n40669, n40670, n40671, n40672, n40673, n40674,
         n40675, n40676, n40677, n40678, n40679, n40680, n40681, n40682,
         n40683, n40684, n40685, n40686, n40687, n40688, n40689, n40690,
         n40691, n40692, n40693, n40694, n40695, n40696, n40697, n40698,
         n40699, n40700, n40701, n40702, n40703, n40704, n40705, n40706,
         n40707, n40708, n40709, n40710, n40711, n40712, n40713, n40714,
         n40715, n40716, n40717, n40718, n40719, n40720, n40721, n40722,
         n40723, n40724, n40725, n40726, n40727, n40728, n40729, n40730,
         n40731, n40732, n40733, n40734, n40735, n40736, n40737, n40738,
         n40739, n40740, n40741, n40742, n40743, n40744, n40745, n40746,
         n40747, n40748, n40749, n40750, n40751, n40752, n40753, n40754,
         n40755, n40756, n40757, n40758, n40759, n40760, n40761, n40762,
         n40763, n40764, n40765, n40766, n40767, n40768, n40769, n40770,
         n40771, n40772, n40773, n40774, n40775, n40776, n40777, n40778,
         n40779, n40780, n40781, n40782, n40783, n40784, n40785, n40786,
         n40787, n40788, n40789, n40790, n40791, n40792, n40793, n40794,
         n40795, n40796, n40797, n40798, n40799, n40800, n40801, n40802,
         n40803, n40804, n40805, n40806, n40807, n40808, n40809, n40810,
         n40811, n40812, n40813, n40814, n40815, n40816, n40817, n40818,
         n40819, n40820, n40821, n40822, n40823, n40824, n40825, n40826,
         n40827, n40828, n40829, n40830, n40831, n40832, n40833, n40834,
         n40835, n40836, n40837, n40838, n40839, n40840, n40841, n40842,
         n40843, n40844, n40845, n40846, n40847, n40848, n40849, n40850,
         n40851, n40852, n40853, n40854, n40855, n40856, n40857, n40858,
         n40859, n40860, n40861, n40862, n40863, n40864, n40865, n40866,
         n40867, n40868, n40869, n40870, n40871, n40872, n40873, n40874,
         n40875, n40876, n40877, n40878, n40879, n40880, n40881, n40882,
         n40883, n40884, n40885, n40886, n40887, n40888, n40889, n40890,
         n40891, n40892, n40893, n40894, n40895, n40896, n40897, n40898,
         n40899, n40900, n40901, n40902, n40903, n40904, n40905, n40906,
         n40907, n40908, n40909, n40910, n40911, n40912, n40913, n40914,
         n40915, n40916, n40917, n40918, n40919, n40920, n40921, n40922,
         n40923, n40924, n40925, n40926, n40927, n40928, n40929, n40930,
         n40931, n40932, n40933, n40934, n40935, n40936, n40937, n40938,
         n40939, n40940, n40941, n40942, n40943, n40944, n40945, n40946,
         n40947, n40948, n40949, n40950, n40951, n40952, n40953, n40954,
         n40955, n40956, n40957, n40958, n40959, n40960, n40961, n40962,
         n40963, n40964, n40965, n40966, n40967, n40968, n40969, n40970,
         n40971, n40972, n40973, n40974, n40975, n40976, n40977, n40978,
         n40979, n40980, n40981, n40982, n40983, n40984, n40985, n40986,
         n40987, n40988, n40989, n40990, n40991, n40992, n40993, n40994,
         n40995, n40996, n40997, n40998, n40999, n41000, n41001, n41002,
         n41003, n41004, n41005, n41006, n41007, n41008, n41009, n41010,
         n41011, n41012, n41013, n41014, n41015, n41016, n41017, n41018,
         n41019, n41020, n41021, n41022, n41023, n41024, n41025, n41026,
         n41027, n41028, n41029, n41030, n41031, n41032, n41033, n41034,
         n41035, n41036, n41037, n41038, n41039, n41040, n41041, n41042,
         n41043, n41044, n41045, n41046, n41047, n41048, n41049, n41050,
         n41051, n41052, n41053, n41054, n41055, n41056, n41057, n41058,
         n41059, n41060, n41061, n41062, n41063, n41064, n41065, n41066,
         n41067, n41068, n41069, n41070, n41071, n41072, n41073, n41074,
         n41075, n41076, n41077, n41078, n41079, n41080, n41081, n41082,
         n41083, n41084, n41085, n41086, n41087, n41088, n41089, n41090,
         n41091, n41092, n41093, n41094, n41095, n41096, n41097, n41098,
         n41099, n41100, n41101, n41102, n41103, n41104, n41105, n41106,
         n41107, n41108, n41109, n41110, n41111, n41112, n41113, n41114,
         n41115, n41116, n41117, n41118, n41119, n41120, n41121, n41122,
         n41123, n41124, n41125, n41126, n41127, n41128, n41129, n41130,
         n41131, n41132, n41133, n41134, n41135, n41136, n41137, n41138,
         n41139, n41140, n41141, n41142, n41143, n41144, n41145, n41146,
         n41147, n41148, n41149, n41150, n41151, n41152, n41153, n41154,
         n41155, n41156, n41157, n41158, n41159, n41160, n41161, n41162,
         n41163, n41164, n41165, n41166, n41167, n41168, n41169, n41170,
         n41171, n41172, n41173, n41174, n41175, n41176, n41177, n41178,
         n41179, n41180, n41181, n41182, n41183, n41184, n41185, n41186,
         n41187, n41188, n41189, n41190, n41191, n41192, n41193, n41194,
         n41195, n41196, n41197, n41198, n41199, n41200, n41201, n41202,
         n41203, n41204, n41205, n41206, n41207, n41208, n41209, n41210,
         n41211, n41212, n41213, n41214, n41215, n41216, n41217, n41218,
         n41219, n41220, n41221, n41222, n41223, n41224, n41225, n41226,
         n41227, n41228, n41229, n41230, n41231, n41232, n41233, n41234,
         n41235, n41236, n41237, n41238, n41239, n41240, n41241, n41242,
         n41243, n41244, n41245, n41246, n41247, n41248, n41249, n41250,
         n41251, n41252, n41253, n41254, n41255, n41256, n41257, n41258,
         n41259, n41260, n41261, n41262, n41263, n41264, n41265, n41266,
         n41267, n41268, n41269, n41270, n41271, n41272, n41273, n41274,
         n41275, n41276, n41277, n41278, n41279, n41280, n41281, n41282,
         n41283, n41284, n41285, n41286, n41287, n41288, n41289, n41290,
         n41291, n41292, n41293, n41294, n41295, n41296, n41297, n41298,
         n41299, n41300, n41301, n41302, n41303, n41304, n41305, n41306,
         n41307, n41308, n41309, n41310, n41311, n41312, n41313, n41314,
         n41315, n41316, n41317, n41318, n41319, n41320, n41321, n41322,
         n41323, n41324, n41325, n41326, n41327, n41328, n41329, n41330,
         n41331, n41332, n41333, n41334, n41335, n41336, n41337, n41338,
         n41339, n41340, n41341, n41342, n41343, n41344, n41345, n41346,
         n41347, n41348, n41349, n41350, n41351, n41352, n41353, n41354,
         n41355, n41356, n41357, n41358, n41359, n41360, n41361, n41362,
         n41363, n41364, n41365, n41366, n41367, n41368, n41369, n41370,
         n41371, n41372, n41373, n41374, n41375, n41376, n41377, n41378,
         n41379, n41380, n41381, n41382, n41383, n41384, n41385, n41386,
         n41387, n41388, n41389, n41390, n41391, n41392, n41393, n41394,
         n41395, n41396, n41397, n41398, n41399, n41400, n41401, n41402,
         n41403, n41404, n41405, n41406, n41407, n41408, n41409, n41410,
         n41411, n41412, n41413, n41414, n41415, n41416, n41417, n41418,
         n41419, n41420, n41421, n41422, n41423, n41424, n41425, n41426,
         n41427, n41428, n41429, n41430, n41431, n41432, n41433, n41434,
         n41435, n41436, n41437, n41438, n41439, n41440, n41441, n41442,
         n41443, n41444, n41445, n41446, n41447, n41448, n41449, n41450,
         n41451, n41452, n41453, n41454, n41455, n41456, n41457, n41458,
         n41459, n41460, n41461, n41462, n41463, n41464, n41465, n41466,
         n41467, n41468, n41469, n41470, n41471, n41472, n41473, n41474,
         n41475, n41476, n41477, n41478, n41479, n41480, n41481, n41482,
         n41483, n41484, n41485, n41486, n41487, n41488, n41489, n41490,
         n41491, n41492, n41493, n41494, n41495, n41496, n41497, n41498,
         n41499, n41500, n41501, n41502, n41503, n41504, n41505, n41506,
         n41507, n41508, n41509, n41510, n41511, n41512, n41513, n41514,
         n41515, n41516, n41517, n41518, n41519, n41520, n41521, n41522,
         n41523, n41524, n41525, n41526, n41527, n41528, n41529, n41530,
         n41531, n41532, n41533, n41534, n41535, n41536, n41537, n41538,
         n41539, n41540, n41541, n41542, n41543, n41544, n41545, n41546,
         n41547, n41548, n41549, n41550, n41551, n41552, n41553, n41554,
         n41555, n41556, n41557, n41558, n41559, n41560, n41561, n41562,
         n41563, n41564, n41565, n41566, n41567, n41568, n41569, n41570,
         n41571, n41572, n41573, n41574, n41575, n41576, n41577, n41578,
         n41579, n41580, n41581, n41582, n41583, n41584, n41585, n41586,
         n41587, n41588, n41589, n41590, n41591, n41592, n41593, n41594,
         n41595, n41596, n41597, n41598, n41599, n41600, n41601, n41602,
         n41603, n41604, n41605, n41606, n41607, n41608, n41609, n41610,
         n41611, n41612, n41613, n41614, n41615, n41616, n41617, n41618,
         n41619, n41620, n41621, n41622, n41623, n41624, n41625, n41626,
         n41627, n41628, n41629, n41630, n41631, n41632, n41633, n41634,
         n41635, n41636, n41637, n41638, n41639, n41640, n41641, n41642,
         n41643, n41644, n41645, n41646, n41647, n41648, n41649, n41650,
         n41651, n41652, n41653, n41654, n41655, n41656, n41657, n41658,
         n41659, n41660, n41661, n41662, n41663, n41664, n41665, n41666,
         n41667, n41668, n41669, n41670, n41671, n41672, n41673, n41674,
         n41675, n41676, n41677, n41678, n41679, n41680, n41681, n41682,
         n41683, n41684, n41685, n41686, n41687, n41688, n41689, n41690,
         n41691, n41692, n41693, n41694, n41695, n41696, n41697, n41698,
         n41699, n41700, n41701, n41702, n41703, n41704, n41705, n41706,
         n41707, n41708, n41709, n41710, n41711, n41712, n41713, n41714,
         n41715, n41716, n41717, n41718, n41719, n41720, n41721, n41722,
         n41723, n41724, n41725, n41726, n41727, n41728, n41729, n41730,
         n41731, n41732, n41733, n41734, n41735, n41736, n41737, n41738,
         n41739, n41740, n41741, n41742, n41743, n41744, n41745, n41746,
         n41747, n41748, n41749, n41750, n41751, n41752, n41753, n41754,
         n41755, n41756, n41757, n41758, n41759, n41760, n41761, n41762,
         n41763, n41764, n41765, n41766, n41767, n41768, n41769, n41770,
         n41771, n41772, n41773, n41774, n41775, n41776, n41777, n41778,
         n41779, n41780, n41781, n41782, n41783, n41784, n41785, n41786,
         n41787, n41788, n41789, n41790, n41791, n41792, n41793, n41794,
         n41795, n41796, n41797, n41798, n41799, n41800, n41801, n41802,
         n41803, n41804, n41805, n41806, n41807, n41808, n41809, n41810,
         n41811, n41812, n41813, n41814, n41815, n41816, n41817, n41818,
         n41819, n41820, n41821, n41822, n41823, n41824, n41825, n41826,
         n41827, n41828, n41829, n41830, n41831, n41832, n41833, n41834,
         n41835, n41836, n41837, n41838, n41839, n41840, n41841, n41842,
         n41843, n41844, n41845, n41846, n41847, n41848, n41849, n41850,
         n41851, n41852, n41853, n41854, n41855, n41856, n41857, n41858,
         n41859, n41860, n41861, n41862, n41863, n41864, n41865, n41866,
         n41867, n41868, n41869, n41870, n41871, n41872, n41873, n41874,
         n41875, n41876, n41877, n41878, n41879, n41880, n41881, n41882,
         n41883, n41884, n41885, n41886, n41887, n41888, n41889, n41890,
         n41891, n41892, n41893, n41894, n41895, n41896, n41897, n41898,
         n41899, n41900, n41901, n41902, n41903, n41904, n41905, n41906,
         n41907, n41908, n41909, n41910, n41911, n41912, n41913, n41914,
         n41915, n41916, n41917, n41918, n41919, n41920, n41921, n41922,
         n41923, n41924, n41925, n41926, n41927, n41928, n41929, n41930,
         n41931, n41932, n41933, n41934, n41935, n41936, n41937, n41938,
         n41939, n41940, n41941, n41942, n41943, n41944, n41945, n41946,
         n41947, n41948, n41949, n41950, n41951, n41952, n41953, n41954,
         n41955, n41956, n41957, n41958, n41959, n41960, n41961, n41962,
         n41963, n41964, n41965, n41966, n41967, n41968, n41969, n41970,
         n41971, n41972, n41973, n41974, n41975, n41976, n41977, n41978,
         n41979, n41980, n41981, n41982, n41983, n41984, n41985, n41986,
         n41987, n41988, n41989, n41990, n41991, n41992, n41993, n41994,
         n41995, n41996, n41997, n41998, n41999, n42000, n42001, n42002,
         n42003, n42004, n42005, n42006, n42007, n42008, n42009, n42010,
         n42011, n42012, n42013, n42014, n42015, n42016, n42017, n42018,
         n42019, n42020, n42021, n42022, n42023, n42024, n42025, n42026,
         n42027, n42028, n42029, n42030, n42031, n42032, n42033, n42034,
         n42035, n42036, n42037, n42038, n42039, n42040, n42041, n42042,
         n42043, n42044, n42045, n42046, n42047, n42048, n42049, n42050,
         n42051, n42052, n42053, n42054, n42055, n42056, n42057, n42058,
         n42059, n42060, n42061, n42062, n42063, n42064, n42065, n42066,
         n42067, n42068, n42069, n42070, n42071, n42072, n42073, n42074,
         n42075, n42076, n42077, n42078, n42079, n42080, n42081, n42082,
         n42083, n42084, n42085, n42086, n42087, n42088, n42089, n42090,
         n42091, n42092, n42093, n42094, n42095, n42096, n42097, n42098,
         n42099, n42100, n42101, n42102, n42103, n42104, n42105, n42106,
         n42107, n42108, n42109, n42110, n42111, n42112, n42113, n42114,
         n42115, n42116, n42117, n42118, n42119, n42120, n42121, n42122,
         n42123, n42124, n42125, n42126, n42127, n42128, n42129, n42130,
         n42131, n42132, n42133, n42134, n42135, n42136, n42137, n42138,
         n42139, n42140, n42141, n42142, n42143, n42144, n42145, n42146,
         n42147, n42148, n42149, n42150, n42151, n42152, n42153, n42154,
         n42155, n42156, n42157, n42158, n42159, n42160, n42161, n42162,
         n42163, n42164, n42165, n42166, n42167, n42168, n42169, n42170,
         n42171, n42172, n42173, n42174, n42175, n42176, n42177, n42178,
         n42179, n42180, n42181, n42182, n42183, n42184, n42185, n42186,
         n42187, n42188, n42189, n42190, n42191, n42192, n42193, n42194,
         n42195, n42196, n42197, n42198, n42199, n42200, n42201, n42202,
         n42203, n42204, n42205, n42206, n42207, n42208, n42209, n42210,
         n42211, n42212, n42213, n42214, n42215, n42216, n42217, n42218,
         n42219, n42220, n42221, n42222, n42223, n42224, n42225, n42226,
         n42227, n42228, n42229, n42230, n42231, n42232, n42233, n42234,
         n42235, n42236, n42237, n42238, n42239, n42240, n42241, n42242,
         n42243, n42244, n42245, n42246, n42247, n42248, n42249, n42250,
         n42251, n42252, n42253, n42254, n42255, n42256, n42257, n42258,
         n42259, n42260, n42261, n42262, n42263, n42264, n42265, n42266,
         n42267, n42268, n42269, n42270, n42271, n42272, n42273, n42274,
         n42275, n42276, n42277, n42278, n42279, n42280, n42281, n42282,
         n42283, n42284, n42285, n42286, n42287, n42288, n42289, n42290,
         n42291, n42292, n42293, n42294, n42295, n42296, n42297, n42298,
         n42299, n42300, n42301, n42302, n42303, n42304, n42305, n42306,
         n42307, n42308, n42309, n42310, n42311, n42312, n42313, n42314,
         n42315, n42316, n42317, n42318, n42319, n42320, n42321, n42322,
         n42323, n42324, n42325, n42326, n42327, n42328, n42329, n42330,
         n42331, n42332, n42333, n42334, n42335, n42336, n42337, n42338,
         n42339, n42340, n42341, n42342, n42343, n42344, n42345, n42346,
         n42347, n42348, n42349, n42350, n42351, n42352, n42353, n42354,
         n42355, n42356, n42357, n42358, n42359, n42360, n42361, n42362,
         n42363, n42364, n42365, n42366, n42367, n42368, n42369, n42370,
         n42371, n42372, n42373, n42374, n42375, n42376, n42377, n42378,
         n42379, n42380, n42381, n42382, n42383, n42384, n42385, n42386,
         n42387, n42388, n42389, n42390, n42391, n42392, n42393, n42394,
         n42395, n42396, n42397, n42398, n42399, n42400, n42401, n42402,
         n42403, n42404, n42405, n42406, n42407, n42408, n42409, n42410,
         n42411, n42412, n42413, n42414, n42415, n42416, n42417, n42418,
         n42419, n42420, n42421, n42422, n42423, n42424, n42425, n42426,
         n42427, n42428, n42429, n42430, n42431, n42432, n42433, n42434,
         n42435, n42436, n42437, n42438, n42439, n42440, n42441, n42442,
         n42443, n42444, n42445, n42446, n42447, n42448, n42449, n42450,
         n42451, n42452, n42453, n42454, n42455, n42456, n42457, n42458,
         n42459, n42460, n42461, n42462, n42463, n42464, n42465, n42466,
         n42467, n42468, n42469, n42470, n42471, n42472, n42473, n42474,
         n42475, n42476, n42477, n42478, n42479, n42480, n42481, n42482,
         n42483, n42484, n42485, n42486, n42487, n42488, n42489, n42490,
         n42491, n42492, n42493, n42494, n42495, n42496, n42497, n42498,
         n42499, n42500, n42501, n42502, n42503, n42504, n42505, n42506,
         n42507, n42508, n42509, n42510, n42511, n42512, n42513, n42514,
         n42515, n42516, n42517, n42518, n42519, n42520, n42521, n42522,
         n42523, n42524, n42525, n42526, n42527, n42528, n42529, n42530,
         n42531, n42532, n42533, n42534, n42535, n42536, n42537, n42538,
         n42539, n42540, n42541, n42542, n42543, n42544, n42545, n42546,
         n42547, n42548, n42549, n42550, n42551, n42552, n42553, n42554,
         n42555, n42556, n42557, n42558, n42559, n42560, n42561, n42562,
         n42563, n42564, n42565, n42566, n42567, n42568, n42569, n42570,
         n42571, n42572, n42573, n42574, n42575, n42576, n42577, n42578,
         n42579, n42580, n42581, n42582, n42583, n42584, n42585, n42586,
         n42587, n42588, n42589, n42590, n42591, n42592, n42593, n42594,
         n42595, n42596, n42597, n42598, n42599, n42600, n42601, n42602,
         n42603, n42604, n42605, n42606, n42607, n42608, n42609, n42610,
         n42611, n42612, n42613, n42614, n42615, n42616, n42617, n42618,
         n42619, n42620, n42621, n42622, n42623, n42624, n42625, n42626,
         n42627, n42628, n42629, n42630, n42631, n42632, n42633, n42634,
         n42635, n42636, n42637, n42638, n42639, n42640, n42641, n42642,
         n42643, n42644, n42645, n42646, n42647, n42648, n42649, n42650,
         n42651, n42652, n42653, n42654, n42655, n42656, n42657, n42658,
         n42659, n42660, n42661, n42662, n42663, n42664, n42665, n42666,
         n42667, n42668, n42669, n42670, n42671, n42672, n42673, n42674,
         n42675, n42676, n42677, n42678, n42679, n42680, n42681, n42682,
         n42683, n42684, n42685, n42686, n42687, n42688, n42689, n42690,
         n42691, n42692, n42693, n42694, n42695, n42696, n42697, n42698,
         n42699, n42700, n42701, n42702, n42703, n42704, n42705, n42706,
         n42707, n42708, n42709, n42710, n42711, n42712, n42713, n42714,
         n42715, n42716, n42717, n42718, n42719, n42720, n42721, n42722,
         n42723, n42724, n42725, n42726, n42727, n42728, n42729, n42730,
         n42731, n42732, n42733, n42734, n42735, n42736, n42737, n42738,
         n42739, n42740, n42741, n42742, n42743, n42744, n42745, n42746,
         n42747, n42748, n42749, n42750, n42751, n42752, n42753, n42754,
         n42755, n42756, n42757, n42758, n42759, n42760, n42761, n42762,
         n42763, n42764, n42765, n42766, n42767, n42768, n42769, n42770,
         n42771, n42772, n42773, n42774, n42775, n42776, n42777, n42778,
         n42779, n42780, n42781, n42782, n42783, n42784, n42785, n42786,
         n42787, n42788, n42789, n42790, n42791, n42792, n42793, n42794,
         n42795, n42796, n42797, n42798, n42799, n42800, n42801, n42802,
         n42803, n42804, n42805, n42806, n42807, n42808, n42809, n42810,
         n42811, n42812, n42813, n42814, n42815, n42816, n42817, n42818,
         n42819, n42820, n42821, n42822, n42823, n42824, n42825, n42826,
         n42827, n42828, n42829, n42830, n42831, n42832, n42833, n42834,
         n42835, n42836, n42837, n42838, n42839, n42840, n42841, n42842,
         n42843, n42844, n42845, n42846, n42847, n42848, n42849, n42850,
         n42851, n42852, n42853, n42854, n42855, n42856, n42857, n42858,
         n42859, n42860, n42861, n42862, n42863, n42864, n42865, n42866,
         n42867, n42868, n42869, n42870, n42871, n42872, n42873, n42874,
         n42875, n42876, n42877, n42878, n42879, n42880, n42881, n42882,
         n42883, n42884, n42885, n42886, n42887, n42888, n42889, n42890,
         n42891, n42892, n42893, n42894, n42895, n42896, n42897, n42898,
         n42899, n42900, n42901, n42902, n42903, n42904, n42905, n42906,
         n42907, n42908, n42909, n42910, n42911, n42912, n42913, n42914,
         n42915, n42916, n42917, n42918, n42919, n42920, n42921, n42922,
         n42923, n42924, n42925, n42926, n42927, n42928, n42929, n42930,
         n42931, n42932, n42933, n42934, n42935, n42936, n42937, n42938,
         n42939, n42940, n42941, n42942, n42943, n42944, n42945, n42946,
         n42947, n42948, n42949, n42950, n42951, n42952, n42953, n42954,
         n42955, n42956, n42957, n42958, n42959, n42960, n42961, n42962,
         n42963, n42964, n42965, n42966, n42967, n42968, n42969, n42970,
         n42971, n42972, n42973, n42974, n42975, n42976, n42977, n42978,
         n42979, n42980, n42981, n42982, n42983, n42984, n42985, n42986,
         n42987, n42988, n42989, n42990, n42991, n42992, n42993, n42994,
         n42995, n42996, n42997, n42998, n42999, n43000, n43001, n43002,
         n43003, n43004, n43005, n43006, n43007, n43008, n43009, n43010,
         n43011, n43012, n43013, n43014, n43015, n43016, n43017, n43018,
         n43019, n43020, n43021, n43022, n43023, n43024, n43025, n43026,
         n43027, n43028, n43029, n43030, n43031, n43032, n43033, n43034,
         n43035, n43036, n43037, n43038, n43039, n43040, n43041, n43042,
         n43043, n43044, n43045, n43046, n43047, n43048, n43049, n43050,
         n43051, n43052, n43053, n43054, n43055, n43056, n43057, n43058,
         n43059, n43060, n43061, n43062, n43063, n43064, n43065, n43066,
         n43067, n43068, n43069, n43070, n43071, n43072, n43073, n43074,
         n43075, n43076, n43077, n43078, n43079, n43080, n43081, n43082,
         n43083, n43084, n43085, n43086, n43087, n43088, n43089, n43090,
         n43091, n43092, n43093, n43094, n43095, n43096, n43097, n43098,
         n43099, n43100, n43101, n43102, n43103, n43104, n43105, n43106,
         n43107, n43108, n43109, n43110, n43111, n43112, n43113, n43114,
         n43115, n43116, n43117, n43118, n43119, n43120, n43121, n43122,
         n43123, n43124, n43125, n43126, n43127, n43128, n43129, n43130,
         n43131, n43132, n43133, n43134, n43135, n43136, n43137, n43138,
         n43139, n43140, n43141, n43142, n43143, n43144, n43145, n43146,
         n43147, n43148, n43149, n43150, n43151, n43152, n43153, n43154,
         n43155, n43156, n43157, n43158, n43159, n43160, n43161, n43162,
         n43163, n43164, n43165, n43166, n43167, n43168, n43169, n43170,
         n43171, n43172, n43173, n43174, n43175, n43176, n43177, n43178,
         n43179, n43180, n43181, n43182, n43183, n43184, n43185, n43186,
         n43187, n43188, n43189, n43190, n43191, n43192, n43193, n43194,
         n43195, n43196, n43197, n43198, n43199, n43200, n43201, n43202,
         n43203, n43204, n43205, n43206, n43207, n43208, n43209, n43210,
         n43211, n43212, n43213, n43214, n43215, n43216, n43217, n43218,
         n43219, n43220, n43221, n43222, n43223, n43224, n43225, n43226,
         n43227, n43228, n43229, n43230, n43231, n43232, n43233, n43234,
         n43235, n43236, n43237, n43238, n43239, n43240, n43241, n43242,
         n43243, n43244, n43245, n43246, n43247, n43248, n43249, n43250,
         n43251, n43252, n43253, n43254, n43255, n43256, n43257, n43258,
         n43259, n43260, n43261, n43262, n43263, n43264, n43265, n43266,
         n43267, n43268, n43269, n43270, n43271, n43272, n43273, n43274,
         n43275, n43276, n43277, n43278, n43279, n43280, n43281, n43282,
         n43283, n43284, n43285, n43286, n43287, n43288, n43289, n43290,
         n43291, n43292, n43293, n43294, n43295, n43296, n43297, n43298,
         n43299, n43300, n43301, n43302, n43303, n43304, n43305, n43306,
         n43307, n43308, n43309, n43310, n43311, n43312, n43313, n43314,
         n43315, n43316, n43317, n43318, n43319, n43320, n43321, n43322,
         n43323, n43324, n43325, n43326, n43327, n43328, n43329, n43330,
         n43331, n43332, n43333, n43334, n43335, n43336, n43337, n43338,
         n43339, n43340, n43341, n43342, n43343, n43344, n43345, n43346,
         n43347, n43348, n43349, n43350, n43351, n43352, n43353, n43354,
         n43355, n43356, n43357, n43358, n43359, n43360, n43361, n43362,
         n43363, n43364, n43365, n43366, n43367, n43368, n43369, n43370,
         n43371, n43372, n43373, n43374, n43375, n43376, n43377, n43378,
         n43379, n43380, n43381, n43382, n43383, n43384, n43385, n43386,
         n43387, n43388, n43389, n43390, n43391, n43392, n43393, n43394,
         n43395, n43396, n43397, n43398, n43399, n43400, n43401, n43402,
         n43403, n43404, n43405, n43406, n43407, n43408, n43409, n43410,
         n43411, n43412, n43413, n43414, n43415, n43416, n43417, n43418,
         n43419, n43420, n43421, n43422, n43423, n43424, n43425, n43426,
         n43427, n43428, n43429, n43430, n43431, n43432, n43433, n43434,
         n43435, n43436, n43437, n43438, n43439, n43440, n43441, n43442,
         n43443, n43444, n43445, n43446, n43447, n43448, n43449, n43450,
         n43451, n43452, n43453, n43454, n43455, n43456, n43457, n43458,
         n43459, n43460, n43461, n43462, n43463, n43464, n43465, n43466,
         n43467, n43468, n43469, n43470, n43471, n43472, n43473, n43474,
         n43475, n43476, n43477, n43478, n43479, n43480, n43481, n43482,
         n43483, n43484, n43485, n43486, n43487, n43488, n43489, n43490,
         n43491, n43492, n43493, n43494, n43495, n43496, n43497, n43498,
         n43499, n43500, n43501, n43502, n43503, n43504, n43505, n43506,
         n43507, n43508, n43509, n43510, n43511, n43512, n43513, n43514,
         n43515, n43516, n43517, n43518, n43519, n43520, n43521, n43522,
         n43523, n43524, n43525, n43526, n43527, n43528, n43529, n43530,
         n43531, n43532, n43533, n43534, n43535, n43536, n43537, n43538,
         n43539, n43540, n43541, n43542, n43543, n43544, n43545, n43546,
         n43547, n43548, n43549, n43550, n43551, n43552, n43553, n43554,
         n43555, n43556, n43557, n43558, n43559, n43560, n43561, n43562,
         n43563, n43564, n43565, n43566, n43567, n43568, n43569, n43570,
         n43571, n43572, n43573, n43574, n43575, n43576, n43577, n43578,
         n43579, n43580, n43581, n43582, n43583, n43584, n43585, n43586,
         n43587, n43588, n43589, n43590, n43591, n43592, n43593, n43594,
         n43595, n43596, n43597, n43598, n43599, n43600, n43601, n43602,
         n43603, n43604, n43605, n43606, n43607, n43608, n43609, n43610,
         n43611, n43612, n43613, n43614, n43615, n43616, n43617, n43618,
         n43619, n43620, n43621, n43622, n43623, n43624, n43625, n43626,
         n43627, n43628, n43629, n43630, n43631, n43632, n43633, n43634,
         n43635, n43636, n43637, n43638, n43639, n43640, n43641, n43642,
         n43643, n43644, n43645, n43646, n43647, n43648, n43649, n43650,
         n43651, n43652, n43653, n43654, n43655, n43656, n43657, n43658,
         n43659, n43660, n43661, n43662, n43663, n43664, n43665, n43666,
         n43667, n43668, n43669, n43670, n43671, n43672, n43673, n43674,
         n43675, n43676, n43677, n43678, n43679, n43680, n43681, n43682,
         n43683, n43684, n43685, n43686, n43687, n43688, n43689, n43690,
         n43691, n43692, n43693, n43694, n43695, n43696, n43697, n43698,
         n43699, n43700, n43701, n43702, n43703, n43704, n43705, n43706,
         n43707, n43708, n43709, n43710, n43711, n43712, n43713, n43714,
         n43715, n43716, n43717, n43718, n43719, n43720, n43721, n43722,
         n43723, n43724, n43725, n43726, n43727, n43728, n43729, n43730,
         n43731, n43732, n43733, n43734, n43735, n43736, n43737, n43738,
         n43739, n43740, n43741, n43742, n43743, n43744, n43745, n43746,
         n43747, n43748, n43749, n43750, n43751, n43752, n43753, n43754,
         n43755, n43756, n43757, n43758, n43759, n43760, n43761, n43762,
         n43763, n43764, n43765, n43766, n43767, n43768, n43769, n43770,
         n43771, n43772, n43773, n43774, n43775, n43776, n43777, n43778,
         n43779, n43780, n43781, n43782, n43783, n43784, n43785, n43786,
         n43787, n43788, n43789, n43790, n43791, n43792, n43793, n43794,
         n43795, n43796, n43797, n43798, n43799, n43800, n43801, n43802,
         n43803, n43804, n43805, n43806, n43807, n43808, n43809, n43810,
         n43811, n43812, n43813, n43814, n43815, n43816, n43817, n43818,
         n43819, n43820, n43821, n43822, n43823, n43824, n43825, n43826,
         n43827, n43828, n43829, n43830, n43831, n43832, n43833, n43834,
         n43835, n43836, n43837, n43838, n43839, n43840, n43841, n43842,
         n43843, n43844, n43845, n43846, n43847, n43848, n43849, n43850,
         n43851, n43852, n43853, n43854, n43855, n43856, n43857, n43858,
         n43859, n43860, n43861, n43862, n43863, n43864, n43865, n43866,
         n43867, n43868, n43869, n43870, n43871, n43872, n43873, n43874,
         n43875, n43876, n43877, n43878, n43879, n43880, n43881, n43882,
         n43883, n43884, n43885, n43886, n43887, n43888, n43889, n43890,
         n43891, n43892, n43893, n43894, n43895, n43896, n43897, n43898,
         n43899, n43900, n43901, n43902, n43903, n43904, n43905, n43906,
         n43907, n43908, n43909, n43910, n43911, n43912, n43913, n43914,
         n43915, n43916, n43917, n43918, n43919, n43920, n43921, n43922,
         n43923, n43924, n43925, n43926, n43927, n43928, n43929, n43930,
         n43931, n43932, n43933, n43934, n43935, n43936, n43937, n43938,
         n43939, n43940, n43941, n43942, n43943, n43944, n43945, n43946,
         n43947, n43948, n43949, n43950, n43951, n43952, n43953, n43954,
         n43955, n43956, n43957, n43958, n43959, n43960, n43961, n43962,
         n43963, n43964, n43965, n43966, n43967, n43968, n43969, n43970,
         n43971, n43972, n43973, n43974, n43975, n43976, n43977, n43978,
         n43979, n43980, n43981, n43982, n43983, n43984, n43985, n43986,
         n43987, n43988, n43989, n43990, n43991, n43992, n43993, n43994,
         n43995, n43996, n43997, n43998, n43999, n44000, n44001, n44002,
         n44003, n44004, n44005, n44006, n44007, n44008, n44009, n44010,
         n44011, n44012, n44013, n44014, n44015, n44016, n44017, n44018,
         n44019, n44020, n44021, n44022, n44023, n44024, n44025, n44026,
         n44027, n44028, n44029, n44030, n44031, n44032, n44033, n44034,
         n44035, n44036, n44037, n44038, n44039, n44040, n44041, n44042,
         n44043, n44044, n44045, n44046, n44047, n44048, n44049, n44050,
         n44051, n44052, n44053, n44054, n44055, n44056, n44057, n44058,
         n44059, n44060, n44061, n44062, n44063, n44064, n44065, n44066,
         n44067, n44068, n44069, n44070, n44071, n44072, n44073, n44074,
         n44075, n44076, n44077, n44078, n44079, n44080, n44081, n44082,
         n44083, n44084, n44085, n44086, n44087, n44088, n44089, n44090,
         n44091, n44092, n44093, n44094, n44095, n44096, n44097, n44098,
         n44099, n44100, n44101, n44102, n44103, n44104, n44105, n44106,
         n44107, n44108, n44109, n44110, n44111, n44112, n44113, n44114,
         n44115, n44116, n44117, n44118, n44119, n44120, n44121, n44122,
         n44123, n44124, n44125, n44126, n44127, n44128, n44129, n44130,
         n44131, n44132, n44133, n44134, n44135, n44136, n44137, n44138,
         n44139, n44140, n44141, n44142, n44143, n44144, n44145, n44146,
         n44147, n44148, n44149, n44150, n44151, n44152, n44153, n44154,
         n44155, n44156, n44157, n44158, n44159, n44160, n44161, n44162,
         n44163, n44164, n44165, n44166, n44167, n44168, n44169, n44170,
         n44171, n44172, n44173, n44174, n44175, n44176, n44177, n44178,
         n44179, n44180, n44181, n44182, n44183, n44184, n44185, n44186,
         n44187, n44188, n44189, n44190, n44191, n44192, n44193, n44194,
         n44195, n44196, n44197, n44198, n44199, n44200, n44201, n44202,
         n44203, n44204, n44205, n44206, n44207, n44208, n44209, n44210,
         n44211, n44212, n44213, n44214, n44215, n44216, n44217, n44218,
         n44219, n44220, n44221, n44222, n44223, n44224, n44225, n44226,
         n44227, n44228, n44229, n44230, n44231, n44232, n44233, n44234,
         n44235, n44236, n44237, n44238, n44239, n44240, n44241, n44242,
         n44243, n44244, n44245, n44246, n44247, n44248, n44249, n44250,
         n44251, n44252, n44253, n44254, n44255, n44256, n44257, n44258,
         n44259, n44260, n44261, n44262, n44263, n44264, n44265, n44266,
         n44267, n44268, n44269, n44270, n44271, n44272, n44273, n44274,
         n44275, n44276, n44277, n44278, n44279, n44280, n44281, n44282,
         n44283, n44284, n44285, n44286, n44287, n44288, n44289, n44290,
         n44291, n44292, n44293, n44294, n44295, n44296, n44297, n44298,
         n44299, n44300, n44301, n44302, n44303, n44304, n44305, n44306,
         n44307, n44308, n44309, n44310, n44311, n44312, n44313, n44314,
         n44315, n44316, n44317, n44318, n44319, n44320, n44321, n44322,
         n44323, n44324, n44325, n44326, n44327, n44328, n44329, n44330,
         n44331, n44332, n44333, n44334, n44335, n44336, n44337, n44338,
         n44339, n44340, n44341, n44342, n44343, n44344, n44345, n44346,
         n44347, n44348, n44349, n44350, n44351, n44352, n44353, n44354,
         n44355, n44356, n44357, n44358, n44359, n44360, n44361, n44362,
         n44363, n44364, n44365, n44366, n44367, n44368, n44369, n44370,
         n44371, n44372, n44373, n44374, n44375, n44376, n44377, n44378,
         n44379, n44380, n44381, n44382, n44383, n44384, n44385, n44386,
         n44387, n44388, n44389, n44390, n44391, n44392, n44393, n44394,
         n44395, n44396, n44397, n44398, n44399, n44400, n44401, n44402,
         n44403, n44404, n44405, n44406, n44407, n44408, n44409, n44410,
         n44411, n44412, n44413, n44414, n44415, n44416, n44417, n44418,
         n44419, n44420, n44421, n44422, n44423, n44424, n44425, n44426,
         n44427, n44428, n44429, n44430, n44431, n44432, n44433, n44434,
         n44435, n44436, n44437, n44438, n44439, n44440, n44441, n44442,
         n44443, n44444, n44445, n44446, n44447, n44448, n44449, n44450,
         n44451, n44452, n44453, n44454, n44455, n44456, n44457, n44458,
         n44459, n44460, n44461, n44462, n44463, n44464, n44465, n44466,
         n44467, n44468, n44469, n44470, n44471, n44472, n44473, n44474,
         n44475, n44476, n44477, n44478, n44479, n44480, n44481, n44482,
         n44483, n44484, n44485, n44486, n44487, n44488, n44489, n44490,
         n44491, n44492, n44493, n44494, n44495, n44496, n44497, n44498,
         n44499, n44500, n44501, n44502, n44503, n44504, n44505, n44506,
         n44507, n44508, n44509, n44510, n44511, n44512, n44513, n44514,
         n44515, n44516, n44517, n44518, n44519, n44520, n44521, n44522,
         n44523, n44524, n44525, n44526, n44527, n44528, n44529, n44530,
         n44531, n44532, n44533, n44534, n44535, n44536, n44537, n44538,
         n44539, n44540, n44541, n44542, n44543, n44544, n44545, n44546,
         n44547, n44548, n44549, n44550, n44551, n44552, n44553, n44554,
         n44555, n44556, n44557, n44558, n44559, n44560, n44561, n44562,
         n44563, n44564, n44565, n44566, n44567, n44568, n44569, n44570,
         n44571, n44572, n44573, n44574, n44575, n44576, n44577, n44578,
         n44579, n44580, n44581, n44582, n44583, n44584, n44585, n44586,
         n44587, n44588, n44589, n44590, n44591, n44592, n44593, n44594,
         n44595, n44596, n44597, n44598, n44599, n44600, n44601, n44602,
         n44603, n44604, n44605, n44606, n44607, n44608, n44609, n44610,
         n44611, n44612, n44613, n44614, n44615, n44616, n44617, n44618,
         n44619, n44620, n44621, n44622, n44623, n44624, n44625, n44626,
         n44627, n44628, n44629, n44630, n44631, n44632, n44633, n44634,
         n44635, n44636, n44637, n44638, n44639, n44640, n44641, n44642,
         n44643, n44644, n44645, n44646, n44647, n44648, n44649, n44650,
         n44651, n44652, n44653, n44654, n44655, n44656, n44657, n44658,
         n44659, n44660, n44661, n44662, n44663, n44664, n44665, n44666,
         n44667, n44668, n44669, n44670, n44671, n44672, n44673, n44674,
         n44675, n44676, n44677, n44678, n44679, n44680, n44681, n44682,
         n44683, n44684, n44685, n44686, n44687, n44688, n44689, n44690,
         n44691, n44692, n44693, n44694, n44695, n44696, n44697, n44698,
         n44699, n44700, n44701, n44702, n44703, n44704, n44705, n44706,
         n44707, n44708, n44709, n44710, n44711, n44712, n44713, n44714,
         n44715, n44716, n44717, n44718, n44719, n44720, n44721, n44722,
         n44723, n44724, n44725, n44726, n44727, n44728, n44729, n44730,
         n44731, n44732, n44733, n44734, n44735, n44736, n44737, n44738,
         n44739, n44740, n44741, n44742, n44743, n44744, n44745, n44746,
         n44747, n44748, n44749, n44750, n44751, n44752, n44753, n44754,
         n44755, n44756, n44757, n44758, n44759, n44760, n44761, n44762,
         n44763, n44764, n44765, n44766, n44767, n44768, n44769, n44770,
         n44771, n44772, n44773, n44774, n44775, n44776, n44777, n44778,
         n44779, n44780, n44781, n44782, n44783, n44784, n44785, n44786,
         n44787, n44788, n44789, n44790, n44791, n44792, n44793, n44794,
         n44795, n44796, n44797, n44798, n44799, n44800, n44801, n44802,
         n44803, n44804, n44805, n44806, n44807, n44808, n44809, n44810,
         n44811, n44812, n44813, n44814, n44815, n44816, n44817, n44818,
         n44819, n44820, n44821, n44822, n44823, n44824, n44825, n44826,
         n44827, n44828, n44829, n44830, n44831, n44832, n44833, n44834,
         n44835, n44836, n44837, n44838, n44839, n44840, n44841, n44842,
         n44843, n44844, n44845, n44846, n44847, n44848, n44849, n44850,
         n44851, n44852, n44853, n44854, n44855, n44856, n44857, n44858,
         n44859, n44860, n44861, n44862, n44863, n44864, n44865, n44866,
         n44867, n44868, n44869, n44870, n44871, n44872, n44873, n44874,
         n44875, n44876, n44877, n44878, n44879, n44880, n44881, n44882,
         n44883, n44884, n44885, n44886, n44887, n44888, n44889, n44890,
         n44891, n44892, n44893, n44894, n44895, n44896, n44897, n44898,
         n44899, n44900, n44901, n44902, n44903, n44904, n44905, n44906,
         n44907, n44908, n44909, n44910, n44911, n44912, n44913, n44914,
         n44915, n44916, n44917, n44918, n44919, n44920, n44921, n44922,
         n44923, n44924, n44925, n44926, n44927, n44928, n44929, n44930,
         n44931, n44932, n44933, n44934, n44935, n44936, n44937, n44938,
         n44939, n44940, n44941, n44942, n44943, n44944, n44945, n44946,
         n44947, n44948, n44949, n44950, n44951, n44952, n44953, n44954,
         n44955, n44956, n44957, n44958, n44959, n44960, n44961, n44962,
         n44963, n44964, n44965, n44966, n44967, n44968, n44969, n44970,
         n44971, n44972, n44973, n44974, n44975, n44976, n44977, n44978,
         n44979, n44980, n44981, n44982, n44983, n44984, n44985, n44986,
         n44987, n44988, n44989, n44990, n44991, n44992, n44993, n44994,
         n44995, n44996, n44997, n44998, n44999, n45000, n45001, n45002,
         n45003, n45004, n45005, n45006, n45007, n45008, n45009, n45010,
         n45011, n45012, n45013, n45014, n45015, n45016, n45017, n45018,
         n45019, n45020, n45021, n45022, n45023, n45024, n45025, n45026,
         n45027, n45028, n45029, n45030, n45031, n45032, n45033, n45034,
         n45035, n45036, n45037, n45038, n45039, n45040, n45041, n45042,
         n45043, n45044, n45045, n45046, n45047, n45048, n45049, n45050,
         n45051, n45052, n45053, n45054, n45055, n45056, n45057, n45058,
         n45059, n45060, n45061, n45062, n45063, n45064, n45065, n45066,
         n45067, n45068, n45069, n45070, n45071, n45072, n45073, n45074,
         n45075, n45076, n45077, n45078, n45079, n45080, n45081, n45082,
         n45083, n45084, n45085, n45086, n45087, n45088, n45089, n45090,
         n45091, n45092, n45093, n45094, n45095, n45096, n45097, n45098,
         n45099, n45100, n45101, n45102, n45103, n45104, n45105, n45106,
         n45107, n45108, n45109, n45110, n45111, n45112, n45113, n45114,
         n45115, n45116, n45117, n45118, n45119, n45120, n45121, n45122,
         n45123, n45124, n45125, n45126, n45127, n45128, n45129, n45130,
         n45131, n45132, n45133, n45134, n45135, n45136, n45137, n45138,
         n45139, n45140, n45141, n45142, n45143, n45144, n45145, n45146,
         n45147, n45148, n45149, n45150, n45151, n45152, n45153, n45154,
         n45155, n45156, n45157, n45158, n45159, n45160, n45161, n45162,
         n45163, n45164, n45165, n45166, n45167, n45168, n45169, n45170,
         n45171, n45172, n45173, n45174, n45175, n45176, n45177, n45178,
         n45179, n45180, n45181, n45182, n45183, n45184, n45185, n45186,
         n45187, n45188, n45189, n45190, n45191, n45192, n45193, n45194,
         n45195, n45196, n45197, n45198, n45199, n45200, n45201, n45202,
         n45203, n45204, n45205, n45206, n45207, n45208, n45209, n45210,
         n45211, n45212, n45213, n45214, n45215, n45216, n45217, n45218,
         n45219, n45220, n45221, n45222, n45223, n45224, n45225, n45226,
         n45227, n45228, n45229, n45230, n45231, n45232, n45233, n45234,
         n45235, n45236, n45237, n45238, n45239, n45240, n45241, n45242,
         n45243, n45244, n45245, n45246, n45247, n45248, n45249, n45250,
         n45251, n45252, n45253, n45254, n45255, n45256, n45257, n45258,
         n45259, n45260, n45261, n45262, n45263, n45264, n45265, n45266,
         n45267, n45268, n45269, n45270, n45271, n45272, n45273, n45274,
         n45275, n45276, n45277, n45278, n45279, n45280, n45281, n45282,
         n45283, n45284, n45285, n45286, n45287, n45288, n45289, n45290,
         n45291, n45292, n45293, n45294, n45295, n45296, n45297, n45298,
         n45299, n45300, n45301, n45302, n45303, n45304, n45305, n45306,
         n45307, n45308, n45309, n45310, n45311, n45312, n45313, n45314,
         n45315, n45316, n45317, n45318, n45319, n45320, n45321, n45322,
         n45323, n45324, n45325, n45326, n45327, n45328, n45329, n45330,
         n45331, n45332, n45333, n45334, n45335, n45336, n45337, n45338,
         n45339, n45340, n45341, n45342, n45343, n45344, n45345, n45346,
         n45347, n45348, n45349, n45350, n45351, n45352, n45353, n45354,
         n45355, n45356, n45357, n45358, n45359, n45360, n45361, n45362,
         n45363, n45364, n45365, n45366, n45367, n45368, n45369, n45370,
         n45371, n45372, n45373, n45374, n45375, n45376, n45377, n45378,
         n45379, n45380, n45381, n45382, n45383, n45384, n45385, n45386,
         n45387, n45388, n45389, n45390, n45391, n45392, n45393, n45394,
         n45395, n45396, n45397, n45398, n45399, n45400, n45401, n45402,
         n45403, n45404, n45405, n45406, n45407, n45408, n45409, n45410,
         n45411, n45412, n45413, n45414, n45415, n45416, n45417, n45418,
         n45419, n45420, n45421, n45422, n45423, n45424, n45425, n45426,
         n45427, n45428, n45429, n45430, n45431, n45432, n45433, n45434,
         n45435, n45436, n45437, n45438, n45439, n45440, n45441, n45442,
         n45443, n45444, n45445, n45446, n45447, n45448, n45449, n45450,
         n45451, n45452, n45453, n45454, n45455, n45456, n45457, n45458,
         n45459, n45460, n45461, n45462, n45463, n45464, n45465, n45466,
         n45467, n45468, n45469, n45470, n45471, n45472, n45473, n45474,
         n45475, n45476, n45477, n45478, n45479, n45480, n45481, n45482,
         n45483, n45484, n45485, n45486, n45487, n45488, n45489, n45490,
         n45491, n45492, n45493, n45494, n45495, n45496, n45497, n45498,
         n45499, n45500, n45501, n45502, n45503, n45504, n45505, n45506,
         n45507, n45508, n45509, n45510, n45511, n45512, n45513, n45514,
         n45515, n45516, n45517, n45518, n45519, n45520, n45521, n45522,
         n45523, n45524, n45525, n45526, n45527, n45528, n45529, n45530,
         n45531, n45532, n45533, n45534, n45535, n45536, n45537, n45538,
         n45539, n45540, n45541, n45542, n45543, n45544, n45545, n45546,
         n45547, n45548, n45549, n45550, n45551, n45552, n45553, n45554,
         n45555, n45556, n45557, n45558, n45559, n45560, n45561, n45562,
         n45563, n45564, n45565, n45566, n45567, n45568, n45569, n45570,
         n45571, n45572, n45573, n45574, n45575, n45576, n45577, n45578,
         n45579, n45580, n45581, n45582, n45583, n45584, n45585, n45586,
         n45587, n45588, n45589, n45590, n45591, n45592, n45593, n45594,
         n45595, n45596, n45597, n45598, n45599, n45600, n45601, n45602,
         n45603, n45604, n45605, n45606, n45607, n45608, n45609, n45610,
         n45611, n45612, n45613, n45614, n45615, n45616, n45617, n45618,
         n45619, n45620, n45621, n45622, n45623, n45624, n45625, n45626,
         n45627, n45628, n45629, n45630, n45631, n45632, n45633, n45634,
         n45635, n45636, n45637, n45638, n45639, n45640, n45641, n45642,
         n45643, n45644, n45645, n45646, n45647, n45648, n45649, n45650,
         n45651, n45652, n45653, n45654, n45655, n45656, n45657, n45658,
         n45659, n45660, n45661, n45662, n45663, n45664, n45665, n45666,
         n45667, n45668, n45669, n45670, n45671, n45672, n45673, n45674,
         n45675, n45676, n45677, n45678, n45679, n45680, n45681, n45682,
         n45683, n45684, n45685, n45686, n45687, n45688, n45689, n45690,
         n45691, n45692, n45693, n45694, n45695, n45696, n45697, n45698,
         n45699, n45700, n45701, n45702, n45703, n45704, n45705, n45706,
         n45707, n45708, n45709, n45710, n45711, n45712, n45713, n45714,
         n45715, n45716, n45717, n45718, n45719, n45720, n45721, n45722,
         n45723, n45724, n45725, n45726, n45727, n45728, n45729, n45730,
         n45731, n45732, n45733, n45734, n45735, n45736, n45737, n45738,
         n45739, n45740, n45741, n45742, n45743, n45744, n45745, n45746,
         n45747, n45748, n45749, n45750, n45751, n45752, n45753, n45754,
         n45755, n45756, n45757, n45758, n45759, n45760, n45761, n45762,
         n45763, n45764, n45765, n45766, n45767, n45768, n45769, n45770,
         n45771, n45772, n45773, n45774, n45775, n45776, n45777, n45778,
         n45779, n45780, n45781, n45782, n45783, n45784, n45785, n45786,
         n45787, n45788, n45789, n45790, n45791, n45792, n45793, n45794,
         n45795, n45796, n45797, n45798, n45799, n45800, n45801, n45802,
         n45803, n45804, n45805, n45806, n45807, n45808, n45809, n45810,
         n45811, n45812, n45813, n45814, n45815, n45816, n45817, n45818,
         n45819, n45820, n45821, n45822, n45823, n45824, n45825, n45826,
         n45827, n45828, n45829, n45830, n45831, n45832, n45833, n45834,
         n45835, n45836, n45837, n45838, n45839, n45840, n45841, n45842,
         n45843, n45844, n45845, n45846, n45847, n45848, n45849, n45850,
         n45851, n45852, n45853, n45854, n45855, n45856, n45857, n45858,
         n45859, n45860, n45861, n45862, n45863, n45864, n45865, n45866,
         n45867, n45868, n45869, n45870, n45871, n45872, n45873, n45874,
         n45875, n45876, n45877, n45878, n45879, n45880, n45881, n45882,
         n45883, n45884, n45885, n45886, n45887, n45888, n45889, n45890,
         n45891, n45892, n45893, n45894, n45895, n45896, n45897, n45898,
         n45899, n45900, n45901, n45902, n45903, n45904, n45905, n45906,
         n45907, n45908, n45909, n45910, n45911, n45912, n45913, n45914,
         n45915, n45916, n45917, n45918, n45919, n45920, n45921, n45922,
         n45923, n45924, n45925, n45926, n45927, n45928, n45929, n45930,
         n45931, n45932, n45933, n45934, n45935, n45936, n45937, n45938,
         n45939, n45940, n45941, n45942, n45943, n45944, n45945, n45946,
         n45947, n45948, n45949, n45950, n45951, n45952, n45953, n45954,
         n45955, n45956, n45957, n45958, n45959, n45960, n45961, n45962,
         n45963, n45964, n45965, n45966, n45967, n45968, n45969, n45970,
         n45971, n45972, n45973, n45974, n45975, n45976, n45977, n45978,
         n45979, n45980, n45981, n45982, n45983, n45984, n45985, n45986,
         n45987, n45988, n45989, n45990, n45991, n45992, n45993, n45994,
         n45995, n45996, n45997, n45998, n45999, n46000, n46001, n46002,
         n46003, n46004, n46005, n46006, n46007, n46008, n46009, n46010,
         n46011, n46012, n46013, n46014, n46015, n46016, n46017, n46018,
         n46019, n46020, n46021, n46022, n46023, n46024, n46025, n46026,
         n46027, n46028, n46029, n46030, n46031, n46032, n46033, n46034,
         n46035, n46036, n46037, n46038, n46039, n46040, n46041, n46042,
         n46043, n46044, n46045, n46046, n46047, n46048, n46049, n46050,
         n46051, n46052, n46053, n46054, n46055, n46056, n46057, n46058,
         n46059, n46060, n46061, n46062, n46063, n46064, n46065, n46066,
         n46067, n46068, n46069, n46070, n46071, n46072, n46073, n46074,
         n46075, n46076, n46077, n46078, n46079, n46080, n46081, n46082,
         n46083, n46084, n46085, n46086, n46087, n46088, n46089, n46090,
         n46091, n46092, n46093, n46094, n46095, n46096, n46097, n46098,
         n46099, n46100, n46101, n46102, n46103, n46104, n46105, n46106,
         n46107, n46108, n46109, n46110, n46111, n46112, n46113, n46114,
         n46115, n46116, n46117, n46118, n46119, n46120, n46121, n46122,
         n46123, n46124, n46125, n46126, n46127, n46128, n46129, n46130,
         n46131, n46132, n46133, n46134, n46135, n46136, n46137, n46138,
         n46139, n46140, n46141, n46142, n46143, n46144, n46145, n46146,
         n46147, n46148, n46149, n46150, n46151, n46152, n46153, n46154,
         n46155, n46156, n46157, n46158, n46159, n46160, n46161, n46162,
         n46163, n46164, n46165, n46166, n46167, n46168, n46169, n46170,
         n46171, n46172, n46173, n46174, n46175, n46176, n46177, n46178,
         n46179, n46180, n46181, n46182, n46183, n46184, n46185, n46186,
         n46187, n46188, n46189, n46190, n46191, n46192, n46193, n46194,
         n46195, n46196, n46197, n46198, n46199, n46200, n46201, n46202,
         n46203, n46204, n46205, n46206, n46207, n46208, n46209, n46210,
         n46211, n46212, n46213, n46214, n46215, n46216, n46217, n46218,
         n46219, n46220, n46221, n46222, n46223, n46224, n46225, n46226,
         n46227, n46228, n46229, n46230, n46231, n46232, n46233, n46234,
         n46235, n46236, n46237, n46238, n46239, n46240, n46241, n46242,
         n46243, n46244, n46245, n46246, n46247, n46248, n46249, n46250,
         n46251, n46252, n46253, n46254, n46255, n46256, n46257, n46258,
         n46259, n46260, n46261, n46262, n46263, n46264, n46265, n46266,
         n46267, n46268, n46269, n46270, n46271, n46272, n46273, n46274,
         n46275, n46276, n46277, n46278, n46279, n46280, n46281, n46282,
         n46283, n46284, n46285, n46286, n46287, n46288, n46289, n46290,
         n46291, n46292, n46293, n46294, n46295, n46296, n46297, n46298,
         n46299, n46300, n46301, n46302, n46303, n46304, n46305, n46306,
         n46307, n46308, n46309, n46310, n46311, n46312, n46313, n46314,
         n46315, n46316, n46317, n46318, n46319, n46320, n46321, n46322,
         n46323, n46324, n46325, n46326, n46327, n46328, n46329, n46330,
         n46331, n46332, n46333, n46334, n46335, n46336, n46337, n46338,
         n46339, n46340, n46341, n46342, n46343, n46344, n46345, n46346,
         n46347, n46348, n46349, n46350, n46351, n46352, n46353, n46354,
         n46355, n46356, n46357, n46358, n46359, n46360, n46361, n46362,
         n46363, n46364, n46365, n46366, n46367, n46368, n46369, n46370,
         n46371, n46372, n46373, n46374, n46375, n46376, n46377, n46378,
         n46379, n46380, n46381, n46382, n46383, n46384, n46385, n46386,
         n46387, n46388, n46389, n46390, n46391, n46392, n46393, n46394,
         n46395, n46396, n46397, n46398, n46399, n46400, n46401, n46402,
         n46403, n46404, n46405, n46406, n46407, n46408, n46409, n46410,
         n46411, n46412, n46413, n46414, n46415, n46416, n46417, n46418,
         n46419, n46420, n46421, n46422, n46423, n46424, n46425, n46426,
         n46427, n46428, n46429, n46430, n46431, n46432, n46433, n46434,
         n46435, n46436, n46437, n46438, n46439, n46440, n46441, n46442,
         n46443, n46444, n46445, n46446, n46447, n46448, n46449, n46450,
         n46451, n46452, n46453, n46454, n46455, n46456, n46457, n46458,
         n46459, n46460, n46461, n46462, n46463, n46464, n46465, n46466,
         n46467, n46468, n46469, n46470, n46471, n46472, n46473, n46474,
         n46475, n46476, n46477, n46478, n46479, n46480, n46481, n46482,
         n46483, n46484, n46485, n46486, n46487, n46488, n46489, n46490,
         n46491, n46492, n46493, n46494, n46495, n46496, n46497, n46498,
         n46499, n46500, n46501, n46502, n46503, n46504, n46505, n46506,
         n46507, n46508, n46509, n46510, n46511, n46512, n46513, n46514,
         n46515, n46516, n46517, n46518, n46519, n46520, n46521, n46522,
         n46523, n46524, n46525, n46526, n46527, n46528, n46529, n46530,
         n46531, n46532, n46533, n46534, n46535, n46536, n46537, n46538,
         n46539, n46540, n46541, n46542, n46543, n46544, n46545, n46546,
         n46547, n46548, n46549, n46550, n46551, n46552, n46553, n46554,
         n46555, n46556, n46557, n46558, n46559, n46560, n46561, n46562,
         n46563, n46564, n46565, n46566, n46567, n46568, n46569, n46570,
         n46571, n46572, n46573, n46574, n46575, n46576, n46577, n46578,
         n46579, n46580, n46581, n46582, n46583, n46584, n46585, n46586,
         n46587, n46588, n46589, n46590, n46591, n46592, n46593, n46594,
         n46595, n46596, n46597, n46598, n46599, n46600, n46601, n46602,
         n46603, n46604, n46605, n46606, n46607, n46608, n46609, n46610,
         n46611, n46612, n46613, n46614, n46615, n46616, n46617, n46618,
         n46619, n46620, n46621, n46622, n46623, n46624, n46625, n46626,
         n46627, n46628, n46629, n46630, n46631, n46632, n46633, n46634,
         n46635, n46636, n46637, n46638, n46639, n46640, n46641, n46642,
         n46643, n46644, n46645, n46646, n46647, n46648, n46649, n46650,
         n46651, n46652, n46653, n46654, n46655, n46656, n46657, n46658,
         n46659, n46660, n46661, n46662, n46663, n46664, n46665, n46666,
         n46667, n46668, n46669, n46670, n46671, n46672, n46673, n46674,
         n46675, n46676, n46677, n46678, n46679, n46680, n46681, n46682,
         n46683, n46684, n46685, n46686, n46687, n46688, n46689, n46690,
         n46691, n46692, n46693, n46694, n46695, n46696, n46697, n46698,
         n46699, n46700, n46701, n46702, n46703, n46704, n46705, n46706,
         n46707, n46708, n46709, n46710, n46711, n46712, n46713, n46714,
         n46715, n46716, n46717, n46718, n46719, n46720, n46721, n46722,
         n46723, n46724, n46725, n46726, n46727, n46728, n46729, n46730,
         n46731, n46732, n46733, n46734, n46735, n46736, n46737, n46738,
         n46739, n46740, n46741, n46742, n46743, n46744, n46745, n46746,
         n46747, n46748, n46749, n46750, n46751, n46752, n46753, n46754,
         n46755, n46756, n46757, n46758, n46759, n46760, n46761, n46762,
         n46763, n46764, n46765, n46766, n46767, n46768, n46769, n46770,
         n46771, n46772, n46773, n46774, n46775, n46776, n46777, n46778,
         n46779, n46780, n46781, n46782, n46783, n46784, n46785, n46786,
         n46787, n46788, n46789, n46790, n46791, n46792, n46793, n46794,
         n46795, n46796, n46797, n46798, n46799, n46800, n46801, n46802,
         n46803, n46804, n46805, n46806, n46807, n46808, n46809, n46810,
         n46811, n46812, n46813, n46814, n46815, n46816, n46817, n46818,
         n46819, n46820, n46821, n46822, n46823, n46824, n46825, n46826,
         n46827, n46828, n46829, n46830, n46831, n46832, n46833, n46834,
         n46835, n46836, n46837, n46838, n46839, n46840, n46841, n46842,
         n46843, n46844, n46845, n46846, n46847, n46848, n46849, n46850,
         n46851, n46852, n46853, n46854, n46855, n46856, n46857, n46858,
         n46859, n46860, n46861, n46862, n46863, n46864, n46865, n46866,
         n46867, n46868, n46869, n46870, n46871, n46872, n46873, n46874,
         n46875, n46876, n46877, n46878, n46879, n46880, n46881, n46882,
         n46883, n46884, n46885, n46886, n46887, n46888, n46889, n46890,
         n46891, n46892, n46893, n46894, n46895, n46896, n46897, n46898,
         n46899, n46900, n46901, n46902, n46903, n46904, n46905, n46906,
         n46907, n46908, n46909, n46910, n46911, n46912, n46913, n46914,
         n46915, n46916, n46917, n46918, n46919, n46920, n46921, n46922,
         n46923, n46924, n46925, n46926, n46927, n46928, n46929, n46930,
         n46931, n46932, n46933, n46934, n46935, n46936, n46937, n46938,
         n46939, n46940, n46941, n46942, n46943, n46944, n46945, n46946,
         n46947, n46948, n46949, n46950, n46951, n46952, n46953, n46954,
         n46955, n46956, n46957, n46958, n46959, n46960, n46961, n46962,
         n46963, n46964, n46965, n46966, n46967, n46968, n46969, n46970,
         n46971, n46972, n46973, n46974, n46975, n46976, n46977, n46978,
         n46979, n46980, n46981, n46982, n46983, n46984, n46985, n46986,
         n46987, n46988, n46989, n46990, n46991, n46992, n46993, n46994,
         n46995, n46996, n46997, n46998, n46999, n47000, n47001, n47002,
         n47003, n47004, n47005, n47006, n47007, n47008, n47009, n47010,
         n47011, n47012, n47013, n47014, n47015, n47016, n47017, n47018,
         n47019, n47020, n47021, n47022, n47023, n47024, n47025, n47026,
         n47027, n47028, n47029, n47030, n47031, n47032, n47033, n47034,
         n47035, n47036, n47037, n47038, n47039, n47040, n47041, n47042,
         n47043, n47044, n47045, n47046, n47047, n47048, n47049, n47050,
         n47051, n47052, n47053, n47054, n47055, n47056, n47057, n47058,
         n47059, n47060, n47061, n47062, n47063, n47064, n47065, n47066,
         n47067, n47068, n47069, n47070, n47071, n47072, n47073, n47074,
         n47075, n47076, n47077, n47078, n47079, n47080, n47081, n47082,
         n47083, n47084, n47085, n47086, n47087, n47088, n47089, n47090,
         n47091, n47092, n47093, n47094, n47095, n47096, n47097, n47098,
         n47099, n47100, n47101, n47102, n47103, n47104, n47105, n47106,
         n47107, n47108, n47109, n47110, n47111, n47112, n47113, n47114,
         n47115, n47116, n47117, n47118, n47119, n47120, n47121, n47122,
         n47123, n47124, n47125, n47126, n47127, n47128, n47129, n47130,
         n47131, n47132, n47133, n47134, n47135, n47136, n47137, n47138,
         n47139, n47140, n47141, n47142, n47143, n47144, n47145, n47146,
         n47147, n47148, n47149, n47150, n47151, n47152, n47153, n47154,
         n47155, n47156, n47157, n47158, n47159, n47160, n47161, n47162,
         n47163, n47164, n47165, n47166, n47167, n47168, n47169, n47170,
         n47171, n47172, n47173, n47174, n47175, n47176, n47177, n47178,
         n47179, n47180, n47181, n47182, n47183, n47184, n47185, n47186,
         n47187, n47188, n47189, n47190, n47191, n47192, n47193, n47194,
         n47195, n47196, n47197, n47198, n47199, n47200, n47201, n47202,
         n47203, n47204, n47205, n47206, n47207, n47208, n47209, n47210,
         n47211, n47212, n47213, n47214, n47215, n47216, n47217, n47218,
         n47219, n47220, n47221, n47222, n47223, n47224, n47225, n47226,
         n47227, n47228, n47229, n47230, n47231, n47232, n47233, n47234,
         n47235, n47236, n47237, n47238, n47239, n47240, n47241, n47242,
         n47243, n47244, n47245, n47246, n47247, n47248, n47249, n47250,
         n47251, n47252, n47253, n47254, n47255, n47256, n47257, n47258,
         n47259, n47260, n47261, n47262, n47263, n47264, n47265, n47266,
         n47267, n47268, n47269, n47270, n47271, n47272, n47273, n47274,
         n47275, n47276, n47277, n47278, n47279, n47280, n47281, n47282,
         n47283, n47284, n47285, n47286, n47287, n47288, n47289, n47290,
         n47291, n47292, n47293, n47294, n47295, n47296, n47297, n47298,
         n47299, n47300, n47301, n47302, n47303, n47304, n47305, n47306,
         n47307, n47308, n47309, n47310, n47311, n47312, n47313, n47314,
         n47315, n47316, n47317, n47318, n47319, n47320, n47321, n47322,
         n47323, n47324, n47325, n47326, n47327, n47328, n47329, n47330,
         n47331, n47332, n47333, n47334, n47335, n47336, n47337, n47338,
         n47339, n47340, n47341, n47342, n47343, n47344, n47345, n47346,
         n47347, n47348, n47349, n47350, n47351, n47352, n47353, n47354,
         n47355, n47356, n47357, n47358, n47359, n47360, n47361, n47362,
         n47363, n47364, n47365, n47366, n47367, n47368, n47369, n47370,
         n47371, n47372, n47373, n47374, n47375, n47376, n47377, n47378,
         n47379, n47380, n47381, n47382, n47383, n47384, n47385, n47386,
         n47387, n47388, n47389, n47390, n47391, n47392, n47393, n47394,
         n47395, n47396, n47397, n47398, n47399, n47400, n47401, n47402,
         n47403, n47404, n47405, n47406, n47407, n47408, n47409, n47410,
         n47411, n47412, n47413, n47414, n47415, n47416, n47417, n47418,
         n47419, n47420, n47421, n47422, n47423, n47424, n47425, n47426,
         n47427, n47428, n47429, n47430, n47431, n47432, n47433, n47434,
         n47435, n47436, n47437, n47438, n47439, n47440, n47441, n47442,
         n47443, n47444, n47445, n47446, n47447, n47448, n47449, n47450,
         n47451, n47452, n47453, n47454, n47455, n47456, n47457, n47458,
         n47459, n47460, n47461, n47462, n47463, n47464, n47465, n47466,
         n47467, n47468, n47469, n47470, n47471, n47472, n47473, n47474,
         n47475, n47476, n47477, n47478, n47479, n47480, n47481, n47482,
         n47483, n47484, n47485, n47486, n47487, n47488, n47489, n47490,
         n47491, n47492, n47493, n47494, n47495, n47496, n47497, n47498,
         n47499, n47500, n47501, n47502, n47503, n47504, n47505, n47506,
         n47507, n47508, n47509, n47510, n47511, n47512, n47513, n47514,
         n47515, n47516, n47517, n47518, n47519, n47520, n47521, n47522,
         n47523, n47524, n47525, n47526, n47527, n47528, n47529, n47530,
         n47531, n47532, n47533, n47534, n47535, n47536, n47537, n47538,
         n47539, n47540, n47541, n47542, n47543, n47544, n47545, n47546,
         n47547, n47548, n47549, n47550, n47551, n47552, n47553, n47554,
         n47555, n47556, n47557, n47558, n47559, n47560, n47561, n47562,
         n47563, n47564, n47565, n47566, n47567, n47568, n47569, n47570,
         n47571, n47572, n47573, n47574, n47575, n47576, n47577, n47578,
         n47579, n47580, n47581, n47582, n47583, n47584, n47585, n47586,
         n47587, n47588, n47589, n47590, n47591, n47592, n47593, n47594,
         n47595, n47596, n47597, n47598, n47599, n47600, n47601, n47602,
         n47603, n47604, n47605, n47606, n47607, n47608, n47609, n47610,
         n47611, n47612, n47613, n47614, n47615, n47616, n47617, n47618,
         n47619, n47620, n47621, n47622, n47623, n47624, n47625, n47626,
         n47627, n47628, n47629, n47630, n47631, n47632, n47633, n47634,
         n47635, n47636, n47637, n47638, n47639, n47640, n47641, n47642,
         n47643, n47644, n47645, n47646, n47647, n47648, n47649, n47650,
         n47651, n47652, n47653, n47654, n47655, n47656, n47657, n47658,
         n47659, n47660, n47661, n47662, n47663, n47664, n47665, n47666,
         n47667, n47668, n47669, n47670, n47671, n47672, n47673, n47674,
         n47675, n47676, n47677, n47678, n47679, n47680, n47681, n47682,
         n47683, n47684, n47685, n47686, n47687, n47688, n47689, n47690,
         n47691, n47692, n47693, n47694, n47695, n47696, n47697, n47698,
         n47699, n47700, n47701, n47702, n47703, n47704, n47705, n47706,
         n47707, n47708, n47709, n47710, n47711, n47712, n47713, n47714,
         n47715, n47716, n47717, n47718, n47719, n47720, n47721, n47722,
         n47723, n47724, n47725, n47726, n47727, n47728, n47729, n47730,
         n47731, n47732, n47733, n47734, n47735, n47736, n47737, n47738,
         n47739, n47740, n47741, n47742, n47743, n47744, n47745, n47746,
         n47747, n47748, n47749, n47750, n47751, n47752, n47753, n47754,
         n47755, n47756, n47757, n47758, n47759, n47760, n47761, n47762,
         n47763, n47764, n47765, n47766, n47767, n47768, n47769, n47770,
         n47771, n47772, n47773, n47774, n47775, n47776, n47777, n47778,
         n47779, n47780, n47781, n47782, n47783, n47784, n47785, n47786,
         n47787, n47788, n47789, n47790, n47791, n47792, n47793, n47794,
         n47795, n47796, n47797, n47798, n47799, n47800, n47801, n47802,
         n47803, n47804, n47805, n47806, n47807, n47808, n47809, n47810,
         n47811, n47812, n47813, n47814, n47815, n47816, n47817, n47818,
         n47819, n47820, n47821, n47822, n47823, n47824, n47825, n47826,
         n47827, n47828, n47829, n47830, n47831, n47832, n47833, n47834,
         n47835, n47836, n47837, n47838, n47839, n47840, n47841, n47842,
         n47843, n47844, n47845, n47846, n47847, n47848, n47849, n47850,
         n47851, n47852, n47853, n47854, n47855, n47856, n47857, n47858,
         n47859, n47860, n47861, n47862, n47863, n47864, n47865, n47866,
         n47867, n47868, n47869, n47870, n47871, n47872, n47873, n47874,
         n47875, n47876, n47877, n47878, n47879, n47880, n47881, n47882,
         n47883, n47884, n47885, n47886, n47887, n47888, n47889, n47890,
         n47891, n47892, n47893, n47894, n47895, n47896, n47897, n47898,
         n47899, n47900, n47901, n47902, n47903, n47904, n47905, n47906,
         n47907, n47908, n47909, n47910, n47911, n47912, n47913, n47914,
         n47915, n47916, n47917, n47918, n47919, n47920, n47921, n47922,
         n47923, n47924, n47925, n47926, n47927, n47928, n47929, n47930,
         n47931, n47932, n47933, n47934, n47935, n47936, n47937, n47938,
         n47939, n47940, n47941, n47942, n47943, n47944, n47945, n47946,
         n47947, n47948, n47949, n47950, n47951, n47952, n47953, n47954,
         n47955, n47956, n47957, n47958, n47959, n47960, n47961, n47962,
         n47963, n47964, n47965, n47966, n47967, n47968, n47969, n47970,
         n47971, n47972, n47973, n47974, n47975, n47976, n47977, n47978,
         n47979, n47980, n47981, n47982, n47983, n47984, n47985, n47986,
         n47987, n47988, n47989, n47990, n47991, n47992, n47993, n47994,
         n47995, n47996, n47997, n47998, n47999, n48000, n48001, n48002,
         n48003, n48004, n48005, n48006, n48007, n48008, n48009, n48010,
         n48011, n48012, n48013, n48014, n48015, n48016, n48017, n48018,
         n48019, n48020, n48021, n48022, n48023, n48024, n48025, n48026,
         n48027, n48028, n48029, n48030, n48031, n48032, n48033, n48034,
         n48035, n48036, n48037, n48038, n48039, n48040, n48041, n48042,
         n48043, n48044, n48045, n48046, n48047, n48048, n48049, n48050,
         n48051, n48052, n48053, n48054, n48055, n48056, n48057, n48058,
         n48059, n48060, n48061, n48062, n48063, n48064, n48065, n48066,
         n48067, n48068, n48069, n48070, n48071, n48072, n48073, n48074,
         n48075, n48076, n48077, n48078, n48079, n48080, n48081, n48082,
         n48083, n48084, n48085, n48086, n48087, n48088, n48089, n48090,
         n48091, n48092, n48093, n48094, n48095, n48096, n48097, n48098,
         n48099, n48100, n48101, n48102, n48103, n48104, n48105, n48106,
         n48107, n48108, n48109, n48110, n48111, n48112, n48113, n48114,
         n48115, n48116, n48117, n48118, n48119, n48120, n48121, n48122,
         n48123, n48124, n48125, n48126, n48127, n48128, n48129, n48130,
         n48131, n48132, n48133, n48134, n48135, n48136, n48137, n48138,
         n48139, n48140, n48141, n48142, n48143, n48144, n48145, n48146,
         n48147, n48148, n48149, n48150, n48151, n48152, n48153, n48154,
         n48155, n48156, n48157, n48158, n48159, n48160, n48161, n48162,
         n48163, n48164, n48165, n48166, n48167, n48168, n48169, n48170,
         n48171, n48172, n48173, n48174, n48175, n48176, n48177, n48178,
         n48179, n48180, n48181, n48182, n48183, n48184, n48185, n48186,
         n48187, n48188, n48189, n48190, n48191, n48192, n48193, n48194,
         n48195, n48196, n48197, n48198, n48199, n48200, n48201, n48202,
         n48203, n48204, n48205, n48206, n48207, n48208, n48209, n48210,
         n48211, n48212, n48213, n48214, n48215, n48216, n48217, n48218,
         n48219, n48220, n48221, n48222, n48223, n48224, n48225, n48226,
         n48227, n48228, n48229, n48230, n48231, n48232, n48233, n48234,
         n48235, n48236, n48237, n48238, n48239, n48240, n48241, n48242,
         n48243, n48244, n48245, n48246, n48247, n48248, n48249, n48250,
         n48251, n48252, n48253, n48254, n48255, n48256, n48257, n48258,
         n48259, n48260, n48261, n48262, n48263, n48264, n48265, n48266,
         n48267, n48268, n48269, n48270, n48271, n48272, n48273, n48274,
         n48275, n48276, n48277, n48278, n48279, n48280, n48281, n48282,
         n48283, n48284, n48285, n48286, n48287, n48288, n48289, n48290,
         n48291, n48292, n48293, n48294, n48295, n48296, n48297, n48298,
         n48299, n48300, n48301, n48302, n48303, n48304, n48305, n48306,
         n48307, n48308, n48309, n48310, n48311, n48312, n48313, n48314,
         n48315, n48316, n48317, n48318, n48319, n48320, n48321, n48322,
         n48323, n48324, n48325, n48326, n48327, n48328, n48329, n48330,
         n48331, n48332, n48333, n48334, n48335, n48336, n48337, n48338,
         n48339, n48340, n48341, n48342, n48343, n48344, n48345, n48346,
         n48347, n48348, n48349, n48350, n48351, n48352, n48353, n48354,
         n48355, n48356, n48357, n48358, n48359, n48360, n48361, n48362,
         n48363, n48364, n48365, n48366, n48367, n48368, n48369, n48370,
         n48371, n48372, n48373, n48374, n48375, n48376, n48377, n48378,
         n48379, n48380, n48381, n48382, n48383, n48384, n48385, n48386,
         n48387, n48388, n48389, n48390, n48391, n48392, n48393, n48394,
         n48395, n48396, n48397, n48398, n48399, n48400, n48401, n48402,
         n48403, n48404, n48405, n48406, n48407, n48408, n48409, n48410,
         n48411, n48412, n48413, n48414, n48415, n48416, n48417, n48418,
         n48419, n48420, n48421, n48422, n48423, n48424, n48425, n48426,
         n48427, n48428, n48429, n48430, n48431, n48432, n48433, n48434,
         n48435, n48436, n48437, n48438, n48439, n48440, n48441, n48442,
         n48443, n48444, n48445, n48446, n48447, n48448, n48449, n48450,
         n48451, n48452, n48453, n48454, n48455, n48456, n48457, n48458,
         n48459, n48460, n48461, n48462, n48463, n48464, n48465, n48466,
         n48467, n48468, n48469, n48470, n48471, n48472, n48473, n48474,
         n48475, n48476, n48477, n48478, n48479, n48480, n48481, n48482,
         n48483, n48484, n48485, n48486, n48487, n48488, n48489, n48490,
         n48491, n48492, n48493, n48494, n48495, n48496, n48497, n48498,
         n48499, n48500, n48501, n48502, n48503, n48504, n48505, n48506,
         n48507, n48508, n48509, n48510, n48511, n48512, n48513, n48514,
         n48515, n48516, n48517, n48518, n48519, n48520, n48521, n48522,
         n48523, n48524, n48525, n48526, n48527, n48528, n48529, n48530,
         n48531, n48532, n48533, n48534, n48535, n48536, n48537, n48538,
         n48539, n48540, n48541, n48542, n48543, n48544, n48545, n48546,
         n48547, n48548, n48549, n48550, n48551, n48552, n48553, n48554,
         n48555, n48556, n48557, n48558, n48559, n48560, n48561, n48562,
         n48563, n48564, n48565, n48566, n48567, n48568, n48569, n48570,
         n48571, n48572, n48573, n48574, n48575, n48576, n48577, n48578,
         n48579, n48580, n48581, n48582, n48583, n48584, n48585, n48586,
         n48587, n48588, n48589, n48590, n48591, n48592, n48593, n48594,
         n48595, n48596, n48597, n48598, n48599, n48600, n48601, n48602,
         n48603, n48604, n48605, n48606, n48607, n48608, n48609, n48610,
         n48611, n48612, n48613, n48614, n48615, n48616, n48617, n48618,
         n48619, n48620, n48621, n48622, n48623, n48624, n48625, n48626,
         n48627, n48628, n48629, n48630, n48631, n48632, n48633, n48634,
         n48635, n48636, n48637, n48638, n48639, n48640, n48641, n48642,
         n48643, n48644, n48645, n48646, n48647, n48648, n48649, n48650,
         n48651, n48652, n48653, n48654, n48655, n48656, n48657, n48658,
         n48659, n48660, n48661, n48662, n48663, n48664, n48665, n48666,
         n48667, n48668, n48669, n48670, n48671, n48672, n48673, n48674,
         n48675, n48676, n48677, n48678, n48679, n48680, n48681, n48682,
         n48683, n48684, n48685, n48686, n48687, n48688, n48689, n48690,
         n48691, n48692, n48693, n48694, n48695, n48696, n48697, n48698,
         n48699, n48700, n48701, n48702, n48703, n48704, n48705, n48706,
         n48707, n48708, n48709, n48710, n48711, n48712, n48713, n48714,
         n48715, n48716, n48717, n48718, n48719, n48720, n48721, n48722,
         n48723, n48724, n48725, n48726, n48727, n48728, n48729, n48730,
         n48731, n48732, n48733, n48734, n48735, n48736, n48737, n48738,
         n48739, n48740, n48741, n48742, n48743, n48744, n48745, n48746,
         n48747, n48748, n48749, n48750, n48751, n48752, n48753, n48754,
         n48755, n48756, n48757, n48758, n48759, n48760, n48761, n48762,
         n48763, n48764, n48765, n48766, n48767, n48768, n48769, n48770,
         n48771, n48772, n48773, n48774, n48775, n48776, n48777, n48778,
         n48779, n48780, n48781, n48782, n48783, n48784, n48785, n48786,
         n48787, n48788, n48789, n48790, n48791, n48792, n48793, n48794,
         n48795, n48796, n48797, n48798, n48799, n48800, n48801, n48802,
         n48803, n48804, n48805, n48806, n48807, n48808, n48809, n48810,
         n48811, n48812, n48813, n48814, n48815, n48816, n48817, n48818,
         n48819, n48820, n48821, n48822, n48823, n48824, n48825, n48826,
         n48827, n48828, n48829, n48830, n48831, n48832, n48833, n48834,
         n48835, n48836, n48837, n48838, n48839, n48840, n48841, n48842,
         n48843, n48844, n48845, n48846, n48847, n48848, n48849, n48850,
         n48851, n48852, n48853, n48854, n48855, n48856, n48857, n48858,
         n48859, n48860, n48861, n48862, n48863, n48864, n48865, n48866,
         n48867, n48868, n48869, n48870, n48871, n48872, n48873, n48874,
         n48875, n48876, n48877, n48878, n48879, n48880, n48881, n48882,
         n48883, n48884, n48885, n48886, n48887, n48888, n48889, n48890,
         n48891, n48892, n48893, n48894, n48895, n48896, n48897, n48898,
         n48899, n48900, n48901, n48902, n48903, n48904, n48905, n48906,
         n48907, n48908, n48909, n48910, n48911, n48912, n48913, n48914,
         n48915, n48916, n48917, n48918, n48919, n48920, n48921, n48922,
         n48923, n48924, n48925, n48926, n48927, n48928, n48929, n48930,
         n48931, n48932, n48933, n48934, n48935, n48936, n48937, n48938,
         n48939, n48940, n48941, n48942, n48943, n48944, n48945, n48946,
         n48947, n48948, n48949, n48950, n48951, n48952, n48953, n48954,
         n48955, n48956, n48957, n48958, n48959, n48960, n48961, n48962,
         n48963, n48964, n48965, n48966, n48967, n48968, n48969, n48970,
         n48971, n48972, n48973, n48974, n48975, n48976, n48977, n48978,
         n48979, n48980, n48981, n48982, n48983, n48984, n48985, n48986,
         n48987, n48988, n48989, n48990, n48991, n48992, n48993, n48994,
         n48995, n48996, n48997, n48998, n48999, n49000, n49001, n49002,
         n49003, n49004, n49005, n49006, n49007, n49008, n49009, n49010,
         n49011, n49012, n49013, n49014, n49015, n49016, n49017, n49018,
         n49019, n49020, n49021, n49022, n49023, n49024, n49025, n49026,
         n49027, n49028, n49029, n49030, n49031, n49032, n49033, n49034,
         n49035, n49036, n49037, n49038, n49039, n49040, n49041, n49042,
         n49043, n49044, n49045, n49046, n49047, n49048, n49049, n49050,
         n49051, n49052, n49053, n49054, n49055, n49056, n49057, n49058,
         n49059, n49060, n49061, n49062, n49063, n49064, n49065, n49066,
         n49067, n49068, n49069, n49070, n49071, n49072, n49073, n49074,
         n49075, n49076, n49077, n49078, n49079, n49080, n49081, n49082,
         n49083, n49084, n49085, n49086, n49087, n49088, n49089, n49090,
         n49091, n49092, n49093, n49094, n49095, n49096, n49097, n49098,
         n49099, n49100, n49101, n49102, n49103, n49104, n49105, n49106,
         n49107, n49108, n49109, n49110, n49111, n49112, n49113, n49114,
         n49115, n49116, n49117, n49118, n49119, n49120, n49121, n49122,
         n49123, n49124, n49125, n49126, n49127, n49128, n49129, n49130,
         n49131, n49132, n49133, n49134, n49135, n49136, n49137, n49138,
         n49139, n49140, n49141, n49142, n49143, n49144, n49145, n49146,
         n49147, n49148, n49149, n49150, n49151, n49152, n49153, n49154,
         n49155, n49156, n49157, n49158, n49159, n49160, n49161, n49162,
         n49163, n49164, n49165, n49166, n49167, n49168, n49169, n49170,
         n49171, n49172, n49173, n49174, n49175, n49176, n49177, n49178,
         n49179, n49180, n49181, n49182, n49183, n49184, n49185, n49186,
         n49187, n49188, n49189, n49190, n49191, n49192, n49193, n49194,
         n49195, n49196, n49197, n49198, n49199, n49200, n49201, n49202,
         n49203, n49204, n49205, n49206, n49207, n49208, n49209, n49210,
         n49211, n49212, n49213, n49214, n49215, n49216, n49217, n49218,
         n49219, n49220, n49221, n49222, n49223, n49224, n49225, n49226,
         n49227, n49228, n49229, n49230, n49231, n49232, n49233, n49234,
         n49235, n49236, n49237, n49238, n49239, n49240, n49241, n49242,
         n49243, n49244, n49245, n49246, n49247, n49248, n49249, n49250,
         n49251, n49252, n49253, n49254, n49255, n49256, n49257, n49258,
         n49259, n49260, n49261, n49262, n49263, n49264, n49265, n49266,
         n49267, n49268, n49269, n49270, n49271, n49272, n49273, n49274,
         n49275, n49276, n49277, n49278, n49279, n49280, n49281, n49282,
         n49283, n49284, n49285, n49286, n49287, n49288, n49289, n49290,
         n49291, n49292, n49293, n49294, n49295, n49296, n49297, n49298,
         n49299, n49300, n49301, n49302, n49303, n49304, n49305, n49306,
         n49307, n49308, n49309, n49310, n49311, n49312, n49313, n49314,
         n49315, n49316, n49317, n49318, n49319, n49320, n49321, n49322,
         n49323, n49324, n49325, n49326, n49327, n49328, n49329, n49330,
         n49331, n49332, n49333, n49334, n49335, n49336, n49337, n49338,
         n49339, n49340, n49341, n49342, n49343, n49344, n49345, n49346,
         n49347, n49348, n49349, n49350, n49351, n49352, n49353, n49354,
         n49355, n49356, n49357, n49358, n49359, n49360, n49361, n49362,
         n49363, n49364, n49365, n49366, n49367, n49368, n49369, n49370,
         n49371, n49372, n49373, n49374, n49375, n49376, n49377, n49378,
         n49379, n49380, n49381, n49382, n49383, n49384, n49385, n49386,
         n49387, n49388, n49389, n49390, n49391, n49392, n49393, n49394,
         n49395, n49396, n49397, n49398, n49399, n49400, n49401, n49402,
         n49403, n49404, n49405, n49406, n49407, n49408, n49409, n49410,
         n49411, n49412, n49413, n49414, n49415, n49416, n49417, n49418,
         n49419, n49420, n49421, n49422, n49423, n49424, n49425, n49426,
         n49427, n49428, n49429, n49430, n49431, n49432, n49433, n49434,
         n49435, n49436, n49437, n49438, n49439, n49440, n49441, n49442,
         n49443, n49444, n49445, n49446, n49447, n49448, n49449, n49450,
         n49451, n49452, n49453, n49454, n49455, n49456, n49457, n49458,
         n49459, n49460, n49461, n49462, n49463, n49464, n49465, n49466,
         n49467, n49468, n49469, n49470, n49471, n49472, n49473, n49474,
         n49475, n49476, n49477, n49478, n49479, n49480, n49481, n49482,
         n49483, n49484, n49485, n49486, n49487, n49488, n49489, n49490,
         n49491, n49492, n49493, n49494, n49495, n49496, n49497, n49498,
         n49499, n49500, n49501, n49502, n49503, n49504, n49505, n49506,
         n49507, n49508, n49509, n49510, n49511, n49512, n49513, n49514,
         n49515, n49516, n49517, n49518, n49519, n49520, n49521, n49522,
         n49523, n49524, n49525, n49526, n49527, n49528, n49529, n49530,
         n49531, n49532, n49533, n49534, n49535, n49536, n49537, n49538,
         n49539, n49540, n49541, n49542, n49543, n49544, n49545, n49546,
         n49547, n49548, n49549, n49550, n49551, n49552, n49553, n49554,
         n49555, n49556, n49557, n49558, n49559, n49560, n49561, n49562,
         n49563, n49564, n49565, n49566, n49567, n49568, n49569, n49570,
         n49571, n49572, n49573, n49574, n49575, n49576, n49577, n49578,
         n49579, n49580, n49581, n49582, n49583, n49584, n49585, n49586,
         n49587, n49588, n49589, n49590, n49591, n49592, n49593, n49594,
         n49595, n49596, n49597, n49598, n49599, n49600, n49601, n49602,
         n49603, n49604, n49605, n49606, n49607, n49608, n49609, n49610,
         n49611, n49612, n49613, n49614, n49615, n49616, n49617, n49618,
         n49619, n49620, n49621, n49622, n49623, n49624, n49625, n49626,
         n49627, n49628, n49629, n49630, n49631, n49632, n49633, n49634,
         n49635, n49636, n49637, n49638, n49639, n49640, n49641, n49642,
         n49643, n49644, n49645, n49646, n49647, n49648, n49649, n49650,
         n49651, n49652, n49653, n49654, n49655, n49656, n49657, n49658,
         n49659, n49660, n49661, n49662, n49663, n49664, n49665, n49666,
         n49667, n49668, n49669, n49670, n49671, n49672, n49673, n49674,
         n49675, n49676, n49677, n49678, n49679, n49680, n49681, n49682,
         n49683, n49684, n49685, n49686, n49687, n49688, n49689, n49690,
         n49691, n49692, n49693, n49694, n49695, n49696, n49697, n49698,
         n49699, n49700, n49701, n49702, n49703, n49704, n49705, n49706,
         n49707, n49708, n49709, n49710, n49711, n49712, n49713, n49714,
         n49715, n49716, n49717, n49718, n49719, n49720, n49721, n49722,
         n49723, n49724, n49725, n49726, n49727, n49728, n49729, n49730,
         n49731, n49732, n49733, n49734, n49735, n49736, n49737, n49738,
         n49739, n49740, n49741, n49742, n49743, n49744, n49745, n49746,
         n49747, n49748, n49749, n49750, n49751, n49752, n49753, n49754,
         n49755, n49756, n49757, n49758, n49759, n49760, n49761, n49762,
         n49763, n49764, n49765, n49766, n49767, n49768, n49769, n49770,
         n49771, n49772, n49773, n49774, n49775, n49776, n49777, n49778,
         n49779, n49780, n49781, n49782, n49783, n49784, n49785, n49786,
         n49787, n49788, n49789, n49790, n49791, n49792, n49793, n49794,
         n49795, n49796, n49797, n49798, n49799, n49800, n49801, n49802,
         n49803, n49804, n49805, n49806, n49807, n49808, n49809, n49810,
         n49811, n49812, n49813, n49814, n49815, n49816, n49817, n49818,
         n49819, n49820, n49821, n49822, n49823, n49824, n49825, n49826,
         n49827, n49828, n49829, n49830, n49831, n49832, n49833, n49834,
         n49835, n49836, n49837, n49838, n49839, n49840, n49841, n49842,
         n49843, n49844, n49845, n49846, n49847, n49848, n49849, n49850,
         n49851, n49852, n49853, n49854, n49855, n49856, n49857, n49858,
         n49859, n49860, n49861, n49862, n49863, n49864, n49865, n49866,
         n49867, n49868, n49869, n49870, n49871, n49872, n49873, n49874,
         n49875, n49876, n49877, n49878, n49879, n49880, n49881, n49882,
         n49883, n49884, n49885, n49886, n49887, n49888, n49889, n49890,
         n49891, n49892, n49893, n49894, n49895, n49896, n49897, n49898,
         n49899, n49900, n49901, n49902, n49903, n49904, n49905, n49906,
         n49907, n49908, n49909, n49910, n49911, n49912, n49913, n49914,
         n49915, n49916, n49917, n49918, n49919, n49920, n49921, n49922,
         n49923, n49924, n49925, n49926, n49927, n49928, n49929, n49930,
         n49931, n49932, n49933, n49934, n49935, n49936, n49937, n49938,
         n49939, n49940, n49941, n49942, n49943, n49944, n49945, n49946,
         n49947, n49948, n49949, n49950, n49951, n49952, n49953, n49954,
         n49955, n49956, n49957, n49958, n49959, n49960, n49961, n49962,
         n49963, n49964, n49965, n49966, n49967, n49968, n49969, n49970,
         n49971, n49972, n49973, n49974, n49975, n49976, n49977, n49978,
         n49979, n49980, n49981, n49982, n49983, n49984, n49985, n49986,
         n49987, n49988, n49989, n49990, n49991, n49992, n49993, n49994,
         n49995, n49996, n49997, n49998, n49999, n50000, n50001, n50002,
         n50003, n50004, n50005, n50006, n50007, n50008, n50009, n50010,
         n50011, n50012, n50013, n50014, n50015, n50016, n50017, n50018,
         n50019, n50020, n50021, n50022, n50023, n50024, n50025, n50026,
         n50027, n50028, n50029, n50030, n50031, n50032, n50033, n50034,
         n50035, n50036, n50037, n50038, n50039, n50040, n50041, n50042,
         n50043, n50044, n50045, n50046, n50047, n50048, n50049, n50050,
         n50051, n50052, n50053, n50054, n50055, n50056, n50057, n50058,
         n50059, n50060, n50061, n50062, n50063, n50064, n50065, n50066,
         n50067, n50068, n50069, n50070, n50071, n50072, n50073, n50074,
         n50075, n50076, n50077, n50078, n50079, n50080, n50081, n50082,
         n50083, n50084, n50085, n50086, n50087, n50088, n50089, n50090,
         n50091, n50092, n50093, n50094, n50095, n50096, n50097, n50098,
         n50099, n50100, n50101, n50102, n50103, n50104, n50105, n50106,
         n50107, n50108, n50109, n50110, n50111, n50112, n50113, n50114,
         n50115, n50116, n50117, n50118, n50119, n50120, n50121, n50122,
         n50123, n50124, n50125, n50126, n50127, n50128, n50129, n50130,
         n50131, n50132, n50133, n50134, n50135, n50136, n50137, n50138,
         n50139, n50140, n50141, n50142, n50143, n50144, n50145, n50146,
         n50147, n50148, n50149, n50150, n50151, n50152, n50153, n50154,
         n50155, n50156, n50157, n50158, n50159, n50160, n50161, n50162,
         n50163, n50164, n50165, n50166, n50167, n50168, n50169, n50170,
         n50171, n50172, n50173, n50174, n50175, n50176, n50177, n50178,
         n50179, n50180, n50181, n50182, n50183, n50184, n50185, n50186,
         n50187, n50188, n50189, n50190, n50191, n50192, n50193, n50194,
         n50195, n50196, n50197, n50198, n50199, n50200, n50201, n50202,
         n50203, n50204, n50205, n50206, n50207, n50208, n50209, n50210,
         n50211, n50212, n50213, n50214, n50215, n50216, n50217, n50218,
         n50219, n50220, n50221, n50222, n50223, n50224, n50225, n50226,
         n50227, n50228, n50229, n50230, n50231, n50232, n50233, n50234,
         n50235, n50236, n50237, n50238, n50239, n50240, n50241, n50242,
         n50243, n50244, n50245, n50246, n50247, n50248, n50249, n50250,
         n50251, n50252, n50253, n50254, n50255, n50256, n50257, n50258,
         n50259, n50260, n50261, n50262, n50263, n50264, n50265, n50266,
         n50267, n50268, n50269, n50270, n50271, n50272, n50273, n50274,
         n50275, n50276, n50277, n50278, n50279, n50280, n50281, n50282,
         n50283, n50284, n50285, n50286, n50287, n50288, n50289, n50290,
         n50291, n50292, n50293, n50294, n50295, n50296, n50297, n50298,
         n50299, n50300, n50301, n50302, n50303, n50304, n50305, n50306,
         n50307, n50308, n50309, n50310, n50311, n50312, n50313, n50314,
         n50315, n50316, n50317, n50318, n50319, n50320, n50321, n50322,
         n50323, n50324, n50325, n50326, n50327, n50328, n50329, n50330,
         n50331, n50332, n50333, n50334, n50335, n50336, n50337, n50338,
         n50339, n50340, n50341, n50342, n50343, n50344, n50345, n50346,
         n50347, n50348, n50349, n50350, n50351, n50352, n50353, n50354,
         n50355, n50356, n50357, n50358, n50359, n50360, n50361, n50362,
         n50363, n50364, n50365, n50366, n50367, n50368, n50369, n50370,
         n50371, n50372, n50373, n50374, n50375, n50376, n50377, n50378,
         n50379, n50380, n50381, n50382, n50383, n50384, n50385, n50386,
         n50387, n50388, n50389, n50390, n50391, n50392, n50393, n50394,
         n50395, n50396, n50397, n50398, n50399, n50400, n50401, n50402,
         n50403, n50404, n50405, n50406, n50407, n50408, n50409, n50410,
         n50411, n50412, n50413, n50414, n50415, n50416, n50417, n50418,
         n50419, n50420, n50421, n50422, n50423, n50424, n50425, n50426,
         n50427, n50428, n50429, n50430, n50431, n50432, n50433, n50434,
         n50435, n50436, n50437, n50438, n50439, n50440, n50441, n50442,
         n50443, n50444, n50445, n50446, n50447, n50448, n50449, n50450,
         n50451, n50452, n50453, n50454, n50455, n50456, n50457, n50458,
         n50459, n50460, n50461, n50462, n50463, n50464, n50465, n50466,
         n50467, n50468, n50469, n50470, n50471, n50472, n50473, n50474,
         n50475, n50476, n50477, n50478, n50479, n50480, n50481, n50482,
         n50483, n50484, n50485, n50486, n50487, n50488, n50489, n50490,
         n50491, n50492, n50493, n50494, n50495, n50496, n50497, n50498,
         n50499, n50500, n50501, n50502, n50503, n50504, n50505, n50506,
         n50507, n50508, n50509, n50510, n50511, n50512, n50513, n50514,
         n50515, n50516, n50517, n50518, n50519, n50520, n50521, n50522,
         n50523, n50524, n50525, n50526, n50527, n50528, n50529, n50530,
         n50531, n50532, n50533, n50534, n50535, n50536, n50537, n50538,
         n50539, n50540, n50541, n50542, n50543, n50544, n50545, n50546,
         n50547, n50548, n50549, n50550, n50551, n50552, n50553, n50554,
         n50555, n50556, n50557, n50558, n50559, n50560, n50561, n50562,
         n50563, n50564, n50565, n50566, n50567, n50568, n50569, n50570,
         n50571, n50572, n50573, n50574, n50575, n50576, n50577, n50578,
         n50579, n50580, n50581, n50582, n50583, n50584, n50585, n50586,
         n50587, n50588, n50589, n50590, n50591, n50592, n50593, n50594,
         n50595, n50596, n50597, n50598, n50599, n50600, n50601, n50602,
         n50603, n50604, n50605, n50606, n50607, n50608, n50609, n50610,
         n50611, n50612, n50613, n50614, n50615, n50616, n50617, n50618,
         n50619, n50620, n50621, n50622, n50623, n50624, n50625, n50626,
         n50627, n50628, n50629, n50630, n50631, n50632, n50633, n50634,
         n50635, n50636, n50637, n50638, n50639, n50640, n50641, n50642,
         n50643, n50644, n50645, n50646, n50647, n50648, n50649, n50650,
         n50651, n50652, n50653, n50654, n50655, n50656, n50657, n50658,
         n50659, n50660, n50661, n50662, n50663, n50664, n50665, n50666,
         n50667, n50668, n50669, n50670, n50671, n50672, n50673, n50674,
         n50675, n50676, n50677, n50678, n50679, n50680, n50681, n50682,
         n50683, n50684, n50685, n50686, n50687, n50688, n50689, n50690,
         n50691, n50692, n50693, n50694, n50695, n50696, n50697, n50698,
         n50699, n50700, n50701, n50702, n50703, n50704, n50705, n50706,
         n50707, n50708, n50709, n50710, n50711, n50712, n50713, n50714,
         n50715, n50716, n50717, n50718, n50719, n50720, n50721, n50722,
         n50723, n50724, n50725, n50726, n50727, n50728, n50729, n50730,
         n50731, n50732, n50733, n50734, n50735, n50736, n50737, n50738,
         n50739, n50740, n50741, n50742, n50743, n50744, n50745, n50746,
         n50747, n50748, n50749, n50750, n50751, n50752, n50753, n50754,
         n50755, n50756, n50757, n50758, n50759, n50760, n50761, n50762,
         n50763, n50764, n50765, n50766, n50767, n50768, n50769, n50770,
         n50771, n50772, n50773, n50774, n50775, n50776, n50777, n50778,
         n50779, n50780, n50781, n50782, n50783, n50784, n50785, n50786,
         n50787, n50788, n50789, n50790, n50791, n50792, n50793, n50794,
         n50795, n50796, n50797, n50798, n50799, n50800, n50801, n50802,
         n50803, n50804, n50805, n50806, n50807, n50808, n50809, n50810,
         n50811, n50812, n50813, n50814, n50815, n50816, n50817, n50818,
         n50819, n50820, n50821, n50822, n50823, n50824, n50825, n50826,
         n50827, n50828, n50829, n50830, n50831, n50832, n50833, n50834,
         n50835, n50836, n50837, n50838, n50839, n50840, n50841, n50842,
         n50843, n50844, n50845, n50846, n50847, n50848, n50849, n50850,
         n50851, n50852, n50853, n50854, n50855, n50856, n50857, n50858,
         n50859, n50860, n50861, n50862, n50863, n50864, n50865, n50866,
         n50867, n50868, n50869, n50870, n50871, n50872, n50873, n50874,
         n50875, n50876, n50877, n50878, n50879, n50880, n50881, n50882,
         n50883, n50884, n50885, n50886, n50887, n50888, n50889, n50890,
         n50891, n50892, n50893, n50894, n50895, n50896, n50897, n50898,
         n50899, n50900, n50901, n50902, n50903, n50904, n50905, n50906,
         n50907, n50908, n50909, n50910, n50911, n50912, n50913, n50914,
         n50915, n50916, n50917, n50918, n50919, n50920, n50921, n50922,
         n50923, n50924, n50925, n50926, n50927, n50928, n50929, n50930,
         n50931, n50932, n50933, n50934, n50935, n50936, n50937, n50938,
         n50939, n50940, n50941, n50942, n50943, n50944, n50945, n50946,
         n50947, n50948, n50949, n50950, n50951, n50952, n50953, n50954,
         n50955, n50956, n50957, n50958, n50959, n50960, n50961, n50962,
         n50963, n50964, n50965, n50966, n50967, n50968, n50969, n50970,
         n50971, n50972, n50973, n50974, n50975, n50976, n50977, n50978,
         n50979, n50980, n50981, n50982, n50983, n50984, n50985, n50986,
         n50987, n50988, n50989, n50990, n50991, n50992, n50993, n50994,
         n50995, n50996, n50997, n50998, n50999, n51000, n51001, n51002,
         n51003, n51004, n51005, n51006, n51007, n51008, n51009, n51010,
         n51011, n51012, n51013, n51014, n51015, n51016, n51017, n51018,
         n51019, n51020, n51021, n51022, n51023, n51024, n51025, n51026,
         n51027, n51028, n51029, n51030, n51031, n51032, n51033, n51034,
         n51035, n51036, n51037, n51038, n51039, n51040, n51041, n51042,
         n51043, n51044, n51045, n51046, n51047, n51048, n51049, n51050,
         n51051, n51052, n51053, n51054, n51055, n51056, n51057, n51058,
         n51059, n51060, n51061, n51062, n51063, n51064, n51065, n51066,
         n51067, n51068, n51069, n51070, n51071, n51072, n51073, n51074,
         n51075, n51076, n51077, n51078, n51079, n51080, n51081, n51082,
         n51083, n51084, n51085, n51086, n51087, n51088, n51089, n51090,
         n51091, n51092, n51093, n51094, n51095, n51096, n51097, n51098,
         n51099, n51100, n51101, n51102, n51103, n51104, n51105, n51106,
         n51107, n51108, n51109, n51110, n51111, n51112, n51113, n51114,
         n51115, n51116, n51117, n51118, n51119, n51120, n51121, n51122,
         n51123, n51124, n51125, n51126, n51127, n51128, n51129, n51130,
         n51131, n51132, n51133, n51134, n51135, n51136, n51137, n51138,
         n51139, n51140, n51141, n51142, n51143, n51144, n51145, n51146,
         n51147, n51148, n51149, n51150, n51151, n51152, n51153, n51154,
         n51155, n51156, n51157, n51158, n51159, n51160, n51161, n51162,
         n51163, n51164, n51165, n51166, n51167, n51168, n51169, n51170,
         n51171, n51172, n51173, n51174, n51175, n51176, n51177, n51178,
         n51179, n51180, n51181, n51182, n51183, n51184, n51185, n51186,
         n51187, n51188, n51189, n51190, n51191, n51192, n51193, n51194,
         n51195, n51196, n51197, n51198, n51199, n51200, n51201, n51202,
         n51203, n51204, n51205, n51206, n51207, n51208, n51209, n51210,
         n51211, n51212, n51213, n51214, n51215, n51216, n51217, n51218,
         n51219, n51220, n51221, n51222, n51223, n51224, n51225, n51226,
         n51227, n51228, n51229, n51230, n51231, n51232, n51233, n51234,
         n51235, n51236, n51237, n51238, n51239, n51240, n51241, n51242,
         n51243, n51244, n51245, n51246, n51247, n51248, n51249, n51250,
         n51251, n51252, n51253, n51254, n51255, n51256, n51257, n51258,
         n51259, n51260, n51261, n51262, n51263, n51264, n51265, n51266,
         n51267, n51268, n51269, n51270, n51271, n51272, n51273, n51274,
         n51275, n51276, n51277, n51278, n51279, n51280, n51281, n51282,
         n51283, n51284, n51285, n51286, n51287, n51288, n51289, n51290,
         n51291, n51292, n51293, n51294, n51295, n51296, n51297, n51298,
         n51299, n51300, n51301, n51302, n51303, n51304, n51305, n51306,
         n51307, n51308, n51309, n51310, n51311, n51312, n51313, n51314,
         n51315, n51316, n51317, n51318, n51319, n51320, n51321, n51322,
         n51323, n51324, n51325, n51326, n51327, n51328, n51329, n51330,
         n51331, n51332, n51333, n51334, n51335, n51336, n51337, n51338,
         n51339, n51340, n51341, n51342, n51343, n51344, n51345, n51346,
         n51347, n51348, n51349, n51350, n51351, n51352, n51353, n51354,
         n51355, n51356, n51357, n51358, n51359, n51360, n51361, n51362,
         n51363, n51364, n51365, n51366, n51367, n51368, n51369, n51370,
         n51371, n51372, n51373, n51374, n51375, n51376, n51377, n51378,
         n51379, n51380, n51381, n51382, n51383, n51384, n51385, n51386,
         n51387, n51388, n51389, n51390, n51391, n51392, n51393, n51394,
         n51395, n51396, n51397, n51398, n51399, n51400, n51401, n51402,
         n51403, n51404, n51405, n51406, n51407, n51408, n51409, n51410,
         n51411, n51412, n51413, n51414, n51415, n51416, n51417, n51418,
         n51419, n51420, n51421, n51422, n51423, n51424, n51425, n51426,
         n51427, n51428, n51429, n51430, n51431, n51432, n51433, n51434,
         n51435, n51436, n51437, n51438, n51439, n51440, n51441, n51442,
         n51443, n51444, n51445, n51446, n51447, n51448, n51449, n51450,
         n51451, n51452, n51453, n51454, n51455, n51456, n51457, n51458,
         n51459, n51460, n51461, n51462, n51463, n51464, n51465, n51466,
         n51467, n51468, n51469, n51470, n51471, n51472, n51473, n51474,
         n51475, n51476, n51477, n51478, n51479, n51480, n51481, n51482,
         n51483, n51484, n51485, n51486, n51487, n51488, n51489, n51490,
         n51491, n51492, n51493, n51494, n51495, n51496, n51497, n51498,
         n51499, n51500, n51501, n51502, n51503, n51504, n51505, n51506,
         n51507, n51508, n51509, n51510, n51511, n51512, n51513, n51514,
         n51515, n51516, n51517, n51518, n51519, n51520, n51521, n51522,
         n51523, n51524, n51525, n51526, n51527, n51528, n51529, n51530,
         n51531, n51532, n51533, n51534, n51535, n51536, n51537, n51538,
         n51539, n51540, n51541, n51542, n51543, n51544, n51545, n51546,
         n51547, n51548, n51549, n51550, n51551, n51552, n51553, n51554,
         n51555, n51556, n51557, n51558, n51559, n51560, n51561, n51562,
         n51563, n51564, n51565, n51566, n51567, n51568, n51569, n51570,
         n51571, n51572, n51573, n51574, n51575, n51576, n51577, n51578,
         n51579, n51580, n51581, n51582, n51583, n51584, n51585, n51586,
         n51587, n51588, n51589, n51590, n51591, n51592, n51593, n51594,
         n51595, n51596, n51597, n51598, n51599, n51600, n51601, n51602,
         n51603, n51604, n51605, n51606, n51607, n51608, n51609, n51610,
         n51611, n51612, n51613, n51614, n51615, n51616, n51617, n51618,
         n51619, n51620, n51621, n51622, n51623, n51624, n51625, n51626,
         n51627, n51628, n51629, n51630, n51631, n51632, n51633, n51634,
         n51635, n51636, n51637, n51638, n51639, n51640, n51641, n51642,
         n51643, n51644, n51645, n51646, n51647, n51648, n51649, n51650,
         n51651, n51652, n51653, n51654, n51655, n51656, n51657, n51658,
         n51659, n51660, n51661, n51662, n51663, n51664, n51665, n51666,
         n51667, n51668, n51669, n51670, n51671, n51672, n51673, n51674,
         n51675, n51676, n51677, n51678, n51679, n51680, n51681, n51682,
         n51683, n51684, n51685, n51686, n51687, n51688, n51689, n51690,
         n51691, n51692, n51693, n51694, n51695, n51696, n51697, n51698,
         n51699, n51700, n51701, n51702, n51703, n51704, n51705, n51706,
         n51707, n51708, n51709, n51710, n51711, n51712, n51713, n51714,
         n51715, n51716, n51717, n51718, n51719, n51720, n51721, n51722,
         n51723, n51724, n51725, n51726, n51727, n51728, n51729, n51730,
         n51731, n51732, n51733, n51734, n51735, n51736, n51737, n51738,
         n51739, n51740, n51741, n51742, n51743, n51744, n51745, n51746,
         n51747, n51748, n51749, n51750, n51751, n51752, n51753, n51754,
         n51755, n51756, n51757, n51758, n51759, n51760, n51761, n51762,
         n51763, n51764, n51765, n51766, n51767, n51768, n51769, n51770,
         n51771, n51772, n51773, n51774, n51775, n51776, n51777, n51778,
         n51779, n51780, n51781, n51782, n51783, n51784, n51785, n51786,
         n51787, n51788, n51789, n51790, n51791, n51792, n51793, n51794,
         n51795, n51796, n51797, n51798, n51799, n51800, n51801, n51802,
         n51803, n51804, n51805, n51806, n51807, n51808, n51809, n51810,
         n51811, n51812, n51813, n51814, n51815, n51816, n51817, n51818,
         n51819, n51820, n51821, n51822, n51823, n51824, n51825, n51826,
         n51827, n51828, n51829, n51830, n51831, n51832, n51833, n51834,
         n51835, n51836, n51837, n51838, n51839, n51840, n51841, n51842,
         n51843, n51844, n51845, n51846, n51847, n51848, n51849, n51850,
         n51851, n51852, n51853, n51854, n51855, n51856, n51857, n51858,
         n51859, n51860, n51861, n51862, n51863, n51864, n51865, n51866,
         n51867, n51868, n51869, n51870, n51871, n51872, n51873, n51874,
         n51875, n51876, n51877, n51878, n51879, n51880, n51881, n51882,
         n51883, n51884, n51885, n51886, n51887, n51888, n51889, n51890,
         n51891, n51892, n51893, n51894, n51895, n51896, n51897, n51898,
         n51899, n51900, n51901, n51902, n51903, n51904, n51905, n51906,
         n51907, n51908, n51909, n51910, n51911, n51912, n51913, n51914,
         n51915, n51916, n51917, n51918, n51919, n51920, n51921, n51922,
         n51923, n51924, n51925, n51926, n51927, n51928, n51929, n51930,
         n51931, n51932, n51933, n51934, n51935, n51936, n51937, n51938,
         n51939, n51940, n51941, n51942, n51943, n51944, n51945, n51946,
         n51947, n51948, n51949, n51950, n51951, n51952, n51953, n51954,
         n51955, n51956, n51957, n51958, n51959, n51960, n51961, n51962,
         n51963, n51964, n51965, n51966, n51967, n51968, n51969, n51970,
         n51971, n51972, n51973, n51974, n51975, n51976, n51977, n51978,
         n51979, n51980, n51981, n51982, n51983, n51984, n51985, n51986,
         n51987, n51988, n51989, n51990, n51991, n51992, n51993, n51994,
         n51995, n51996, n51997, n51998, n51999, n52000, n52001, n52002,
         n52003, n52004, n52005, n52006, n52007, n52008, n52009, n52010,
         n52011, n52012, n52013, n52014, n52015, n52016, n52017, n52018,
         n52019, n52020, n52021, n52022, n52023, n52024, n52025, n52026,
         n52027, n52028, n52029, n52030, n52031, n52032, n52033, n52034,
         n52035, n52036, n52037, n52038, n52039, n52040, n52041, n52042,
         n52043, n52044, n52045, n52046, n52047, n52048, n52049, n52050,
         n52051, n52052, n52053, n52054, n52055, n52056, n52057, n52058,
         n52059, n52060, n52061, n52062, n52063, n52064, n52065, n52066,
         n52067, n52068, n52069, n52070, n52071, n52072, n52073, n52074,
         n52075, n52076, n52077, n52078, n52079, n52080, n52081, n52082,
         n52083, n52084, n52085, n52086, n52087, n52088, n52089, n52090,
         n52091, n52092, n52093, n52094, n52095, n52096, n52097, n52098,
         n52099, n52100, n52101, n52102, n52103, n52104, n52105, n52106,
         n52107, n52108, n52109, n52110, n52111, n52112, n52113, n52114,
         n52115, n52116, n52117, n52118, n52119, n52120, n52121, n52122,
         n52123, n52124, n52125, n52126, n52127, n52128, n52129, n52130,
         n52131, n52132, n52133, n52134, n52135, n52136, n52137, n52138,
         n52139, n52140, n52141, n52142, n52143, n52144, n52145, n52146,
         n52147, n52148, n52149, n52150, n52151, n52152, n52153, n52154,
         n52155, n52156, n52157, n52158, n52159, n52160, n52161, n52162,
         n52163, n52164, n52165, n52166, n52167, n52168, n52169, n52170,
         n52171, n52172, n52173, n52174, n52175, n52176, n52177, n52178,
         n52179, n52180, n52181, n52182, n52183, n52184, n52185, n52186,
         n52187, n52188, n52189, n52190, n52191, n52192, n52193, n52194,
         n52195, n52196, n52197, n52198, n52199, n52200, n52201, n52202,
         n52203, n52204, n52205, n52206, n52207, n52208, n52209, n52210,
         n52211, n52212, n52213, n52214, n52215, n52216, n52217, n52218,
         n52219, n52220, n52221, n52222, n52223, n52224, n52225, n52226,
         n52227, n52228, n52229, n52230, n52231, n52232, n52233, n52234,
         n52235, n52236, n52237, n52238, n52239, n52240, n52241, n52242,
         n52243, n52244, n52245, n52246, n52247, n52248, n52249, n52250,
         n52251, n52252, n52253, n52254, n52255, n52256, n52257, n52258,
         n52259, n52260, n52261, n52262, n52263, n52264, n52265, n52266,
         n52267, n52268, n52269, n52270, n52271, n52272, n52273, n52274,
         n52275, n52276, n52277, n52278, n52279, n52280, n52281, n52282,
         n52283, n52284, n52285, n52286, n52287, n52288, n52289, n52290,
         n52291, n52292, n52293, n52294, n52295, n52296, n52297, n52298,
         n52299, n52300, n52301, n52302, n52303, n52304, n52305, n52306,
         n52307, n52308, n52309, n52310, n52311, n52312, n52313, n52314,
         n52315, n52316, n52317, n52318, n52319, n52320, n52321, n52322,
         n52323, n52324, n52325, n52326, n52327, n52328, n52329, n52330,
         n52331, n52332, n52333, n52334, n52335, n52336, n52337, n52338,
         n52339, n52340, n52341, n52342, n52343, n52344, n52345, n52346,
         n52347, n52348, n52349, n52350, n52351, n52352, n52353, n52354,
         n52355, n52356, n52357, n52358, n52359, n52360, n52361, n52362,
         n52363, n52364, n52365, n52366, n52367, n52368, n52369, n52370,
         n52371, n52372, n52373, n52374, n52375, n52376, n52377, n52378,
         n52379, n52380, n52381, n52382, n52383, n52384, n52385, n52386,
         n52387, n52388, n52389, n52390, n52391, n52392, n52393, n52394,
         n52395, n52396, n52397, n52398, n52399, n52400, n52401, n52402,
         n52403, n52404, n52405, n52406, n52407, n52408, n52409, n52410,
         n52411, n52412, n52413, n52414, n52415, n52416, n52417, n52418,
         n52419, n52420, n52421, n52422, n52423, n52424, n52425, n52426,
         n52427, n52428, n52429, n52430, n52431, n52432, n52433, n52434,
         n52435, n52436, n52437, n52438, n52439, n52440, n52441, n52442,
         n52443, n52444, n52445, n52446, n52447, n52448, n52449, n52450,
         n52451, n52452, n52453, n52454, n52455, n52456, n52457, n52458,
         n52459, n52460, n52461, n52462, n52463, n52464, n52465, n52466,
         n52467, n52468, n52469, n52470, n52471, n52472, n52473, n52474,
         n52475, n52476, n52477, n52478, n52479, n52480, n52481, n52482,
         n52483, n52484, n52485, n52486, n52487, n52488, n52489, n52490,
         n52491, n52492, n52493, n52494, n52495, n52496, n52497, n52498,
         n52499, n52500, n52501, n52502, n52503, n52504, n52505, n52506,
         n52507, n52508, n52509, n52510, n52511, n52512, n52513, n52514,
         n52515, n52516, n52517, n52518, n52519, n52520, n52521, n52522,
         n52523, n52524, n52525, n52526, n52527, n52528, n52529, n52530,
         n52531, n52532, n52533, n52534, n52535, n52536, n52537, n52538,
         n52539, n52540, n52541, n52542, n52543, n52544, n52545, n52546,
         n52547, n52548, n52549, n52550, n52551, n52552, n52553, n52554,
         n52555, n52556, n52557, n52558, n52559, n52560, n52561, n52562,
         n52563, n52564, n52565, n52566, n52567, n52568, n52569, n52570,
         n52571, n52572, n52573, n52574, n52575, n52576, n52577, n52578,
         n52579, n52580, n52581, n52582, n52583, n52584, n52585, n52586,
         n52587, n52588, n52589, n52590, n52591, n52592, n52593, n52594,
         n52595, n52596, n52597, n52598, n52599, n52600, n52601, n52602,
         n52603, n52604, n52605, n52606, n52607, n52608, n52609, n52610,
         n52611, n52612, n52613, n52614, n52615, n52616, n52617, n52618,
         n52619, n52620, n52621, n52622, n52623, n52624, n52625, n52626,
         n52627, n52628, n52629, n52630, n52631, n52632, n52633, n52634,
         n52635, n52636, n52637, n52638, n52639, n52640, n52641, n52642,
         n52643, n52644, n52645, n52646, n52647, n52648, n52649, n52650,
         n52651, n52652, n52653, n52654, n52655, n52656, n52657, n52658,
         n52659, n52660, n52661, n52662, n52663, n52664, n52665, n52666,
         n52667, n52668, n52669, n52670, n52671, n52672, n52673, n52674,
         n52675, n52676, n52677, n52678, n52679, n52680, n52681, n52682,
         n52683, n52684, n52685, n52686, n52687, n52688, n52689, n52690,
         n52691, n52692, n52693, n52694, n52695, n52696, n52697, n52698,
         n52699, n52700, n52701, n52702, n52703, n52704, n52705, n52706,
         n52707, n52708, n52709, n52710, n52711, n52712, n52713, n52714,
         n52715, n52716, n52717, n52718, n52719, n52720, n52721, n52722,
         n52723, n52724, n52725, n52726, n52727, n52728, n52729, n52730,
         n52731, n52732, n52733, n52734, n52735, n52736, n52737, n52738,
         n52739, n52740, n52741, n52742, n52743, n52744, n52745, n52746,
         n52747, n52748, n52749, n52750, n52751, n52752, n52753, n52754,
         n52755, n52756, n52757, n52758, n52759, n52760, n52761, n52762,
         n52763, n52764, n52765, n52766, n52767, n52768, n52769, n52770,
         n52771, n52772, n52773, n52774, n52775, n52776, n52777, n52778,
         n52779, n52780, n52781, n52782, n52783, n52784, n52785, n52786,
         n52787, n52788, n52789, n52790, n52791, n52792, n52793, n52794,
         n52795, n52796, n52797, n52798, n52799, n52800, n52801, n52802,
         n52803, n52804, n52805, n52806, n52807, n52808, n52809, n52810,
         n52811, n52812, n52813, n52814, n52815, n52816, n52817, n52818,
         n52819, n52820, n52821, n52822, n52823, n52824, n52825, n52826,
         n52827, n52828, n52829, n52830, n52831, n52832, n52833, n52834,
         n52835, n52836, n52837, n52838, n52839, n52840, n52841, n52842,
         n52843, n52844, n52845, n52846, n52847, n52848, n52849, n52850,
         n52851, n52852, n52853, n52854, n52855, n52856, n52857, n52858,
         n52859, n52860, n52861, n52862, n52863, n52864, n52865, n52866,
         n52867, n52868, n52869, n52870, n52871, n52872, n52873, n52874,
         n52875, n52876, n52877, n52878, n52879, n52880, n52881, n52882,
         n52883, n52884, n52885, n52886, n52887, n52888, n52889, n52890,
         n52891, n52892, n52893, n52894, n52895, n52896, n52897, n52898,
         n52899, n52900, n52901, n52902, n52903, n52904, n52905, n52906,
         n52907, n52908, n52909, n52910, n52911, n52912, n52913, n52914,
         n52915, n52916, n52917, n52918, n52919, n52920, n52921, n52922,
         n52923, n52924, n52925, n52926, n52927, n52928, n52929, n52930,
         n52931, n52932, n52933, n52934, n52935, n52936, n52937, n52938,
         n52939, n52940, n52941, n52942, n52943, n52944, n52945, n52946,
         n52947, n52948, n52949, n52950, n52951, n52952, n52953, n52954,
         n52955, n52956, n52957, n52958, n52959, n52960, n52961, n52962,
         n52963, n52964, n52965, n52966, n52967, n52968, n52969, n52970,
         n52971, n52972, n52973, n52974, n52975, n52976, n52977, n52978,
         n52979, n52980, n52981, n52982, n52983, n52984, n52985, n52986,
         n52987, n52988, n52989, n52990, n52991, n52992, n52993, n52994,
         n52995, n52996, n52997, n52998, n52999, n53000, n53001, n53002,
         n53003, n53004, n53005, n53006, n53007, n53008, n53009, n53010,
         n53011, n53012, n53013, n53014, n53015, n53016, n53017, n53018,
         n53019, n53020, n53021, n53022, n53023, n53024, n53025, n53026,
         n53027, n53028, n53029, n53030, n53031, n53032, n53033, n53034,
         n53035, n53036, n53037, n53038, n53039, n53040, n53041, n53042,
         n53043, n53044, n53045, n53046, n53047, n53048, n53049, n53050,
         n53051, n53052, n53053, n53054, n53055, n53056, n53057, n53058,
         n53059, n53060, n53061, n53062, n53063, n53064, n53065, n53066,
         n53067, n53068, n53069, n53070, n53071, n53072, n53073, n53074,
         n53075, n53076, n53077, n53078, n53079, n53080, n53081, n53082,
         n53083, n53084, n53085, n53086, n53087, n53088, n53089, n53090,
         n53091, n53092, n53093, n53094, n53095, n53096, n53097, n53098,
         n53099, n53100, n53101, n53102, n53103, n53104, n53105, n53106,
         n53107, n53108, n53109, n53110, n53111, n53112, n53113, n53114,
         n53115, n53116, n53117, n53118, n53119, n53120, n53121, n53122,
         n53123, n53124, n53125, n53126, n53127, n53128, n53129, n53130,
         n53131, n53132, n53133, n53134, n53135, n53136, n53137, n53138,
         n53139, n53140, n53141, n53142, n53143, n53144, n53145, n53146,
         n53147, n53148, n53149, n53150, n53151, n53152, n53153, n53154,
         n53155, n53156, n53157, n53158, n53159, n53160, n53161, n53162,
         n53163, n53164, n53165, n53166, n53167, n53168, n53169, n53170,
         n53171, n53172, n53173, n53174, n53175, n53176, n53177, n53178,
         n53179, n53180, n53181, n53182, n53183, n53184, n53185, n53186,
         n53187, n53188, n53189, n53190, n53191, n53192, n53193, n53194,
         n53195, n53196, n53197, n53198, n53199, n53200, n53201, n53202,
         n53203, n53204, n53205, n53206, n53207, n53208, n53209, n53210,
         n53211, n53212, n53213, n53214, n53215, n53216, n53217, n53218,
         n53219, n53220, n53221, n53222, n53223, n53224, n53225, n53226,
         n53227, n53228, n53229, n53230, n53231, n53232, n53233, n53234,
         n53235, n53236, n53237, n53238, n53239, n53240, n53241, n53242,
         n53243, n53244, n53245, n53246, n53247, n53248, n53249, n53250,
         n53251, n53252, n53253, n53254, n53255, n53256, n53257, n53258,
         n53259, n53260, n53261, n53262, n53263, n53264, n53265, n53266,
         n53267, n53268, n53269, n53270, n53271, n53272, n53273, n53274,
         n53275, n53276, n53277, n53278, n53279, n53280, n53281, n53282,
         n53283, n53284, n53285, n53286, n53287, n53288, n53289, n53290,
         n53291, n53292, n53293, n53294, n53295, n53296, n53297, n53298,
         n53299, n53300, n53301, n53302, n53303, n53304, n53305, n53306,
         n53307, n53308, n53309, n53310, n53311, n53312, n53313, n53314,
         n53315, n53316, n53317, n53318, n53319, n53320, n53321, n53322,
         n53323, n53324, n53325, n53326, n53327, n53328, n53329, n53330,
         n53331, n53332, n53333, n53334, n53335, n53336, n53337, n53338,
         n53339, n53340, n53341, n53342, n53343, n53344, n53345, n53346,
         n53347, n53348, n53349, n53350, n53351, n53352, n53353, n53354,
         n53355, n53356, n53357, n53358, n53359, n53360, n53361, n53362,
         n53363, n53364, n53365, n53366, n53367, n53368, n53369, n53370,
         n53371, n53372, n53373, n53374, n53375, n53376, n53377, n53378,
         n53379, n53380, n53381, n53382, n53383, n53384, n53385, n53386,
         n53387, n53388, n53389, n53390, n53391, n53392, n53393, n53394,
         n53395, n53396, n53397, n53398, n53399, n53400, n53401, n53402,
         n53403, n53404, n53405, n53406, n53407, n53408, n53409, n53410,
         n53411, n53412, n53413, n53414, n53415, n53416, n53417, n53418,
         n53419, n53420, n53421, n53422, n53423, n53424, n53425, n53426,
         n53427, n53428, n53429, n53430, n53431, n53432, n53433, n53434,
         n53435, n53436, n53437, n53438, n53439, n53440, n53441, n53442,
         n53443, n53444, n53445, n53446, n53447, n53448, n53449, n53450,
         n53451, n53452, n53453, n53454, n53455, n53456, n53457, n53458,
         n53459, n53460, n53461, n53462, n53463, n53464, n53465, n53466,
         n53467, n53468, n53469, n53470, n53471, n53472, n53473, n53474,
         n53475, n53476, n53477, n53478, n53479, n53480, n53481, n53482,
         n53483, n53484, n53485, n53486, n53487, n53488, n53489, n53490,
         n53491, n53492, n53493, n53494, n53495, n53496, n53497, n53498,
         n53499, n53500, n53501, n53502, n53503, n53504, n53505, n53506,
         n53507, n53508, n53509, n53510, n53511, n53512, n53513, n53514,
         n53515, n53516, n53517, n53518, n53519, n53520, n53521, n53522,
         n53523, n53524, n53525, n53526, n53527, n53528, n53529, n53530,
         n53531, n53532, n53533, n53534, n53535, n53536, n53537, n53538,
         n53539, n53540, n53541, n53542, n53543, n53544, n53545, n53546,
         n53547, n53548, n53549, n53550, n53551, n53552, n53553, n53554,
         n53555, n53556, n53557, n53558, n53559, n53560, n53561, n53562,
         n53563, n53564, n53565, n53566, n53567, n53568, n53569, n53570,
         n53571, n53572, n53573, n53574, n53575, n53576, n53577, n53578,
         n53579, n53580, n53581, n53582, n53583, n53584, n53585, n53586,
         n53587, n53588, n53589, n53590, n53591, n53592, n53593, n53594,
         n53595, n53596, n53597, n53598, n53599, n53600, n53601, n53602,
         n53603, n53604, n53605, n53606, n53607, n53608, n53609, n53610,
         n53611, n53612, n53613, n53614, n53615, n53616, n53617, n53618,
         n53619, n53620, n53621, n53622, n53623, n53624, n53625, n53626,
         n53627, n53628, n53629, n53630, n53631, n53632, n53633, n53634,
         n53635, n53636, n53637, n53638, n53639, n53640, n53641, n53642,
         n53643, n53644, n53645, n53646, n53647, n53648, n53649, n53650,
         n53651, n53652, n53653, n53654, n53655, n53656, n53657, n53658,
         n53659, n53660, n53661, n53662, n53663, n53664, n53665, n53666,
         n53667, n53668, n53669, n53670, n53671, n53672, n53673, n53674,
         n53675, n53676, n53677, n53678, n53679, n53680, n53681, n53682,
         n53683, n53684, n53685, n53686, n53687, n53688, n53689, n53690,
         n53691, n53692, n53693, n53694, n53695, n53696, n53697, n53698,
         n53699, n53700, n53701, n53702, n53703, n53704, n53705, n53706,
         n53707, n53708, n53709, n53710, n53711, n53712, n53713, n53714,
         n53715, n53716, n53717, n53718, n53719, n53720, n53721, n53722,
         n53723, n53724, n53725, n53726, n53727, n53728, n53729, n53730,
         n53731, n53732, n53733, n53734, n53735, n53736, n53737, n53738,
         n53739, n53740, n53741, n53742, n53743, n53744, n53745, n53746,
         n53747, n53748, n53749, n53750, n53751, n53752, n53753, n53754,
         n53755, n53756, n53757, n53758, n53759, n53760, n53761, n53762,
         n53763, n53764, n53765, n53766, n53767, n53768, n53769, n53770,
         n53771, n53772, n53773, n53774, n53775, n53776, n53777, n53778,
         n53779, n53780, n53781, n53782, n53783, n53784, n53785, n53786,
         n53787, n53788, n53789, n53790, n53791, n53792, n53793, n53794,
         n53795, n53796, n53797, n53798, n53799, n53800, n53801, n53802,
         n53803, n53804, n53805, n53806, n53807, n53808, n53809, n53810,
         n53811, n53812, n53813, n53814, n53815, n53816, n53817, n53818,
         n53819, n53820, n53821, n53822, n53823, n53824, n53825, n53826,
         n53827, n53828, n53829, n53830, n53831, n53832, n53833, n53834,
         n53835, n53836, n53837, n53838, n53839, n53840, n53841, n53842,
         n53843, n53844, n53845, n53846, n53847, n53848, n53849, n53850,
         n53851, n53852, n53853, n53854, n53855, n53856, n53857, n53858,
         n53859, n53860, n53861, n53862, n53863, n53864, n53865, n53866,
         n53867, n53868, n53869, n53870, n53871, n53872, n53873, n53874,
         n53875, n53876, n53877, n53878, n53879, n53880, n53881, n53882,
         n53883, n53884, n53885, n53886, n53887, n53888, n53889, n53890,
         n53891, n53892, n53893, n53894, n53895, n53896, n53897, n53898,
         n53899, n53900, n53901, n53902, n53903, n53904, n53905, n53906,
         n53907, n53908, n53909, n53910, n53911, n53912, n53913, n53914,
         n53915, n53916, n53917, n53918, n53919, n53920, n53921, n53922,
         n53923, n53924, n53925, n53926, n53927, n53928, n53929, n53930,
         n53931, n53932, n53933, n53934, n53935, n53936, n53937, n53938,
         n53939, n53940, n53941, n53942, n53943, n53944, n53945, n53946,
         n53947, n53948, n53949, n53950, n53951, n53952, n53953, n53954,
         n53955, n53956, n53957, n53958, n53959, n53960, n53961, n53962,
         n53963, n53964, n53965, n53966, n53967, n53968, n53969, n53970,
         n53971, n53972, n53973, n53974, n53975, n53976, n53977, n53978,
         n53979, n53980, n53981, n53982, n53983, n53984, n53985, n53986,
         n53987, n53988, n53989, n53990, n53991, n53992, n53993, n53994,
         n53995, n53996, n53997, n53998, n53999, n54000, n54001, n54002,
         n54003, n54004, n54005, n54006, n54007, n54008, n54009, n54010,
         n54011, n54012, n54013, n54014, n54015, n54016, n54017, n54018,
         n54019, n54020, n54021, n54022, n54023, n54024, n54025, n54026,
         n54027, n54028, n54029, n54030, n54031, n54032, n54033, n54034,
         n54035, n54036, n54037, n54038, n54039, n54040, n54041, n54042,
         n54043, n54044, n54045, n54046, n54047, n54048, n54049, n54050,
         n54051, n54052, n54053, n54054, n54055, n54056, n54057, n54058,
         n54059, n54060, n54061, n54062, n54063, n54064, n54065, n54066,
         n54067, n54068, n54069, n54070, n54071, n54072, n54073, n54074,
         n54075, n54076, n54077, n54078, n54079, n54080, n54081, n54082,
         n54083, n54084, n54085, n54086, n54087, n54088, n54089, n54090,
         n54091, n54092, n54093, n54094, n54095, n54096, n54097, n54098,
         n54099, n54100, n54101, n54102, n54103, n54104, n54105, n54106,
         n54107, n54108, n54109, n54110, n54111, n54112, n54113, n54114,
         n54115, n54116, n54117, n54118, n54119, n54120, n54121, n54122,
         n54123, n54124, n54125, n54126, n54127, n54128, n54129, n54130,
         n54131, n54132, n54133, n54134, n54135, n54136, n54137, n54138,
         n54139, n54140, n54141, n54142, n54143, n54144, n54145, n54146,
         n54147, n54148, n54149, n54150, n54151, n54152, n54153, n54154,
         n54155, n54156, n54157, n54158, n54159, n54160, n54161, n54162,
         n54163, n54164, n54165, n54166, n54167, n54168, n54169, n54170,
         n54171, n54172, n54173, n54174, n54175, n54176, n54177, n54178,
         n54179, n54180, n54181, n54182, n54183, n54184, n54185, n54186,
         n54187, n54188, n54189, n54190, n54191, n54192, n54193, n54194,
         n54195, n54196, n54197, n54198, n54199, n54200, n54201, n54202,
         n54203, n54204, n54205, n54206, n54207, n54208, n54209, n54210,
         n54211, n54212, n54213, n54214, n54215, n54216, n54217, n54218,
         n54219, n54220, n54221, n54222, n54223, n54224, n54225, n54226,
         n54227, n54228, n54229, n54230, n54231, n54232, n54233, n54234,
         n54235, n54236, n54237, n54238, n54239, n54240, n54241, n54242,
         n54243, n54244, n54245, n54246, n54247, n54248, n54249, n54250,
         n54251, n54252, n54253, n54254, n54255, n54256, n54257, n54258,
         n54259, n54260, n54261, n54262, n54263, n54264, n54265, n54266,
         n54267, n54268, n54269, n54270, n54271, n54272, n54273, n54274,
         n54275, n54276, n54277, n54278, n54279, n54280, n54281, n54282,
         n54283, n54284, n54285, n54286, n54287, n54288, n54289, n54290,
         n54291, n54292, n54293, n54294, n54295, n54296, n54297, n54298,
         n54299, n54300, n54301, n54302, n54303, n54304, n54305, n54306,
         n54307, n54308, n54309, n54310, n54311, n54312, n54313, n54314,
         n54315, n54316, n54317, n54318, n54319, n54320, n54321, n54322,
         n54323, n54324, n54325, n54326, n54327, n54328, n54329, n54330,
         n54331, n54332, n54333, n54334, n54335, n54336, n54337, n54338,
         n54339, n54340, n54341, n54342, n54343, n54344, n54345, n54346,
         n54347, n54348, n54349, n54350, n54351, n54352, n54353, n54354,
         n54355, n54356, n54357, n54358, n54359, n54360, n54361, n54362,
         n54363, n54364, n54365, n54366, n54367, n54368, n54369, n54370,
         n54371, n54372, n54373, n54374, n54375, n54376, n54377, n54378,
         n54379, n54380, n54381, n54382, n54383, n54384, n54385, n54386,
         n54387, n54388, n54389, n54390, n54391, n54392, n54393, n54394,
         n54395, n54396, n54397, n54398, n54399, n54400, n54401, n54402,
         n54403, n54404, n54405, n54406, n54407, n54408, n54409, n54410,
         n54411, n54412, n54413, n54414, n54415, n54416, n54417, n54418,
         n54419, n54420, n54421, n54422, n54423, n54424, n54425, n54426,
         n54427, n54428, n54429, n54430, n54431, n54432, n54433, n54434,
         n54435, n54436, n54437, n54438, n54439, n54440, n54441, n54442,
         n54443, n54444, n54445, n54446, n54447, n54448, n54449, n54450,
         n54451, n54452, n54453, n54454, n54455, n54456, n54457, n54458,
         n54459, n54460, n54461, n54462, n54463, n54464, n54465, n54466,
         n54467, n54468, n54469, n54470, n54471, n54472, n54473, n54474,
         n54475, n54476, n54477, n54478, n54479, n54480, n54481, n54482,
         n54483, n54484, n54485, n54486, n54487, n54488, n54489, n54490,
         n54491, n54492, n54493, n54494, n54495, n54496, n54497, n54498,
         n54499, n54500, n54501, n54502, n54503, n54504, n54505, n54506,
         n54507, n54508, n54509, n54510, n54511, n54512, n54513, n54514,
         n54515, n54516, n54517, n54518, n54519, n54520, n54521, n54522,
         n54523, n54524, n54525, n54526, n54527, n54528, n54529, n54530,
         n54531, n54532, n54533, n54534, n54535, n54536, n54537, n54538,
         n54539, n54540, n54541, n54542, n54543, n54544, n54545, n54546,
         n54547, n54548, n54549, n54550, n54551, n54552, n54553, n54554,
         n54555, n54556, n54557, n54558, n54559, n54560, n54561, n54562,
         n54563, n54564, n54565, n54566, n54567, n54568, n54569, n54570,
         n54571, n54572, n54573, n54574, n54575, n54576, n54577, n54578,
         n54579, n54580, n54581, n54582, n54583, n54584, n54585, n54586,
         n54587, n54588, n54589, n54590, n54591, n54592, n54593, n54594,
         n54595, n54596, n54597, n54598, n54599, n54600, n54601, n54602,
         n54603, n54604, n54605, n54606, n54607, n54608, n54609, n54610,
         n54611, n54612, n54613, n54614, n54615, n54616, n54617, n54618,
         n54619, n54620, n54621, n54622, n54623, n54624, n54625, n54626,
         n54627, n54628, n54629, n54630, n54631, n54632, n54633, n54634,
         n54635, n54636, n54637, n54638, n54639, n54640, n54641, n54642,
         n54643, n54644, n54645, n54646, n54647, n54648, n54649, n54650,
         n54651, n54652, n54653, n54654, n54655, n54656, n54657, n54658,
         n54659, n54660, n54661, n54662, n54663, n54664, n54665, n54666,
         n54667, n54668, n54669, n54670, n54671, n54672, n54673, n54674,
         n54675, n54676, n54677, n54678, n54679, n54680, n54681, n54682,
         n54683, n54684, n54685, n54686, n54687, n54688, n54689, n54690,
         n54691, n54692, n54693, n54694, n54695, n54696, n54697, n54698,
         n54699, n54700, n54701, n54702, n54703, n54704, n54705, n54706,
         n54707, n54708, n54709, n54710, n54711, n54712, n54713, n54714,
         n54715, n54716, n54717, n54718, n54719, n54720, n54721, n54722,
         n54723, n54724, n54725, n54726, n54727, n54728, n54729, n54730,
         n54731, n54732, n54733, n54734, n54735, n54736, n54737, n54738,
         n54739, n54740, n54741, n54742, n54743, n54744, n54745, n54746,
         n54747, n54748, n54749, n54750, n54751, n54752, n54753, n54754,
         n54755, n54756, n54757, n54758, n54759, n54760, n54761, n54762,
         n54763, n54764, n54765, n54766, n54767, n54768, n54769, n54770,
         n54771, n54772, n54773, n54774, n54775, n54776, n54777, n54778,
         n54779, n54780, n54781, n54782, n54783, n54784, n54785, n54786,
         n54787, n54788, n54789, n54790, n54791, n54792, n54793, n54794,
         n54795, n54796, n54797, n54798, n54799, n54800, n54801, n54802,
         n54803, n54804, n54805, n54806, n54807, n54808, n54809, n54810,
         n54811, n54812, n54813, n54814, n54815, n54816, n54817, n54818,
         n54819, n54820, n54821, n54822, n54823, n54824, n54825, n54826,
         n54827, n54828, n54829, n54830, n54831, n54832, n54833, n54834,
         n54835, n54836, n54837, n54838, n54839, n54840, n54841, n54842,
         n54843, n54844, n54845, n54846, n54847, n54848, n54849, n54850,
         n54851, n54852, n54853, n54854, n54855, n54856, n54857, n54858,
         n54859, n54860, n54861, n54862, n54863, n54864, n54865, n54866,
         n54867, n54868, n54869, n54870, n54871, n54872, n54873, n54874,
         n54875, n54876, n54877, n54878, n54879, n54880, n54881, n54882,
         n54883, n54884, n54885, n54886, n54887, n54888, n54889, n54890,
         n54891, n54892, n54893, n54894, n54895, n54896, n54897, n54898,
         n54899, n54900, n54901, n54902, n54903, n54904, n54905, n54906,
         n54907, n54908, n54909, n54910, n54911, n54912, n54913, n54914,
         n54915, n54916, n54917, n54918, n54919, n54920, n54921, n54922,
         n54923, n54924, n54925, n54926, n54927, n54928, n54929, n54930,
         n54931, n54932, n54933, n54934, n54935, n54936, n54937, n54938,
         n54939, n54940, n54941, n54942, n54943, n54944, n54945, n54946,
         n54947, n54948, n54949, n54950, n54951, n54952, n54953, n54954,
         n54955, n54956, n54957, n54958, n54959, n54960, n54961, n54962,
         n54963, n54964, n54965, n54966, n54967, n54968, n54969, n54970,
         n54971, n54972, n54973, n54974, n54975, n54976, n54977, n54978,
         n54979, n54980, n54981, n54982, n54983, n54984, n54985, n54986,
         n54987, n54988, n54989, n54990, n54991, n54992, n54993, n54994,
         n54995, n54996, n54997, n54998, n54999, n55000, n55001, n55002,
         n55003, n55004, n55005, n55006, n55007, n55008, n55009, n55010,
         n55011, n55012, n55013, n55014, n55015, n55016, n55017, n55018,
         n55019, n55020, n55021, n55022, n55023, n55024, n55025, n55026,
         n55027, n55028, n55029, n55030, n55031, n55032, n55033, n55034,
         n55035, n55036, n55037, n55038, n55039, n55040, n55041, n55042,
         n55043, n55044, n55045, n55046, n55047, n55048, n55049, n55050,
         n55051, n55052, n55053, n55054, n55055, n55056, n55057, n55058,
         n55059, n55060, n55061, n55062, n55063, n55064, n55065, n55066,
         n55067, n55068, n55069, n55070, n55071, n55072, n55073, n55074,
         n55075, n55076, n55077, n55078, n55079, n55080, n55081, n55082,
         n55083, n55084, n55085, n55086, n55087, n55088, n55089, n55090,
         n55091, n55092, n55093, n55094, n55095, n55096, n55097, n55098,
         n55099, n55100, n55101, n55102, n55103, n55104, n55105, n55106,
         n55107, n55108, n55109, n55110, n55111, n55112, n55113, n55114,
         n55115, n55116, n55117, n55118, n55119, n55120, n55121, n55122,
         n55123, n55124, n55125, n55126, n55127, n55128, n55129, n55130,
         n55131, n55132, n55133, n55134, n55135, n55136, n55137, n55138,
         n55139, n55140, n55141, n55142, n55143, n55144, n55145, n55146,
         n55147, n55148, n55149, n55150, n55151, n55152, n55153, n55154,
         n55155, n55156, n55157, n55158, n55159, n55160, n55161, n55162,
         n55163, n55164, n55165, n55166, n55167, n55168, n55169, n55170,
         n55171, n55172, n55173, n55174, n55175, n55176, n55177, n55178,
         n55179, n55180, n55181, n55182, n55183, n55184, n55185, n55186,
         n55187, n55188, n55189, n55190, n55191, n55192, n55193, n55194,
         n55195, n55196, n55197, n55198, n55199, n55200, n55201, n55202,
         n55203, n55204, n55205, n55206, n55207, n55208, n55209, n55210,
         n55211, n55212, n55213, n55214, n55215, n55216, n55217, n55218,
         n55219, n55220, n55221, n55222, n55223, n55224, n55225, n55226,
         n55227, n55228, n55229, n55230, n55231, n55232, n55233, n55234,
         n55235, n55236, n55237, n55238, n55239, n55240, n55241, n55242,
         n55243, n55244, n55245, n55246, n55247, n55248, n55249, n55250,
         n55251, n55252, n55253, n55254, n55255, n55256, n55257, n55258,
         n55259, n55260, n55261, n55262, n55263, n55264, n55265, n55266,
         n55267, n55268, n55269, n55270, n55271, n55272, n55273, n55274,
         n55275, n55276, n55277, n55278, n55279, n55280, n55281, n55282,
         n55283, n55284, n55285, n55286, n55287, n55288, n55289, n55290,
         n55291, n55292, n55293, n55294, n55295, n55296, n55297, n55298,
         n55299, n55300, n55301, n55302, n55303, n55304, n55305, n55306,
         n55307, n55308, n55309, n55310, n55311, n55312, n55313, n55314,
         n55315, n55316, n55317, n55318, n55319, n55320, n55321, n55322,
         n55323, n55324, n55325, n55326, n55327, n55328, n55329, n55330,
         n55331, n55332, n55333, n55334, n55335, n55336, n55337, n55338,
         n55339, n55340, n55341, n55342, n55343, n55344, n55345, n55346,
         n55347, n55348, n55349, n55350, n55351, n55352, n55353, n55354,
         n55355, n55356, n55357, n55358, n55359, n55360, n55361, n55362,
         n55363, n55364, n55365, n55366, n55367, n55368, n55369, n55370,
         n55371, n55372, n55373, n55374, n55375, n55376, n55377, n55378,
         n55379, n55380, n55381, n55382, n55383, n55384, n55385, n55386,
         n55387, n55388, n55389, n55390, n55391, n55392, n55393, n55394,
         n55395, n55396, n55397, n55398, n55399, n55400, n55401, n55402,
         n55403, n55404, n55405, n55406, n55407, n55408, n55409, n55410,
         n55411, n55412, n55413, n55414, n55415, n55416, n55417, n55418,
         n55419, n55420, n55421, n55422, n55423, n55424, n55425, n55426,
         n55427, n55428, n55429, n55430, n55431, n55432, n55433, n55434,
         n55435, n55436, n55437, n55438, n55439, n55440, n55441, n55442,
         n55443, n55444, n55445, n55446, n55447, n55448, n55449, n55450,
         n55451, n55452, n55453, n55454, n55455, n55456, n55457, n55458,
         n55459, n55460, n55461, n55462, n55463, n55464, n55465, n55466,
         n55467, n55468, n55469, n55470, n55471, n55472, n55473, n55474,
         n55475, n55476, n55477, n55478, n55479, n55480, n55481, n55482,
         n55483, n55484, n55485, n55486, n55487, n55488, n55489, n55490,
         n55491, n55492, n55493, n55494, n55495, n55496, n55497, n55498,
         n55499, n55500, n55501, n55502, n55503, n55504, n55505, n55506,
         n55507, n55508, n55509, n55510, n55511, n55512, n55513, n55514,
         n55515, n55516, n55517, n55518, n55519, n55520, n55521, n55522,
         n55523, n55524, n55525, n55526, n55527, n55528, n55529, n55530,
         n55531, n55532, n55533, n55534, n55535, n55536, n55537, n55538,
         n55539, n55540, n55541, n55542, n55543, n55544, n55545, n55546,
         n55547, n55548, n55549, n55550, n55551, n55552, n55553, n55554,
         n55555, n55556, n55557, n55558, n55559, n55560, n55561, n55562,
         n55563, n55564, n55565, n55566, n55567, n55568, n55569, n55570,
         n55571, n55572, n55573, n55574, n55575, n55576, n55577, n55578,
         n55579, n55580, n55581, n55582, n55583, n55584, n55585, n55586,
         n55587, n55588, n55589, n55590, n55591, n55592, n55593, n55594,
         n55595, n55596, n55597, n55598, n55599, n55600, n55601, n55602,
         n55603, n55604, n55605, n55606, n55607, n55608, n55609, n55610,
         n55611, n55612, n55613, n55614, n55615, n55616, n55617, n55618,
         n55619, n55620, n55621, n55622, n55623, n55624, n55625, n55626,
         n55627, n55628, n55629, n55630, n55631, n55632, n55633, n55634,
         n55635, n55636, n55637, n55638, n55639, n55640, n55641, n55642,
         n55643, n55644, n55645, n55646, n55647, n55648, n55649, n55650,
         n55651, n55652, n55653, n55654, n55655, n55656, n55657, n55658,
         n55659, n55660, n55661, n55662, n55663, n55664, n55665, n55666,
         n55667, n55668, n55669, n55670, n55671, n55672, n55673, n55674,
         n55675, n55676, n55677, n55678, n55679, n55680, n55681, n55682,
         n55683, n55684, n55685, n55686, n55687, n55688, n55689, n55690,
         n55691, n55692, n55693, n55694, n55695, n55696, n55697, n55698,
         n55699, n55700, n55701, n55702, n55703, n55704, n55705, n55706,
         n55707, n55708, n55709, n55710, n55711, n55712, n55713, n55714,
         n55715, n55716, n55717, n55718, n55719, n55720, n55721, n55722,
         n55723, n55724, n55725, n55726, n55727, n55728, n55729, n55730,
         n55731, n55732, n55733, n55734, n55735, n55736, n55737, n55738,
         n55739, n55740, n55741, n55742, n55743, n55744, n55745, n55746,
         n55747, n55748, n55749, n55750, n55751, n55752, n55753, n55754,
         n55755, n55756, n55757, n55758, n55759, n55760, n55761, n55762,
         n55763, n55764, n55765, n55766, n55767, n55768, n55769, n55770,
         n55771, n55772, n55773, n55774, n55775, n55776, n55777, n55778,
         n55779, n55780, n55781, n55782, n55783, n55784, n55785, n55786,
         n55787, n55788, n55789, n55790, n55791, n55792, n55793, n55794,
         n55795, n55796, n55797, n55798, n55799, n55800, n55801, n55802,
         n55803, n55804, n55805, n55806, n55807, n55808, n55809, n55810,
         n55811, n55812, n55813, n55814, n55815, n55816, n55817, n55818,
         n55819, n55820, n55821, n55822, n55823, n55824, n55825, n55826,
         n55827, n55828, n55829, n55830, n55831, n55832, n55833, n55834,
         n55835, n55836, n55837, n55838, n55839, n55840, n55841, n55842,
         n55843, n55844, n55845, n55846, n55847, n55848, n55849, n55850,
         n55851, n55852, n55853, n55854, n55855, n55856, n55857, n55858,
         n55859, n55860, n55861, n55862, n55863, n55864, n55865, n55866,
         n55867, n55868, n55869, n55870, n55871, n55872, n55873, n55874,
         n55875, n55876, n55877, n55878, n55879, n55880, n55881, n55882,
         n55883, n55884, n55885, n55886, n55887, n55888, n55889, n55890,
         n55891, n55892, n55893, n55894, n55895, n55896, n55897, n55898,
         n55899, n55900, n55901, n55902, n55903, n55904, n55905, n55906,
         n55907, n55908, n55909, n55910, n55911, n55912, n55913, n55914,
         n55915, n55916, n55917, n55918, n55919, n55920, n55921, n55922,
         n55923, n55924, n55925, n55926, n55927, n55928, n55929, n55930,
         n55931, n55932, n55933, n55934, n55935, n55936, n55937, n55938,
         n55939, n55940, n55941, n55942, n55943, n55944, n55945, n55946,
         n55947, n55948, n55949, n55950, n55951, n55952, n55953, n55954,
         n55955, n55956, n55957, n55958, n55959, n55960, n55961, n55962,
         n55963, n55964, n55965, n55966, n55967, n55968, n55969, n55970,
         n55971, n55972, n55973, n55974, n55975, n55976, n55977, n55978,
         n55979, n55980, n55981, n55982, n55983, n55984, n55985, n55986,
         n55987, n55988, n55989, n55990, n55991, n55992, n55993, n55994,
         n55995, n55996, n55997, n55998, n55999, n56000, n56001, n56002,
         n56003, n56004, n56005, n56006, n56007, n56008, n56009, n56010,
         n56011, n56012, n56013, n56014, n56015, n56016, n56017, n56018,
         n56019, n56020, n56021, n56022, n56023, n56024, n56025, n56026,
         n56027, n56028, n56029, n56030, n56031, n56032, n56033, n56034,
         n56035, n56036, n56037, n56038, n56039, n56040, n56041, n56042,
         n56043, n56044, n56045, n56046, n56047, n56048, n56049, n56050,
         n56051, n56052, n56053, n56054, n56055, n56056, n56057, n56058,
         n56059, n56060, n56061, n56062, n56063, n56064, n56065, n56066,
         n56067, n56068, n56069, n56070, n56071, n56072, n56073, n56074,
         n56075, n56076, n56077, n56078, n56079, n56080, n56081, n56082,
         n56083, n56084, n56085, n56086, n56087, n56088, n56089, n56090,
         n56091, n56092, n56093, n56094, n56095, n56096, n56097, n56098,
         n56099, n56100, n56101, n56102, n56103, n56104, n56105, n56106,
         n56107, n56108, n56109, n56110, n56111, n56112, n56113, n56114,
         n56115, n56116, n56117, n56118, n56119, n56120, n56121, n56122,
         n56123, n56124, n56125, n56126, n56127, n56128, n56129, n56130,
         n56131, n56132, n56133, n56134, n56135, n56136, n56137, n56138,
         n56139, n56140, n56141, n56142, n56143, n56144, n56145, n56146,
         n56147, n56148, n56149, n56150, n56151, n56152, n56153, n56154,
         n56155, n56156, n56157, n56158, n56159, n56160, n56161, n56162,
         n56163, n56164, n56165, n56166, n56167, n56168, n56169, n56170,
         n56171, n56172, n56173, n56174, n56175, n56176, n56177, n56178,
         n56179, n56180, n56181, n56182, n56183, n56184, n56185, n56186,
         n56187, n56188, n56189, n56190, n56191, n56192, n56193, n56194,
         n56195, n56196, n56197, n56198, n56199, n56200, n56201, n56202,
         n56203, n56204, n56205, n56206, n56207, n56208, n56209, n56210,
         n56211, n56212, n56213, n56214, n56215, n56216, n56217, n56218,
         n56219, n56220, n56221, n56222, n56223, n56224, n56225, n56226,
         n56227, n56228, n56229, n56230, n56231, n56232, n56233, n56234,
         n56235, n56236, n56237, n56238, n56239, n56240, n56241, n56242,
         n56243, n56244, n56245, n56246, n56247, n56248, n56249, n56250,
         n56251, n56252, n56253, n56254, n56255, n56256, n56257, n56258,
         n56259, n56260, n56261, n56262, n56263, n56264, n56265, n56266,
         n56267, n56268, n56269, n56270, n56271, n56272, n56273, n56274,
         n56275, n56276, n56277, n56278, n56279, n56280, n56281, n56282,
         n56283, n56284, n56285, n56286, n56287, n56288, n56289, n56290,
         n56291, n56292, n56293, n56294, n56295, n56296, n56297, n56298,
         n56299, n56300, n56301, n56302, n56303, n56304, n56305, n56306,
         n56307, n56308, n56309, n56310, n56311, n56312, n56313, n56314,
         n56315, n56316, n56317, n56318, n56319, n56320, n56321, n56322,
         n56323, n56324, n56325, n56326, n56327, n56328, n56329, n56330,
         n56331, n56332, n56333, n56334, n56335, n56336, n56337, n56338,
         n56339, n56340, n56341, n56342, n56343, n56344, n56345, n56346,
         n56347, n56348, n56349, n56350, n56351, n56352, n56353, n56354,
         n56355, n56356, n56357, n56358, n56359, n56360, n56361, n56362,
         n56363, n56364, n56365, n56366, n56367, n56368, n56369, n56370,
         n56371, n56372, n56373, n56374, n56375, n56376, n56377, n56378,
         n56379, n56380, n56381, n56382, n56383, n56384, n56385, n56386,
         n56387, n56388, n56389, n56390, n56391, n56392, n56393, n56394,
         n56395, n56396, n56397, n56398, n56399, n56400, n56401, n56402,
         n56403, n56404, n56405, n56406, n56407, n56408, n56409, n56410,
         n56411, n56412, n56413, n56414, n56415, n56416, n56417, n56418,
         n56419, n56420, n56421, n56422, n56423, n56424, n56425, n56426,
         n56427, n56428, n56429, n56430, n56431, n56432, n56433, n56434,
         n56435, n56436, n56437, n56438, n56439, n56440, n56441, n56442,
         n56443, n56444, n56445, n56446, n56447, n56448, n56449, n56450,
         n56451, n56452, n56453, n56454, n56455, n56456, n56457, n56458,
         n56459, n56460, n56461, n56462, n56463, n56464, n56465, n56466,
         n56467, n56468, n56469, n56470, n56471, n56472, n56473, n56474,
         n56475, n56476, n56477, n56478, n56479, n56480, n56481, n56482,
         n56483, n56484, n56485, n56486, n56487, n56488, n56489, n56490,
         n56491, n56492, n56493, n56494, n56495, n56496, n56497, n56498,
         n56499, n56500, n56501, n56502, n56503, n56504, n56505, n56506,
         n56507, n56508, n56509, n56510, n56511, n56512, n56513, n56514,
         n56515, n56516, n56517, n56518, n56519, n56520, n56521, n56522,
         n56523, n56524, n56525, n56526, n56527, n56528, n56529, n56530,
         n56531, n56532, n56533, n56534, n56535, n56536, n56537, n56538,
         n56539, n56540, n56541, n56542, n56543, n56544, n56545, n56546,
         n56547, n56548, n56549, n56550, n56551, n56552, n56553, n56554,
         n56555, n56556, n56557, n56558, n56559, n56560, n56561, n56562,
         n56563, n56564, n56565, n56566, n56567, n56568, n56569, n56570,
         n56571, n56572, n56573, n56574, n56575, n56576, n56577, n56578,
         n56579, n56580, n56581, n56582, n56583, n56584, n56585, n56586,
         n56587, n56588, n56589, n56590, n56591, n56592, n56593, n56594,
         n56595, n56596, n56597, n56598, n56599, n56600, n56601, n56602,
         n56603, n56604, n56605, n56606, n56607, n56608, n56609, n56610,
         n56611, n56612, n56613, n56614, n56615, n56616, n56617, n56618,
         n56619, n56620, n56621, n56622, n56623, n56624, n56625, n56626,
         n56627, n56628, n56629, n56630, n56631, n56632, n56633, n56634,
         n56635, n56636, n56637, n56638, n56639, n56640, n56641, n56642,
         n56643, n56644, n56645, n56646, n56647, n56648, n56649, n56650,
         n56651, n56652, n56653, n56654, n56655, n56656, n56657, n56658,
         n56659, n56660, n56661, n56662, n56663, n56664, n56665, n56666,
         n56667, n56668, n56669, n56670, n56671, n56672, n56673, n56674,
         n56675, n56676, n56677, n56678, n56679, n56680, n56681, n56682,
         n56683, n56684, n56685, n56686, n56687, n56688, n56689, n56690,
         n56691, n56692, n56693, n56694, n56695, n56696, n56697, n56698,
         n56699, n56700, n56701, n56702, n56703, n56704, n56705, n56706,
         n56707, n56708, n56709, n56710, n56711, n56712, n56713, n56714,
         n56715, n56716, n56717, n56718, n56719, n56720, n56721, n56722,
         n56723, n56724, n56725, n56726, n56727, n56728, n56729, n56730,
         n56731, n56732, n56733, n56734, n56735, n56736, n56737, n56738,
         n56739, n56740, n56741, n56742, n56743, n56744, n56745, n56746,
         n56747, n56748, n56749, n56750, n56751, n56752, n56753, n56754,
         n56755, n56756, n56757, n56758, n56759, n56760, n56761, n56762,
         n56763, n56764, n56765, n56766, n56767, n56768, n56769, n56770,
         n56771, n56772, n56773, n56774, n56775, n56776, n56777, n56778,
         n56779, n56780, n56781, n56782, n56783, n56784, n56785, n56786,
         n56787, n56788, n56789, n56790, n56791, n56792, n56793, n56794,
         n56795, n56796, n56797, n56798, n56799, n56800, n56801, n56802,
         n56803, n56804, n56805, n56806, n56807, n56808, n56809, n56810,
         n56811, n56812, n56813, n56814, n56815, n56816, n56817, n56818,
         n56819, n56820, n56821, n56822, n56823, n56824, n56825, n56826,
         n56827, n56828, n56829, n56830, n56831, n56832, n56833, n56834,
         n56835, n56836, n56837, n56838, n56839, n56840, n56841, n56842,
         n56843, n56844, n56845, n56846, n56847, n56848, n56849, n56850,
         n56851, n56852, n56853, n56854, n56855, n56856, n56857, n56858,
         n56859, n56860, n56861, n56862, n56863, n56864, n56865, n56866,
         n56867, n56868, n56869, n56870, n56871, n56872, n56873, n56874,
         n56875, n56876, n56877, n56878, n56879, n56880, n56881, n56882,
         n56883, n56884, n56885, n56886, n56887, n56888, n56889, n56890,
         n56891, n56892, n56893, n56894, n56895, n56896, n56897, n56898,
         n56899, n56900, n56901, n56902, n56903, n56904, n56905, n56906,
         n56907, n56908, n56909, n56910, n56911, n56912, n56913, n56914,
         n56915, n56916, n56917, n56918, n56919, n56920, n56921, n56922,
         n56923, n56924, n56925, n56926, n56927, n56928, n56929, n56930,
         n56931, n56932, n56933, n56934, n56935, n56936, n56937, n56938,
         n56939, n56940, n56941, n56942, n56943, n56944, n56945, n56946,
         n56947, n56948, n56949, n56950, n56951, n56952, n56953, n56954,
         n56955, n56956, n56957, n56958, n56959, n56960, n56961, n56962,
         n56963, n56964, n56965, n56966, n56967, n56968, n56969, n56970,
         n56971, n56972, n56973, n56974, n56975, n56976, n56977, n56978,
         n56979, n56980, n56981, n56982, n56983, n56984, n56985, n56986,
         n56987, n56988, n56989, n56990, n56991, n56992, n56993, n56994,
         n56995, n56996, n56997, n56998, n56999, n57000, n57001, n57002,
         n57003, n57004, n57005, n57006, n57007, n57008, n57009, n57010,
         n57011, n57012, n57013, n57014, n57015, n57016, n57017, n57018,
         n57019, n57020, n57021, n57022, n57023, n57024, n57025, n57026,
         n57027, n57028, n57029, n57030, n57031, n57032, n57033, n57034,
         n57035, n57036, n57037, n57038, n57039, n57040, n57041, n57042,
         n57043, n57044, n57045, n57046, n57047, n57048, n57049, n57050,
         n57051, n57052, n57053, n57054, n57055, n57056, n57057, n57058,
         n57059, n57060, n57061, n57062, n57063, n57064, n57065, n57066,
         n57067, n57068, n57069, n57070, n57071, n57072, n57073, n57074,
         n57075, n57076, n57077, n57078, n57079, n57080, n57081, n57082,
         n57083, n57084, n57085, n57086, n57087, n57088, n57089, n57090,
         n57091, n57092, n57093, n57094, n57095, n57096, n57097, n57098,
         n57099, n57100, n57101, n57102, n57103, n57104, n57105, n57106,
         n57107, n57108, n57109, n57110, n57111, n57112, n57113, n57114,
         n57115, n57116, n57117, n57118, n57119, n57120, n57121, n57122,
         n57123, n57124, n57125, n57126, n57127, n57128, n57129, n57130,
         n57131, n57132, n57133, n57134, n57135, n57136, n57137, n57138,
         n57139, n57140, n57141, n57142, n57143, n57144, n57145, n57146,
         n57147, n57148, n57149, n57150, n57151, n57152, n57153, n57154,
         n57155, n57156, n57157, n57158, n57159, n57160, n57161, n57162,
         n57163, n57164, n57165, n57166, n57167, n57168, n57169, n57170,
         n57171, n57172, n57173, n57174, n57175, n57176, n57177, n57178,
         n57179, n57180, n57181, n57182, n57183, n57184, n57185, n57186,
         n57187, n57188, n57189, n57190, n57191, n57192, n57193, n57194,
         n57195, n57196, n57197, n57198, n57199, n57200, n57201, n57202,
         n57203, n57204, n57205, n57206, n57207, n57208, n57209, n57210,
         n57211, n57212, n57213, n57214, n57215, n57216, n57217, n57218,
         n57219, n57220, n57221, n57222, n57223, n57224, n57225, n57226,
         n57227, n57228, n57229, n57230, n57231, n57232, n57233, n57234,
         n57235, n57236, n57237, n57238, n57239, n57240, n57241, n57242,
         n57243, n57244, n57245, n57246, n57247, n57248, n57249, n57250,
         n57251, n57252, n57253, n57254, n57255, n57256, n57257, n57258,
         n57259, n57260, n57261, n57262, n57263, n57264, n57265, n57266,
         n57267, n57268, n57269, n57270, n57271, n57272, n57273, n57274,
         n57275, n57276, n57277, n57278, n57279, n57280, n57281, n57282,
         n57283, n57284, n57285, n57286, n57287, n57288, n57289, n57290,
         n57291, n57292, n57293, n57294, n57295, n57296, n57297, n57298,
         n57299, n57300, n57301, n57302, n57303, n57304, n57305, n57306,
         n57307, n57308, n57309, n57310, n57311, n57312, n57313, n57314,
         n57315, n57316, n57317, n57318, n57319, n57320, n57321, n57322,
         n57323, n57324, n57325, n57326, n57327, n57328, n57329, n57330,
         n57331, n57332, n57333, n57334, n57335, n57336, n57337, n57338,
         n57339, n57340, n57341, n57342, n57343, n57344, n57345, n57346,
         n57347, n57348, n57349, n57350, n57351, n57352, n57353, n57354,
         n57355, n57356, n57357, n57358, n57359, n57360, n57361, n57362,
         n57363, n57364, n57365, n57366, n57367, n57368, n57369, n57370,
         n57371, n57372, n57373, n57374, n57375, n57376, n57377, n57378,
         n57379, n57380, n57381, n57382, n57383, n57384, n57385, n57386,
         n57387, n57388, n57389, n57390, n57391, n57392, n57393, n57394,
         n57395, n57396, n57397, n57398, n57399, n57400, n57401, n57402,
         n57403, n57404, n57405, n57406, n57407, n57408, n57409, n57410,
         n57411, n57412, n57413, n57414, n57415, n57416, n57417, n57418,
         n57419, n57420, n57421, n57422, n57423, n57424, n57425, n57426,
         n57427, n57428, n57429, n57430, n57431, n57432, n57433, n57434,
         n57435, n57436, n57437, n57438, n57439, n57440, n57441, n57442,
         n57443, n57444, n57445, n57446, n57447, n57448, n57449, n57450,
         n57451, n57452, n57453, n57454, n57455, n57456, n57457, n57458,
         n57459, n57460, n57461, n57462, n57463, n57464, n57465, n57466,
         n57467, n57468, n57469, n57470, n57471, n57472, n57473, n57474,
         n57475, n57476, n57477, n57478, n57479, n57480, n57481, n57482,
         n57483, n57484, n57485, n57486, n57487, n57488, n57489, n57490,
         n57491, n57492, n57493, n57494, n57495, n57496, n57497, n57498,
         n57499, n57500, n57501, n57502, n57503, n57504, n57505, n57506,
         n57507, n57508, n57509, n57510, n57511, n57512, n57513, n57514,
         n57515, n57516, n57517, n57518, n57519, n57520, n57521, n57522,
         n57523, n57524, n57525, n57526, n57527, n57528, n57529, n57530,
         n57531, n57532, n57533, n57534, n57535, n57536, n57537, n57538,
         n57539, n57540, n57541, n57542, n57543, n57544, n57545, n57546,
         n57547, n57548, n57549, n57550, n57551, n57552, n57553, n57554,
         n57555, n57556, n57557, n57558, n57559, n57560, n57561, n57562,
         n57563, n57564, n57565, n57566, n57567, n57568, n57569, n57570,
         n57571, n57572, n57573, n57574, n57575, n57576, n57577, n57578,
         n57579, n57580, n57581, n57582, n57583, n57584, n57585, n57586,
         n57587, n57588, n57589, n57590, n57591, n57592, n57593, n57594,
         n57595, n57596, n57597, n57598, n57599, n57600, n57601, n57602,
         n57603, n57604, n57605, n57606, n57607, n57608, n57609, n57610,
         n57611, n57612, n57613, n57614, n57615, n57616, n57617, n57618,
         n57619, n57620, n57621, n57622, n57623, n57624, n57625, n57626,
         n57627, n57628, n57629, n57630, n57631, n57632, n57633, n57634,
         n57635, n57636, n57637, n57638, n57639, n57640, n57641, n57642,
         n57643, n57644, n57645, n57646, n57647, n57648, n57649, n57650,
         n57651, n57652, n57653, n57654, n57655, n57656, n57657, n57658,
         n57659, n57660, n57661, n57662, n57663, n57664, n57665, n57666,
         n57667, n57668, n57669, n57670, n57671, n57672, n57673, n57674,
         n57675, n57676, n57677, n57678, n57679, n57680, n57681, n57682,
         n57683, n57684, n57685, n57686, n57687, n57688, n57689, n57690,
         n57691, n57692, n57693, n57694, n57695, n57696, n57697, n57698,
         n57699, n57700, n57701, n57702, n57703, n57704, n57705, n57706,
         n57707, n57708, n57709, n57710, n57711, n57712, n57713, n57714,
         n57715, n57716, n57717, n57718, n57719, n57720, n57721, n57722,
         n57723, n57724, n57725, n57726, n57727, n57728, n57729, n57730,
         n57731, n57732, n57733, n57734, n57735, n57736, n57737, n57738,
         n57739, n57740, n57741, n57742, n57743, n57744, n57745, n57746,
         n57747, n57748, n57749, n57750, n57751, n57752, n57753, n57754,
         n57755, n57756, n57757, n57758, n57759, n57760, n57761, n57762,
         n57763, n57764, n57765, n57766, n57767, n57768, n57769, n57770,
         n57771, n57772, n57773, n57774, n57775, n57776, n57777, n57778,
         n57779, n57780, n57781, n57782, n57783, n57784, n57785, n57786,
         n57787, n57788, n57789, n57790, n57791, n57792, n57793, n57794,
         n57795, n57796, n57797, n57798, n57799, n57800, n57801, n57802,
         n57803, n57804, n57805, n57806, n57807, n57808, n57809, n57810,
         n57811, n57812, n57813, n57814, n57815, n57816, n57817, n57818,
         n57819, n57820, n57821, n57822, n57823, n57824, n57825, n57826,
         n57827, n57828, n57829, n57830, n57831, n57832, n57833, n57834,
         n57835, n57836, n57837, n57838, n57839, n57840, n57841, n57842,
         n57843, n57844, n57845, n57846, n57847, n57848, n57849, n57850,
         n57851, n57852, n57853, n57854, n57855, n57856, n57857, n57858,
         n57859, n57860, n57861, n57862, n57863, n57864, n57865, n57866,
         n57867, n57868, n57869, n57870, n57871, n57872, n57873, n57874,
         n57875, n57876, n57877, n57878, n57879, n57880, n57881, n57882,
         n57883, n57884, n57885, n57886, n57887, n57888, n57889, n57890,
         n57891, n57892, n57893, n57894, n57895, n57896, n57897, n57898,
         n57899, n57900, n57901, n57902, n57903, n57904, n57905, n57906,
         n57907, n57908, n57909, n57910, n57911, n57912, n57913, n57914,
         n57915, n57916, n57917, n57918, n57919, n57920, n57921, n57922,
         n57923, n57924, n57925, n57926, n57927, n57928, n57929, n57930,
         n57931, n57932, n57933, n57934, n57935, n57936, n57937, n57938,
         n57939, n57940, n57941, n57942, n57943, n57944, n57945, n57946,
         n57947, n57948, n57949, n57950, n57951, n57952, n57953, n57954,
         n57955, n57956, n57957, n57958, n57959, n57960, n57961, n57962,
         n57963, n57964, n57965, n57966, n57967, n57968, n57969, n57970,
         n57971, n57972, n57973, n57974, n57975, n57976, n57977, n57978,
         n57979, n57980, n57981, n57982, n57983, n57984, n57985, n57986,
         n57987, n57988, n57989, n57990, n57991, n57992, n57993, n57994,
         n57995, n57996, n57997, n57998, n57999, n58000, n58001, n58002,
         n58003, n58004, n58005, n58006, n58007, n58008, n58009, n58010,
         n58011, n58012, n58013, n58014, n58015, n58016, n58017, n58018,
         n58019, n58020, n58021, n58022, n58023, n58024, n58025, n58026,
         n58027, n58028, n58029, n58030, n58031, n58032, n58033, n58034,
         n58035, n58036, n58037, n58038, n58039, n58040, n58041, n58042,
         n58043, n58044, n58045, n58046, n58047, n58048, n58049, n58050,
         n58051, n58052, n58053, n58054, n58055, n58056, n58057, n58058,
         n58059, n58060, n58061, n58062, n58063, n58064, n58065, n58066,
         n58067, n58068, n58069, n58070, n58071, n58072, n58073, n58074,
         n58075, n58076, n58077, n58078, n58079, n58080, n58081, n58082,
         n58083, n58084, n58085, n58086, n58087, n58088, n58089, n58090,
         n58091, n58092, n58093, n58094, n58095, n58096, n58097, n58098,
         n58099, n58100, n58101, n58102, n58103, n58104, n58105, n58106,
         n58107, n58108, n58109, n58110, n58111, n58112, n58113, n58114,
         n58115, n58116, n58117, n58118, n58119, n58120, n58121, n58122,
         n58123, n58124, n58125, n58126, n58127, n58128, n58129, n58130,
         n58131, n58132, n58133, n58134, n58135, n58136, n58137, n58138,
         n58139, n58140, n58141, n58142, n58143, n58144, n58145, n58146,
         n58147, n58148, n58149, n58150, n58151, n58152, n58153, n58154,
         n58155, n58156, n58157, n58158, n58159, n58160, n58161, n58162,
         n58163, n58164, n58165, n58166, n58167, n58168, n58169, n58170,
         n58171, n58172, n58173, n58174, n58175, n58176, n58177, n58178,
         n58179, n58180, n58181, n58182, n58183, n58184, n58185, n58186,
         n58187, n58188, n58189, n58190, n58191, n58192, n58193, n58194,
         n58195, n58196, n58197, n58198, n58199, n58200, n58201, n58202,
         n58203, n58204, n58205, n58206, n58207, n58208, n58209, n58210,
         n58211, n58212, n58213, n58214, n58215, n58216, n58217, n58218,
         n58219, n58220, n58221, n58222, n58223, n58224, n58225, n58226,
         n58227, n58228, n58229, n58230, n58231, n58232, n58233, n58234,
         n58235, n58236, n58237, n58238, n58239, n58240, n58241, n58242,
         n58243, n58244, n58245, n58246, n58247, n58248, n58249, n58250,
         n58251, n58252, n58253, n58254, n58255, n58256, n58257, n58258,
         n58259, n58260, n58261, n58262, n58263, n58264, n58265, n58266,
         n58267, n58268, n58269, n58270, n58271, n58272, n58273, n58274,
         n58275, n58276, n58277, n58278, n58279, n58280, n58281, n58282,
         n58283, n58284, n58285, n58286, n58287, n58288, n58289, n58290,
         n58291, n58292, n58293, n58294, n58295, n58296, n58297, n58298,
         n58299, n58300, n58301, n58302, n58303, n58304, n58305, n58306,
         n58307, n58308, n58309, n58310, n58311, n58312, n58313, n58314,
         n58315, n58316, n58317, n58318, n58319, n58320, n58321, n58322,
         n58323, n58324, n58325, n58326, n58327, n58328, n58329, n58330,
         n58331, n58332, n58333, n58334, n58335, n58336, n58337, n58338,
         n58339, n58340, n58341, n58342, n58343, n58344, n58345, n58346,
         n58347, n58348, n58349, n58350, n58351, n58352, n58353, n58354,
         n58355, n58356, n58357, n58358, n58359, n58360, n58361, n58362,
         n58363, n58364, n58365, n58366, n58367, n58368, n58369, n58370,
         n58371, n58372, n58373, n58374, n58375, n58376, n58377, n58378,
         n58379, n58380, n58381, n58382, n58383, n58384, n58385, n58386,
         n58387, n58388, n58389, n58390, n58391, n58392, n58393, n58394,
         n58395, n58396, n58397, n58398, n58399, n58400, n58401, n58402,
         n58403, n58404, n58405, n58406, n58407, n58408, n58409, n58410,
         n58411, n58412, n58413, n58414, n58415, n58416, n58417, n58418,
         n58419, n58420, n58421, n58422, n58423, n58424, n58425, n58426,
         n58427, n58428, n58429, n58430, n58431, n58432, n58433, n58434,
         n58435, n58436, n58437, n58438, n58439, n58440, n58441, n58442,
         n58443, n58444, n58445, n58446, n58447, n58448, n58449, n58450,
         n58451, n58452, n58453, n58454, n58455, n58456, n58457, n58458,
         n58459, n58460, n58461, n58462, n58463, n58464, n58465, n58466,
         n58467, n58468, n58469, n58470, n58471, n58472, n58473, n58474,
         n58475, n58476, n58477, n58478, n58479, n58480, n58481, n58482,
         n58483, n58484, n58485, n58486, n58487, n58488, n58489, n58490,
         n58491, n58492, n58493, n58494, n58495, n58496, n58497, n58498,
         n58499, n58500, n58501, n58502, n58503, n58504, n58505, n58506,
         n58507, n58508, n58509, n58510, n58511, n58512, n58513, n58514,
         n58515, n58516, n58517, n58518, n58519, n58520, n58521, n58522,
         n58523, n58524, n58525, n58526, n58527, n58528, n58529, n58530,
         n58531, n58532, n58533, n58534, n58535, n58536, n58537, n58538,
         n58539, n58540, n58541, n58542, n58543, n58544, n58545, n58546,
         n58547, n58548, n58549, n58550, n58551, n58552, n58553, n58554,
         n58555, n58556, n58557, n58558, n58559, n58560, n58561, n58562,
         n58563, n58564, n58565, n58566, n58567, n58568, n58569, n58570,
         n58571, n58572, n58573, n58574, n58575, n58576, n58577, n58578,
         n58579, n58580, n58581, n58582, n58583, n58584, n58585, n58586,
         n58587, n58588, n58589, n58590, n58591, n58592, n58593, n58594,
         n58595, n58596, n58597, n58598, n58599, n58600, n58601, n58602,
         n58603, n58604, n58605, n58606, n58607, n58608, n58609, n58610,
         n58611, n58612, n58613, n58614, n58615, n58616, n58617, n58618,
         n58619, n58620, n58621, n58622, n58623, n58624, n58625, n58626,
         n58627, n58628, n58629, n58630, n58631, n58632, n58633, n58634,
         n58635, n58636, n58637, n58638, n58639, n58640, n58641, n58642,
         n58643, n58644, n58645, n58646, n58647, n58648, n58649, n58650,
         n58651, n58652, n58653, n58654, n58655, n58656, n58657, n58658,
         n58659, n58660, n58661, n58662, n58663, n58664, n58665, n58666,
         n58667, n58668, n58669, n58670, n58671, n58672, n58673, n58674,
         n58675, n58676, n58677, n58678, n58679, n58680, n58681, n58682,
         n58683, n58684, n58685, n58686, n58687, n58688, n58689, n58690,
         n58691, n58692, n58693, n58694, n58695, n58696, n58697, n58698,
         n58699, n58700, n58701, n58702, n58703, n58704, n58705, n58706,
         n58707, n58708, n58709, n58710, n58711, n58712, n58713, n58714,
         n58715, n58716, n58717, n58718, n58719, n58720, n58721, n58722,
         n58723, n58724, n58725, n58726, n58727, n58728, n58729, n58730,
         n58731, n58732, n58733, n58734, n58735, n58736, n58737, n58738,
         n58739, n58740, n58741, n58742, n58743, n58744, n58745, n58746,
         n58747, n58748, n58749, n58750, n58751, n58752, n58753, n58754,
         n58755, n58756, n58757, n58758, n58759, n58760, n58761, n58762,
         n58763, n58764, n58765, n58766, n58767, n58768, n58769, n58770,
         n58771, n58772, n58773, n58774, n58775, n58776, n58777, n58778,
         n58779, n58780, n58781, n58782, n58783, n58784, n58785, n58786,
         n58787, n58788, n58789, n58790, n58791, n58792, n58793, n58794,
         n58795, n58796, n58797, n58798, n58799, n58800, n58801, n58802,
         n58803, n58804, n58805, n58806, n58807, n58808, n58809, n58810,
         n58811, n58812, n58813, n58814, n58815, n58816, n58817, n58818,
         n58819, n58820, n58821, n58822, n58823, n58824, n58825, n58826,
         n58827, n58828, n58829, n58830, n58831, n58832, n58833, n58834,
         n58835, n58836, n58837, n58838, n58839, n58840, n58841, n58842,
         n58843, n58844, n58845, n58846, n58847, n58848, n58849, n58850,
         n58851, n58852, n58853, n58854, n58855, n58856, n58857, n58858,
         n58859, n58860, n58861, n58862, n58863, n58864, n58865, n58866,
         n58867, n58868, n58869, n58870, n58871, n58872, n58873, n58874,
         n58875, n58876, n58877, n58878, n58879, n58880, n58881, n58882,
         n58883, n58884, n58885, n58886, n58887, n58888, n58889, n58890,
         n58891, n58892, n58893, n58894, n58895, n58896, n58897, n58898,
         n58899, n58900, n58901, n58902, n58903, n58904, n58905, n58906,
         n58907, n58908, n58909, n58910, n58911, n58912, n58913, n58914,
         n58915, n58916, n58917, n58918, n58919, n58920, n58921, n58922,
         n58923, n58924, n58925, n58926, n58927, n58928, n58929, n58930,
         n58931, n58932, n58933, n58934, n58935, n58936, n58937, n58938,
         n58939, n58940, n58941, n58942, n58943, n58944, n58945, n58946,
         n58947, n58948, n58949, n58950, n58951, n58952, n58953, n58954,
         n58955, n58956, n58957, n58958, n58959, n58960, n58961, n58962,
         n58963, n58964, n58965, n58966, n58967, n58968, n58969, n58970,
         n58971, n58972, n58973, n58974, n58975, n58976, n58977, n58978,
         n58979, n58980, n58981, n58982, n58983, n58984, n58985, n58986,
         n58987, n58988, n58989, n58990, n58991, n58992, n58993, n58994,
         n58995, n58996, n58997, n58998, n58999, n59000, n59001, n59002,
         n59003, n59004, n59005, n59006, n59007, n59008, n59009, n59010,
         n59011, n59012, n59013, n59014, n59015, n59016, n59017, n59018,
         n59019, n59020, n59021, n59022, n59023, n59024, n59025, n59026,
         n59027, n59028, n59029, n59030, n59031, n59032, n59033, n59034,
         n59035, n59036, n59037, n59038, n59039, n59040, n59041, n59042,
         n59043, n59044, n59045, n59046, n59047, n59048, n59049, n59050,
         n59051, n59052, n59053, n59054, n59055, n59056, n59057, n59058,
         n59059, n59060, n59061, n59062, n59063, n59064, n59065, n59066,
         n59067, n59068, n59069, n59070, n59071, n59072, n59073, n59074,
         n59075, n59076, n59077, n59078, n59079, n59080, n59081, n59082,
         n59083, n59084, n59085, n59086, n59087, n59088, n59089, n59090,
         n59091, n59092, n59093, n59094, n59095, n59096, n59097, n59098,
         n59099, n59100, n59101, n59102, n59103, n59104, n59105, n59106,
         n59107, n59108, n59109, n59110, n59111, n59112, n59113, n59114,
         n59115, n59116, n59117, n59118, n59119, n59120, n59121, n59122,
         n59123, n59124, n59125, n59126, n59127, n59128, n59129, n59130,
         n59131, n59132, n59133, n59134, n59135, n59136, n59137, n59138,
         n59139, n59140, n59141, n59142, n59143, n59144, n59145, n59146,
         n59147, n59148, n59149, n59150, n59151, n59152, n59153, n59154,
         n59155, n59156, n59157, n59158, n59159, n59160, n59161, n59162,
         n59163, n59164, n59165, n59166, n59167, n59168, n59169, n59170,
         n59171, n59172, n59173, n59174, n59175, n59176, n59177, n59178,
         n59179, n59180, n59181, n59182, n59183, n59184, n59185, n59186,
         n59187, n59188, n59189, n59190, n59191, n59192, n59193, n59194,
         n59195, n59196, n59197, n59198, n59199, n59200, n59201, n59202,
         n59203, n59204, n59205, n59206, n59207, n59208, n59209, n59210,
         n59211, n59212, n59213, n59214, n59215, n59216, n59217, n59218,
         n59219, n59220, n59221, n59222, n59223, n59224, n59225, n59226,
         n59227, n59228, n59229, n59230, n59231, n59232, n59233, n59234,
         n59235, n59236, n59237, n59238, n59239, n59240, n59241, n59242,
         n59243, n59244, n59245, n59246, n59247, n59248, n59249, n59250,
         n59251, n59252, n59253, n59254, n59255, n59256, n59257, n59258,
         n59259, n59260, n59261, n59262, n59263, n59264, n59265, n59266,
         n59267, n59268, n59269, n59270, n59271, n59272, n59273, n59274,
         n59275, n59276, n59277, n59278, n59279, n59280, n59281, n59282,
         n59283, n59284, n59285, n59286, n59287, n59288, n59289, n59290,
         n59291, n59292, n59293, n59294, n59295, n59296, n59297, n59298,
         n59299, n59300, n59301, n59302, n59303, n59304, n59305, n59306,
         n59307, n59308, n59309, n59310, n59311, n59312, n59313, n59314,
         n59315, n59316, n59317, n59318, n59319, n59320, n59321, n59322,
         n59323, n59324, n59325, n59326, n59327, n59328, n59329, n59330,
         n59331, n59332, n59333, n59334, n59335, n59336, n59337, n59338,
         n59339, n59340, n59341, n59342, n59343, n59344, n59345, n59346,
         n59347, n59348, n59349, n59350, n59351, n59352, n59353, n59354,
         n59355, n59356, n59357, n59358, n59359, n59360, n59361, n59362,
         n59363, n59364, n59365, n59366, n59367, n59368, n59369, n59370,
         n59371, n59372, n59373, n59374, n59375, n59376, n59377, n59378,
         n59379, n59380, n59381, n59382, n59383, n59384, n59385, n59386,
         n59387, n59388, n59389, n59390, n59391, n59392, n59393, n59394,
         n59395, n59396, n59397, n59398, n59399, n59400, n59401, n59402,
         n59403, n59404, n59405, n59406, n59407, n59408, n59409, n59410,
         n59411, n59412, n59413, n59414, n59415, n59416, n59417, n59418,
         n59419, n59420, n59421, n59422, n59423, n59424, n59425, n59426,
         n59427, n59428, n59429, n59430, n59431, n59432, n59433, n59434,
         n59435, n59436, n59437, n59438, n59439, n59440, n59441, n59442,
         n59443, n59444, n59445, n59446, n59447, n59448, n59449, n59450,
         n59451, n59452, n59453, n59454, n59455, n59456, n59457, n59458,
         n59459, n59460, n59461, n59462, n59463, n59464, n59465, n59466,
         n59467, n59468, n59469, n59470, n59471, n59472, n59473, n59474,
         n59475, n59476, n59477, n59478, n59479, n59480, n59481, n59482,
         n59483, n59484, n59485, n59486, n59487, n59488, n59489, n59490,
         n59491, n59492, n59493, n59494, n59495, n59496, n59497, n59498,
         n59499, n59500, n59501, n59502, n59503, n59504, n59505, n59506,
         n59507, n59508, n59509, n59510, n59511, n59512, n59513, n59514,
         n59515, n59516, n59517, n59518, n59519, n59520, n59521, n59522,
         n59523, n59524, n59525, n59526, n59527, n59528, n59529, n59530,
         n59531, n59532, n59533, n59534, n59535, n59536, n59537, n59538,
         n59539, n59540, n59541, n59542, n59543, n59544, n59545, n59546,
         n59547, n59548, n59549, n59550, n59551, n59552, n59553, n59554,
         n59555, n59556, n59557, n59558, n59559, n59560, n59561, n59562,
         n59563, n59564, n59565, n59566, n59567, n59568, n59569, n59570,
         n59571, n59572, n59573, n59574, n59575, n59576, n59577, n59578,
         n59579, n59580, n59581, n59582, n59583, n59584, n59585, n59586,
         n59587, n59588, n59589, n59590, n59591, n59592, n59593, n59594,
         n59595, n59596, n59597, n59598, n59599, n59600, n59601, n59602,
         n59603, n59604, n59605, n59606, n59607, n59608, n59609, n59610,
         n59611, n59612, n59613, n59614, n59615, n59616, n59617, n59618,
         n59619, n59620, n59621, n59622, n59623, n59624, n59625, n59626,
         n59627, n59628, n59629, n59630, n59631, n59632, n59633, n59634,
         n59635, n59636, n59637, n59638, n59639, n59640, n59641, n59642,
         n59643, n59644, n59645, n59646, n59647, n59648, n59649, n59650,
         n59651, n59652, n59653, n59654, n59655, n59656, n59657, n59658,
         n59659, n59660, n59661, n59662, n59663, n59664, n59665, n59666,
         n59667, n59668, n59669, n59670, n59671, n59672, n59673, n59674,
         n59675, n59676, n59677, n59678, n59679, n59680, n59681, n59682,
         n59683, n59684, n59685, n59686, n59687, n59688, n59689, n59690,
         n59691, n59692, n59693, n59694, n59695, n59696, n59697, n59698,
         n59699, n59700, n59701, n59702, n59703, n59704, n59705, n59706,
         n59707, n59708, n59709, n59710, n59711, n59712, n59713, n59714,
         n59715, n59716, n59717, n59718, n59719, n59720, n59721, n59722,
         n59723, n59724, n59725, n59726, n59727, n59728, n59729, n59730,
         n59731, n59732, n59733, n59734, n59735, n59736, n59737, n59738,
         n59739, n59740, n59741, n59742, n59743, n59744, n59745, n59746,
         n59747, n59748, n59749, n59750, n59751, n59752, n59753, n59754,
         n59755, n59756, n59757, n59758, n59759, n59760, n59761, n59762,
         n59763, n59764, n59765, n59766, n59767, n59768, n59769, n59770,
         n59771, n59772, n59773, n59774, n59775, n59776, n59777, n59778,
         n59779, n59780, n59781, n59782, n59783, n59784, n59785, n59786,
         n59787, n59788, n59789, n59790, n59791, n59792, n59793, n59794,
         n59795, n59796, n59797, n59798, n59799, n59800, n59801, n59802,
         n59803, n59804, n59805, n59806, n59807, n59808, n59809, n59810,
         n59811, n59812, n59813, n59814, n59815, n59816, n59817, n59818,
         n59819, n59820, n59821, n59822, n59823, n59824, n59825, n59826,
         n59827, n59828, n59829, n59830, n59831, n59832, n59833, n59834,
         n59835, n59836, n59837, n59838, n59839, n59840, n59841, n59842,
         n59843, n59844, n59845, n59846, n59847, n59848, n59849, n59850,
         n59851, n59852, n59853, n59854, n59855, n59856, n59857, n59858,
         n59859, n59860, n59861, n59862, n59863, n59864, n59865, n59866,
         n59867, n59868, n59869, n59870, n59871, n59872, n59873, n59874,
         n59875, n59876, n59877, n59878, n59879, n59880, n59881, n59882,
         n59883, n59884, n59885, n59886, n59887, n59888, n59889, n59890,
         n59891, n59892, n59893, n59894, n59895, n59896, n59897, n59898,
         n59899, n59900, n59901, n59902, n59903, n59904, n59905, n59906,
         n59907, n59908, n59909, n59910, n59911, n59912, n59913, n59914,
         n59915, n59916, n59917, n59918, n59919, n59920, n59921, n59922,
         n59923, n59924, n59925, n59926, n59927, n59928, n59929, n59930,
         n59931, n59932, n59933, n59934, n59935, n59936, n59937, n59938,
         n59939, n59940, n59941, n59942, n59943, n59944, n59945, n59946,
         n59947, n59948, n59949, n59950, n59951, n59952, n59953, n59954,
         n59955, n59956, n59957, n59958, n59959, n59960, n59961, n59962,
         n59963, n59964, n59965, n59966, n59967, n59968, n59969, n59970,
         n59971, n59972, n59973, n59974, n59975, n59976, n59977, n59978,
         n59979, n59980, n59981, n59982, n59983, n59984, n59985, n59986,
         n59987, n59988, n59989, n59990, n59991, n59992, n59993, n59994,
         n59995, n59996, n59997, n59998, n59999, n60000, n60001, n60002,
         n60003, n60004, n60005, n60006, n60007, n60008, n60009, n60010,
         n60011, n60012, n60013, n60014, n60015, n60016, n60017, n60018,
         n60019, n60020, n60021, n60022, n60023, n60024, n60025, n60026,
         n60027, n60028, n60029, n60030, n60031, n60032, n60033, n60034,
         n60035, n60036, n60037, n60038, n60039, n60040, n60041, n60042,
         n60043, n60044, n60045, n60046, n60047, n60048, n60049, n60050,
         n60051, n60052, n60053, n60054, n60055, n60056, n60057, n60058,
         n60059, n60060, n60061, n60062, n60063, n60064, n60065, n60066,
         n60067, n60068, n60069, n60070, n60071, n60072, n60073, n60074,
         n60075, n60076, n60077, n60078, n60079, n60080, n60081, n60082,
         n60083, n60084, n60085, n60086, n60087, n60088, n60089, n60090,
         n60091, n60092, n60093, n60094, n60095, n60096, n60097, n60098,
         n60099, n60100, n60101, n60102, n60103, n60104, n60105, n60106,
         n60107, n60108, n60109, n60110, n60111, n60112, n60113, n60114,
         n60115, n60116, n60117, n60118, n60119, n60120, n60121, n60122,
         n60123, n60124, n60125, n60126, n60127, n60128, n60129, n60130,
         n60131, n60132, n60133, n60134, n60135, n60136, n60137, n60138,
         n60139, n60140, n60141, n60142, n60143, n60144, n60145, n60146,
         n60147, n60148, n60149, n60150, n60151, n60152, n60153, n60154,
         n60155, n60156, n60157, n60158, n60159, n60160, n60161, n60162,
         n60163, n60164, n60165, n60166, n60167, n60168, n60169, n60170,
         n60171, n60172, n60173, n60174, n60175, n60176, n60177, n60178,
         n60179, n60180, n60181, n60182, n60183, n60184, n60185, n60186,
         n60187, n60188, n60189, n60190, n60191, n60192, n60193, n60194,
         n60195, n60196, n60197, n60198, n60199, n60200, n60201, n60202,
         n60203, n60204, n60205, n60206, n60207, n60208, n60209, n60210,
         n60211, n60212, n60213, n60214, n60215, n60216, n60217, n60218,
         n60219, n60220, n60221, n60222, n60223, n60224, n60225, n60226,
         n60227, n60228, n60229, n60230, n60231, n60232, n60233, n60234,
         n60235, n60236, n60237, n60238, n60239, n60240, n60241, n60242,
         n60243, n60244, n60245, n60246, n60247, n60248, n60249, n60250,
         n60251, n60252, n60253, n60254, n60255, n60256, n60257, n60258,
         n60259, n60260, n60261, n60262, n60263, n60264, n60265, n60266,
         n60267, n60268, n60269, n60270, n60271, n60272, n60273, n60274,
         n60275, n60276, n60277, n60278, n60279, n60280, n60281, n60282,
         n60283, n60284, n60285, n60286, n60287, n60288, n60289, n60290,
         n60291, n60292, n60293, n60294, n60295, n60296, n60297, n60298,
         n60299, n60300, n60301, n60302, n60303, n60304, n60305, n60306,
         n60307, n60308, n60309, n60310, n60311, n60312, n60313, n60314,
         n60315, n60316, n60317, n60318, n60319, n60320, n60321, n60322,
         n60323, n60324, n60325, n60326, n60327, n60328, n60329, n60330,
         n60331, n60332, n60333, n60334, n60335, n60336, n60337, n60338,
         n60339, n60340, n60341, n60342, n60343, n60344, n60345, n60346,
         n60347, n60348, n60349, n60350, n60351, n60352, n60353, n60354,
         n60355, n60356, n60357, n60358, n60359, n60360, n60361, n60362,
         n60363, n60364, n60365, n60366, n60367, n60368, n60369, n60370,
         n60371, n60372, n60373, n60374, n60375, n60376, n60377, n60378,
         n60379, n60380, n60381, n60382, n60383, n60384, n60385, n60386,
         n60387, n60388, n60389, n60390, n60391, n60392, n60393, n60394,
         n60395, n60396, n60397, n60398, n60399, n60400, n60401, n60402,
         n60403, n60404, n60405, n60406, n60407, n60408, n60409, n60410,
         n60411, n60412, n60413, n60414, n60415, n60416, n60417, n60418,
         n60419, n60420, n60421, n60422, n60423, n60424, n60425, n60426,
         n60427, n60428, n60429, n60430, n60431, n60432, n60433, n60434,
         n60435, n60436, n60437, n60438, n60439, n60440, n60441, n60442,
         n60443, n60444, n60445, n60446, n60447, n60448, n60449, n60450,
         n60451, n60452, n60453, n60454, n60455, n60456, n60457, n60458,
         n60459, n60460, n60461, n60462, n60463, n60464, n60465, n60466,
         n60467, n60468, n60469, n60470, n60471, n60472, n60473, n60474,
         n60475, n60476, n60477, n60478, n60479, n60480, n60481, n60482,
         n60483, n60484, n60485, n60486, n60487, n60488, n60489, n60490,
         n60491, n60492, n60493, n60494, n60495, n60496, n60497, n60498,
         n60499, n60500, n60501, n60502, n60503, n60504, n60505, n60506,
         n60507, n60508, n60509, n60510, n60511, n60512, n60513, n60514,
         n60515, n60516, n60517, n60518, n60519, n60520, n60521, n60522,
         n60523, n60524, n60525, n60526, n60527, n60528, n60529, n60530,
         n60531, n60532, n60533, n60534, n60535, n60536, n60537, n60538,
         n60539, n60540, n60541, n60542, n60543, n60544, n60545, n60546,
         n60547, n60548, n60549, n60550, n60551, n60552, n60553, n60554,
         n60555, n60556, n60557, n60558, n60559, n60560, n60561, n60562,
         n60563, n60564, n60565, n60566, n60567, n60568, n60569, n60570,
         n60571, n60572, n60573, n60574, n60575, n60576, n60577, n60578,
         n60579, n60580, n60581, n60582, n60583, n60584, n60585, n60586,
         n60587, n60588, n60589, n60590, n60591, n60592, n60593, n60594,
         n60595, n60596, n60597, n60598, n60599, n60600, n60601, n60602,
         n60603, n60604, n60605, n60606, n60607, n60608, n60609, n60610,
         n60611, n60612, n60613, n60614, n60615, n60616, n60617, n60618,
         n60619, n60620, n60621, n60622, n60623, n60624, n60625, n60626,
         n60627, n60628, n60629, n60630, n60631, n60632, n60633, n60634,
         n60635, n60636, n60637, n60638, n60639, n60640, n60641, n60642,
         n60643, n60644, n60645, n60646, n60647, n60648, n60649, n60650,
         n60651, n60652, n60653, n60654, n60655, n60656, n60657, n60658,
         n60659, n60660, n60661, n60662, n60663, n60664, n60665, n60666,
         n60667, n60668, n60669, n60670, n60671, n60672, n60673, n60674,
         n60675, n60676, n60677, n60678, n60679, n60680, n60681, n60682,
         n60683, n60684, n60685, n60686, n60687, n60688, n60689, n60690,
         n60691, n60692, n60693, n60694, n60695, n60696, n60697, n60698,
         n60699, n60700, n60701, n60702, n60703, n60704, n60705, n60706,
         n60707, n60708, n60709, n60710, n60711, n60712, n60713, n60714,
         n60715, n60716, n60717, n60718, n60719, n60720, n60721, n60722,
         n60723, n60724, n60725, n60726, n60727, n60728, n60729, n60730,
         n60731, n60732, n60733, n60734, n60735, n60736, n60737, n60738,
         n60739, n60740, n60741, n60742, n60743, n60744, n60745, n60746,
         n60747, n60748, n60749, n60750, n60751, n60752, n60753, n60754,
         n60755, n60756, n60757, n60758, n60759, n60760, n60761, n60762,
         n60763, n60764, n60765, n60766, n60767, n60768, n60769, n60770,
         n60771, n60772, n60773, n60774, n60775, n60776, n60777, n60778,
         n60779, n60780, n60781, n60782, n60783, n60784, n60785, n60786,
         n60787, n60788, n60789, n60790, n60791, n60792, n60793, n60794,
         n60795, n60796, n60797, n60798, n60799, n60800, n60801, n60802,
         n60803, n60804, n60805, n60806, n60807, n60808, n60809, n60810,
         n60811, n60812, n60813, n60814, n60815, n60816, n60817, n60818,
         n60819, n60820, n60821, n60822, n60823, n60824, n60825, n60826,
         n60827, n60828, n60829, n60830, n60831, n60832, n60833, n60834,
         n60835, n60836, n60837, n60838, n60839, n60840, n60841, n60842,
         n60843, n60844, n60845, n60846, n60847, n60848, n60849, n60850,
         n60851, n60852, n60853, n60854, n60855, n60856, n60857, n60858,
         n60859, n60860, n60861, n60862, n60863, n60864, n60865, n60866,
         n60867, n60868, n60869, n60870, n60871, n60872, n60873, n60874,
         n60875, n60876, n60877, n60878, n60879, n60880, n60881, n60882,
         n60883, n60884, n60885, n60886, n60887, n60888, n60889, n60890,
         n60891, n60892, n60893, n60894, n60895, n60896, n60897, n60898,
         n60899, n60900, n60901, n60902, n60903, n60904, n60905, n60906,
         n60907, n60908, n60909, n60910, n60911, n60912, n60913, n60914,
         n60915, n60916, n60917, n60918, n60919, n60920, n60921, n60922,
         n60923, n60924, n60925, n60926, n60927, n60928, n60929, n60930,
         n60931, n60932, n60933, n60934, n60935, n60936, n60937, n60938,
         n60939, n60940, n60941, n60942, n60943, n60944, n60945, n60946,
         n60947, n60948, n60949, n60950, n60951, n60952, n60953, n60954,
         n60955, n60956, n60957, n60958, n60959, n60960, n60961, n60962,
         n60963, n60964, n60965, n60966, n60967, n60968, n60969, n60970,
         n60971, n60972, n60973, n60974, n60975, n60976, n60977, n60978,
         n60979, n60980, n60981, n60982, n60983, n60984, n60985, n60986,
         n60987, n60988, n60989, n60990, n60991, n60992, n60993, n60994,
         n60995, n60996, n60997, n60998, n60999, n61000, n61001, n61002,
         n61003, n61004, n61005, n61006, n61007, n61008, n61009, n61010,
         n61011, n61012, n61013, n61014, n61015, n61016, n61017, n61018,
         n61019, n61020, n61021, n61022, n61023, n61024, n61025, n61026,
         n61027, n61028, n61029, n61030, n61031, n61032, n61033, n61034,
         n61035, n61036, n61037, n61038, n61039, n61040, n61041, n61042,
         n61043, n61044, n61045, n61046, n61047, n61048, n61049, n61050,
         n61051, n61052, n61053, n61054, n61055, n61056, n61057, n61058,
         n61059, n61060, n61061, n61062, n61063, n61064, n61065, n61066,
         n61067, n61068, n61069, n61070, n61071, n61072, n61073, n61074,
         n61075, n61076, n61077, n61078, n61079, n61080, n61081, n61082,
         n61083, n61084, n61085, n61086, n61087, n61088, n61089, n61090,
         n61091, n61092, n61093, n61094, n61095, n61096, n61097, n61098,
         n61099, n61100, n61101, n61102, n61103, n61104, n61105, n61106,
         n61107, n61108, n61109, n61110, n61111, n61112, n61113, n61114,
         n61115, n61116, n61117, n61118, n61119, n61120, n61121, n61122,
         n61123, n61124, n61125, n61126, n61127, n61128, n61129, n61130,
         n61131, n61132, n61133, n61134, n61135, n61136, n61137, n61138,
         n61139, n61140, n61141, n61142, n61143, n61144, n61145, n61146,
         n61147, n61148, n61149, n61150, n61151, n61152, n61153, n61154,
         n61155, n61156, n61157, n61158, n61159, n61160, n61161, n61162,
         n61163, n61164, n61165, n61166, n61167, n61168, n61169, n61170,
         n61171, n61172, n61173, n61174, n61175, n61176, n61177, n61178,
         n61179, n61180, n61181, n61182, n61183, n61184, n61185, n61186,
         n61187, n61188, n61189, n61190, n61191, n61192, n61193, n61194,
         n61195, n61196, n61197, n61198, n61199, n61200, n61201, n61202,
         n61203, n61204, n61205, n61206, n61207, n61208, n61209, n61210,
         n61211, n61212, n61213, n61214, n61215, n61216, n61217, n61218,
         n61219, n61220, n61221, n61222, n61223, n61224, n61225, n61226,
         n61227, n61228, n61229, n61230, n61231, n61232, n61233, n61234,
         n61235, n61236, n61237, n61238, n61239, n61240, n61241, n61242,
         n61243, n61244, n61245, n61246, n61247, n61248, n61249, n61250,
         n61251, n61252, n61253, n61254, n61255, n61256, n61257, n61258,
         n61259, n61260, n61261, n61262, n61263, n61264, n61265, n61266,
         n61267, n61268, n61269, n61270, n61271, n61272, n61273, n61274,
         n61275, n61276, n61277, n61278, n61279, n61280, n61281, n61282,
         n61283, n61284, n61285, n61286, n61287, n61288, n61289, n61290,
         n61291, n61292, n61293, n61294, n61295, n61296, n61297, n61298,
         n61299, n61300, n61301, n61302, n61303, n61304, n61305, n61306,
         n61307, n61308, n61309, n61310, n61311, n61312, n61313, n61314,
         n61315, n61316, n61317, n61318, n61319, n61320, n61321, n61322,
         n61323, n61324, n61325, n61326, n61327, n61328, n61329, n61330,
         n61331, n61332, n61333, n61334, n61335, n61336, n61337, n61338,
         n61339, n61340, n61341, n61342, n61343, n61344, n61345, n61346,
         n61347, n61348, n61349, n61350, n61351, n61352, n61353, n61354,
         n61355, n61356, n61357, n61358, n61359, n61360, n61361, n61362,
         n61363, n61364, n61365, n61366, n61367, n61368, n61369, n61370,
         n61371, n61372, n61373, n61374, n61375, n61376, n61377, n61378,
         n61379, n61380, n61381, n61382, n61383, n61384, n61385, n61386,
         n61387, n61388, n61389, n61390, n61391, n61392, n61393, n61394,
         n61395, n61396, n61397, n61398, n61399, n61400, n61401, n61402,
         n61403, n61404, n61405, n61406, n61407, n61408, n61409, n61410,
         n61411, n61412, n61413, n61414, n61415, n61416, n61417, n61418,
         n61419, n61420, n61421, n61422, n61423, n61424, n61425, n61426,
         n61427, n61428, n61429, n61430, n61431, n61432, n61433, n61434,
         n61435, n61436, n61437, n61438, n61439, n61440, n61441, n61442,
         n61443, n61444, n61445, n61446, n61447, n61448, n61449, n61450,
         n61451, n61452, n61453, n61454, n61455, n61456, n61457, n61458,
         n61459, n61460, n61461, n61462, n61463, n61464, n61465, n61466,
         n61467, n61468, n61469, n61470, n61471, n61472, n61473, n61474,
         n61475, n61476, n61477, n61478, n61479, n61480, n61481, n61482,
         n61483, n61484, n61485, n61486, n61487, n61488, n61489, n61490,
         n61491, n61492, n61493, n61494, n61495, n61496, n61497, n61498,
         n61499, n61500, n61501, n61502, n61503, n61504, n61505, n61506,
         n61507, n61508, n61509, n61510, n61511, n61512, n61513, n61514,
         n61515, n61516, n61517, n61518, n61519, n61520, n61521, n61522,
         n61523, n61524, n61525, n61526, n61527, n61528, n61529, n61530,
         n61531, n61532, n61533, n61534, n61535, n61536, n61537, n61538,
         n61539, n61540, n61541, n61542, n61543, n61544, n61545, n61546,
         n61547, n61548, n61549, n61550, n61551, n61552, n61553, n61554,
         n61555, n61556, n61557, n61558, n61559, n61560, n61561, n61562,
         n61563, n61564, n61565, n61566, n61567, n61568, n61569, n61570,
         n61571, n61572, n61573, n61574, n61575, n61576, n61577, n61578,
         n61579, n61580, n61581, n61582, n61583, n61584, n61585, n61586,
         n61587, n61588, n61589, n61590, n61591, n61592, n61593, n61594,
         n61595, n61596, n61597, n61598, n61599, n61600, n61601, n61602,
         n61603, n61604, n61605, n61606, n61607, n61608, n61609, n61610,
         n61611, n61612, n61613, n61614, n61615, n61616, n61617, n61618,
         n61619, n61620, n61621, n61622, n61623, n61624, n61625, n61626,
         n61627, n61628, n61629, n61630, n61631, n61632, n61633, n61634,
         n61635, n61636, n61637, n61638, n61639, n61640, n61641, n61642,
         n61643, n61644, n61645, n61646, n61647, n61648, n61649, n61650,
         n61651, n61652, n61653, n61654, n61655, n61656, n61657, n61658,
         n61659, n61660, n61661, n61662, n61663, n61664, n61665, n61666,
         n61667, n61668, n61669, n61670, n61671, n61672, n61673, n61674,
         n61675, n61676, n61677, n61678, n61679, n61680, n61681, n61682,
         n61683, n61684, n61685, n61686, n61687, n61688, n61689, n61690,
         n61691, n61692, n61693, n61694, n61695, n61696, n61697, n61698,
         n61699, n61700, n61701, n61702, n61703, n61704, n61705, n61706,
         n61707, n61708, n61709, n61710, n61711, n61712, n61713, n61714,
         n61715, n61716, n61717, n61718, n61719, n61720, n61721, n61722,
         n61723, n61724, n61725, n61726, n61727, n61728, n61729, n61730,
         n61731, n61732, n61733, n61734, n61735, n61736, n61737, n61738,
         n61739, n61740, n61741, n61742, n61743, n61744, n61745, n61746,
         n61747, n61748, n61749, n61750, n61751, n61752, n61753, n61754,
         n61755, n61756, n61757, n61758, n61759, n61760, n61761, n61762,
         n61763, n61764, n61765, n61766, n61767, n61768, n61769, n61770,
         n61771, n61772, n61773, n61774, n61775, n61776, n61777, n61778,
         n61779, n61780, n61781, n61782, n61783, n61784, n61785, n61786,
         n61787, n61788, n61789, n61790, n61791, n61792, n61793, n61794,
         n61795, n61796, n61797, n61798, n61799, n61800, n61801, n61802,
         n61803, n61804, n61805, n61806, n61807, n61808, n61809, n61810,
         n61811, n61812, n61813, n61814, n61815, n61816, n61817, n61818,
         n61819, n61820, n61821, n61822, n61823, n61824, n61825, n61826,
         n61827, n61828, n61829, n61830, n61831, n61832, n61833, n61834,
         n61835, n61836, n61837, n61838, n61839, n61840, n61841, n61842,
         n61843, n61844, n61845, n61846, n61847, n61848, n61849, n61850,
         n61851, n61852, n61853, n61854, n61855, n61856, n61857, n61858,
         n61859, n61860, n61861, n61862, n61863, n61864, n61865, n61866,
         n61867, n61868, n61869, n61870, n61871, n61872, n61873, n61874,
         n61875, n61876, n61877, n61878, n61879, n61880, n61881, n61882,
         n61883, n61884, n61885, n61886, n61887, n61888, n61889, n61890,
         n61891, n61892, n61893, n61894, n61895, n61896, n61897, n61898,
         n61899, n61900, n61901, n61902, n61903, n61904, n61905, n61906,
         n61907, n61908, n61909, n61910, n61911, n61912, n61913, n61914,
         n61915, n61916, n61917, n61918, n61919, n61920, n61921, n61922,
         n61923, n61924, n61925, n61926, n61927, n61928, n61929, n61930,
         n61931, n61932, n61933, n61934, n61935, n61936, n61937, n61938,
         n61939, n61940, n61941, n61942, n61943, n61944, n61945, n61946,
         n61947, n61948, n61949, n61950, n61951, n61952, n61953, n61954,
         n61955, n61956, n61957, n61958, n61959, n61960, n61961, n61962,
         n61963, n61964, n61965, n61966, n61967, n61968, n61969, n61970,
         n61971, n61972, n61973, n61974, n61975, n61976, n61977, n61978,
         n61979, n61980, n61981, n61982, n61983, n61984, n61985, n61986,
         n61987, n61988, n61989, n61990, n61991, n61992, n61993, n61994,
         n61995, n61996, n61997, n61998, n61999, n62000, n62001, n62002,
         n62003, n62004, n62005, n62006, n62007, n62008, n62009, n62010,
         n62011, n62012, n62013, n62014, n62015, n62016, n62017, n62018,
         n62019, n62020, n62021, n62022, n62023, n62024, n62025, n62026,
         n62027, n62028, n62029, n62030, n62031, n62032, n62033, n62034,
         n62035, n62036, n62037, n62038, n62039, n62040, n62041, n62042,
         n62043, n62044, n62045, n62046, n62047, n62048, n62049, n62050,
         n62051, n62052, n62053, n62054, n62055, n62056, n62057, n62058,
         n62059, n62060, n62061, n62062, n62063, n62064, n62065, n62066,
         n62067, n62068, n62069, n62070, n62071, n62072, n62073, n62074,
         n62075, n62076, n62077, n62078, n62079, n62080, n62081, n62082,
         n62083, n62084, n62085, n62086, n62087, n62088, n62089, n62090,
         n62091, n62092, n62093, n62094, n62095, n62096, n62097, n62098,
         n62099, n62100, n62101, n62102, n62103, n62104, n62105, n62106,
         n62107, n62108, n62109, n62110, n62111, n62112, n62113, n62114,
         n62115, n62116, n62117, n62118, n62119, n62120, n62121, n62122,
         n62123, n62124, n62125, n62126, n62127, n62128, n62129, n62130,
         n62131, n62132, n62133, n62134, n62135, n62136, n62137, n62138,
         n62139, n62140, n62141, n62142, n62143, n62144, n62145, n62146,
         n62147, n62148, n62149, n62150, n62151, n62152, n62153, n62154,
         n62155, n62156, n62157, n62158, n62159, n62160, n62161, n62162,
         n62163, n62164, n62165, n62166, n62167, n62168, n62169, n62170,
         n62171, n62172, n62173, n62174, n62175, n62176, n62177, n62178,
         n62179, n62180, n62181, n62182, n62183, n62184, n62185, n62186,
         n62187, n62188, n62189, n62190, n62191, n62192, n62193, n62194,
         n62195, n62196, n62197, n62198, n62199, n62200, n62201, n62202,
         n62203, n62204, n62205, n62206, n62207, n62208, n62209, n62210,
         n62211, n62212, n62213, n62214, n62215, n62216, n62217, n62218,
         n62219, n62220, n62221, n62222, n62223, n62224, n62225, n62226,
         n62227, n62228, n62229, n62230, n62231, n62232, n62233, n62234,
         n62235, n62236, n62237, n62238, n62239, n62240, n62241, n62242,
         n62243, n62244, n62245, n62246, n62247, n62248, n62249, n62250,
         n62251, n62252, n62253, n62254, n62255, n62256, n62257, n62258,
         n62259, n62260, n62261, n62262, n62263, n62264, n62265, n62266,
         n62267, n62268, n62269, n62270, n62271, n62272, n62273, n62274,
         n62275, n62276, n62277, n62278, n62279, n62280, n62281, n62282,
         n62283, n62284, n62285, n62286, n62287, n62288, n62289, n62290,
         n62291, n62292, n62293, n62294, n62295, n62296, n62297, n62298,
         n62299, n62300, n62301, n62302, n62303, n62304, n62305, n62306,
         n62307, n62308, n62309, n62310, n62311, n62312, n62313, n62314,
         n62315, n62316, n62317, n62318, n62319, n62320, n62321, n62322,
         n62323, n62324, n62325, n62326, n62327, n62328, n62329, n62330,
         n62331, n62332, n62333, n62334, n62335, n62336, n62337, n62338,
         n62339, n62340, n62341, n62342, n62343, n62344, n62345, n62346,
         n62347, n62348, n62349, n62350, n62351, n62352, n62353, n62354,
         n62355, n62356, n62357, n62358, n62359, n62360, n62361, n62362,
         n62363, n62364, n62365, n62366, n62367, n62368, n62369, n62370,
         n62371, n62372, n62373, n62374, n62375, n62376, n62377, n62378,
         n62379, n62380, n62381, n62382, n62383, n62384, n62385, n62386,
         n62387, n62388, n62389, n62390, n62391, n62392, n62393, n62394,
         n62395, n62396, n62397, n62398, n62399, n62400, n62401, n62402,
         n62403, n62404, n62405, n62406, n62407, n62408, n62409, n62410,
         n62411, n62412, n62413, n62414, n62415, n62416, n62417, n62418,
         n62419, n62420, n62421, n62422, n62423, n62424, n62425, n62426,
         n62427, n62428, n62429, n62430, n62431, n62432, n62433, n62434,
         n62435, n62436, n62437, n62438, n62439, n62440, n62441, n62442,
         n62443, n62444, n62445, n62446, n62447, n62448, n62449, n62450,
         n62451, n62452, n62453, n62454, n62455, n62456, n62457, n62458,
         n62459, n62460, n62461, n62462, n62463, n62464, n62465, n62466,
         n62467, n62468, n62469, n62470, n62471, n62472, n62473, n62474,
         n62475, n62476, n62477, n62478, n62479, n62480, n62481, n62482,
         n62483, n62484, n62485, n62486, n62487, n62488, n62489, n62490,
         n62491, n62492, n62493, n62494, n62495, n62496, n62497, n62498,
         n62499, n62500, n62501, n62502, n62503, n62504, n62505, n62506,
         n62507, n62508, n62509, n62510, n62511, n62512, n62513, n62514,
         n62515, n62516, n62517, n62518, n62519, n62520, n62521, n62522,
         n62523, n62524, n62525, n62526, n62527, n62528, n62529, n62530,
         n62531, n62532, n62533, n62534, n62535, n62536, n62537, n62538,
         n62539, n62540, n62541, n62542, n62543, n62544, n62545, n62546,
         n62547, n62548, n62549, n62550, n62551, n62552, n62553, n62554,
         n62555, n62556, n62557, n62558, n62559, n62560, n62561, n62562,
         n62563, n62564, n62565, n62566, n62567, n62568, n62569, n62570,
         n62571, n62572, n62573, n62574, n62575, n62576, n62577, n62578,
         n62579, n62580, n62581, n62582, n62583, n62584, n62585, n62586,
         n62587, n62588, n62589, n62590, n62591, n62592, n62593, n62594,
         n62595, n62596, n62597, n62598, n62599, n62600, n62601, n62602,
         n62603, n62604, n62605, n62606, n62607, n62608, n62609, n62610,
         n62611, n62612, n62613, n62614, n62615, n62616, n62617, n62618,
         n62619, n62620, n62621, n62622, n62623, n62624, n62625, n62626,
         n62627, n62628, n62629, n62630, n62631, n62632, n62633, n62634,
         n62635, n62636, n62637, n62638, n62639, n62640, n62641, n62642,
         n62643, n62644, n62645, n62646, n62647, n62648, n62649, n62650,
         n62651, n62652, n62653, n62654, n62655, n62656, n62657, n62658,
         n62659, n62660, n62661, n62662, n62663, n62664, n62665, n62666,
         n62667, n62668, n62669, n62670, n62671, n62672, n62673, n62674,
         n62675, n62676, n62677, n62678, n62679, n62680, n62681, n62682,
         n62683, n62684, n62685, n62686, n62687, n62688, n62689, n62690,
         n62691, n62692, n62693, n62694, n62695, n62696, n62697, n62698,
         n62699, n62700, n62701, n62702, n62703, n62704, n62705, n62706,
         n62707, n62708, n62709, n62710, n62711, n62712, n62713, n62714,
         n62715, n62716, n62717, n62718, n62719, n62720, n62721, n62722,
         n62723, n62724, n62725, n62726, n62727, n62728, n62729, n62730,
         n62731, n62732, n62733, n62734, n62735, n62736, n62737, n62738,
         n62739, n62740, n62741, n62742, n62743, n62744, n62745, n62746,
         n62747, n62748, n62749, n62750, n62751, n62752, n62753, n62754,
         n62755, n62756, n62757, n62758, n62759, n62760, n62761, n62762,
         n62763, n62764, n62765, n62766, n62767, n62768, n62769, n62770,
         n62771, n62772, n62773, n62774, n62775, n62776, n62777, n62778,
         n62779, n62780, n62781, n62782, n62783, n62784, n62785, n62786,
         n62787, n62788, n62789, n62790, n62791, n62792, n62793, n62794,
         n62795, n62796, n62797, n62798, n62799, n62800, n62801, n62802,
         n62803, n62804, n62805, n62806, n62807, n62808, n62809, n62810,
         n62811, n62812, n62813, n62814, n62815, n62816, n62817, n62818,
         n62819, n62820, n62821, n62822, n62823, n62824, n62825, n62826,
         n62827, n62828, n62829, n62830, n62831, n62832, n62833, n62834,
         n62835, n62836, n62837, n62838, n62839, n62840, n62841, n62842,
         n62843, n62844, n62845, n62846, n62847, n62848, n62849, n62850,
         n62851, n62852, n62853, n62854, n62855, n62856, n62857, n62858,
         n62859, n62860, n62861, n62862, n62863, n62864, n62865, n62866,
         n62867, n62868, n62869, n62870, n62871, n62872, n62873, n62874,
         n62875, n62876, n62877, n62878, n62879, n62880, n62881, n62882,
         n62883, n62884, n62885, n62886, n62887, n62888, n62889, n62890,
         n62891, n62892, n62893, n62894, n62895, n62896, n62897, n62898,
         n62899, n62900, n62901, n62902, n62903, n62904, n62905, n62906,
         n62907, n62908, n62909, n62910, n62911, n62912, n62913, n62914,
         n62915, n62916, n62917, n62918, n62919, n62920, n62921, n62922,
         n62923, n62924, n62925, n62926, n62927, n62928, n62929, n62930,
         n62931, n62932, n62933, n62934, n62935, n62936, n62937, n62938,
         n62939, n62940, n62941, n62942, n62943, n62944, n62945, n62946,
         n62947, n62948, n62949, n62950, n62951, n62952, n62953, n62954,
         n62955, n62956, n62957, n62958, n62959, n62960, n62961, n62962,
         n62963, n62964, n62965, n62966, n62967, n62968, n62969, n62970,
         n62971, n62972, n62973, n62974, n62975, n62976, n62977, n62978,
         n62979, n62980, n62981, n62982, n62983, n62984, n62985, n62986,
         n62987, n62988, n62989, n62990, n62991, n62992, n62993, n62994,
         n62995, n62996, n62997, n62998, n62999, n63000, n63001, n63002,
         n63003, n63004, n63005, n63006, n63007, n63008, n63009, n63010,
         n63011, n63012, n63013, n63014, n63015, n63016, n63017, n63018,
         n63019, n63020, n63021, n63022, n63023, n63024, n63025, n63026,
         n63027, n63028, n63029, n63030, n63031, n63032, n63033, n63034,
         n63035, n63036, n63037, n63038, n63039, n63040, n63041, n63042,
         n63043, n63044, n63045, n63046, n63047, n63048, n63049, n63050,
         n63051, n63052, n63053, n63054, n63055, n63056, n63057, n63058,
         n63059, n63060, n63061, n63062, n63063, n63064, n63065, n63066,
         n63067, n63068, n63069, n63070, n63071, n63072, n63073, n63074,
         n63075, n63076, n63077, n63078, n63079, n63080, n63081, n63082,
         n63083, n63084, n63085, n63086, n63087, n63088, n63089, n63090,
         n63091, n63092, n63093, n63094, n63095, n63096, n63097, n63098,
         n63099, n63100, n63101, n63102, n63103, n63104, n63105, n63106,
         n63107, n63108, n63109, n63110, n63111, n63112, n63113, n63114,
         n63115, n63116, n63117, n63118, n63119, n63120, n63121, n63122,
         n63123, n63124, n63125, n63126, n63127, n63128, n63129, n63130,
         n63131, n63132, n63133, n63134, n63135, n63136, n63137, n63138,
         n63139, n63140, n63141, n63142, n63143, n63144, n63145, n63146,
         n63147, n63148, n63149, n63150, n63151, n63152, n63153, n63154,
         n63155, n63156, n63157, n63158, n63159, n63160, n63161, n63162,
         n63163, n63164, n63165, n63166, n63167, n63168, n63169, n63170,
         n63171, n63172, n63173, n63174, n63175, n63176, n63177, n63178,
         n63179, n63180, n63181, n63182, n63183, n63184, n63185, n63186,
         n63187, n63188, n63189, n63190, n63191, n63192, n63193, n63194,
         n63195, n63196, n63197, n63198, n63199, n63200, n63201, n63202,
         n63203, n63204, n63205, n63206, n63207, n63208, n63209, n63210,
         n63211, n63212, n63213, n63214, n63215, n63216, n63217, n63218,
         n63219, n63220, n63221, n63222, n63223, n63224, n63225, n63226,
         n63227, n63228, n63229, n63230, n63231, n63232, n63233, n63234,
         n63235, n63236, n63237, n63238, n63239, n63240, n63241, n63242,
         n63243, n63244, n63245, n63246, n63247, n63248, n63249, n63250,
         n63251, n63252, n63253, n63254, n63255, n63256, n63257, n63258,
         n63259, n63260, n63261, n63262, n63263, n63264, n63265, n63266,
         n63267, n63268, n63269, n63270, n63271, n63272, n63273, n63274,
         n63275, n63276, n63277, n63278, n63279, n63280, n63281, n63282,
         n63283, n63284, n63285, n63286, n63287, n63288, n63289, n63290,
         n63291, n63292, n63293, n63294, n63295, n63296, n63297, n63298,
         n63299, n63300, n63301, n63302, n63303, n63304, n63305, n63306,
         n63307, n63308, n63309, n63310, n63311, n63312, n63313, n63314,
         n63315, n63316, n63317, n63318, n63319, n63320, n63321, n63322,
         n63323, n63324, n63325, n63326, n63327, n63328, n63329, n63330,
         n63331, n63332, n63333, n63334, n63335, n63336, n63337, n63338,
         n63339, n63340, n63341, n63342, n63343, n63344, n63345, n63346,
         n63347, n63348, n63349, n63350, n63351, n63352, n63353, n63354,
         n63355, n63356, n63357, n63358, n63359, n63360, n63361, n63362,
         n63363, n63364, n63365, n63366, n63367, n63368, n63369, n63370,
         n63371, n63372, n63373, n63374, n63375, n63376, n63377, n63378,
         n63379, n63380, n63381, n63382, n63383, n63384, n63385, n63386,
         n63387, n63388, n63389, n63390, n63391, n63392, n63393, n63394,
         n63395, n63396, n63397, n63398, n63399, n63400, n63401, n63402,
         n63403, n63404, n63405, n63406, n63407, n63408, n63409, n63410,
         n63411, n63412, n63413, n63414, n63415, n63416, n63417, n63418,
         n63419, n63420, n63421, n63422, n63423, n63424, n63425, n63426,
         n63427, n63428, n63429, n63430, n63431, n63432, n63433, n63434,
         n63435, n63436, n63437, n63438, n63439, n63440, n63441, n63442,
         n63443, n63444, n63445, n63446, n63447, n63448, n63449, n63450,
         n63451, n63452, n63453, n63454, n63455, n63456, n63457, n63458,
         n63459, n63460, n63461, n63462, n63463, n63464, n63465, n63466,
         n63467, n63468, n63469, n63470, n63471, n63472, n63473, n63474,
         n63475, n63476, n63477, n63478, n63479, n63480, n63481, n63482,
         n63483, n63484, n63485, n63486, n63487, n63488, n63489, n63490,
         n63491, n63492, n63493, n63494, n63495, n63496, n63497, n63498,
         n63499, n63500, n63501, n63502, n63503, n63504, n63505, n63506,
         n63507, n63508, n63509, n63510, n63511, n63512, n63513, n63514,
         n63515, n63516, n63517, n63518, n63519, n63520, n63521, n63522,
         n63523, n63524, n63525, n63526, n63527, n63528, n63529, n63530,
         n63531, n63532, n63533, n63534, n63535, n63536, n63537, n63538,
         n63539, n63540, n63541, n63542, n63543, n63544, n63545, n63546,
         n63547, n63548, n63549, n63550, n63551, n63552, n63553, n63554,
         n63555, n63556, n63557, n63558, n63559, n63560, n63561, n63562,
         n63563, n63564, n63565, n63566, n63567, n63568, n63569, n63570,
         n63571, n63572, n63573, n63574, n63575, n63576, n63577, n63578,
         n63579, n63580, n63581, n63582, n63583, n63584, n63585, n63586,
         n63587, n63588, n63589, n63590, n63591, n63592, n63593, n63594,
         n63595, n63596, n63597, n63598, n63599, n63600, n63601, n63602,
         n63603, n63604, n63605, n63606, n63607, n63608, n63609, n63610,
         n63611, n63612, n63613, n63614, n63615, n63616, n63617, n63618,
         n63619, n63620, n63621, n63622, n63623, n63624, n63625, n63626,
         n63627, n63628, n63629, n63630, n63631, n63632, n63633, n63634,
         n63635, n63636, n63637, n63638, n63639, n63640, n63641, n63642,
         n63643, n63644, n63645, n63646, n63647, n63648, n63649, n63650,
         n63651, n63652, n63653, n63654, n63655, n63656, n63657, n63658,
         n63659, n63660, n63661, n63662, n63663, n63664, n63665, n63666,
         n63667, n63668, n63669, n63670, n63671, n63672, n63673, n63674,
         n63675, n63676, n63677, n63678, n63679, n63680, n63681, n63682,
         n63683, n63684, n63685, n63686, n63687, n63688, n63689, n63690,
         n63691, n63692, n63693, n63694, n63695, n63696, n63697, n63698,
         n63699, n63700, n63701, n63702, n63703, n63704, n63705, n63706,
         n63707, n63708, n63709, n63710, n63711, n63712, n63713, n63714,
         n63715, n63716, n63717, n63718, n63719, n63720, n63721, n63722,
         n63723, n63724, n63725, n63726, n63727, n63728, n63729, n63730,
         n63731, n63732, n63733, n63734, n63735, n63736, n63737, n63738,
         n63739, n63740, n63741, n63742, n63743, n63744, n63745, n63746,
         n63747, n63748, n63749, n63750, n63751, n63752, n63753, n63754,
         n63755, n63756, n63757, n63758, n63759, n63760, n63761, n63762,
         n63763, n63764, n63765, n63766, n63767, n63768, n63769, n63770,
         n63771, n63772, n63773, n63774, n63775, n63776, n63777, n63778,
         n63779, n63780, n63781, n63782, n63783, n63784, n63785, n63786,
         n63787, n63788, n63789, n63790, n63791, n63792, n63793, n63794,
         n63795, n63796, n63797, n63798, n63799, n63800, n63801, n63802,
         n63803, n63804, n63805, n63806, n63807, n63808, n63809, n63810,
         n63811, n63812, n63813, n63814, n63815, n63816, n63817, n63818,
         n63819, n63820, n63821, n63822, n63823, n63824, n63825, n63826,
         n63827, n63828, n63829, n63830, n63831, n63832, n63833, n63834,
         n63835, n63836, n63837, n63838, n63839, n63840, n63841, n63842,
         n63843, n63844, n63845, n63846, n63847, n63848, n63849, n63850,
         n63851, n63852, n63853, n63854, n63855, n63856, n63857, n63858,
         n63859, n63860, n63861, n63862, n63863, n63864, n63865, n63866,
         n63867, n63868, n63869, n63870, n63871, n63872, n63873, n63874,
         n63875, n63876, n63877, n63878, n63879, n63880, n63881, n63882,
         n63883, n63884, n63885, n63886, n63887, n63888, n63889, n63890,
         n63891, n63892, n63893, n63894, n63895, n63896, n63897, n63898,
         n63899, n63900, n63901, n63902, n63903, n63904, n63905, n63906,
         n63907, n63908, n63909, n63910, n63911, n63912, n63913, n63914,
         n63915, n63916, n63917, n63918, n63919, n63920, n63921, n63922,
         n63923, n63924, n63925, n63926, n63927, n63928, n63929, n63930,
         n63931, n63932, n63933, n63934, n63935, n63936, n63937, n63938,
         n63939, n63940, n63941, n63942, n63943, n63944, n63945, n63946,
         n63947, n63948, n63949, n63950, n63951, n63952, n63953, n63954,
         n63955, n63956, n63957, n63958, n63959, n63960, n63961, n63962,
         n63963, n63964, n63965, n63966, n63967, n63968, n63969, n63970,
         n63971, n63972, n63973, n63974, n63975, n63976, n63977, n63978,
         n63979, n63980, n63981, n63982, n63983, n63984, n63985, n63986,
         n63987, n63988, n63989, n63990, n63991, n63992, n63993, n63994,
         n63995, n63996, n63997, n63998, n63999, n64000, n64001, n64002,
         n64003, n64004, n64005, n64006, n64007, n64008, n64009, n64010,
         n64011, n64012, n64013, n64014, n64015, n64016, n64017, n64018,
         n64019, n64020, n64021, n64022, n64023, n64024, n64025, n64026,
         n64027, n64028, n64029, n64030, n64031, n64032, n64033, n64034,
         n64035, n64036, n64037, n64038, n64039, n64040, n64041, n64042,
         n64043, n64044, n64045, n64046, n64047, n64048, n64049, n64050,
         n64051, n64052, n64053, n64054, n64055, n64056, n64057, n64058,
         n64059, n64060, n64061, n64062, n64063, n64064, n64065, n64066,
         n64067, n64068, n64069, n64070, n64071, n64072, n64073, n64074,
         n64075, n64076, n64077, n64078, n64079, n64080, n64081, n64082,
         n64083, n64084, n64085, n64086, n64087, n64088, n64089, n64090,
         n64091, n64092, n64093, n64094, n64095, n64096, n64097, n64098,
         n64099, n64100, n64101, n64102, n64103, n64104, n64105, n64106,
         n64107, n64108, n64109, n64110, n64111, n64112, n64113, n64114,
         n64115, n64116, n64117, n64118, n64119, n64120, n64121, n64122,
         n64123, n64124, n64125, n64126, n64127, n64128, n64129, n64130,
         n64131, n64132, n64133, n64134, n64135, n64136, n64137, n64138,
         n64139, n64140, n64141, n64142, n64143, n64144, n64145, n64146,
         n64147, n64148, n64149, n64150, n64151, n64152, n64153, n64154,
         n64155, n64156, n64157, n64158, n64159, n64160, n64161, n64162,
         n64163, n64164, n64165, n64166, n64167, n64168, n64169, n64170,
         n64171, n64172, n64173, n64174, n64175, n64176, n64177, n64178,
         n64179, n64180, n64181, n64182, n64183, n64184, n64185, n64186,
         n64187, n64188, n64189, n64190, n64191, n64192, n64193, n64194,
         n64195, n64196, n64197, n64198, n64199, n64200, n64201, n64202,
         n64203, n64204, n64205, n64206, n64207, n64208, n64209, n64210,
         n64211, n64212, n64213, n64214, n64215, n64216, n64217, n64218,
         n64219, n64220, n64221, n64222, n64223, n64224, n64225, n64226,
         n64227, n64228, n64229, n64230, n64231, n64232, n64233, n64234,
         n64235, n64236, n64237, n64238, n64239, n64240, n64241, n64242,
         n64243, n64244, n64245, n64246, n64247, n64248, n64249, n64250,
         n64251, n64252, n64253, n64254, n64255, n64256, n64257, n64258,
         n64259, n64260, n64261, n64262, n64263, n64264, n64265, n64266,
         n64267, n64268, n64269, n64270, n64271, n64272, n64273, n64274,
         n64275, n64276, n64277, n64278, n64279, n64280, n64281, n64282,
         n64283, n64284, n64285, n64286, n64287, n64288, n64289, n64290,
         n64291, n64292, n64293, n64294, n64295, n64296, n64297, n64298,
         n64299, n64300, n64301, n64302, n64303, n64304, n64305, n64306,
         n64307, n64308, n64309, n64310, n64311, n64312, n64313, n64314,
         n64315, n64316, n64317, n64318, n64319, n64320, n64321, n64322,
         n64323, n64324, n64325, n64326, n64327, n64328, n64329, n64330,
         n64331, n64332, n64333, n64334, n64335, n64336, n64337, n64338,
         n64339, n64340, n64341, n64342, n64343, n64344, n64345, n64346,
         n64347, n64348, n64349, n64350, n64351, n64352, n64353, n64354,
         n64355, n64356, n64357, n64358, n64359, n64360, n64361, n64362,
         n64363, n64364, n64365, n64366, n64367, n64368, n64369, n64370,
         n64371, n64372, n64373, n64374, n64375, n64376, n64377, n64378,
         n64379, n64380, n64381, n64382, n64383, n64384, n64385, n64386,
         n64387, n64388, n64389, n64390, n64391, n64392, n64393, n64394,
         n64395, n64396, n64397, n64398, n64399, n64400, n64401, n64402,
         n64403, n64404, n64405, n64406, n64407, n64408, n64409, n64410,
         n64411, n64412, n64413, n64414, n64415, n64416, n64417, n64418,
         n64419, n64420, n64421, n64422, n64423, n64424, n64425, n64426,
         n64427, n64428, n64429, n64430, n64431, n64432, n64433, n64434,
         n64435, n64436, n64437, n64438, n64439, n64440, n64441, n64442,
         n64443, n64444, n64445, n64446, n64447, n64448, n64449, n64450,
         n64451, n64452, n64453, n64454, n64455, n64456, n64457, n64458,
         n64459, n64460, n64461, n64462, n64463, n64464, n64465, n64466,
         n64467, n64468, n64469, n64470, n64471, n64472, n64473, n64474,
         n64475, n64476, n64477, n64478, n64479, n64480, n64481, n64482,
         n64483, n64484, n64485, n64486, n64487, n64488, n64489, n64490,
         n64491, n64492, n64493, n64494, n64495, n64496, n64497, n64498,
         n64499, n64500, n64501, n64502, n64503, n64504, n64505, n64506,
         n64507, n64508, n64509, n64510, n64511, n64512, n64513, n64514,
         n64515, n64516, n64517, n64518, n64519, n64520, n64521, n64522,
         n64523, n64524, n64525, n64526, n64527, n64528, n64529, n64530,
         n64531, n64532, n64533, n64534, n64535, n64536, n64537, n64538,
         n64539, n64540, n64541, n64542, n64543, n64544, n64545, n64546,
         n64547, n64548, n64549, n64550, n64551, n64552, n64553, n64554,
         n64555, n64556, n64557, n64558, n64559, n64560, n64561, n64562,
         n64563, n64564, n64565, n64566, n64567, n64568, n64569, n64570,
         n64571, n64572, n64573, n64574, n64575, n64576, n64577, n64578,
         n64579, n64580, n64581, n64582, n64583, n64584, n64585, n64586,
         n64587, n64588, n64589, n64590, n64591, n64592, n64593, n64594,
         n64595, n64596, n64597, n64598, n64599, n64600, n64601, n64602,
         n64603, n64604, n64605, n64606, n64607, n64608, n64609, n64610,
         n64611, n64612, n64613, n64614, n64615, n64616, n64617, n64618,
         n64619, n64620, n64621, n64622, n64623, n64624, n64625, n64626,
         n64627, n64628, n64629, n64630, n64631, n64632, n64633, n64634,
         n64635, n64636, n64637, n64638, n64639, n64640, n64641, n64642,
         n64643, n64644, n64645, n64646, n64647, n64648, n64649, n64650,
         n64651, n64652, n64653, n64654, n64655, n64656, n64657, n64658,
         n64659, n64660, n64661, n64662, n64663, n64664, n64665, n64666,
         n64667, n64668, n64669, n64670, n64671, n64672, n64673, n64674,
         n64675, n64676, n64677, n64678, n64679, n64680, n64681, n64682,
         n64683, n64684, n64685, n64686, n64687, n64688, n64689, n64690,
         n64691, n64692, n64693, n64694, n64695, n64696, n64697, n64698,
         n64699, n64700, n64701, n64702, n64703, n64704, n64705, n64706,
         n64707, n64708, n64709, n64710, n64711, n64712, n64713, n64714,
         n64715, n64716, n64717, n64718, n64719, n64720, n64721, n64722,
         n64723, n64724, n64725, n64726, n64727, n64728, n64729, n64730,
         n64731, n64732, n64733, n64734, n64735, n64736, n64737, n64738,
         n64739, n64740, n64741, n64742, n64743, n64744, n64745, n64746,
         n64747, n64748, n64749, n64750, n64751, n64752, n64753, n64754,
         n64755, n64756, n64757, n64758, n64759, n64760, n64761, n64762,
         n64763, n64764, n64765, n64766, n64767, n64768, n64769, n64770,
         n64771, n64772, n64773, n64774, n64775, n64776, n64777, n64778,
         n64779, n64780, n64781, n64782, n64783, n64784, n64785, n64786,
         n64787, n64788, n64789, n64790, n64791, n64792, n64793, n64794,
         n64795, n64796, n64797, n64798, n64799, n64800, n64801, n64802,
         n64803, n64804, n64805, n64806, n64807, n64808, n64809, n64810,
         n64811, n64812, n64813, n64814, n64815, n64816, n64817, n64818,
         n64819, n64820, n64821, n64822, n64823, n64824, n64825, n64826,
         n64827, n64828, n64829, n64830, n64831, n64832, n64833, n64834,
         n64835, n64836, n64837, n64838, n64839, n64840, n64841, n64842,
         n64843, n64844, n64845, n64846, n64847, n64848, n64849, n64850,
         n64851, n64852, n64853, n64854, n64855, n64856, n64857, n64858,
         n64859, n64860, n64861, n64862, n64863, n64864, n64865, n64866,
         n64867, n64868, n64869, n64870, n64871, n64872, n64873, n64874,
         n64875, n64876, n64877, n64878, n64879, n64880, n64881, n64882,
         n64883, n64884, n64885, n64886, n64887, n64888, n64889, n64890,
         n64891, n64892, n64893, n64894, n64895, n64896, n64897, n64898,
         n64899, n64900, n64901, n64902, n64903, n64904, n64905, n64906,
         n64907, n64908, n64909, n64910, n64911, n64912, n64913, n64914,
         n64915, n64916, n64917, n64918, n64919, n64920, n64921, n64922,
         n64923, n64924, n64925, n64926, n64927, n64928, n64929, n64930,
         n64931, n64932, n64933, n64934, n64935, n64936, n64937, n64938,
         n64939, n64940, n64941, n64942, n64943, n64944, n64945, n64946,
         n64947, n64948, n64949, n64950, n64951, n64952, n64953, n64954,
         n64955, n64956, n64957, n64958, n64959, n64960, n64961, n64962,
         n64963, n64964, n64965, n64966, n64967, n64968, n64969, n64970,
         n64971, n64972, n64973, n64974, n64975, n64976, n64977, n64978,
         n64979, n64980, n64981, n64982, n64983, n64984, n64985, n64986,
         n64987, n64988, n64989, n64990, n64991, n64992, n64993, n64994,
         n64995, n64996, n64997, n64998, n64999, n65000, n65001, n65002,
         n65003, n65004, n65005, n65006, n65007, n65008, n65009, n65010,
         n65011, n65012, n65013, n65014, n65015, n65016, n65017, n65018,
         n65019, n65020, n65021, n65022, n65023, n65024, n65025, n65026,
         n65027, n65028, n65029, n65030, n65031, n65032, n65033, n65034,
         n65035, n65036, n65037, n65038, n65039, n65040, n65041, n65042,
         n65043, n65044, n65045, n65046, n65047, n65048, n65049, n65050,
         n65051, n65052, n65053, n65054, n65055, n65056, n65057, n65058,
         n65059, n65060, n65061, n65062, n65063, n65064, n65065, n65066,
         n65067, n65068, n65069, n65070, n65071, n65072, n65073, n65074,
         n65075, n65076, n65077, n65078, n65079, n65080, n65081, n65082,
         n65083, n65084, n65085, n65086, n65087, n65088, n65089, n65090,
         n65091, n65092, n65093, n65094, n65095, n65096, n65097, n65098,
         n65099, n65100, n65101, n65102, n65103, n65104, n65105, n65106,
         n65107, n65108, n65109, n65110, n65111, n65112, n65113, n65114,
         n65115, n65116, n65117, n65118, n65119, n65120, n65121, n65122,
         n65123, n65124, n65125, n65126, n65127, n65128, n65129, n65130,
         n65131, n65132, n65133, n65134, n65135, n65136, n65137, n65138,
         n65139, n65140, n65141, n65142, n65143, n65144, n65145, n65146,
         n65147, n65148, n65149, n65150, n65151, n65152, n65153, n65154,
         n65155, n65156, n65157, n65158, n65159, n65160, n65161, n65162,
         n65163, n65164, n65165, n65166, n65167, n65168, n65169, n65170,
         n65171, n65172, n65173, n65174, n65175, n65176, n65177, n65178,
         n65179, n65180, n65181, n65182, n65183, n65184, n65185, n65186,
         n65187, n65188, n65189, n65190, n65191, n65192, n65193, n65194,
         n65195, n65196, n65197, n65198, n65199, n65200, n65201, n65202,
         n65203, n65204, n65205, n65206, n65207, n65208, n65209, n65210,
         n65211, n65212, n65213, n65214, n65215, n65216, n65217, n65218,
         n65219, n65220, n65221, n65222, n65223, n65224, n65225, n65226,
         n65227, n65228, n65229, n65230, n65231, n65232, n65233, n65234,
         n65235, n65236, n65237, n65238, n65239, n65240, n65241, n65242,
         n65243, n65244, n65245, n65246, n65247, n65248, n65249, n65250,
         n65251, n65252, n65253, n65254, n65255, n65256, n65257, n65258,
         n65259, n65260, n65261, n65262, n65263, n65264, n65265, n65266,
         n65267, n65268, n65269, n65270, n65271, n65272, n65273, n65274,
         n65275, n65276, n65277, n65278, n65279, n65280, n65281, n65282,
         n65283, n65284, n65285, n65286, n65287, n65288, n65289, n65290,
         n65291, n65292, n65293, n65294, n65295, n65296, n65297, n65298,
         n65299, n65300, n65301, n65302, n65303, n65304, n65305, n65306,
         n65307, n65308, n65309, n65310, n65311, n65312, n65313, n65314,
         n65315, n65316, n65317, n65318, n65319, n65320, n65321, n65322,
         n65323, n65324, n65325, n65326, n65327, n65328, n65329, n65330,
         n65331, n65332, n65333, n65334, n65335, n65336, n65337, n65338,
         n65339, n65340, n65341, n65342, n65343, n65344, n65345, n65346,
         n65347, n65348, n65349, n65350, n65351, n65352, n65353, n65354,
         n65355, n65356, n65357, n65358, n65359, n65360, n65361, n65362,
         n65363, n65364, n65365, n65366, n65367, n65368, n65369, n65370,
         n65371, n65372, n65373, n65374, n65375, n65376, n65377, n65378,
         n65379, n65380, n65381, n65382, n65383, n65384, n65385, n65386,
         n65387, n65388, n65389, n65390, n65391, n65392, n65393, n65394,
         n65395, n65396, n65397, n65398, n65399, n65400, n65401, n65402,
         n65403, n65404, n65405, n65406, n65407, n65408, n65409, n65410,
         n65411, n65412, n65413, n65414, n65415, n65416, n65417, n65418,
         n65419, n65420, n65421, n65422, n65423, n65424, n65425, n65426,
         n65427, n65428, n65429, n65430, n65431, n65432, n65433, n65434,
         n65435, n65436, n65437, n65438, n65439, n65440, n65441, n65442,
         n65443, n65444, n65445, n65446, n65447, n65448, n65449, n65450,
         n65451, n65452, n65453, n65454, n65455, n65456, n65457, n65458,
         n65459, n65460, n65461, n65462, n65463, n65464, n65465, n65466,
         n65467, n65468, n65469, n65470, n65471, n65472, n65473, n65474,
         n65475, n65476, n65477, n65478, n65479, n65480, n65481, n65482,
         n65483, n65484, n65485, n65486, n65487, n65488, n65489, n65490,
         n65491, n65492, n65493, n65494, n65495, n65496, n65497, n65498,
         n65499, n65500, n65501, n65502, n65503, n65504, n65505, n65506,
         n65507, n65508, n65509, n65510, n65511, n65512, n65513, n65514,
         n65515, n65516, n65517, n65518, n65519, n65520, n65521, n65522,
         n65523, n65524, n65525, n65526, n65527, n65528, n65529, n65530,
         n65531, n65532, n65533, n65534, n65535, n65536, n65537, n65538,
         n65539, n65540, n65541, n65542, n65543, n65544, n65545, n65546,
         n65547, n65548, n65549, n65550, n65551, n65552, n65553, n65554,
         n65555, n65556, n65557, n65558, n65559, n65560, n65561, n65562,
         n65563, n65564, n65565, n65566, n65567, n65568, n65569, n65570,
         n65571, n65572, n65573, n65574, n65575, n65576, n65577, n65578,
         n65579, n65580, n65581, n65582, n65583, n65584, n65585, n65586,
         n65587, n65588, n65589, n65590, n65591, n65592, n65593, n65594,
         n65595, n65596, n65597, n65598, n65599, n65600, n65601, n65602,
         n65603, n65604, n65605, n65606, n65607, n65608, n65609, n65610,
         n65611, n65612, n65613, n65614, n65615, n65616, n65617, n65618,
         n65619, n65620, n65621, n65622, n65623, n65624, n65625, n65626,
         n65627, n65628, n65629, n65630, n65631, n65632, n65633, n65634,
         n65635, n65636, n65637, n65638, n65639, n65640, n65641, n65642,
         n65643, n65644, n65645, n65646, n65647, n65648, n65649, n65650,
         n65651, n65652, n65653, n65654, n65655, n65656, n65657, n65658,
         n65659, n65660, n65661, n65662, n65663, n65664, n65665, n65666,
         n65667, n65668, n65669, n65670, n65671, n65672, n65673, n65674,
         n65675, n65676, n65677, n65678, n65679, n65680, n65681, n65682,
         n65683, n65684, n65685, n65686, n65687, n65688, n65689, n65690,
         n65691, n65692, n65693, n65694, n65695, n65696, n65697, n65698,
         n65699, n65700, n65701, n65702, n65703, n65704, n65705, n65706,
         n65707, n65708, n65709, n65710, n65711, n65712, n65713, n65714,
         n65715, n65716, n65717, n65718, n65719, n65720, n65721, n65722,
         n65723, n65724, n65725, n65726, n65727, n65728, n65729, n65730,
         n65731, n65732, n65733, n65734, n65735, n65736, n65737, n65738,
         n65739, n65740, n65741, n65742, n65743, n65744, n65745, n65746,
         n65747, n65748, n65749, n65750, n65751, n65752, n65753, n65754,
         n65755, n65756, n65757, n65758, n65759, n65760, n65761, n65762,
         n65763, n65764, n65765, n65766, n65767, n65768, n65769, n65770,
         n65771, n65772, n65773, n65774, n65775, n65776, n65777, n65778,
         n65779, n65780, n65781, n65782, n65783, n65784, n65785, n65786,
         n65787, n65788, n65789, n65790, n65791, n65792, n65793, n65794,
         n65795, n65796, n65797, n65798, n65799, n65800, n65801, n65802,
         n65803, n65804, n65805, n65806, n65807, n65808, n65809, n65810,
         n65811, n65812, n65813, n65814, n65815, n65816, n65817, n65818,
         n65819, n65820, n65821, n65822, n65823, n65824, n65825, n65826,
         n65827, n65828, n65829, n65830, n65831, n65832, n65833, n65834,
         n65835, n65836, n65837, n65838, n65839, n65840, n65841, n65842,
         n65843, n65844, n65845, n65846, n65847, n65848, n65849, n65850,
         n65851, n65852, n65853, n65854, n65855, n65856, n65857, n65858,
         n65859, n65860, n65861, n65862, n65863, n65864, n65865, n65866,
         n65867, n65868, n65869, n65870, n65871, n65872, n65873, n65874,
         n65875, n65876, n65877, n65878, n65879, n65880, n65881, n65882,
         n65883, n65884, n65885, n65886, n65887, n65888, n65889, n65890,
         n65891, n65892, n65893, n65894, n65895, n65896, n65897, n65898,
         n65899, n65900, n65901, n65902, n65903, n65904, n65905, n65906,
         n65907, n65908, n65909, n65910, n65911, n65912, n65913, n65914,
         n65915, n65916, n65917, n65918, n65919, n65920, n65921, n65922,
         n65923, n65924, n65925, n65926, n65927, n65928, n65929, n65930,
         n65931, n65932, n65933, n65934, n65935, n65936, n65937, n65938,
         n65939, n65940, n65941, n65942, n65943, n65944, n65945, n65946,
         n65947, n65948, n65949, n65950, n65951, n65952, n65953, n65954,
         n65955, n65956, n65957, n65958, n65959, n65960, n65961, n65962,
         n65963, n65964, n65965, n65966, n65967, n65968, n65969, n65970,
         n65971, n65972, n65973, n65974, n65975, n65976, n65977, n65978,
         n65979, n65980, n65981, n65982, n65983, n65984, n65985, n65986,
         n65987, n65988, n65989, n65990, n65991, n65992, n65993, n65994,
         n65995, n65996, n65997, n65998, n65999, n66000, n66001, n66002,
         n66003, n66004, n66005, n66006, n66007, n66008, n66009, n66010,
         n66011, n66012, n66013, n66014, n66015, n66016, n66017, n66018,
         n66019, n66020, n66021, n66022, n66023, n66024, n66025, n66026,
         n66027, n66028, n66029, n66030, n66031, n66032, n66033, n66034,
         n66035, n66036, n66037, n66038, n66039, n66040, n66041, n66042,
         n66043, n66044, n66045, n66046, n66047, n66048, n66049, n66050,
         n66051, n66052, n66053, n66054, n66055, n66056, n66057, n66058,
         n66059, n66060, n66061, n66062, n66063, n66064, n66065, n66066,
         n66067, n66068, n66069, n66070, n66071, n66072, n66073, n66074,
         n66075, n66076, n66077, n66078, n66079, n66080, n66081, n66082,
         n66083, n66084, n66085, n66086, n66087, n66088, n66089, n66090,
         n66091, n66092, n66093, n66094, n66095, n66096, n66097, n66098,
         n66099, n66100, n66101, n66102, n66103, n66104, n66105, n66106,
         n66107, n66108, n66109, n66110, n66111, n66112, n66113, n66114,
         n66115, n66116, n66117, n66118, n66119, n66120, n66121, n66122,
         n66123, n66124, n66125, n66126, n66127, n66128, n66129, n66130,
         n66131, n66132, n66133, n66134, n66135, n66136, n66137, n66138,
         n66139, n66140, n66141, n66142, n66143, n66144, n66145, n66146,
         n66147, n66148, n66149, n66150, n66151, n66152, n66153, n66154,
         n66155, n66156, n66157, n66158, n66159, n66160, n66161, n66162,
         n66163, n66164, n66165, n66166, n66167, n66168, n66169, n66170,
         n66171, n66172, n66173, n66174, n66175, n66176, n66177, n66178,
         n66179, n66180, n66181, n66182, n66183, n66184, n66185, n66186,
         n66187, n66188, n66189, n66190, n66191, n66192, n66193, n66194,
         n66195, n66196, n66197, n66198, n66199, n66200, n66201, n66202,
         n66203, n66204, n66205, n66206, n66207, n66208, n66209, n66210,
         n66211, n66212, n66213, n66214, n66215, n66216, n66217, n66218,
         n66219, n66220, n66221, n66222, n66223, n66224, n66225, n66226,
         n66227, n66228, n66229, n66230, n66231, n66232, n66233, n66234,
         n66235, n66236, n66237, n66238, n66239, n66240, n66241, n66242,
         n66243, n66244, n66245, n66246, n66247, n66248, n66249, n66250,
         n66251, n66252, n66253, n66254, n66255, n66256, n66257, n66258,
         n66259, n66260, n66261, n66262, n66263, n66264, n66265, n66266,
         n66267, n66268, n66269, n66270, n66271, n66272, n66273, n66274,
         n66275, n66276, n66277, n66278, n66279, n66280, n66281, n66282,
         n66283, n66284, n66285, n66286, n66287, n66288, n66289, n66290,
         n66291, n66292, n66293, n66294, n66295, n66296, n66297, n66298,
         n66299, n66300, n66301, n66302, n66303, n66304, n66305, n66306,
         n66307, n66308, n66309, n66310, n66311, n66312, n66313, n66314,
         n66315, n66316, n66317, n66318, n66319, n66320, n66321, n66322,
         n66323, n66324, n66325, n66326, n66327, n66328, n66329, n66330,
         n66331, n66332, n66333, n66334, n66335, n66336, n66337, n66338,
         n66339, n66340, n66341, n66342, n66343, n66344, n66345, n66346,
         n66347, n66348, n66349, n66350, n66351, n66352, n66353, n66354,
         n66355, n66356, n66357, n66358, n66359, n66360, n66361, n66362,
         n66363, n66364, n66365, n66366, n66367, n66368, n66369, n66370,
         n66371, n66372, n66373, n66374, n66375, n66376, n66377, n66378,
         n66379, n66380, n66381, n66382, n66383, n66384, n66385, n66386,
         n66387, n66388, n66389, n66390, n66391, n66392, n66393, n66394,
         n66395, n66396, n66397, n66398, n66399, n66400, n66401, n66402,
         n66403, n66404, n66405, n66406, n66407, n66408, n66409, n66410,
         n66411, n66412, n66413, n66414, n66415, n66416, n66417, n66418,
         n66419, n66420, n66421, n66422, n66423, n66424, n66425, n66426,
         n66427, n66428, n66429, n66430, n66431, n66432, n66433, n66434,
         n66435, n66436, n66437, n66438, n66439, n66440, n66441, n66442,
         n66443, n66444, n66445, n66446, n66447, n66448, n66449, n66450,
         n66451, n66452, n66453, n66454, n66455, n66456, n66457, n66458,
         n66459, n66460, n66461, n66462, n66463, n66464, n66465, n66466,
         n66467, n66468, n66469, n66470, n66471, n66472, n66473, n66474,
         n66475, n66476, n66477, n66478, n66479, n66480, n66481, n66482,
         n66483, n66484, n66485, n66486, n66487, n66488, n66489, n66490,
         n66491, n66492, n66493, n66494, n66495, n66496, n66497, n66498,
         n66499, n66500, n66501, n66502, n66503, n66504, n66505, n66506,
         n66507, n66508, n66509, n66510, n66511, n66512, n66513, n66514,
         n66515, n66516, n66517, n66518, n66519, n66520, n66521, n66522,
         n66523, n66524, n66525, n66526, n66527, n66528, n66529, n66530,
         n66531, n66532, n66533, n66534, n66535, n66536, n66537, n66538,
         n66539, n66540, n66541, n66542, n66543, n66544, n66545, n66546,
         n66547, n66548, n66549, n66550, n66551, n66552, n66553, n66554,
         n66555, n66556, n66557, n66558, n66559, n66560, n66561, n66562,
         n66563, n66564, n66565, n66566, n66567, n66568, n66569, n66570,
         n66571, n66572, n66573, n66574, n66575, n66576, n66577, n66578,
         n66579, n66580, n66581, n66582, n66583, n66584, n66585, n66586,
         n66587, n66588, n66589, n66590, n66591, n66592, n66593, n66594,
         n66595, n66596, n66597, n66598, n66599, n66600, n66601, n66602,
         n66603, n66604, n66605, n66606, n66607, n66608, n66609, n66610,
         n66611, n66612, n66613, n66614, n66615, n66616, n66617, n66618,
         n66619, n66620, n66621, n66622, n66623, n66624, n66625, n66626,
         n66627, n66628, n66629, n66630, n66631, n66632, n66633, n66634,
         n66635, n66636, n66637, n66638, n66639, n66640, n66641, n66642,
         n66643, n66644, n66645, n66646, n66647, n66648, n66649, n66650,
         n66651, n66652, n66653, n66654, n66655, n66656, n66657, n66658,
         n66659, n66660, n66661, n66662, n66663, n66664, n66665, n66666,
         n66667, n66668, n66669, n66670, n66671, n66672, n66673, n66674,
         n66675, n66676, n66677, n66678, n66679, n66680, n66681, n66682,
         n66683, n66684, n66685, n66686, n66687, n66688, n66689, n66690,
         n66691, n66692, n66693, n66694, n66695, n66696, n66697, n66698,
         n66699, n66700, n66701, n66702, n66703, n66704, n66705, n66706,
         n66707, n66708, n66709, n66710, n66711, n66712, n66713, n66714,
         n66715, n66716, n66717, n66718, n66719, n66720, n66721, n66722,
         n66723, n66724, n66725, n66726, n66727, n66728, n66729, n66730,
         n66731, n66732, n66733, n66734, n66735, n66736, n66737, n66738,
         n66739, n66740, n66741, n66742, n66743, n66744, n66745, n66746,
         n66747, n66748, n66749, n66750, n66751, n66752, n66753, n66754,
         n66755, n66756, n66757, n66758, n66759, n66760, n66761, n66762,
         n66763, n66764, n66765, n66766, n66767, n66768, n66769, n66770,
         n66771, n66772, n66773, n66774, n66775, n66776, n66777, n66778,
         n66779, n66780, n66781, n66782, n66783, n66784, n66785, n66786,
         n66787, n66788, n66789, n66790, n66791, n66792, n66793, n66794,
         n66795, n66796, n66797, n66798, n66799, n66800, n66801, n66802,
         n66803, n66804, n66805, n66806, n66807, n66808, n66809, n66810,
         n66811, n66812, n66813, n66814, n66815, n66816, n66817, n66818,
         n66819, n66820, n66821, n66822, n66823, n66824, n66825, n66826,
         n66827, n66828, n66829, n66830, n66831, n66832, n66833, n66834,
         n66835, n66836, n66837, n66838, n66839, n66840, n66841, n66842,
         n66843, n66844, n66845, n66846, n66847, n66848, n66849, n66850,
         n66851, n66852, n66853, n66854, n66855, n66856, n66857, n66858,
         n66859, n66860, n66861, n66862, n66863, n66864, n66865, n66866,
         n66867, n66868, n66869, n66870, n66871, n66872, n66873, n66874,
         n66875, n66876, n66877, n66878, n66879, n66880, n66881, n66882,
         n66883, n66884, n66885, n66886, n66887, n66888, n66889, n66890,
         n66891, n66892, n66893, n66894, n66895, n66896, n66897, n66898,
         n66899, n66900, n66901, n66902, n66903, n66904, n66905, n66906,
         n66907, n66908, n66909, n66910, n66911, n66912, n66913, n66914,
         n66915, n66916, n66917, n66918, n66919, n66920, n66921, n66922,
         n66923, n66924, n66925, n66926, n66927, n66928, n66929, n66930,
         n66931, n66932, n66933, n66934, n66935, n66936, n66937, n66938,
         n66939, n66940, n66941, n66942, n66943, n66944, n66945, n66946,
         n66947, n66948, n66949, n66950, n66951, n66952, n66953, n66954,
         n66955, n66956, n66957, n66958, n66959, n66960, n66961, n66962,
         n66963, n66964, n66965, n66966, n66967, n66968, n66969, n66970,
         n66971, n66972, n66973, n66974, n66975, n66976, n66977, n66978,
         n66979, n66980, n66981, n66982, n66983, n66984, n66985, n66986,
         n66987, n66988, n66989, n66990, n66991, n66992, n66993, n66994,
         n66995, n66996, n66997, n66998, n66999, n67000, n67001, n67002,
         n67003, n67004, n67005, n67006, n67007, n67008, n67009, n67010,
         n67011, n67012, n67013, n67014, n67015, n67016, n67017, n67018,
         n67019, n67020, n67021, n67022, n67023, n67024, n67025, n67026,
         n67027, n67028, n67029, n67030, n67031, n67032, n67033, n67034,
         n67035, n67036, n67037, n67038, n67039, n67040, n67041, n67042,
         n67043, n67044, n67045, n67046, n67047, n67048, n67049, n67050,
         n67051, n67052, n67053, n67054, n67055, n67056, n67057, n67058,
         n67059, n67060, n67061, n67062, n67063, n67064, n67065, n67066,
         n67067, n67068, n67069, n67070, n67071, n67072, n67073, n67074,
         n67075, n67076, n67077, n67078, n67079, n67080, n67081, n67082,
         n67083, n67084, n67085, n67086, n67087, n67088, n67089, n67090,
         n67091, n67092, n67093, n67094, n67095, n67096, n67097, n67098,
         n67099, n67100, n67101, n67102, n67103, n67104, n67105, n67106,
         n67107, n67108, n67109, n67110, n67111, n67112, n67113, n67114,
         n67115, n67116, n67117, n67118, n67119, n67120, n67121, n67122,
         n67123, n67124, n67125, n67126, n67127, n67128, n67129, n67130,
         n67131, n67132, n67133, n67134, n67135, n67136, n67137, n67138,
         n67139, n67140, n67141, n67142, n67143, n67144, n67145, n67146,
         n67147, n67148, n67149, n67150, n67151, n67152, n67153, n67154,
         n67155, n67156, n67157, n67158, n67159, n67160, n67161, n67162,
         n67163, n67164, n67165, n67166, n67167, n67168, n67169, n67170,
         n67171, n67172, n67173, n67174, n67175, n67176, n67177, n67178,
         n67179, n67180, n67181, n67182, n67183, n67184, n67185, n67186,
         n67187, n67188, n67189, n67190, n67191, n67192, n67193, n67194,
         n67195, n67196, n67197, n67198, n67199, n67200, n67201, n67202,
         n67203, n67204, n67205, n67206, n67207, n67208, n67209, n67210,
         n67211, n67212, n67213, n67214, n67215, n67216, n67217, n67218,
         n67219, n67220, n67221, n67222, n67223, n67224, n67225, n67226,
         n67227, n67228, n67229, n67230, n67231, n67232, n67233, n67234,
         n67235, n67236, n67237, n67238, n67239, n67240, n67241, n67242,
         n67243, n67244, n67245, n67246, n67247, n67248, n67249, n67250,
         n67251, n67252, n67253, n67254, n67255, n67256, n67257, n67258,
         n67259, n67260, n67261, n67262, n67263, n67264, n67265, n67266,
         n67267, n67268, n67269, n67270, n67271, n67272, n67273, n67274,
         n67275, n67276, n67277, n67278, n67279, n67280, n67281, n67282,
         n67283, n67284, n67285, n67286, n67287, n67288, n67289, n67290,
         n67291, n67292, n67293, n67294, n67295, n67296, n67297, n67298,
         n67299, n67300, n67301, n67302, n67303, n67304, n67305, n67306,
         n67307, n67308, n67309, n67310, n67311, n67312, n67313, n67314,
         n67315, n67316, n67317, n67318, n67319, n67320, n67321, n67322,
         n67323, n67324, n67325, n67326, n67327, n67328, n67329, n67330,
         n67331, n67332, n67333, n67334, n67335, n67336, n67337, n67338,
         n67339, n67340, n67341, n67342, n67343, n67344, n67345, n67346,
         n67347, n67348, n67349, n67350, n67351, n67352, n67353, n67354,
         n67355, n67356, n67357, n67358, n67359, n67360, n67361, n67362,
         n67363, n67364, n67365, n67366, n67367, n67368, n67369, n67370,
         n67371, n67372, n67373, n67374, n67375, n67376, n67377, n67378,
         n67379, n67380, n67381, n67382, n67383, n67384, n67385, n67386,
         n67387, n67388, n67389, n67390, n67391, n67392, n67393, n67394,
         n67395, n67396, n67397, n67398, n67399, n67400, n67401, n67402,
         n67403, n67404, n67405, n67406, n67407, n67408, n67409, n67410,
         n67411, n67412, n67413, n67414, n67415, n67416, n67417, n67418,
         n67419, n67420, n67421, n67422, n67423, n67424, n67425, n67426,
         n67427, n67428, n67429, n67430, n67431, n67432, n67433, n67434,
         n67435, n67436, n67437, n67438, n67439, n67440, n67441, n67442,
         n67443, n67444, n67445, n67446, n67447, n67448, n67449, n67450,
         n67451, n67452, n67453, n67454, n67455, n67456, n67457, n67458,
         n67459, n67460, n67461, n67462, n67463, n67464, n67465, n67466,
         n67467, n67468, n67469, n67470, n67471, n67472, n67473, n67474,
         n67475, n67476, n67477, n67478, n67479, n67480, n67481, n67482,
         n67483, n67484, n67485, n67486, n67487, n67488, n67489, n67490,
         n67491, n67492, n67493, n67494, n67495, n67496, n67497, n67498,
         n67499, n67500, n67501, n67502, n67503, n67504, n67505, n67506,
         n67507, n67508, n67509, n67510, n67511, n67512, n67513, n67514,
         n67515, n67516, n67517, n67518, n67519, n67520, n67521, n67522,
         n67523, n67524, n67525, n67526, n67527, n67528, n67529, n67530,
         n67531, n67532, n67533, n67534, n67535, n67536, n67537, n67538,
         n67539, n67540, n67541, n67542, n67543, n67544, n67545, n67546,
         n67547, n67548, n67549, n67550, n67551, n67552, n67553, n67554,
         n67555, n67556, n67557, n67558, n67559, n67560, n67561, n67562,
         n67563, n67564, n67565, n67566, n67567, n67568, n67569, n67570,
         n67571, n67572, n67573, n67574, n67575, n67576, n67577, n67578,
         n67579, n67580, n67581, n67582, n67583, n67584, n67585, n67586,
         n67587, n67588, n67589, n67590, n67591, n67592, n67593, n67594,
         n67595, n67596, n67597, n67598, n67599, n67600, n67601, n67602,
         n67603, n67604, n67605, n67606, n67607, n67608, n67609, n67610,
         n67611, n67612, n67613, n67614, n67615, n67616, n67617, n67618,
         n67619, n67620, n67621, n67622, n67623, n67624, n67625, n67626,
         n67627, n67628, n67629, n67630, n67631, n67632, n67633, n67634,
         n67635, n67636, n67637, n67638, n67639, n67640, n67641, n67642,
         n67643, n67644, n67645, n67646, n67647, n67648, n67649, n67650,
         n67651, n67652, n67653, n67654, n67655, n67656, n67657, n67658,
         n67659, n67660, n67661, n67662, n67663, n67664, n67665, n67666,
         n67667, n67668, n67669, n67670, n67671, n67672, n67673, n67674,
         n67675, n67676, n67677, n67678, n67679, n67680, n67681, n67682,
         n67683, n67684, n67685, n67686, n67687, n67688, n67689, n67690,
         n67691, n67692, n67693, n67694, n67695, n67696, n67697, n67698,
         n67699, n67700, n67701, n67702, n67703, n67704, n67705, n67706,
         n67707, n67708, n67709, n67710, n67711, n67712, n67713, n67714,
         n67715, n67716, n67717, n67718, n67719, n67720, n67721, n67722,
         n67723, n67724, n67725, n67726, n67727, n67728, n67729, n67730,
         n67731, n67732, n67733, n67734, n67735, n67736, n67737, n67738,
         n67739, n67740, n67741, n67742, n67743, n67744, n67745, n67746,
         n67747, n67748, n67749, n67750, n67751, n67752, n67753, n67754,
         n67755, n67756, n67757, n67758, n67759, n67760, n67761, n67762,
         n67763, n67764, n67765, n67766, n67767, n67768, n67769, n67770,
         n67771, n67772, n67773, n67774, n67775, n67776, n67777, n67778,
         n67779, n67780, n67781, n67782, n67783, n67784, n67785, n67786,
         n67787, n67788, n67789, n67790, n67791, n67792, n67793, n67794,
         n67795, n67796, n67797, n67798, n67799, n67800, n67801, n67802,
         n67803, n67804, n67805, n67806, n67807, n67808, n67809, n67810,
         n67811, n67812, n67813, n67814, n67815, n67816, n67817, n67818,
         n67819, n67820, n67821, n67822, n67823, n67824, n67825, n67826,
         n67827, n67828, n67829, n67830, n67831, n67832, n67833, n67834,
         n67835, n67836, n67837, n67838, n67839, n67840, n67841, n67842,
         n67843, n67844, n67845, n67846, n67847, n67848, n67849, n67850,
         n67851, n67852, n67853, n67854, n67855, n67856, n67857, n67858,
         n67859, n67860, n67861, n67862, n67863, n67864, n67865, n67866,
         n67867, n67868, n67869, n67870, n67871, n67872, n67873, n67874,
         n67875, n67876, n67877, n67878, n67879, n67880, n67881, n67882,
         n67883, n67884, n67885, n67886, n67887, n67888, n67889, n67890,
         n67891, n67892, n67893, n67894, n67895, n67896, n67897, n67898,
         n67899, n67900, n67901, n67902, n67903, n67904, n67905, n67906,
         n67907, n67908, n67909, n67910, n67911, n67912, n67913, n67914,
         n67915, n67916, n67917, n67918, n67919, n67920, n67921, n67922,
         n67923, n67924, n67925, n67926, n67927, n67928, n67929, n67930,
         n67931, n67932, n67933, n67934, n67935, n67936, n67937, n67938,
         n67939, n67940, n67941, n67942, n67943, n67944, n67945, n67946,
         n67947, n67948, n67949, n67950, n67951, n67952, n67953, n67954,
         n67955, n67956, n67957, n67958, n67959, n67960, n67961, n67962,
         n67963, n67964, n67965, n67966, n67967, n67968, n67969, n67970,
         n67971, n67972, n67973, n67974, n67975, n67976, n67977, n67978,
         n67979, n67980, n67981, n67982, n67983, n67984, n67985, n67986,
         n67987, n67988, n67989, n67990, n67991, n67992, n67993, n67994,
         n67995, n67996, n67997, n67998, n67999, n68000, n68001, n68002,
         n68003, n68004, n68005, n68006, n68007, n68008, n68009, n68010,
         n68011, n68012, n68013, n68014, n68015, n68016, n68017, n68018,
         n68019, n68020, n68021, n68022, n68023, n68024, n68025, n68026,
         n68027, n68028, n68029, n68030, n68031, n68032, n68033, n68034,
         n68035, n68036, n68037, n68038, n68039, n68040, n68041, n68042,
         n68043, n68044, n68045, n68046, n68047, n68048, n68049, n68050,
         n68051, n68052, n68053, n68054, n68055, n68056, n68057, n68058,
         n68059, n68060, n68061, n68062, n68063, n68064, n68065, n68066,
         n68067, n68068, n68069, n68070, n68071, n68072, n68073, n68074,
         n68075, n68076, n68077, n68078, n68079, n68080, n68081, n68082,
         n68083, n68084, n68085, n68086, n68087, n68088, n68089, n68090,
         n68091, n68092, n68093, n68094, n68095, n68096, n68097, n68098,
         n68099, n68100, n68101, n68102, n68103, n68104, n68105, n68106,
         n68107, n68108, n68109, n68110, n68111, n68112, n68113, n68114,
         n68115, n68116, n68117, n68118, n68119, n68120, n68121, n68122,
         n68123, n68124, n68125, n68126, n68127, n68128, n68129, n68130,
         n68131, n68132, n68133, n68134, n68135, n68136, n68137, n68138,
         n68139, n68140, n68141, n68142, n68143, n68144, n68145, n68146,
         n68147, n68148, n68149, n68150, n68151, n68152, n68153, n68154,
         n68155, n68156, n68157, n68158, n68159, n68160, n68161, n68162,
         n68163, n68164, n68165, n68166, n68167, n68168, n68169, n68170,
         n68171, n68172, n68173, n68174, n68175, n68176, n68177, n68178,
         n68179, n68180, n68181, n68182, n68183, n68184, n68185, n68186,
         n68187, n68188, n68189, n68190, n68191, n68192, n68193, n68194,
         n68195, n68196, n68197, n68198, n68199, n68200, n68201, n68202,
         n68203, n68204, n68205, n68206, n68207, n68208, n68209, n68210,
         n68211, n68212, n68213, n68214, n68215, n68216, n68217, n68218,
         n68219, n68220, n68221, n68222, n68223, n68224, n68225, n68226,
         n68227, n68228, n68229, n68230, n68231, n68232, n68233, n68234,
         n68235, n68236, n68237, n68238, n68239, n68240, n68241, n68242,
         n68243, n68244, n68245, n68246, n68247, n68248, n68249, n68250,
         n68251, n68252, n68253, n68254, n68255, n68256, n68257, n68258,
         n68259, n68260, n68261, n68262, n68263, n68264, n68265, n68266,
         n68267, n68268, n68269, n68270, n68271, n68272, n68273, n68274,
         n68275, n68276, n68277, n68278, n68279, n68280, n68281, n68282,
         n68283, n68284, n68285, n68286, n68287, n68288, n68289, n68290,
         n68291, n68292, n68293, n68294, n68295, n68296, n68297, n68298,
         n68299, n68300, n68301, n68302, n68303, n68304, n68305, n68306,
         n68307, n68308, n68309, n68310, n68311, n68312, n68313, n68314,
         n68315, n68316, n68317, n68318, n68319, n68320, n68321, n68322,
         n68323, n68324, n68325, n68326, n68327, n68328, n68329, n68330,
         n68331, n68332, n68333, n68334, n68335, n68336, n68337, n68338,
         n68339, n68340, n68341, n68342, n68343, n68344, n68345, n68346,
         n68347, n68348, n68349, n68350, n68351, n68352, n68353, n68354,
         n68355, n68356, n68357, n68358, n68359, n68360, n68361, n68362,
         n68363, n68364, n68365, n68366, n68367, n68368, n68369, n68370,
         n68371, n68372, n68373, n68374, n68375, n68376, n68377, n68378,
         n68379, n68380, n68381, n68382, n68383, n68384, n68385, n68386,
         n68387, n68388, n68389, n68390, n68391, n68392, n68393, n68394,
         n68395, n68396, n68397, n68398, n68399, n68400, n68401, n68402,
         n68403, n68404, n68405, n68406, n68407, n68408, n68409, n68410,
         n68411, n68412, n68413, n68414, n68415, n68416, n68417, n68418,
         n68419, n68420, n68421, n68422, n68423, n68424, n68425, n68426,
         n68427, n68428, n68429, n68430, n68431, n68432, n68433, n68434,
         n68435, n68436, n68437, n68438, n68439, n68440, n68441, n68442,
         n68443, n68444, n68445, n68446, n68447, n68448, n68449, n68450,
         n68451, n68452, n68453, n68454, n68455, n68456, n68457, n68458,
         n68459, n68460, n68461, n68462, n68463, n68464, n68465, n68466,
         n68467, n68468, n68469, n68470, n68471, n68472, n68473, n68474,
         n68475, n68476, n68477, n68478, n68479, n68480, n68481, n68482,
         n68483, n68484, n68485, n68486, n68487, n68488, n68489, n68490,
         n68491, n68492, n68493, n68494, n68495, n68496, n68497, n68498,
         n68499, n68500, n68501, n68502, n68503, n68504, n68505, n68506,
         n68507, n68508, n68509, n68510, n68511, n68512, n68513, n68514,
         n68515, n68516, n68517, n68518, n68519, n68520, n68521, n68522,
         n68523, n68524, n68525, n68526, n68527, n68528, n68529, n68530,
         n68531, n68532, n68533, n68534, n68535, n68536, n68537, n68538,
         n68539, n68540, n68541, n68542, n68543, n68544, n68545, n68546,
         n68547, n68548, n68549, n68550, n68551, n68552, n68553, n68554,
         n68555, n68556, n68557, n68558, n68559, n68560, n68561, n68562,
         n68563, n68564, n68565, n68566, n68567, n68568, n68569, n68570,
         n68571, n68572, n68573, n68574, n68575, n68576, n68577, n68578,
         n68579, n68580, n68581, n68582, n68583, n68584, n68585, n68586,
         n68587, n68588, n68589, n68590, n68591, n68592, n68593, n68594,
         n68595, n68596, n68597, n68598, n68599, n68600, n68601, n68602,
         n68603, n68604, n68605, n68606, n68607, n68608, n68609, n68610,
         n68611, n68612, n68613, n68614, n68615, n68616, n68617, n68618,
         n68619, n68620, n68621, n68622, n68623, n68624, n68625, n68626,
         n68627, n68628, n68629, n68630, n68631, n68632, n68633, n68634,
         n68635, n68636, n68637, n68638, n68639, n68640, n68641, n68642,
         n68643, n68644, n68645, n68646, n68647, n68648, n68649, n68650,
         n68651, n68652, n68653, n68654, n68655, n68656, n68657, n68658,
         n68659, n68660, n68661, n68662, n68663, n68664, n68665, n68666,
         n68667, n68668, n68669, n68670, n68671, n68672, n68673, n68674,
         n68675, n68676, n68677, n68678, n68679, n68680, n68681, n68682,
         n68683, n68684, n68685, n68686, n68687, n68688, n68689, n68690,
         n68691, n68692, n68693, n68694, n68695, n68696, n68697, n68698,
         n68699, n68700, n68701, n68702, n68703, n68704, n68705, n68706,
         n68707, n68708, n68709, n68710, n68711, n68712, n68713, n68714,
         n68715, n68716, n68717, n68718, n68719, n68720, n68721, n68722,
         n68723, n68724, n68725, n68726, n68727, n68728, n68729, n68730,
         n68731, n68732, n68733, n68734, n68735, n68736, n68737, n68738,
         n68739, n68740, n68741, n68742, n68743, n68744, n68745, n68746,
         n68747, n68748, n68749, n68750, n68751, n68752, n68753, n68754,
         n68755, n68756, n68757, n68758, n68759, n68760, n68761, n68762,
         n68763, n68764, n68765, n68766, n68767, n68768, n68769, n68770,
         n68771, n68772, n68773, n68774, n68775, n68776, n68777, n68778,
         n68779, n68780, n68781, n68782, n68783, n68784, n68785, n68786,
         n68787, n68788, n68789, n68790, n68791, n68792, n68793, n68794,
         n68795, n68796, n68797, n68798, n68799, n68800, n68801, n68802,
         n68803, n68804, n68805, n68806, n68807, n68808, n68809, n68810,
         n68811, n68812, n68813, n68814, n68815, n68816, n68817, n68818,
         n68819, n68820, n68821, n68822, n68823, n68824, n68825, n68826,
         n68827, n68828, n68829, n68830, n68831, n68832, n68833, n68834,
         n68835, n68836, n68837, n68838, n68839, n68840, n68841, n68842,
         n68843, n68844, n68845, n68846, n68847, n68848, n68849, n68850,
         n68851, n68852, n68853, n68854, n68855, n68856, n68857, n68858,
         n68859, n68860, n68861, n68862, n68863, n68864, n68865, n68866,
         n68867, n68868, n68869, n68870, n68871, n68872, n68873, n68874,
         n68875, n68876, n68877, n68878, n68879, n68880, n68881, n68882,
         n68883, n68884, n68885, n68886, n68887, n68888, n68889, n68890,
         n68891, n68892, n68893, n68894, n68895, n68896, n68897, n68898,
         n68899, n68900, n68901, n68902, n68903, n68904, n68905, n68906,
         n68907, n68908, n68909, n68910, n68911, n68912, n68913, n68914,
         n68915, n68916, n68917, n68918, n68919, n68920, n68921, n68922,
         n68923, n68924, n68925, n68926, n68927, n68928, n68929, n68930,
         n68931, n68932, n68933, n68934, n68935, n68936, n68937, n68938,
         n68939, n68940, n68941, n68942, n68943, n68944, n68945, n68946,
         n68947, n68948, n68949, n68950, n68951, n68952, n68953, n68954,
         n68955, n68956, n68957, n68958, n68959, n68960, n68961, n68962,
         n68963, n68964, n68965, n68966, n68967, n68968, n68969, n68970,
         n68971, n68972, n68973, n68974, n68975, n68976, n68977, n68978,
         n68979, n68980, n68981, n68982, n68983, n68984, n68985, n68986,
         n68987, n68988, n68989, n68990, n68991, n68992, n68993, n68994,
         n68995, n68996, n68997, n68998, n68999, n69000, n69001, n69002,
         n69003, n69004, n69005, n69006, n69007, n69008, n69009, n69010,
         n69011, n69012, n69013, n69014, n69015, n69016, n69017, n69018,
         n69019, n69020, n69021, n69022, n69023, n69024, n69025, n69026,
         n69027, n69028, n69029, n69030, n69031, n69032, n69033, n69034,
         n69035, n69036, n69037, n69038, n69039, n69040, n69041, n69042,
         n69043, n69044, n69045, n69046, n69047, n69048, n69049, n69050,
         n69051, n69052, n69053, n69054, n69055, n69056, n69057, n69058,
         n69059, n69060, n69061, n69062, n69063, n69064, n69065, n69066,
         n69067, n69068, n69069, n69070, n69071, n69072, n69073, n69074,
         n69075, n69076, n69077, n69078, n69079, n69080, n69081, n69082,
         n69083, n69084, n69085, n69086, n69087, n69088, n69089, n69090,
         n69091, n69092, n69093, n69094, n69095, n69096, n69097, n69098,
         n69099, n69100, n69101, n69102, n69103, n69104, n69105, n69106,
         n69107, n69108, n69109, n69110, n69111, n69112, n69113, n69114,
         n69115, n69116, n69117, n69118, n69119, n69120, n69121, n69122,
         n69123, n69124, n69125, n69126, n69127, n69128, n69129, n69130,
         n69131, n69132, n69133, n69134, n69135, n69136, n69137, n69138,
         n69139, n69140, n69141, n69142, n69143, n69144, n69145, n69146,
         n69147, n69148, n69149, n69150, n69151, n69152, n69153, n69154,
         n69155, n69156, n69157, n69158, n69159, n69160, n69161, n69162,
         n69163, n69164, n69165, n69166, n69167, n69168, n69169, n69170,
         n69171, n69172, n69173, n69174, n69175, n69176, n69177, n69178,
         n69179, n69180, n69181, n69182, n69183, n69184, n69185, n69186,
         n69187, n69188, n69189, n69190, n69191, n69192, n69193, n69194,
         n69195, n69196, n69197, n69198, n69199, n69200, n69201, n69202,
         n69203, n69204, n69205, n69206, n69207, n69208, n69209, n69210,
         n69211, n69212, n69213, n69214, n69215, n69216, n69217, n69218,
         n69219, n69220, n69221, n69222, n69223, n69224, n69225, n69226,
         n69227, n69228, n69229, n69230, n69231, n69232, n69233, n69234,
         n69235, n69236, n69237, n69238, n69239, n69240, n69241, n69242,
         n69243, n69244, n69245, n69246, n69247, n69248, n69249, n69250,
         n69251, n69252, n69253, n69254, n69255, n69256, n69257, n69258,
         n69259, n69260, n69261, n69262, n69263, n69264, n69265, n69266,
         n69267, n69268, n69269, n69270, n69271, n69272, n69273, n69274,
         n69275, n69276, n69277, n69278, n69279, n69280, n69281, n69282,
         n69283, n69284, n69285, n69286, n69287, n69288, n69289, n69290,
         n69291, n69292, n69293, n69294, n69295, n69296, n69297, n69298,
         n69299, n69300, n69301, n69302, n69303, n69304, n69305, n69306,
         n69307, n69308, n69309, n69310, n69311, n69312, n69313, n69314,
         n69315, n69316, n69317, n69318, n69319, n69320, n69321, n69322,
         n69323, n69324, n69325, n69326, n69327, n69328, n69329, n69330,
         n69331, n69332, n69333, n69334, n69335, n69336, n69337, n69338,
         n69339, n69340, n69341, n69342, n69343, n69344, n69345, n69346,
         n69347, n69348, n69349, n69350, n69351, n69352, n69353, n69354,
         n69355, n69356, n69357, n69358, n69359, n69360, n69361, n69362,
         n69363, n69364, n69365, n69366, n69367, n69368, n69369, n69370,
         n69371, n69372, n69373, n69374, n69375, n69376, n69377, n69378,
         n69379, n69380, n69381, n69382, n69383, n69384, n69385, n69386,
         n69387, n69388, n69389, n69390, n69391, n69392, n69393, n69394,
         n69395, n69396, n69397, n69398, n69399, n69400, n69401, n69402,
         n69403, n69404, n69405, n69406, n69407, n69408, n69409, n69410,
         n69411, n69412, n69413, n69414, n69415, n69416, n69417, n69418,
         n69419, n69420, n69421, n69422, n69423, n69424, n69425, n69426,
         n69427, n69428, n69429, n69430, n69431, n69432, n69433, n69434,
         n69435, n69436, n69437, n69438, n69439, n69440, n69441, n69442,
         n69443, n69444, n69445, n69446, n69447, n69448, n69449, n69450,
         n69451, n69452, n69453, n69454, n69455, n69456, n69457, n69458,
         n69459, n69460, n69461, n69462, n69463, n69464, n69465, n69466,
         n69467, n69468, n69469, n69470, n69471, n69472, n69473, n69474,
         n69475, n69476, n69477, n69478, n69479, n69480, n69481, n69482,
         n69483, n69484, n69485, n69486, n69487, n69488, n69489, n69490,
         n69491, n69492, n69493, n69494, n69495, n69496, n69497, n69498,
         n69499, n69500, n69501, n69502, n69503, n69504, n69505, n69506,
         n69507, n69508, n69509, n69510, n69511, n69512, n69513, n69514,
         n69515, n69516, n69517, n69518, n69519, n69520, n69521, n69522,
         n69523, n69524, n69525, n69526, n69527, n69528, n69529, n69530,
         n69531, n69532, n69533, n69534, n69535, n69536, n69537, n69538,
         n69539, n69540, n69541, n69542, n69543, n69544, n69545, n69546,
         n69547, n69548, n69549, n69550, n69551, n69552, n69553, n69554,
         n69555, n69556, n69557, n69558, n69559, n69560, n69561, n69562,
         n69563, n69564, n69565, n69566, n69567, n69568, n69569, n69570,
         n69571, n69572, n69573, n69574, n69575, n69576, n69577, n69578,
         n69579, n69580, n69581, n69582, n69583, n69584, n69585, n69586,
         n69587, n69588, n69589, n69590, n69591, n69592, n69593, n69594,
         n69595, n69596, n69597, n69598, n69599, n69600, n69601, n69602,
         n69603, n69604, n69605, n69606, n69607, n69608, n69609, n69610,
         n69611, n69612, n69613, n69614, n69615, n69616, n69617, n69618,
         n69619, n69620, n69621, n69622, n69623, n69624, n69625, n69626,
         n69627, n69628, n69629, n69630, n69631, n69632, n69633, n69634,
         n69635, n69636, n69637, n69638, n69639, n69640, n69641, n69642,
         n69643, n69644, n69645, n69646, n69647, n69648, n69649, n69650,
         n69651, n69652, n69653, n69654, n69655, n69656, n69657, n69658,
         n69659, n69660, n69661, n69662, n69663, n69664, n69665, n69666,
         n69667, n69668, n69669, n69670, n69671, n69672, n69673, n69674,
         n69675, n69676, n69677, n69678, n69679, n69680, n69681, n69682,
         n69683, n69684, n69685, n69686, n69687, n69688, n69689, n69690,
         n69691, n69692, n69693, n69694, n69695, n69696, n69697, n69698,
         n69699, n69700, n69701, n69702, n69703, n69704, n69705, n69706,
         n69707, n69708, n69709, n69710, n69711, n69712, n69713, n69714,
         n69715, n69716, n69717, n69718, n69719, n69720, n69721, n69722,
         n69723, n69724, n69725, n69726, n69727, n69728, n69729, n69730,
         n69731, n69732, n69733, n69734, n69735, n69736, n69737, n69738,
         n69739, n69740, n69741, n69742, n69743, n69744, n69745, n69746,
         n69747, n69748, n69749, n69750, n69751, n69752, n69753, n69754,
         n69755, n69756, n69757, n69758, n69759, n69760, n69761, n69762,
         n69763, n69764, n69765, n69766, n69767, n69768, n69769, n69770,
         n69771, n69772, n69773, n69774, n69775, n69776, n69777, n69778,
         n69779, n69780, n69781, n69782, n69783, n69784, n69785, n69786,
         n69787, n69788, n69789, n69790, n69791, n69792, n69793, n69794,
         n69795, n69796, n69797, n69798, n69799, n69800, n69801, n69802,
         n69803, n69804, n69805, n69806, n69807, n69808, n69809, n69810,
         n69811, n69812, n69813, n69814, n69815, n69816, n69817, n69818,
         n69819, n69820, n69821, n69822, n69823, n69824, n69825, n69826,
         n69827, n69828, n69829, n69830, n69831, n69832, n69833, n69834,
         n69835, n69836, n69837, n69838, n69839, n69840, n69841, n69842,
         n69843, n69844, n69845, n69846, n69847, n69848, n69849, n69850,
         n69851, n69852, n69853, n69854, n69855, n69856, n69857, n69858,
         n69859, n69860, n69861, n69862, n69863, n69864, n69865, n69866,
         n69867, n69868, n69869, n69870, n69871, n69872, n69873, n69874,
         n69875, n69876, n69877, n69878, n69879, n69880, n69881, n69882,
         n69883, n69884, n69885, n69886, n69887, n69888, n69889, n69890,
         n69891, n69892, n69893, n69894, n69895, n69896, n69897, n69898,
         n69899, n69900, n69901, n69902, n69903, n69904, n69905, n69906,
         n69907, n69908, n69909, n69910, n69911, n69912, n69913, n69914,
         n69915, n69916, n69917, n69918, n69919, n69920, n69921, n69922,
         n69923, n69924, n69925, n69926, n69927, n69928, n69929, n69930,
         n69931, n69932, n69933, n69934, n69935, n69936, n69937, n69938,
         n69939, n69940, n69941, n69942, n69943, n69944, n69945, n69946,
         n69947, n69948, n69949, n69950, n69951, n69952, n69953, n69954,
         n69955, n69956, n69957, n69958, n69959, n69960, n69961, n69962,
         n69963, n69964, n69965, n69966, n69967, n69968, n69969, n69970,
         n69971, n69972, n69973, n69974, n69975, n69976, n69977, n69978,
         n69979, n69980, n69981, n69982, n69983, n69984, n69985, n69986,
         n69987, n69988, n69989, n69990, n69991, n69992, n69993, n69994,
         n69995, n69996, n69997, n69998, n69999, n70000, n70001, n70002,
         n70003, n70004, n70005, n70006, n70007, n70008, n70009, n70010,
         n70011, n70012, n70013, n70014, n70015, n70016, n70017, n70018,
         n70019, n70020, n70021, n70022, n70023, n70024, n70025, n70026,
         n70027, n70028, n70029, n70030, n70031, n70032, n70033, n70034,
         n70035, n70036, n70037, n70038, n70039, n70040, n70041, n70042,
         n70043, n70044, n70045, n70046, n70047, n70048, n70049, n70050,
         n70051, n70052, n70053, n70054, n70055, n70056, n70057, n70058,
         n70059, n70060, n70061, n70062, n70063, n70064, n70065, n70066,
         n70067, n70068, n70069, n70070, n70071, n70072, n70073, n70074,
         n70075, n70076, n70077, n70078, n70079, n70080, n70081, n70082,
         n70083, n70084, n70085, n70086, n70087, n70088, n70089, n70090,
         n70091, n70092, n70093, n70094, n70095, n70096, n70097, n70098,
         n70099, n70100, n70101, n70102, n70103, n70104, n70105, n70106,
         n70107, n70108, n70109, n70110, n70111, n70112, n70113, n70114,
         n70115, n70116, n70117, n70118, n70119, n70120, n70121, n70122,
         n70123, n70124, n70125, n70126, n70127, n70128, n70129, n70130,
         n70131, n70132, n70133, n70134, n70135, n70136, n70137, n70138,
         n70139, n70140, n70141, n70142, n70143, n70144, n70145, n70146,
         n70147, n70148, n70149, n70150, n70151, n70152, n70153, n70154,
         n70155, n70156, n70157, n70158, n70159, n70160, n70161, n70162,
         n70163, n70164, n70165, n70166, n70167, n70168, n70169, n70170,
         n70171, n70172, n70173, n70174, n70175, n70176, n70177, n70178,
         n70179, n70180, n70181, n70182, n70183, n70184, n70185, n70186,
         n70187, n70188, n70189, n70190, n70191, n70192, n70193, n70194,
         n70195, n70196, n70197, n70198, n70199, n70200, n70201, n70202,
         n70203, n70204, n70205, n70206, n70207, n70208, n70209, n70210,
         n70211, n70212, n70213, n70214, n70215, n70216, n70217, n70218,
         n70219, n70220, n70221, n70222, n70223, n70224, n70225, n70226,
         n70227, n70228, n70229, n70230, n70231, n70232, n70233, n70234,
         n70235, n70236, n70237, n70238, n70239, n70240, n70241, n70242,
         n70243, n70244, n70245, n70246, n70247, n70248, n70249, n70250,
         n70251, n70252, n70253, n70254, n70255, n70256, n70257, n70258,
         n70259, n70260, n70261, n70262, n70263, n70264, n70265, n70266,
         n70267, n70268, n70269, n70270, n70271, n70272, n70273, n70274,
         n70275, n70276, n70277, n70278, n70279, n70280, n70281, n70282,
         n70283, n70284, n70285, n70286, n70287, n70288, n70289, n70290,
         n70291, n70292, n70293, n70294, n70295, n70296, n70297, n70298,
         n70299, n70300, n70301, n70302, n70303, n70304, n70305, n70306,
         n70307, n70308, n70309, n70310, n70311, n70312, n70313, n70314,
         n70315, n70316, n70317, n70318, n70319, n70320, n70321, n70322,
         n70323, n70324, n70325, n70326, n70327, n70328, n70329, n70330,
         n70331, n70332, n70333, n70334, n70335, n70336, n70337, n70338,
         n70339, n70340, n70341, n70342, n70343, n70344, n70345, n70346,
         n70347, n70348, n70349, n70350, n70351, n70352, n70353, n70354,
         n70355, n70356, n70357, n70358, n70359, n70360, n70361, n70362,
         n70363, n70364, n70365, n70366, n70367, n70368, n70369, n70370,
         n70371, n70372, n70373, n70374, n70375, n70376, n70377, n70378,
         n70379, n70380, n70381, n70382, n70383, n70384, n70385, n70386,
         n70387, n70388, n70389, n70390, n70391, n70392, n70393, n70394,
         n70395, n70396, n70397, n70398, n70399, n70400, n70401, n70402,
         n70403, n70404, n70405, n70406, n70407, n70408, n70409, n70410,
         n70411, n70412, n70413, n70414, n70415, n70416, n70417, n70418,
         n70419, n70420, n70421, n70422, n70423, n70424, n70425, n70426,
         n70427, n70428, n70429, n70430, n70431, n70432, n70433, n70434,
         n70435, n70436, n70437, n70438, n70439, n70440, n70441, n70442,
         n70443, n70444, n70445, n70446, n70447, n70448, n70449, n70450,
         n70451, n70452, n70453, n70454, n70455, n70456, n70457, n70458,
         n70459, n70460, n70461, n70462, n70463, n70464, n70465, n70466,
         n70467, n70468, n70469, n70470, n70471, n70472, n70473, n70474,
         n70475, n70476, n70477, n70478, n70479, n70480, n70481, n70482,
         n70483, n70484, n70485, n70486, n70487, n70488, n70489, n70490,
         n70491, n70492, n70493, n70494, n70495, n70496, n70497, n70498,
         n70499, n70500, n70501, n70502, n70503, n70504, n70505, n70506,
         n70507, n70508, n70509, n70510, n70511, n70512, n70513, n70514,
         n70515, n70516, n70517, n70518, n70519, n70520, n70521, n70522,
         n70523, n70524, n70525, n70526, n70527, n70528, n70529, n70530,
         n70531, n70532, n70533, n70534, n70535, n70536, n70537, n70538,
         n70539, n70540, n70541, n70542, n70543, n70544, n70545, n70546,
         n70547, n70548, n70549, n70550, n70551, n70552, n70553, n70554,
         n70555, n70556, n70557, n70558, n70559, n70560, n70561, n70562,
         n70563, n70564, n70565, n70566, n70567, n70568, n70569, n70570,
         n70571, n70572, n70573, n70574, n70575, n70576, n70577, n70578,
         n70579, n70580, n70581, n70582, n70583, n70584, n70585, n70586,
         n70587, n70588, n70589, n70590, n70591, n70592, n70593, n70594,
         n70595, n70596, n70597, n70598, n70599, n70600, n70601, n70602,
         n70603, n70604, n70605, n70606, n70607, n70608, n70609, n70610,
         n70611, n70612, n70613, n70614, n70615, n70616, n70617, n70618,
         n70619, n70620, n70621, n70622, n70623, n70624, n70625, n70626,
         n70627, n70628, n70629, n70630, n70631, n70632, n70633, n70634,
         n70635, n70636, n70637, n70638, n70639, n70640, n70641, n70642,
         n70643, n70644, n70645, n70646, n70647, n70648, n70649, n70650,
         n70651, n70652, n70653, n70654, n70655, n70656, n70657, n70658,
         n70659, n70660, n70661, n70662, n70663, n70664, n70665, n70666,
         n70667, n70668, n70669, n70670, n70671, n70672, n70673, n70674,
         n70675, n70676, n70677, n70678, n70679, n70680, n70681, n70682,
         n70683, n70684, n70685, n70686, n70687, n70688, n70689, n70690,
         n70691, n70692, n70693, n70694, n70695, n70696, n70697, n70698,
         n70699, n70700, n70701, n70702, n70703, n70704, n70705, n70706,
         n70707, n70708, n70709, n70710, n70711, n70712, n70713, n70714,
         n70715, n70716, n70717, n70718, n70719, n70720, n70721, n70722,
         n70723, n70724, n70725, n70726, n70727, n70728, n70729, n70730,
         n70731, n70732, n70733, n70734, n70735, n70736, n70737, n70738,
         n70739, n70740, n70741, n70742, n70743, n70744, n70745, n70746,
         n70747, n70748, n70749, n70750, n70751, n70752, n70753, n70754,
         n70755, n70756, n70757, n70758, n70759, n70760, n70761, n70762,
         n70763, n70764, n70765, n70766, n70767, n70768, n70769, n70770,
         n70771, n70772, n70773, n70774, n70775, n70776, n70777, n70778,
         n70779, n70780, n70781, n70782, n70783, n70784, n70785, n70786,
         n70787, n70788, n70789, n70790, n70791, n70792, n70793, n70794,
         n70795, n70796, n70797, n70798, n70799, n70800, n70801, n70802,
         n70803, n70804, n70805, n70806, n70807, n70808, n70809, n70810,
         n70811, n70812, n70813, n70814, n70815, n70816, n70817, n70818,
         n70819, n70820, n70821, n70822, n70823, n70824, n70825, n70826,
         n70827, n70828, n70829, n70830, n70831, n70832, n70833, n70834,
         n70835, n70836, n70837, n70838, n70839, n70840, n70841, n70842,
         n70843, n70844, n70845, n70846, n70847, n70848, n70849, n70850,
         n70851, n70852, n70853, n70854, n70855, n70856, n70857, n70858,
         n70859, n70860, n70861, n70862, n70863, n70864, n70865, n70866,
         n70867, n70868, n70869, n70870, n70871, n70872, n70873, n70874,
         n70875, n70876, n70877, n70878, n70879, n70880, n70881, n70882,
         n70883, n70884, n70885, n70886, n70887, n70888, n70889, n70890,
         n70891, n70892, n70893, n70894, n70895, n70896, n70897, n70898,
         n70899, n70900, n70901, n70902, n70903, n70904, n70905, n70906,
         n70907, n70908, n70909, n70910, n70911, n70912, n70913, n70914,
         n70915, n70916, n70917, n70918, n70919, n70920, n70921, n70922,
         n70923, n70924, n70925, n70926, n70927, n70928, n70929, n70930,
         n70931, n70932, n70933, n70934, n70935, n70936, n70937, n70938,
         n70939, n70940, n70941, n70942, n70943, n70944, n70945, n70946,
         n70947, n70948, n70949, n70950, n70951, n70952, n70953, n70954,
         n70955, n70956, n70957, n70958, n70959, n70960, n70961, n70962,
         n70963, n70964, n70965, n70966, n70967, n70968, n70969, n70970,
         n70971, n70972, n70973, n70974, n70975, n70976, n70977, n70978,
         n70979, n70980, n70981, n70982, n70983, n70984, n70985, n70986,
         n70987, n70988, n70989, n70990, n70991, n70992, n70993, n70994,
         n70995, n70996, n70997, n70998, n70999, n71000, n71001, n71002,
         n71003, n71004, n71005, n71006, n71007, n71008, n71009, n71010,
         n71011, n71012, n71013, n71014, n71015, n71016, n71017, n71018,
         n71019, n71020, n71021, n71022, n71023, n71024, n71025, n71026,
         n71027, n71028, n71029, n71030, n71031, n71032, n71033, n71034,
         n71035, n71036, n71037, n71038, n71039, n71040, n71041, n71042,
         n71043, n71044, n71045, n71046, n71047, n71048, n71049, n71050,
         n71051, n71052, n71053, n71054, n71055, n71056, n71057, n71058,
         n71059, n71060, n71061, n71062, n71063, n71064, n71065, n71066,
         n71067, n71068, n71069, n71070, n71071, n71072, n71073, n71074,
         n71075, n71076, n71077, n71078, n71079, n71080, n71081, n71082,
         n71083, n71084, n71085, n71086, n71087, n71088, n71089, n71090,
         n71091, n71092, n71093, n71094, n71095, n71096, n71097, n71098,
         n71099, n71100, n71101, n71102, n71103, n71104, n71105, n71106,
         n71107, n71108, n71109, n71110, n71111, n71112, n71113, n71114,
         n71115, n71116, n71117, n71118, n71119, n71120, n71121, n71122,
         n71123, n71124, n71125, n71126, n71127, n71128, n71129, n71130,
         n71131, n71132, n71133, n71134, n71135, n71136, n71137, n71138,
         n71139, n71140, n71141, n71142, n71143, n71144, n71145, n71146,
         n71147, n71148, n71149, n71150, n71151, n71152, n71153, n71154,
         n71155, n71156, n71157, n71158, n71159, n71160, n71161, n71162,
         n71163, n71164, n71165, n71166, n71167, n71168, n71169, n71170,
         n71171, n71172, n71173, n71174, n71175, n71176, n71177, n71178,
         n71179, n71180, n71181, n71182, n71183, n71184, n71185, n71186,
         n71187, n71188, n71189, n71190, n71191, n71192, n71193, n71194,
         n71195, n71196, n71197, n71198, n71199, n71200, n71201, n71202,
         n71203, n71204, n71205, n71206, n71207, n71208, n71209, n71210,
         n71211, n71212, n71213, n71214, n71215, n71216, n71217, n71218,
         n71219, n71220, n71221, n71222, n71223, n71224, n71225, n71226,
         n71227, n71228, n71229, n71230, n71231, n71232, n71233, n71234,
         n71235, n71236, n71237, n71238, n71239, n71240, n71241, n71242,
         n71243, n71244, n71245, n71246, n71247, n71248, n71249, n71250,
         n71251, n71252, n71253, n71254, n71255, n71256, n71257, n71258,
         n71259, n71260, n71261, n71262, n71263, n71264, n71265, n71266,
         n71267, n71268, n71269, n71270, n71271, n71272, n71273, n71274,
         n71275, n71276, n71277, n71278, n71279, n71280, n71281, n71282,
         n71283, n71284, n71285, n71286, n71287, n71288, n71289, n71290,
         n71291, n71292, n71293, n71294, n71295, n71296, n71297, n71298,
         n71299, n71300, n71301, n71302, n71303, n71304, n71305, n71306,
         n71307, n71308, n71309, n71310, n71311, n71312, n71313, n71314,
         n71315, n71316, n71317, n71318, n71319, n71320, n71321, n71322,
         n71323, n71324, n71325, n71326, n71327, n71328, n71329, n71330,
         n71331, n71332, n71333, n71334, n71335, n71336, n71337, n71338,
         n71339, n71340, n71341, n71342, n71343, n71344, n71345, n71346,
         n71347, n71348, n71349, n71350, n71351, n71352, n71353, n71354,
         n71355, n71356, n71357, n71358, n71359, n71360, n71361, n71362,
         n71363, n71364, n71365, n71366, n71367, n71368, n71369, n71370,
         n71371, n71372, n71373, n71374, n71375, n71376, n71377, n71378,
         n71379, n71380, n71381, n71382, n71383, n71384, n71385, n71386,
         n71387, n71388, n71389, n71390, n71391, n71392, n71393, n71394,
         n71395, n71396, n71397, n71398, n71399, n71400, n71401, n71402,
         n71403, n71404, n71405, n71406, n71407, n71408, n71409, n71410,
         n71411, n71412, n71413, n71414, n71415, n71416, n71417, n71418,
         n71419, n71420, n71421, n71422, n71423, n71424, n71425, n71426,
         n71427, n71428, n71429, n71430, n71431, n71432, n71433, n71434,
         n71435, n71436, n71437, n71438, n71439, n71440, n71441, n71442,
         n71443, n71444, n71445, n71446, n71447, n71448, n71449, n71450,
         n71451, n71452, n71453, n71454, n71455, n71456, n71457, n71458,
         n71459, n71460, n71461, n71462, n71463, n71464, n71465, n71466,
         n71467, n71468, n71469, n71470, n71471, n71472, n71473, n71474,
         n71475, n71476, n71477, n71478, n71479, n71480, n71481, n71482,
         n71483, n71484, n71485, n71486, n71487, n71488, n71489, n71490,
         n71491, n71492, n71493, n71494, n71495, n71496, n71497, n71498,
         n71499, n71500, n71501, n71502, n71503, n71504, n71505, n71506,
         n71507, n71508, n71509, n71510, n71511, n71512, n71513, n71514,
         n71515, n71516, n71517, n71518, n71519, n71520, n71521, n71522,
         n71523, n71524, n71525, n71526, n71527, n71528, n71529, n71530,
         n71531, n71532, n71533, n71534, n71535, n71536, n71537, n71538,
         n71539, n71540, n71541, n71542, n71543, n71544, n71545, n71546,
         n71547, n71548, n71549, n71550, n71551, n71552, n71553, n71554,
         n71555, n71556, n71557, n71558, n71559, n71560, n71561, n71562,
         n71563, n71564, n71565, n71566, n71567, n71568, n71569, n71570,
         n71571, n71572, n71573, n71574, n71575, n71576, n71577, n71578,
         n71579, n71580, n71581, n71582, n71583, n71584, n71585, n71586,
         n71587, n71588, n71589, n71590, n71591, n71592, n71593, n71594,
         n71595, n71596, n71597, n71598, n71599, n71600, n71601, n71602,
         n71603, n71604, n71605, n71606, n71607, n71608, n71609, n71610,
         n71611, n71612, n71613, n71614, n71615, n71616, n71617, n71618,
         n71619, n71620, n71621, n71622, n71623, n71624, n71625, n71626,
         n71627, n71628, n71629, n71630, n71631, n71632, n71633, n71634,
         n71635, n71636, n71637, n71638, n71639, n71640, n71641, n71642,
         n71643, n71644, n71645, n71646, n71647, n71648, n71649, n71650,
         n71651, n71652, n71653, n71654, n71655, n71656, n71657, n71658,
         n71659, n71660, n71661, n71662, n71663, n71664, n71665, n71666,
         n71667, n71668, n71669, n71670, n71671, n71672, n71673, n71674,
         n71675, n71676, n71677, n71678, n71679, n71680, n71681, n71682,
         n71683, n71684, n71685, n71686, n71687, n71688, n71689, n71690,
         n71691, n71692, n71693, n71694, n71695, n71696, n71697, n71698,
         n71699, n71700, n71701, n71702, n71703, n71704, n71705, n71706,
         n71707, n71708, n71709, n71710, n71711, n71712, n71713, n71714,
         n71715, n71716, n71717, n71718, n71719, n71720, n71721, n71722,
         n71723, n71724, n71725, n71726, n71727, n71728, n71729, n71730,
         n71731, n71732, n71733, n71734, n71735, n71736, n71737, n71738,
         n71739, n71740, n71741, n71742, n71743, n71744, n71745, n71746,
         n71747, n71748, n71749, n71750, n71751, n71752, n71753, n71754,
         n71755, n71756, n71757, n71758, n71759, n71760, n71761, n71762,
         n71763, n71764, n71765, n71766, n71767, n71768, n71769, n71770,
         n71771, n71772, n71773, n71774, n71775, n71776, n71777, n71778,
         n71779, n71780, n71781, n71782, n71783, n71784, n71785, n71786,
         n71787, n71788, n71789, n71790, n71791, n71792, n71793, n71794,
         n71795, n71796, n71797, n71798, n71799, n71800, n71801, n71802,
         n71803, n71804, n71805, n71806, n71807, n71808, n71809, n71810,
         n71811, n71812, n71813, n71814, n71815, n71816, n71817, n71818,
         n71819, n71820, n71821, n71822, n71823, n71824, n71825, n71826,
         n71827, n71828, n71829, n71830, n71831, n71832, n71833, n71834,
         n71835, n71836, n71837, n71838, n71839, n71840, n71841, n71842,
         n71843, n71844, n71845, n71846, n71847, n71848, n71849, n71850,
         n71851, n71852, n71853, n71854, n71855, n71856, n71857, n71858,
         n71859, n71860, n71861, n71862, n71863, n71864, n71865, n71866,
         n71867, n71868, n71869, n71870, n71871, n71872, n71873, n71874,
         n71875, n71876, n71877, n71878, n71879, n71880, n71881, n71882,
         n71883, n71884, n71885, n71886, n71887, n71888, n71889, n71890,
         n71891, n71892, n71893, n71894, n71895, n71896, n71897, n71898,
         n71899, n71900, n71901, n71902, n71903, n71904, n71905, n71906,
         n71907, n71908, n71909, n71910, n71911, n71912, n71913, n71914,
         n71915, n71916, n71917, n71918, n71919, n71920, n71921, n71922,
         n71923, n71924, n71925, n71926, n71927, n71928, n71929, n71930,
         n71931, n71932, n71933, n71934, n71935, n71936, n71937, n71938,
         n71939, n71940, n71941, n71942, n71943, n71944, n71945, n71946,
         n71947, n71948, n71949, n71950, n71951, n71952, n71953, n71954,
         n71955, n71956, n71957, n71958, n71959, n71960, n71961, n71962,
         n71963, n71964, n71965, n71966, n71967, n71968, n71969, n71970,
         n71971, n71972, n71973, n71974, n71975, n71976, n71977, n71978,
         n71979, n71980, n71981, n71982, n71983, n71984, n71985, n71986,
         n71987, n71988, n71989, n71990, n71991, n71992, n71993, n71994,
         n71995, n71996, n71997, n71998, n71999, n72000, n72001, n72002,
         n72003, n72004, n72005, n72006, n72007, n72008, n72009, n72010,
         n72011, n72012, n72013, n72014, n72015, n72016, n72017, n72018,
         n72019, n72020, n72021, n72022, n72023, n72024, n72025, n72026,
         n72027, n72028, n72029, n72030, n72031, n72032, n72033, n72034,
         n72035, n72036, n72037, n72038, n72039, n72040, n72041, n72042,
         n72043, n72044, n72045, n72046, n72047, n72048, n72049, n72050,
         n72051, n72052, n72053, n72054, n72055, n72056, n72057, n72058,
         n72059, n72060, n72061, n72062, n72063, n72064, n72065, n72066,
         n72067, n72068, n72069, n72070, n72071, n72072, n72073, n72074,
         n72075, n72076, n72077, n72078, n72079, n72080, n72081, n72082,
         n72083, n72084, n72085, n72086, n72087, n72088, n72089, n72090,
         n72091, n72092, n72093, n72094, n72095, n72096, n72097, n72098,
         n72099, n72100, n72101, n72102, n72103, n72104, n72105, n72106,
         n72107, n72108, n72109, n72110, n72111, n72112, n72113, n72114,
         n72115, n72116, n72117, n72118, n72119, n72120, n72121, n72122,
         n72123, n72124, n72125, n72126, n72127, n72128, n72129, n72130,
         n72131, n72132, n72133, n72134, n72135, n72136, n72137, n72138,
         n72139, n72140, n72141, n72142, n72143, n72144, n72145, n72146,
         n72147, n72148, n72149, n72150, n72151, n72152, n72153, n72154,
         n72155, n72156, n72157, n72158, n72159, n72160, n72161, n72162,
         n72163, n72164, n72165, n72166, n72167, n72168, n72169, n72170,
         n72171, n72172, n72173, n72174, n72175, n72176, n72177, n72178,
         n72179, n72180, n72181, n72182, n72183, n72184, n72185, n72186,
         n72187, n72188, n72189, n72190, n72191, n72192, n72193, n72194,
         n72195, n72196, n72197, n72198, n72199, n72200, n72201, n72202,
         n72203, n72204, n72205, n72206, n72207, n72208, n72209, n72210,
         n72211, n72212, n72213, n72214, n72215, n72216, n72217, n72218,
         n72219, n72220, n72221, n72222, n72223, n72224, n72225, n72226,
         n72227, n72228, n72229, n72230, n72231, n72232, n72233, n72234,
         n72235, n72236, n72237, n72238, n72239, n72240, n72241, n72242,
         n72243, n72244, n72245, n72246, n72247, n72248, n72249, n72250,
         n72251, n72252, n72253, n72254, n72255, n72256, n72257, n72258,
         n72259, n72260, n72261, n72262, n72263, n72264, n72265, n72266,
         n72267, n72268, n72269, n72270, n72271, n72272, n72273, n72274,
         n72275, n72276, n72277, n72278, n72279, n72280, n72281, n72282,
         n72283, n72284, n72285, n72286, n72287, n72288, n72289, n72290,
         n72291, n72292, n72293, n72294, n72295, n72296, n72297, n72298,
         n72299, n72300, n72301, n72302, n72303, n72304, n72305, n72306,
         n72307, n72308, n72309, n72310, n72311, n72312, n72313, n72314,
         n72315, n72316, n72317, n72318, n72319, n72320, n72321, n72322,
         n72323, n72324, n72325, n72326, n72327, n72328, n72329, n72330,
         n72331, n72332, n72333, n72334, n72335, n72336, n72337, n72338,
         n72339, n72340, n72341, n72342, n72343, n72344, n72345, n72346,
         n72347, n72348, n72349, n72350, n72351, n72352, n72353, n72354,
         n72355, n72356, n72357, n72358, n72359, n72360, n72361, n72362,
         n72363, n72364, n72365, n72366, n72367, n72368, n72369, n72370,
         n72371, n72372, n72373, n72374, n72375, n72376, n72377, n72378,
         n72379, n72380, n72381, n72382, n72383, n72384, n72385, n72386,
         n72387, n72388, n72389, n72390, n72391, n72392, n72393, n72394,
         n72395, n72396, n72397, n72398, n72399, n72400, n72401, n72402,
         n72403, n72404, n72405, n72406, n72407, n72408, n72409, n72410,
         n72411, n72412, n72413, n72414, n72415, n72416, n72417, n72418,
         n72419, n72420, n72421, n72422, n72423, n72424, n72425, n72426,
         n72427, n72428, n72429, n72430, n72431, n72432, n72433, n72434,
         n72435, n72436, n72437, n72438, n72439, n72440, n72441, n72442,
         n72443, n72444, n72445, n72446, n72447, n72448, n72449, n72450,
         n72451, n72452, n72453, n72454, n72455, n72456, n72457, n72458,
         n72459, n72460, n72461, n72462, n72463, n72464, n72465, n72466,
         n72467, n72468, n72469, n72470, n72471, n72472, n72473, n72474,
         n72475, n72476, n72477, n72478, n72479, n72480, n72481, n72482,
         n72483, n72484, n72485, n72486, n72487, n72488, n72489, n72490,
         n72491, n72492, n72493, n72494, n72495, n72496, n72497, n72498,
         n72499, n72500, n72501, n72502, n72503, n72504, n72505, n72506,
         n72507, n72508, n72509, n72510, n72511, n72512, n72513, n72514,
         n72515, n72516, n72517, n72518, n72519, n72520, n72521, n72522,
         n72523, n72524, n72525, n72526, n72527, n72528, n72529, n72530,
         n72531, n72532, n72533, n72534, n72535, n72536, n72537, n72538,
         n72539, n72540, n72541, n72542, n72543, n72544, n72545, n72546,
         n72547, n72548, n72549, n72550, n72551, n72552, n72553, n72554,
         n72555, n72556, n72557, n72558, n72559, n72560, n72561, n72562,
         n72563, n72564, n72565, n72566, n72567, n72568, n72569, n72570,
         n72571, n72572, n72573, n72574, n72575, n72576, n72577, n72578,
         n72579, n72580, n72581, n72582, n72583, n72584, n72585, n72586,
         n72587, n72588, n72589, n72590, n72591, n72592, n72593, n72594,
         n72595, n72596, n72597, n72598, n72599, n72600, n72601, n72602,
         n72603, n72604, n72605, n72606, n72607, n72608, n72609, n72610,
         n72611, n72612, n72613, n72614, n72615, n72616, n72617, n72618,
         n72619, n72620, n72621, n72622, n72623, n72624, n72625, n72626,
         n72627, n72628, n72629, n72630, n72631, n72632, n72633, n72634,
         n72635, n72636, n72637, n72638, n72639, n72640, n72641, n72642,
         n72643, n72644, n72645, n72646, n72647, n72648, n72649, n72650,
         n72651, n72652, n72653, n72654, n72655, n72656, n72657, n72658,
         n72659, n72660, n72661, n72662, n72663, n72664, n72665, n72666,
         n72667, n72668, n72669, n72670, n72671, n72672, n72673, n72674,
         n72675, n72676, n72677, n72678, n72679, n72680, n72681, n72682,
         n72683, n72684, n72685, n72686, n72687, n72688, n72689, n72690,
         n72691, n72692, n72693, n72694, n72695, n72696, n72697, n72698,
         n72699, n72700, n72701, n72702, n72703, n72704, n72705, n72706,
         n72707, n72708, n72709, n72710, n72711, n72712, n72713, n72714,
         n72715, n72716, n72717, n72718, n72719, n72720, n72721, n72722,
         n72723, n72724, n72725, n72726, n72727, n72728, n72729, n72730,
         n72731, n72732, n72733, n72734, n72735, n72736, n72737, n72738,
         n72739, n72740, n72741, n72742, n72743, n72744, n72745, n72746,
         n72747, n72748, n72749, n72750, n72751, n72752, n72753, n72754,
         n72755, n72756, n72757, n72758, n72759, n72760, n72761, n72762,
         n72763, n72764, n72765, n72766, n72767, n72768, n72769, n72770,
         n72771, n72772, n72773, n72774, n72775, n72776, n72777, n72778,
         n72779, n72780, n72781, n72782, n72783, n72784, n72785, n72786,
         n72787, n72788, n72789, n72790, n72791, n72792, n72793, n72794,
         n72795, n72796, n72797, n72798, n72799, n72800, n72801, n72802,
         n72803, n72804, n72805, n72806, n72807, n72808, n72809, n72810,
         n72811, n72812, n72813, n72814, n72815, n72816, n72817, n72818,
         n72819, n72820, n72821, n72822, n72823, n72824, n72825, n72826,
         n72827, n72828, n72829, n72830, n72831, n72832, n72833, n72834,
         n72835, n72836, n72837, n72838, n72839, n72840, n72841, n72842,
         n72843, n72844, n72845, n72846, n72847, n72848, n72849, n72850,
         n72851, n72852, n72853, n72854, n72855, n72856, n72857, n72858,
         n72859, n72860, n72861, n72862, n72863, n72864, n72865, n72866,
         n72867, n72868, n72869, n72870, n72871, n72872, n72873, n72874,
         n72875, n72876, n72877, n72878, n72879, n72880, n72881, n72882,
         n72883, n72884, n72885, n72886, n72887, n72888, n72889, n72890,
         n72891, n72892, n72893, n72894, n72895, n72896, n72897, n72898,
         n72899, n72900, n72901, n72902, n72903, n72904, n72905, n72906,
         n72907, n72908, n72909, n72910, n72911, n72912, n72913, n72914,
         n72915, n72916, n72917, n72918, n72919, n72920, n72921, n72922,
         n72923, n72924, n72925, n72926, n72927, n72928, n72929, n72930,
         n72931, n72932, n72933, n72934, n72935, n72936, n72937, n72938,
         n72939, n72940, n72941, n72942, n72943, n72944, n72945, n72946,
         n72947, n72948, n72949, n72950, n72951, n72952, n72953, n72954,
         n72955, n72956, n72957, n72958, n72959, n72960, n72961, n72962,
         n72963, n72964, n72965, n72966, n72967, n72968, n72969, n72970,
         n72971, n72972, n72973, n72974, n72975, n72976, n72977, n72978,
         n72979, n72980, n72981, n72982, n72983, n72984, n72985, n72986,
         n72987, n72988, n72989, n72990, n72991, n72992, n72993, n72994,
         n72995, n72996, n72997, n72998, n72999, n73000, n73001, n73002,
         n73003, n73004, n73005, n73006, n73007, n73008, n73009, n73010,
         n73011, n73012, n73013, n73014, n73015, n73016, n73017, n73018,
         n73019, n73020, n73021, n73022, n73023, n73024, n73025, n73026,
         n73027, n73028, n73029, n73030, n73031, n73032, n73033, n73034,
         n73035, n73036, n73037, n73038, n73039, n73040, n73041, n73042,
         n73043, n73044, n73045, n73046, n73047, n73048, n73049, n73050,
         n73051, n73052, n73053, n73054, n73055, n73056, n73057, n73058,
         n73059, n73060, n73061, n73062, n73063, n73064, n73065, n73066,
         n73067, n73068, n73069, n73070, n73071, n73072, n73073, n73074,
         n73075, n73076, n73077, n73078, n73079, n73080, n73081, n73082,
         n73083, n73084, n73085, n73086, n73087, n73088, n73089, n73090,
         n73091, n73092, n73093, n73094, n73095, n73096, n73097, n73098,
         n73099, n73100, n73101, n73102, n73103, n73104, n73105, n73106,
         n73107, n73108, n73109, n73110, n73111, n73112, n73113, n73114,
         n73115, n73116, n73117, n73118, n73119, n73120, n73121, n73122,
         n73123, n73124, n73125, n73126, n73127, n73128, n73129, n73130,
         n73131, n73132, n73133, n73134, n73135, n73136, n73137, n73138,
         n73139, n73140, n73141, n73142, n73143, n73144, n73145, n73146,
         n73147, n73148, n73149, n73150, n73151, n73152, n73153, n73154,
         n73155, n73156, n73157, n73158, n73159, n73160, n73161, n73162,
         n73163, n73164, n73165, n73166, n73167, n73168, n73169, n73170,
         n73171, n73172, n73173, n73174, n73175, n73176, n73177, n73178,
         n73179, n73180, n73181, n73182, n73183, n73184, n73185, n73186,
         n73187, n73188, n73189, n73190, n73191, n73192, n73193, n73194,
         n73195, n73196, n73197, n73198, n73199, n73200, n73201, n73202,
         n73203, n73204, n73205, n73206, n73207, n73208, n73209, n73210,
         n73211, n73212, n73213, n73214, n73215, n73216, n73217, n73218,
         n73219, n73220, n73221, n73222, n73223, n73224, n73225, n73226,
         n73227, n73228, n73229, n73230, n73231, n73232, n73233, n73234,
         n73235, n73236, n73237, n73238, n73239, n73240, n73241, n73242,
         n73243, n73244, n73245, n73246, n73247, n73248, n73249, n73250,
         n73251, n73252, n73253, n73254, n73255, n73256, n73257, n73258,
         n73259, n73260, n73261, n73262, n73263, n73264, n73265, n73266,
         n73267, n73268, n73269, n73270, n73271, n73272, n73273, n73274,
         n73275, n73276, n73277, n73278, n73279, n73280, n73281, n73282,
         n73283, n73284, n73285, n73286, n73287, n73288, n73289, n73290,
         n73291, n73292, n73293, n73294, n73295, n73296, n73297, n73298,
         n73299, n73300, n73301, n73302, n73303, n73304, n73305, n73306,
         n73307, n73308, n73309, n73310, n73311, n73312, n73313, n73314,
         n73315, n73316, n73317, n73318, n73319, n73320, n73321, n73322,
         n73323, n73324, n73325, n73326, n73327, n73328, n73329, n73330,
         n73331, n73332, n73333, n73334, n73335, n73336, n73337, n73338,
         n73339, n73340, n73341, n73342, n73343, n73344, n73345, n73346,
         n73347, n73348, n73349, n73350, n73351, n73352, n73353, n73354,
         n73355, n73356, n73357, n73358, n73359, n73360, n73361, n73362,
         n73363, n73364, n73365, n73366, n73367, n73368, n73369, n73370,
         n73371, n73372, n73373, n73374, n73375, n73376, n73377, n73378,
         n73379, n73380, n73381, n73382, n73383, n73384, n73385, n73386,
         n73387, n73388, n73389, n73390, n73391, n73392, n73393, n73394,
         n73395, n73396, n73397, n73398, n73399, n73400, n73401, n73402,
         n73403, n73404, n73405, n73406, n73407, n73408, n73409, n73410,
         n73411, n73412, n73413, n73414, n73415, n73416, n73417, n73418,
         n73419, n73420, n73421, n73422, n73423, n73424, n73425, n73426,
         n73427, n73428, n73429, n73430, n73431, n73432, n73433, n73434,
         n73435, n73436, n73437, n73438, n73439, n73440, n73441, n73442,
         n73443, n73444, n73445, n73446, n73447, n73448, n73449, n73450,
         n73451, n73452, n73453, n73454, n73455, n73456, n73457, n73458,
         n73459, n73460, n73461, n73462, n73463, n73464, n73465, n73466,
         n73467, n73468, n73469, n73470, n73471, n73472, n73473, n73474,
         n73475, n73476, n73477, n73478, n73479, n73480, n73481, n73482,
         n73483, n73484, n73485, n73486, n73487, n73488, n73489, n73490,
         n73491, n73492, n73493, n73494, n73495, n73496, n73497, n73498,
         n73499, n73500, n73501, n73502, n73503, n73504, n73505, n73506,
         n73507, n73508, n73509, n73510, n73511, n73512, n73513, n73514,
         n73515, n73516, n73517, n73518, n73519, n73520, n73521, n73522,
         n73523, n73524, n73525, n73526, n73527, n73528, n73529, n73530,
         n73531, n73532, n73533, n73534, n73535, n73536, n73537, n73538,
         n73539, n73540, n73541, n73542, n73543, n73544, n73545, n73546,
         n73547, n73548, n73549, n73550, n73551, n73552, n73553, n73554,
         n73555, n73556, n73557, n73558, n73559, n73560, n73561, n73562,
         n73563, n73564, n73565, n73566, n73567, n73568, n73569, n73570,
         n73571, n73572, n73573, n73574, n73575, n73576, n73577, n73578,
         n73579, n73580, n73581, n73582, n73583, n73584, n73585, n73586,
         n73587, n73588, n73589, n73590, n73591, n73592, n73593, n73594,
         n73595, n73596, n73597, n73598, n73599, n73600, n73601, n73602,
         n73603, n73604, n73605, n73606, n73607, n73608, n73609, n73610,
         n73611, n73612, n73613, n73614, n73615, n73616, n73617, n73618,
         n73619, n73620, n73621, n73622, n73623, n73624, n73625, n73626,
         n73627, n73628, n73629, n73630, n73631, n73632, n73633, n73634,
         n73635, n73636, n73637, n73638, n73639, n73640, n73641, n73642,
         n73643, n73644, n73645, n73646, n73647, n73648, n73649, n73650,
         n73651, n73652, n73653, n73654, n73655, n73656, n73657, n73658,
         n73659, n73660, n73661, n73662, n73663, n73664, n73665, n73666,
         n73667, n73668, n73669, n73670, n73671, n73672, n73673, n73674,
         n73675, n73676, n73677, n73678, n73679, n73680, n73681, n73682,
         n73683, n73684, n73685, n73686, n73687, n73688, n73689, n73690,
         n73691, n73692, n73693, n73694, n73695, n73696, n73697, n73698,
         n73699, n73700, n73701, n73702, n73703, n73704, n73705, n73706,
         n73707, n73708, n73709, n73710, n73711, n73712, n73713, n73714,
         n73715, n73716, n73717, n73718, n73719, n73720, n73721, n73722,
         n73723, n73724, n73725, n73726, n73727, n73728, n73729, n73730,
         n73731, n73732, n73733, n73734, n73735, n73736, n73737, n73738,
         n73739, n73740, n73741, n73742, n73743, n73744, n73745, n73746,
         n73747, n73748, n73749, n73750, n73751, n73752, n73753, n73754,
         n73755, n73756, n73757, n73758, n73759, n73760, n73761, n73762,
         n73763, n73764, n73765, n73766, n73767, n73768, n73769, n73770,
         n73771, n73772, n73773, n73774, n73775, n73776, n73777, n73778,
         n73779, n73780, n73781, n73782, n73783, n73784, n73785, n73786,
         n73787, n73788, n73789, n73790, n73791, n73792, n73793, n73794,
         n73795, n73796, n73797, n73798, n73799, n73800, n73801, n73802,
         n73803, n73804, n73805, n73806, n73807, n73808, n73809, n73810,
         n73811, n73812, n73813, n73814, n73815, n73816, n73817, n73818,
         n73819, n73820, n73821, n73822, n73823, n73824, n73825, n73826,
         n73827, n73828, n73829, n73830, n73831, n73832, n73833, n73834,
         n73835, n73836, n73837, n73838, n73839, n73840, n73841, n73842,
         n73843, n73844, n73845, n73846, n73847, n73848, n73849, n73850,
         n73851, n73852, n73853, n73854, n73855, n73856, n73857, n73858,
         n73859, n73860, n73861, n73862, n73863, n73864, n73865, n73866,
         n73867, n73868, n73869, n73870, n73871, n73872, n73873, n73874,
         n73875, n73876, n73877, n73878, n73879, n73880, n73881, n73882,
         n73883, n73884, n73885, n73886, n73887, n73888, n73889, n73890,
         n73891, n73892, n73893, n73894, n73895, n73896, n73897, n73898,
         n73899, n73900, n73901, n73902, n73903, n73904, n73905, n73906,
         n73907, n73908, n73909, n73910, n73911, n73912, n73913, n73914,
         n73915, n73916, n73917, n73918, n73919, n73920, n73921, n73922,
         n73923, n73924, n73925, n73926, n73927, n73928, n73929, n73930,
         n73931, n73932, n73933, n73934, n73935, n73936, n73937, n73938,
         n73939, n73940, n73941, n73942, n73943, n73944, n73945, n73946,
         n73947, n73948, n73949, n73950, n73951, n73952, n73953, n73954,
         n73955, n73956, n73957, n73958, n73959, n73960, n73961, n73962,
         n73963, n73964, n73965, n73966, n73967, n73968, n73969, n73970,
         n73971, n73972, n73973, n73974, n73975, n73976, n73977, n73978,
         n73979, n73980, n73981, n73982, n73983, n73984, n73985, n73986,
         n73987, n73988, n73989, n73990, n73991, n73992, n73993, n73994,
         n73995, n73996, n73997, n73998, n73999, n74000, n74001, n74002,
         n74003, n74004, n74005, n74006, n74007, n74008, n74009, n74010,
         n74011, n74012, n74013, n74014, n74015, n74016, n74017, n74018,
         n74019, n74020, n74021, n74022, n74023, n74024, n74025, n74026,
         n74027, n74028, n74029, n74030, n74031, n74032, n74033, n74034,
         n74035, n74036, n74037, n74038, n74039, n74040, n74041, n74042,
         n74043, n74044, n74045, n74046, n74047, n74048, n74049, n74050,
         n74051, n74052, n74053, n74054, n74055, n74056, n74057, n74058,
         n74059, n74060, n74061, n74062, n74063, n74064, n74065, n74066,
         n74067, n74068, n74069, n74070, n74071, n74072, n74073, n74074,
         n74075, n74076, n74077, n74078, n74079, n74080, n74081, n74082,
         n74083, n74084, n74085, n74086, n74087, n74088, n74089, n74090,
         n74091, n74092, n74093, n74094, n74095, n74096, n74097, n74098,
         n74099, n74100, n74101, n74102, n74103, n74104, n74105, n74106,
         n74107, n74108, n74109, n74110, n74111, n74112, n74113, n74114,
         n74115, n74116, n74117, n74118, n74119, n74120, n74121, n74122,
         n74123, n74124, n74125, n74126, n74127, n74128, n74129, n74130,
         n74131, n74132, n74133, n74134, n74135, n74136, n74137, n74138,
         n74139, n74140, n74141, n74142, n74143, n74144, n74145, n74146,
         n74147, n74148, n74149, n74150, n74151, n74152, n74153, n74154,
         n74155, n74156, n74157, n74158, n74159, n74160, n74161, n74162,
         n74163, n74164, n74165, n74166, n74167, n74168, n74169, n74170,
         n74171, n74172, n74173, n74174, n74175, n74176, n74177, n74178,
         n74179, n74180, n74181, n74182, n74183, n74184, n74185, n74186,
         n74187, n74188, n74189, n74190, n74191, n74192, n74193, n74194,
         n74195, n74196, n74197, n74198, n74199, n74200, n74201, n74202,
         n74203, n74204, n74205, n74206, n74207, n74208, n74209, n74210,
         n74211, n74212, n74213, n74214, n74215, n74216, n74217, n74218,
         n74219, n74220, n74221, n74222, n74223, n74224, n74225, n74226,
         n74227, n74228, n74229, n74230, n74231, n74232, n74233, n74234,
         n74235, n74236, n74237, n74238, n74239, n74240, n74241, n74242,
         n74243, n74244, n74245, n74246, n74247, n74248, n74249, n74250,
         n74251, n74252, n74253, n74254, n74255, n74256, n74257, n74258,
         n74259, n74260, n74261, n74262, n74263, n74264, n74265, n74266,
         n74267, n74268, n74269, n74270, n74271, n74272, n74273, n74274,
         n74275, n74276, n74277, n74278, n74279, n74280, n74281, n74282,
         n74283, n74284, n74285, n74286, n74287, n74288, n74289, n74290,
         n74291, n74292, n74293, n74294, n74295, n74296, n74297, n74298,
         n74299, n74300, n74301, n74302, n74303, n74304, n74305, n74306,
         n74307, n74308, n74309, n74310, n74311, n74312, n74313, n74314,
         n74315, n74316, n74317, n74318, n74319, n74320, n74321, n74322,
         n74323, n74324, n74325, n74326, n74327, n74328, n74329, n74330,
         n74331, n74332, n74333, n74334, n74335, n74336, n74337, n74338,
         n74339, n74340, n74341, n74342, n74343, n74344, n74345, n74346,
         n74347, n74348, n74349, n74350, n74351, n74352, n74353, n74354,
         n74355, n74356, n74357, n74358, n74359, n74360, n74361, n74362,
         n74363, n74364, n74365, n74366, n74367, n74368, n74369, n74370,
         n74371, n74372, n74373, n74374, n74375, n74376, n74377, n74378,
         n74379, n74380, n74381, n74382, n74383, n74384, n74385, n74386,
         n74387, n74388, n74389, n74390, n74391, n74392, n74393, n74394,
         n74395, n74396, n74397, n74398, n74399, n74400, n74401, n74402,
         n74403, n74404, n74405, n74406, n74407, n74408, n74409, n74410,
         n74411, n74412, n74413, n74414, n74415, n74416, n74417, n74418,
         n74419, n74420, n74421, n74422, n74423, n74424, n74425, n74426,
         n74427, n74428, n74429, n74430, n74431, n74432, n74433, n74434,
         n74435, n74436, n74437, n74438, n74439, n74440, n74441, n74442,
         n74443, n74444, n74445, n74446, n74447, n74448, n74449, n74450,
         n74451, n74452, n74453, n74454, n74455, n74456, n74457, n74458,
         n74459, n74460, n74461, n74462, n74463, n74464, n74465, n74466,
         n74467, n74468, n74469, n74470, n74471, n74472, n74473, n74474,
         n74475, n74476, n74477, n74478, n74479, n74480, n74481, n74482,
         n74483, n74484, n74485, n74486, n74487, n74488, n74489, n74490,
         n74491, n74492, n74493, n74494, n74495, n74496, n74497, n74498,
         n74499, n74500, n74501, n74502, n74503, n74504, n74505, n74506,
         n74507, n74508, n74509, n74510, n74511, n74512, n74513, n74514,
         n74515, n74516, n74517, n74518, n74519, n74520, n74521, n74522,
         n74523, n74524, n74525, n74526, n74527, n74528, n74529, n74530,
         n74531, n74532, n74533, n74534, n74535, n74536, n74537, n74538,
         n74539, n74540, n74541, n74542, n74543, n74544, n74545, n74546,
         n74547, n74548, n74549, n74550, n74551, n74552, n74553, n74554,
         n74555, n74556, n74557, n74558, n74559, n74560, n74561, n74562,
         n74563, n74564, n74565, n74566, n74567, n74568, n74569, n74570,
         n74571, n74572, n74573, n74574, n74575, n74576, n74577, n74578,
         n74579, n74580, n74581, n74582, n74583, n74584, n74585, n74586,
         n74587, n74588, n74589, n74590, n74591, n74592, n74593, n74594,
         n74595, n74596, n74597, n74598, n74599, n74600, n74601, n74602,
         n74603, n74604, n74605, n74606, n74607, n74608, n74609, n74610,
         n74611, n74612, n74613, n74614, n74615, n74616, n74617, n74618,
         n74619, n74620, n74621, n74622, n74623, n74624, n74625, n74626,
         n74627, n74628, n74629, n74630, n74631, n74632, n74633, n74634,
         n74635, n74636, n74637, n74638, n74639, n74640, n74641, n74642,
         n74643, n74644, n74645, n74646, n74647, n74648, n74649, n74650,
         n74651, n74652, n74653, n74654, n74655, n74656, n74657, n74658,
         n74659, n74660, n74661, n74662, n74663, n74664, n74665, n74666,
         n74667, n74668, n74669, n74670, n74671, n74672, n74673, n74674,
         n74675, n74676, n74677, n74678, n74679, n74680, n74681, n74682,
         n74683, n74684, n74685, n74686, n74687, n74688, n74689, n74690,
         n74691, n74692, n74693, n74694, n74695, n74696, n74697, n74698,
         n74699, n74700, n74701, n74702, n74703, n74704, n74705, n74706,
         n74707, n74708, n74709, n74710, n74711, n74712, n74713, n74714,
         n74715, n74716, n74717, n74718, n74719, n74720, n74721, n74722,
         n74723, n74724, n74725, n74726, n74727, n74728, n74729, n74730,
         n74731, n74732, n74733, n74734, n74735, n74736, n74737, n74738,
         n74739, n74740, n74741, n74742, n74743, n74744, n74745, n74746,
         n74747, n74748, n74749, n74750, n74751, n74752, n74753, n74754,
         n74755, n74756, n74757, n74758, n74759, n74760, n74761, n74762,
         n74763, n74764, n74765, n74766, n74767, n74768, n74769, n74770,
         n74771, n74772, n74773, n74774, n74775, n74776, n74777, n74778,
         n74779, n74780, n74781, n74782, n74783, n74784, n74785, n74786,
         n74787, n74788, n74789, n74790, n74791, n74792, n74793, n74794,
         n74795, n74796, n74797, n74798, n74799, n74800, n74801, n74802,
         n74803, n74804, n74805, n74806, n74807, n74808, n74809, n74810,
         n74811, n74812, n74813, n74814, n74815, n74816, n74817, n74818,
         n74819, n74820, n74821, n74822, n74823, n74824, n74825, n74826,
         n74827, n74828, n74829, n74830, n74831, n74832, n74833, n74834,
         n74835, n74836, n74837, n74838, n74839, n74840, n74841, n74842,
         n74843, n74844, n74845, n74846, n74847, n74848, n74849, n74850,
         n74851, n74852, n74853, n74854, n74855, n74856, n74857, n74858,
         n74859, n74860, n74861, n74862, n74863, n74864, n74865, n74866,
         n74867, n74868, n74869, n74870, n74871, n74872, n74873, n74874,
         n74875, n74876, n74877, n74878, n74879, n74880, n74881, n74882,
         n74883, n74884, n74885, n74886, n74887, n74888, n74889, n74890,
         n74891, n74892, n74893, n74894, n74895, n74896, n74897, n74898,
         n74899, n74900, n74901, n74902, n74903, n74904, n74905, n74906,
         n74907, n74908, n74909, n74910, n74911, n74912, n74913, n74914,
         n74915, n74916, n74917, n74918, n74919, n74920, n74921, n74922,
         n74923, n74924, n74925, n74926, n74927, n74928, n74929, n74930,
         n74931, n74932, n74933, n74934, n74935, n74936, n74937, n74938,
         n74939, n74940, n74941, n74942, n74943, n74944, n74945, n74946,
         n74947, n74948, n74949, n74950, n74951, n74952, n74953, n74954,
         n74955, n74956, n74957, n74958, n74959, n74960, n74961, n74962,
         n74963, n74964, n74965, n74966, n74967, n74968, n74969, n74970,
         n74971, n74972, n74973, n74974, n74975, n74976, n74977, n74978,
         n74979, n74980, n74981, n74982, n74983, n74984, n74985, n74986,
         n74987, n74988, n74989, n74990, n74991, n74992, n74993, n74994,
         n74995, n74996, n74997, n74998, n74999, n75000, n75001, n75002,
         n75003, n75004, n75005, n75006, n75007, n75008, n75009, n75010,
         n75011, n75012, n75013, n75014, n75015, n75016, n75017, n75018,
         n75019, n75020, n75021, n75022, n75023, n75024, n75025, n75026,
         n75027, n75028, n75029, n75030, n75031, n75032, n75033, n75034,
         n75035, n75036, n75037, n75038, n75039, n75040, n75041, n75042,
         n75043, n75044, n75045, n75046, n75047, n75048, n75049, n75050,
         n75051, n75052, n75053, n75054, n75055, n75056, n75057, n75058,
         n75059, n75060, n75061, n75062, n75063, n75064, n75065, n75066,
         n75067, n75068, n75069, n75070, n75071, n75072, n75073, n75074,
         n75075, n75076, n75077, n75078, n75079, n75080, n75081, n75082,
         n75083, n75084, n75085, n75086, n75087, n75088, n75089, n75090,
         n75091, n75092, n75093, n75094, n75095, n75096, n75097, n75098,
         n75099, n75100, n75101, n75102, n75103, n75104, n75105, n75106,
         n75107, n75108, n75109, n75110, n75111, n75112, n75113, n75114,
         n75115, n75116, n75117, n75118, n75119, n75120, n75121, n75122,
         n75123, n75124, n75125, n75126, n75127, n75128, n75129, n75130,
         n75131, n75132, n75133, n75134, n75135, n75136, n75137, n75138,
         n75139, n75140, n75141, n75142, n75143, n75144, n75145, n75146,
         n75147, n75148, n75149, n75150, n75151, n75152, n75153, n75154,
         n75155, n75156, n75157, n75158, n75159, n75160, n75161, n75162,
         n75163, n75164, n75165, n75166, n75167, n75168, n75169, n75170,
         n75171, n75172, n75173, n75174, n75175, n75176, n75177, n75178,
         n75179, n75180, n75181, n75182, n75183, n75184, n75185, n75186,
         n75187, n75188, n75189, n75190, n75191, n75192, n75193, n75194,
         n75195, n75196, n75197, n75198, n75199, n75200, n75201, n75202,
         n75203, n75204, n75205, n75206, n75207, n75208, n75209, n75210,
         n75211, n75212, n75213, n75214, n75215, n75216, n75217, n75218,
         n75219, n75220, n75221, n75222, n75223, n75224, n75225, n75226,
         n75227, n75228, n75229, n75230, n75231, n75232, n75233, n75234,
         n75235, n75236, n75237, n75238, n75239, n75240, n75241, n75242,
         n75243, n75244, n75245, n75246, n75247, n75248, n75249, n75250,
         n75251, n75252, n75253, n75254, n75255, n75256, n75257, n75258,
         n75259, n75260, n75261, n75262, n75263, n75264, n75265, n75266,
         n75267, n75268, n75269, n75270, n75271, n75272, n75273, n75274,
         n75275, n75276, n75277, n75278, n75279, n75280, n75281, n75282,
         n75283, n75284, n75285, n75286, n75287, n75288, n75289, n75290,
         n75291, n75292, n75293, n75294, n75295, n75296, n75297, n75298,
         n75299, n75300, n75301, n75302, n75303, n75304, n75305, n75306,
         n75307, n75308, n75309, n75310, n75311, n75312, n75313, n75314,
         n75315, n75316, n75317, n75318, n75319, n75320, n75321, n75322,
         n75323, n75324, n75325, n75326, n75327, n75328, n75329, n75330,
         n75331, n75332, n75333, n75334, n75335, n75336, n75337, n75338,
         n75339, n75340, n75341, n75342, n75343, n75344, n75345, n75346,
         n75347, n75348, n75349, n75350, n75351, n75352, n75353, n75354,
         n75355, n75356, n75357, n75358, n75359, n75360, n75361, n75362,
         n75363, n75364, n75365, n75366, n75367, n75368, n75369, n75370,
         n75371, n75372, n75373, n75374, n75375, n75376, n75377, n75378,
         n75379, n75380, n75381, n75382, n75383, n75384, n75385, n75386,
         n75387, n75388, n75389, n75390, n75391, n75392, n75393, n75394,
         n75395, n75396, n75397, n75398, n75399, n75400, n75401, n75402,
         n75403, n75404, n75405, n75406, n75407, n75408, n75409, n75410,
         n75411, n75412, n75413, n75414, n75415, n75416, n75417, n75418,
         n75419, n75420, n75421, n75422, n75423, n75424, n75425, n75426,
         n75427, n75428, n75429, n75430, n75431, n75432, n75433, n75434,
         n75435, n75436, n75437, n75438, n75439, n75440, n75441, n75442,
         n75443, n75444, n75445, n75446, n75447, n75448, n75449, n75450,
         n75451, n75452, n75453, n75454, n75455, n75456, n75457, n75458,
         n75459, n75460, n75461, n75462, n75463, n75464, n75465, n75466,
         n75467, n75468, n75469, n75470, n75471, n75472, n75473, n75474,
         n75475, n75476, n75477, n75478, n75479, n75480, n75481, n75482,
         n75483, n75484, n75485, n75486, n75487, n75488, n75489, n75490,
         n75491, n75492, n75493, n75494, n75495, n75496, n75497, n75498,
         n75499, n75500, n75501, n75502, n75503, n75504, n75505, n75506,
         n75507, n75508, n75509, n75510, n75511, n75512, n75513, n75514,
         n75515, n75516, n75517, n75518, n75519, n75520, n75521, n75522,
         n75523, n75524, n75525, n75526, n75527, n75528, n75529, n75530,
         n75531, n75532, n75533, n75534, n75535, n75536, n75537, n75538,
         n75539, n75540, n75541, n75542, n75543, n75544, n75545, n75546,
         n75547, n75548, n75549, n75550, n75551, n75552, n75553, n75554,
         n75555, n75556, n75557, n75558, n75559, n75560, n75561, n75562,
         n75563, n75564, n75565, n75566, n75567, n75568, n75569, n75570,
         n75571, n75572, n75573, n75574, n75575, n75576, n75577, n75578,
         n75579, n75580, n75581, n75582, n75583, n75584, n75585, n75586,
         n75587, n75588, n75589, n75590, n75591, n75592, n75593, n75594,
         n75595, n75596, n75597, n75598, n75599, n75600, n75601, n75602,
         n75603, n75604, n75605, n75606, n75607, n75608, n75609, n75610,
         n75611, n75612, n75613, n75614, n75615, n75616, n75617, n75618,
         n75619, n75620, n75621, n75622, n75623, n75624, n75625, n75626,
         n75627, n75628, n75629, n75630, n75631, n75632, n75633, n75634,
         n75635, n75636, n75637, n75638, n75639, n75640, n75641, n75642,
         n75643, n75644, n75645, n75646, n75647, n75648, n75649, n75650,
         n75651, n75652, n75653, n75654, n75655, n75656, n75657, n75658,
         n75659, n75660, n75661, n75662, n75663, n75664, n75665, n75666,
         n75667, n75668, n75669, n75670, n75671, n75672, n75673, n75674,
         n75675, n75676, n75677, n75678, n75679, n75680, n75681, n75682,
         n75683, n75684, n75685, n75686, n75687, n75688, n75689, n75690,
         n75691, n75692, n75693, n75694, n75695, n75696, n75697, n75698,
         n75699, n75700, n75701, n75702, n75703, n75704, n75705, n75706,
         n75707, n75708, n75709, n75710, n75711, n75712, n75713, n75714,
         n75715, n75716, n75717, n75718, n75719, n75720, n75721, n75722,
         n75723, n75724, n75725, n75726, n75727, n75728, n75729, n75730,
         n75731, n75732, n75733, n75734, n75735, n75736, n75737, n75738,
         n75739, n75740, n75741, n75742, n75743, n75744, n75745, n75746,
         n75747, n75748, n75749, n75750, n75751, n75752, n75753, n75754,
         n75755, n75756, n75757, n75758, n75759, n75760, n75761, n75762,
         n75763, n75764, n75765, n75766, n75767, n75768, n75769, n75770,
         n75771, n75772, n75773, n75774, n75775, n75776, n75777, n75778,
         n75779, n75780, n75781, n75782, n75783, n75784, n75785, n75786,
         n75787, n75788, n75789, n75790, n75791, n75792, n75793, n75794,
         n75795, n75796, n75797, n75798, n75799, n75800, n75801, n75802,
         n75803, n75804, n75805, n75806, n75807, n75808, n75809, n75810,
         n75811, n75812, n75813, n75814, n75815, n75816, n75817, n75818,
         n75819, n75820, n75821, n75822, n75823, n75824, n75825, n75826,
         n75827, n75828, n75829, n75830, n75831, n75832, n75833, n75834,
         n75835, n75836, n75837, n75838, n75839, n75840, n75841, n75842,
         n75843, n75844, n75845, n75846, n75847, n75848, n75849, n75850,
         n75851, n75852, n75853, n75854, n75855, n75856, n75857, n75858,
         n75859, n75860, n75861, n75862, n75863, n75864, n75865, n75866,
         n75867, n75868, n75869, n75870, n75871, n75872, n75873, n75874,
         n75875, n75876, n75877, n75878, n75879, n75880, n75881, n75882,
         n75883, n75884, n75885, n75886, n75887, n75888, n75889, n75890,
         n75891, n75892, n75893, n75894, n75895, n75896, n75897, n75898,
         n75899, n75900, n75901, n75902, n75903, n75904, n75905, n75906,
         n75907, n75908, n75909, n75910, n75911, n75912, n75913, n75914,
         n75915, n75916, n75917, n75918, n75919, n75920, n75921, n75922,
         n75923, n75924, n75925, n75926, n75927, n75928, n75929, n75930,
         n75931, n75932, n75933, n75934, n75935, n75936, n75937, n75938,
         n75939, n75940, n75941, n75942, n75943, n75944, n75945, n75946,
         n75947, n75948, n75949, n75950, n75951, n75952, n75953, n75954,
         n75955, n75956, n75957, n75958, n75959, n75960, n75961, n75962,
         n75963, n75964, n75965, n75966, n75967, n75968, n75969, n75970,
         n75971, n75972, n75973, n75974, n75975, n75976, n75977, n75978,
         n75979, n75980, n75981, n75982, n75983, n75984, n75985, n75986,
         n75987, n75988, n75989, n75990, n75991, n75992, n75993, n75994,
         n75995, n75996, n75997, n75998, n75999, n76000, n76001, n76002,
         n76003, n76004, n76005, n76006, n76007, n76008, n76009, n76010,
         n76011, n76012, n76013, n76014, n76015, n76016, n76017, n76018,
         n76019, n76020, n76021, n76022, n76023, n76024, n76025, n76026,
         n76027, n76028, n76029, n76030, n76031, n76032, n76033, n76034,
         n76035, n76036, n76037, n76038, n76039, n76040, n76041, n76042,
         n76043, n76044, n76045, n76046, n76047, n76048, n76049, n76050,
         n76051, n76052, n76053, n76054, n76055, n76056, n76057, n76058,
         n76059, n76060, n76061, n76062, n76063, n76064, n76065, n76066,
         n76067, n76068, n76069, n76070, n76071, n76072, n76073, n76074,
         n76075, n76076, n76077, n76078, n76079, n76080, n76081, n76082,
         n76083, n76084, n76085, n76086, n76087, n76088, n76089, n76090,
         n76091, n76092, n76093, n76094, n76095, n76096, n76097, n76098,
         n76099, n76100, n76101, n76102, n76103, n76104, n76105, n76106,
         n76107, n76108, n76109, n76110, n76111, n76112, n76113, n76114,
         n76115, n76116, n76117, n76118, n76119, n76120, n76121, n76122,
         n76123, n76124, n76125, n76126, n76127, n76128, n76129, n76130,
         n76131, n76132, n76133, n76134, n76135, n76136, n76137, n76138,
         n76139, n76140, n76141, n76142, n76143, n76144, n76145, n76146,
         n76147, n76148, n76149, n76150, n76151, n76152, n76153, n76154,
         n76155, n76156, n76157, n76158, n76159, n76160, n76161, n76162,
         n76163, n76164, n76165, n76166, n76167, n76168, n76169, n76170,
         n76171, n76172, n76173, n76174, n76175, n76176, n76177, n76178,
         n76179, n76180, n76181, n76182, n76183, n76184, n76185, n76186,
         n76187, n76188, n76189, n76190, n76191, n76192, n76193, n76194,
         n76195, n76196, n76197, n76198, n76199, n76200, n76201, n76202,
         n76203, n76204, n76205, n76206, n76207, n76208, n76209, n76210,
         n76211, n76212, n76213, n76214, n76215, n76216, n76217, n76218,
         n76219, n76220, n76221, n76222, n76223, n76224, n76225, n76226,
         n76227, n76228, n76229, n76230, n76231, n76232, n76233, n76234,
         n76235, n76236, n76237, n76238, n76239, n76240, n76241, n76242,
         n76243, n76244, n76245, n76246, n76247, n76248, n76249, n76250,
         n76251, n76252, n76253, n76254, n76255, n76256, n76257, n76258,
         n76259, n76260, n76261, n76262, n76263, n76264, n76265, n76266,
         n76267, n76268, n76269, n76270, n76271, n76272, n76273, n76274,
         n76275, n76276, n76277, n76278, n76279, n76280, n76281, n76282,
         n76283, n76284, n76285, n76286, n76287, n76288, n76289, n76290,
         n76291, n76292, n76293, n76294, n76295, n76296, n76297, n76298,
         n76299, n76300, n76301, n76302, n76303, n76304, n76305, n76306,
         n76307, n76308, n76309, n76310, n76311, n76312, n76313, n76314,
         n76315, n76316, n76317, n76318, n76319, n76320, n76321, n76322,
         n76323, n76324, n76325, n76326, n76327, n76328, n76329, n76330,
         n76331, n76332, n76333, n76334, n76335, n76336, n76337, n76338,
         n76339, n76340, n76341, n76342, n76343, n76344, n76345, n76346,
         n76347, n76348, n76349, n76350, n76351, n76352, n76353, n76354,
         n76355, n76356, n76357, n76358, n76359, n76360, n76361, n76362,
         n76363, n76364, n76365, n76366, n76367, n76368, n76369, n76370,
         n76371, n76372, n76373, n76374, n76375, n76376, n76377, n76378,
         n76379, n76380, n76381, n76382, n76383, n76384, n76385, n76386,
         n76387, n76388, n76389, n76390, n76391, n76392, n76393, n76394,
         n76395, n76396, n76397, n76398, n76399, n76400, n76401, n76402,
         n76403, n76404, n76405, n76406, n76407, n76408, n76409, n76410,
         n76411, n76412, n76413, n76414, n76415, n76416, n76417, n76418,
         n76419, n76420, n76421, n76422, n76423, n76424, n76425, n76426,
         n76427, n76428, n76429, n76430, n76431, n76432, n76433, n76434,
         n76435, n76436, n76437, n76438, n76439, n76440, n76441, n76442,
         n76443, n76444, n76445, n76446, n76447, n76448, n76449, n76450,
         n76451, n76452, n76453, n76454, n76455, n76456, n76457, n76458,
         n76459, n76460, n76461, n76462, n76463, n76464, n76465, n76466,
         n76467, n76468, n76469, n76470, n76471, n76472, n76473, n76474,
         n76475, n76476, n76477, n76478, n76479, n76480, n76481, n76482,
         n76483, n76484, n76485, n76486, n76487, n76488, n76489, n76490,
         n76491, n76492, n76493, n76494, n76495, n76496, n76497, n76498,
         n76499, n76500, n76501, n76502, n76503, n76504, n76505, n76506,
         n76507, n76508, n76509, n76510, n76511, n76512, n76513, n76514,
         n76515, n76516, n76517, n76518, n76519, n76520, n76521, n76522,
         n76523, n76524, n76525, n76526, n76527, n76528, n76529, n76530,
         n76531, n76532, n76533, n76534, n76535, n76536, n76537, n76538,
         n76539, n76540, n76541, n76542, n76543, n76544, n76545, n76546,
         n76547, n76548, n76549, n76550, n76551, n76552, n76553, n76554,
         n76555, n76556, n76557, n76558, n76559, n76560, n76561, n76562,
         n76563, n76564, n76565, n76566, n76567, n76568, n76569, n76570,
         n76571, n76572, n76573, n76574, n76575, n76576, n76577, n76578,
         n76579, n76580, n76581, n76582, n76583, n76584, n76585, n76586,
         n76587, n76588, n76589, n76590, n76591, n76592, n76593, n76594,
         n76595, n76596, n76597, n76598, n76599, n76600, n76601, n76602,
         n76603, n76604, n76605, n76606, n76607, n76608, n76609, n76610,
         n76611, n76612, n76613, n76614, n76615, n76616, n76617, n76618,
         n76619, n76620, n76621, n76622, n76623, n76624, n76625, n76626,
         n76627, n76628, n76629, n76630, n76631, n76632, n76633, n76634,
         n76635, n76636, n76637, n76638, n76639, n76640, n76641, n76642,
         n76643, n76644, n76645, n76646, n76647, n76648, n76649, n76650,
         n76651, n76652, n76653, n76654, n76655, n76656, n76657, n76658,
         n76659, n76660, n76661, n76662, n76663, n76664, n76665, n76666,
         n76667, n76668, n76669, n76670, n76671, n76672, n76673, n76674,
         n76675, n76676, n76677, n76678, n76679, n76680, n76681, n76682,
         n76683, n76684, n76685, n76686, n76687, n76688, n76689, n76690,
         n76691, n76692, n76693, n76694, n76695, n76696, n76697, n76698,
         n76699, n76700, n76701, n76702, n76703, n76704, n76705, n76706,
         n76707, n76708, n76709, n76710, n76711, n76712, n76713, n76714,
         n76715, n76716, n76717, n76718, n76719, n76720, n76721, n76722,
         n76723, n76724, n76725, n76726, n76727, n76728, n76729, n76730,
         n76731, n76732, n76733, n76734, n76735, n76736, n76737, n76738,
         n76739, n76740, n76741, n76742, n76743, n76744, n76745, n76746,
         n76747, n76748, n76749, n76750, n76751, n76752, n76753, n76754,
         n76755, n76756, n76757, n76758, n76759, n76760, n76761, n76762,
         n76763, n76764, n76765, n76766, n76767, n76768, n76769, n76770,
         n76771, n76772, n76773, n76774, n76775, n76776, n76777, n76778,
         n76779, n76780, n76781, n76782, n76783, n76784, n76785, n76786,
         n76787, n76788, n76789, n76790, n76791, n76792, n76793, n76794,
         n76795, n76796, n76797, n76798, n76799, n76800, n76801, n76802,
         n76803, n76804, n76805, n76806, n76807, n76808, n76809, n76810,
         n76811, n76812, n76813, n76814, n76815, n76816, n76817, n76818,
         n76819, n76820, n76821, n76822, n76823, n76824, n76825, n76826,
         n76827, n76828, n76829, n76830, n76831, n76832, n76833, n76834,
         n76835, n76836, n76837, n76838, n76839, n76840, n76841, n76842,
         n76843, n76844, n76845, n76846, n76847, n76848, n76849, n76850,
         n76851, n76852, n76853, n76854, n76855, n76856, n76857, n76858,
         n76859, n76860, n76861, n76862, n76863, n76864, n76865, n76866,
         n76867, n76868, n76869, n76870, n76871, n76872, n76873, n76874,
         n76875, n76876, n76877, n76878, n76879, n76880, n76881, n76882,
         n76883, n76884, n76885, n76886, n76887, n76888, n76889, n76890,
         n76891, n76892, n76893, n76894, n76895, n76896, n76897, n76898,
         n76899, n76900, n76901, n76902, n76903, n76904, n76905, n76906,
         n76907, n76908, n76909, n76910, n76911, n76912, n76913, n76914,
         n76915, n76916, n76917, n76918, n76919, n76920, n76921, n76922,
         n76923, n76924, n76925, n76926, n76927, n76928, n76929, n76930,
         n76931, n76932, n76933, n76934, n76935, n76936, n76937, n76938,
         n76939, n76940, n76941, n76942, n76943, n76944, n76945, n76946,
         n76947, n76948, n76949, n76950, n76951, n76952, n76953, n76954,
         n76955, n76956, n76957, n76958, n76959, n76960, n76961, n76962,
         n76963, n76964, n76965, n76966, n76967, n76968, n76969, n76970,
         n76971, n76972, n76973, n76974, n76975, n76976, n76977, n76978,
         n76979, n76980, n76981, n76982, n76983, n76984, n76985, n76986,
         n76987, n76988, n76989, n76990, n76991, n76992, n76993, n76994,
         n76995, n76996, n76997, n76998, n76999, n77000, n77001, n77002,
         n77003, n77004, n77005, n77006, n77007, n77008, n77009, n77010,
         n77011, n77012, n77013, n77014, n77015, n77016, n77017, n77018,
         n77019, n77020, n77021, n77022, n77023, n77024, n77025, n77026,
         n77027, n77028, n77029, n77030, n77031, n77032, n77033, n77034,
         n77035, n77036, n77037, n77038, n77039, n77040, n77041, n77042,
         n77043, n77044, n77045, n77046, n77047, n77048, n77049, n77050,
         n77051, n77052, n77053, n77054, n77055, n77056, n77057, n77058,
         n77059, n77060, n77061, n77062, n77063, n77064, n77065, n77066,
         n77067, n77068, n77069, n77070, n77071, n77072, n77073, n77074,
         n77075, n77076, n77077, n77078, n77079, n77080, n77081, n77082,
         n77083, n77084, n77085, n77086, n77087, n77088, n77089, n77090,
         n77091, n77092, n77093, n77094, n77095, n77096, n77097, n77098,
         n77099, n77100, n77101, n77102, n77103, n77104, n77105, n77106,
         n77107, n77108, n77109, n77110, n77111, n77112, n77113, n77114,
         n77115, n77116, n77117, n77118, n77119, n77120, n77121, n77122,
         n77123, n77124, n77125, n77126, n77127, n77128, n77129, n77130,
         n77131, n77132, n77133, n77134, n77135, n77136, n77137, n77138,
         n77139, n77140, n77141, n77142, n77143, n77144, n77145, n77146,
         n77147, n77148, n77149, n77150, n77151, n77152, n77153, n77154,
         n77155, n77156, n77157, n77158, n77159, n77160, n77161, n77162,
         n77163, n77164, n77165, n77166, n77167, n77168, n77169, n77170,
         n77171, n77172, n77173, n77174, n77175, n77176, n77177, n77178,
         n77179, n77180, n77181, n77182, n77183, n77184, n77185, n77186,
         n77187, n77188, n77189, n77190, n77191, n77192, n77193, n77194,
         n77195, n77196, n77197, n77198, n77199, n77200, n77201, n77202,
         n77203, n77204, n77205, n77206, n77207, n77208, n77209, n77210,
         n77211, n77212, n77213, n77214, n77215, n77216, n77217, n77218,
         n77219, n77220, n77221, n77222, n77223, n77224, n77225, n77226,
         n77227, n77228, n77229, n77230, n77231, n77232, n77233, n77234,
         n77235, n77236, n77237, n77238, n77239, n77240, n77241, n77242,
         n77243, n77244, n77245, n77246, n77247, n77248, n77249, n77250,
         n77251, n77252, n77253, n77254, n77255, n77256, n77257, n77258,
         n77259, n77260, n77261, n77262, n77263, n77264, n77265, n77266,
         n77267, n77268, n77269, n77270, n77271, n77272, n77273, n77274,
         n77275, n77276, n77277, n77278, n77279, n77280, n77281, n77282,
         n77283, n77284, n77285, n77286, n77287, n77288, n77289, n77290,
         n77291, n77292, n77293, n77294, n77295, n77296, n77297, n77298,
         n77299, n77300, n77301, n77302, n77303, n77304, n77305, n77306,
         n77307, n77308, n77309, n77310, n77311, n77312, n77313, n77314,
         n77315, n77316, n77317, n77318, n77319, n77320, n77321, n77322,
         n77323, n77324, n77325, n77326, n77327, n77328, n77329, n77330,
         n77331, n77332, n77333, n77334, n77335, n77336, n77337, n77338,
         n77339, n77340, n77341, n77342, n77343, n77344, n77345, n77346,
         n77347, n77348, n77349, n77350, n77351, n77352, n77353, n77354,
         n77355, n77356, n77357, n77358, n77359, n77360, n77361, n77362,
         n77363, n77364, n77365, n77366, n77367, n77368, n77369, n77370,
         n77371, n77372, n77373, n77374, n77375, n77376, n77377, n77378,
         n77379, n77380, n77381, n77382, n77383, n77384, n77385, n77386,
         n77387, n77388, n77389, n77390, n77391, n77392, n77393, n77394,
         n77395, n77396, n77397, n77398, n77399, n77400, n77401, n77402,
         n77403, n77404, n77405, n77406, n77407, n77408, n77409, n77410,
         n77411, n77412, n77413, n77414, n77415, n77416, n77417, n77418,
         n77419, n77420, n77421, n77422, n77423, n77424, n77425, n77426,
         n77427, n77428, n77429, n77430, n77431, n77432, n77433, n77434,
         n77435, n77436, n77437, n77438, n77439, n77440, n77441, n77442,
         n77443, n77444, n77445, n77446, n77447, n77448, n77449, n77450,
         n77451, n77452, n77453, n77454, n77455, n77456, n77457, n77458,
         n77459, n77460, n77461, n77462, n77463, n77464, n77465, n77466,
         n77467, n77468, n77469, n77470, n77471, n77472, n77473, n77474,
         n77475, n77476, n77477, n77478, n77479, n77480, n77481, n77482,
         n77483, n77484, n77485, n77486, n77487, n77488, n77489, n77490,
         n77491, n77492, n77493, n77494, n77495, n77496, n77497, n77498,
         n77499, n77500, n77501, n77502, n77503, n77504, n77505, n77506,
         n77507, n77508, n77509, n77510, n77511, n77512, n77513, n77514,
         n77515, n77516, n77517, n77518, n77519, n77520, n77521, n77522,
         n77523, n77524, n77525, n77526, n77527, n77528, n77529, n77530,
         n77531, n77532, n77533, n77534, n77535, n77536, n77537, n77538,
         n77539, n77540, n77541, n77542, n77543, n77544, n77545, n77546,
         n77547, n77548, n77549, n77550, n77551, n77552, n77553, n77554,
         n77555, n77556, n77557, n77558, n77559, n77560, n77561, n77562,
         n77563, n77564, n77565, n77566, n77567, n77568, n77569, n77570,
         n77571, n77572, n77573, n77574, n77575, n77576, n77577, n77578,
         n77579, n77580, n77581, n77582, n77583, n77584, n77585, n77586,
         n77587, n77588, n77589, n77590, n77591, n77592, n77593, n77594,
         n77595, n77596, n77597, n77598, n77599, n77600, n77601, n77602,
         n77603, n77604, n77605, n77606, n77607, n77608, n77609, n77610,
         n77611, n77612, n77613, n77614, n77615, n77616, n77617, n77618,
         n77619, n77620, n77621, n77622, n77623, n77624, n77625, n77626,
         n77627, n77628, n77629, n77630, n77631, n77632, n77633, n77634,
         n77635, n77636, n77637, n77638, n77639, n77640, n77641, n77642,
         n77643, n77644, n77645, n77646, n77647, n77648, n77649, n77650,
         n77651, n77652, n77653, n77654, n77655, n77656, n77657, n77658,
         n77659, n77660, n77661, n77662, n77663, n77664, n77665, n77666,
         n77667, n77668, n77669, n77670, n77671, n77672, n77673, n77674,
         n77675, n77676, n77677, n77678, n77679, n77680, n77681, n77682,
         n77683, n77684, n77685, n77686, n77687, n77688, n77689, n77690,
         n77691, n77692, n77693, n77694, n77695, n77696, n77697, n77698,
         n77699, n77700, n77701, n77702, n77703, n77704, n77705, n77706,
         n77707, n77708, n77709, n77710, n77711, n77712, n77713, n77714,
         n77715, n77716, n77717, n77718, n77719, n77720, n77721, n77722,
         n77723, n77724, n77725, n77726, n77727, n77728, n77729, n77730,
         n77731, n77732, n77733, n77734, n77735, n77736, n77737, n77738,
         n77739, n77740, n77741, n77742, n77743, n77744, n77745, n77746,
         n77747, n77748, n77749, n77750, n77751, n77752, n77753, n77754,
         n77755, n77756, n77757, n77758, n77759, n77760, n77761, n77762,
         n77763, n77764, n77765, n77766, n77767, n77768, n77769, n77770,
         n77771, n77772, n77773, n77774, n77775, n77776, n77777, n77778,
         n77779, n77780, n77781, n77782, n77783, n77784, n77785, n77786,
         n77787, n77788, n77789, n77790, n77791, n77792, n77793, n77794,
         n77795, n77796, n77797, n77798, n77799, n77800, n77801, n77802,
         n77803, n77804, n77805, n77806, n77807, n77808, n77809, n77810,
         n77811, n77812, n77813, n77814, n77815, n77816, n77817, n77818,
         n77819, n77820, n77821, n77822, n77823, n77824, n77825, n77826,
         n77827, n77828, n77829, n77830, n77831, n77832, n77833, n77834,
         n77835, n77836, n77837, n77838, n77839, n77840, n77841, n77842,
         n77843, n77844, n77845, n77846, n77847, n77848, n77849, n77850,
         n77851, n77852, n77853, n77854, n77855, n77856, n77857, n77858,
         n77859, n77860, n77861, n77862, n77863, n77864, n77865, n77866,
         n77867, n77868, n77869, n77870, n77871, n77872, n77873, n77874,
         n77875, n77876, n77877, n77878, n77879, n77880, n77881, n77882,
         n77883, n77884, n77885, n77886, n77887, n77888, n77889, n77890,
         n77891, n77892, n77893, n77894, n77895, n77896, n77897, n77898,
         n77899, n77900, n77901, n77902, n77903, n77904, n77905, n77906,
         n77907, n77908, n77909, n77910, n77911, n77912, n77913, n77914,
         n77915, n77916, n77917, n77918, n77919, n77920, n77921, n77922,
         n77923, n77924, n77925, n77926, n77927, n77928, n77929, n77930,
         n77931, n77932, n77933, n77934, n77935, n77936, n77937, n77938,
         n77939, n77940, n77941, n77942, n77943, n77944, n77945, n77946,
         n77947, n77948, n77949, n77950, n77951, n77952, n77953, n77954,
         n77955, n77956, n77957, n77958, n77959, n77960, n77961, n77962,
         n77963, n77964, n77965, n77966, n77967, n77968, n77969, n77970,
         n77971, n77972, n77973, n77974, n77975, n77976, n77977, n77978,
         n77979, n77980, n77981, n77982, n77983, n77984, n77985, n77986,
         n77987, n77988, n77989, n77990, n77991, n77992, n77993, n77994,
         n77995, n77996, n77997, n77998, n77999, n78000, n78001, n78002,
         n78003, n78004, n78005, n78006, n78007, n78008, n78009, n78010,
         n78011, n78012, n78013, n78014, n78015, n78016, n78017, n78018,
         n78019, n78020, n78021, n78022, n78023, n78024, n78025, n78026,
         n78027, n78028, n78029, n78030, n78031, n78032, n78033, n78034,
         n78035, n78036, n78037, n78038, n78039, n78040, n78041, n78042,
         n78043, n78044, n78045, n78046, n78047, n78048, n78049, n78050,
         n78051, n78052, n78053, n78054, n78055, n78056, n78057, n78058,
         n78059, n78060, n78061, n78062, n78063, n78064, n78065, n78066,
         n78067, n78068, n78069, n78070, n78071, n78072, n78073, n78074,
         n78075, n78076, n78077, n78078, n78079, n78080, n78081, n78082,
         n78083, n78084, n78085, n78086, n78087, n78088, n78089, n78090,
         n78091, n78092, n78093, n78094, n78095, n78096, n78097, n78098,
         n78099, n78100, n78101, n78102, n78103, n78104, n78105, n78106,
         n78107, n78108, n78109, n78110, n78111, n78112, n78113, n78114,
         n78115, n78116, n78117, n78118, n78119, n78120, n78121, n78122,
         n78123, n78124, n78125, n78126, n78127, n78128, n78129, n78130,
         n78131, n78132, n78133, n78134, n78135, n78136, n78137, n78138,
         n78139, n78140, n78141, n78142, n78143, n78144, n78145, n78146,
         n78147, n78148, n78149, n78150, n78151, n78152, n78153, n78154,
         n78155, n78156, n78157, n78158, n78159, n78160, n78161, n78162,
         n78163, n78164, n78165, n78166, n78167, n78168, n78169, n78170,
         n78171, n78172, n78173, n78174, n78175, n78176, n78177, n78178,
         n78179, n78180, n78181, n78182, n78183, n78184, n78185, n78186,
         n78187, n78188, n78189, n78190, n78191, n78192, n78193, n78194,
         n78195, n78196, n78197, n78198, n78199, n78200, n78201, n78202,
         n78203, n78204, n78205, n78206, n78207, n78208, n78209, n78210,
         n78211, n78212, n78213, n78214, n78215, n78216, n78217, n78218,
         n78219, n78220, n78221, n78222, n78223, n78224, n78225, n78226,
         n78227, n78228, n78229, n78230, n78231, n78232, n78233, n78234,
         n78235, n78236, n78237, n78238, n78239, n78240, n78241, n78242,
         n78243, n78244, n78245, n78246, n78247, n78248, n78249, n78250,
         n78251, n78252, n78253, n78254, n78255, n78256, n78257, n78258,
         n78259, n78260, n78261, n78262, n78263, n78264, n78265, n78266,
         n78267, n78268, n78269, n78270, n78271, n78272, n78273, n78274,
         n78275, n78276, n78277, n78278, n78279, n78280, n78281, n78282,
         n78283, n78284, n78285, n78286, n78287, n78288, n78289, n78290,
         n78291, n78292, n78293, n78294, n78295, n78296, n78297, n78298,
         n78299, n78300, n78301, n78302, n78303, n78304, n78305, n78306,
         n78307, n78308, n78309, n78310, n78311, n78312, n78313, n78314,
         n78315, n78316, n78317, n78318, n78319, n78320, n78321, n78322,
         n78323, n78324, n78325, n78326, n78327, n78328, n78329, n78330,
         n78331, n78332, n78333, n78334, n78335, n78336, n78337, n78338,
         n78339, n78340, n78341, n78342, n78343, n78344, n78345, n78346,
         n78347, n78348, n78349, n78350, n78351, n78352, n78353, n78354,
         n78355, n78356, n78357, n78358, n78359, n78360, n78361, n78362,
         n78363, n78364, n78365, n78366, n78367, n78368, n78369, n78370,
         n78371, n78372, n78373, n78374, n78375, n78376, n78377, n78378,
         n78379, n78380, n78381, n78382, n78383, n78384, n78385, n78386,
         n78387, n78388, n78389, n78390, n78391, n78392, n78393, n78394,
         n78395, n78396, n78397, n78398, n78399, n78400, n78401, n78402,
         n78403, n78404, n78405, n78406, n78407, n78408, n78409, n78410,
         n78411, n78412, n78413, n78414, n78415, n78416, n78417, n78418,
         n78419, n78420, n78421, n78422, n78423, n78424, n78425, n78426,
         n78427, n78428, n78429, n78430, n78431, n78432, n78433, n78434,
         n78435, n78436, n78437, n78438, n78439, n78440, n78441, n78442,
         n78443, n78444, n78445, n78446, n78447, n78448, n78449, n78450,
         n78451, n78452, n78453, n78454, n78455, n78456, n78457, n78458,
         n78459, n78460, n78461, n78462, n78463, n78464, n78465, n78466,
         n78467, n78468, n78469, n78470, n78471, n78472, n78473, n78474,
         n78475, n78476, n78477, n78478, n78479, n78480, n78481, n78482,
         n78483, n78484, n78485, n78486, n78487, n78488, n78489, n78490,
         n78491, n78492, n78493, n78494, n78495, n78496, n78497, n78498,
         n78499, n78500, n78501, n78502, n78503, n78504, n78505, n78506,
         n78507, n78508, n78509, n78510, n78511, n78512, n78513, n78514,
         n78515, n78516, n78517, n78518, n78519, n78520, n78521, n78522,
         n78523, n78524, n78525, n78526, n78527, n78528, n78529, n78530,
         n78531, n78532, n78533, n78534, n78535, n78536, n78537, n78538,
         n78539, n78540, n78541, n78542, n78543, n78544, n78545, n78546,
         n78547, n78548, n78549, n78550, n78551, n78552, n78553, n78554,
         n78555, n78556, n78557, n78558, n78559, n78560, n78561, n78562,
         n78563, n78564, n78565, n78566, n78567, n78568, n78569, n78570,
         n78571, n78572, n78573, n78574, n78575, n78576, n78577, n78578,
         n78579, n78580, n78581, n78582, n78583, n78584, n78585, n78586,
         n78587, n78588, n78589, n78590, n78591, n78592, n78593, n78594,
         n78595, n78596, n78597, n78598, n78599, n78600, n78601, n78602,
         n78603, n78604, n78605, n78606, n78607, n78608, n78609, n78610,
         n78611, n78612, n78613, n78614, n78615, n78616, n78617, n78618,
         n78619, n78620, n78621, n78622, n78623, n78624, n78625, n78626,
         n78627, n78628, n78629, n78630, n78631, n78632, n78633, n78634,
         n78635, n78636, n78637, n78638, n78639, n78640, n78641, n78642,
         n78643, n78644, n78645, n78646, n78647, n78648, n78649, n78650,
         n78651, n78652, n78653, n78654, n78655, n78656, n78657, n78658,
         n78659, n78660, n78661, n78662, n78663, n78664, n78665, n78666,
         n78667, n78668, n78669, n78670, n78671, n78672, n78673, n78674,
         n78675, n78676, n78677, n78678, n78679, n78680, n78681, n78682,
         n78683, n78684, n78685, n78686, n78687, n78688, n78689, n78690,
         n78691, n78692, n78693, n78694, n78695, n78696, n78697, n78698,
         n78699, n78700, n78701, n78702, n78703, n78704, n78705, n78706,
         n78707, n78708, n78709, n78710, n78711, n78712, n78713, n78714,
         n78715, n78716, n78717, n78718, n78719, n78720, n78721, n78722,
         n78723, n78724, n78725, n78726, n78727, n78728, n78729, n78730,
         n78731, n78732, n78733, n78734, n78735, n78736, n78737, n78738,
         n78739, n78740, n78741, n78742, n78743, n78744, n78745, n78746,
         n78747, n78748, n78749, n78750, n78751, n78752, n78753, n78754,
         n78755, n78756, n78757, n78758, n78759, n78760, n78761, n78762,
         n78763, n78764, n78765, n78766, n78767, n78768, n78769, n78770,
         n78771, n78772, n78773, n78774, n78775, n78776, n78777, n78778,
         n78779, n78780, n78781, n78782, n78783, n78784, n78785, n78786,
         n78787, n78788, n78789, n78790, n78791, n78792, n78793, n78794,
         n78795, n78796, n78797, n78798, n78799, n78800, n78801, n78802,
         n78803, n78804, n78805, n78806, n78807, n78808, n78809, n78810,
         n78811, n78812, n78813, n78814, n78815, n78816, n78817, n78818,
         n78819, n78820, n78821, n78822, n78823, n78824, n78825, n78826,
         n78827, n78828, n78829, n78830, n78831, n78832, n78833, n78834,
         n78835, n78836, n78837, n78838, n78839, n78840, n78841, n78842,
         n78843, n78844, n78845, n78846, n78847, n78848, n78849, n78850,
         n78851, n78852, n78853, n78854, n78855, n78856, n78857, n78858,
         n78859, n78860, n78861, n78862, n78863, n78864, n78865, n78866,
         n78867, n78868, n78869, n78870, n78871, n78872, n78873, n78874,
         n78875, n78876, n78877, n78878, n78879, n78880, n78881, n78882,
         n78883, n78884, n78885, n78886, n78887, n78888, n78889, n78890,
         n78891, n78892, n78893, n78894, n78895, n78896, n78897, n78898,
         n78899, n78900, n78901, n78902, n78903, n78904, n78905, n78906,
         n78907, n78908, n78909, n78910, n78911, n78912, n78913, n78914,
         n78915, n78916, n78917, n78918, n78919, n78920, n78921, n78922,
         n78923, n78924, n78925, n78926, n78927, n78928, n78929, n78930,
         n78931, n78932, n78933, n78934, n78935, n78936, n78937, n78938,
         n78939, n78940, n78941, n78942, n78943, n78944, n78945, n78946,
         n78947, n78948, n78949, n78950, n78951, n78952, n78953, n78954,
         n78955, n78956, n78957, n78958, n78959, n78960, n78961, n78962,
         n78963, n78964, n78965, n78966, n78967, n78968, n78969, n78970,
         n78971, n78972, n78973, n78974, n78975, n78976, n78977, n78978,
         n78979, n78980, n78981, n78982, n78983, n78984, n78985, n78986,
         n78987, n78988, n78989, n78990, n78991, n78992, n78993, n78994,
         n78995, n78996, n78997, n78998, n78999, n79000, n79001, n79002,
         n79003, n79004, n79005, n79006, n79007, n79008, n79009, n79010,
         n79011, n79012, n79013, n79014, n79015, n79016, n79017, n79018,
         n79019, n79020, n79021, n79022, n79023, n79024, n79025, n79026,
         n79027, n79028, n79029, n79030, n79031, n79032, n79033, n79034,
         n79035, n79036, n79037, n79038, n79039, n79040, n79041, n79042,
         n79043, n79044, n79045, n79046, n79047, n79048, n79049, n79050,
         n79051, n79052, n79053, n79054, n79055, n79056, n79057, n79058,
         n79059, n79060, n79061, n79062, n79063, n79064, n79065, n79066,
         n79067, n79068, n79069, n79070, n79071, n79072, n79073, n79074,
         n79075, n79076, n79077, n79078, n79079, n79080, n79081, n79082,
         n79083, n79084, n79085, n79086, n79087, n79088, n79089, n79090,
         n79091, n79092, n79093, n79094, n79095, n79096, n79097, n79098,
         n79099, n79100, n79101, n79102, n79103, n79104, n79105, n79106,
         n79107, n79108, n79109, n79110, n79111, n79112, n79113, n79114,
         n79115, n79116, n79117, n79118, n79119, n79120, n79121, n79122,
         n79123, n79124, n79125, n79126, n79127, n79128, n79129, n79130,
         n79131, n79132, n79133, n79134, n79135, n79136, n79137, n79138,
         n79139, n79140, n79141, n79142, n79143, n79144, n79145, n79146,
         n79147, n79148, n79149, n79150, n79151, n79152, n79153, n79154,
         n79155, n79156, n79157, n79158, n79159, n79160, n79161, n79162,
         n79163, n79164, n79165, n79166, n79167, n79168, n79169, n79170,
         n79171, n79172, n79173, n79174, n79175, n79176, n79177, n79178,
         n79179, n79180, n79181, n79182, n79183, n79184, n79185, n79186,
         n79187, n79188, n79189, n79190, n79191, n79192, n79193, n79194,
         n79195, n79196, n79197, n79198, n79199, n79200, n79201, n79202,
         n79203, n79204, n79205, n79206, n79207, n79208, n79209, n79210,
         n79211, n79212, n79213, n79214, n79215, n79216, n79217, n79218,
         n79219, n79220, n79221, n79222, n79223, n79224, n79225, n79226,
         n79227, n79228, n79229, n79230, n79231, n79232, n79233, n79234,
         n79235, n79236, n79237, n79238, n79239, n79240, n79241, n79242,
         n79243, n79244, n79245, n79246, n79247, n79248, n79249, n79250,
         n79251, n79252, n79253, n79254, n79255, n79256, n79257, n79258,
         n79259, n79260, n79261, n79262, n79263, n79264, n79265, n79266,
         n79267, n79268, n79269, n79270, n79271, n79272, n79273, n79274,
         n79275, n79276, n79277, n79278, n79279, n79280, n79281, n79282,
         n79283, n79284, n79285, n79286, n79287, n79288, n79289, n79290,
         n79291, n79292, n79293, n79294, n79295, n79296, n79297, n79298,
         n79299, n79300, n79301, n79302, n79303, n79304, n79305, n79306,
         n79307, n79308, n79309, n79310, n79311, n79312, n79313, n79314,
         n79315, n79316, n79317, n79318, n79319, n79320, n79321, n79322,
         n79323, n79324, n79325, n79326, n79327, n79328, n79329, n79330,
         n79331, n79332, n79333, n79334, n79335, n79336, n79337, n79338,
         n79339, n79340, n79341, n79342, n79343, n79344, n79345, n79346,
         n79347, n79348, n79349, n79350, n79351, n79352, n79353, n79354,
         n79355, n79356, n79357, n79358, n79359, n79360, n79361, n79362,
         n79363, n79364, n79365, n79366, n79367, n79368, n79369, n79370,
         n79371, n79372, n79373, n79374, n79375, n79376, n79377, n79378,
         n79379, n79380, n79381, n79382, n79383, n79384, n79385, n79386,
         n79387, n79388, n79389, n79390, n79391, n79392, n79393, n79394,
         n79395, n79396, n79397, n79398, n79399, n79400, n79401, n79402,
         n79403, n79404, n79405, n79406, n79407, n79408, n79409, n79410,
         n79411, n79412, n79413, n79414, n79415, n79416, n79417, n79418,
         n79419, n79420, n79421, n79422, n79423, n79424, n79425, n79426,
         n79427, n79428, n79429, n79430, n79431, n79432, n79433, n79434,
         n79435, n79436, n79437, n79438, n79439, n79440, n79441, n79442,
         n79443, n79444, n79445, n79446, n79447, n79448, n79449, n79450,
         n79451, n79452, n79453, n79454, n79455, n79456, n79457, n79458,
         n79459, n79460, n79461, n79462, n79463, n79464, n79465, n79466,
         n79467, n79468, n79469, n79470, n79471, n79472, n79473, n79474,
         n79475, n79476, n79477, n79478, n79479, n79480, n79481, n79482,
         n79483, n79484, n79485, n79486, n79487, n79488, n79489, n79490,
         n79491, n79492, n79493, n79494, n79495, n79496, n79497, n79498,
         n79499, n79500, n79501, n79502, n79503, n79504, n79505, n79506,
         n79507, n79508, n79509, n79510, n79511, n79512, n79513, n79514,
         n79515, n79516, n79517, n79518, n79519, n79520, n79521, n79522,
         n79523, n79524, n79525, n79526, n79527, n79528, n79529, n79530,
         n79531, n79532, n79533, n79534, n79535, n79536, n79537, n79538,
         n79539, n79540, n79541, n79542, n79543, n79544, n79545, n79546,
         n79547, n79548, n79549, n79550, n79551, n79552, n79553, n79554,
         n79555, n79556, n79557, n79558, n79559, n79560, n79561, n79562,
         n79563, n79564, n79565, n79566, n79567, n79568, n79569, n79570,
         n79571, n79572, n79573, n79574, n79575, n79576, n79577, n79578,
         n79579, n79580, n79581, n79582, n79583, n79584, n79585, n79586,
         n79587, n79588, n79589, n79590, n79591, n79592, n79593, n79594,
         n79595, n79596, n79597, n79598, n79599, n79600, n79601, n79602,
         n79603, n79604, n79605, n79606, n79607, n79608, n79609, n79610,
         n79611, n79612, n79613, n79614, n79615, n79616, n79617, n79618,
         n79619, n79620, n79621, n79622, n79623, n79624, n79625, n79626,
         n79627, n79628, n79629, n79630, n79631, n79632, n79633, n79634,
         n79635, n79636, n79637, n79638, n79639, n79640, n79641, n79642,
         n79643, n79644, n79645, n79646, n79647, n79648, n79649, n79650,
         n79651, n79652, n79653, n79654, n79655, n79656, n79657, n79658,
         n79659, n79660, n79661, n79662, n79663, n79664, n79665, n79666,
         n79667, n79668, n79669, n79670, n79671, n79672, n79673, n79674,
         n79675, n79676, n79677, n79678, n79679, n79680, n79681, n79682,
         n79683, n79684, n79685, n79686, n79687, n79688, n79689, n79690,
         n79691, n79692, n79693, n79694, n79695, n79696, n79697, n79698,
         n79699, n79700, n79701, n79702, n79703, n79704, n79705, n79706,
         n79707, n79708, n79709, n79710, n79711, n79712, n79713, n79714,
         n79715, n79716, n79717, n79718, n79719, n79720, n79721, n79722,
         n79723, n79724, n79725, n79726, n79727, n79728, n79729, n79730,
         n79731, n79732, n79733, n79734, n79735, n79736, n79737, n79738,
         n79739, n79740, n79741, n79742, n79743, n79744, n79745, n79746,
         n79747, n79748, n79749, n79750, n79751, n79752, n79753, n79754,
         n79755, n79756, n79757, n79758, n79759, n79760, n79761, n79762,
         n79763, n79764, n79765, n79766, n79767, n79768, n79769, n79770,
         n79771, n79772, n79773, n79774, n79775, n79776, n79777, n79778,
         n79779, n79780, n79781, n79782, n79783, n79784, n79785, n79786,
         n79787, n79788, n79789, n79790, n79791, n79792, n79793, n79794,
         n79795, n79796, n79797, n79798, n79799, n79800, n79801, n79802,
         n79803, n79804, n79805, n79806, n79807, n79808, n79809, n79810,
         n79811, n79812, n79813, n79814, n79815, n79816, n79817, n79818,
         n79819, n79820, n79821, n79822, n79823, n79824, n79825, n79826,
         n79827, n79828, n79829, n79830, n79831, n79832, n79833, n79834,
         n79835, n79836, n79837, n79838, n79839, n79840, n79841, n79842,
         n79843, n79844, n79845, n79846, n79847, n79848, n79849, n79850,
         n79851, n79852, n79853, n79854, n79855, n79856, n79857, n79858,
         n79859, n79860, n79861, n79862, n79863, n79864, n79865, n79866,
         n79867, n79868, n79869, n79870, n79871, n79872, n79873, n79874,
         n79875, n79876, n79877, n79878, n79879, n79880, n79881, n79882,
         n79883, n79884, n79885, n79886, n79887, n79888, n79889, n79890,
         n79891, n79892, n79893, n79894, n79895, n79896, n79897, n79898,
         n79899, n79900, n79901, n79902, n79903, n79904, n79905, n79906,
         n79907, n79908, n79909, n79910, n79911, n79912, n79913, n79914,
         n79915, n79916, n79917, n79918, n79919, n79920, n79921, n79922,
         n79923, n79924, n79925, n79926, n79927, n79928, n79929, n79930,
         n79931, n79932, n79933, n79934, n79935, n79936, n79937, n79938,
         n79939, n79940, n79941, n79942, n79943, n79944, n79945, n79946,
         n79947, n79948, n79949, n79950, n79951, n79952, n79953, n79954,
         n79955, n79956, n79957, n79958, n79959, n79960, n79961, n79962,
         n79963, n79964, n79965, n79966, n79967, n79968, n79969, n79970,
         n79971, n79972, n79973, n79974, n79975, n79976, n79977, n79978,
         n79979, n79980, n79981, n79982, n79983, n79984, n79985, n79986,
         n79987, n79988, n79989, n79990, n79991, n79992, n79993, n79994,
         n79995, n79996, n79997, n79998, n79999, n80000, n80001, n80002,
         n80003, n80004, n80005, n80006, n80007, n80008, n80009, n80010,
         n80011, n80012, n80013, n80014, n80015, n80016, n80017, n80018,
         n80019, n80020, n80021, n80022, n80023, n80024, n80025, n80026,
         n80027, n80028, n80029, n80030, n80031, n80032, n80033, n80034,
         n80035, n80036, n80037, n80038, n80039, n80040, n80041, n80042,
         n80043, n80044, n80045, n80046, n80047, n80048, n80049, n80050,
         n80051, n80052, n80053, n80054, n80055, n80056, n80057, n80058,
         n80059, n80060, n80061, n80062, n80063, n80064, n80065, n80066,
         n80067, n80068, n80069, n80070, n80071, n80072, n80073, n80074,
         n80075, n80076, n80077, n80078, n80079, n80080, n80081, n80082,
         n80083, n80084, n80085, n80086, n80087, n80088, n80089, n80090,
         n80091, n80092, n80093, n80094, n80095, n80096, n80097, n80098,
         n80099, n80100, n80101, n80102, n80103, n80104, n80105, n80106,
         n80107, n80108, n80109, n80110, n80111, n80112, n80113, n80114,
         n80115, n80116, n80117, n80118, n80119, n80120, n80121, n80122,
         n80123, n80124, n80125, n80126, n80127, n80128, n80129, n80130,
         n80131, n80132, n80133, n80134, n80135, n80136, n80137, n80138,
         n80139, n80140, n80141, n80142, n80143, n80144, n80145, n80146,
         n80147, n80148, n80149, n80150, n80151, n80152, n80153, n80154,
         n80155, n80156, n80157, n80158, n80159, n80160, n80161, n80162,
         n80163, n80164, n80165, n80166, n80167, n80168, n80169, n80170,
         n80171, n80172, n80173, n80174, n80175, n80176, n80177, n80178,
         n80179, n80180, n80181, n80182, n80183, n80184, n80185, n80186,
         n80187, n80188, n80189, n80190, n80191, n80192, n80193, n80194,
         n80195, n80196, n80197, n80198, n80199, n80200, n80201, n80202,
         n80203, n80204, n80205, n80206, n80207, n80208, n80209, n80210,
         n80211, n80212, n80213, n80214, n80215, n80216, n80217, n80218,
         n80219, n80220, n80221, n80222, n80223, n80224, n80225, n80226,
         n80227, n80228, n80229, n80230, n80231, n80232, n80233, n80234,
         n80235, n80236, n80237, n80238, n80239, n80240, n80241, n80242,
         n80243, n80244, n80245, n80246, n80247, n80248, n80249, n80250,
         n80251, n80252, n80253, n80254, n80255, n80256, n80257, n80258,
         n80259, n80260, n80261, n80262, n80263, n80264, n80265, n80266,
         n80267, n80268, n80269, n80270, n80271, n80272, n80273, n80274,
         n80275, n80276, n80277, n80278, n80279, n80280, n80281, n80282,
         n80283, n80284, n80285, n80286, n80287, n80288, n80289, n80290,
         n80291, n80292, n80293, n80294, n80295, n80296, n80297, n80298,
         n80299, n80300, n80301, n80302, n80303, n80304, n80305, n80306,
         n80307, n80308, n80309, n80310, n80311, n80312, n80313, n80314,
         n80315, n80316, n80317, n80318, n80319, n80320, n80321, n80322,
         n80323, n80324, n80325, n80326, n80327, n80328, n80329, n80330,
         n80331, n80332, n80333, n80334, n80335, n80336, n80337, n80338,
         n80339, n80340, n80341, n80342, n80343, n80344, n80345, n80346,
         n80347, n80348, n80349, n80350, n80351, n80352, n80353, n80354,
         n80355, n80356, n80357, n80358, n80359, n80360, n80361, n80362,
         n80363, n80364, n80365, n80366, n80367, n80368, n80369, n80370,
         n80371, n80372, n80373, n80374, n80375, n80376, n80377, n80378,
         n80379, n80380, n80381, n80382, n80383, n80384, n80385, n80386,
         n80387, n80388, n80389, n80390, n80391, n80392, n80393, n80394,
         n80395, n80396, n80397, n80398, n80399, n80400, n80401, n80402,
         n80403, n80404, n80405, n80406, n80407, n80408, n80409, n80410,
         n80411, n80412, n80413, n80414, n80415, n80416, n80417, n80418,
         n80419, n80420, n80421, n80422, n80423, n80424, n80425, n80426,
         n80427, n80428, n80429, n80430, n80431, n80432, n80433, n80434,
         n80435, n80436, n80437, n80438, n80439, n80440, n80441, n80442,
         n80443, n80444, n80445, n80446, n80447, n80448, n80449, n80450,
         n80451, n80452, n80453, n80454, n80455, n80456, n80457, n80458,
         n80459, n80460, n80461, n80462, n80463, n80464, n80465, n80466,
         n80467, n80468, n80469, n80470, n80471, n80472, n80473, n80474,
         n80475, n80476, n80477, n80478, n80479, n80480, n80481, n80482,
         n80483, n80484, n80485, n80486, n80487, n80488, n80489, n80490,
         n80491, n80492, n80493, n80494, n80495, n80496, n80497, n80498,
         n80499, n80500, n80501, n80502, n80503, n80504, n80505, n80506,
         n80507, n80508, n80509, n80510, n80511, n80512, n80513, n80514,
         n80515, n80516, n80517, n80518, n80519, n80520, n80521, n80522,
         n80523, n80524, n80525, n80526, n80527, n80528, n80529, n80530,
         n80531, n80532, n80533, n80534, n80535, n80536, n80537, n80538,
         n80539, n80540, n80541, n80542, n80543, n80544, n80545, n80546,
         n80547, n80548, n80549, n80550, n80551, n80552, n80553, n80554,
         n80555, n80556, n80557, n80558, n80559, n80560, n80561, n80562,
         n80563, n80564, n80565, n80566, n80567, n80568, n80569, n80570,
         n80571, n80572, n80573, n80574, n80575, n80576, n80577, n80578,
         n80579, n80580, n80581, n80582, n80583, n80584, n80585, n80586,
         n80587, n80588, n80589, n80590, n80591, n80592, n80593, n80594,
         n80595, n80596, n80597, n80598, n80599, n80600, n80601, n80602,
         n80603, n80604, n80605, n80606, n80607, n80608, n80609, n80610,
         n80611, n80612, n80613, n80614, n80615, n80616, n80617, n80618,
         n80619, n80620, n80621, n80622, n80623, n80624, n80625, n80626,
         n80627, n80628, n80629, n80630, n80631, n80632, n80633, n80634,
         n80635, n80636, n80637, n80638, n80639, n80640, n80641, n80642,
         n80643, n80644, n80645, n80646, n80647, n80648, n80649, n80650,
         n80651, n80652, n80653, n80654, n80655, n80656, n80657, n80658,
         n80659, n80660, n80661, n80662, n80663, n80664, n80665, n80666,
         n80667, n80668, n80669, n80670, n80671, n80672, n80673, n80674,
         n80675, n80676, n80677, n80678, n80679, n80680, n80681, n80682,
         n80683, n80684, n80685, n80686, n80687, n80688, n80689, n80690,
         n80691, n80692, n80693, n80694, n80695, n80696, n80697, n80698,
         n80699, n80700, n80701, n80702, n80703, n80704, n80705, n80706,
         n80707, n80708, n80709, n80710, n80711, n80712, n80713, n80714,
         n80715, n80716, n80717, n80718, n80719, n80720, n80721, n80722,
         n80723, n80724, n80725, n80726, n80727, n80728, n80729, n80730,
         n80731, n80732, n80733, n80734, n80735, n80736, n80737, n80738,
         n80739, n80740, n80741, n80742, n80743, n80744, n80745, n80746,
         n80747, n80748, n80749, n80750, n80751, n80752, n80753, n80754,
         n80755, n80756, n80757, n80758, n80759, n80760, n80761, n80762,
         n80763, n80764, n80765, n80766, n80767, n80768, n80769, n80770,
         n80771, n80772, n80773, n80774, n80775, n80776, n80777, n80778,
         n80779, n80780, n80781, n80782, n80783, n80784, n80785, n80786,
         n80787, n80788, n80789, n80790, n80791, n80792, n80793, n80794,
         n80795, n80796, n80797, n80798, n80799, n80800, n80801, n80802,
         n80803, n80804, n80805, n80806, n80807, n80808, n80809, n80810,
         n80811, n80812, n80813, n80814, n80815, n80816, n80817, n80818,
         n80819, n80820, n80821, n80822, n80823, n80824, n80825, n80826,
         n80827, n80828, n80829, n80830, n80831, n80832, n80833, n80834,
         n80835, n80836, n80837, n80838, n80839, n80840, n80841, n80842,
         n80843, n80844, n80845, n80846, n80847, n80848, n80849, n80850,
         n80851, n80852, n80853, n80854, n80855, n80856, n80857, n80858,
         n80859, n80860, n80861, n80862, n80863, n80864, n80865, n80866,
         n80867, n80868, n80869, n80870, n80871, n80872, n80873, n80874,
         n80875, n80876, n80877, n80878, n80879, n80880, n80881, n80882,
         n80883, n80884, n80885, n80886, n80887, n80888, n80889, n80890,
         n80891, n80892, n80893, n80894, n80895, n80896, n80897, n80898,
         n80899, n80900, n80901, n80902, n80903, n80904, n80905, n80906,
         n80907, n80908, n80909, n80910, n80911, n80912, n80913, n80914,
         n80915, n80916, n80917, n80918, n80919, n80920, n80921, n80922,
         n80923, n80924, n80925, n80926, n80927, n80928, n80929, n80930,
         n80931, n80932, n80933, n80934, n80935, n80936, n80937, n80938,
         n80939, n80940, n80941, n80942, n80943, n80944, n80945, n80946,
         n80947, n80948, n80949, n80950, n80951, n80952, n80953, n80954,
         n80955, n80956, n80957, n80958, n80959, n80960, n80961, n80962,
         n80963, n80964, n80965, n80966, n80967, n80968, n80969, n80970,
         n80971, n80972, n80973, n80974, n80975, n80976, n80977, n80978,
         n80979, n80980, n80981, n80982, n80983, n80984, n80985, n80986,
         n80987, n80988, n80989, n80990, n80991, n80992, n80993, n80994,
         n80995, n80996, n80997, n80998, n80999, n81000, n81001, n81002,
         n81003, n81004, n81005, n81006, n81007, n81008, n81009, n81010,
         n81011, n81012, n81013, n81014, n81015, n81016, n81017, n81018,
         n81019, n81020, n81021, n81022, n81023, n81024, n81025, n81026,
         n81027, n81028, n81029, n81030, n81031, n81032, n81033, n81034,
         n81035, n81036, n81037, n81038, n81039, n81040, n81041, n81042,
         n81043, n81044, n81045, n81046, n81047, n81048, n81049, n81050,
         n81051, n81052, n81053, n81054, n81055, n81056, n81057, n81058,
         n81059, n81060, n81061, n81062, n81063, n81064, n81065, n81066,
         n81067, n81068, n81069, n81070, n81071, n81072, n81073, n81074,
         n81075, n81076, n81077, n81078, n81079, n81080, n81081, n81082,
         n81083, n81084, n81085, n81086, n81087, n81088, n81089, n81090,
         n81091, n81092, n81093, n81094, n81095, n81096, n81097, n81098,
         n81099, n81100, n81101, n81102, n81103, n81104, n81105, n81106,
         n81107, n81108, n81109, n81110, n81111, n81112, n81113, n81114,
         n81115, n81116, n81117, n81118, n81119, n81120, n81121, n81122,
         n81123, n81124, n81125, n81126, n81127, n81128, n81129, n81130,
         n81131, n81132, n81133, n81134, n81135, n81136, n81137, n81138,
         n81139, n81140, n81141, n81142, n81143, n81144, n81145, n81146,
         n81147, n81148, n81149, n81150, n81151, n81152, n81153, n81154,
         n81155, n81156, n81157, n81158, n81159, n81160, n81161, n81162,
         n81163, n81164, n81165, n81166, n81167, n81168, n81169, n81170,
         n81171, n81172, n81173, n81174, n81175, n81176, n81177, n81178,
         n81179, n81180, n81181, n81182, n81183, n81184, n81185, n81186,
         n81187, n81188, n81189, n81190, n81191, n81192, n81193, n81194,
         n81195, n81196, n81197, n81198, n81199, n81200, n81201, n81202,
         n81203, n81204, n81205, n81206, n81207, n81208, n81209, n81210,
         n81211, n81212, n81213, n81214, n81215, n81216, n81217, n81218,
         n81219, n81220, n81221, n81222, n81223, n81224, n81225, n81226,
         n81227, n81228, n81229, n81230, n81231, n81232, n81233, n81234,
         n81235, n81236, n81237, n81238, n81239, n81240, n81241, n81242,
         n81243, n81244, n81245, n81246, n81247, n81248, n81249, n81250,
         n81251, n81252, n81253, n81254, n81255, n81256, n81257, n81258,
         n81259, n81260, n81261, n81262, n81263, n81264, n81265, n81266,
         n81267, n81268, n81269, n81270, n81271, n81272, n81273, n81274,
         n81275, n81276, n81277, n81278, n81279, n81280, n81281, n81282,
         n81283, n81284, n81285, n81286, n81287, n81288, n81289, n81290,
         n81291, n81292, n81293, n81294, n81295, n81296, n81297, n81298,
         n81299, n81300, n81301, n81302, n81303, n81304, n81305, n81306,
         n81307, n81308, n81309, n81310, n81311, n81312, n81313, n81314,
         n81315, n81316, n81317, n81318, n81319, n81320, n81321, n81322,
         n81323, n81324, n81325, n81326, n81327, n81328, n81329, n81330,
         n81331, n81332, n81333, n81334, n81335, n81336, n81337, n81338,
         n81339, n81340, n81341, n81342, n81343, n81344, n81345, n81346,
         n81347, n81348, n81349, n81350, n81351, n81352, n81353, n81354,
         n81355, n81356, n81357, n81358, n81359, n81360, n81361, n81362,
         n81363, n81364, n81365, n81366, n81367, n81368, n81369, n81370,
         n81371, n81372, n81373, n81374, n81375, n81376, n81377, n81378,
         n81379, n81380, n81381, n81382, n81383, n81384, n81385, n81386,
         n81387, n81388, n81389, n81390, n81391, n81392, n81393, n81394,
         n81395, n81396, n81397, n81398, n81399, n81400, n81401, n81402,
         n81403, n81404, n81405, n81406, n81407, n81408, n81409, n81410,
         n81411, n81412, n81413, n81414, n81415, n81416, n81417, n81418,
         n81419, n81420, n81421, n81422, n81423, n81424, n81425, n81426,
         n81427, n81428, n81429, n81430, n81431, n81432, n81433, n81434,
         n81435, n81436, n81437, n81438, n81439, n81440, n81441, n81442,
         n81443, n81444, n81445, n81446, n81447, n81448, n81449, n81450,
         n81451, n81452, n81453, n81454, n81455, n81456, n81457, n81458,
         n81459, n81460, n81461, n81462, n81463, n81464, n81465, n81466,
         n81467, n81468, n81469, n81470, n81471, n81472, n81473, n81474,
         n81475, n81476, n81477, n81478, n81479, n81480, n81481, n81482,
         n81483, n81484, n81485, n81486, n81487, n81488, n81489, n81490,
         n81491, n81492, n81493, n81494, n81495, n81496, n81497, n81498,
         n81499, n81500, n81501, n81502, n81503, n81504, n81505, n81506,
         n81507, n81508, n81509, n81510, n81511, n81512, n81513, n81514,
         n81515, n81516, n81517, n81518, n81519, n81520, n81521, n81522,
         n81523, n81524, n81525, n81526, n81527, n81528, n81529, n81530,
         n81531, n81532, n81533, n81534, n81535, n81536, n81537, n81538,
         n81539, n81540, n81541, n81542, n81543, n81544, n81545, n81546,
         n81547, n81548, n81549, n81550, n81551, n81552, n81553, n81554,
         n81555, n81556, n81557, n81558, n81559, n81560, n81561, n81562,
         n81563, n81564, n81565, n81566, n81567, n81568, n81569, n81570,
         n81571, n81572, n81573, n81574, n81575, n81576, n81577, n81578,
         n81579, n81580, n81581, n81582, n81583, n81584, n81585, n81586,
         n81587, n81588, n81589, n81590, n81591, n81592, n81593, n81594,
         n81595, n81596, n81597, n81598, n81599, n81600, n81601, n81602,
         n81603, n81604, n81605, n81606, n81607, n81608, n81609, n81610,
         n81611, n81612, n81613, n81614, n81615, n81616, n81617, n81618,
         n81619, n81620, n81621, n81622, n81623, n81624, n81625, n81626,
         n81627, n81628, n81629, n81630, n81631, n81632, n81633, n81634,
         n81635, n81636, n81637, n81638, n81639, n81640, n81641, n81642,
         n81643, n81644, n81645, n81646, n81647, n81648, n81649, n81650,
         n81651, n81652, n81653, n81654, n81655, n81656, n81657, n81658,
         n81659, n81660, n81661, n81662, n81663, n81664, n81665, n81666,
         n81667, n81668, n81669, n81670, n81671, n81672, n81673, n81674,
         n81675, n81676, n81677, n81678, n81679, n81680, n81681, n81682,
         n81683, n81684, n81685, n81686, n81687, n81688, n81689, n81690,
         n81691, n81692, n81693, n81694, n81695, n81696, n81697, n81698,
         n81699, n81700, n81701, n81702, n81703, n81704, n81705, n81706,
         n81707, n81708, n81709, n81710, n81711, n81712, n81713, n81714,
         n81715, n81716, n81717, n81718, n81719, n81720, n81721, n81722,
         n81723, n81724, n81725, n81726, n81727, n81728, n81729, n81730,
         n81731, n81732, n81733, n81734, n81735, n81736, n81737, n81738,
         n81739, n81740, n81741, n81742, n81743, n81744, n81745, n81746,
         n81747, n81748, n81749, n81750, n81751, n81752, n81753, n81754,
         n81755, n81756, n81757, n81758, n81759, n81760, n81761, n81762,
         n81763, n81764, n81765, n81766, n81767, n81768, n81769, n81770,
         n81771, n81772, n81773, n81774, n81775, n81776, n81777, n81778,
         n81779, n81780, n81781, n81782, n81783, n81784, n81785, n81786,
         n81787, n81788, n81789, n81790, n81791, n81792, n81793, n81794,
         n81795, n81796, n81797, n81798, n81799, n81800, n81801, n81802,
         n81803, n81804, n81805, n81806, n81807, n81808, n81809, n81810,
         n81811, n81812, n81813, n81814, n81815, n81816, n81817, n81818,
         n81819, n81820, n81821, n81822, n81823, n81824, n81825, n81826,
         n81827, n81828, n81829, n81830, n81831, n81832, n81833, n81834,
         n81835, n81836, n81837, n81838, n81839, n81840, n81841, n81842,
         n81843, n81844, n81845, n81846, n81847, n81848, n81849, n81850,
         n81851, n81852, n81853, n81854, n81855, n81856, n81857, n81858,
         n81859, n81860, n81861, n81862, n81863, n81864, n81865, n81866,
         n81867, n81868, n81869, n81870, n81871, n81872, n81873, n81874,
         n81875, n81876, n81877, n81878, n81879, n81880, n81881, n81882,
         n81883, n81884, n81885, n81886, n81887, n81888, n81889, n81890,
         n81891, n81892, n81893, n81894, n81895, n81896, n81897, n81898,
         n81899, n81900, n81901, n81902, n81903, n81904, n81905, n81906,
         n81907, n81908, n81909, n81910, n81911, n81912, n81913, n81914,
         n81915, n81916, n81917, n81918, n81919, n81920, n81921, n81922,
         n81923, n81924, n81925, n81926, n81927, n81928, n81929, n81930,
         n81931, n81932, n81933, n81934, n81935, n81936, n81937, n81938,
         n81939, n81940, n81941, n81942, n81943, n81944, n81945, n81946,
         n81947, n81948, n81949, n81950, n81951, n81952, n81953, n81954,
         n81955, n81956, n81957, n81958, n81959, n81960, n81961, n81962,
         n81963, n81964, n81965, n81966, n81967, n81968, n81969, n81970,
         n81971, n81972, n81973, n81974, n81975, n81976, n81977, n81978,
         n81979, n81980, n81981, n81982, n81983, n81984, n81985, n81986,
         n81987, n81988, n81989, n81990, n81991, n81992, n81993, n81994,
         n81995, n81996, n81997, n81998, n81999, n82000, n82001, n82002,
         n82003, n82004, n82005, n82006, n82007, n82008, n82009, n82010,
         n82011, n82012, n82013, n82014, n82015, n82016, n82017, n82018,
         n82019, n82020, n82021, n82022, n82023, n82024, n82025, n82026,
         n82027, n82028, n82029, n82030, n82031, n82032, n82033, n82034,
         n82035, n82036, n82037, n82038, n82039, n82040, n82041, n82042,
         n82043, n82044, n82045, n82046, n82047, n82048, n82049, n82050,
         n82051, n82052, n82053, n82054, n82055, n82056, n82057, n82058,
         n82059, n82060, n82061, n82062, n82063, n82064, n82065, n82066,
         n82067, n82068, n82069, n82070, n82071, n82072, n82073, n82074,
         n82075, n82076, n82077, n82078, n82079, n82080, n82081, n82082,
         n82083, n82084, n82085, n82086, n82087, n82088, n82089, n82090,
         n82091, n82092, n82093, n82094, n82095, n82096, n82097, n82098,
         n82099, n82100, n82101, n82102, n82103, n82104, n82105, n82106,
         n82107, n82108, n82109, n82110, n82111, n82112, n82113, n82114,
         n82115, n82116, n82117, n82118, n82119, n82120, n82121, n82122,
         n82123, n82124, n82125, n82126, n82127, n82128, n82129, n82130,
         n82131, n82132, n82133, n82134, n82135, n82136, n82137, n82138,
         n82139, n82140, n82141, n82142, n82143, n82144, n82145, n82146,
         n82147, n82148, n82149, n82150, n82151, n82152, n82153, n82154,
         n82155, n82156, n82157, n82158, n82159, n82160, n82161, n82162,
         n82163, n82164, n82165, n82166, n82167, n82168, n82169, n82170,
         n82171, n82172, n82173, n82174, n82175, n82176, n82177, n82178,
         n82179, n82180, n82181, n82182, n82183, n82184, n82185, n82186,
         n82187, n82188, n82189, n82190, n82191, n82192, n82193, n82194,
         n82195, n82196, n82197, n82198, n82199, n82200, n82201, n82202,
         n82203, n82204, n82205, n82206, n82207, n82208, n82209, n82210,
         n82211, n82212, n82213, n82214, n82215, n82216, n82217, n82218,
         n82219, n82220, n82221, n82222, n82223, n82224, n82225, n82226,
         n82227, n82228, n82229, n82230, n82231, n82232, n82233, n82234,
         n82235, n82236, n82237, n82238, n82239, n82240, n82241, n82242,
         n82243, n82244, n82245, n82246, n82247, n82248, n82249, n82250,
         n82251, n82252, n82253, n82254, n82255, n82256, n82257, n82258,
         n82259, n82260, n82261, n82262, n82263, n82264, n82265, n82266,
         n82267, n82268, n82269, n82270, n82271, n82272, n82273, n82274,
         n82275, n82276, n82277, n82278, n82279, n82280, n82281, n82282,
         n82283, n82284, n82285, n82286, n82287, n82288, n82289, n82290,
         n82291, n82292, n82293, n82294, n82295, n82296, n82297, n82298,
         n82299, n82300, n82301, n82302, n82303, n82304, n82305, n82306,
         n82307, n82308, n82309, n82310, n82311, n82312, n82313, n82314,
         n82315, n82316, n82317, n82318, n82319, n82320, n82321, n82322,
         n82323, n82324, n82325, n82326, n82327, n82328, n82329, n82330,
         n82331, n82332, n82333, n82334, n82335, n82336, n82337, n82338,
         n82339, n82340, n82341, n82342, n82343, n82344, n82345, n82346,
         n82347, n82348, n82349, n82350, n82351, n82352, n82353, n82354,
         n82355, n82356, n82357, n82358, n82359, n82360, n82361, n82362,
         n82363, n82364, n82365, n82366, n82367, n82368, n82369, n82370,
         n82371, n82372, n82373, n82374, n82375, n82376, n82377, n82378,
         n82379, n82380, n82381, n82382, n82383, n82384, n82385, n82386,
         n82387, n82388, n82389, n82390, n82391, n82392, n82393, n82394,
         n82395, n82396, n82397, n82398, n82399, n82400, n82401, n82402,
         n82403, n82404, n82405, n82406, n82407, n82408, n82409, n82410,
         n82411, n82412, n82413, n82414, n82415, n82416, n82417, n82418,
         n82419, n82420, n82421, n82422, n82423, n82424, n82425, n82426,
         n82427, n82428, n82429, n82430, n82431, n82432, n82433, n82434,
         n82435, n82436, n82437, n82438, n82439, n82440, n82441, n82442,
         n82443, n82444, n82445, n82446, n82447, n82448, n82449, n82450,
         n82451, n82452, n82453, n82454, n82455, n82456, n82457, n82458,
         n82459, n82460, n82461, n82462, n82463, n82464, n82465, n82466,
         n82467, n82468, n82469, n82470, n82471, n82472, n82473, n82474,
         n82475, n82476, n82477, n82478, n82479, n82480, n82481, n82482,
         n82483, n82484, n82485, n82486, n82487, n82488, n82489, n82490,
         n82491, n82492, n82493, n82494, n82495, n82496, n82497, n82498,
         n82499, n82500, n82501, n82502, n82503, n82504, n82505, n82506,
         n82507, n82508, n82509, n82510, n82511, n82512, n82513, n82514,
         n82515, n82516, n82517, n82518, n82519, n82520, n82521, n82522,
         n82523, n82524, n82525, n82526, n82527, n82528, n82529, n82530,
         n82531, n82532, n82533, n82534, n82535, n82536, n82537, n82538,
         n82539, n82540, n82541, n82542, n82543, n82544, n82545, n82546,
         n82547, n82548, n82549, n82550, n82551, n82552, n82553, n82554,
         n82555, n82556, n82557, n82558, n82559, n82560, n82561, n82562,
         n82563, n82564, n82565, n82566, n82567, n82568, n82569, n82570,
         n82571, n82572, n82573, n82574, n82575, n82576, n82577, n82578,
         n82579, n82580, n82581, n82582, n82583, n82584, n82585, n82586,
         n82587, n82588, n82589, n82590, n82591, n82592, n82593, n82594,
         n82595, n82596, n82597, n82598, n82599, n82600, n82601, n82602,
         n82603, n82604, n82605, n82606, n82607, n82608, n82609, n82610,
         n82611, n82612, n82613, n82614, n82615, n82616, n82617, n82618,
         n82619, n82620, n82621, n82622, n82623, n82624, n82625, n82626,
         n82627, n82628, n82629, n82630, n82631, n82632, n82633, n82634,
         n82635, n82636, n82637, n82638, n82639, n82640, n82641, n82642,
         n82643, n82644, n82645, n82646, n82647, n82648, n82649, n82650,
         n82651, n82652, n82653, n82654, n82655, n82656, n82657, n82658,
         n82659, n82660, n82661, n82662, n82663, n82664, n82665, n82666,
         n82667, n82668, n82669, n82670, n82671, n82672, n82673, n82674,
         n82675, n82676, n82677, n82678, n82679, n82680, n82681, n82682,
         n82683, n82684, n82685, n82686, n82687, n82688, n82689, n82690,
         n82691, n82692, n82693, n82694, n82695, n82696, n82697, n82698,
         n82699, n82700, n82701, n82702, n82703, n82704, n82705, n82706,
         n82707, n82708, n82709, n82710, n82711, n82712, n82713, n82714,
         n82715, n82716, n82717, n82718, n82719, n82720, n82721, n82722,
         n82723, n82724, n82725, n82726, n82727, n82728, n82729, n82730,
         n82731, n82732, n82733, n82734, n82735, n82736, n82737, n82738,
         n82739, n82740, n82741, n82742, n82743, n82744, n82745, n82746,
         n82747, n82748, n82749, n82750, n82751, n82752, n82753, n82754,
         n82755, n82756, n82757, n82758, n82759, n82760, n82761, n82762,
         n82763, n82764, n82765, n82766, n82767, n82768, n82769, n82770,
         n82771, n82772, n82773, n82774, n82775, n82776, n82777, n82778,
         n82779, n82780, n82781, n82782, n82783, n82784, n82785, n82786,
         n82787, n82788, n82789, n82790, n82791, n82792, n82793, n82794,
         n82795, n82796, n82797, n82798, n82799, n82800, n82801, n82802,
         n82803, n82804, n82805, n82806, n82807, n82808, n82809, n82810,
         n82811, n82812, n82813, n82814, n82815, n82816, n82817, n82818,
         n82819, n82820, n82821, n82822, n82823, n82824, n82825, n82826,
         n82827, n82828, n82829, n82830, n82831, n82832, n82833, n82834,
         n82835, n82836, n82837, n82838, n82839, n82840, n82841, n82842,
         n82843, n82844, n82845, n82846, n82847, n82848, n82849, n82850,
         n82851, n82852, n82853, n82854, n82855, n82856, n82857, n82858,
         n82859, n82860, n82861, n82862, n82863, n82864, n82865, n82866,
         n82867, n82868, n82869, n82870, n82871, n82872, n82873, n82874,
         n82875, n82876, n82877, n82878, n82879, n82880, n82881, n82882,
         n82883, n82884, n82885, n82886, n82887, n82888, n82889, n82890,
         n82891, n82892, n82893, n82894, n82895, n82896, n82897, n82898,
         n82899, n82900, n82901, n82902, n82903, n82904, n82905, n82906,
         n82907, n82908, n82909, n82910, n82911, n82912, n82913, n82914,
         n82915, n82916, n82917, n82918, n82919, n82920, n82921, n82922,
         n82923, n82924, n82925, n82926, n82927, n82928, n82929, n82930,
         n82931, n82932, n82933, n82934, n82935, n82936, n82937, n82938,
         n82939, n82940, n82941, n82942, n82943, n82944, n82945, n82946,
         n82947, n82948, n82949, n82950, n82951, n82952, n82953, n82954,
         n82955, n82956, n82957, n82958, n82959, n82960, n82961, n82962,
         n82963, n82964, n82965, n82966, n82967, n82968, n82969, n82970,
         n82971, n82972, n82973, n82974, n82975, n82976, n82977, n82978,
         n82979, n82980, n82981, n82982, n82983, n82984, n82985, n82986,
         n82987, n82988, n82989, n82990, n82991, n82992, n82993, n82994,
         n82995, n82996, n82997, n82998, n82999, n83000, n83001, n83002,
         n83003, n83004, n83005, n83006, n83007, n83008, n83009, n83010,
         n83011, n83012, n83013, n83014, n83015, n83016, n83017, n83018,
         n83019, n83020, n83021, n83022, n83023, n83024, n83025, n83026,
         n83027, n83028, n83029, n83030, n83031, n83032, n83033, n83034,
         n83035, n83036, n83037, n83038, n83039, n83040, n83041, n83042,
         n83043, n83044, n83045, n83046, n83047, n83048, n83049, n83050,
         n83051, n83052, n83053, n83054, n83055, n83056, n83057, n83058,
         n83059, n83060, n83061, n83062, n83063, n83064, n83065, n83066,
         n83067, n83068, n83069, n83070, n83071, n83072, n83073, n83074,
         n83075, n83076, n83077, n83078, n83079, n83080, n83081, n83082,
         n83083, n83084, n83085, n83086, n83087, n83088, n83089, n83090,
         n83091, n83092, n83093, n83094, n83095, n83096, n83097, n83098,
         n83099, n83100, n83101, n83102, n83103, n83104, n83105, n83106,
         n83107, n83108, n83109, n83110, n83111, n83112, n83113, n83114,
         n83115, n83116, n83117, n83118, n83119, n83120, n83121, n83122,
         n83123, n83124, n83125, n83126, n83127, n83128, n83129, n83130,
         n83131, n83132, n83133, n83134, n83135, n83136, n83137, n83138,
         n83139, n83140, n83141, n83142, n83143, n83144, n83145, n83146,
         n83147, n83148, n83149, n83150, n83151, n83152, n83153, n83154,
         n83155, n83156, n83157, n83158, n83159, n83160, n83161, n83162,
         n83163, n83164, n83165, n83166, n83167, n83168, n83169, n83170,
         n83171, n83172, n83173, n83174, n83175, n83176, n83177, n83178,
         n83179, n83180, n83181, n83182, n83183, n83184, n83185, n83186,
         n83187, n83188, n83189, n83190, n83191, n83192, n83193, n83194,
         n83195, n83196, n83197, n83198, n83199, n83200, n83201, n83202,
         n83203, n83204, n83205, n83206, n83207, n83208, n83209, n83210,
         n83211, n83212, n83213, n83214, n83215, n83216, n83217, n83218,
         n83219, n83220, n83221, n83222, n83223, n83224, n83225, n83226,
         n83227, n83228, n83229, n83230, n83231, n83232, n83233, n83234,
         n83235, n83236, n83237, n83238, n83239, n83240, n83241, n83242,
         n83243, n83244, n83245, n83246, n83247, n83248, n83249, n83250,
         n83251, n83252, n83253, n83254, n83255, n83256, n83257, n83258,
         n83259, n83260, n83261, n83262, n83263, n83264, n83265, n83266,
         n83267, n83268, n83269, n83270, n83271, n83272, n83273, n83274,
         n83275, n83276, n83277, n83278, n83279, n83280, n83281, n83282,
         n83283, n83284, n83285, n83286, n83287, n83288, n83289, n83290,
         n83291, n83292, n83293, n83294, n83295, n83296, n83297, n83298,
         n83299, n83300, n83301, n83302, n83303, n83304, n83305, n83306,
         n83307, n83308, n83309, n83310, n83311, n83312, n83313, n83314,
         n83315, n83316, n83317, n83318, n83319, n83320, n83321, n83322,
         n83323, n83324, n83325, n83326, n83327, n83328, n83329, n83330,
         n83331, n83332, n83333, n83334, n83335, n83336, n83337, n83338,
         n83339, n83340, n83341, n83342, n83343, n83344, n83345, n83346,
         n83347, n83348, n83349, n83350, n83351, n83352, n83353, n83354,
         n83355, n83356, n83357, n83358, n83359, n83360, n83361, n83362,
         n83363, n83364, n83365, n83366, n83367, n83368, n83369, n83370,
         n83371, n83372, n83373, n83374, n83375, n83376, n83377, n83378,
         n83379, n83380, n83381, n83382, n83383, n83384, n83385, n83386,
         n83387, n83388, n83389, n83390, n83391, n83392, n83393, n83394,
         n83395, n83396, n83397, n83398, n83399, n83400, n83401, n83402,
         n83403, n83404, n83405, n83406, n83407, n83408, n83409, n83410,
         n83411, n83412, n83413, n83414, n83415, n83416, n83417, n83418,
         n83419, n83420, n83421, n83422, n83423, n83424, n83425, n83426,
         n83427, n83428, n83429, n83430, n83431, n83432, n83433, n83434,
         n83435, n83436, n83437, n83438, n83439, n83440, n83441, n83442,
         n83443, n83444, n83445, n83446, n83447, n83448, n83449, n83450,
         n83451, n83452, n83453, n83454, n83455, n83456, n83457, n83458,
         n83459, n83460, n83461, n83462, n83463, n83464, n83465, n83466,
         n83467, n83468, n83469, n83470, n83471, n83472, n83473, n83474,
         n83475, n83476, n83477, n83478, n83479, n83480, n83481, n83482,
         n83483, n83484, n83485, n83486, n83487, n83488, n83489, n83490,
         n83491, n83492, n83493, n83494, n83495, n83496, n83497, n83498,
         n83499, n83500, n83501, n83502, n83503, n83504, n83505, n83506,
         n83507, n83508, n83509, n83510, n83511, n83512, n83513, n83514,
         n83515, n83516, n83517, n83518, n83519, n83520, n83521, n83522,
         n83523, n83524, n83525, n83526, n83527, n83528, n83529, n83530,
         n83531, n83532, n83533, n83534, n83535, n83536, n83537, n83538,
         n83539, n83540, n83541, n83542, n83543, n83544, n83545, n83546,
         n83547, n83548, n83549, n83550, n83551, n83552, n83553, n83554,
         n83555, n83556, n83557, n83558, n83559, n83560, n83561, n83562,
         n83563, n83564, n83565, n83566, n83567, n83568, n83569, n83570,
         n83571, n83572, n83573, n83574, n83575, n83576, n83577, n83578,
         n83579, n83580, n83581, n83582, n83583, n83584, n83585, n83586,
         n83587, n83588, n83589, n83590, n83591, n83592, n83593, n83594,
         n83595, n83596, n83597, n83598, n83599, n83600, n83601, n83602,
         n83603, n83604, n83605, n83606, n83607, n83608, n83609, n83610,
         n83611, n83612, n83613, n83614, n83615, n83616, n83617, n83618,
         n83619, n83620, n83621, n83622, n83623, n83624, n83625, n83626,
         n83627, n83628, n83629, n83630, n83631, n83632, n83633, n83634,
         n83635, n83636, n83637, n83638, n83639, n83640, n83641, n83642,
         n83643, n83644, n83645, n83646, n83647, n83648, n83649, n83650,
         n83651, n83652, n83653, n83654, n83655, n83656, n83657, n83658,
         n83659, n83660, n83661, n83662, n83663, n83664, n83665, n83666,
         n83667, n83668, n83669, n83670, n83671, n83672, n83673, n83674,
         n83675, n83676, n83677, n83678, n83679, n83680, n83681, n83682,
         n83683, n83684, n83685, n83686, n83687, n83688, n83689, n83690,
         n83691, n83692, n83693, n83694, n83695, n83696, n83697, n83698,
         n83699, n83700, n83701, n83702, n83703, n83704, n83705, n83706,
         n83707, n83708, n83709, n83710, n83711, n83712, n83713, n83714,
         n83715, n83716, n83717, n83718, n83719, n83720, n83721, n83722,
         n83723, n83724, n83725, n83726, n83727, n83728, n83729, n83730,
         n83731, n83732, n83733, n83734, n83735, n83736, n83737, n83738,
         n83739, n83740, n83741, n83742, n83743, n83744, n83745, n83746,
         n83747, n83748, n83749, n83750, n83751, n83752, n83753, n83754,
         n83755, n83756, n83757, n83758, n83759, n83760, n83761, n83762,
         n83763, n83764, n83765, n83766, n83767, n83768, n83769, n83770,
         n83771, n83772, n83773, n83774, n83775, n83776, n83777, n83778,
         n83779, n83780, n83781, n83782, n83783, n83784, n83785, n83786,
         n83787, n83788, n83789, n83790, n83791, n83792, n83793, n83794,
         n83795, n83796, n83797, n83798, n83799, n83800, n83801, n83802,
         n83803, n83804, n83805, n83806, n83807, n83808, n83809, n83810,
         n83811, n83812, n83813, n83814, n83815, n83816, n83817, n83818,
         n83819, n83820, n83821, n83822, n83823, n83824, n83825, n83826,
         n83827, n83828, n83829, n83830, n83831, n83832, n83833, n83834,
         n83835, n83836, n83837, n83838, n83839, n83840, n83841, n83842,
         n83843, n83844, n83845, n83846, n83847, n83848, n83849, n83850,
         n83851, n83852, n83853, n83854, n83855, n83856, n83857, n83858,
         n83859, n83860, n83861, n83862, n83863, n83864, n83865, n83866,
         n83867, n83868, n83869, n83870, n83871, n83872, n83873, n83874,
         n83875, n83876, n83877, n83878, n83879, n83880, n83881, n83882,
         n83883, n83884, n83885, n83886, n83887, n83888, n83889, n83890,
         n83891, n83892, n83893, n83894, n83895, n83896, n83897, n83898,
         n83899, n83900, n83901, n83902, n83903, n83904, n83905, n83906,
         n83907, n83908, n83909, n83910, n83911, n83912, n83913, n83914,
         n83915, n83916, n83917, n83918, n83919, n83920, n83921, n83922,
         n83923, n83924, n83925, n83926, n83927, n83928, n83929, n83930,
         n83931, n83932, n83933, n83934, n83935, n83936, n83937, n83938,
         n83939, n83940, n83941, n83942, n83943, n83944, n83945, n83946,
         n83947, n83948, n83949, n83950, n83951, n83952, n83953, n83954,
         n83955, n83956, n83957, n83958, n83959, n83960, n83961, n83962,
         n83963, n83964, n83965, n83966, n83967, n83968, n83969, n83970,
         n83971, n83972, n83973, n83974, n83975, n83976, n83977, n83978,
         n83979, n83980, n83981, n83982, n83983, n83984, n83985, n83986,
         n83987, n83988, n83989, n83990, n83991, n83992, n83993, n83994,
         n83995, n83996, n83997, n83998, n83999, n84000, n84001, n84002,
         n84003, n84004, n84005, n84006, n84007, n84008, n84009, n84010,
         n84011, n84012, n84013, n84014, n84015, n84016, n84017, n84018,
         n84019, n84020, n84021, n84022, n84023, n84024, n84025, n84026,
         n84027, n84028, n84029, n84030, n84031, n84032, n84033, n84034,
         n84035, n84036, n84037, n84038, n84039, n84040, n84041, n84042,
         n84043, n84044, n84045, n84046, n84047, n84048, n84049, n84050,
         n84051, n84052, n84053, n84054, n84055, n84056, n84057, n84058,
         n84059, n84060, n84061, n84062, n84063, n84064, n84065, n84066,
         n84067, n84068, n84069, n84070, n84071, n84072, n84073, n84074,
         n84075, n84076, n84077, n84078, n84079, n84080, n84081, n84082,
         n84083, n84084, n84085, n84086, n84087, n84088, n84089, n84090,
         n84091, n84092, n84093, n84094, n84095, n84096, n84097, n84098,
         n84099, n84100, n84101, n84102, n84103, n84104, n84105, n84106,
         n84107, n84108, n84109, n84110, n84111, n84112, n84113, n84114,
         n84115, n84116, n84117, n84118, n84119, n84120, n84121, n84122,
         n84123, n84124, n84125, n84126, n84127, n84128, n84129, n84130,
         n84131, n84132, n84133, n84134, n84135, n84136, n84137, n84138,
         n84139, n84140, n84141, n84142, n84143, n84144, n84145, n84146,
         n84147, n84148, n84149, n84150, n84151, n84152, n84153, n84154,
         n84155, n84156, n84157, n84158, n84159, n84160, n84161, n84162,
         n84163, n84164, n84165, n84166, n84167, n84168, n84169, n84170,
         n84171, n84172, n84173, n84174, n84175, n84176, n84177, n84178,
         n84179, n84180, n84181, n84182, n84183, n84184, n84185, n84186,
         n84187, n84188, n84189, n84190, n84191, n84192, n84193, n84194,
         n84195, n84196, n84197, n84198, n84199, n84200, n84201, n84202,
         n84203, n84204, n84205, n84206, n84207, n84208, n84209, n84210,
         n84211, n84212, n84213, n84214, n84215, n84216, n84217, n84218,
         n84219, n84220, n84221, n84222, n84223, n84224, n84225, n84226,
         n84227, n84228, n84229, n84230, n84231, n84232, n84233, n84234,
         n84235, n84236, n84237, n84238, n84239, n84240, n84241, n84242,
         n84243, n84244, n84245, n84246, n84247, n84248, n84249, n84250,
         n84251, n84252, n84253, n84254, n84255, n84256, n84257, n84258,
         n84259, n84260, n84261, n84262, n84263, n84264, n84265, n84266,
         n84267, n84268, n84269, n84270, n84271, n84272, n84273, n84274,
         n84275, n84276, n84277, n84278, n84279, n84280, n84281, n84282,
         n84283, n84284, n84285, n84286, n84287, n84288, n84289, n84290,
         n84291, n84292, n84293, n84294, n84295, n84296, n84297, n84298,
         n84299, n84300, n84301, n84302, n84303, n84304, n84305, n84306,
         n84307, n84308, n84309, n84310, n84311, n84312, n84313, n84314,
         n84315, n84316, n84317, n84318, n84319, n84320, n84321, n84322,
         n84323, n84324, n84325, n84326, n84327, n84328, n84329, n84330,
         n84331, n84332, n84333, n84334, n84335, n84336, n84337, n84338,
         n84339, n84340, n84341, n84342, n84343, n84344, n84345, n84346,
         n84347, n84348, n84349, n84350, n84351, n84352, n84353, n84354,
         n84355, n84356, n84357, n84358, n84359, n84360, n84361, n84362,
         n84363, n84364, n84365, n84366, n84367, n84368, n84369, n84370,
         n84371, n84372, n84373, n84374, n84375, n84376, n84377, n84378,
         n84379, n84380, n84381, n84382, n84383, n84384, n84385, n84386,
         n84387, n84388, n84389, n84390, n84391, n84392, n84393, n84394,
         n84395, n84396, n84397, n84398, n84399, n84400, n84401, n84402,
         n84403, n84404, n84405, n84406, n84407, n84408, n84409, n84410,
         n84411, n84412, n84413, n84414, n84415, n84416, n84417, n84418,
         n84419, n84420, n84421, n84422, n84423, n84424, n84425, n84426,
         n84427, n84428, n84429, n84430, n84431, n84432, n84433, n84434,
         n84435, n84436, n84437, n84438, n84439, n84440, n84441, n84442,
         n84443, n84444, n84445, n84446, n84447, n84448, n84449, n84450,
         n84451, n84452, n84453, n84454, n84455, n84456, n84457, n84458,
         n84459, n84460, n84461, n84462, n84463, n84464, n84465, n84466,
         n84467, n84468, n84469, n84470, n84471, n84472, n84473, n84474,
         n84475, n84476, n84477, n84478, n84479, n84480, n84481, n84482,
         n84483, n84484, n84485, n84486, n84487, n84488, n84489, n84490,
         n84491, n84492, n84493, n84494, n84495, n84496, n84497, n84498,
         n84499, n84500, n84501, n84502, n84503, n84504, n84505, n84506,
         n84507, n84508, n84509, n84510, n84511, n84512, n84513, n84514,
         n84515, n84516, n84517, n84518, n84519, n84520, n84521, n84522,
         n84523, n84524, n84525, n84526, n84527, n84528, n84529, n84530,
         n84531, n84532, n84533, n84534, n84535, n84536, n84537, n84538,
         n84539, n84540, n84541, n84542, n84543, n84544, n84545, n84546,
         n84547, n84548, n84549, n84550, n84551, n84552, n84553, n84554,
         n84555, n84556, n84557, n84558, n84559, n84560, n84561, n84562,
         n84563, n84564, n84565, n84566, n84567, n84568, n84569, n84570,
         n84571, n84572, n84573, n84574, n84575, n84576, n84577, n84578,
         n84579, n84580, n84581, n84582, n84583, n84584, n84585, n84586,
         n84587, n84588, n84589, n84590, n84591, n84592, n84593, n84594,
         n84595, n84596, n84597, n84598, n84599, n84600, n84601, n84602,
         n84603, n84604, n84605, n84606, n84607, n84608, n84609, n84610,
         n84611, n84612, n84613, n84614, n84615, n84616, n84617, n84618,
         n84619, n84620, n84621, n84622, n84623, n84624, n84625, n84626,
         n84627, n84628, n84629, n84630, n84631, n84632, n84633, n84634,
         n84635, n84636, n84637, n84638, n84639, n84640, n84641, n84642,
         n84643, n84644, n84645, n84646, n84647, n84648, n84649, n84650,
         n84651, n84652, n84653, n84654, n84655, n84656, n84657, n84658,
         n84659, n84660, n84661, n84662, n84663, n84664, n84665, n84666,
         n84667, n84668, n84669, n84670, n84671, n84672, n84673, n84674,
         n84675, n84676, n84677, n84678, n84679, n84680, n84681, n84682,
         n84683, n84684, n84685, n84686, n84687, n84688, n84689, n84690,
         n84691, n84692, n84693, n84694, n84695, n84696, n84697, n84698,
         n84699, n84700, n84701, n84702, n84703, n84704, n84705, n84706,
         n84707, n84708, n84709, n84710, n84711, n84712, n84713, n84714,
         n84715, n84716, n84717, n84718, n84719, n84720, n84721, n84722,
         n84723, n84724, n84725, n84726, n84727, n84728, n84729, n84730,
         n84731, n84732, n84733, n84734, n84735, n84736, n84737, n84738,
         n84739, n84740, n84741, n84742, n84743, n84744, n84745, n84746,
         n84747, n84748, n84749, n84750, n84751, n84752, n84753, n84754,
         n84755, n84756, n84757, n84758, n84759, n84760, n84761, n84762,
         n84763, n84764, n84765, n84766, n84767, n84768, n84769, n84770,
         n84771, n84772, n84773, n84774, n84775, n84776, n84777, n84778,
         n84779, n84780, n84781, n84782, n84783, n84784, n84785, n84786,
         n84787, n84788, n84789, n84790, n84791, n84792, n84793, n84794,
         n84795, n84796, n84797, n84798, n84799, n84800, n84801, n84802,
         n84803, n84804, n84805, n84806, n84807, n84808, n84809, n84810,
         n84811, n84812, n84813, n84814, n84815, n84816, n84817, n84818,
         n84819, n84820, n84821, n84822, n84823, n84824, n84825, n84826,
         n84827, n84828, n84829, n84830, n84831, n84832, n84833, n84834,
         n84835, n84836, n84837, n84838, n84839, n84840, n84841, n84842,
         n84843, n84844, n84845, n84846, n84847, n84848, n84849, n84850,
         n84851, n84852, n84853, n84854, n84855, n84856, n84857, n84858,
         n84859, n84860, n84861, n84862, n84863, n84864, n84865, n84866,
         n84867, n84868, n84869, n84870, n84871, n84872, n84873, n84874,
         n84875, n84876, n84877, n84878, n84879, n84880, n84881, n84882,
         n84883, n84884, n84885, n84886, n84887, n84888, n84889, n84890,
         n84891, n84892, n84893, n84894, n84895, n84896, n84897, n84898,
         n84899, n84900, n84901, n84902, n84903, n84904, n84905, n84906,
         n84907, n84908, n84909, n84910, n84911, n84912, n84913, n84914,
         n84915, n84916, n84917, n84918, n84919, n84920, n84921, n84922,
         n84923, n84924, n84925, n84926, n84927, n84928, n84929, n84930,
         n84931, n84932, n84933, n84934, n84935, n84936, n84937, n84938,
         n84939, n84940, n84941, n84942, n84943, n84944, n84945, n84946,
         n84947, n84948, n84949, n84950, n84951, n84952, n84953, n84954,
         n84955, n84956, n84957, n84958, n84959, n84960, n84961, n84962,
         n84963, n84964, n84965, n84966, n84967, n84968, n84969, n84970,
         n84971, n84972, n84973, n84974, n84975, n84976, n84977, n84978,
         n84979, n84980, n84981, n84982, n84983, n84984, n84985, n84986,
         n84987, n84988, n84989, n84990, n84991, n84992, n84993, n84994,
         n84995, n84996, n84997, n84998, n84999, n85000, n85001, n85002,
         n85003, n85004, n85005, n85006, n85007, n85008, n85009, n85010,
         n85011, n85012, n85013, n85014, n85015, n85016, n85017, n85018,
         n85019, n85020, n85021, n85022, n85023, n85024, n85025, n85026,
         n85027, n85028, n85029, n85030, n85031, n85032, n85033, n85034,
         n85035, n85036, n85037, n85038, n85039, n85040, n85041, n85042,
         n85043, n85044, n85045, n85046, n85047, n85048, n85049, n85050,
         n85051, n85052, n85053, n85054, n85055, n85056, n85057, n85058,
         n85059, n85060, n85061, n85062, n85063, n85064, n85065, n85066,
         n85067, n85068, n85069, n85070, n85071, n85072, n85073, n85074,
         n85075, n85076, n85077, n85078, n85079, n85080, n85081, n85082,
         n85083, n85084, n85085, n85086, n85087, n85088, n85089, n85090,
         n85091, n85092, n85093, n85094, n85095, n85096, n85097, n85098,
         n85099, n85100, n85101, n85102, n85103, n85104, n85105, n85106,
         n85107, n85108, n85109, n85110, n85111, n85112, n85113, n85114,
         n85115, n85116, n85117, n85118, n85119, n85120, n85121, n85122,
         n85123, n85124, n85125, n85126, n85127, n85128, n85129, n85130,
         n85131, n85132, n85133, n85134, n85135, n85136, n85137, n85138,
         n85139, n85140, n85141, n85142, n85143, n85144, n85145, n85146,
         n85147, n85148, n85149, n85150, n85151, n85152, n85153, n85154,
         n85155, n85156, n85157, n85158, n85159, n85160, n85161, n85162,
         n85163, n85164, n85165, n85166, n85167, n85168, n85169, n85170,
         n85171, n85172, n85173, n85174, n85175, n85176, n85177, n85178,
         n85179, n85180, n85181, n85182, n85183, n85184, n85185, n85186,
         n85187, n85188, n85189, n85190, n85191, n85192, n85193, n85194,
         n85195, n85196, n85197, n85198, n85199, n85200, n85201, n85202,
         n85203, n85204, n85205, n85206, n85207, n85208, n85209, n85210,
         n85211, n85212, n85213, n85214, n85215, n85216, n85217, n85218,
         n85219, n85220, n85221, n85222, n85223, n85224, n85225, n85226,
         n85227, n85228, n85229, n85230, n85231, n85232, n85233, n85234,
         n85235, n85236, n85237, n85238, n85239, n85240, n85241, n85242,
         n85243, n85244, n85245, n85246, n85247, n85248, n85249, n85250,
         n85251, n85252, n85253, n85254, n85255, n85256, n85257, n85258,
         n85259, n85260, n85261, n85262, n85263, n85264, n85265, n85266,
         n85267, n85268, n85269, n85270, n85271, n85272, n85273, n85274,
         n85275, n85276, n85277, n85278, n85279, n85280, n85281, n85282,
         n85283, n85284, n85285, n85286, n85287, n85288, n85289, n85290,
         n85291, n85292, n85293, n85294, n85295, n85296, n85297, n85298,
         n85299, n85300, n85301, n85302, n85303, n85304, n85305, n85306,
         n85307, n85308, n85309, n85310, n85311, n85312, n85313, n85314,
         n85315, n85316, n85317, n85318, n85319, n85320, n85321, n85322,
         n85323, n85324, n85325, n85326, n85327, n85328, n85329, n85330,
         n85331, n85332, n85333, n85334, n85335, n85336, n85337, n85338,
         n85339, n85340, n85341, n85342, n85343, n85344, n85345, n85346,
         n85347, n85348, n85349, n85350, n85351, n85352, n85353, n85354,
         n85355, n85356, n85357, n85358, n85359, n85360, n85361, n85362,
         n85363, n85364, n85365, n85366, n85367, n85368, n85369, n85370,
         n85371, n85372, n85373, n85374, n85375, n85376, n85377, n85378,
         n85379, n85380, n85381, n85382, n85383, n85384, n85385, n85386,
         n85387, n85388, n85389, n85390, n85391, n85392, n85393, n85394,
         n85395, n85396, n85397, n85398, n85399, n85400, n85401, n85402,
         n85403, n85404, n85405, n85406, n85407, n85408, n85409, n85410,
         n85411, n85412, n85413, n85414, n85415, n85416, n85417, n85418,
         n85419, n85420, n85421, n85422, n85423, n85424, n85425, n85426,
         n85427, n85428, n85429, n85430, n85431, n85432, n85433, n85434,
         n85435, n85436, n85437, n85438, n85439, n85440, n85441, n85442,
         n85443, n85444, n85445, n85446, n85447, n85448, n85449, n85450,
         n85451, n85452, n85453, n85454, n85455, n85456, n85457, n85458,
         n85459, n85460, n85461, n85462, n85463, n85464, n85465, n85466,
         n85467, n85468, n85469, n85470, n85471, n85472, n85473, n85474,
         n85475, n85476, n85477, n85478, n85479, n85480, n85481, n85482,
         n85483, n85484, n85485, n85486, n85487, n85488, n85489, n85490,
         n85491, n85492, n85493, n85494, n85495, n85496, n85497, n85498,
         n85499, n85500, n85501, n85502, n85503, n85504, n85505, n85506,
         n85507, n85508, n85509, n85510, n85511, n85512, n85513, n85514,
         n85515, n85516, n85517, n85518, n85519, n85520, n85521, n85522,
         n85523, n85524, n85525, n85526, n85527, n85528, n85529, n85530,
         n85531, n85532, n85533, n85534, n85535, n85536, n85537, n85538,
         n85539, n85540, n85541, n85542, n85543, n85544, n85545, n85546,
         n85547, n85548, n85549, n85550, n85551, n85552, n85553, n85554,
         n85555, n85556, n85557, n85558, n85559, n85560, n85561, n85562,
         n85563, n85564, n85565, n85566, n85567, n85568, n85569, n85570,
         n85571, n85572, n85573, n85574, n85575, n85576, n85577, n85578,
         n85579, n85580, n85581, n85582, n85583, n85584, n85585, n85586,
         n85587, n85588, n85589, n85590, n85591, n85592, n85593, n85594,
         n85595, n85596, n85597, n85598, n85599, n85600, n85601, n85602,
         n85603, n85604, n85605, n85606, n85607, n85608, n85609, n85610,
         n85611, n85612, n85613, n85614, n85615, n85616, n85617, n85618,
         n85619, n85620, n85621, n85622, n85623, n85624, n85625, n85626,
         n85627, n85628, n85629, n85630, n85631, n85632, n85633, n85634,
         n85635, n85636, n85637, n85638, n85639, n85640, n85641, n85642,
         n85643, n85644, n85645, n85646, n85647, n85648, n85649, n85650,
         n85651, n85652, n85653, n85654, n85655, n85656, n85657, n85658,
         n85659, n85660, n85661, n85662, n85663, n85664, n85665, n85666,
         n85667, n85668, n85669, n85670, n85671, n85672, n85673, n85674,
         n85675, n85676, n85677, n85678, n85679, n85680, n85681, n85682,
         n85683, n85684, n85685, n85686, n85687, n85688, n85689, n85690,
         n85691, n85692, n85693, n85694, n85695, n85696, n85697, n85698,
         n85699, n85700, n85701, n85702, n85703, n85704, n85705, n85706,
         n85707, n85708, n85709, n85710, n85711, n85712, n85713, n85714,
         n85715, n85716, n85717, n85718, n85719, n85720, n85721, n85722,
         n85723, n85724, n85725, n85726, n85727, n85728, n85729, n85730,
         n85731, n85732, n85733, n85734, n85735, n85736, n85737, n85738,
         n85739, n85740, n85741, n85742, n85743, n85744, n85745, n85746,
         n85747, n85748, n85749, n85750, n85751, n85752, n85753, n85754,
         n85755, n85756, n85757, n85758, n85759, n85760, n85761, n85762,
         n85763, n85764, n85765, n85766, n85767, n85768, n85769, n85770,
         n85771, n85772, n85773, n85774, n85775, n85776, n85777, n85778,
         n85779, n85780, n85781, n85782, n85783, n85784, n85785, n85786,
         n85787, n85788, n85789, n85790, n85791, n85792, n85793, n85794,
         n85795, n85796, n85797, n85798, n85799, n85800, n85801, n85802,
         n85803, n85804, n85805, n85806, n85807, n85808, n85809, n85810,
         n85811, n85812, n85813, n85814, n85815, n85816, n85817, n85818,
         n85819, n85820, n85821, n85822, n85823, n85824, n85825, n85826,
         n85827, n85828, n85829, n85830, n85831, n85832, n85833, n85834,
         n85835, n85836, n85837, n85838, n85839, n85840, n85841, n85842,
         n85843, n85844, n85845, n85846, n85847, n85848, n85849, n85850,
         n85851, n85852, n85853, n85854, n85855, n85856, n85857, n85858,
         n85859, n85860, n85861, n85862, n85863, n85864, n85865, n85866,
         n85867, n85868, n85869, n85870, n85871, n85872, n85873, n85874,
         n85875, n85876, n85877, n85878, n85879, n85880, n85881, n85882,
         n85883, n85884, n85885, n85886, n85887, n85888, n85889, n85890,
         n85891, n85892, n85893, n85894, n85895, n85896, n85897, n85898,
         n85899, n85900, n85901, n85902, n85903, n85904, n85905, n85906,
         n85907, n85908, n85909, n85910, n85911, n85912, n85913, n85914,
         n85915, n85916, n85917, n85918, n85919, n85920, n85921, n85922,
         n85923, n85924, n85925, n85926, n85927, n85928, n85929, n85930,
         n85931, n85932, n85933, n85934, n85935, n85936, n85937, n85938,
         n85939, n85940, n85941, n85942, n85943, n85944, n85945, n85946,
         n85947, n85948, n85949, n85950, n85951, n85952, n85953, n85954,
         n85955, n85956, n85957, n85958, n85959, n85960, n85961, n85962,
         n85963, n85964, n85965, n85966, n85967, n85968, n85969, n85970,
         n85971, n85972, n85973, n85974, n85975, n85976, n85977, n85978,
         n85979, n85980, n85981, n85982, n85983, n85984, n85985, n85986,
         n85987, n85988, n85989, n85990, n85991, n85992, n85993, n85994,
         n85995, n85996, n85997, n85998, n85999, n86000, n86001, n86002,
         n86003, n86004, n86005, n86006, n86007, n86008, n86009, n86010,
         n86011, n86012, n86013, n86014, n86015, n86016, n86017, n86018,
         n86019, n86020, n86021, n86022, n86023, n86024, n86025, n86026,
         n86027, n86028, n86029, n86030, n86031, n86032, n86033, n86034,
         n86035, n86036, n86037, n86038, n86039, n86040, n86041, n86042,
         n86043, n86044, n86045, n86046, n86047, n86048, n86049, n86050,
         n86051, n86052, n86053, n86054, n86055, n86056, n86057, n86058,
         n86059, n86060, n86061, n86062, n86063, n86064, n86065, n86066,
         n86067, n86068, n86069, n86070, n86071, n86072, n86073, n86074,
         n86075, n86076, n86077, n86078, n86079, n86080, n86081, n86082,
         n86083, n86084, n86085, n86086, n86087, n86088, n86089, n86090,
         n86091, n86092, n86093, n86094, n86095, n86096, n86097, n86098,
         n86099, n86100, n86101, n86102, n86103, n86104, n86105, n86106,
         n86107, n86108, n86109, n86110, n86111, n86112, n86113, n86114,
         n86115, n86116, n86117, n86118, n86119, n86120, n86121, n86122,
         n86123, n86124, n86125, n86126, n86127, n86128, n86129, n86130,
         n86131, n86132, n86133, n86134, n86135, n86136, n86137, n86138,
         n86139, n86140, n86141, n86142, n86143, n86144, n86145, n86146,
         n86147, n86148, n86149, n86150, n86151, n86152, n86153, n86154,
         n86155, n86156, n86157, n86158, n86159, n86160, n86161, n86162,
         n86163, n86164, n86165, n86166, n86167, n86168, n86169, n86170,
         n86171, n86172, n86173, n86174, n86175, n86176, n86177, n86178,
         n86179, n86180, n86181, n86182, n86183, n86184, n86185, n86186,
         n86187, n86188, n86189, n86190, n86191, n86192, n86193, n86194,
         n86195, n86196, n86197, n86198, n86199, n86200, n86201, n86202,
         n86203, n86204, n86205, n86206, n86207, n86208, n86209, n86210,
         n86211, n86212, n86213, n86214, n86215, n86216, n86217, n86218,
         n86219, n86220, n86221, n86222, n86223, n86224, n86225, n86226,
         n86227, n86228, n86229, n86230, n86231, n86232, n86233, n86234,
         n86235, n86236, n86237, n86238, n86239, n86240, n86241, n86242,
         n86243, n86244, n86245, n86246, n86247, n86248, n86249, n86250,
         n86251, n86252, n86253, n86254, n86255, n86256, n86257, n86258,
         n86259, n86260, n86261, n86262, n86263, n86264, n86265, n86266,
         n86267, n86268, n86269, n86270, n86271, n86272, n86273, n86274,
         n86275, n86276, n86277, n86278, n86279, n86280, n86281, n86282,
         n86283, n86284, n86285, n86286, n86287, n86288, n86289, n86290,
         n86291, n86292, n86293, n86294, n86295, n86296, n86297, n86298,
         n86299, n86300, n86301, n86302, n86303, n86304, n86305, n86306,
         n86307, n86308, n86309, n86310, n86311, n86312, n86313, n86314,
         n86315, n86316, n86317, n86318, n86319, n86320, n86321, n86322,
         n86323, n86324, n86325, n86326, n86327, n86328, n86329, n86330,
         n86331, n86332, n86333, n86334, n86335, n86336, n86337, n86338,
         n86339, n86340, n86341, n86342, n86343, n86344, n86345, n86346,
         n86347, n86348, n86349, n86350, n86351, n86352, n86353, n86354,
         n86355, n86356, n86357, n86358, n86359, n86360, n86361, n86362,
         n86363, n86364, n86365, n86366, n86367, n86368, n86369, n86370,
         n86371, n86372, n86373, n86374, n86375, n86376, n86377, n86378,
         n86379, n86380, n86381, n86382, n86383, n86384, n86385, n86386,
         n86387, n86388, n86389, n86390, n86391, n86392, n86393, n86394,
         n86395, n86396, n86397, n86398, n86399, n86400, n86401, n86402,
         n86403, n86404, n86405, n86406, n86407, n86408, n86409, n86410,
         n86411, n86412, n86413, n86414, n86415, n86416, n86417, n86418,
         n86419, n86420, n86421, n86422, n86423, n86424, n86425, n86426,
         n86427, n86428, n86429, n86430, n86431, n86432, n86433, n86434,
         n86435, n86436, n86437, n86438, n86439, n86440, n86441, n86442,
         n86443, n86444, n86445, n86446, n86447, n86448, n86449, n86450,
         n86451, n86452, n86453, n86454, n86455, n86456, n86457, n86458,
         n86459, n86460, n86461, n86462, n86463, n86464, n86465, n86466,
         n86467, n86468, n86469, n86470, n86471, n86472, n86473, n86474,
         n86475, n86476, n86477, n86478, n86479, n86480, n86481, n86482,
         n86483, n86484, n86485, n86486, n86487, n86488, n86489, n86490,
         n86491, n86492, n86493, n86494, n86495, n86496, n86497, n86498,
         n86499, n86500, n86501, n86502, n86503, n86504, n86505, n86506,
         n86507, n86508, n86509, n86510, n86511, n86512, n86513, n86514,
         n86515, n86516, n86517, n86518, n86519, n86520, n86521, n86522,
         n86523, n86524, n86525, n86526, n86527, n86528, n86529, n86530,
         n86531, n86532, n86533, n86534, n86535, n86536, n86537, n86538,
         n86539, n86540, n86541, n86542, n86543, n86544, n86545, n86546,
         n86547, n86548, n86549, n86550, n86551, n86552, n86553, n86554,
         n86555, n86556, n86557, n86558, n86559, n86560, n86561, n86562,
         n86563, n86564, n86565, n86566, n86567, n86568, n86569, n86570,
         n86571, n86572, n86573, n86574, n86575, n86576, n86577, n86578,
         n86579, n86580, n86581, n86582, n86583, n86584, n86585, n86586,
         n86587, n86588, n86589, n86590, n86591, n86592, n86593, n86594,
         n86595, n86596, n86597, n86598, n86599, n86600, n86601, n86602,
         n86603, n86604, n86605, n86606, n86607, n86608, n86609, n86610,
         n86611, n86612, n86613, n86614, n86615, n86616, n86617, n86618,
         n86619, n86620, n86621, n86622, n86623, n86624, n86625, n86626,
         n86627, n86628, n86629, n86630, n86631, n86632, n86633, n86634,
         n86635, n86636, n86637, n86638, n86639, n86640, n86641, n86642,
         n86643, n86644, n86645, n86646, n86647, n86648, n86649, n86650,
         n86651, n86652, n86653, n86654, n86655, n86656, n86657, n86658,
         n86659, n86660, n86661, n86662, n86663, n86664, n86665, n86666,
         n86667, n86668, n86669, n86670, n86671, n86672, n86673, n86674,
         n86675, n86676, n86677, n86678, n86679, n86680, n86681, n86682,
         n86683, n86684, n86685, n86686, n86687, n86688, n86689, n86690,
         n86691, n86692, n86693, n86694, n86695, n86696, n86697, n86698,
         n86699, n86700, n86701, n86702, n86703, n86704, n86705, n86706,
         n86707, n86708, n86709, n86710, n86711, n86712, n86713, n86714,
         n86715, n86716, n86717, n86718, n86719, n86720, n86721, n86722,
         n86723, n86724, n86725, n86726, n86727, n86728, n86729, n86730,
         n86731, n86732, n86733, n86734, n86735, n86736, n86737, n86738,
         n86739, n86740, n86741, n86742, n86743, n86744, n86745, n86746,
         n86747, n86748, n86749, n86750, n86751, n86752, n86753, n86754,
         n86755, n86756, n86757, n86758, n86759, n86760, n86761, n86762,
         n86763, n86764, n86765, n86766, n86767, n86768, n86769, n86770,
         n86771, n86772, n86773, n86774, n86775, n86776, n86777, n86778,
         n86779, n86780, n86781, n86782, n86783, n86784, n86785, n86786,
         n86787, n86788, n86789, n86790, n86791, n86792, n86793, n86794,
         n86795, n86796, n86797, n86798, n86799, n86800, n86801, n86802,
         n86803, n86804, n86805, n86806, n86807, n86808, n86809, n86810,
         n86811, n86812, n86813, n86814, n86815, n86816, n86817, n86818,
         n86819, n86820, n86821, n86822, n86823, n86824, n86825, n86826,
         n86827, n86828, n86829, n86830, n86831, n86832, n86833, n86834,
         n86835, n86836, n86837, n86838, n86839, n86840, n86841, n86842,
         n86843, n86844, n86845, n86846, n86847, n86848, n86849, n86850,
         n86851, n86852, n86853, n86854, n86855, n86856, n86857, n86858,
         n86859, n86860, n86861, n86862, n86863, n86864, n86865, n86866,
         n86867, n86868, n86869, n86870, n86871, n86872, n86873, n86874,
         n86875, n86876, n86877, n86878, n86879, n86880, n86881, n86882,
         n86883, n86884, n86885, n86886, n86887, n86888, n86889, n86890,
         n86891, n86892, n86893, n86894, n86895, n86896, n86897, n86898,
         n86899, n86900, n86901, n86902, n86903, n86904, n86905, n86906,
         n86907, n86908, n86909, n86910, n86911, n86912, n86913, n86914,
         n86915, n86916, n86917, n86918, n86919, n86920, n86921, n86922,
         n86923, n86924, n86925, n86926, n86927, n86928, n86929, n86930,
         n86931, n86932, n86933, n86934, n86935, n86936, n86937, n86938,
         n86939, n86940, n86941, n86942, n86943, n86944, n86945, n86946,
         n86947, n86948, n86949, n86950, n86951, n86952, n86953, n86954,
         n86955, n86956, n86957, n86958, n86959, n86960, n86961, n86962,
         n86963, n86964, n86965, n86966, n86967, n86968, n86969, n86970,
         n86971, n86972, n86973, n86974, n86975, n86976, n86977, n86978,
         n86979, n86980, n86981, n86982, n86983, n86984, n86985, n86986,
         n86987, n86988, n86989, n86990, n86991, n86992, n86993, n86994,
         n86995, n86996, n86997, n86998, n86999, n87000, n87001, n87002,
         n87003, n87004, n87005, n87006, n87007, n87008, n87009, n87010,
         n87011, n87012, n87013, n87014, n87015, n87016, n87017, n87018,
         n87019, n87020, n87021, n87022, n87023, n87024, n87025, n87026,
         n87027, n87028, n87029, n87030, n87031, n87032, n87033, n87034,
         n87035, n87036, n87037, n87038, n87039, n87040, n87041, n87042,
         n87043, n87044, n87045, n87046, n87047, n87048, n87049, n87050,
         n87051, n87052, n87053, n87054, n87055, n87056, n87057, n87058,
         n87059, n87060, n87061, n87062, n87063, n87064, n87065, n87066,
         n87067, n87068, n87069, n87070, n87071, n87072, n87073, n87074,
         n87075, n87076, n87077, n87078, n87079, n87080, n87081, n87082,
         n87083, n87084, n87085, n87086, n87087, n87088, n87089, n87090,
         n87091, n87092, n87093, n87094, n87095, n87096, n87097, n87098,
         n87099, n87100, n87101, n87102, n87103, n87104, n87105, n87106,
         n87107, n87108, n87109, n87110, n87111, n87112, n87113, n87114,
         n87115, n87116, n87117, n87118, n87119, n87120, n87121, n87122,
         n87123, n87124, n87125, n87126, n87127, n87128, n87129, n87130,
         n87131, n87132, n87133, n87134, n87135, n87136, n87137, n87138,
         n87139, n87140, n87141, n87142, n87143, n87144, n87145, n87146,
         n87147, n87148, n87149, n87150, n87151, n87152, n87153, n87154,
         n87155, n87156, n87157, n87158, n87159, n87160, n87161, n87162,
         n87163, n87164, n87165, n87166, n87167, n87168, n87169, n87170,
         n87171, n87172, n87173, n87174, n87175, n87176, n87177, n87178,
         n87179, n87180, n87181, n87182, n87183, n87184, n87185, n87186,
         n87187, n87188, n87189, n87190, n87191, n87192, n87193, n87194,
         n87195, n87196, n87197, n87198, n87199, n87200, n87201, n87202,
         n87203, n87204, n87205, n87206, n87207, n87208, n87209, n87210,
         n87211, n87212, n87213, n87214, n87215, n87216, n87217, n87218,
         n87219, n87220, n87221, n87222, n87223, n87224, n87225, n87226,
         n87227, n87228, n87229, n87230, n87231, n87232, n87233, n87234,
         n87235, n87236, n87237, n87238, n87239, n87240, n87241, n87242,
         n87243, n87244, n87245, n87246, n87247, n87248, n87249, n87250,
         n87251, n87252, n87253, n87254, n87255, n87256, n87257, n87258,
         n87259, n87260, n87261, n87262, n87263, n87264, n87265, n87266,
         n87267, n87268, n87269, n87270, n87271, n87272, n87273, n87274,
         n87275, n87276, n87277, n87278, n87279, n87280, n87281, n87282,
         n87283, n87284, n87285, n87286, n87287, n87288, n87289, n87290,
         n87291, n87292, n87293, n87294, n87295, n87296, n87297, n87298,
         n87299, n87300, n87301, n87302, n87303, n87304, n87305, n87306,
         n87307, n87308, n87309, n87310, n87311, n87312, n87313, n87314,
         n87315, n87316, n87317, n87318, n87319, n87320, n87321, n87322,
         n87323, n87324, n87325, n87326, n87327, n87328, n87329, n87330,
         n87331, n87332, n87333, n87334, n87335, n87336, n87337, n87338,
         n87339, n87340, n87341, n87342, n87343, n87344, n87345, n87346,
         n87347, n87348, n87349, n87350, n87351, n87352, n87353, n87354,
         n87355, n87356, n87357, n87358, n87359, n87360, n87361, n87362,
         n87363, n87364, n87365, n87366, n87367, n87368, n87369, n87370,
         n87371, n87372, n87373, n87374, n87375, n87376, n87377, n87378,
         n87379, n87380, n87381, n87382, n87383, n87384, n87385, n87386,
         n87387, n87388, n87389, n87390, n87391, n87392, n87393, n87394,
         n87395, n87396, n87397, n87398, n87399, n87400, n87401, n87402,
         n87403, n87404, n87405, n87406, n87407, n87408, n87409, n87410,
         n87411, n87412, n87413, n87414, n87415, n87416, n87417, n87418,
         n87419, n87420, n87421, n87422, n87423, n87424, n87425, n87426,
         n87427, n87428, n87429, n87430, n87431, n87432, n87433, n87434,
         n87435, n87436, n87437, n87438, n87439, n87440, n87441, n87442,
         n87443, n87444, n87445, n87446, n87447, n87448, n87449, n87450,
         n87451, n87452, n87453, n87454, n87455, n87456, n87457, n87458,
         n87459, n87460, n87461, n87462, n87463, n87464, n87465, n87466,
         n87467, n87468, n87469, n87470, n87471, n87472, n87473, n87474,
         n87475, n87476, n87477, n87478, n87479, n87480, n87481, n87482,
         n87483, n87484, n87485, n87486, n87487, n87488, n87489, n87490,
         n87491, n87492, n87493, n87494, n87495, n87496, n87497, n87498,
         n87499, n87500, n87501, n87502, n87503, n87504, n87505, n87506,
         n87507, n87508, n87509, n87510, n87511, n87512, n87513, n87514,
         n87515, n87516, n87517, n87518, n87519, n87520, n87521, n87522,
         n87523, n87524, n87525, n87526, n87527, n87528, n87529, n87530,
         n87531, n87532, n87533, n87534, n87535, n87536, n87537, n87538,
         n87539, n87540, n87541, n87542, n87543, n87544, n87545, n87546,
         n87547, n87548, n87549, n87550, n87551, n87552, n87553, n87554,
         n87555, n87556, n87557, n87558, n87559, n87560, n87561, n87562,
         n87563, n87564, n87565, n87566, n87567, n87568, n87569, n87570,
         n87571, n87572, n87573, n87574, n87575, n87576, n87577, n87578,
         n87579, n87580, n87581, n87582, n87583, n87584, n87585, n87586,
         n87587, n87588, n87589, n87590, n87591, n87592, n87593, n87594,
         n87595, n87596, n87597, n87598, n87599, n87600, n87601, n87602,
         n87603, n87604, n87605, n87606, n87607, n87608, n87609, n87610,
         n87611, n87612, n87613, n87614, n87615, n87616, n87617, n87618,
         n87619, n87620, n87621, n87622, n87623, n87624, n87625, n87626,
         n87627, n87628, n87629, n87630, n87631, n87632, n87633, n87634,
         n87635, n87636, n87637, n87638, n87639, n87640, n87641, n87642,
         n87643, n87644, n87645, n87646, n87647, n87648, n87649, n87650,
         n87651, n87652, n87653, n87654, n87655, n87656, n87657, n87658,
         n87659, n87660, n87661, n87662, n87663, n87664, n87665, n87666,
         n87667, n87668, n87669, n87670, n87671, n87672, n87673, n87674,
         n87675, n87676, n87677, n87678, n87679, n87680, n87681, n87682,
         n87683, n87684, n87685, n87686, n87687, n87688, n87689, n87690,
         n87691, n87692, n87693, n87694, n87695, n87696, n87697, n87698,
         n87699, n87700, n87701, n87702, n87703, n87704, n87705, n87706,
         n87707, n87708, n87709, n87710, n87711, n87712, n87713, n87714,
         n87715, n87716, n87717, n87718, n87719, n87720, n87721, n87722,
         n87723, n87724, n87725, n87726, n87727, n87728, n87729, n87730,
         n87731, n87732, n87733, n87734, n87735, n87736, n87737, n87738,
         n87739, n87740, n87741, n87742, n87743, n87744, n87745, n87746,
         n87747, n87748, n87749, n87750, n87751, n87752, n87753, n87754,
         n87755, n87756, n87757, n87758, n87759, n87760, n87761, n87762,
         n87763, n87764, n87765, n87766, n87767, n87768, n87769, n87770,
         n87771, n87772, n87773, n87774, n87775, n87776, n87777, n87778,
         n87779, n87780, n87781, n87782, n87783, n87784, n87785, n87786,
         n87787, n87788, n87789, n87790, n87791, n87792, n87793, n87794,
         n87795, n87796, n87797, n87798, n87799, n87800, n87801, n87802,
         n87803, n87804, n87805, n87806, n87807, n87808, n87809, n87810,
         n87811, n87812, n87813, n87814, n87815, n87816, n87817, n87818,
         n87819, n87820, n87821, n87822, n87823, n87824, n87825, n87826,
         n87827, n87828, n87829, n87830, n87831, n87832, n87833, n87834,
         n87835, n87836, n87837, n87838, n87839, n87840, n87841, n87842,
         n87843, n87844, n87845, n87846, n87847, n87848, n87849, n87850,
         n87851, n87852, n87853, n87854, n87855, n87856, n87857, n87858,
         n87859, n87860, n87861, n87862, n87863, n87864, n87865, n87866,
         n87867, n87868, n87869, n87870, n87871, n87872, n87873, n87874,
         n87875, n87876, n87877, n87878, n87879, n87880, n87881, n87882,
         n87883, n87884, n87885, n87886, n87887, n87888, n87889, n87890,
         n87891, n87892, n87893, n87894, n87895, n87896, n87897, n87898,
         n87899, n87900, n87901, n87902, n87903, n87904, n87905, n87906,
         n87907, n87908, n87909, n87910, n87911, n87912, n87913, n87914,
         n87915, n87916, n87917, n87918, n87919, n87920, n87921, n87922,
         n87923, n87924, n87925, n87926, n87927, n87928, n87929, n87930,
         n87931, n87932, n87933, n87934, n87935, n87936, n87937, n87938,
         n87939, n87940, n87941, n87942, n87943, n87944, n87945, n87946,
         n87947, n87948, n87949, n87950, n87951, n87952, n87953, n87954,
         n87955, n87956, n87957, n87958, n87959, n87960, n87961, n87962,
         n87963, n87964, n87965, n87966, n87967, n87968, n87969, n87970,
         n87971, n87972, n87973, n87974, n87975, n87976, n87977, n87978,
         n87979, n87980, n87981, n87982, n87983, n87984, n87985, n87986,
         n87987, n87988, n87989, n87990, n87991, n87992, n87993, n87994,
         n87995, n87996, n87997, n87998, n87999, n88000, n88001, n88002,
         n88003, n88004, n88005, n88006, n88007, n88008, n88009, n88010,
         n88011, n88012, n88013, n88014, n88015, n88016, n88017, n88018,
         n88019, n88020, n88021, n88022, n88023, n88024, n88025, n88026,
         n88027, n88028, n88029, n88030, n88031, n88032, n88033, n88034,
         n88035, n88036, n88037, n88038, n88039, n88040, n88041, n88042,
         n88043, n88044, n88045, n88046, n88047, n88048, n88049, n88050,
         n88051, n88052, n88053, n88054, n88055, n88056, n88057, n88058,
         n88059, n88060, n88061, n88062, n88063, n88064, n88065, n88066,
         n88067, n88068, n88069, n88070, n88071, n88072, n88073, n88074,
         n88075, n88076, n88077, n88078, n88079, n88080, n88081, n88082,
         n88083, n88084, n88085, n88086, n88087, n88088, n88089, n88090,
         n88091, n88092, n88093, n88094, n88095, n88096, n88097, n88098,
         n88099, n88100, n88101, n88102, n88103, n88104, n88105, n88106,
         n88107, n88108, n88109, n88110, n88111, n88112, n88113, n88114,
         n88115, n88116, n88117, n88118, n88119, n88120, n88121, n88122,
         n88123, n88124, n88125, n88126, n88127, n88128, n88129, n88130,
         n88131, n88132, n88133, n88134, n88135, n88136, n88137, n88138,
         n88139, n88140, n88141, n88142, n88143, n88144, n88145, n88146,
         n88147, n88148, n88149, n88150, n88151, n88152, n88153, n88154,
         n88155, n88156, n88157, n88158, n88159, n88160, n88161, n88162,
         n88163, n88164, n88165, n88166, n88167, n88168, n88169, n88170,
         n88171, n88172, n88173, n88174, n88175, n88176, n88177, n88178,
         n88179, n88180, n88181, n88182, n88183, n88184, n88185, n88186,
         n88187, n88188, n88189, n88190, n88191, n88192, n88193, n88194,
         n88195, n88196, n88197, n88198, n88199, n88200, n88201, n88202,
         n88203, n88204, n88205, n88206, n88207, n88208, n88209, n88210,
         n88211, n88212, n88213, n88214, n88215, n88216, n88217, n88218,
         n88219, n88220, n88221, n88222, n88223, n88224, n88225, n88226,
         n88227, n88228, n88229, n88230, n88231, n88232, n88233, n88234,
         n88235, n88236, n88237, n88238, n88239, n88240, n88241, n88242,
         n88243, n88244, n88245, n88246, n88247, n88248, n88249, n88250,
         n88251, n88252, n88253, n88254, n88255, n88256, n88257, n88258,
         n88259, n88260, n88261, n88262, n88263, n88264, n88265, n88266,
         n88267, n88268, n88269, n88270, n88271, n88272, n88273, n88274,
         n88275, n88276, n88277, n88278, n88279, n88280, n88281, n88282,
         n88283, n88284, n88285, n88286, n88287, n88288, n88289, n88290,
         n88291, n88292, n88293, n88294, n88295, n88296, n88297, n88298,
         n88299, n88300, n88301, n88302, n88303, n88304, n88305, n88306,
         n88307, n88308, n88309, n88310, n88311, n88312, n88313, n88314,
         n88315, n88316, n88317, n88318, n88319, n88320, n88321, n88322,
         n88323, n88324, n88325, n88326, n88327, n88328, n88329, n88330,
         n88331, n88332, n88333, n88334, n88335, n88336, n88337, n88338,
         n88339, n88340, n88341, n88342, n88343, n88344, n88345, n88346,
         n88347, n88348, n88349, n88350, n88351, n88352, n88353, n88354,
         n88355, n88356, n88357, n88358, n88359, n88360, n88361, n88362,
         n88363, n88364, n88365, n88366, n88367, n88368, n88369, n88370,
         n88371, n88372, n88373, n88374, n88375, n88376, n88377, n88378,
         n88379, n88380, n88381, n88382, n88383, n88384, n88385, n88386,
         n88387, n88388, n88389, n88390, n88391, n88392, n88393, n88394,
         n88395, n88396, n88397, n88398, n88399, n88400, n88401, n88402,
         n88403, n88404, n88405, n88406, n88407, n88408, n88409, n88410,
         n88411, n88412, n88413, n88414, n88415, n88416, n88417, n88418,
         n88419, n88420, n88421, n88422, n88423, n88424, n88425, n88426,
         n88427, n88428, n88429, n88430, n88431, n88432, n88433, n88434,
         n88435, n88436, n88437, n88438, n88439, n88440, n88441, n88442,
         n88443, n88444, n88445, n88446, n88447, n88448, n88449, n88450,
         n88451, n88452, n88453, n88454, n88455, n88456, n88457, n88458,
         n88459, n88460, n88461, n88462, n88463, n88464, n88465, n88466,
         n88467, n88468, n88469, n88470, n88471, n88472, n88473, n88474,
         n88475, n88476, n88477, n88478, n88479, n88480, n88481, n88482,
         n88483, n88484, n88485, n88486, n88487, n88488, n88489, n88490,
         n88491, n88492, n88493, n88494, n88495, n88496, n88497, n88498,
         n88499, n88500, n88501, n88502, n88503, n88504, n88505, n88506,
         n88507, n88508, n88509, n88510, n88511, n88512, n88513, n88514,
         n88515, n88516, n88517, n88518, n88519, n88520, n88521, n88522,
         n88523, n88524, n88525, n88526, n88527, n88528, n88529, n88530,
         n88531, n88532, n88533, n88534, n88535, n88536, n88537, n88538,
         n88539, n88540, n88541, n88542, n88543, n88544, n88545, n88546,
         n88547, n88548, n88549, n88550, n88551, n88552, n88553, n88554,
         n88555, n88556, n88557, n88558, n88559, n88560, n88561, n88562,
         n88563, n88564, n88565, n88566, n88567, n88568, n88569, n88570,
         n88571, n88572, n88573, n88574, n88575, n88576, n88577, n88578,
         n88579, n88580, n88581, n88582, n88583, n88584, n88585, n88586,
         n88587, n88588, n88589, n88590, n88591, n88592, n88593, n88594,
         n88595, n88596, n88597, n88598, n88599, n88600, n88601, n88602,
         n88603, n88604, n88605, n88606, n88607, n88608, n88609, n88610,
         n88611, n88612, n88613, n88614, n88615, n88616, n88617, n88618,
         n88619, n88620, n88621, n88622, n88623, n88624, n88625, n88626,
         n88627, n88628, n88629, n88630, n88631, n88632, n88633, n88634,
         n88635, n88636, n88637, n88638, n88639, n88640, n88641, n88642,
         n88643, n88644, n88645, n88646, n88647, n88648, n88649, n88650,
         n88651, n88652, n88653, n88654, n88655, n88656, n88657, n88658,
         n88659, n88660, n88661, n88662, n88663, n88664, n88665, n88666,
         n88667, n88668, n88669, n88670, n88671, n88672, n88673, n88674,
         n88675, n88676, n88677, n88678, n88679, n88680, n88681, n88682,
         n88683, n88684, n88685, n88686, n88687, n88688, n88689, n88690,
         n88691, n88692, n88693, n88694, n88695, n88696, n88697, n88698,
         n88699, n88700, n88701, n88702, n88703, n88704, n88705, n88706,
         n88707, n88708, n88709, n88710, n88711, n88712, n88713, n88714,
         n88715, n88716, n88717, n88718, n88719, n88720, n88721, n88722,
         n88723, n88724, n88725, n88726, n88727, n88728, n88729, n88730,
         n88731, n88732, n88733, n88734, n88735, n88736, n88737, n88738,
         n88739, n88740, n88741, n88742, n88743, n88744, n88745, n88746,
         n88747, n88748, n88749, n88750, n88751, n88752, n88753, n88754,
         n88755, n88756, n88757, n88758, n88759, n88760, n88761, n88762,
         n88763, n88764, n88765, n88766, n88767, n88768, n88769, n88770,
         n88771, n88772, n88773, n88774, n88775, n88776, n88777, n88778,
         n88779, n88780, n88781, n88782, n88783, n88784, n88785, n88786,
         n88787, n88788, n88789, n88790, n88791, n88792, n88793, n88794,
         n88795, n88796, n88797, n88798, n88799, n88800, n88801, n88802,
         n88803, n88804, n88805, n88806, n88807, n88808, n88809, n88810,
         n88811, n88812, n88813, n88814, n88815, n88816, n88817, n88818,
         n88819, n88820, n88821, n88822, n88823, n88824, n88825, n88826,
         n88827, n88828, n88829, n88830, n88831, n88832, n88833, n88834,
         n88835, n88836, n88837, n88838, n88839, n88840, n88841, n88842,
         n88843, n88844, n88845, n88846, n88847, n88848, n88849, n88850,
         n88851, n88852, n88853, n88854, n88855, n88856, n88857, n88858,
         n88859, n88860, n88861, n88862, n88863, n88864, n88865, n88866,
         n88867, n88868, n88869, n88870, n88871, n88872, n88873, n88874,
         n88875, n88876, n88877, n88878, n88879, n88880, n88881, n88882,
         n88883, n88884, n88885, n88886, n88887, n88888, n88889, n88890,
         n88891, n88892, n88893, n88894, n88895, n88896, n88897, n88898,
         n88899, n88900, n88901, n88902, n88903, n88904, n88905, n88906,
         n88907, n88908, n88909, n88910, n88911, n88912, n88913, n88914,
         n88915, n88916, n88917, n88918, n88919, n88920, n88921, n88922,
         n88923, n88924, n88925, n88926, n88927, n88928, n88929, n88930,
         n88931, n88932, n88933, n88934, n88935, n88936, n88937, n88938,
         n88939, n88940, n88941, n88942, n88943, n88944, n88945, n88946,
         n88947, n88948, n88949, n88950, n88951, n88952, n88953, n88954,
         n88955, n88956, n88957, n88958, n88959, n88960, n88961, n88962,
         n88963, n88964, n88965, n88966, n88967, n88968, n88969, n88970,
         n88971, n88972, n88973, n88974, n88975, n88976, n88977, n88978,
         n88979, n88980, n88981, n88982, n88983, n88984, n88985, n88986,
         n88987, n88988, n88989, n88990, n88991, n88992, n88993, n88994,
         n88995, n88996, n88997, n88998, n88999, n89000, n89001, n89002,
         n89003, n89004, n89005, n89006, n89007, n89008, n89009, n89010,
         n89011, n89012, n89013, n89014, n89015, n89016, n89017, n89018,
         n89019, n89020, n89021, n89022, n89023, n89024, n89025, n89026,
         n89027, n89028, n89029, n89030, n89031, n89032, n89033, n89034,
         n89035, n89036, n89037, n89038, n89039, n89040, n89041, n89042,
         n89043, n89044, n89045, n89046, n89047, n89048, n89049, n89050,
         n89051, n89052, n89053, n89054, n89055, n89056, n89057, n89058,
         n89059, n89060, n89061, n89062, n89063, n89064, n89065, n89066,
         n89067, n89068, n89069, n89070, n89071, n89072, n89073, n89074,
         n89075, n89076, n89077, n89078, n89079, n89080, n89081, n89082,
         n89083, n89084, n89085, n89086, n89087, n89088, n89089, n89090,
         n89091, n89092, n89093, n89094, n89095, n89096, n89097, n89098,
         n89099, n89100, n89101, n89102, n89103, n89104, n89105, n89106,
         n89107, n89108, n89109, n89110, n89111, n89112, n89113, n89114,
         n89115, n89116, n89117, n89118, n89119, n89120, n89121, n89122,
         n89123, n89124, n89125, n89126, n89127, n89128, n89129, n89130,
         n89131, n89132, n89133, n89134, n89135, n89136, n89137, n89138,
         n89139, n89140, n89141, n89142, n89143, n89144, n89145, n89146,
         n89147, n89148, n89149, n89150, n89151, n89152, n89153, n89154,
         n89155, n89156, n89157, n89158, n89159, n89160, n89161, n89162,
         n89163, n89164, n89165, n89166, n89167, n89168, n89169, n89170,
         n89171, n89172, n89173, n89174, n89175, n89176, n89177, n89178,
         n89179, n89180, n89181, n89182, n89183, n89184, n89185, n89186,
         n89187, n89188, n89189, n89190, n89191, n89192, n89193, n89194,
         n89195, n89196, n89197, n89198, n89199, n89200, n89201, n89202,
         n89203, n89204, n89205, n89206, n89207, n89208, n89209, n89210,
         n89211, n89212, n89213, n89214, n89215, n89216, n89217, n89218,
         n89219, n89220, n89221, n89222, n89223, n89224, n89225, n89226,
         n89227, n89228, n89229, n89230, n89231, n89232, n89233, n89234,
         n89235, n89236, n89237, n89238, n89239, n89240, n89241, n89242,
         n89243, n89244, n89245, n89246, n89247, n89248, n89249, n89250,
         n89251, n89252, n89253, n89254, n89255, n89256, n89257, n89258,
         n89259, n89260, n89261, n89262, n89263, n89264, n89265, n89266,
         n89267, n89268, n89269, n89270, n89271, n89272, n89273, n89274,
         n89275, n89276, n89277, n89278, n89279, n89280, n89281, n89282,
         n89283, n89284, n89285, n89286, n89287, n89288, n89289, n89290,
         n89291, n89292, n89293, n89294, n89295, n89296, n89297, n89298,
         n89299, n89300, n89301, n89302, n89303, n89304, n89305, n89306,
         n89307, n89308, n89309, n89310, n89311, n89312, n89313, n89314,
         n89315, n89316, n89317, n89318, n89319, n89320, n89321, n89322,
         n89323, n89324, n89325, n89326, n89327, n89328, n89329, n89330,
         n89331, n89332, n89333, n89334, n89335, n89336, n89337, n89338,
         n89339, n89340, n89341, n89342, n89343, n89344, n89345, n89346,
         n89347, n89348, n89349, n89350, n89351, n89352, n89353, n89354,
         n89355, n89356, n89357, n89358, n89359, n89360, n89361, n89362,
         n89363, n89364, n89365, n89366, n89367, n89368, n89369, n89370,
         n89371, n89372, n89373, n89374, n89375, n89376, n89377, n89378,
         n89379, n89380, n89381, n89382, n89383, n89384, n89385, n89386,
         n89387, n89388, n89389, n89390, n89391, n89392, n89393, n89394,
         n89395, n89396, n89397, n89398, n89399, n89400, n89401, n89402,
         n89403, n89404, n89405, n89406, n89407, n89408, n89409, n89410,
         n89411, n89412, n89413, n89414, n89415, n89416, n89417, n89418,
         n89419, n89420, n89421, n89422, n89423, n89424, n89425, n89426,
         n89427, n89428, n89429, n89430, n89431, n89432, n89433, n89434,
         n89435, n89436, n89437, n89438, n89439, n89440, n89441, n89442,
         n89443, n89444, n89445, n89446, n89447, n89448, n89449, n89450,
         n89451, n89452, n89453, n89454, n89455, n89456, n89457, n89458,
         n89459, n89460, n89461, n89462, n89463, n89464, n89465, n89466,
         n89467, n89468, n89469, n89470, n89471, n89472, n89473, n89474,
         n89475, n89476, n89477, n89478, n89479, n89480, n89481, n89482,
         n89483, n89484, n89485, n89486, n89487, n89488, n89489, n89490,
         n89491, n89492, n89493, n89494, n89495, n89496, n89497, n89498,
         n89499, n89500, n89501, n89502, n89503, n89504, n89505, n89506,
         n89507, n89508, n89509, n89510, n89511, n89512, n89513, n89514,
         n89515, n89516, n89517, n89518, n89519, n89520, n89521, n89522,
         n89523, n89524, n89525, n89526, n89527, n89528, n89529, n89530,
         n89531, n89532, n89533, n89534, n89535, n89536, n89537, n89538,
         n89539, n89540, n89541, n89542, n89543, n89544, n89545, n89546,
         n89547, n89548, n89549, n89550, n89551, n89552, n89553, n89554,
         n89555, n89556, n89557, n89558, n89559, n89560, n89561, n89562,
         n89563, n89564, n89565, n89566, n89567, n89568, n89569, n89570,
         n89571, n89572, n89573, n89574, n89575, n89576, n89577, n89578,
         n89579, n89580, n89581, n89582, n89583, n89584, n89585, n89586,
         n89587, n89588, n89589, n89590, n89591, n89592, n89593, n89594,
         n89595, n89596, n89597, n89598, n89599, n89600, n89601, n89602,
         n89603, n89604, n89605, n89606, n89607, n89608, n89609, n89610,
         n89611, n89612, n89613, n89614, n89615, n89616, n89617, n89618,
         n89619, n89620, n89621, n89622, n89623, n89624, n89625, n89626,
         n89627, n89628, n89629, n89630, n89631, n89632, n89633, n89634,
         n89635, n89636, n89637, n89638, n89639, n89640, n89641, n89642,
         n89643, n89644, n89645, n89646, n89647, n89648, n89649, n89650,
         n89651, n89652, n89653, n89654, n89655, n89656, n89657, n89658,
         n89659, n89660, n89661, n89662, n89663, n89664, n89665, n89666,
         n89667, n89668, n89669, n89670, n89671, n89672, n89673, n89674,
         n89675, n89676, n89677, n89678, n89679, n89680, n89681, n89682,
         n89683, n89684, n89685, n89686, n89687, n89688, n89689, n89690,
         n89691, n89692, n89693, n89694, n89695, n89696, n89697, n89698,
         n89699, n89700, n89701, n89702, n89703, n89704, n89705, n89706,
         n89707, n89708, n89709, n89710, n89711, n89712, n89713, n89714,
         n89715, n89716, n89717, n89718, n89719, n89720, n89721, n89722,
         n89723, n89724, n89725, n89726, n89727, n89728, n89729, n89730,
         n89731, n89732, n89733, n89734, n89735, n89736, n89737, n89738,
         n89739, n89740, n89741, n89742, n89743, n89744, n89745, n89746,
         n89747, n89748, n89749, n89750, n89751, n89752, n89753, n89754,
         n89755, n89756, n89757, n89758, n89759, n89760, n89761, n89762,
         n89763, n89764, n89765, n89766, n89767, n89768, n89769, n89770,
         n89771, n89772, n89773, n89774, n89775, n89776, n89777, n89778,
         n89779, n89780, n89781, n89782, n89783, n89784, n89785, n89786,
         n89787, n89788, n89789, n89790, n89791, n89792, n89793, n89794,
         n89795, n89796, n89797, n89798, n89799, n89800, n89801, n89802,
         n89803, n89804, n89805, n89806, n89807, n89808, n89809, n89810,
         n89811, n89812, n89813, n89814, n89815, n89816, n89817, n89818,
         n89819, n89820, n89821, n89822, n89823, n89824, n89825, n89826,
         n89827, n89828, n89829, n89830, n89831, n89832, n89833, n89834,
         n89835, n89836, n89837, n89838, n89839, n89840, n89841, n89842,
         n89843, n89844, n89845, n89846, n89847, n89848, n89849, n89850,
         n89851, n89852, n89853, n89854, n89855, n89856, n89857, n89858,
         n89859, n89860, n89861, n89862, n89863, n89864, n89865, n89866,
         n89867, n89868, n89869, n89870, n89871, n89872, n89873, n89874,
         n89875, n89876, n89877, n89878, n89879, n89880, n89881, n89882,
         n89883, n89884, n89885, n89886, n89887, n89888, n89889, n89890,
         n89891, n89892, n89893, n89894, n89895, n89896, n89897, n89898,
         n89899, n89900, n89901, n89902, n89903, n89904, n89905, n89906,
         n89907, n89908, n89909, n89910, n89911, n89912, n89913, n89914,
         n89915, n89916, n89917, n89918, n89919, n89920, n89921, n89922,
         n89923, n89924, n89925, n89926, n89927, n89928, n89929, n89930,
         n89931, n89932, n89933, n89934, n89935, n89936, n89937, n89938,
         n89939, n89940, n89941, n89942, n89943, n89944, n89945, n89946,
         n89947, n89948, n89949, n89950, n89951, n89952, n89953, n89954,
         n89955, n89956, n89957, n89958, n89959, n89960, n89961, n89962,
         n89963, n89964, n89965, n89966, n89967, n89968, n89969, n89970,
         n89971, n89972, n89973, n89974, n89975, n89976, n89977, n89978,
         n89979, n89980, n89981, n89982, n89983, n89984, n89985, n89986,
         n89987, n89988, n89989, n89990, n89991, n89992, n89993, n89994,
         n89995, n89996, n89997, n89998, n89999, n90000, n90001, n90002,
         n90003, n90004, n90005, n90006, n90007, n90008, n90009, n90010,
         n90011, n90012, n90013, n90014, n90015, n90016, n90017, n90018,
         n90019, n90020, n90021, n90022, n90023, n90024, n90025, n90026,
         n90027, n90028, n90029, n90030, n90031, n90032, n90033, n90034,
         n90035, n90036, n90037, n90038, n90039, n90040, n90041, n90042,
         n90043, n90044, n90045, n90046, n90047, n90048, n90049, n90050,
         n90051, n90052, n90053, n90054, n90055, n90056, n90057, n90058,
         n90059, n90060, n90061, n90062, n90063, n90064, n90065, n90066,
         n90067, n90068, n90069, n90070, n90071, n90072, n90073, n90074,
         n90075, n90076, n90077, n90078, n90079, n90080, n90081, n90082,
         n90083, n90084, n90085, n90086, n90087, n90088, n90089, n90090,
         n90091, n90092, n90093, n90094, n90095, n90096, n90097, n90098,
         n90099, n90100, n90101, n90102, n90103, n90104, n90105, n90106,
         n90107, n90108, n90109, n90110, n90111, n90112, n90113, n90114,
         n90115, n90116, n90117, n90118, n90119, n90120, n90121, n90122,
         n90123, n90124, n90125, n90126, n90127, n90128, n90129, n90130,
         n90131, n90132, n90133, n90134, n90135, n90136, n90137, n90138,
         n90139, n90140, n90141, n90142, n90143, n90144, n90145, n90146,
         n90147, n90148, n90149, n90150, n90151, n90152, n90153, n90154,
         n90155, n90156, n90157, n90158, n90159, n90160, n90161, n90162,
         n90163, n90164, n90165, n90166, n90167, n90168, n90169, n90170,
         n90171, n90172, n90173, n90174, n90175, n90176, n90177, n90178,
         n90179, n90180, n90181, n90182, n90183, n90184, n90185, n90186,
         n90187, n90188, n90189, n90190, n90191, n90192, n90193, n90194,
         n90195, n90196, n90197, n90198, n90199, n90200, n90201, n90202,
         n90203, n90204, n90205, n90206, n90207, n90208, n90209, n90210,
         n90211, n90212, n90213, n90214, n90215, n90216, n90217, n90218,
         n90219, n90220, n90221, n90222, n90223, n90224, n90225, n90226,
         n90227, n90228, n90229, n90230, n90231, n90232, n90233, n90234,
         n90235, n90236, n90237, n90238, n90239, n90240, n90241, n90242,
         n90243, n90244, n90245, n90246, n90247, n90248, n90249, n90250,
         n90251, n90252, n90253, n90254, n90255, n90256, n90257, n90258,
         n90259, n90260, n90261, n90262, n90263, n90264, n90265, n90266,
         n90267, n90268, n90269, n90270, n90271, n90272, n90273, n90274,
         n90275, n90276, n90277, n90278, n90279, n90280, n90281, n90282,
         n90283, n90284, n90285, n90286, n90287, n90288, n90289, n90290,
         n90291, n90292, n90293, n90294, n90295, n90296, n90297, n90298,
         n90299, n90300, n90301, n90302, n90303, n90304, n90305, n90306,
         n90307, n90308, n90309, n90310, n90311, n90312, n90313, n90314,
         n90315, n90316, n90317, n90318, n90319, n90320, n90321, n90322,
         n90323, n90324, n90325, n90326, n90327, n90328, n90329, n90330,
         n90331, n90332, n90333, n90334, n90335, n90336, n90337, n90338,
         n90339, n90340, n90341, n90342, n90343, n90344, n90345, n90346,
         n90347, n90348, n90349, n90350, n90351, n90352, n90353, n90354,
         n90355, n90356, n90357, n90358, n90359, n90360, n90361, n90362,
         n90363, n90364, n90365, n90366, n90367, n90368, n90369, n90370,
         n90371, n90372, n90373, n90374, n90375, n90376, n90377, n90378,
         n90379, n90380, n90381, n90382, n90383, n90384, n90385, n90386,
         n90387, n90388, n90389, n90390, n90391, n90392, n90393, n90394,
         n90395, n90396, n90397, n90398, n90399, n90400, n90401, n90402,
         n90403, n90404, n90405, n90406, n90407, n90408, n90409, n90410,
         n90411, n90412, n90413, n90414, n90415, n90416, n90417, n90418,
         n90419, n90420, n90421, n90422, n90423, n90424, n90425, n90426,
         n90427, n90428, n90429, n90430, n90431, n90432, n90433, n90434,
         n90435, n90436, n90437, n90438, n90439, n90440, n90441, n90442,
         n90443, n90444, n90445, n90446, n90447, n90448, n90449, n90450,
         n90451, n90452, n90453, n90454, n90455, n90456, n90457, n90458,
         n90459, n90460, n90461, n90462, n90463, n90464, n90465, n90466,
         n90467, n90468, n90469, n90470, n90471, n90472, n90473, n90474,
         n90475, n90476, n90477, n90478, n90479, n90480, n90481, n90482,
         n90483, n90484, n90485, n90486, n90487, n90488, n90489, n90490,
         n90491, n90492, n90493, n90494, n90495, n90496, n90497, n90498,
         n90499, n90500, n90501, n90502, n90503, n90504, n90505, n90506,
         n90507, n90508, n90509, n90510, n90511, n90512, n90513, n90514,
         n90515, n90516, n90517, n90518, n90519, n90520, n90521, n90522,
         n90523, n90524, n90525, n90526, n90527, n90528, n90529, n90530,
         n90531, n90532, n90533, n90534, n90535, n90536, n90537, n90538,
         n90539, n90540, n90541, n90542, n90543, n90544, n90545, n90546,
         n90547, n90548, n90549, n90550, n90551, n90552, n90553, n90554,
         n90555, n90556, n90557, n90558, n90559, n90560, n90561, n90562,
         n90563, n90564, n90565, n90566, n90567, n90568, n90569, n90570,
         n90571, n90572, n90573, n90574, n90575, n90576, n90577, n90578,
         n90579, n90580, n90581, n90582, n90583, n90584, n90585, n90586,
         n90587, n90588, n90589, n90590, n90591, n90592, n90593, n90594,
         n90595, n90596, n90597, n90598, n90599, n90600, n90601, n90602,
         n90603, n90604, n90605, n90606, n90607, n90608, n90609, n90610,
         n90611, n90612, n90613, n90614, n90615, n90616, n90617, n90618,
         n90619, n90620, n90621, n90622, n90623, n90624, n90625, n90626,
         n90627, n90628, n90629, n90630, n90631, n90632, n90633, n90634,
         n90635, n90636, n90637, n90638, n90639, n90640, n90641, n90642,
         n90643, n90644, n90645, n90646, n90647, n90648, n90649, n90650,
         n90651, n90652, n90653, n90654, n90655, n90656, n90657, n90658,
         n90659, n90660, n90661, n90662, n90663, n90664, n90665, n90666,
         n90667, n90668, n90669, n90670, n90671, n90672, n90673, n90674,
         n90675, n90676, n90677, n90678, n90679, n90680, n90681, n90682,
         n90683, n90684, n90685, n90686, n90687, n90688, n90689, n90690,
         n90691, n90692, n90693, n90694, n90695, n90696, n90697, n90698,
         n90699, n90700, n90701, n90702, n90703, n90704, n90705, n90706,
         n90707, n90708, n90709, n90710, n90711, n90712, n90713, n90714,
         n90715, n90716, n90717, n90718, n90719, n90720, n90721, n90722,
         n90723, n90724, n90725, n90726, n90727, n90728, n90729, n90730,
         n90731, n90732, n90733, n90734, n90735, n90736, n90737, n90738,
         n90739, n90740, n90741, n90742, n90743, n90744, n90745, n90746,
         n90747, n90748, n90749, n90750, n90751, n90752, n90753, n90754,
         n90755, n90756, n90757, n90758, n90759, n90760, n90761, n90762,
         n90763, n90764, n90765, n90766, n90767, n90768, n90769, n90770,
         n90771, n90772, n90773, n90774, n90775, n90776, n90777, n90778,
         n90779, n90780, n90781, n90782, n90783, n90784, n90785, n90786,
         n90787, n90788, n90789, n90790, n90791, n90792, n90793, n90794,
         n90795, n90796, n90797, n90798, n90799, n90800, n90801, n90802,
         n90803, n90804, n90805, n90806, n90807, n90808, n90809, n90810,
         n90811, n90812, n90813, n90814, n90815, n90816, n90817, n90818,
         n90819, n90820, n90821, n90822, n90823, n90824, n90825, n90826,
         n90827, n90828, n90829, n90830, n90831, n90832, n90833, n90834,
         n90835, n90836, n90837, n90838, n90839, n90840, n90841, n90842,
         n90843, n90844, n90845, n90846, n90847, n90848, n90849, n90850,
         n90851, n90852, n90853, n90854, n90855, n90856, n90857, n90858,
         n90859, n90860, n90861, n90862, n90863, n90864, n90865, n90866,
         n90867, n90868, n90869, n90870, n90871, n90872, n90873, n90874,
         n90875, n90876, n90877, n90878, n90879, n90880, n90881, n90882,
         n90883, n90884, n90885, n90886, n90887, n90888, n90889, n90890,
         n90891, n90892, n90893, n90894, n90895, n90896, n90897, n90898,
         n90899, n90900, n90901, n90902, n90903, n90904, n90905, n90906,
         n90907, n90908, n90909, n90910, n90911, n90912, n90913, n90914,
         n90915, n90916, n90917, n90918, n90919, n90920, n90921, n90922,
         n90923, n90924, n90925, n90926, n90927, n90928, n90929, n90930,
         n90931, n90932, n90933, n90934, n90935, n90936, n90937, n90938,
         n90939, n90940, n90941, n90942, n90943, n90944, n90945, n90946,
         n90947, n90948, n90949, n90950, n90951, n90952, n90953, n90954,
         n90955, n90956, n90957, n90958, n90959, n90960, n90961, n90962,
         n90963, n90964, n90965, n90966, n90967, n90968, n90969, n90970,
         n90971, n90972, n90973, n90974, n90975, n90976, n90977, n90978,
         n90979, n90980, n90981, n90982, n90983, n90984, n90985, n90986,
         n90987, n90988, n90989, n90990, n90991, n90992, n90993, n90994,
         n90995, n90996, n90997, n90998, n90999, n91000, n91001, n91002,
         n91003, n91004, n91005, n91006, n91007, n91008, n91009, n91010,
         n91011, n91012, n91013, n91014, n91015, n91016, n91017, n91018,
         n91019, n91020, n91021, n91022, n91023, n91024, n91025, n91026,
         n91027, n91028, n91029, n91030, n91031, n91032, n91033, n91034,
         n91035, n91036, n91037, n91038, n91039, n91040, n91041, n91042,
         n91043, n91044, n91045, n91046, n91047, n91048, n91049, n91050,
         n91051, n91052, n91053, n91054, n91055, n91056, n91057, n91058,
         n91059, n91060, n91061, n91062, n91063, n91064, n91065, n91066,
         n91067, n91068, n91069, n91070, n91071, n91072, n91073, n91074,
         n91075, n91076, n91077, n91078, n91079, n91080, n91081, n91082,
         n91083, n91084, n91085, n91086, n91087, n91088, n91089, n91090,
         n91091, n91092, n91093, n91094, n91095, n91096, n91097, n91098,
         n91099, n91100, n91101, n91102, n91103, n91104, n91105, n91106,
         n91107, n91108, n91109, n91110, n91111, n91112, n91113, n91114,
         n91115, n91116, n91117, n91118, n91119, n91120, n91121, n91122,
         n91123, n91124, n91125, n91126, n91127, n91128, n91129, n91130,
         n91131, n91132, n91133, n91134, n91135, n91136, n91137, n91138,
         n91139, n91140, n91141, n91142, n91143, n91144, n91145, n91146,
         n91147, n91148, n91149, n91150, n91151, n91152, n91153, n91154,
         n91155, n91156, n91157, n91158, n91159, n91160, n91161, n91162,
         n91163, n91164, n91165, n91166, n91167, n91168, n91169, n91170,
         n91171, n91172, n91173, n91174, n91175, n91176, n91177, n91178,
         n91179, n91180, n91181, n91182, n91183, n91184, n91185, n91186,
         n91187, n91188, n91189, n91190, n91191, n91192, n91193, n91194,
         n91195, n91196, n91197, n91198, n91199, n91200, n91201, n91202,
         n91203, n91204, n91205, n91206, n91207, n91208, n91209, n91210,
         n91211, n91212, n91213, n91214, n91215, n91216, n91217, n91218,
         n91219, n91220, n91221, n91222, n91223, n91224, n91225, n91226,
         n91227, n91228, n91229, n91230, n91231, n91232, n91233, n91234,
         n91235, n91236, n91237, n91238, n91239, n91240, n91241, n91242,
         n91243, n91244, n91245, n91246, n91247, n91248, n91249, n91250,
         n91251, n91252, n91253, n91254, n91255, n91256, n91257, n91258,
         n91259, n91260, n91261, n91262, n91263, n91264, n91265, n91266,
         n91267, n91268, n91269, n91270, n91271, n91272, n91273, n91274,
         n91275, n91276, n91277, n91278, n91279, n91280, n91281, n91282,
         n91283, n91284, n91285, n91286, n91287, n91288, n91289, n91290,
         n91291, n91292, n91293, n91294, n91295, n91296, n91297, n91298,
         n91299, n91300, n91301, n91302, n91303, n91304, n91305, n91306,
         n91307, n91308, n91309, n91310, n91311, n91312, n91313, n91314,
         n91315, n91316, n91317, n91318, n91319, n91320, n91321, n91322,
         n91323, n91324, n91325, n91326, n91327, n91328, n91329, n91330,
         n91331, n91332, n91333, n91334, n91335, n91336, n91337, n91338,
         n91339, n91340, n91341, n91342, n91343, n91344, n91345, n91346,
         n91347, n91348, n91349, n91350, n91351, n91352, n91353, n91354,
         n91355, n91356, n91357, n91358, n91359, n91360, n91361, n91362,
         n91363, n91364, n91365, n91366, n91367, n91368, n91369, n91370,
         n91371, n91372, n91373, n91374, n91375, n91376, n91377, n91378,
         n91379, n91380, n91381, n91382, n91383, n91384, n91385, n91386,
         n91387, n91388, n91389, n91390, n91391, n91392, n91393, n91394,
         n91395, n91396, n91397, n91398, n91399, n91400, n91401, n91402,
         n91403, n91404, n91405, n91406, n91407, n91408, n91409, n91410,
         n91411, n91412, n91413, n91414, n91415, n91416, n91417, n91418,
         n91419, n91420, n91421, n91422, n91423, n91424, n91425, n91426,
         n91427, n91428, n91429, n91430, n91431, n91432, n91433, n91434,
         n91435, n91436, n91437, n91438, n91439, n91440, n91441, n91442,
         n91443, n91444, n91445, n91446, n91447, n91448, n91449, n91450,
         n91451, n91452, n91453, n91454, n91455, n91456, n91457, n91458,
         n91459, n91460, n91461, n91462, n91463, n91464, n91465, n91466,
         n91467, n91468, n91469, n91470, n91471, n91472, n91473, n91474,
         n91475, n91476, n91477, n91478, n91479, n91480, n91481, n91482,
         n91483, n91484, n91485, n91486, n91487, n91488, n91489, n91490,
         n91491, n91492, n91493, n91494, n91495, n91496, n91497, n91498,
         n91499, n91500, n91501, n91502, n91503, n91504, n91505, n91506,
         n91507, n91508, n91509, n91510, n91511, n91512, n91513, n91514,
         n91515, n91516, n91517, n91518, n91519, n91520, n91521, n91522,
         n91523, n91524, n91525, n91526, n91527, n91528, n91529, n91530,
         n91531, n91532, n91533, n91534, n91535, n91536, n91537, n91538,
         n91539, n91540, n91541, n91542, n91543, n91544, n91545, n91546,
         n91547, n91548, n91549, n91550, n91551, n91552, n91553, n91554,
         n91555, n91556, n91557, n91558, n91559, n91560, n91561, n91562,
         n91563, n91564, n91565, n91566, n91567, n91568, n91569, n91570,
         n91571, n91572, n91573, n91574, n91575, n91576, n91577, n91578,
         n91579, n91580, n91581, n91582, n91583, n91584, n91585, n91586,
         n91587, n91588, n91589, n91590, n91591, n91592, n91593, n91594,
         n91595, n91596, n91597, n91598, n91599, n91600, n91601, n91602,
         n91603, n91604, n91605, n91606, n91607, n91608, n91609, n91610,
         n91611, n91612, n91613, n91614, n91615, n91616, n91617, n91618,
         n91619, n91620, n91621, n91622, n91623, n91624, n91625, n91626,
         n91627, n91628, n91629, n91630, n91631, n91632, n91633, n91634,
         n91635, n91636, n91637, n91638, n91639, n91640, n91641, n91642,
         n91643, n91644, n91645, n91646, n91647, n91648, n91649, n91650,
         n91651, n91652, n91653, n91654, n91655, n91656, n91657, n91658,
         n91659, n91660, n91661, n91662, n91663, n91664, n91665, n91666,
         n91667, n91668, n91669, n91670, n91671, n91672, n91673, n91674,
         n91675, n91676, n91677, n91678, n91679, n91680, n91681, n91682,
         n91683, n91684, n91685, n91686, n91687, n91688, n91689, n91690,
         n91691, n91692, n91693, n91694, n91695, n91696, n91697, n91698,
         n91699, n91700, n91701, n91702, n91703, n91704, n91705, n91706,
         n91707, n91708, n91709, n91710, n91711, n91712, n91713, n91714,
         n91715, n91716, n91717, n91718, n91719, n91720, n91721, n91722,
         n91723, n91724, n91725, n91726, n91727, n91728, n91729, n91730,
         n91731, n91732, n91733, n91734, n91735, n91736, n91737, n91738,
         n91739, n91740, n91741, n91742, n91743, n91744, n91745, n91746,
         n91747, n91748, n91749, n91750, n91751, n91752, n91753, n91754,
         n91755, n91756, n91757, n91758, n91759, n91760, n91761, n91762,
         n91763, n91764, n91765, n91766, n91767, n91768, n91769, n91770,
         n91771, n91772, n91773, n91774, n91775, n91776, n91777, n91778,
         n91779, n91780, n91781, n91782, n91783, n91784, n91785, n91786,
         n91787, n91788, n91789, n91790, n91791, n91792, n91793, n91794,
         n91795, n91796, n91797, n91798, n91799, n91800, n91801, n91802,
         n91803, n91804, n91805, n91806, n91807, n91808, n91809, n91810,
         n91811, n91812, n91813, n91814, n91815, n91816, n91817, n91818,
         n91819, n91820, n91821, n91822, n91823, n91824, n91825, n91826,
         n91827, n91828, n91829, n91830, n91831, n91832, n91833, n91834,
         n91835, n91836, n91837, n91838, n91839, n91840, n91841, n91842,
         n91843, n91844, n91845, n91846, n91847, n91848, n91849, n91850,
         n91851, n91852, n91853, n91854, n91855, n91856, n91857, n91858,
         n91859, n91860, n91861, n91862, n91863, n91864, n91865, n91866,
         n91867, n91868, n91869, n91870, n91871, n91872, n91873, n91874,
         n91875, n91876, n91877, n91878, n91879, n91880, n91881, n91882,
         n91883, n91884, n91885, n91886, n91887, n91888, n91889, n91890,
         n91891, n91892, n91893, n91894, n91895, n91896, n91897, n91898,
         n91899, n91900, n91901, n91902, n91903, n91904, n91905, n91906,
         n91907, n91908, n91909, n91910, n91911, n91912, n91913, n91914,
         n91915, n91916, n91917, n91918, n91919, n91920, n91921, n91922,
         n91923, n91924, n91925, n91926, n91927, n91928, n91929, n91930,
         n91931, n91932, n91933, n91934, n91935, n91936, n91937, n91938,
         n91939, n91940, n91941, n91942, n91943, n91944, n91945, n91946,
         n91947, n91948, n91949, n91950, n91951, n91952, n91953, n91954,
         n91955, n91956, n91957, n91958, n91959, n91960, n91961, n91962,
         n91963, n91964, n91965, n91966, n91967, n91968, n91969, n91970,
         n91971, n91972, n91973, n91974, n91975, n91976, n91977, n91978,
         n91979, n91980, n91981, n91982, n91983, n91984, n91985, n91986,
         n91987, n91988, n91989, n91990, n91991, n91992, n91993, n91994,
         n91995, n91996, n91997, n91998, n91999, n92000, n92001, n92002,
         n92003, n92004, n92005, n92006, n92007, n92008, n92009, n92010,
         n92011, n92012, n92013, n92014, n92015, n92016, n92017, n92018,
         n92019, n92020, n92021, n92022, n92023, n92024, n92025, n92026,
         n92027, n92028, n92029, n92030, n92031, n92032, n92033, n92034,
         n92035, n92036, n92037, n92038, n92039, n92040, n92041, n92042,
         n92043, n92044, n92045, n92046, n92047, n92048, n92049, n92050,
         n92051, n92052, n92053, n92054, n92055, n92056, n92057, n92058,
         n92059, n92060, n92061, n92062, n92063, n92064, n92065, n92066,
         n92067, n92068, n92069, n92070, n92071, n92072, n92073, n92074,
         n92075, n92076, n92077, n92078, n92079, n92080, n92081, n92082,
         n92083, n92084, n92085, n92086, n92087, n92088, n92089, n92090,
         n92091, n92092, n92093, n92094, n92095, n92096, n92097, n92098,
         n92099, n92100, n92101, n92102, n92103, n92104, n92105, n92106,
         n92107, n92108, n92109, n92110, n92111, n92112, n92113, n92114,
         n92115, n92116, n92117, n92118, n92119, n92120, n92121, n92122,
         n92123, n92124, n92125, n92126, n92127, n92128, n92129, n92130,
         n92131, n92132, n92133, n92134, n92135, n92136, n92137, n92138,
         n92139, n92140, n92141, n92142, n92143, n92144, n92145, n92146,
         n92147, n92148, n92149, n92150, n92151, n92152, n92153, n92154,
         n92155, n92156, n92157, n92158, n92159, n92160, n92161, n92162,
         n92163, n92164, n92165, n92166, n92167, n92168, n92169, n92170,
         n92171, n92172, n92173, n92174, n92175, n92176, n92177, n92178,
         n92179, n92180, n92181, n92182, n92183, n92184, n92185, n92186,
         n92187, n92188, n92189, n92190, n92191, n92192, n92193, n92194,
         n92195, n92196, n92197, n92198, n92199, n92200, n92201, n92202,
         n92203, n92204, n92205, n92206, n92207, n92208, n92209, n92210,
         n92211, n92212, n92213, n92214, n92215, n92216, n92217, n92218,
         n92219, n92220, n92221, n92222, n92223, n92224, n92225, n92226,
         n92227, n92228, n92229, n92230, n92231, n92232, n92233, n92234,
         n92235, n92236, n92237, n92238, n92239, n92240, n92241, n92242,
         n92243, n92244, n92245, n92246, n92247, n92248, n92249, n92250,
         n92251, n92252, n92253, n92254, n92255, n92256, n92257, n92258,
         n92259, n92260, n92261, n92262, n92263, n92264, n92265, n92266,
         n92267, n92268, n92269, n92270, n92271, n92272, n92273, n92274,
         n92275, n92276, n92277, n92278, n92279, n92280, n92281, n92282,
         n92283, n92284, n92285, n92286, n92287, n92288, n92289, n92290,
         n92291, n92292, n92293, n92294, n92295, n92296, n92297, n92298,
         n92299, n92300, n92301, n92302, n92303, n92304, n92305, n92306,
         n92307, n92308, n92309, n92310, n92311, n92312, n92313, n92314,
         n92315, n92316, n92317, n92318, n92319, n92320, n92321, n92322,
         n92323, n92324, n92325, n92326, n92327, n92328, n92329, n92330,
         n92331, n92332, n92333, n92334, n92335, n92336, n92337, n92338,
         n92339, n92340, n92341, n92342, n92343, n92344, n92345, n92346,
         n92347, n92348;

  NOR U55792 ( .A(n77753), .B(n83554), .Z(n38259) );
  XOR U55793 ( .A(n83639), .B(n38259), .Z(n38260) );
  NOR U55794 ( .A(n83549), .B(n83551), .Z(n38261) );
  IV U55795 ( .A(n38261), .Z(n38262) );
  NOR U55796 ( .A(n38260), .B(n38262), .Z(n38263) );
  NOR U55797 ( .A(n38261), .B(n83553), .Z(n38264) );
  NOR U55798 ( .A(n38263), .B(n38264), .Z(n38265) );
  IV U55799 ( .A(n38265), .Z(n83647) );
  NOR U55800 ( .A(n88227), .B(n88226), .Z(n38266) );
  NOR U55801 ( .A(n88228), .B(n38266), .Z(n38267) );
  IV U55802 ( .A(n88229), .Z(n38268) );
  NOR U55803 ( .A(n88230), .B(n38268), .Z(n38269) );
  NOR U55804 ( .A(n38269), .B(n88231), .Z(n38270) );
  XOR U55805 ( .A(n38270), .B(n38267), .Z(n38271) );
  IV U55806 ( .A(n38271), .Z(n88232) );
  NOR U55807 ( .A(n90704), .B(n90705), .Z(n38272) );
  NOR U55808 ( .A(n90706), .B(n38272), .Z(n38273) );
  IV U55809 ( .A(n38273), .Z(n90707) );
  NOR U55810 ( .A(n91765), .B(n91766), .Z(n38274) );
  NOR U55811 ( .A(n91767), .B(n38274), .Z(n38275) );
  IV U55812 ( .A(n38275), .Z(n91777) );
  NOR U55813 ( .A(n83546), .B(n83547), .Z(n38276) );
  NOR U55814 ( .A(n83548), .B(n38276), .Z(n38277) );
  IV U55815 ( .A(n38277), .Z(n89284) );
  NOR U55816 ( .A(n51450), .B(n46486), .Z(n38278) );
  NOR U55817 ( .A(n46483), .B(n51983), .Z(n38279) );
  IV U55818 ( .A(n51449), .Z(n38280) );
  IV U55819 ( .A(n38278), .Z(n38281) );
  IV U55820 ( .A(n38279), .Z(n38282) );
  IV U55821 ( .A(n51982), .Z(n38283) );
  NOR U55822 ( .A(n38283), .B(n38282), .Z(n38284) );
  NOR U55823 ( .A(n51982), .B(n38278), .Z(n38285) );
  NOR U55824 ( .A(n38281), .B(n38280), .Z(n38286) );
  NOR U55825 ( .A(n38285), .B(n38286), .Z(n38287) );
  NOR U55826 ( .A(n38279), .B(n38287), .Z(n38288) );
  NOR U55827 ( .A(n38284), .B(n38288), .Z(n51988) );
  XOR U55828 ( .A(n38289), .B(n51411), .Z(n38290) );
  NOR U55829 ( .A(n46526), .B(n56693), .Z(n38291) );
  NOR U55830 ( .A(n38291), .B(n38290), .Z(n38292) );
  NOR U55831 ( .A(n38292), .B(n46533), .Z(n38293) );
  NOR U55832 ( .A(n56690), .B(n38293), .Z(n46539) );
  IV U55833 ( .A(n51410), .Z(n38289) );
  NOR U55834 ( .A(n67216), .B(n67632), .Z(n38294) );
  NOR U55835 ( .A(n67634), .B(n38294), .Z(n38295) );
  IV U55836 ( .A(n67634), .Z(n38296) );
  IV U55837 ( .A(n62183), .Z(n38297) );
  NOR U55838 ( .A(n38296), .B(n38297), .Z(n38298) );
  NOR U55839 ( .A(n72049), .B(n38298), .Z(n38299) );
  IV U55840 ( .A(n38294), .Z(n38300) );
  NOR U55841 ( .A(n38299), .B(n38300), .Z(n38301) );
  NOR U55842 ( .A(n38295), .B(n38301), .Z(n38302) );
  IV U55843 ( .A(n38302), .Z(n67631) );
  IV U55844 ( .A(n88789), .Z(n38303) );
  NOR U55845 ( .A(n88791), .B(n88790), .Z(n38304) );
  NOR U55846 ( .A(n38303), .B(n88793), .Z(n38305) );
  NOR U55847 ( .A(n38304), .B(n38305), .Z(n38306) );
  IV U55848 ( .A(n88788), .Z(n38307) );
  IV U55849 ( .A(n88786), .Z(n38308) );
  NOR U55850 ( .A(n88787), .B(n38308), .Z(n38309) );
  NOR U55851 ( .A(n88786), .B(n88785), .Z(n38310) );
  NOR U55852 ( .A(n38310), .B(n38307), .Z(n38311) );
  NOR U55853 ( .A(n38309), .B(n38311), .Z(n38312) );
  NOR U55854 ( .A(n88782), .B(n88783), .Z(n38313) );
  NOR U55855 ( .A(n88784), .B(n38313), .Z(n38314) );
  XOR U55856 ( .A(n38312), .B(n38314), .Z(n38315) );
  NOR U55857 ( .A(n88780), .B(n88781), .Z(n38316) );
  XOR U55858 ( .A(n38306), .B(n38315), .Z(n38317) );
  XOR U55859 ( .A(n38316), .B(n38317), .Z(n89789) );
  NOR U55860 ( .A(n84192), .B(n84193), .Z(n38318) );
  NOR U55861 ( .A(n84194), .B(n38318), .Z(n38319) );
  IV U55862 ( .A(n38319), .Z(n89998) );
  XOR U55863 ( .A(n38320), .B(n77192), .Z(n38321) );
  NOR U55864 ( .A(n73017), .B(n82898), .Z(n38322) );
  NOR U55865 ( .A(n38322), .B(n38321), .Z(n38323) );
  NOR U55866 ( .A(n38323), .B(n73024), .Z(n38324) );
  NOR U55867 ( .A(n82892), .B(n38324), .Z(n38325) );
  IV U55868 ( .A(n38325), .Z(n78526) );
  IV U55869 ( .A(n77191), .Z(n38320) );
  IV U55870 ( .A(n88670), .Z(n38326) );
  NOR U55871 ( .A(n88669), .B(n88672), .Z(n38327) );
  NOR U55872 ( .A(n88673), .B(n38327), .Z(n38328) );
  NOR U55873 ( .A(n38326), .B(n88671), .Z(n38329) );
  NOR U55874 ( .A(n88674), .B(n38328), .Z(n38330) );
  IV U55875 ( .A(n38330), .Z(n38331) );
  NOR U55876 ( .A(n38329), .B(n38331), .Z(n38332) );
  IV U55877 ( .A(n88675), .Z(n38333) );
  NOR U55878 ( .A(n88678), .B(n88677), .Z(n38334) );
  NOR U55879 ( .A(n38333), .B(n88676), .Z(n38335) );
  NOR U55880 ( .A(n38334), .B(n38335), .Z(n38336) );
  XOR U55881 ( .A(n38332), .B(n38336), .Z(n88687) );
  XOR U55882 ( .A(n38337), .B(n78681), .Z(n38338) );
  NOR U55883 ( .A(n73293), .B(n78681), .Z(n38339) );
  NOR U55884 ( .A(n38339), .B(n38338), .Z(n38340) );
  NOR U55885 ( .A(n38340), .B(n82629), .Z(n38341) );
  IV U55886 ( .A(n38341), .Z(n78694) );
  IV U55887 ( .A(n78682), .Z(n38337) );
  IV U55888 ( .A(n84456), .Z(n38342) );
  NOR U55889 ( .A(n84456), .B(n84455), .Z(n38343) );
  NOR U55890 ( .A(n84454), .B(n38342), .Z(n38344) );
  NOR U55891 ( .A(n84457), .B(n38344), .Z(n38345) );
  NOR U55892 ( .A(n38343), .B(n38345), .Z(n90260) );
  NOR U55893 ( .A(n88471), .B(n88508), .Z(n38346) );
  NOR U55894 ( .A(n88466), .B(n88467), .Z(n38347) );
  NOR U55895 ( .A(n38346), .B(n38347), .Z(n38348) );
  IV U55896 ( .A(n88473), .Z(n38349) );
  NOR U55897 ( .A(n88486), .B(n88485), .Z(n38350) );
  NOR U55898 ( .A(n88483), .B(n88482), .Z(n38351) );
  NOR U55899 ( .A(n38350), .B(n38351), .Z(n38352) );
  IV U55900 ( .A(n88478), .Z(n38353) );
  IV U55901 ( .A(n88481), .Z(n38354) );
  NOR U55902 ( .A(n38354), .B(n38353), .Z(n38355) );
  NOR U55903 ( .A(n88480), .B(n38355), .Z(n38356) );
  XOR U55904 ( .A(n38356), .B(n38352), .Z(n38357) );
  NOR U55905 ( .A(n88493), .B(n88494), .Z(n38358) );
  IV U55906 ( .A(n38358), .Z(n38359) );
  NOR U55907 ( .A(n88492), .B(n38359), .Z(n38360) );
  XOR U55908 ( .A(n38357), .B(n38360), .Z(n38361) );
  NOR U55909 ( .A(n38349), .B(n88474), .Z(n38362) );
  NOR U55910 ( .A(n88475), .B(n38362), .Z(n38363) );
  XOR U55911 ( .A(n38361), .B(n38363), .Z(n38364) );
  XOR U55912 ( .A(n88472), .B(n38348), .Z(n38365) );
  XOR U55913 ( .A(n38366), .B(n38365), .Z(n90236) );
  IV U55914 ( .A(n38364), .Z(n38366) );
  NOR U55915 ( .A(n88333), .B(n88332), .Z(n38367) );
  NOR U55916 ( .A(n88334), .B(n38367), .Z(n88335) );
  IV U55917 ( .A(n88214), .Z(n38368) );
  IV U55918 ( .A(n88212), .Z(n38369) );
  NOR U55919 ( .A(n38369), .B(n88213), .Z(n38370) );
  NOR U55920 ( .A(n38368), .B(n88215), .Z(n38371) );
  NOR U55921 ( .A(n38370), .B(n38371), .Z(n38372) );
  IV U55922 ( .A(n88216), .Z(n38373) );
  IV U55923 ( .A(n88218), .Z(n38374) );
  NOR U55924 ( .A(n38374), .B(n88219), .Z(n38375) );
  NOR U55925 ( .A(n38373), .B(n88217), .Z(n38376) );
  NOR U55926 ( .A(n38375), .B(n38376), .Z(n38377) );
  IV U55927 ( .A(n88221), .Z(n38378) );
  NOR U55928 ( .A(n88222), .B(n38378), .Z(n38379) );
  IV U55929 ( .A(n88225), .Z(n38380) );
  NOR U55930 ( .A(n88220), .B(n38380), .Z(n38381) );
  NOR U55931 ( .A(n88224), .B(n38381), .Z(n38382) );
  NOR U55932 ( .A(n38379), .B(n38382), .Z(n38383) );
  XOR U55933 ( .A(n38372), .B(n38377), .Z(n38384) );
  XOR U55934 ( .A(n38383), .B(n38384), .Z(n88233) );
  NOR U55935 ( .A(n87976), .B(n87975), .Z(n38385) );
  XOR U55936 ( .A(n87965), .B(n87966), .Z(n38386) );
  XOR U55937 ( .A(n38385), .B(n38386), .Z(n38387) );
  NOR U55938 ( .A(n87954), .B(n87953), .Z(n38388) );
  XOR U55939 ( .A(n87940), .B(n87941), .Z(n38389) );
  XOR U55940 ( .A(n38388), .B(n38389), .Z(n38390) );
  IV U55941 ( .A(n87977), .Z(n38391) );
  NOR U55942 ( .A(n87978), .B(n38391), .Z(n38392) );
  XOR U55943 ( .A(n90724), .B(n90723), .Z(n38393) );
  XOR U55944 ( .A(n38392), .B(n38393), .Z(n38394) );
  NOR U55945 ( .A(n90737), .B(n90736), .Z(n38395) );
  NOR U55946 ( .A(n90732), .B(n90731), .Z(n38396) );
  XOR U55947 ( .A(n38395), .B(n38396), .Z(n38397) );
  IV U55948 ( .A(n90739), .Z(n38398) );
  IV U55949 ( .A(n90742), .Z(n38399) );
  NOR U55950 ( .A(n38399), .B(n38398), .Z(n38400) );
  NOR U55951 ( .A(n90741), .B(n38400), .Z(n38401) );
  XOR U55952 ( .A(n38401), .B(n38397), .Z(n38402) );
  XOR U55953 ( .A(n38394), .B(n38402), .Z(n38403) );
  XOR U55954 ( .A(n38387), .B(n38390), .Z(n38404) );
  XOR U55955 ( .A(n38403), .B(n38404), .Z(n38405) );
  IV U55956 ( .A(n38405), .Z(n90743) );
  NOR U55957 ( .A(n48144), .B(n49953), .Z(n38406) );
  NOR U55958 ( .A(n53325), .B(n48145), .Z(n38407) );
  IV U55959 ( .A(n38406), .Z(n38408) );
  IV U55960 ( .A(n38407), .Z(n38409) );
  IV U55961 ( .A(n49952), .Z(n38410) );
  NOR U55962 ( .A(n38410), .B(n38408), .Z(n38411) );
  NOR U55963 ( .A(n48146), .B(n38409), .Z(n38412) );
  NOR U55964 ( .A(n49952), .B(n38407), .Z(n38413) );
  NOR U55965 ( .A(n38412), .B(n38413), .Z(n38414) );
  NOR U55966 ( .A(n38406), .B(n38414), .Z(n38415) );
  NOR U55967 ( .A(n38411), .B(n38415), .Z(n53339) );
  IV U55968 ( .A(n87652), .Z(n38416) );
  NOR U55969 ( .A(n87655), .B(n87654), .Z(n38417) );
  NOR U55970 ( .A(n38416), .B(n87653), .Z(n38418) );
  NOR U55971 ( .A(n38417), .B(n38418), .Z(n38419) );
  IV U55972 ( .A(n87657), .Z(n38420) );
  IV U55973 ( .A(n87660), .Z(n38421) );
  NOR U55974 ( .A(n38420), .B(n38421), .Z(n38422) );
  NOR U55975 ( .A(n87659), .B(n38422), .Z(n38423) );
  XOR U55976 ( .A(n87671), .B(n90893), .Z(n38424) );
  XOR U55977 ( .A(n90892), .B(n38424), .Z(n38425) );
  IV U55978 ( .A(n90910), .Z(n38426) );
  NOR U55979 ( .A(n90922), .B(n90921), .Z(n38427) );
  NOR U55980 ( .A(n90915), .B(n90914), .Z(n38428) );
  XOR U55981 ( .A(n38427), .B(n38428), .Z(n38429) );
  NOR U55982 ( .A(n90905), .B(n90904), .Z(n38430) );
  NOR U55983 ( .A(n38430), .B(n38426), .Z(n38431) );
  XOR U55984 ( .A(n38429), .B(n38431), .Z(n38432) );
  XOR U55985 ( .A(n38425), .B(n38432), .Z(n38433) );
  XOR U55986 ( .A(n38423), .B(n87672), .Z(n38434) );
  XOR U55987 ( .A(n38433), .B(n38434), .Z(n38435) );
  XOR U55988 ( .A(n38419), .B(n38435), .Z(n38436) );
  IV U55989 ( .A(n38436), .Z(n90923) );
  NOR U55990 ( .A(n85276), .B(n85277), .Z(n38437) );
  NOR U55991 ( .A(n85278), .B(n38437), .Z(n38438) );
  IV U55992 ( .A(n38438), .Z(n87595) );
  NOR U55993 ( .A(n76083), .B(n76084), .Z(n38439) );
  NOR U55994 ( .A(n76085), .B(n38439), .Z(n38440) );
  IV U55995 ( .A(n38440), .Z(n85529) );
  NOR U55996 ( .A(n75971), .B(n75968), .Z(n38441) );
  IV U55997 ( .A(n74469), .Z(n38442) );
  IV U55998 ( .A(n75970), .Z(n38443) );
  IV U55999 ( .A(n38441), .Z(n38444) );
  NOR U56000 ( .A(n75970), .B(n38441), .Z(n38445) );
  NOR U56001 ( .A(n38443), .B(n38442), .Z(n38446) );
  NOR U56002 ( .A(n85620), .B(n38446), .Z(n38447) );
  NOR U56003 ( .A(n38447), .B(n38444), .Z(n38448) );
  NOR U56004 ( .A(n38445), .B(n38448), .Z(n38449) );
  IV U56005 ( .A(n38449), .Z(n75964) );
  NOR U56006 ( .A(n87271), .B(n87270), .Z(n38450) );
  NOR U56007 ( .A(n87272), .B(n38450), .Z(n38451) );
  IV U56008 ( .A(n87274), .Z(n38452) );
  NOR U56009 ( .A(n87275), .B(n38452), .Z(n38453) );
  NOR U56010 ( .A(n87276), .B(n87273), .Z(n38454) );
  NOR U56011 ( .A(n87277), .B(n38454), .Z(n38455) );
  NOR U56012 ( .A(n38453), .B(n38455), .Z(n38456) );
  NOR U56013 ( .A(n87268), .B(n87269), .Z(n38457) );
  NOR U56014 ( .A(n38451), .B(n38457), .Z(n38458) );
  XOR U56015 ( .A(n38456), .B(n38458), .Z(n87285) );
  NOR U56016 ( .A(n85892), .B(n85893), .Z(n38459) );
  NOR U56017 ( .A(n85894), .B(n38459), .Z(n38460) );
  IV U56018 ( .A(n38460), .Z(n85896) );
  IV U56019 ( .A(n86886), .Z(n38461) );
  NOR U56020 ( .A(n86888), .B(n86887), .Z(n38462) );
  NOR U56021 ( .A(n38462), .B(n38461), .Z(n38463) );
  NOR U56022 ( .A(n86889), .B(n86890), .Z(n38464) );
  NOR U56023 ( .A(n86891), .B(n38464), .Z(n38465) );
  NOR U56024 ( .A(n38463), .B(n38465), .Z(n86901) );
  IV U56025 ( .A(n86658), .Z(n38466) );
  NOR U56026 ( .A(n86658), .B(n86657), .Z(n38467) );
  NOR U56027 ( .A(n86656), .B(n38466), .Z(n38468) );
  NOR U56028 ( .A(n86659), .B(n38468), .Z(n38469) );
  NOR U56029 ( .A(n38467), .B(n38469), .Z(n38470) );
  NOR U56030 ( .A(n86654), .B(n86653), .Z(n38471) );
  NOR U56031 ( .A(n86655), .B(n38471), .Z(n38472) );
  XOR U56032 ( .A(n38470), .B(n38472), .Z(n38473) );
  IV U56033 ( .A(n86650), .Z(n38474) );
  NOR U56034 ( .A(n91855), .B(n91854), .Z(n38475) );
  XOR U56035 ( .A(n91846), .B(n91847), .Z(n38476) );
  XOR U56036 ( .A(n38475), .B(n38476), .Z(n38477) );
  NOR U56037 ( .A(n38474), .B(n86651), .Z(n38478) );
  NOR U56038 ( .A(n86652), .B(n38478), .Z(n38479) );
  XOR U56039 ( .A(n38477), .B(n38479), .Z(n38480) );
  XOR U56040 ( .A(n38473), .B(n38480), .Z(n91856) );
  IV U56041 ( .A(n86505), .Z(n38481) );
  NOR U56042 ( .A(n86512), .B(n86511), .Z(n38482) );
  NOR U56043 ( .A(n86509), .B(n86508), .Z(n38483) );
  NOR U56044 ( .A(n38482), .B(n38483), .Z(n38484) );
  IV U56045 ( .A(n38484), .Z(n38485) );
  IV U56046 ( .A(n86501), .Z(n38486) );
  IV U56047 ( .A(n86503), .Z(n38487) );
  NOR U56048 ( .A(n38487), .B(n86504), .Z(n38488) );
  NOR U56049 ( .A(n38486), .B(n86502), .Z(n38489) );
  NOR U56050 ( .A(n38488), .B(n38489), .Z(n38490) );
  NOR U56051 ( .A(n38481), .B(n86506), .Z(n38491) );
  NOR U56052 ( .A(n38491), .B(n38485), .Z(n38492) );
  XOR U56053 ( .A(n38490), .B(n38492), .Z(n38493) );
  IV U56054 ( .A(n86516), .Z(n38494) );
  NOR U56055 ( .A(n86513), .B(n38494), .Z(n38495) );
  NOR U56056 ( .A(n86515), .B(n38495), .Z(n38496) );
  NOR U56057 ( .A(n86517), .B(n38496), .Z(n38497) );
  XOR U56058 ( .A(n38493), .B(n38497), .Z(n86552) );
  IV U56059 ( .A(x[1599]), .Z(n38498) );
  XOR U56060 ( .A(n38498), .B(y[1599]), .Z(n92272) );
  XOR U56061 ( .A(x[1598]), .B(y[1598]), .Z(n92217) );
  XOR U56062 ( .A(x[1597]), .B(y[1597]), .Z(n92184) );
  XOR U56063 ( .A(x[1596]), .B(y[1596]), .Z(n92157) );
  XOR U56064 ( .A(x[1595]), .B(y[1595]), .Z(n92147) );
  XOR U56065 ( .A(x[1594]), .B(y[1594]), .Z(n92122) );
  XOR U56066 ( .A(x[1593]), .B(y[1593]), .Z(n86392) );
  XOR U56067 ( .A(x[1592]), .B(y[1592]), .Z(n86364) );
  XOR U56068 ( .A(x[1591]), .B(y[1591]), .Z(n80655) );
  XOR U56069 ( .A(x[1590]), .B(y[1590]), .Z(n75320) );
  XOR U56070 ( .A(x[1589]), .B(y[1589]), .Z(n70018) );
  XOR U56071 ( .A(x[1588]), .B(y[1588]), .Z(n64859) );
  XOR U56072 ( .A(x[1587]), .B(y[1587]), .Z(n64842) );
  XOR U56073 ( .A(x[1586]), .B(y[1586]), .Z(n38499) );
  IV U56074 ( .A(n38499), .Z(n59649) );
  IV U56075 ( .A(x[1585]), .Z(n38500) );
  XOR U56076 ( .A(n38500), .B(y[1585]), .Z(n59626) );
  XOR U56077 ( .A(x[1584]), .B(y[1584]), .Z(n59617) );
  XOR U56078 ( .A(x[1583]), .B(y[1583]), .Z(n59604) );
  XOR U56079 ( .A(x[1582]), .B(y[1582]), .Z(n38501) );
  IV U56080 ( .A(n38501), .Z(n59581) );
  IV U56081 ( .A(x[1581]), .Z(n38502) );
  XOR U56082 ( .A(n38502), .B(y[1581]), .Z(n59565) );
  XOR U56083 ( .A(x[1580]), .B(y[1580]), .Z(n59561) );
  XOR U56084 ( .A(x[1579]), .B(y[1579]), .Z(n54253) );
  XOR U56085 ( .A(x[1578]), .B(y[1578]), .Z(n38503) );
  IV U56086 ( .A(n38503), .Z(n54246) );
  IV U56087 ( .A(x[1577]), .Z(n38504) );
  XOR U56088 ( .A(n38504), .B(y[1577]), .Z(n49126) );
  XOR U56089 ( .A(x[1576]), .B(y[1576]), .Z(n44380) );
  XOR U56090 ( .A(x[1575]), .B(y[1575]), .Z(n44384) );
  XOR U56091 ( .A(x[1574]), .B(y[1574]), .Z(n38505) );
  IV U56092 ( .A(n38505), .Z(n44378) );
  IV U56093 ( .A(x[1573]), .Z(n38506) );
  XOR U56094 ( .A(n38506), .B(y[1573]), .Z(n44375) );
  XOR U56095 ( .A(x[1572]), .B(y[1572]), .Z(n44370) );
  XOR U56096 ( .A(x[1571]), .B(y[1571]), .Z(n44367) );
  XOR U56097 ( .A(x[1570]), .B(y[1570]), .Z(n38507) );
  IV U56098 ( .A(n38507), .Z(n44365) );
  IV U56099 ( .A(x[1569]), .Z(n38508) );
  XOR U56100 ( .A(n38508), .B(y[1569]), .Z(n44362) );
  XOR U56101 ( .A(x[1568]), .B(y[1568]), .Z(n38645) );
  XOR U56102 ( .A(x[1567]), .B(y[1567]), .Z(n44357) );
  XOR U56103 ( .A(x[1566]), .B(y[1566]), .Z(n38509) );
  IV U56104 ( .A(n38509), .Z(n44355) );
  IV U56105 ( .A(x[1565]), .Z(n38510) );
  XOR U56106 ( .A(n38510), .B(y[1565]), .Z(n38651) );
  XOR U56107 ( .A(x[1564]), .B(y[1564]), .Z(n38648) );
  XOR U56108 ( .A(x[1563]), .B(y[1563]), .Z(n38656) );
  XOR U56109 ( .A(x[1562]), .B(y[1562]), .Z(n38511) );
  IV U56110 ( .A(n38511), .Z(n38654) );
  IV U56111 ( .A(x[1561]), .Z(n38512) );
  XOR U56112 ( .A(n38512), .B(y[1561]), .Z(n38660) );
  XOR U56113 ( .A(x[1560]), .B(y[1560]), .Z(n44350) );
  XOR U56114 ( .A(x[1559]), .B(y[1559]), .Z(n44347) );
  XOR U56115 ( .A(x[1558]), .B(y[1558]), .Z(n38513) );
  IV U56116 ( .A(n38513), .Z(n38665) );
  IV U56117 ( .A(x[1557]), .Z(n38514) );
  XOR U56118 ( .A(n38514), .B(y[1557]), .Z(n38663) );
  XOR U56119 ( .A(x[1556]), .B(y[1556]), .Z(n44341) );
  XOR U56120 ( .A(x[1555]), .B(y[1555]), .Z(n44338) );
  XOR U56121 ( .A(x[1554]), .B(y[1554]), .Z(n38515) );
  IV U56122 ( .A(n38515), .Z(n38670) );
  IV U56123 ( .A(x[1553]), .Z(n38516) );
  XOR U56124 ( .A(n38516), .B(y[1553]), .Z(n38668) );
  XOR U56125 ( .A(x[1552]), .B(y[1552]), .Z(n38675) );
  XOR U56126 ( .A(x[1551]), .B(y[1551]), .Z(n38672) );
  XOR U56127 ( .A(x[1550]), .B(y[1550]), .Z(n38517) );
  IV U56128 ( .A(n38517), .Z(n44335) );
  IV U56129 ( .A(x[1549]), .Z(n38518) );
  XOR U56130 ( .A(n38518), .B(y[1549]), .Z(n44333) );
  XOR U56131 ( .A(x[1548]), .B(y[1548]), .Z(n44328) );
  XOR U56132 ( .A(x[1547]), .B(y[1547]), .Z(n44325) );
  XOR U56133 ( .A(x[1546]), .B(y[1546]), .Z(n38681) );
  XOR U56134 ( .A(x[1545]), .B(y[1545]), .Z(n38678) );
  XOR U56135 ( .A(x[1544]), .B(y[1544]), .Z(n38684) );
  XOR U56136 ( .A(x[1543]), .B(y[1543]), .Z(n44319) );
  XOR U56137 ( .A(x[1542]), .B(y[1542]), .Z(n44316) );
  XOR U56138 ( .A(x[1541]), .B(y[1541]), .Z(n38519) );
  IV U56139 ( .A(n38519), .Z(n38691) );
  IV U56140 ( .A(x[1540]), .Z(n38520) );
  XOR U56141 ( .A(n38520), .B(y[1540]), .Z(n38687) );
  XOR U56142 ( .A(x[1539]), .B(y[1539]), .Z(n44311) );
  XOR U56143 ( .A(x[1538]), .B(y[1538]), .Z(n44308) );
  XOR U56144 ( .A(x[1537]), .B(y[1537]), .Z(n44304) );
  XOR U56145 ( .A(x[1536]), .B(y[1536]), .Z(n44301) );
  XOR U56146 ( .A(x[1535]), .B(y[1535]), .Z(n44297) );
  XOR U56147 ( .A(x[1534]), .B(y[1534]), .Z(n44294) );
  XOR U56148 ( .A(x[1533]), .B(y[1533]), .Z(n38695) );
  XOR U56149 ( .A(x[1532]), .B(y[1532]), .Z(n38692) );
  XOR U56150 ( .A(x[1531]), .B(y[1531]), .Z(n38701) );
  XOR U56151 ( .A(x[1530]), .B(y[1530]), .Z(n38698) );
  XOR U56152 ( .A(x[1529]), .B(y[1529]), .Z(n38707) );
  XOR U56153 ( .A(x[1528]), .B(y[1528]), .Z(n38704) );
  XOR U56154 ( .A(x[1527]), .B(y[1527]), .Z(n44290) );
  XOR U56155 ( .A(x[1526]), .B(y[1526]), .Z(n44287) );
  XOR U56156 ( .A(x[1525]), .B(y[1525]), .Z(n38713) );
  XOR U56157 ( .A(x[1524]), .B(y[1524]), .Z(n38710) );
  XOR U56158 ( .A(x[1523]), .B(y[1523]), .Z(n38719) );
  XOR U56159 ( .A(x[1522]), .B(y[1522]), .Z(n38716) );
  XOR U56160 ( .A(x[1521]), .B(y[1521]), .Z(n38521) );
  IV U56161 ( .A(n38521), .Z(n44283) );
  IV U56162 ( .A(x[1520]), .Z(n38522) );
  XOR U56163 ( .A(n38522), .B(y[1520]), .Z(n44280) );
  XOR U56164 ( .A(x[1519]), .B(y[1519]), .Z(n38523) );
  IV U56165 ( .A(n38523), .Z(n38724) );
  IV U56166 ( .A(x[1518]), .Z(n38524) );
  XOR U56167 ( .A(n38524), .B(y[1518]), .Z(n44273) );
  XOR U56168 ( .A(x[1517]), .B(y[1517]), .Z(n38725) );
  XOR U56169 ( .A(x[1516]), .B(y[1516]), .Z(n44260) );
  XOR U56170 ( .A(x[1515]), .B(y[1515]), .Z(n44256) );
  XOR U56171 ( .A(x[1514]), .B(y[1514]), .Z(n44263) );
  XOR U56172 ( .A(x[1513]), .B(y[1513]), .Z(n44251) );
  XOR U56173 ( .A(x[1512]), .B(y[1512]), .Z(n44248) );
  XOR U56174 ( .A(x[1511]), .B(y[1511]), .Z(n38728) );
  XOR U56175 ( .A(x[1510]), .B(y[1510]), .Z(n38735) );
  XOR U56176 ( .A(x[1509]), .B(y[1509]), .Z(n38732) );
  XOR U56177 ( .A(x[1508]), .B(y[1508]), .Z(n44245) );
  XOR U56178 ( .A(x[1507]), .B(y[1507]), .Z(n44459) );
  XOR U56179 ( .A(x[1506]), .B(y[1506]), .Z(n44234) );
  XOR U56180 ( .A(x[1505]), .B(y[1505]), .Z(n38738) );
  XOR U56181 ( .A(x[1504]), .B(y[1504]), .Z(n38744) );
  XOR U56182 ( .A(x[1503]), .B(y[1503]), .Z(n38741) );
  XOR U56183 ( .A(x[1502]), .B(y[1502]), .Z(n44228) );
  XOR U56184 ( .A(x[1501]), .B(y[1501]), .Z(n44225) );
  XOR U56185 ( .A(x[1500]), .B(y[1500]), .Z(n38750) );
  XOR U56186 ( .A(x[1499]), .B(y[1499]), .Z(n38747) );
  XOR U56187 ( .A(x[1498]), .B(y[1498]), .Z(n44222) );
  XOR U56188 ( .A(x[1497]), .B(y[1497]), .Z(n44219) );
  XOR U56189 ( .A(x[1496]), .B(y[1496]), .Z(n44216) );
  XOR U56190 ( .A(x[1495]), .B(y[1495]), .Z(n44213) );
  XOR U56191 ( .A(x[1494]), .B(y[1494]), .Z(n44209) );
  XOR U56192 ( .A(x[1493]), .B(y[1493]), .Z(n44206) );
  XOR U56193 ( .A(x[1492]), .B(y[1492]), .Z(n38753) );
  XOR U56194 ( .A(x[1491]), .B(y[1491]), .Z(n44202) );
  XOR U56195 ( .A(x[1490]), .B(y[1490]), .Z(n44199) );
  XOR U56196 ( .A(x[1489]), .B(y[1489]), .Z(n44195) );
  XOR U56197 ( .A(x[1488]), .B(y[1488]), .Z(n44192) );
  XOR U56198 ( .A(x[1487]), .B(y[1487]), .Z(n38756) );
  XOR U56199 ( .A(x[1486]), .B(y[1486]), .Z(n44188) );
  XOR U56200 ( .A(x[1485]), .B(y[1485]), .Z(n44185) );
  XOR U56201 ( .A(x[1484]), .B(y[1484]), .Z(n44181) );
  XOR U56202 ( .A(x[1483]), .B(y[1483]), .Z(n44178) );
  XOR U56203 ( .A(x[1482]), .B(y[1482]), .Z(n38759) );
  XOR U56204 ( .A(x[1481]), .B(y[1481]), .Z(n44164) );
  XOR U56205 ( .A(x[1480]), .B(y[1480]), .Z(n44161) );
  XOR U56206 ( .A(x[1479]), .B(y[1479]), .Z(n38762) );
  XOR U56207 ( .A(x[1478]), .B(y[1478]), .Z(n44157) );
  XOR U56208 ( .A(x[1477]), .B(y[1477]), .Z(n44154) );
  XOR U56209 ( .A(x[1476]), .B(y[1476]), .Z(n44150) );
  XOR U56210 ( .A(x[1475]), .B(y[1475]), .Z(n44147) );
  XOR U56211 ( .A(x[1474]), .B(y[1474]), .Z(n38765) );
  XOR U56212 ( .A(x[1473]), .B(y[1473]), .Z(n44140) );
  XOR U56213 ( .A(x[1472]), .B(y[1472]), .Z(n38768) );
  XOR U56214 ( .A(x[1471]), .B(y[1471]), .Z(n38774) );
  XOR U56215 ( .A(x[1470]), .B(y[1470]), .Z(n38771) );
  XOR U56216 ( .A(x[1469]), .B(y[1469]), .Z(n38780) );
  XOR U56217 ( .A(x[1468]), .B(y[1468]), .Z(n38777) );
  XOR U56218 ( .A(x[1467]), .B(y[1467]), .Z(n38783) );
  XOR U56219 ( .A(x[1466]), .B(y[1466]), .Z(n44133) );
  XOR U56220 ( .A(x[1465]), .B(y[1465]), .Z(n44130) );
  XOR U56221 ( .A(x[1464]), .B(y[1464]), .Z(n38789) );
  XOR U56222 ( .A(x[1463]), .B(y[1463]), .Z(n38786) );
  XOR U56223 ( .A(x[1462]), .B(y[1462]), .Z(n44127) );
  XOR U56224 ( .A(x[1461]), .B(y[1461]), .Z(n44124) );
  XOR U56225 ( .A(x[1460]), .B(y[1460]), .Z(n38795) );
  XOR U56226 ( .A(x[1459]), .B(y[1459]), .Z(n38792) );
  XOR U56227 ( .A(x[1458]), .B(y[1458]), .Z(n38799) );
  XOR U56228 ( .A(x[1457]), .B(y[1457]), .Z(n44120) );
  XOR U56229 ( .A(x[1456]), .B(y[1456]), .Z(n44117) );
  XOR U56230 ( .A(x[1455]), .B(y[1455]), .Z(n38805) );
  XOR U56231 ( .A(x[1454]), .B(y[1454]), .Z(n38802) );
  XOR U56232 ( .A(x[1453]), .B(y[1453]), .Z(n44113) );
  XOR U56233 ( .A(x[1452]), .B(y[1452]), .Z(n44110) );
  XOR U56234 ( .A(x[1451]), .B(y[1451]), .Z(n38811) );
  XOR U56235 ( .A(x[1450]), .B(y[1450]), .Z(n38808) );
  XOR U56236 ( .A(x[1449]), .B(y[1449]), .Z(n38814) );
  XOR U56237 ( .A(x[1448]), .B(y[1448]), .Z(n44096) );
  XOR U56238 ( .A(x[1447]), .B(y[1447]), .Z(n44093) );
  XOR U56239 ( .A(x[1446]), .B(y[1446]), .Z(n44089) );
  XOR U56240 ( .A(x[1445]), .B(y[1445]), .Z(n44086) );
  XOR U56241 ( .A(x[1444]), .B(y[1444]), .Z(n44075) );
  XOR U56242 ( .A(x[1443]), .B(y[1443]), .Z(n38817) );
  XOR U56243 ( .A(x[1442]), .B(y[1442]), .Z(n44078) );
  XOR U56244 ( .A(x[1441]), .B(y[1441]), .Z(n38823) );
  XOR U56245 ( .A(x[1440]), .B(y[1440]), .Z(n38820) );
  XOR U56246 ( .A(x[1439]), .B(y[1439]), .Z(n38829) );
  XOR U56247 ( .A(x[1438]), .B(y[1438]), .Z(n38826) );
  XOR U56248 ( .A(x[1437]), .B(y[1437]), .Z(n38832) );
  XOR U56249 ( .A(x[1436]), .B(y[1436]), .Z(n38839) );
  XOR U56250 ( .A(x[1435]), .B(y[1435]), .Z(n38838) );
  XOR U56251 ( .A(x[1434]), .B(y[1434]), .Z(n38845) );
  XOR U56252 ( .A(x[1433]), .B(y[1433]), .Z(n38842) );
  XOR U56253 ( .A(x[1432]), .B(y[1432]), .Z(n38848) );
  XOR U56254 ( .A(x[1431]), .B(y[1431]), .Z(n44068) );
  XOR U56255 ( .A(x[1430]), .B(y[1430]), .Z(n44065) );
  XOR U56256 ( .A(x[1429]), .B(y[1429]), .Z(n38854) );
  XOR U56257 ( .A(x[1428]), .B(y[1428]), .Z(n38851) );
  XOR U56258 ( .A(x[1427]), .B(y[1427]), .Z(n38860) );
  XOR U56259 ( .A(x[1426]), .B(y[1426]), .Z(n38857) );
  XOR U56260 ( .A(x[1425]), .B(y[1425]), .Z(n38866) );
  XOR U56261 ( .A(x[1424]), .B(y[1424]), .Z(n38863) );
  XOR U56262 ( .A(x[1423]), .B(y[1423]), .Z(n38869) );
  XOR U56263 ( .A(x[1422]), .B(y[1422]), .Z(n44057) );
  XOR U56264 ( .A(x[1421]), .B(y[1421]), .Z(n38872) );
  XOR U56265 ( .A(x[1420]), .B(y[1420]), .Z(n44050) );
  XOR U56266 ( .A(x[1419]), .B(y[1419]), .Z(n44047) );
  XOR U56267 ( .A(x[1418]), .B(y[1418]), .Z(n48838) );
  XOR U56268 ( .A(x[1417]), .B(y[1417]), .Z(n44041) );
  XOR U56269 ( .A(x[1416]), .B(y[1416]), .Z(n38878) );
  XOR U56270 ( .A(x[1415]), .B(y[1415]), .Z(n38875) );
  XOR U56271 ( .A(x[1414]), .B(y[1414]), .Z(n44035) );
  XOR U56272 ( .A(x[1413]), .B(y[1413]), .Z(n44032) );
  XOR U56273 ( .A(x[1412]), .B(y[1412]), .Z(n48827) );
  XOR U56274 ( .A(x[1411]), .B(y[1411]), .Z(n44027) );
  IV U56275 ( .A(n44027), .Z(n48814) );
  XOR U56276 ( .A(x[1410]), .B(y[1410]), .Z(n38881) );
  XOR U56277 ( .A(x[1409]), .B(y[1409]), .Z(n38887) );
  XOR U56278 ( .A(x[1408]), .B(y[1408]), .Z(n38884) );
  XOR U56279 ( .A(x[1407]), .B(y[1407]), .Z(n44024) );
  XOR U56280 ( .A(x[1406]), .B(y[1406]), .Z(n44021) );
  XOR U56281 ( .A(x[1405]), .B(y[1405]), .Z(n44018) );
  XOR U56282 ( .A(x[1404]), .B(y[1404]), .Z(n44015) );
  XOR U56283 ( .A(x[1403]), .B(y[1403]), .Z(n44011) );
  XOR U56284 ( .A(x[1402]), .B(y[1402]), .Z(n44008) );
  XOR U56285 ( .A(x[1401]), .B(y[1401]), .Z(n38890) );
  XOR U56286 ( .A(x[1400]), .B(y[1400]), .Z(n43997) );
  XOR U56287 ( .A(x[1399]), .B(y[1399]), .Z(n43991) );
  XOR U56288 ( .A(x[1398]), .B(y[1398]), .Z(n43988) );
  XOR U56289 ( .A(x[1397]), .B(y[1397]), .Z(n43984) );
  XOR U56290 ( .A(x[1396]), .B(y[1396]), .Z(n43981) );
  XOR U56291 ( .A(x[1395]), .B(y[1395]), .Z(n43977) );
  XOR U56292 ( .A(x[1394]), .B(y[1394]), .Z(n43974) );
  XOR U56293 ( .A(x[1393]), .B(y[1393]), .Z(n43971) );
  XOR U56294 ( .A(x[1392]), .B(y[1392]), .Z(n43968) );
  XOR U56295 ( .A(x[1391]), .B(y[1391]), .Z(n43964) );
  XOR U56296 ( .A(x[1390]), .B(y[1390]), .Z(n43961) );
  XOR U56297 ( .A(x[1389]), .B(y[1389]), .Z(n38893) );
  XOR U56298 ( .A(x[1388]), .B(y[1388]), .Z(n43958) );
  XOR U56299 ( .A(x[1387]), .B(y[1387]), .Z(n43955) );
  XOR U56300 ( .A(x[1386]), .B(y[1386]), .Z(n48789) );
  XOR U56301 ( .A(x[1385]), .B(y[1385]), .Z(n43949) );
  XOR U56302 ( .A(x[1384]), .B(y[1384]), .Z(n43944) );
  XOR U56303 ( .A(x[1383]), .B(y[1383]), .Z(n43941) );
  XOR U56304 ( .A(x[1382]), .B(y[1382]), .Z(n38900) );
  XOR U56305 ( .A(x[1381]), .B(y[1381]), .Z(n38897) );
  XOR U56306 ( .A(x[1380]), .B(y[1380]), .Z(n59205) );
  XOR U56307 ( .A(x[1379]), .B(y[1379]), .Z(n38903) );
  IV U56308 ( .A(n38903), .Z(n38906) );
  XOR U56309 ( .A(x[1378]), .B(y[1378]), .Z(n38910) );
  IV U56310 ( .A(n38910), .Z(n48765) );
  XOR U56311 ( .A(x[1377]), .B(y[1377]), .Z(n38912) );
  XOR U56312 ( .A(x[1376]), .B(y[1376]), .Z(n43936) );
  XOR U56313 ( .A(x[1375]), .B(y[1375]), .Z(n43933) );
  XOR U56314 ( .A(x[1374]), .B(y[1374]), .Z(n43929) );
  XOR U56315 ( .A(x[1373]), .B(y[1373]), .Z(n43926) );
  XOR U56316 ( .A(x[1372]), .B(y[1372]), .Z(n43921) );
  XOR U56317 ( .A(x[1371]), .B(y[1371]), .Z(n43918) );
  XOR U56318 ( .A(x[1370]), .B(y[1370]), .Z(n38916) );
  XOR U56319 ( .A(x[1369]), .B(y[1369]), .Z(n38922) );
  XOR U56320 ( .A(x[1368]), .B(y[1368]), .Z(n38525) );
  IV U56321 ( .A(n38525), .Z(n38921) );
  IV U56322 ( .A(x[1367]), .Z(n38526) );
  XOR U56323 ( .A(n38526), .B(y[1367]), .Z(n43904) );
  XOR U56324 ( .A(x[1366]), .B(y[1366]), .Z(n38925) );
  XOR U56325 ( .A(x[1365]), .B(y[1365]), .Z(n43905) );
  XOR U56326 ( .A(x[1364]), .B(y[1364]), .Z(n38931) );
  XOR U56327 ( .A(x[1363]), .B(y[1363]), .Z(n38928) );
  XOR U56328 ( .A(x[1362]), .B(y[1362]), .Z(n38937) );
  XOR U56329 ( .A(x[1361]), .B(y[1361]), .Z(n38934) );
  XOR U56330 ( .A(x[1360]), .B(y[1360]), .Z(n43895) );
  XOR U56331 ( .A(x[1359]), .B(y[1359]), .Z(n43892) );
  XOR U56332 ( .A(x[1358]), .B(y[1358]), .Z(n38943) );
  XOR U56333 ( .A(x[1357]), .B(y[1357]), .Z(n38940) );
  XOR U56334 ( .A(x[1356]), .B(y[1356]), .Z(n43888) );
  XOR U56335 ( .A(x[1355]), .B(y[1355]), .Z(n43885) );
  XOR U56336 ( .A(x[1354]), .B(y[1354]), .Z(n43881) );
  XOR U56337 ( .A(x[1353]), .B(y[1353]), .Z(n43878) );
  XOR U56338 ( .A(x[1352]), .B(y[1352]), .Z(n43874) );
  XOR U56339 ( .A(x[1351]), .B(y[1351]), .Z(n43871) );
  XOR U56340 ( .A(x[1350]), .B(y[1350]), .Z(n43867) );
  XOR U56341 ( .A(x[1349]), .B(y[1349]), .Z(n43864) );
  XOR U56342 ( .A(x[1346]), .B(y[1346]), .Z(n38949) );
  XOR U56343 ( .A(x[1345]), .B(y[1345]), .Z(n38946) );
  XOR U56344 ( .A(x[1344]), .B(y[1344]), .Z(n38955) );
  XOR U56345 ( .A(x[1343]), .B(y[1343]), .Z(n38952) );
  XOR U56346 ( .A(x[1342]), .B(y[1342]), .Z(n38961) );
  XOR U56347 ( .A(x[1341]), .B(y[1341]), .Z(n38958) );
  XOR U56348 ( .A(x[1340]), .B(y[1340]), .Z(n38967) );
  XOR U56349 ( .A(x[1339]), .B(y[1339]), .Z(n38964) );
  XOR U56350 ( .A(x[1338]), .B(y[1338]), .Z(n38970) );
  XOR U56351 ( .A(x[1337]), .B(y[1337]), .Z(n43852) );
  XOR U56352 ( .A(x[1336]), .B(y[1336]), .Z(n43849) );
  XOR U56353 ( .A(x[1335]), .B(y[1335]), .Z(n43845) );
  XOR U56354 ( .A(x[1334]), .B(y[1334]), .Z(n43842) );
  XOR U56355 ( .A(x[1333]), .B(y[1333]), .Z(n38973) );
  XOR U56356 ( .A(x[1332]), .B(y[1332]), .Z(n43834) );
  XOR U56357 ( .A(x[1331]), .B(y[1331]), .Z(n43831) );
  XOR U56358 ( .A(x[1330]), .B(y[1330]), .Z(n43826) );
  XOR U56359 ( .A(x[1329]), .B(y[1329]), .Z(n43823) );
  XOR U56360 ( .A(x[1328]), .B(y[1328]), .Z(n38976) );
  XOR U56361 ( .A(x[1327]), .B(y[1327]), .Z(n38982) );
  XOR U56362 ( .A(x[1326]), .B(y[1326]), .Z(n38979) );
  XOR U56363 ( .A(x[1325]), .B(y[1325]), .Z(n43818) );
  XOR U56364 ( .A(x[1324]), .B(y[1324]), .Z(n43815) );
  XOR U56365 ( .A(x[1323]), .B(y[1323]), .Z(n38988) );
  XOR U56366 ( .A(x[1322]), .B(y[1322]), .Z(n38985) );
  XOR U56367 ( .A(x[1321]), .B(y[1321]), .Z(n43811) );
  XOR U56368 ( .A(x[1320]), .B(y[1320]), .Z(n43808) );
  XOR U56369 ( .A(x[1319]), .B(y[1319]), .Z(n43805) );
  XOR U56370 ( .A(x[1318]), .B(y[1318]), .Z(n43802) );
  XOR U56371 ( .A(x[1317]), .B(y[1317]), .Z(n43798) );
  XOR U56372 ( .A(x[1316]), .B(y[1316]), .Z(n43795) );
  XOR U56373 ( .A(x[1315]), .B(y[1315]), .Z(n38991) );
  XOR U56374 ( .A(x[1314]), .B(y[1314]), .Z(n44665) );
  XOR U56375 ( .A(x[1313]), .B(y[1313]), .Z(n48598) );
  XOR U56376 ( .A(x[1312]), .B(y[1312]), .Z(n38994) );
  XOR U56377 ( .A(x[1311]), .B(y[1311]), .Z(n43787) );
  XOR U56378 ( .A(x[1310]), .B(y[1310]), .Z(n43784) );
  XOR U56379 ( .A(x[1309]), .B(y[1309]), .Z(n43780) );
  XOR U56380 ( .A(x[1308]), .B(y[1308]), .Z(n43778) );
  IV U56381 ( .A(n43778), .Z(n43776) );
  XOR U56382 ( .A(x[1307]), .B(y[1307]), .Z(n38997) );
  XOR U56383 ( .A(x[1306]), .B(y[1306]), .Z(n39003) );
  XOR U56384 ( .A(x[1305]), .B(y[1305]), .Z(n39000) );
  XOR U56385 ( .A(x[1304]), .B(y[1304]), .Z(n39009) );
  XOR U56386 ( .A(x[1303]), .B(y[1303]), .Z(n39006) );
  XOR U56387 ( .A(x[1302]), .B(y[1302]), .Z(n39015) );
  XOR U56388 ( .A(x[1301]), .B(y[1301]), .Z(n39012) );
  XOR U56389 ( .A(x[1300]), .B(y[1300]), .Z(n39021) );
  XOR U56390 ( .A(x[1299]), .B(y[1299]), .Z(n38527) );
  IV U56391 ( .A(n38527), .Z(n39020) );
  IV U56392 ( .A(x[1298]), .Z(n38528) );
  XOR U56393 ( .A(n38528), .B(y[1298]), .Z(n39029) );
  XOR U56394 ( .A(x[1297]), .B(y[1297]), .Z(n39025) );
  XOR U56395 ( .A(x[1296]), .B(y[1296]), .Z(n39030) );
  XOR U56396 ( .A(x[1295]), .B(y[1295]), .Z(n39036) );
  XOR U56397 ( .A(x[1294]), .B(y[1294]), .Z(n39033) );
  XOR U56398 ( .A(x[1293]), .B(y[1293]), .Z(n39042) );
  XOR U56399 ( .A(x[1292]), .B(y[1292]), .Z(n39039) );
  XOR U56400 ( .A(x[1291]), .B(y[1291]), .Z(n39045) );
  XOR U56401 ( .A(x[1290]), .B(y[1290]), .Z(n43770) );
  XOR U56402 ( .A(x[1289]), .B(y[1289]), .Z(n43767) );
  XOR U56403 ( .A(x[1288]), .B(y[1288]), .Z(n39051) );
  XOR U56404 ( .A(x[1287]), .B(y[1287]), .Z(n39048) );
  XOR U56405 ( .A(x[1286]), .B(y[1286]), .Z(n39057) );
  XOR U56406 ( .A(x[1285]), .B(y[1285]), .Z(n39054) );
  XOR U56407 ( .A(x[1282]), .B(y[1282]), .Z(n39065) );
  XOR U56408 ( .A(x[1281]), .B(y[1281]), .Z(n43754) );
  XOR U56409 ( .A(x[1280]), .B(y[1280]), .Z(n43748) );
  XOR U56410 ( .A(x[1279]), .B(y[1279]), .Z(n43745) );
  XOR U56411 ( .A(x[1278]), .B(y[1278]), .Z(n43741) );
  XOR U56412 ( .A(x[1277]), .B(y[1277]), .Z(n43738) );
  XOR U56413 ( .A(x[1276]), .B(y[1276]), .Z(n43734) );
  XOR U56414 ( .A(x[1275]), .B(y[1275]), .Z(n43731) );
  XOR U56415 ( .A(x[1274]), .B(y[1274]), .Z(n39071) );
  XOR U56416 ( .A(x[1273]), .B(y[1273]), .Z(n39068) );
  XOR U56417 ( .A(x[1272]), .B(y[1272]), .Z(n39077) );
  XOR U56418 ( .A(x[1271]), .B(y[1271]), .Z(n39074) );
  XOR U56419 ( .A(x[1270]), .B(y[1270]), .Z(n39083) );
  XOR U56420 ( .A(x[1269]), .B(y[1269]), .Z(n39080) );
  XOR U56421 ( .A(x[1268]), .B(y[1268]), .Z(n39086) );
  XOR U56422 ( .A(x[1267]), .B(y[1267]), .Z(n39092) );
  XOR U56423 ( .A(x[1266]), .B(y[1266]), .Z(n39089) );
  XOR U56424 ( .A(x[1265]), .B(y[1265]), .Z(n39098) );
  XOR U56425 ( .A(x[1264]), .B(y[1264]), .Z(n39095) );
  XOR U56426 ( .A(x[1263]), .B(y[1263]), .Z(n43725) );
  XOR U56427 ( .A(x[1262]), .B(y[1262]), .Z(n43722) );
  XOR U56428 ( .A(x[1261]), .B(y[1261]), .Z(n39104) );
  XOR U56429 ( .A(x[1260]), .B(y[1260]), .Z(n39101) );
  XOR U56430 ( .A(x[1259]), .B(y[1259]), .Z(n39110) );
  XOR U56431 ( .A(x[1258]), .B(y[1258]), .Z(n39107) );
  XOR U56432 ( .A(x[1257]), .B(y[1257]), .Z(n43717) );
  XOR U56433 ( .A(x[1256]), .B(y[1256]), .Z(n43714) );
  XOR U56434 ( .A(x[1255]), .B(y[1255]), .Z(n39113) );
  XOR U56435 ( .A(x[1254]), .B(y[1254]), .Z(n43709) );
  XOR U56436 ( .A(x[1253]), .B(y[1253]), .Z(n43706) );
  XOR U56437 ( .A(x[1252]), .B(y[1252]), .Z(n39120) );
  XOR U56438 ( .A(x[1251]), .B(y[1251]), .Z(n39119) );
  IV U56439 ( .A(n39119), .Z(n39117) );
  XOR U56440 ( .A(x[1250]), .B(y[1250]), .Z(n39123) );
  XOR U56441 ( .A(x[1249]), .B(y[1249]), .Z(n43702) );
  XOR U56442 ( .A(x[1248]), .B(y[1248]), .Z(n43699) );
  XOR U56443 ( .A(x[1247]), .B(y[1247]), .Z(n39126) );
  XOR U56444 ( .A(x[1246]), .B(y[1246]), .Z(n39132) );
  XOR U56445 ( .A(x[1245]), .B(y[1245]), .Z(n39129) );
  XOR U56446 ( .A(x[1244]), .B(y[1244]), .Z(n43696) );
  XOR U56447 ( .A(x[1243]), .B(y[1243]), .Z(n43693) );
  XOR U56448 ( .A(x[1242]), .B(y[1242]), .Z(n38529) );
  IV U56449 ( .A(n38529), .Z(n43691) );
  IV U56450 ( .A(x[1241]), .Z(n38530) );
  XOR U56451 ( .A(n38530), .B(y[1241]), .Z(n43688) );
  XOR U56452 ( .A(x[1240]), .B(y[1240]), .Z(n43684) );
  XOR U56453 ( .A(x[1239]), .B(y[1239]), .Z(n43681) );
  XOR U56454 ( .A(x[1238]), .B(y[1238]), .Z(n39138) );
  XOR U56455 ( .A(x[1237]), .B(y[1237]), .Z(n39135) );
  XOR U56456 ( .A(x[1236]), .B(y[1236]), .Z(n43677) );
  XOR U56457 ( .A(x[1235]), .B(y[1235]), .Z(n43674) );
  XOR U56458 ( .A(x[1234]), .B(y[1234]), .Z(n39145) );
  XOR U56459 ( .A(x[1233]), .B(y[1233]), .Z(n39142) );
  XOR U56460 ( .A(x[1232]), .B(y[1232]), .Z(n43670) );
  XOR U56461 ( .A(x[1231]), .B(y[1231]), .Z(n43667) );
  XOR U56462 ( .A(x[1230]), .B(y[1230]), .Z(n38531) );
  IV U56463 ( .A(n38531), .Z(n43665) );
  IV U56464 ( .A(x[1229]), .Z(n38532) );
  XOR U56465 ( .A(n38532), .B(y[1229]), .Z(n43662) );
  XOR U56466 ( .A(x[1228]), .B(y[1228]), .Z(n43658) );
  XOR U56467 ( .A(x[1227]), .B(y[1227]), .Z(n43655) );
  XOR U56468 ( .A(x[1226]), .B(y[1226]), .Z(n39148) );
  XOR U56469 ( .A(x[1225]), .B(y[1225]), .Z(n43645) );
  XOR U56470 ( .A(x[1224]), .B(y[1224]), .Z(n39154) );
  XOR U56471 ( .A(x[1223]), .B(y[1223]), .Z(n39151) );
  XOR U56472 ( .A(x[1222]), .B(y[1222]), .Z(n43638) );
  XOR U56473 ( .A(x[1221]), .B(y[1221]), .Z(n43635) );
  XOR U56474 ( .A(x[1220]), .B(y[1220]), .Z(n39157) );
  XOR U56475 ( .A(x[1219]), .B(y[1219]), .Z(n43627) );
  XOR U56476 ( .A(x[1218]), .B(y[1218]), .Z(n38533) );
  IV U56477 ( .A(n38533), .Z(n39162) );
  IV U56478 ( .A(x[1217]), .Z(n38534) );
  XOR U56479 ( .A(n38534), .B(y[1217]), .Z(n43622) );
  XOR U56480 ( .A(x[1216]), .B(y[1216]), .Z(n43619) );
  XOR U56481 ( .A(x[1215]), .B(y[1215]), .Z(n39163) );
  XOR U56482 ( .A(x[1214]), .B(y[1214]), .Z(n43614) );
  XOR U56483 ( .A(x[1213]), .B(y[1213]), .Z(n43611) );
  XOR U56484 ( .A(x[1212]), .B(y[1212]), .Z(n43607) );
  XOR U56485 ( .A(x[1211]), .B(y[1211]), .Z(n43604) );
  XOR U56486 ( .A(x[1210]), .B(y[1210]), .Z(n39166) );
  XOR U56487 ( .A(x[1209]), .B(y[1209]), .Z(n43593) );
  XOR U56488 ( .A(x[1208]), .B(y[1208]), .Z(n39169) );
  XOR U56489 ( .A(x[1207]), .B(y[1207]), .Z(n43585) );
  XOR U56490 ( .A(x[1206]), .B(y[1206]), .Z(n38535) );
  IV U56491 ( .A(n38535), .Z(n39174) );
  IV U56492 ( .A(x[1205]), .Z(n38536) );
  XOR U56493 ( .A(n38536), .B(y[1205]), .Z(n43580) );
  XOR U56494 ( .A(x[1204]), .B(y[1204]), .Z(n43577) );
  XOR U56495 ( .A(x[1203]), .B(y[1203]), .Z(n43573) );
  XOR U56496 ( .A(x[1202]), .B(y[1202]), .Z(n43570) );
  XOR U56497 ( .A(x[1201]), .B(y[1201]), .Z(n43566) );
  XOR U56498 ( .A(x[1200]), .B(y[1200]), .Z(n43563) );
  XOR U56499 ( .A(x[1199]), .B(y[1199]), .Z(n39175) );
  XOR U56500 ( .A(x[1198]), .B(y[1198]), .Z(n43558) );
  XOR U56501 ( .A(x[1197]), .B(y[1197]), .Z(n43555) );
  XOR U56502 ( .A(x[1196]), .B(y[1196]), .Z(n43551) );
  XOR U56503 ( .A(x[1195]), .B(y[1195]), .Z(n43548) );
  XOR U56504 ( .A(x[1194]), .B(y[1194]), .Z(n43544) );
  XOR U56505 ( .A(x[1193]), .B(y[1193]), .Z(n43541) );
  XOR U56506 ( .A(x[1192]), .B(y[1192]), .Z(n43537) );
  XOR U56507 ( .A(x[1191]), .B(y[1191]), .Z(n43534) );
  XOR U56508 ( .A(x[1190]), .B(y[1190]), .Z(n39181) );
  XOR U56509 ( .A(x[1189]), .B(y[1189]), .Z(n39178) );
  XOR U56510 ( .A(x[1184]), .B(y[1184]), .Z(n39192) );
  XOR U56511 ( .A(x[1183]), .B(y[1183]), .Z(n39189) );
  XOR U56512 ( .A(x[1182]), .B(y[1182]), .Z(n39198) );
  XOR U56513 ( .A(x[1181]), .B(y[1181]), .Z(n39195) );
  XOR U56514 ( .A(x[1180]), .B(y[1180]), .Z(n39201) );
  XOR U56515 ( .A(x[1179]), .B(y[1179]), .Z(n39207) );
  XOR U56516 ( .A(x[1178]), .B(y[1178]), .Z(n39204) );
  XOR U56517 ( .A(x[1177]), .B(y[1177]), .Z(n39213) );
  XOR U56518 ( .A(x[1176]), .B(y[1176]), .Z(n38537) );
  IV U56519 ( .A(n38537), .Z(n39211) );
  IV U56520 ( .A(x[1175]), .Z(n38538) );
  XOR U56521 ( .A(n38538), .B(y[1175]), .Z(n39217) );
  XOR U56522 ( .A(x[1174]), .B(y[1174]), .Z(n43523) );
  XOR U56523 ( .A(x[1173]), .B(y[1173]), .Z(n43520) );
  XOR U56524 ( .A(x[1172]), .B(y[1172]), .Z(n39221) );
  XOR U56525 ( .A(x[1171]), .B(y[1171]), .Z(n39218) );
  XOR U56526 ( .A(x[1170]), .B(y[1170]), .Z(n43517) );
  XOR U56527 ( .A(x[1169]), .B(y[1169]), .Z(n43514) );
  XOR U56528 ( .A(x[1168]), .B(y[1168]), .Z(n43510) );
  XOR U56529 ( .A(x[1167]), .B(y[1167]), .Z(n43507) );
  XOR U56530 ( .A(x[1166]), .B(y[1166]), .Z(n43492) );
  XOR U56531 ( .A(x[1165]), .B(y[1165]), .Z(n43498) );
  XOR U56532 ( .A(x[1164]), .B(y[1164]), .Z(n38539) );
  IV U56533 ( .A(n38539), .Z(n43497) );
  IV U56534 ( .A(x[1163]), .Z(n38540) );
  XOR U56535 ( .A(n38540), .B(y[1163]), .Z(n43489) );
  XOR U56536 ( .A(x[1162]), .B(y[1162]), .Z(n43486) );
  XOR U56537 ( .A(x[1161]), .B(y[1161]), .Z(n39224) );
  XOR U56538 ( .A(x[1160]), .B(y[1160]), .Z(n43480) );
  XOR U56539 ( .A(x[1159]), .B(y[1159]), .Z(n39227) );
  XOR U56540 ( .A(x[1158]), .B(y[1158]), .Z(n43475) );
  XOR U56541 ( .A(x[1157]), .B(y[1157]), .Z(n43472) );
  XOR U56542 ( .A(x[1156]), .B(y[1156]), .Z(n39233) );
  XOR U56543 ( .A(x[1155]), .B(y[1155]), .Z(n39230) );
  XOR U56544 ( .A(x[1154]), .B(y[1154]), .Z(n43469) );
  XOR U56545 ( .A(x[1153]), .B(y[1153]), .Z(n43466) );
  XOR U56546 ( .A(x[1152]), .B(y[1152]), .Z(n38541) );
  IV U56547 ( .A(n38541), .Z(n39238) );
  IV U56548 ( .A(x[1151]), .Z(n38542) );
  XOR U56549 ( .A(n38542), .B(y[1151]), .Z(n43460) );
  XOR U56550 ( .A(x[1150]), .B(y[1150]), .Z(n39239) );
  XOR U56551 ( .A(x[1149]), .B(y[1149]), .Z(n43454) );
  XOR U56552 ( .A(x[1148]), .B(y[1148]), .Z(n43451) );
  XOR U56553 ( .A(x[1147]), .B(y[1147]), .Z(n39245) );
  XOR U56554 ( .A(x[1146]), .B(y[1146]), .Z(n39242) );
  XOR U56555 ( .A(x[1145]), .B(y[1145]), .Z(n39248) );
  XOR U56556 ( .A(x[1144]), .B(y[1144]), .Z(n43441) );
  XOR U56557 ( .A(x[1143]), .B(y[1143]), .Z(n43438) );
  XOR U56558 ( .A(x[1142]), .B(y[1142]), .Z(n39254) );
  XOR U56559 ( .A(x[1141]), .B(y[1141]), .Z(n39251) );
  XOR U56560 ( .A(x[1140]), .B(y[1140]), .Z(n38543) );
  IV U56561 ( .A(n38543), .Z(n39260) );
  IV U56562 ( .A(x[1139]), .Z(n38544) );
  XOR U56563 ( .A(n38544), .B(y[1139]), .Z(n39258) );
  XOR U56564 ( .A(x[1138]), .B(y[1138]), .Z(n39262) );
  XOR U56565 ( .A(x[1137]), .B(y[1137]), .Z(n43432) );
  XOR U56566 ( .A(x[1136]), .B(y[1136]), .Z(n43429) );
  XOR U56567 ( .A(x[1135]), .B(y[1135]), .Z(n43425) );
  XOR U56568 ( .A(x[1134]), .B(y[1134]), .Z(n43422) );
  XOR U56569 ( .A(x[1133]), .B(y[1133]), .Z(n39268) );
  XOR U56570 ( .A(x[1132]), .B(y[1132]), .Z(n39265) );
  XOR U56571 ( .A(x[1131]), .B(y[1131]), .Z(n39275) );
  XOR U56572 ( .A(x[1130]), .B(y[1130]), .Z(n39272) );
  XOR U56573 ( .A(x[1129]), .B(y[1129]), .Z(n43418) );
  XOR U56574 ( .A(x[1128]), .B(y[1128]), .Z(n43415) );
  XOR U56575 ( .A(x[1127]), .B(y[1127]), .Z(n38545) );
  IV U56576 ( .A(n38545), .Z(n39280) );
  IV U56577 ( .A(x[1126]), .Z(n38546) );
  XOR U56578 ( .A(n38546), .B(y[1126]), .Z(n43412) );
  XOR U56579 ( .A(x[1125]), .B(y[1125]), .Z(n43409) );
  XOR U56580 ( .A(x[1124]), .B(y[1124]), .Z(n39281) );
  XOR U56581 ( .A(x[1123]), .B(y[1123]), .Z(n43401) );
  XOR U56582 ( .A(x[1122]), .B(y[1122]), .Z(n39284) );
  XOR U56583 ( .A(x[1121]), .B(y[1121]), .Z(n43395) );
  XOR U56584 ( .A(x[1120]), .B(y[1120]), .Z(n43392) );
  XOR U56585 ( .A(x[1119]), .B(y[1119]), .Z(n39287) );
  XOR U56586 ( .A(x[1118]), .B(y[1118]), .Z(n39294) );
  XOR U56587 ( .A(x[1117]), .B(y[1117]), .Z(n39291) );
  XOR U56588 ( .A(x[1116]), .B(y[1116]), .Z(n39300) );
  XOR U56589 ( .A(x[1115]), .B(y[1115]), .Z(n39297) );
  XOR U56590 ( .A(x[1114]), .B(y[1114]), .Z(n39303) );
  XOR U56591 ( .A(x[1113]), .B(y[1113]), .Z(n43381) );
  XOR U56592 ( .A(x[1112]), .B(y[1112]), .Z(n39306) );
  XOR U56593 ( .A(x[1111]), .B(y[1111]), .Z(n43360) );
  XOR U56594 ( .A(x[1110]), .B(y[1110]), .Z(n43357) );
  XOR U56595 ( .A(x[1109]), .B(y[1109]), .Z(n43353) );
  XOR U56596 ( .A(x[1108]), .B(y[1108]), .Z(n43350) );
  XOR U56597 ( .A(x[1107]), .B(y[1107]), .Z(n43346) );
  XOR U56598 ( .A(x[1106]), .B(y[1106]), .Z(n43343) );
  XOR U56599 ( .A(x[1105]), .B(y[1105]), .Z(n43339) );
  XOR U56600 ( .A(x[1104]), .B(y[1104]), .Z(n43336) );
  XOR U56601 ( .A(x[1103]), .B(y[1103]), .Z(n43332) );
  XOR U56602 ( .A(x[1102]), .B(y[1102]), .Z(n43329) );
  XOR U56603 ( .A(x[1101]), .B(y[1101]), .Z(n39309) );
  XOR U56604 ( .A(x[1100]), .B(y[1100]), .Z(n43323) );
  XOR U56605 ( .A(x[1099]), .B(y[1099]), .Z(n39312) );
  XOR U56606 ( .A(x[1096]), .B(y[1096]), .Z(n43313) );
  XOR U56607 ( .A(x[1095]), .B(y[1095]), .Z(n43310) );
  XOR U56608 ( .A(x[1094]), .B(y[1094]), .Z(n43306) );
  XOR U56609 ( .A(x[1093]), .B(y[1093]), .Z(n43303) );
  XOR U56610 ( .A(x[1092]), .B(y[1092]), .Z(n43299) );
  XOR U56611 ( .A(x[1091]), .B(y[1091]), .Z(n43296) );
  XOR U56612 ( .A(x[1090]), .B(y[1090]), .Z(n43292) );
  XOR U56613 ( .A(x[1089]), .B(y[1089]), .Z(n43289) );
  XOR U56614 ( .A(x[1088]), .B(y[1088]), .Z(n38547) );
  IV U56615 ( .A(n38547), .Z(n43287) );
  IV U56616 ( .A(x[1087]), .Z(n38548) );
  XOR U56617 ( .A(n38548), .B(y[1087]), .Z(n43285) );
  XOR U56618 ( .A(x[1086]), .B(y[1086]), .Z(n43280) );
  XOR U56619 ( .A(x[1085]), .B(y[1085]), .Z(n43277) );
  XOR U56620 ( .A(x[1084]), .B(y[1084]), .Z(n39315) );
  XOR U56621 ( .A(x[1083]), .B(y[1083]), .Z(n39322) );
  XOR U56622 ( .A(x[1082]), .B(y[1082]), .Z(n39319) );
  XOR U56623 ( .A(x[1081]), .B(y[1081]), .Z(n43272) );
  XOR U56624 ( .A(x[1080]), .B(y[1080]), .Z(n43269) );
  XOR U56625 ( .A(x[1079]), .B(y[1079]), .Z(n39328) );
  XOR U56626 ( .A(x[1078]), .B(y[1078]), .Z(n39325) );
  XOR U56627 ( .A(x[1077]), .B(y[1077]), .Z(n39331) );
  XOR U56628 ( .A(x[1076]), .B(y[1076]), .Z(n38549) );
  IV U56629 ( .A(n38549), .Z(n43265) );
  IV U56630 ( .A(x[1075]), .Z(n38550) );
  XOR U56631 ( .A(n38550), .B(y[1075]), .Z(n43263) );
  XOR U56632 ( .A(x[1074]), .B(y[1074]), .Z(n39337) );
  XOR U56633 ( .A(x[1073]), .B(y[1073]), .Z(n39334) );
  XOR U56634 ( .A(x[1072]), .B(y[1072]), .Z(n43250) );
  XOR U56635 ( .A(x[1071]), .B(y[1071]), .Z(n39340) );
  XOR U56636 ( .A(x[1070]), .B(y[1070]), .Z(n43253) );
  XOR U56637 ( .A(x[1069]), .B(y[1069]), .Z(n43246) );
  XOR U56638 ( .A(x[1068]), .B(y[1068]), .Z(n43243) );
  XOR U56639 ( .A(x[1067]), .B(y[1067]), .Z(n39347) );
  XOR U56640 ( .A(x[1066]), .B(y[1066]), .Z(n39344) );
  XOR U56641 ( .A(x[1065]), .B(y[1065]), .Z(n39353) );
  XOR U56642 ( .A(x[1064]), .B(y[1064]), .Z(n39350) );
  XOR U56643 ( .A(x[1063]), .B(y[1063]), .Z(n43238) );
  XOR U56644 ( .A(x[1062]), .B(y[1062]), .Z(n43235) );
  XOR U56645 ( .A(x[1061]), .B(y[1061]), .Z(n39356) );
  XOR U56646 ( .A(x[1058]), .B(y[1058]), .Z(n39362) );
  XOR U56647 ( .A(x[1057]), .B(y[1057]), .Z(n39359) );
  XOR U56648 ( .A(x[1056]), .B(y[1056]), .Z(n43225) );
  XOR U56649 ( .A(x[1055]), .B(y[1055]), .Z(n43222) );
  XOR U56650 ( .A(x[1054]), .B(y[1054]), .Z(n39369) );
  XOR U56651 ( .A(x[1053]), .B(y[1053]), .Z(n39366) );
  XOR U56652 ( .A(x[1052]), .B(y[1052]), .Z(n43219) );
  XOR U56653 ( .A(x[1051]), .B(y[1051]), .Z(n43216) );
  XOR U56654 ( .A(x[1050]), .B(y[1050]), .Z(n39375) );
  XOR U56655 ( .A(x[1049]), .B(y[1049]), .Z(n39372) );
  XOR U56656 ( .A(x[1048]), .B(y[1048]), .Z(n43212) );
  XOR U56657 ( .A(x[1047]), .B(y[1047]), .Z(n43209) );
  XOR U56658 ( .A(x[1046]), .B(y[1046]), .Z(n39381) );
  XOR U56659 ( .A(x[1045]), .B(y[1045]), .Z(n39378) );
  XOR U56660 ( .A(x[1044]), .B(y[1044]), .Z(n39387) );
  XOR U56661 ( .A(x[1043]), .B(y[1043]), .Z(n39384) );
  XOR U56662 ( .A(x[1042]), .B(y[1042]), .Z(n39393) );
  XOR U56663 ( .A(x[1041]), .B(y[1041]), .Z(n39390) );
  XOR U56664 ( .A(x[1040]), .B(y[1040]), .Z(n39399) );
  XOR U56665 ( .A(x[1039]), .B(y[1039]), .Z(n39396) );
  XOR U56666 ( .A(x[1038]), .B(y[1038]), .Z(n43204) );
  XOR U56667 ( .A(x[1037]), .B(y[1037]), .Z(n43201) );
  XOR U56668 ( .A(x[1036]), .B(y[1036]), .Z(n39405) );
  XOR U56669 ( .A(x[1035]), .B(y[1035]), .Z(n39402) );
  XOR U56670 ( .A(x[1034]), .B(y[1034]), .Z(n39411) );
  XOR U56671 ( .A(x[1033]), .B(y[1033]), .Z(n39408) );
  XOR U56672 ( .A(x[1032]), .B(y[1032]), .Z(n43197) );
  XOR U56673 ( .A(x[1031]), .B(y[1031]), .Z(n43194) );
  XOR U56674 ( .A(x[1030]), .B(y[1030]), .Z(n39417) );
  XOR U56675 ( .A(x[1029]), .B(y[1029]), .Z(n39414) );
  XOR U56676 ( .A(x[1028]), .B(y[1028]), .Z(n43182) );
  XOR U56677 ( .A(x[1027]), .B(y[1027]), .Z(n39420) );
  XOR U56678 ( .A(x[1026]), .B(y[1026]), .Z(n43185) );
  XOR U56679 ( .A(x[1025]), .B(y[1025]), .Z(n39424) );
  XOR U56680 ( .A(x[1024]), .B(y[1024]), .Z(n43178) );
  XOR U56681 ( .A(x[1023]), .B(y[1023]), .Z(n43175) );
  XOR U56682 ( .A(x[1022]), .B(y[1022]), .Z(n39430) );
  XOR U56683 ( .A(x[1021]), .B(y[1021]), .Z(n39427) );
  XOR U56684 ( .A(x[1020]), .B(y[1020]), .Z(n39436) );
  XOR U56685 ( .A(x[1019]), .B(y[1019]), .Z(n39433) );
  XOR U56686 ( .A(x[1018]), .B(y[1018]), .Z(n39442) );
  XOR U56687 ( .A(x[1017]), .B(y[1017]), .Z(n39439) );
  XOR U56688 ( .A(x[1016]), .B(y[1016]), .Z(n39445) );
  XOR U56689 ( .A(x[1015]), .B(y[1015]), .Z(n39451) );
  XOR U56690 ( .A(x[1014]), .B(y[1014]), .Z(n39448) );
  XOR U56691 ( .A(x[1013]), .B(y[1013]), .Z(n39457) );
  XOR U56692 ( .A(x[1012]), .B(y[1012]), .Z(n39454) );
  XOR U56693 ( .A(x[1011]), .B(y[1011]), .Z(n39460) );
  XOR U56694 ( .A(x[1010]), .B(y[1010]), .Z(n39466) );
  XOR U56695 ( .A(x[1009]), .B(y[1009]), .Z(n39463) );
  XOR U56696 ( .A(x[1008]), .B(y[1008]), .Z(n39472) );
  XOR U56697 ( .A(x[1007]), .B(y[1007]), .Z(n39469) );
  XOR U56698 ( .A(x[1006]), .B(y[1006]), .Z(n39476) );
  XOR U56699 ( .A(x[1005]), .B(y[1005]), .Z(n43168) );
  XOR U56700 ( .A(x[1004]), .B(y[1004]), .Z(n43165) );
  XOR U56701 ( .A(x[1003]), .B(y[1003]), .Z(n39482) );
  XOR U56702 ( .A(x[1002]), .B(y[1002]), .Z(n39479) );
  XOR U56703 ( .A(x[1001]), .B(y[1001]), .Z(n39485) );
  XOR U56704 ( .A(x[1000]), .B(y[1000]), .Z(n43159) );
  XOR U56705 ( .A(x[999]), .B(y[999]), .Z(n43156) );
  XOR U56706 ( .A(x[998]), .B(y[998]), .Z(n39491) );
  XOR U56707 ( .A(x[997]), .B(y[997]), .Z(n39488) );
  XOR U56708 ( .A(x[996]), .B(y[996]), .Z(n39500) );
  XOR U56709 ( .A(x[995]), .B(y[995]), .Z(n39497) );
  XOR U56710 ( .A(x[994]), .B(y[994]), .Z(n39494) );
  XOR U56711 ( .A(x[993]), .B(y[993]), .Z(n39506) );
  XOR U56712 ( .A(x[992]), .B(y[992]), .Z(n39503) );
  XOR U56713 ( .A(x[991]), .B(y[991]), .Z(n39512) );
  XOR U56714 ( .A(x[990]), .B(y[990]), .Z(n39509) );
  XOR U56715 ( .A(x[989]), .B(y[989]), .Z(n39515) );
  XOR U56716 ( .A(x[988]), .B(y[988]), .Z(n43145) );
  XOR U56717 ( .A(x[987]), .B(y[987]), .Z(n43142) );
  XOR U56718 ( .A(x[986]), .B(y[986]), .Z(n43138) );
  XOR U56719 ( .A(x[985]), .B(y[985]), .Z(n43135) );
  XOR U56720 ( .A(x[984]), .B(y[984]), .Z(n43131) );
  XOR U56721 ( .A(x[983]), .B(y[983]), .Z(n43128) );
  XOR U56722 ( .A(x[982]), .B(y[982]), .Z(n43124) );
  XOR U56723 ( .A(x[981]), .B(y[981]), .Z(n43121) );
  XOR U56724 ( .A(x[980]), .B(y[980]), .Z(n43117) );
  XOR U56725 ( .A(x[979]), .B(y[979]), .Z(n43114) );
  XOR U56726 ( .A(x[978]), .B(y[978]), .Z(n39521) );
  XOR U56727 ( .A(x[977]), .B(y[977]), .Z(n39518) );
  XOR U56728 ( .A(x[976]), .B(y[976]), .Z(n43108) );
  XOR U56729 ( .A(x[975]), .B(y[975]), .Z(n43105) );
  XOR U56730 ( .A(x[974]), .B(y[974]), .Z(n39527) );
  XOR U56731 ( .A(x[973]), .B(y[973]), .Z(n39524) );
  XOR U56732 ( .A(x[972]), .B(y[972]), .Z(n39530) );
  XOR U56733 ( .A(x[971]), .B(y[971]), .Z(n39533) );
  XOR U56734 ( .A(x[970]), .B(y[970]), .Z(n43093) );
  XOR U56735 ( .A(x[969]), .B(y[969]), .Z(n39536) );
  XOR U56736 ( .A(x[968]), .B(y[968]), .Z(n39542) );
  XOR U56737 ( .A(x[967]), .B(y[967]), .Z(n39539) );
  XOR U56738 ( .A(x[966]), .B(y[966]), .Z(n39549) );
  XOR U56739 ( .A(x[965]), .B(y[965]), .Z(n39546) );
  XOR U56740 ( .A(x[964]), .B(y[964]), .Z(n43086) );
  XOR U56741 ( .A(x[963]), .B(y[963]), .Z(n43083) );
  XOR U56742 ( .A(x[962]), .B(y[962]), .Z(n43079) );
  XOR U56743 ( .A(x[961]), .B(y[961]), .Z(n43078) );
  XOR U56744 ( .A(x[960]), .B(y[960]), .Z(n43071) );
  XOR U56745 ( .A(x[959]), .B(y[959]), .Z(n43068) );
  XOR U56746 ( .A(x[958]), .B(y[958]), .Z(n39552) );
  XOR U56747 ( .A(x[957]), .B(y[957]), .Z(n39558) );
  XOR U56748 ( .A(x[956]), .B(y[956]), .Z(n39555) );
  XOR U56749 ( .A(x[955]), .B(y[955]), .Z(n39564) );
  XOR U56750 ( .A(x[954]), .B(y[954]), .Z(n39561) );
  XOR U56751 ( .A(x[953]), .B(y[953]), .Z(n39571) );
  XOR U56752 ( .A(x[952]), .B(y[952]), .Z(n39568) );
  XOR U56753 ( .A(x[951]), .B(y[951]), .Z(n39574) );
  XOR U56754 ( .A(x[950]), .B(y[950]), .Z(n39580) );
  XOR U56755 ( .A(x[949]), .B(y[949]), .Z(n39577) );
  XOR U56756 ( .A(x[948]), .B(y[948]), .Z(n39586) );
  XOR U56757 ( .A(x[947]), .B(y[947]), .Z(n39583) );
  XOR U56758 ( .A(x[946]), .B(y[946]), .Z(n39589) );
  XOR U56759 ( .A(x[945]), .B(y[945]), .Z(n43057) );
  XOR U56760 ( .A(x[944]), .B(y[944]), .Z(n43054) );
  XOR U56761 ( .A(x[943]), .B(y[943]), .Z(n39595) );
  XOR U56762 ( .A(x[942]), .B(y[942]), .Z(n39592) );
  XOR U56763 ( .A(x[941]), .B(y[941]), .Z(n39598) );
  XOR U56764 ( .A(x[940]), .B(y[940]), .Z(n43048) );
  XOR U56765 ( .A(x[939]), .B(y[939]), .Z(n43045) );
  XOR U56766 ( .A(x[938]), .B(y[938]), .Z(n39601) );
  XOR U56767 ( .A(x[937]), .B(y[937]), .Z(n39604) );
  XOR U56768 ( .A(x[936]), .B(y[936]), .Z(n43033) );
  XOR U56769 ( .A(x[935]), .B(y[935]), .Z(n39607) );
  XOR U56770 ( .A(x[934]), .B(y[934]), .Z(n39614) );
  XOR U56771 ( .A(x[933]), .B(y[933]), .Z(n39611) );
  XOR U56772 ( .A(x[932]), .B(y[932]), .Z(n39620) );
  XOR U56773 ( .A(x[931]), .B(y[931]), .Z(n39617) );
  XOR U56774 ( .A(x[930]), .B(y[930]), .Z(n39623) );
  XOR U56775 ( .A(x[929]), .B(y[929]), .Z(n43025) );
  XOR U56776 ( .A(x[928]), .B(y[928]), .Z(n43022) );
  XOR U56777 ( .A(x[927]), .B(y[927]), .Z(n39629) );
  XOR U56778 ( .A(x[926]), .B(y[926]), .Z(n39626) );
  XOR U56779 ( .A(x[925]), .B(y[925]), .Z(n39635) );
  XOR U56780 ( .A(x[924]), .B(y[924]), .Z(n39632) );
  XOR U56781 ( .A(x[923]), .B(y[923]), .Z(n43018) );
  XOR U56782 ( .A(x[922]), .B(y[922]), .Z(n43015) );
  XOR U56783 ( .A(x[921]), .B(y[921]), .Z(n39638) );
  XOR U56784 ( .A(x[920]), .B(y[920]), .Z(n43011) );
  XOR U56785 ( .A(x[919]), .B(y[919]), .Z(n43008) );
  XOR U56786 ( .A(x[918]), .B(y[918]), .Z(n39645) );
  XOR U56787 ( .A(x[917]), .B(y[917]), .Z(n39642) );
  XOR U56788 ( .A(x[916]), .B(y[916]), .Z(n43004) );
  XOR U56789 ( .A(x[915]), .B(y[915]), .Z(n43001) );
  XOR U56790 ( .A(x[914]), .B(y[914]), .Z(n42990) );
  XOR U56791 ( .A(x[913]), .B(y[913]), .Z(n39648) );
  XOR U56792 ( .A(x[912]), .B(y[912]), .Z(n42993) );
  XOR U56793 ( .A(x[911]), .B(y[911]), .Z(n42986) );
  XOR U56794 ( .A(x[910]), .B(y[910]), .Z(n42975) );
  XOR U56795 ( .A(x[909]), .B(y[909]), .Z(n39652) );
  XOR U56796 ( .A(x[908]), .B(y[908]), .Z(n42978) );
  XOR U56797 ( .A(x[907]), .B(y[907]), .Z(n39659) );
  XOR U56798 ( .A(x[906]), .B(y[906]), .Z(n39656) );
  XOR U56799 ( .A(x[905]), .B(y[905]), .Z(n42971) );
  XOR U56800 ( .A(x[904]), .B(y[904]), .Z(n42968) );
  XOR U56801 ( .A(x[903]), .B(y[903]), .Z(n39662) );
  XOR U56802 ( .A(x[902]), .B(y[902]), .Z(n39666) );
  XOR U56803 ( .A(x[901]), .B(y[901]), .Z(n42956) );
  XOR U56804 ( .A(x[900]), .B(y[900]), .Z(n39669) );
  XOR U56805 ( .A(x[899]), .B(y[899]), .Z(n42946) );
  XOR U56806 ( .A(x[898]), .B(y[898]), .Z(n39672) );
  XOR U56807 ( .A(x[897]), .B(y[897]), .Z(n42940) );
  XOR U56808 ( .A(x[896]), .B(y[896]), .Z(n42937) );
  XOR U56809 ( .A(x[895]), .B(y[895]), .Z(n42933) );
  XOR U56810 ( .A(x[894]), .B(y[894]), .Z(n42930) );
  XOR U56811 ( .A(x[893]), .B(y[893]), .Z(n42926) );
  XOR U56812 ( .A(x[892]), .B(y[892]), .Z(n42923) );
  XOR U56813 ( .A(x[891]), .B(y[891]), .Z(n42919) );
  XOR U56814 ( .A(x[890]), .B(y[890]), .Z(n42916) );
  XOR U56815 ( .A(x[889]), .B(y[889]), .Z(n42912) );
  XOR U56816 ( .A(x[888]), .B(y[888]), .Z(n42909) );
  XOR U56817 ( .A(x[887]), .B(y[887]), .Z(n42906) );
  XOR U56818 ( .A(x[886]), .B(y[886]), .Z(n42903) );
  XOR U56819 ( .A(x[885]), .B(y[885]), .Z(n42889) );
  XOR U56820 ( .A(x[884]), .B(y[884]), .Z(n42886) );
  XOR U56821 ( .A(x[883]), .B(y[883]), .Z(n39675) );
  XOR U56822 ( .A(x[882]), .B(y[882]), .Z(n39681) );
  XOR U56823 ( .A(x[881]), .B(y[881]), .Z(n39678) );
  XOR U56824 ( .A(x[880]), .B(y[880]), .Z(n42881) );
  XOR U56825 ( .A(x[879]), .B(y[879]), .Z(n42878) );
  XOR U56826 ( .A(x[878]), .B(y[878]), .Z(n39687) );
  XOR U56827 ( .A(x[877]), .B(y[877]), .Z(n39684) );
  XOR U56828 ( .A(x[876]), .B(y[876]), .Z(n42874) );
  XOR U56829 ( .A(x[875]), .B(y[875]), .Z(n42871) );
  XOR U56830 ( .A(x[874]), .B(y[874]), .Z(n42868) );
  XOR U56831 ( .A(x[873]), .B(y[873]), .Z(n42865) );
  XOR U56832 ( .A(x[872]), .B(y[872]), .Z(n42861) );
  XOR U56833 ( .A(x[871]), .B(y[871]), .Z(n42858) );
  XOR U56834 ( .A(x[870]), .B(y[870]), .Z(n39693) );
  XOR U56835 ( .A(x[869]), .B(y[869]), .Z(n39690) );
  XOR U56836 ( .A(x[868]), .B(y[868]), .Z(n42853) );
  XOR U56837 ( .A(x[867]), .B(y[867]), .Z(n42850) );
  XOR U56838 ( .A(x[866]), .B(y[866]), .Z(n55409) );
  XOR U56839 ( .A(x[865]), .B(y[865]), .Z(n42845) );
  XOR U56840 ( .A(x[864]), .B(y[864]), .Z(n39699) );
  XOR U56841 ( .A(x[863]), .B(y[863]), .Z(n39696) );
  XOR U56842 ( .A(x[862]), .B(y[862]), .Z(n42840) );
  XOR U56843 ( .A(x[861]), .B(y[861]), .Z(n42837) );
  XOR U56844 ( .A(x[860]), .B(y[860]), .Z(n42833) );
  XOR U56845 ( .A(x[859]), .B(y[859]), .Z(n42830) );
  XOR U56846 ( .A(x[858]), .B(y[858]), .Z(n42826) );
  XOR U56847 ( .A(x[857]), .B(y[857]), .Z(n42823) );
  XOR U56848 ( .A(x[856]), .B(y[856]), .Z(n42820) );
  XOR U56849 ( .A(x[855]), .B(y[855]), .Z(n42817) );
  XOR U56850 ( .A(x[854]), .B(y[854]), .Z(n42813) );
  XOR U56851 ( .A(x[853]), .B(y[853]), .Z(n42810) );
  XOR U56852 ( .A(x[852]), .B(y[852]), .Z(n39702) );
  XOR U56853 ( .A(x[851]), .B(y[851]), .Z(n39708) );
  XOR U56854 ( .A(x[850]), .B(y[850]), .Z(n39705) );
  XOR U56855 ( .A(x[849]), .B(y[849]), .Z(n42805) );
  XOR U56856 ( .A(x[848]), .B(y[848]), .Z(n42802) );
  XOR U56857 ( .A(x[847]), .B(y[847]), .Z(n39711) );
  XOR U56858 ( .A(x[846]), .B(y[846]), .Z(n42796) );
  XOR U56859 ( .A(x[845]), .B(y[845]), .Z(n39714) );
  XOR U56860 ( .A(x[844]), .B(y[844]), .Z(n42789) );
  XOR U56861 ( .A(x[843]), .B(y[843]), .Z(n42786) );
  XOR U56862 ( .A(x[842]), .B(y[842]), .Z(n39720) );
  XOR U56863 ( .A(x[841]), .B(y[841]), .Z(n39717) );
  XOR U56864 ( .A(x[840]), .B(y[840]), .Z(n42782) );
  XOR U56865 ( .A(x[839]), .B(y[839]), .Z(n42779) );
  XOR U56866 ( .A(x[838]), .B(y[838]), .Z(n42775) );
  XOR U56867 ( .A(x[837]), .B(y[837]), .Z(n42772) );
  XOR U56868 ( .A(x[836]), .B(y[836]), .Z(n42768) );
  XOR U56869 ( .A(x[835]), .B(y[835]), .Z(n42765) );
  XOR U56870 ( .A(x[834]), .B(y[834]), .Z(n47599) );
  XOR U56871 ( .A(x[833]), .B(y[833]), .Z(n47586) );
  XOR U56872 ( .A(x[832]), .B(y[832]), .Z(n39723) );
  XOR U56873 ( .A(x[831]), .B(y[831]), .Z(n39729) );
  XOR U56874 ( .A(x[830]), .B(y[830]), .Z(n39726) );
  XOR U56875 ( .A(x[829]), .B(y[829]), .Z(n42756) );
  XOR U56876 ( .A(x[828]), .B(y[828]), .Z(n42753) );
  XOR U56877 ( .A(x[827]), .B(y[827]), .Z(n39736) );
  XOR U56878 ( .A(x[826]), .B(y[826]), .Z(n39733) );
  XOR U56879 ( .A(x[825]), .B(y[825]), .Z(n39742) );
  XOR U56880 ( .A(x[824]), .B(y[824]), .Z(n39739) );
  XOR U56881 ( .A(x[823]), .B(y[823]), .Z(n39748) );
  XOR U56882 ( .A(x[822]), .B(y[822]), .Z(n39745) );
  XOR U56883 ( .A(x[821]), .B(y[821]), .Z(n39751) );
  XOR U56884 ( .A(x[820]), .B(y[820]), .Z(n38551) );
  IV U56885 ( .A(n38551), .Z(n39757) );
  IV U56886 ( .A(x[819]), .Z(n38552) );
  XOR U56887 ( .A(n38552), .B(y[819]), .Z(n39754) );
  XOR U56888 ( .A(x[818]), .B(y[818]), .Z(n39762) );
  XOR U56889 ( .A(x[817]), .B(y[817]), .Z(n39759) );
  XOR U56890 ( .A(x[816]), .B(y[816]), .Z(n38553) );
  IV U56891 ( .A(n38553), .Z(n39767) );
  IV U56892 ( .A(x[815]), .Z(n38554) );
  XOR U56893 ( .A(n38554), .B(y[815]), .Z(n39772) );
  XOR U56894 ( .A(x[814]), .B(y[814]), .Z(n39768) );
  XOR U56895 ( .A(x[813]), .B(y[813]), .Z(n42742) );
  XOR U56896 ( .A(x[812]), .B(y[812]), .Z(n38555) );
  IV U56897 ( .A(n38555), .Z(n42740) );
  IV U56898 ( .A(x[811]), .Z(n38556) );
  XOR U56899 ( .A(n38556), .B(y[811]), .Z(n42736) );
  XOR U56900 ( .A(x[810]), .B(y[810]), .Z(n42733) );
  XOR U56901 ( .A(x[809]), .B(y[809]), .Z(n42729) );
  XOR U56902 ( .A(x[808]), .B(y[808]), .Z(n38557) );
  IV U56903 ( .A(n38557), .Z(n42727) );
  IV U56904 ( .A(x[807]), .Z(n38558) );
  XOR U56905 ( .A(n38558), .B(y[807]), .Z(n42723) );
  XOR U56906 ( .A(x[806]), .B(y[806]), .Z(n42720) );
  XOR U56907 ( .A(x[805]), .B(y[805]), .Z(n42715) );
  XOR U56908 ( .A(x[804]), .B(y[804]), .Z(n38559) );
  IV U56909 ( .A(n38559), .Z(n42713) );
  IV U56910 ( .A(x[803]), .Z(n38560) );
  XOR U56911 ( .A(n38560), .B(y[803]), .Z(n39773) );
  XOR U56912 ( .A(x[802]), .B(y[802]), .Z(n39778) );
  XOR U56913 ( .A(x[801]), .B(y[801]), .Z(n39775) );
  XOR U56914 ( .A(x[800]), .B(y[800]), .Z(n38561) );
  IV U56915 ( .A(n38561), .Z(n39784) );
  IV U56916 ( .A(x[799]), .Z(n38562) );
  XOR U56917 ( .A(n38562), .B(y[799]), .Z(n42708) );
  XOR U56918 ( .A(x[798]), .B(y[798]), .Z(n42704) );
  XOR U56919 ( .A(x[797]), .B(y[797]), .Z(n39785) );
  XOR U56920 ( .A(x[796]), .B(y[796]), .Z(n38563) );
  IV U56921 ( .A(n38563), .Z(n42700) );
  IV U56922 ( .A(x[795]), .Z(n38564) );
  XOR U56923 ( .A(n38564), .B(y[795]), .Z(n42698) );
  XOR U56924 ( .A(x[794]), .B(y[794]), .Z(n42693) );
  XOR U56925 ( .A(x[793]), .B(y[793]), .Z(n42690) );
  XOR U56926 ( .A(x[792]), .B(y[792]), .Z(n38565) );
  IV U56927 ( .A(n38565), .Z(n39790) );
  IV U56928 ( .A(x[791]), .Z(n38566) );
  XOR U56929 ( .A(n38566), .B(y[791]), .Z(n42682) );
  XOR U56930 ( .A(x[790]), .B(y[790]), .Z(n42675) );
  XOR U56931 ( .A(x[789]), .B(y[789]), .Z(n42672) );
  XOR U56932 ( .A(x[788]), .B(y[788]), .Z(n38567) );
  IV U56933 ( .A(n38567), .Z(n39794) );
  IV U56934 ( .A(x[787]), .Z(n38568) );
  XOR U56935 ( .A(n38568), .B(y[787]), .Z(n39791) );
  XOR U56936 ( .A(x[786]), .B(y[786]), .Z(n38569) );
  IV U56937 ( .A(n38569), .Z(n42669) );
  IV U56938 ( .A(x[785]), .Z(n38570) );
  XOR U56939 ( .A(n38570), .B(y[785]), .Z(n42666) );
  XOR U56940 ( .A(x[784]), .B(y[784]), .Z(n38571) );
  IV U56941 ( .A(n38571), .Z(n39800) );
  IV U56942 ( .A(x[783]), .Z(n38572) );
  XOR U56943 ( .A(n38572), .B(y[783]), .Z(n39797) );
  XOR U56944 ( .A(x[782]), .B(y[782]), .Z(n38573) );
  IV U56945 ( .A(n38573), .Z(n42664) );
  IV U56946 ( .A(x[781]), .Z(n38574) );
  XOR U56947 ( .A(n38574), .B(y[781]), .Z(n42661) );
  XOR U56948 ( .A(x[780]), .B(y[780]), .Z(n38575) );
  IV U56949 ( .A(n38575), .Z(n39805) );
  IV U56950 ( .A(x[779]), .Z(n38576) );
  XOR U56951 ( .A(n38576), .B(y[779]), .Z(n39803) );
  XOR U56952 ( .A(x[778]), .B(y[778]), .Z(n39810) );
  XOR U56953 ( .A(x[777]), .B(y[777]), .Z(n39807) );
  XOR U56954 ( .A(x[776]), .B(y[776]), .Z(n42657) );
  XOR U56955 ( .A(x[775]), .B(y[775]), .Z(n42654) );
  XOR U56956 ( .A(x[774]), .B(y[774]), .Z(n42650) );
  XOR U56957 ( .A(x[773]), .B(y[773]), .Z(n42647) );
  XOR U56958 ( .A(x[772]), .B(y[772]), .Z(n39816) );
  XOR U56959 ( .A(x[771]), .B(y[771]), .Z(n39813) );
  XOR U56960 ( .A(x[770]), .B(y[770]), .Z(n42643) );
  XOR U56961 ( .A(x[769]), .B(y[769]), .Z(n47479) );
  XOR U56962 ( .A(x[768]), .B(y[768]), .Z(n42636) );
  XOR U56963 ( .A(x[767]), .B(y[767]), .Z(n42633) );
  XOR U56964 ( .A(x[766]), .B(y[766]), .Z(n39822) );
  XOR U56965 ( .A(x[765]), .B(y[765]), .Z(n39819) );
  XOR U56966 ( .A(x[764]), .B(y[764]), .Z(n39828) );
  XOR U56967 ( .A(x[763]), .B(y[763]), .Z(n39825) );
  XOR U56968 ( .A(x[762]), .B(y[762]), .Z(n39834) );
  XOR U56969 ( .A(x[761]), .B(y[761]), .Z(n39831) );
  XOR U56970 ( .A(x[760]), .B(y[760]), .Z(n39837) );
  XOR U56971 ( .A(x[759]), .B(y[759]), .Z(n39844) );
  XOR U56972 ( .A(x[758]), .B(y[758]), .Z(n39841) );
  XOR U56973 ( .A(x[757]), .B(y[757]), .Z(n39850) );
  XOR U56974 ( .A(x[756]), .B(y[756]), .Z(n38577) );
  IV U56975 ( .A(n38577), .Z(n39849) );
  IV U56976 ( .A(x[755]), .Z(n38578) );
  XOR U56977 ( .A(n38578), .B(y[755]), .Z(n42627) );
  XOR U56978 ( .A(x[754]), .B(y[754]), .Z(n42624) );
  XOR U56979 ( .A(x[753]), .B(y[753]), .Z(n42621) );
  XOR U56980 ( .A(x[752]), .B(y[752]), .Z(n38579) );
  IV U56981 ( .A(n38579), .Z(n42620) );
  IV U56982 ( .A(x[751]), .Z(n38580) );
  XOR U56983 ( .A(n38580), .B(y[751]), .Z(n42617) );
  XOR U56984 ( .A(x[750]), .B(y[750]), .Z(n38581) );
  IV U56985 ( .A(n38581), .Z(n42614) );
  IV U56986 ( .A(x[749]), .Z(n38582) );
  XOR U56987 ( .A(n38582), .B(y[749]), .Z(n39857) );
  XOR U56988 ( .A(x[748]), .B(y[748]), .Z(n39853) );
  XOR U56989 ( .A(x[747]), .B(y[747]), .Z(n42609) );
  XOR U56990 ( .A(x[746]), .B(y[746]), .Z(n42606) );
  XOR U56991 ( .A(x[745]), .B(y[745]), .Z(n42603) );
  XOR U56992 ( .A(x[744]), .B(y[744]), .Z(n42600) );
  XOR U56993 ( .A(x[743]), .B(y[743]), .Z(n42596) );
  XOR U56994 ( .A(x[742]), .B(y[742]), .Z(n42593) );
  XOR U56995 ( .A(x[741]), .B(y[741]), .Z(n39858) );
  XOR U56996 ( .A(x[740]), .B(y[740]), .Z(n42589) );
  XOR U56997 ( .A(x[739]), .B(y[739]), .Z(n42586) );
  IV U56998 ( .A(n42586), .Z(n45258) );
  XOR U56999 ( .A(x[738]), .B(y[738]), .Z(n39861) );
  XOR U57000 ( .A(x[737]), .B(y[737]), .Z(n42575) );
  XOR U57001 ( .A(x[736]), .B(y[736]), .Z(n39864) );
  XOR U57002 ( .A(x[735]), .B(y[735]), .Z(n42563) );
  XOR U57003 ( .A(x[734]), .B(y[734]), .Z(n42557) );
  XOR U57004 ( .A(x[733]), .B(y[733]), .Z(n42554) );
  XOR U57005 ( .A(x[732]), .B(y[732]), .Z(n39870) );
  XOR U57006 ( .A(x[731]), .B(y[731]), .Z(n39867) );
  XOR U57007 ( .A(x[730]), .B(y[730]), .Z(n42551) );
  XOR U57008 ( .A(x[729]), .B(y[729]), .Z(n42548) );
  XOR U57009 ( .A(x[728]), .B(y[728]), .Z(n42544) );
  XOR U57010 ( .A(x[727]), .B(y[727]), .Z(n42541) );
  XOR U57011 ( .A(x[726]), .B(y[726]), .Z(n42537) );
  XOR U57012 ( .A(x[725]), .B(y[725]), .Z(n42534) );
  XOR U57013 ( .A(x[724]), .B(y[724]), .Z(n39873) );
  XOR U57014 ( .A(x[723]), .B(y[723]), .Z(n39879) );
  XOR U57015 ( .A(x[722]), .B(y[722]), .Z(n39876) );
  XOR U57016 ( .A(x[721]), .B(y[721]), .Z(n39883) );
  XOR U57017 ( .A(x[720]), .B(y[720]), .Z(n42529) );
  XOR U57018 ( .A(x[719]), .B(y[719]), .Z(n42526) );
  XOR U57019 ( .A(x[718]), .B(y[718]), .Z(n39889) );
  XOR U57020 ( .A(x[717]), .B(y[717]), .Z(n39886) );
  XOR U57021 ( .A(x[716]), .B(y[716]), .Z(n42523) );
  XOR U57022 ( .A(x[715]), .B(y[715]), .Z(n42520) );
  XOR U57023 ( .A(x[714]), .B(y[714]), .Z(n42517) );
  XOR U57024 ( .A(x[713]), .B(y[713]), .Z(n42514) );
  XOR U57025 ( .A(x[712]), .B(y[712]), .Z(n42510) );
  XOR U57026 ( .A(x[711]), .B(y[711]), .Z(n42507) );
  XOR U57027 ( .A(x[710]), .B(y[710]), .Z(n42503) );
  XOR U57028 ( .A(x[709]), .B(y[709]), .Z(n42500) );
  XOR U57029 ( .A(x[708]), .B(y[708]), .Z(n42496) );
  XOR U57030 ( .A(x[707]), .B(y[707]), .Z(n42493) );
  XOR U57031 ( .A(x[706]), .B(y[706]), .Z(n39895) );
  XOR U57032 ( .A(x[705]), .B(y[705]), .Z(n39892) );
  XOR U57033 ( .A(x[704]), .B(y[704]), .Z(n42489) );
  XOR U57034 ( .A(x[703]), .B(y[703]), .Z(n42486) );
  XOR U57035 ( .A(x[702]), .B(y[702]), .Z(n39901) );
  XOR U57036 ( .A(x[701]), .B(y[701]), .Z(n39898) );
  XOR U57037 ( .A(x[700]), .B(y[700]), .Z(n39907) );
  XOR U57038 ( .A(x[699]), .B(y[699]), .Z(n39904) );
  XOR U57039 ( .A(x[698]), .B(y[698]), .Z(n39913) );
  XOR U57040 ( .A(x[697]), .B(y[697]), .Z(n39910) );
  XOR U57041 ( .A(x[696]), .B(y[696]), .Z(n39916) );
  XOR U57042 ( .A(x[695]), .B(y[695]), .Z(n42481) );
  XOR U57043 ( .A(x[694]), .B(y[694]), .Z(n42478) );
  XOR U57044 ( .A(x[693]), .B(y[693]), .Z(n39922) );
  XOR U57045 ( .A(x[692]), .B(y[692]), .Z(n39919) );
  XOR U57046 ( .A(x[691]), .B(y[691]), .Z(n39925) );
  XOR U57047 ( .A(x[690]), .B(y[690]), .Z(n42474) );
  XOR U57048 ( .A(x[689]), .B(y[689]), .Z(n42471) );
  XOR U57049 ( .A(x[688]), .B(y[688]), .Z(n42467) );
  XOR U57050 ( .A(x[687]), .B(y[687]), .Z(n42464) );
  XOR U57051 ( .A(x[686]), .B(y[686]), .Z(n42459) );
  XOR U57052 ( .A(x[685]), .B(y[685]), .Z(n42456) );
  XOR U57053 ( .A(x[684]), .B(y[684]), .Z(n39931) );
  XOR U57054 ( .A(x[683]), .B(y[683]), .Z(n39928) );
  XOR U57055 ( .A(x[682]), .B(y[682]), .Z(n39937) );
  XOR U57056 ( .A(x[681]), .B(y[681]), .Z(n39934) );
  XOR U57057 ( .A(x[680]), .B(y[680]), .Z(n42451) );
  XOR U57058 ( .A(x[679]), .B(y[679]), .Z(n42448) );
  XOR U57059 ( .A(x[678]), .B(y[678]), .Z(n39943) );
  XOR U57060 ( .A(x[677]), .B(y[677]), .Z(n39940) );
  XOR U57061 ( .A(x[676]), .B(y[676]), .Z(n39949) );
  XOR U57062 ( .A(x[675]), .B(y[675]), .Z(n39946) );
  XOR U57063 ( .A(x[674]), .B(y[674]), .Z(n39955) );
  XOR U57064 ( .A(x[673]), .B(y[673]), .Z(n39952) );
  XOR U57065 ( .A(x[672]), .B(y[672]), .Z(n39961) );
  XOR U57066 ( .A(x[671]), .B(y[671]), .Z(n39958) );
  XOR U57067 ( .A(x[670]), .B(y[670]), .Z(n39967) );
  XOR U57068 ( .A(x[669]), .B(y[669]), .Z(n39964) );
  XOR U57069 ( .A(x[668]), .B(y[668]), .Z(n42440) );
  XOR U57070 ( .A(x[667]), .B(y[667]), .Z(n42437) );
  XOR U57071 ( .A(x[666]), .B(y[666]), .Z(n42433) );
  XOR U57072 ( .A(x[665]), .B(y[665]), .Z(n42430) );
  XOR U57073 ( .A(x[664]), .B(y[664]), .Z(n39973) );
  XOR U57074 ( .A(x[663]), .B(y[663]), .Z(n39970) );
  XOR U57075 ( .A(x[662]), .B(y[662]), .Z(n39979) );
  XOR U57076 ( .A(x[661]), .B(y[661]), .Z(n39976) );
  XOR U57077 ( .A(x[660]), .B(y[660]), .Z(n42424) );
  XOR U57078 ( .A(x[659]), .B(y[659]), .Z(n42421) );
  XOR U57079 ( .A(x[658]), .B(y[658]), .Z(n42417) );
  XOR U57080 ( .A(x[657]), .B(y[657]), .Z(n42414) );
  XOR U57081 ( .A(x[656]), .B(y[656]), .Z(n42411) );
  XOR U57082 ( .A(x[655]), .B(y[655]), .Z(n42408) );
  XOR U57083 ( .A(x[654]), .B(y[654]), .Z(n42404) );
  XOR U57084 ( .A(x[653]), .B(y[653]), .Z(n42401) );
  XOR U57085 ( .A(x[652]), .B(y[652]), .Z(n39982) );
  XOR U57086 ( .A(x[651]), .B(y[651]), .Z(n39988) );
  XOR U57087 ( .A(x[650]), .B(y[650]), .Z(n39985) );
  XOR U57088 ( .A(x[649]), .B(y[649]), .Z(n39991) );
  XOR U57089 ( .A(x[648]), .B(y[648]), .Z(n39998) );
  XOR U57090 ( .A(x[647]), .B(y[647]), .Z(n39995) );
  XOR U57091 ( .A(x[646]), .B(y[646]), .Z(n42395) );
  XOR U57092 ( .A(x[645]), .B(y[645]), .Z(n42392) );
  XOR U57093 ( .A(x[644]), .B(y[644]), .Z(n42388) );
  XOR U57094 ( .A(x[643]), .B(y[643]), .Z(n42385) );
  XOR U57095 ( .A(x[642]), .B(y[642]), .Z(n40004) );
  XOR U57096 ( .A(x[641]), .B(y[641]), .Z(n40001) );
  XOR U57097 ( .A(x[640]), .B(y[640]), .Z(n42381) );
  XOR U57098 ( .A(x[639]), .B(y[639]), .Z(n42378) );
  XOR U57099 ( .A(x[638]), .B(y[638]), .Z(n40007) );
  XOR U57100 ( .A(x[637]), .B(y[637]), .Z(n40014) );
  XOR U57101 ( .A(x[636]), .B(y[636]), .Z(n40011) );
  XOR U57102 ( .A(x[635]), .B(y[635]), .Z(n40017) );
  XOR U57103 ( .A(x[634]), .B(y[634]), .Z(n40023) );
  XOR U57104 ( .A(x[633]), .B(y[633]), .Z(n40020) );
  XOR U57105 ( .A(x[632]), .B(y[632]), .Z(n42373) );
  XOR U57106 ( .A(x[631]), .B(y[631]), .Z(n42370) );
  XOR U57107 ( .A(x[630]), .B(y[630]), .Z(n40026) );
  XOR U57108 ( .A(x[629]), .B(y[629]), .Z(n42366) );
  XOR U57109 ( .A(x[628]), .B(y[628]), .Z(n42363) );
  XOR U57110 ( .A(x[627]), .B(y[627]), .Z(n40032) );
  XOR U57111 ( .A(x[626]), .B(y[626]), .Z(n40029) );
  XOR U57112 ( .A(x[625]), .B(y[625]), .Z(n40035) );
  XOR U57113 ( .A(x[624]), .B(y[624]), .Z(n40041) );
  XOR U57114 ( .A(x[623]), .B(y[623]), .Z(n40038) );
  XOR U57115 ( .A(x[622]), .B(y[622]), .Z(n40047) );
  XOR U57116 ( .A(x[621]), .B(y[621]), .Z(n40044) );
  XOR U57117 ( .A(x[620]), .B(y[620]), .Z(n42341) );
  XOR U57118 ( .A(x[619]), .B(y[619]), .Z(n42338) );
  XOR U57119 ( .A(x[618]), .B(y[618]), .Z(n42334) );
  XOR U57120 ( .A(x[617]), .B(y[617]), .Z(n42331) );
  XOR U57121 ( .A(x[616]), .B(y[616]), .Z(n42327) );
  XOR U57122 ( .A(x[615]), .B(y[615]), .Z(n42324) );
  XOR U57123 ( .A(x[614]), .B(y[614]), .Z(n42320) );
  XOR U57124 ( .A(x[613]), .B(y[613]), .Z(n42317) );
  XOR U57125 ( .A(x[612]), .B(y[612]), .Z(n40050) );
  XOR U57126 ( .A(x[611]), .B(y[611]), .Z(n42313) );
  XOR U57127 ( .A(x[610]), .B(y[610]), .Z(n42310) );
  XOR U57128 ( .A(x[609]), .B(y[609]), .Z(n42306) );
  XOR U57129 ( .A(x[608]), .B(y[608]), .Z(n42303) );
  XOR U57130 ( .A(x[607]), .B(y[607]), .Z(n40053) );
  XOR U57131 ( .A(x[606]), .B(y[606]), .Z(n42299) );
  XOR U57132 ( .A(x[605]), .B(y[605]), .Z(n42296) );
  XOR U57133 ( .A(x[604]), .B(y[604]), .Z(n42292) );
  XOR U57134 ( .A(x[603]), .B(y[603]), .Z(n42289) );
  XOR U57135 ( .A(x[602]), .B(y[602]), .Z(n40056) );
  XOR U57136 ( .A(x[601]), .B(y[601]), .Z(n42284) );
  XOR U57137 ( .A(x[600]), .B(y[600]), .Z(n42281) );
  XOR U57138 ( .A(x[599]), .B(y[599]), .Z(n42278) );
  XOR U57139 ( .A(x[598]), .B(y[598]), .Z(n42275) );
  XOR U57140 ( .A(x[597]), .B(y[597]), .Z(n42262) );
  XOR U57141 ( .A(x[596]), .B(y[596]), .Z(n40059) );
  XOR U57142 ( .A(x[595]), .B(y[595]), .Z(n42265) );
  XOR U57143 ( .A(x[594]), .B(y[594]), .Z(n40063) );
  XOR U57144 ( .A(x[593]), .B(y[593]), .Z(n42257) );
  XOR U57145 ( .A(x[592]), .B(y[592]), .Z(n42254) );
  XOR U57146 ( .A(x[591]), .B(y[591]), .Z(n40066) );
  XOR U57147 ( .A(x[590]), .B(y[590]), .Z(n42250) );
  XOR U57148 ( .A(x[589]), .B(y[589]), .Z(n42247) );
  XOR U57149 ( .A(x[588]), .B(y[588]), .Z(n42243) );
  XOR U57150 ( .A(x[587]), .B(y[587]), .Z(n42240) );
  XOR U57151 ( .A(x[586]), .B(y[586]), .Z(n40069) );
  XOR U57152 ( .A(x[585]), .B(y[585]), .Z(n40075) );
  XOR U57153 ( .A(x[584]), .B(y[584]), .Z(n40072) );
  XOR U57154 ( .A(x[583]), .B(y[583]), .Z(n40078) );
  XOR U57155 ( .A(x[582]), .B(y[582]), .Z(n42233) );
  XOR U57156 ( .A(x[581]), .B(y[581]), .Z(n40081) );
  XOR U57157 ( .A(x[580]), .B(y[580]), .Z(n45507) );
  XOR U57158 ( .A(x[579]), .B(y[579]), .Z(n40086) );
  XOR U57159 ( .A(x[578]), .B(y[578]), .Z(n40090) );
  XOR U57160 ( .A(x[577]), .B(y[577]), .Z(n40093) );
  XOR U57161 ( .A(x[576]), .B(y[576]), .Z(n42222) );
  XOR U57162 ( .A(x[575]), .B(y[575]), .Z(n40096) );
  XOR U57163 ( .A(x[574]), .B(y[574]), .Z(n42216) );
  XOR U57164 ( .A(x[573]), .B(y[573]), .Z(n42213) );
  XOR U57165 ( .A(x[572]), .B(y[572]), .Z(n40102) );
  XOR U57166 ( .A(x[571]), .B(y[571]), .Z(n40099) );
  XOR U57167 ( .A(x[570]), .B(y[570]), .Z(n38583) );
  IV U57168 ( .A(n38583), .Z(n40109) );
  IV U57169 ( .A(x[569]), .Z(n38584) );
  XOR U57170 ( .A(n38584), .B(y[569]), .Z(n40106) );
  XOR U57171 ( .A(x[568]), .B(y[568]), .Z(n40113) );
  XOR U57172 ( .A(x[567]), .B(y[567]), .Z(n40110) );
  XOR U57173 ( .A(x[566]), .B(y[566]), .Z(n40116) );
  XOR U57174 ( .A(x[565]), .B(y[565]), .Z(n42206) );
  XOR U57175 ( .A(x[564]), .B(y[564]), .Z(n42203) );
  XOR U57176 ( .A(x[563]), .B(y[563]), .Z(n40122) );
  XOR U57177 ( .A(x[562]), .B(y[562]), .Z(n40119) );
  XOR U57178 ( .A(x[561]), .B(y[561]), .Z(n40128) );
  XOR U57179 ( .A(x[560]), .B(y[560]), .Z(n40125) );
  XOR U57180 ( .A(x[559]), .B(y[559]), .Z(n40132) );
  XOR U57181 ( .A(x[558]), .B(y[558]), .Z(n38585) );
  IV U57182 ( .A(n38585), .Z(n42199) );
  IV U57183 ( .A(x[557]), .Z(n38586) );
  XOR U57184 ( .A(n38586), .B(y[557]), .Z(n42196) );
  XOR U57185 ( .A(x[556]), .B(y[556]), .Z(n42193) );
  XOR U57186 ( .A(x[555]), .B(y[555]), .Z(n42190) );
  XOR U57187 ( .A(x[554]), .B(y[554]), .Z(n40138) );
  XOR U57188 ( .A(x[553]), .B(y[553]), .Z(n40135) );
  XOR U57189 ( .A(x[552]), .B(y[552]), .Z(n42185) );
  XOR U57190 ( .A(x[551]), .B(y[551]), .Z(n42182) );
  XOR U57191 ( .A(x[550]), .B(y[550]), .Z(n42178) );
  XOR U57192 ( .A(x[549]), .B(y[549]), .Z(n42175) );
  XOR U57193 ( .A(x[548]), .B(y[548]), .Z(n40144) );
  XOR U57194 ( .A(x[547]), .B(y[547]), .Z(n40141) );
  XOR U57195 ( .A(x[546]), .B(y[546]), .Z(n38587) );
  IV U57196 ( .A(n38587), .Z(n40151) );
  IV U57197 ( .A(x[545]), .Z(n38588) );
  XOR U57198 ( .A(n38588), .B(y[545]), .Z(n40147) );
  XOR U57199 ( .A(x[544]), .B(y[544]), .Z(n40152) );
  XOR U57200 ( .A(x[543]), .B(y[543]), .Z(n42161) );
  XOR U57201 ( .A(x[542]), .B(y[542]), .Z(n40155) );
  XOR U57202 ( .A(x[541]), .B(y[541]), .Z(n42153) );
  XOR U57203 ( .A(x[540]), .B(y[540]), .Z(n40158) );
  XOR U57204 ( .A(x[539]), .B(y[539]), .Z(n40164) );
  XOR U57205 ( .A(x[538]), .B(y[538]), .Z(n40161) );
  XOR U57206 ( .A(x[537]), .B(y[537]), .Z(n40170) );
  XOR U57207 ( .A(x[536]), .B(y[536]), .Z(n40167) );
  XOR U57208 ( .A(x[535]), .B(y[535]), .Z(n40173) );
  XOR U57209 ( .A(x[534]), .B(y[534]), .Z(n38589) );
  IV U57210 ( .A(n38589), .Z(n42145) );
  IV U57211 ( .A(x[533]), .Z(n38590) );
  XOR U57212 ( .A(n38590), .B(y[533]), .Z(n42142) );
  XOR U57213 ( .A(x[532]), .B(y[532]), .Z(n40179) );
  XOR U57214 ( .A(x[531]), .B(y[531]), .Z(n40176) );
  XOR U57215 ( .A(x[530]), .B(y[530]), .Z(n40182) );
  XOR U57216 ( .A(x[529]), .B(y[529]), .Z(n42131) );
  XOR U57217 ( .A(x[528]), .B(y[528]), .Z(n40185) );
  XOR U57218 ( .A(x[527]), .B(y[527]), .Z(n42118) );
  XOR U57219 ( .A(x[526]), .B(y[526]), .Z(n40188) );
  XOR U57220 ( .A(x[525]), .B(y[525]), .Z(n42108) );
  XOR U57221 ( .A(x[524]), .B(y[524]), .Z(n42105) );
  XOR U57222 ( .A(x[523]), .B(y[523]), .Z(n42100) );
  XOR U57223 ( .A(x[522]), .B(y[522]), .Z(n42097) );
  XOR U57224 ( .A(x[521]), .B(y[521]), .Z(n38591) );
  IV U57225 ( .A(n38591), .Z(n40192) );
  IV U57226 ( .A(x[520]), .Z(n38592) );
  XOR U57227 ( .A(n38592), .B(y[520]), .Z(n40198) );
  XOR U57228 ( .A(x[519]), .B(y[519]), .Z(n40194) );
  XOR U57229 ( .A(x[518]), .B(y[518]), .Z(n40202) );
  XOR U57230 ( .A(x[517]), .B(y[517]), .Z(n40199) );
  XOR U57231 ( .A(x[516]), .B(y[516]), .Z(n40206) );
  XOR U57232 ( .A(x[515]), .B(y[515]), .Z(n42093) );
  XOR U57233 ( .A(x[514]), .B(y[514]), .Z(n42090) );
  XOR U57234 ( .A(x[513]), .B(y[513]), .Z(n42086) );
  XOR U57235 ( .A(x[512]), .B(y[512]), .Z(n42083) );
  XOR U57236 ( .A(x[511]), .B(y[511]), .Z(n40209) );
  XOR U57237 ( .A(x[510]), .B(y[510]), .Z(n42078) );
  XOR U57238 ( .A(x[509]), .B(y[509]), .Z(n42075) );
  XOR U57239 ( .A(x[508]), .B(y[508]), .Z(n42071) );
  XOR U57240 ( .A(x[507]), .B(y[507]), .Z(n42068) );
  XOR U57241 ( .A(x[506]), .B(y[506]), .Z(n40215) );
  XOR U57242 ( .A(x[505]), .B(y[505]), .Z(n40212) );
  XOR U57243 ( .A(x[504]), .B(y[504]), .Z(n40218) );
  XOR U57244 ( .A(x[503]), .B(y[503]), .Z(n42062) );
  XOR U57245 ( .A(x[502]), .B(y[502]), .Z(n42059) );
  XOR U57246 ( .A(x[501]), .B(y[501]), .Z(n40224) );
  XOR U57247 ( .A(x[500]), .B(y[500]), .Z(n40221) );
  XOR U57248 ( .A(x[499]), .B(y[499]), .Z(n40227) );
  XOR U57249 ( .A(x[498]), .B(y[498]), .Z(n42052) );
  XOR U57250 ( .A(x[497]), .B(y[497]), .Z(n40230) );
  XOR U57251 ( .A(x[496]), .B(y[496]), .Z(n42046) );
  XOR U57252 ( .A(x[495]), .B(y[495]), .Z(n42043) );
  XOR U57253 ( .A(x[494]), .B(y[494]), .Z(n40233) );
  XOR U57254 ( .A(x[493]), .B(y[493]), .Z(n42032) );
  XOR U57255 ( .A(x[492]), .B(y[492]), .Z(n40239) );
  XOR U57256 ( .A(x[491]), .B(y[491]), .Z(n40236) );
  XOR U57257 ( .A(x[490]), .B(y[490]), .Z(n42025) );
  XOR U57258 ( .A(x[489]), .B(y[489]), .Z(n42022) );
  XOR U57259 ( .A(x[488]), .B(y[488]), .Z(n42018) );
  XOR U57260 ( .A(x[487]), .B(y[487]), .Z(n42015) );
  XOR U57261 ( .A(x[486]), .B(y[486]), .Z(n40245) );
  XOR U57262 ( .A(x[485]), .B(y[485]), .Z(n40242) );
  XOR U57263 ( .A(x[484]), .B(y[484]), .Z(n40248) );
  XOR U57264 ( .A(x[483]), .B(y[483]), .Z(n42005) );
  XOR U57265 ( .A(x[482]), .B(y[482]), .Z(n42002) );
  XOR U57266 ( .A(x[481]), .B(y[481]), .Z(n41997) );
  XOR U57267 ( .A(x[480]), .B(y[480]), .Z(n41994) );
  XOR U57268 ( .A(x[479]), .B(y[479]), .Z(n40251) );
  XOR U57269 ( .A(x[478]), .B(y[478]), .Z(n41991) );
  XOR U57270 ( .A(x[477]), .B(y[477]), .Z(n41988) );
  XOR U57271 ( .A(x[476]), .B(y[476]), .Z(n41984) );
  XOR U57272 ( .A(x[475]), .B(y[475]), .Z(n41981) );
  XOR U57273 ( .A(x[474]), .B(y[474]), .Z(n40254) );
  XOR U57274 ( .A(x[473]), .B(y[473]), .Z(n40261) );
  XOR U57275 ( .A(x[472]), .B(y[472]), .Z(n40258) );
  XOR U57276 ( .A(x[471]), .B(y[471]), .Z(n41977) );
  XOR U57277 ( .A(x[470]), .B(y[470]), .Z(n41974) );
  XOR U57278 ( .A(x[469]), .B(y[469]), .Z(n41970) );
  XOR U57279 ( .A(x[468]), .B(y[468]), .Z(n41967) );
  XOR U57280 ( .A(x[467]), .B(y[467]), .Z(n41963) );
  XOR U57281 ( .A(x[466]), .B(y[466]), .Z(n41960) );
  XOR U57282 ( .A(x[465]), .B(y[465]), .Z(n40267) );
  XOR U57283 ( .A(x[464]), .B(y[464]), .Z(n40264) );
  XOR U57284 ( .A(x[463]), .B(y[463]), .Z(n41956) );
  XOR U57285 ( .A(x[462]), .B(y[462]), .Z(n41953) );
  XOR U57286 ( .A(x[461]), .B(y[461]), .Z(n41950) );
  XOR U57287 ( .A(x[460]), .B(y[460]), .Z(n41947) );
  XOR U57288 ( .A(x[459]), .B(y[459]), .Z(n41943) );
  XOR U57289 ( .A(x[458]), .B(y[458]), .Z(n41940) );
  XOR U57290 ( .A(x[457]), .B(y[457]), .Z(n40271) );
  XOR U57291 ( .A(x[456]), .B(y[456]), .Z(n41934) );
  XOR U57292 ( .A(x[455]), .B(y[455]), .Z(n40274) );
  XOR U57293 ( .A(x[454]), .B(y[454]), .Z(n41927) );
  XOR U57294 ( .A(x[453]), .B(y[453]), .Z(n41924) );
  XOR U57295 ( .A(x[452]), .B(y[452]), .Z(n41920) );
  XOR U57296 ( .A(x[451]), .B(y[451]), .Z(n41917) );
  XOR U57297 ( .A(x[450]), .B(y[450]), .Z(n41913) );
  XOR U57298 ( .A(x[449]), .B(y[449]), .Z(n41910) );
  XOR U57299 ( .A(x[448]), .B(y[448]), .Z(n40277) );
  XOR U57300 ( .A(x[447]), .B(y[447]), .Z(n40284) );
  XOR U57301 ( .A(x[446]), .B(y[446]), .Z(n40281) );
  XOR U57302 ( .A(x[445]), .B(y[445]), .Z(n40287) );
  XOR U57303 ( .A(x[444]), .B(y[444]), .Z(n41904) );
  XOR U57304 ( .A(x[443]), .B(y[443]), .Z(n41901) );
  XOR U57305 ( .A(x[442]), .B(y[442]), .Z(n40293) );
  XOR U57306 ( .A(x[441]), .B(y[441]), .Z(n40290) );
  XOR U57307 ( .A(x[440]), .B(y[440]), .Z(n41897) );
  XOR U57308 ( .A(x[439]), .B(y[439]), .Z(n41894) );
  XOR U57309 ( .A(x[436]), .B(y[436]), .Z(n40303) );
  XOR U57310 ( .A(x[435]), .B(y[435]), .Z(n40300) );
  XOR U57311 ( .A(x[434]), .B(y[434]), .Z(n40309) );
  XOR U57312 ( .A(x[433]), .B(y[433]), .Z(n40306) );
  XOR U57313 ( .A(x[432]), .B(y[432]), .Z(n41890) );
  XOR U57314 ( .A(x[431]), .B(y[431]), .Z(n41887) );
  XOR U57315 ( .A(x[430]), .B(y[430]), .Z(n41883) );
  XOR U57316 ( .A(x[429]), .B(y[429]), .Z(n41880) );
  XOR U57317 ( .A(x[428]), .B(y[428]), .Z(n41876) );
  XOR U57318 ( .A(x[427]), .B(y[427]), .Z(n41873) );
  XOR U57319 ( .A(x[426]), .B(y[426]), .Z(n40315) );
  XOR U57320 ( .A(x[425]), .B(y[425]), .Z(n40312) );
  XOR U57321 ( .A(x[424]), .B(y[424]), .Z(n41868) );
  XOR U57322 ( .A(x[423]), .B(y[423]), .Z(n41865) );
  XOR U57323 ( .A(x[422]), .B(y[422]), .Z(n41862) );
  XOR U57324 ( .A(x[421]), .B(y[421]), .Z(n41859) );
  XOR U57325 ( .A(x[420]), .B(y[420]), .Z(n41855) );
  XOR U57326 ( .A(x[419]), .B(y[419]), .Z(n41852) );
  XOR U57327 ( .A(x[418]), .B(y[418]), .Z(n40318) );
  XOR U57328 ( .A(x[417]), .B(y[417]), .Z(n40325) );
  XOR U57329 ( .A(x[416]), .B(y[416]), .Z(n40322) );
  XOR U57330 ( .A(x[415]), .B(y[415]), .Z(n40328) );
  XOR U57331 ( .A(x[414]), .B(y[414]), .Z(n40334) );
  XOR U57332 ( .A(x[413]), .B(y[413]), .Z(n40331) );
  XOR U57333 ( .A(x[412]), .B(y[412]), .Z(n40340) );
  XOR U57334 ( .A(x[411]), .B(y[411]), .Z(n40337) );
  XOR U57335 ( .A(x[410]), .B(y[410]), .Z(n40346) );
  XOR U57336 ( .A(x[409]), .B(y[409]), .Z(n40343) );
  XOR U57337 ( .A(x[408]), .B(y[408]), .Z(n41847) );
  XOR U57338 ( .A(x[407]), .B(y[407]), .Z(n41844) );
  XOR U57339 ( .A(x[406]), .B(y[406]), .Z(n40349) );
  XOR U57340 ( .A(x[405]), .B(y[405]), .Z(n41829) );
  XOR U57341 ( .A(x[404]), .B(y[404]), .Z(n40353) );
  XOR U57342 ( .A(x[403]), .B(y[403]), .Z(n41832) );
  XOR U57343 ( .A(x[402]), .B(y[402]), .Z(n40360) );
  XOR U57344 ( .A(x[401]), .B(y[401]), .Z(n40357) );
  XOR U57345 ( .A(x[400]), .B(y[400]), .Z(n40366) );
  XOR U57346 ( .A(x[399]), .B(y[399]), .Z(n40363) );
  XOR U57347 ( .A(x[398]), .B(y[398]), .Z(n40372) );
  XOR U57348 ( .A(x[397]), .B(y[397]), .Z(n40369) );
  XOR U57349 ( .A(x[396]), .B(y[396]), .Z(n41821) );
  XOR U57350 ( .A(x[395]), .B(y[395]), .Z(n41818) );
  XOR U57351 ( .A(x[394]), .B(y[394]), .Z(n40378) );
  XOR U57352 ( .A(x[393]), .B(y[393]), .Z(n40375) );
  XOR U57353 ( .A(x[392]), .B(y[392]), .Z(n40384) );
  XOR U57354 ( .A(x[391]), .B(y[391]), .Z(n40381) );
  XOR U57355 ( .A(x[390]), .B(y[390]), .Z(n40387) );
  XOR U57356 ( .A(x[389]), .B(y[389]), .Z(n41812) );
  XOR U57357 ( .A(x[388]), .B(y[388]), .Z(n41809) );
  XOR U57358 ( .A(x[387]), .B(y[387]), .Z(n40390) );
  XOR U57359 ( .A(x[386]), .B(y[386]), .Z(n40396) );
  XOR U57360 ( .A(x[385]), .B(y[385]), .Z(n40393) );
  XOR U57361 ( .A(x[384]), .B(y[384]), .Z(n41804) );
  XOR U57362 ( .A(x[383]), .B(y[383]), .Z(n41801) );
  XOR U57363 ( .A(x[382]), .B(y[382]), .Z(n40402) );
  XOR U57364 ( .A(x[381]), .B(y[381]), .Z(n40399) );
  XOR U57365 ( .A(x[380]), .B(y[380]), .Z(n40408) );
  XOR U57366 ( .A(x[379]), .B(y[379]), .Z(n40405) );
  XOR U57367 ( .A(x[378]), .B(y[378]), .Z(n46826) );
  XOR U57368 ( .A(x[377]), .B(y[377]), .Z(n40414) );
  XOR U57369 ( .A(x[376]), .B(y[376]), .Z(n40420) );
  XOR U57370 ( .A(x[375]), .B(y[375]), .Z(n40417) );
  XOR U57371 ( .A(x[374]), .B(y[374]), .Z(n40424) );
  XOR U57372 ( .A(x[373]), .B(y[373]), .Z(n40430) );
  XOR U57373 ( .A(x[372]), .B(y[372]), .Z(n40427) );
  XOR U57374 ( .A(x[371]), .B(y[371]), .Z(n40436) );
  XOR U57375 ( .A(x[370]), .B(y[370]), .Z(n40433) );
  XOR U57376 ( .A(x[369]), .B(y[369]), .Z(n41794) );
  XOR U57377 ( .A(x[368]), .B(y[368]), .Z(n41791) );
  XOR U57378 ( .A(x[367]), .B(y[367]), .Z(n41787) );
  XOR U57379 ( .A(x[366]), .B(y[366]), .Z(n41784) );
  XOR U57380 ( .A(x[365]), .B(y[365]), .Z(n41780) );
  XOR U57381 ( .A(x[364]), .B(y[364]), .Z(n38593) );
  IV U57382 ( .A(n38593), .Z(n41778) );
  IV U57383 ( .A(x[363]), .Z(n38594) );
  XOR U57384 ( .A(n38594), .B(y[363]), .Z(n40444) );
  XOR U57385 ( .A(x[362]), .B(y[362]), .Z(n40440) );
  XOR U57386 ( .A(x[361]), .B(y[361]), .Z(n41772) );
  XOR U57387 ( .A(x[360]), .B(y[360]), .Z(n38595) );
  IV U57388 ( .A(n38595), .Z(n41771) );
  IV U57389 ( .A(x[359]), .Z(n38596) );
  XOR U57390 ( .A(n38596), .B(y[359]), .Z(n40449) );
  XOR U57391 ( .A(x[358]), .B(y[358]), .Z(n40445) );
  XOR U57392 ( .A(x[357]), .B(y[357]), .Z(n40453) );
  XOR U57393 ( .A(x[356]), .B(y[356]), .Z(n38597) );
  IV U57394 ( .A(n38597), .Z(n40451) );
  IV U57395 ( .A(x[355]), .Z(n38598) );
  XOR U57396 ( .A(n38598), .B(y[355]), .Z(n40459) );
  XOR U57397 ( .A(x[354]), .B(y[354]), .Z(n40456) );
  XOR U57398 ( .A(x[353]), .B(y[353]), .Z(n40461) );
  XOR U57399 ( .A(x[352]), .B(y[352]), .Z(n38599) );
  IV U57400 ( .A(n38599), .Z(n41764) );
  IV U57401 ( .A(x[351]), .Z(n38600) );
  XOR U57402 ( .A(n38600), .B(y[351]), .Z(n41761) );
  XOR U57403 ( .A(x[350]), .B(y[350]), .Z(n38601) );
  IV U57404 ( .A(n38601), .Z(n40468) );
  IV U57405 ( .A(x[349]), .Z(n38602) );
  XOR U57406 ( .A(n38602), .B(y[349]), .Z(n40465) );
  XOR U57407 ( .A(x[348]), .B(y[348]), .Z(n41757) );
  XOR U57408 ( .A(x[347]), .B(y[347]), .Z(n41754) );
  XOR U57409 ( .A(x[346]), .B(y[346]), .Z(n40473) );
  XOR U57410 ( .A(x[345]), .B(y[345]), .Z(n40470) );
  XOR U57411 ( .A(x[344]), .B(y[344]), .Z(n41750) );
  XOR U57412 ( .A(x[343]), .B(y[343]), .Z(n41747) );
  XOR U57413 ( .A(x[342]), .B(y[342]), .Z(n40479) );
  XOR U57414 ( .A(x[341]), .B(y[341]), .Z(n40476) );
  XOR U57415 ( .A(x[340]), .B(y[340]), .Z(n41744) );
  XOR U57416 ( .A(x[339]), .B(y[339]), .Z(n41741) );
  XOR U57417 ( .A(x[338]), .B(y[338]), .Z(n41738) );
  XOR U57418 ( .A(x[337]), .B(y[337]), .Z(n57399) );
  XOR U57419 ( .A(x[336]), .B(y[336]), .Z(n40485) );
  XOR U57420 ( .A(x[335]), .B(y[335]), .Z(n40482) );
  XOR U57421 ( .A(x[334]), .B(y[334]), .Z(n40492) );
  XOR U57422 ( .A(x[333]), .B(y[333]), .Z(n40489) );
  XOR U57423 ( .A(x[332]), .B(y[332]), .Z(n41731) );
  XOR U57424 ( .A(x[331]), .B(y[331]), .Z(n41728) );
  XOR U57425 ( .A(x[330]), .B(y[330]), .Z(n41724) );
  XOR U57426 ( .A(x[329]), .B(y[329]), .Z(n41721) );
  XOR U57427 ( .A(x[328]), .B(y[328]), .Z(n38603) );
  IV U57428 ( .A(n38603), .Z(n41718) );
  IV U57429 ( .A(x[327]), .Z(n38604) );
  XOR U57430 ( .A(n38604), .B(y[327]), .Z(n41716) );
  XOR U57431 ( .A(x[326]), .B(y[326]), .Z(n41701) );
  XOR U57432 ( .A(x[325]), .B(y[325]), .Z(n41698) );
  XOR U57433 ( .A(x[324]), .B(y[324]), .Z(n40498) );
  XOR U57434 ( .A(x[323]), .B(y[323]), .Z(n40495) );
  XOR U57435 ( .A(x[322]), .B(y[322]), .Z(n40504) );
  XOR U57436 ( .A(x[321]), .B(y[321]), .Z(n40501) );
  XOR U57437 ( .A(x[320]), .B(y[320]), .Z(n40510) );
  XOR U57438 ( .A(x[319]), .B(y[319]), .Z(n40507) );
  XOR U57439 ( .A(x[318]), .B(y[318]), .Z(n41693) );
  XOR U57440 ( .A(x[317]), .B(y[317]), .Z(n41690) );
  XOR U57441 ( .A(x[316]), .B(y[316]), .Z(n38605) );
  IV U57442 ( .A(n38605), .Z(n41688) );
  IV U57443 ( .A(x[315]), .Z(n38606) );
  XOR U57444 ( .A(n38606), .B(y[315]), .Z(n41685) );
  XOR U57445 ( .A(x[314]), .B(y[314]), .Z(n41681) );
  XOR U57446 ( .A(x[313]), .B(y[313]), .Z(n41678) );
  XOR U57447 ( .A(x[312]), .B(y[312]), .Z(n41674) );
  XOR U57448 ( .A(x[311]), .B(y[311]), .Z(n41671) );
  XOR U57449 ( .A(x[310]), .B(y[310]), .Z(n41667) );
  XOR U57450 ( .A(x[309]), .B(y[309]), .Z(n41664) );
  XOR U57451 ( .A(x[308]), .B(y[308]), .Z(n41653) );
  XOR U57452 ( .A(x[307]), .B(y[307]), .Z(n41649) );
  XOR U57453 ( .A(x[306]), .B(y[306]), .Z(n41656) );
  XOR U57454 ( .A(x[305]), .B(y[305]), .Z(n41644) );
  XOR U57455 ( .A(x[304]), .B(y[304]), .Z(n38607) );
  IV U57456 ( .A(n38607), .Z(n41642) );
  IV U57457 ( .A(x[303]), .Z(n38608) );
  XOR U57458 ( .A(n38608), .B(y[303]), .Z(n40514) );
  XOR U57459 ( .A(x[302]), .B(y[302]), .Z(n40518) );
  XOR U57460 ( .A(x[301]), .B(y[301]), .Z(n40515) );
  XOR U57461 ( .A(x[300]), .B(y[300]), .Z(n41638) );
  XOR U57462 ( .A(x[299]), .B(y[299]), .Z(n41635) );
  XOR U57463 ( .A(x[298]), .B(y[298]), .Z(n40521) );
  XOR U57464 ( .A(x[297]), .B(y[297]), .Z(n40528) );
  XOR U57465 ( .A(x[296]), .B(y[296]), .Z(n40525) );
  XOR U57466 ( .A(x[295]), .B(y[295]), .Z(n40534) );
  XOR U57467 ( .A(x[294]), .B(y[294]), .Z(n40531) );
  XOR U57468 ( .A(x[293]), .B(y[293]), .Z(n40540) );
  XOR U57469 ( .A(x[292]), .B(y[292]), .Z(n38609) );
  IV U57470 ( .A(n38609), .Z(n40538) );
  IV U57471 ( .A(x[291]), .Z(n38610) );
  XOR U57472 ( .A(n38610), .B(y[291]), .Z(n41632) );
  XOR U57473 ( .A(x[290]), .B(y[290]), .Z(n41629) );
  XOR U57474 ( .A(x[289]), .B(y[289]), .Z(n40546) );
  XOR U57475 ( .A(x[288]), .B(y[288]), .Z(n40543) );
  XOR U57476 ( .A(x[287]), .B(y[287]), .Z(n40552) );
  XOR U57477 ( .A(x[286]), .B(y[286]), .Z(n40549) );
  XOR U57478 ( .A(x[285]), .B(y[285]), .Z(n41625) );
  XOR U57479 ( .A(x[284]), .B(y[284]), .Z(n41622) );
  XOR U57480 ( .A(x[283]), .B(y[283]), .Z(n41619) );
  XOR U57481 ( .A(x[282]), .B(y[282]), .Z(n41616) );
  XOR U57482 ( .A(x[281]), .B(y[281]), .Z(n40555) );
  XOR U57483 ( .A(x[280]), .B(y[280]), .Z(n41608) );
  XOR U57484 ( .A(x[279]), .B(y[279]), .Z(n41605) );
  XOR U57485 ( .A(x[278]), .B(y[278]), .Z(n41601) );
  XOR U57486 ( .A(x[277]), .B(y[277]), .Z(n41598) );
  XOR U57487 ( .A(x[276]), .B(y[276]), .Z(n41594) );
  XOR U57488 ( .A(x[275]), .B(y[275]), .Z(n41591) );
  XOR U57489 ( .A(x[272]), .B(y[272]), .Z(n41588) );
  XOR U57490 ( .A(x[271]), .B(y[271]), .Z(n41585) );
  XOR U57491 ( .A(x[270]), .B(y[270]), .Z(n41581) );
  XOR U57492 ( .A(x[269]), .B(y[269]), .Z(n41578) );
  XOR U57493 ( .A(x[268]), .B(y[268]), .Z(n40563) );
  XOR U57494 ( .A(x[267]), .B(y[267]), .Z(n41573) );
  XOR U57495 ( .A(x[266]), .B(y[266]), .Z(n41570) );
  XOR U57496 ( .A(x[265]), .B(y[265]), .Z(n40566) );
  XOR U57497 ( .A(x[264]), .B(y[264]), .Z(n41566) );
  XOR U57498 ( .A(x[263]), .B(y[263]), .Z(n41563) );
  XOR U57499 ( .A(x[262]), .B(y[262]), .Z(n40572) );
  XOR U57500 ( .A(x[261]), .B(y[261]), .Z(n40569) );
  XOR U57501 ( .A(x[260]), .B(y[260]), .Z(n41560) );
  XOR U57502 ( .A(x[259]), .B(y[259]), .Z(n41557) );
  XOR U57503 ( .A(x[258]), .B(y[258]), .Z(n40578) );
  XOR U57504 ( .A(x[257]), .B(y[257]), .Z(n40575) );
  XOR U57505 ( .A(x[256]), .B(y[256]), .Z(n41553) );
  XOR U57506 ( .A(x[255]), .B(y[255]), .Z(n41550) );
  XOR U57507 ( .A(x[254]), .B(y[254]), .Z(n40582) );
  XOR U57508 ( .A(x[253]), .B(y[253]), .Z(n40589) );
  XOR U57509 ( .A(x[252]), .B(y[252]), .Z(n40586) );
  XOR U57510 ( .A(x[251]), .B(y[251]), .Z(n40592) );
  XOR U57511 ( .A(x[250]), .B(y[250]), .Z(n41545) );
  XOR U57512 ( .A(x[249]), .B(y[249]), .Z(n41542) );
  XOR U57513 ( .A(x[248]), .B(y[248]), .Z(n40598) );
  XOR U57514 ( .A(x[247]), .B(y[247]), .Z(n40595) );
  XOR U57515 ( .A(x[246]), .B(y[246]), .Z(n56527) );
  XOR U57516 ( .A(x[245]), .B(y[245]), .Z(n40602) );
  XOR U57517 ( .A(x[244]), .B(y[244]), .Z(n38611) );
  IV U57518 ( .A(n38611), .Z(n41540) );
  XOR U57519 ( .A(x[243]), .B(y[243]), .Z(n41536) );
  XOR U57520 ( .A(x[242]), .B(y[242]), .Z(n51315) );
  XOR U57521 ( .A(x[241]), .B(y[241]), .Z(n41531) );
  IV U57522 ( .A(n41531), .Z(n41533) );
  XOR U57523 ( .A(x[240]), .B(y[240]), .Z(n38612) );
  IV U57524 ( .A(n38612), .Z(n40610) );
  IV U57525 ( .A(x[239]), .Z(n38613) );
  XOR U57526 ( .A(n38613), .B(y[239]), .Z(n40608) );
  XOR U57527 ( .A(x[238]), .B(y[238]), .Z(n41526) );
  XOR U57528 ( .A(x[237]), .B(y[237]), .Z(n41523) );
  XOR U57529 ( .A(x[236]), .B(y[236]), .Z(n40612) );
  XOR U57530 ( .A(x[235]), .B(y[235]), .Z(n40619) );
  XOR U57531 ( .A(x[234]), .B(y[234]), .Z(n40616) );
  XOR U57532 ( .A(x[233]), .B(y[233]), .Z(n41520) );
  XOR U57533 ( .A(x[232]), .B(y[232]), .Z(n41517) );
  XOR U57534 ( .A(x[231]), .B(y[231]), .Z(n40625) );
  XOR U57535 ( .A(x[230]), .B(y[230]), .Z(n40622) );
  XOR U57536 ( .A(x[229]), .B(y[229]), .Z(n40628) );
  XOR U57537 ( .A(x[228]), .B(y[228]), .Z(n38614) );
  IV U57538 ( .A(n38614), .Z(n40635) );
  IV U57539 ( .A(x[227]), .Z(n38615) );
  XOR U57540 ( .A(n38615), .B(y[227]), .Z(n40633) );
  XOR U57541 ( .A(x[226]), .B(y[226]), .Z(n40641) );
  XOR U57542 ( .A(x[225]), .B(y[225]), .Z(n40638) );
  XOR U57543 ( .A(x[224]), .B(y[224]), .Z(n41512) );
  XOR U57544 ( .A(x[223]), .B(y[223]), .Z(n41509) );
  XOR U57545 ( .A(x[222]), .B(y[222]), .Z(n40647) );
  XOR U57546 ( .A(x[221]), .B(y[221]), .Z(n40644) );
  XOR U57547 ( .A(x[220]), .B(y[220]), .Z(n41506) );
  XOR U57548 ( .A(x[219]), .B(y[219]), .Z(n41503) );
  XOR U57549 ( .A(x[218]), .B(y[218]), .Z(n40653) );
  XOR U57550 ( .A(x[217]), .B(y[217]), .Z(n40650) );
  XOR U57551 ( .A(x[216]), .B(y[216]), .Z(n38616) );
  IV U57552 ( .A(n38616), .Z(n41489) );
  IV U57553 ( .A(x[215]), .Z(n38617) );
  XOR U57554 ( .A(n38617), .B(y[215]), .Z(n41486) );
  XOR U57555 ( .A(x[214]), .B(y[214]), .Z(n40656) );
  XOR U57556 ( .A(x[213]), .B(y[213]), .Z(n41475) );
  XOR U57557 ( .A(x[212]), .B(y[212]), .Z(n38618) );
  IV U57558 ( .A(n38618), .Z(n40660) );
  IV U57559 ( .A(x[211]), .Z(n38619) );
  XOR U57560 ( .A(n38619), .B(y[211]), .Z(n41468) );
  XOR U57561 ( .A(x[210]), .B(y[210]), .Z(n40662) );
  XOR U57562 ( .A(x[209]), .B(y[209]), .Z(n41462) );
  XOR U57563 ( .A(x[208]), .B(y[208]), .Z(n38620) );
  IV U57564 ( .A(n38620), .Z(n41461) );
  IV U57565 ( .A(x[207]), .Z(n38621) );
  XOR U57566 ( .A(n38621), .B(y[207]), .Z(n40666) );
  XOR U57567 ( .A(x[206]), .B(y[206]), .Z(n41453) );
  XOR U57568 ( .A(x[205]), .B(y[205]), .Z(n40667) );
  XOR U57569 ( .A(x[204]), .B(y[204]), .Z(n38622) );
  IV U57570 ( .A(n38622), .Z(n40673) );
  IV U57571 ( .A(x[203]), .Z(n38623) );
  XOR U57572 ( .A(n38623), .B(y[203]), .Z(n40671) );
  XOR U57573 ( .A(x[202]), .B(y[202]), .Z(n40678) );
  XOR U57574 ( .A(x[201]), .B(y[201]), .Z(n40675) );
  XOR U57575 ( .A(x[200]), .B(y[200]), .Z(n38624) );
  IV U57576 ( .A(n38624), .Z(n41447) );
  IV U57577 ( .A(x[199]), .Z(n38625) );
  XOR U57578 ( .A(n38625), .B(y[199]), .Z(n41445) );
  XOR U57579 ( .A(x[198]), .B(y[198]), .Z(n41441) );
  XOR U57580 ( .A(x[197]), .B(y[197]), .Z(n41438) );
  XOR U57581 ( .A(x[196]), .B(y[196]), .Z(n38626) );
  IV U57582 ( .A(n38626), .Z(n40684) );
  IV U57583 ( .A(x[195]), .Z(n38627) );
  XOR U57584 ( .A(n38627), .B(y[195]), .Z(n40681) );
  XOR U57585 ( .A(x[194]), .B(y[194]), .Z(n40686) );
  XOR U57586 ( .A(x[193]), .B(y[193]), .Z(n41429) );
  XOR U57587 ( .A(x[192]), .B(y[192]), .Z(n40689) );
  XOR U57588 ( .A(x[191]), .B(y[191]), .Z(n41423) );
  XOR U57589 ( .A(x[190]), .B(y[190]), .Z(n41420) );
  XOR U57590 ( .A(x[189]), .B(y[189]), .Z(n40692) );
  XOR U57591 ( .A(x[188]), .B(y[188]), .Z(n40698) );
  XOR U57592 ( .A(x[187]), .B(y[187]), .Z(n40695) );
  XOR U57593 ( .A(x[186]), .B(y[186]), .Z(n41416) );
  XOR U57594 ( .A(x[185]), .B(y[185]), .Z(n41413) );
  XOR U57595 ( .A(x[184]), .B(y[184]), .Z(n40704) );
  XOR U57596 ( .A(x[183]), .B(y[183]), .Z(n40701) );
  XOR U57597 ( .A(x[182]), .B(y[182]), .Z(n41409) );
  XOR U57598 ( .A(x[181]), .B(y[181]), .Z(n41406) );
  XOR U57599 ( .A(x[180]), .B(y[180]), .Z(n41395) );
  XOR U57600 ( .A(x[179]), .B(y[179]), .Z(n40707) );
  XOR U57601 ( .A(x[178]), .B(y[178]), .Z(n41398) );
  XOR U57602 ( .A(x[177]), .B(y[177]), .Z(n40711) );
  XOR U57603 ( .A(x[176]), .B(y[176]), .Z(n41382) );
  XOR U57604 ( .A(x[175]), .B(y[175]), .Z(n40714) );
  XOR U57605 ( .A(x[174]), .B(y[174]), .Z(n40720) );
  XOR U57606 ( .A(x[173]), .B(y[173]), .Z(n40717) );
  XOR U57607 ( .A(x[172]), .B(y[172]), .Z(n41370) );
  XOR U57608 ( .A(x[171]), .B(y[171]), .Z(n41367) );
  XOR U57609 ( .A(x[170]), .B(y[170]), .Z(n40723) );
  XOR U57610 ( .A(x[169]), .B(y[169]), .Z(n40730) );
  XOR U57611 ( .A(x[168]), .B(y[168]), .Z(n40727) );
  XOR U57612 ( .A(x[167]), .B(y[167]), .Z(n40733) );
  XOR U57613 ( .A(x[166]), .B(y[166]), .Z(n41362) );
  XOR U57614 ( .A(x[165]), .B(y[165]), .Z(n41359) );
  XOR U57615 ( .A(x[164]), .B(y[164]), .Z(n40739) );
  XOR U57616 ( .A(x[163]), .B(y[163]), .Z(n40736) );
  XOR U57617 ( .A(x[162]), .B(y[162]), .Z(n40745) );
  XOR U57618 ( .A(x[161]), .B(y[161]), .Z(n40742) );
  XOR U57619 ( .A(x[160]), .B(y[160]), .Z(n40751) );
  XOR U57620 ( .A(x[159]), .B(y[159]), .Z(n40748) );
  XOR U57621 ( .A(x[158]), .B(y[158]), .Z(n40754) );
  XOR U57622 ( .A(x[157]), .B(y[157]), .Z(n41353) );
  XOR U57623 ( .A(x[156]), .B(y[156]), .Z(n41350) );
  XOR U57624 ( .A(x[155]), .B(y[155]), .Z(n40760) );
  XOR U57625 ( .A(x[154]), .B(y[154]), .Z(n40757) );
  XOR U57626 ( .A(x[153]), .B(y[153]), .Z(n40763) );
  XOR U57627 ( .A(x[152]), .B(y[152]), .Z(n40769) );
  XOR U57628 ( .A(x[151]), .B(y[151]), .Z(n40766) );
  XOR U57629 ( .A(x[150]), .B(y[150]), .Z(n40776) );
  XOR U57630 ( .A(x[149]), .B(y[149]), .Z(n40773) );
  XOR U57631 ( .A(x[148]), .B(y[148]), .Z(n41347) );
  XOR U57632 ( .A(x[147]), .B(y[147]), .Z(n41344) );
  XOR U57633 ( .A(x[146]), .B(y[146]), .Z(n40782) );
  XOR U57634 ( .A(x[145]), .B(y[145]), .Z(n40779) );
  XOR U57635 ( .A(x[144]), .B(y[144]), .Z(n40788) );
  XOR U57636 ( .A(x[143]), .B(y[143]), .Z(n40785) );
  XOR U57637 ( .A(x[142]), .B(y[142]), .Z(n40794) );
  XOR U57638 ( .A(x[141]), .B(y[141]), .Z(n40791) );
  XOR U57639 ( .A(x[140]), .B(y[140]), .Z(n40800) );
  XOR U57640 ( .A(x[139]), .B(y[139]), .Z(n40797) );
  XOR U57641 ( .A(x[138]), .B(y[138]), .Z(n40806) );
  XOR U57642 ( .A(x[137]), .B(y[137]), .Z(n40803) );
  XOR U57643 ( .A(x[136]), .B(y[136]), .Z(n40809) );
  XOR U57644 ( .A(x[135]), .B(y[135]), .Z(n41335) );
  XOR U57645 ( .A(x[134]), .B(y[134]), .Z(n41332) );
  XOR U57646 ( .A(x[133]), .B(y[133]), .Z(n41329) );
  XOR U57647 ( .A(x[132]), .B(y[132]), .Z(n41326) );
  XOR U57648 ( .A(x[131]), .B(y[131]), .Z(n40815) );
  XOR U57649 ( .A(x[130]), .B(y[130]), .Z(n40812) );
  XOR U57650 ( .A(x[129]), .B(y[129]), .Z(n40821) );
  XOR U57651 ( .A(x[128]), .B(y[128]), .Z(n40818) );
  XOR U57652 ( .A(x[127]), .B(y[127]), .Z(n41313) );
  XOR U57653 ( .A(x[126]), .B(y[126]), .Z(n41310) );
  XOR U57654 ( .A(x[125]), .B(y[125]), .Z(n40827) );
  XOR U57655 ( .A(x[124]), .B(y[124]), .Z(n40824) );
  XOR U57656 ( .A(x[123]), .B(y[123]), .Z(n41306) );
  XOR U57657 ( .A(x[122]), .B(y[122]), .Z(n41303) );
  XOR U57658 ( .A(x[121]), .B(y[121]), .Z(n41299) );
  XOR U57659 ( .A(x[120]), .B(y[120]), .Z(n41296) );
  XOR U57660 ( .A(x[119]), .B(y[119]), .Z(n40830) );
  XOR U57661 ( .A(x[118]), .B(y[118]), .Z(n41292) );
  XOR U57662 ( .A(x[117]), .B(y[117]), .Z(n41289) );
  XOR U57663 ( .A(x[116]), .B(y[116]), .Z(n40833) );
  XOR U57664 ( .A(x[115]), .B(y[115]), .Z(n41283) );
  XOR U57665 ( .A(x[114]), .B(y[114]), .Z(n40836) );
  XOR U57666 ( .A(x[113]), .B(y[113]), .Z(n40842) );
  XOR U57667 ( .A(x[112]), .B(y[112]), .Z(n40839) );
  XOR U57668 ( .A(x[111]), .B(y[111]), .Z(n40848) );
  XOR U57669 ( .A(x[110]), .B(y[110]), .Z(n40845) );
  XOR U57670 ( .A(x[109]), .B(y[109]), .Z(n40851) );
  XOR U57671 ( .A(x[108]), .B(y[108]), .Z(n41275) );
  XOR U57672 ( .A(x[107]), .B(y[107]), .Z(n41272) );
  XOR U57673 ( .A(x[106]), .B(y[106]), .Z(n40857) );
  XOR U57674 ( .A(x[105]), .B(y[105]), .Z(n40854) );
  XOR U57675 ( .A(x[104]), .B(y[104]), .Z(n40863) );
  XOR U57676 ( .A(x[103]), .B(y[103]), .Z(n40860) );
  XOR U57677 ( .A(x[102]), .B(y[102]), .Z(n40869) );
  XOR U57678 ( .A(x[101]), .B(y[101]), .Z(n40866) );
  XOR U57679 ( .A(x[100]), .B(y[100]), .Z(n40875) );
  XOR U57680 ( .A(x[99]), .B(y[99]), .Z(n40872) );
  XOR U57681 ( .A(x[98]), .B(y[98]), .Z(n41264) );
  XOR U57682 ( .A(x[97]), .B(y[97]), .Z(n41261) );
  XOR U57683 ( .A(x[96]), .B(y[96]), .Z(n40881) );
  XOR U57684 ( .A(x[95]), .B(y[95]), .Z(n40878) );
  XOR U57685 ( .A(x[94]), .B(y[94]), .Z(n40887) );
  XOR U57686 ( .A(x[93]), .B(y[93]), .Z(n40884) );
  XOR U57687 ( .A(x[92]), .B(y[92]), .Z(n41256) );
  XOR U57688 ( .A(x[91]), .B(y[91]), .Z(n41253) );
  XOR U57689 ( .A(x[90]), .B(y[90]), .Z(n41249) );
  XOR U57690 ( .A(x[89]), .B(y[89]), .Z(n41246) );
  XOR U57691 ( .A(x[88]), .B(y[88]), .Z(n41242) );
  XOR U57692 ( .A(x[87]), .B(y[87]), .Z(n41239) );
  XOR U57693 ( .A(x[86]), .B(y[86]), .Z(n40893) );
  XOR U57694 ( .A(x[85]), .B(y[85]), .Z(n40890) );
  XOR U57695 ( .A(x[84]), .B(y[84]), .Z(n40899) );
  XOR U57696 ( .A(x[83]), .B(y[83]), .Z(n40896) );
  XOR U57697 ( .A(x[82]), .B(y[82]), .Z(n41235) );
  XOR U57698 ( .A(x[81]), .B(y[81]), .Z(n41232) );
  XOR U57699 ( .A(x[80]), .B(y[80]), .Z(n40906) );
  XOR U57700 ( .A(x[79]), .B(y[79]), .Z(n40903) );
  XOR U57701 ( .A(x[78]), .B(y[78]), .Z(n40912) );
  XOR U57702 ( .A(x[77]), .B(y[77]), .Z(n40909) );
  XOR U57703 ( .A(x[76]), .B(y[76]), .Z(n40915) );
  XOR U57704 ( .A(x[75]), .B(y[75]), .Z(n41225) );
  XOR U57705 ( .A(x[74]), .B(y[74]), .Z(n41222) );
  XOR U57706 ( .A(x[73]), .B(y[73]), .Z(n41219) );
  XOR U57707 ( .A(x[72]), .B(y[72]), .Z(n41216) );
  XOR U57708 ( .A(x[71]), .B(y[71]), .Z(n41212) );
  XOR U57709 ( .A(x[70]), .B(y[70]), .Z(n41209) );
  XOR U57710 ( .A(x[69]), .B(y[69]), .Z(n41205) );
  XOR U57711 ( .A(x[68]), .B(y[68]), .Z(n41202) );
  XOR U57712 ( .A(x[67]), .B(y[67]), .Z(n41198) );
  XOR U57713 ( .A(x[66]), .B(y[66]), .Z(n41195) );
  XOR U57714 ( .A(x[65]), .B(y[65]), .Z(n40918) );
  XOR U57715 ( .A(x[64]), .B(y[64]), .Z(n41191) );
  XOR U57716 ( .A(x[63]), .B(y[63]), .Z(n41188) );
  XOR U57717 ( .A(x[62]), .B(y[62]), .Z(n41184) );
  XOR U57718 ( .A(x[61]), .B(y[61]), .Z(n41181) );
  XOR U57719 ( .A(x[60]), .B(y[60]), .Z(n40921) );
  XOR U57720 ( .A(x[59]), .B(y[59]), .Z(n41178) );
  XOR U57721 ( .A(x[58]), .B(y[58]), .Z(n41175) );
  XOR U57722 ( .A(x[57]), .B(y[57]), .Z(n41171) );
  XOR U57723 ( .A(x[56]), .B(y[56]), .Z(n41168) );
  XOR U57724 ( .A(x[55]), .B(y[55]), .Z(n40927) );
  XOR U57725 ( .A(x[54]), .B(y[54]), .Z(n40924) );
  XOR U57726 ( .A(x[53]), .B(y[53]), .Z(n41157) );
  XOR U57727 ( .A(x[52]), .B(y[52]), .Z(n40930) );
  XOR U57728 ( .A(x[51]), .B(y[51]), .Z(n41160) );
  XOR U57729 ( .A(x[50]), .B(y[50]), .Z(n40934) );
  XOR U57730 ( .A(x[49]), .B(y[49]), .Z(n40940) );
  XOR U57731 ( .A(x[48]), .B(y[48]), .Z(n40937) );
  XOR U57732 ( .A(x[47]), .B(y[47]), .Z(n40947) );
  XOR U57733 ( .A(x[46]), .B(y[46]), .Z(n40944) );
  XOR U57734 ( .A(x[45]), .B(y[45]), .Z(n40953) );
  XOR U57735 ( .A(x[44]), .B(y[44]), .Z(n40950) );
  XOR U57736 ( .A(x[43]), .B(y[43]), .Z(n41152) );
  XOR U57737 ( .A(x[42]), .B(y[42]), .Z(n41149) );
  XOR U57738 ( .A(x[41]), .B(y[41]), .Z(n41145) );
  XOR U57739 ( .A(x[40]), .B(y[40]), .Z(n41142) );
  XOR U57740 ( .A(x[39]), .B(y[39]), .Z(n40956) );
  XOR U57741 ( .A(x[38]), .B(y[38]), .Z(n40963) );
  XOR U57742 ( .A(x[37]), .B(y[37]), .Z(n40960) );
  XOR U57743 ( .A(x[36]), .B(y[36]), .Z(n40969) );
  XOR U57744 ( .A(x[35]), .B(y[35]), .Z(n40966) );
  XOR U57745 ( .A(x[34]), .B(y[34]), .Z(n40973) );
  XOR U57746 ( .A(x[33]), .B(y[33]), .Z(n41130) );
  XOR U57747 ( .A(x[32]), .B(y[32]), .Z(n40976) );
  XOR U57748 ( .A(x[31]), .B(y[31]), .Z(n41117) );
  XOR U57749 ( .A(x[30]), .B(y[30]), .Z(n40979) );
  XOR U57750 ( .A(x[29]), .B(y[29]), .Z(n41109) );
  XOR U57751 ( .A(x[28]), .B(y[28]), .Z(n40982) );
  XOR U57752 ( .A(x[27]), .B(y[27]), .Z(n40988) );
  XOR U57753 ( .A(x[26]), .B(y[26]), .Z(n40985) );
  XOR U57754 ( .A(x[25]), .B(y[25]), .Z(n40995) );
  XOR U57755 ( .A(x[24]), .B(y[24]), .Z(n40992) );
  XOR U57756 ( .A(x[23]), .B(y[23]), .Z(n40998) );
  XOR U57757 ( .A(x[22]), .B(y[22]), .Z(n41094) );
  XOR U57758 ( .A(x[21]), .B(y[21]), .Z(n41001) );
  XOR U57759 ( .A(x[20]), .B(y[20]), .Z(n41082) );
  XOR U57760 ( .A(x[19]), .B(y[19]), .Z(n41074) );
  XOR U57761 ( .A(x[18]), .B(y[18]), .Z(n41071) );
  XOR U57762 ( .A(x[17]), .B(y[17]), .Z(n41007) );
  XOR U57763 ( .A(x[16]), .B(y[16]), .Z(n41004) );
  XOR U57764 ( .A(x[15]), .B(y[15]), .Z(n41010) );
  XOR U57765 ( .A(x[14]), .B(y[14]), .Z(n41064) );
  XOR U57766 ( .A(x[13]), .B(y[13]), .Z(n41013) );
  XOR U57767 ( .A(x[12]), .B(y[12]), .Z(n41019) );
  XOR U57768 ( .A(x[11]), .B(y[11]), .Z(n41016) );
  XOR U57769 ( .A(x[10]), .B(y[10]), .Z(n41025) );
  XOR U57770 ( .A(x[9]), .B(y[9]), .Z(n41022) );
  XOR U57771 ( .A(x[8]), .B(y[8]), .Z(n41031) );
  XOR U57772 ( .A(x[7]), .B(y[7]), .Z(n41028) );
  IV U57773 ( .A(x[6]), .Z(n38628) );
  XOR U57774 ( .A(n38628), .B(y[6]), .Z(n41057) );
  XOR U57775 ( .A(x[5]), .B(y[5]), .Z(n41053) );
  XOR U57776 ( .A(x[4]), .B(y[4]), .Z(n41035) );
  XOR U57777 ( .A(y[3]), .B(x[3]), .Z(n41038) );
  XOR U57778 ( .A(x[2]), .B(y[2]), .Z(n41047) );
  XOR U57779 ( .A(x[1]), .B(y[1]), .Z(n38629) );
  IV U57780 ( .A(n38629), .Z(n41044) );
  XOR U57781 ( .A(y[0]), .B(x[0]), .Z(n41042) );
  XOR U57782 ( .A(n41044), .B(n41042), .Z(n41048) );
  XOR U57783 ( .A(n41047), .B(n41048), .Z(n41039) );
  XOR U57784 ( .A(n41038), .B(n41039), .Z(n41036) );
  XOR U57785 ( .A(n41035), .B(n41036), .Z(n41054) );
  XOR U57786 ( .A(n41053), .B(n41054), .Z(n41056) );
  XOR U57787 ( .A(n41057), .B(n41056), .Z(n41029) );
  XOR U57788 ( .A(n41028), .B(n41029), .Z(n38630) );
  IV U57789 ( .A(n38630), .Z(n41030) );
  XOR U57790 ( .A(n41031), .B(n41030), .Z(n41024) );
  XOR U57791 ( .A(n41022), .B(n41024), .Z(n41027) );
  XOR U57792 ( .A(n41025), .B(n41027), .Z(n41018) );
  XOR U57793 ( .A(n41016), .B(n41018), .Z(n41021) );
  XOR U57794 ( .A(n41019), .B(n41021), .Z(n41015) );
  XOR U57795 ( .A(n41013), .B(n41015), .Z(n41066) );
  XOR U57796 ( .A(n41064), .B(n41066), .Z(n41012) );
  XOR U57797 ( .A(n41010), .B(n41012), .Z(n41006) );
  XOR U57798 ( .A(n41004), .B(n41006), .Z(n41009) );
  XOR U57799 ( .A(n41007), .B(n41009), .Z(n41072) );
  XOR U57800 ( .A(n41071), .B(n41072), .Z(n41076) );
  XOR U57801 ( .A(n41074), .B(n41076), .Z(n41084) );
  XOR U57802 ( .A(n41082), .B(n41084), .Z(n41003) );
  XOR U57803 ( .A(n41001), .B(n41003), .Z(n41096) );
  XOR U57804 ( .A(n41094), .B(n41096), .Z(n41000) );
  XOR U57805 ( .A(n40998), .B(n41000), .Z(n40994) );
  XOR U57806 ( .A(n40992), .B(n40994), .Z(n40996) );
  XOR U57807 ( .A(n40995), .B(n40996), .Z(n40986) );
  XOR U57808 ( .A(n40985), .B(n40986), .Z(n40989) );
  XOR U57809 ( .A(n40988), .B(n40989), .Z(n40984) );
  XOR U57810 ( .A(n40982), .B(n40984), .Z(n41111) );
  XOR U57811 ( .A(n41109), .B(n41111), .Z(n40981) );
  XOR U57812 ( .A(n40979), .B(n40981), .Z(n41118) );
  XOR U57813 ( .A(n41117), .B(n41118), .Z(n40977) );
  XOR U57814 ( .A(n40976), .B(n40977), .Z(n41132) );
  XOR U57815 ( .A(n41130), .B(n41132), .Z(n40975) );
  XOR U57816 ( .A(n40973), .B(n40975), .Z(n40967) );
  XOR U57817 ( .A(n40966), .B(n40967), .Z(n40971) );
  XOR U57818 ( .A(n40969), .B(n40971), .Z(n40962) );
  XOR U57819 ( .A(n40960), .B(n40962), .Z(n40964) );
  XOR U57820 ( .A(n40963), .B(n40964), .Z(n40957) );
  XOR U57821 ( .A(n40956), .B(n40957), .Z(n41143) );
  XOR U57822 ( .A(n41142), .B(n41143), .Z(n41147) );
  XOR U57823 ( .A(n41145), .B(n41147), .Z(n41151) );
  XOR U57824 ( .A(n41149), .B(n41151), .Z(n41153) );
  XOR U57825 ( .A(n41152), .B(n41153), .Z(n40952) );
  XOR U57826 ( .A(n40950), .B(n40952), .Z(n40955) );
  XOR U57827 ( .A(n40953), .B(n40955), .Z(n40946) );
  XOR U57828 ( .A(n40944), .B(n40946), .Z(n40948) );
  XOR U57829 ( .A(n40947), .B(n40948), .Z(n40939) );
  XOR U57830 ( .A(n40937), .B(n40939), .Z(n40941) );
  XOR U57831 ( .A(n40940), .B(n40941), .Z(n40935) );
  XOR U57832 ( .A(n40934), .B(n40935), .Z(n41162) );
  XOR U57833 ( .A(n41160), .B(n41162), .Z(n40932) );
  XOR U57834 ( .A(n40930), .B(n40932), .Z(n41159) );
  XOR U57835 ( .A(n41157), .B(n41159), .Z(n40926) );
  XOR U57836 ( .A(n40924), .B(n40926), .Z(n40928) );
  XOR U57837 ( .A(n40927), .B(n40928), .Z(n41169) );
  XOR U57838 ( .A(n41168), .B(n41169), .Z(n41173) );
  XOR U57839 ( .A(n41171), .B(n41173), .Z(n41177) );
  XOR U57840 ( .A(n41175), .B(n41177), .Z(n41179) );
  XOR U57841 ( .A(n41178), .B(n41179), .Z(n40923) );
  XOR U57842 ( .A(n40921), .B(n40923), .Z(n41183) );
  XOR U57843 ( .A(n41181), .B(n41183), .Z(n41186) );
  XOR U57844 ( .A(n41184), .B(n41186), .Z(n41189) );
  XOR U57845 ( .A(n41188), .B(n41189), .Z(n41192) );
  XOR U57846 ( .A(n41191), .B(n41192), .Z(n40920) );
  XOR U57847 ( .A(n40918), .B(n40920), .Z(n41196) );
  XOR U57848 ( .A(n41195), .B(n41196), .Z(n41199) );
  XOR U57849 ( .A(n41198), .B(n41199), .Z(n41204) );
  XOR U57850 ( .A(n41202), .B(n41204), .Z(n41207) );
  XOR U57851 ( .A(n41205), .B(n41207), .Z(n41210) );
  XOR U57852 ( .A(n41209), .B(n41210), .Z(n41213) );
  XOR U57853 ( .A(n41212), .B(n41213), .Z(n41218) );
  XOR U57854 ( .A(n41216), .B(n41218), .Z(n41221) );
  XOR U57855 ( .A(n41219), .B(n41221), .Z(n41224) );
  XOR U57856 ( .A(n41222), .B(n41224), .Z(n41226) );
  XOR U57857 ( .A(n41225), .B(n41226), .Z(n40917) );
  XOR U57858 ( .A(n40915), .B(n40917), .Z(n40911) );
  XOR U57859 ( .A(n40909), .B(n40911), .Z(n40913) );
  XOR U57860 ( .A(n40912), .B(n40913), .Z(n40904) );
  XOR U57861 ( .A(n40903), .B(n40904), .Z(n40908) );
  XOR U57862 ( .A(n40906), .B(n40908), .Z(n41233) );
  XOR U57863 ( .A(n41232), .B(n41233), .Z(n41236) );
  XOR U57864 ( .A(n41235), .B(n41236), .Z(n40898) );
  XOR U57865 ( .A(n40896), .B(n40898), .Z(n40900) );
  XOR U57866 ( .A(n40899), .B(n40900), .Z(n40892) );
  XOR U57867 ( .A(n40890), .B(n40892), .Z(n40894) );
  XOR U57868 ( .A(n40893), .B(n40894), .Z(n41240) );
  XOR U57869 ( .A(n41239), .B(n41240), .Z(n41243) );
  XOR U57870 ( .A(n41242), .B(n41243), .Z(n41247) );
  XOR U57871 ( .A(n41246), .B(n41247), .Z(n41250) );
  XOR U57872 ( .A(n41249), .B(n41250), .Z(n41255) );
  XOR U57873 ( .A(n41253), .B(n41255), .Z(n41258) );
  XOR U57874 ( .A(n41256), .B(n41258), .Z(n40885) );
  XOR U57875 ( .A(n40884), .B(n40885), .Z(n40889) );
  XOR U57876 ( .A(n40887), .B(n40889), .Z(n40879) );
  XOR U57877 ( .A(n40878), .B(n40879), .Z(n40882) );
  XOR U57878 ( .A(n40881), .B(n40882), .Z(n41263) );
  XOR U57879 ( .A(n41261), .B(n41263), .Z(n41266) );
  XOR U57880 ( .A(n41264), .B(n41266), .Z(n40873) );
  XOR U57881 ( .A(n40872), .B(n40873), .Z(n40877) );
  XOR U57882 ( .A(n40875), .B(n40877), .Z(n40868) );
  XOR U57883 ( .A(n40866), .B(n40868), .Z(n40871) );
  XOR U57884 ( .A(n40869), .B(n40871), .Z(n40861) );
  XOR U57885 ( .A(n40860), .B(n40861), .Z(n40864) );
  XOR U57886 ( .A(n40863), .B(n40864), .Z(n40856) );
  XOR U57887 ( .A(n40854), .B(n40856), .Z(n40858) );
  XOR U57888 ( .A(n40857), .B(n40858), .Z(n41273) );
  XOR U57889 ( .A(n41272), .B(n41273), .Z(n41277) );
  XOR U57890 ( .A(n41275), .B(n41277), .Z(n40852) );
  XOR U57891 ( .A(n40851), .B(n40852), .Z(n40847) );
  XOR U57892 ( .A(n40845), .B(n40847), .Z(n40849) );
  XOR U57893 ( .A(n40848), .B(n40849), .Z(n40841) );
  XOR U57894 ( .A(n40839), .B(n40841), .Z(n40843) );
  XOR U57895 ( .A(n40842), .B(n40843), .Z(n40837) );
  XOR U57896 ( .A(n40836), .B(n40837), .Z(n41285) );
  XOR U57897 ( .A(n41283), .B(n41285), .Z(n40835) );
  XOR U57898 ( .A(n40833), .B(n40835), .Z(n41291) );
  XOR U57899 ( .A(n41289), .B(n41291), .Z(n41294) );
  XOR U57900 ( .A(n41292), .B(n41294), .Z(n40832) );
  XOR U57901 ( .A(n40830), .B(n40832), .Z(n41298) );
  XOR U57902 ( .A(n41296), .B(n41298), .Z(n41300) );
  XOR U57903 ( .A(n41299), .B(n41300), .Z(n41305) );
  XOR U57904 ( .A(n41303), .B(n41305), .Z(n41308) );
  XOR U57905 ( .A(n41306), .B(n41308), .Z(n40826) );
  XOR U57906 ( .A(n40824), .B(n40826), .Z(n40828) );
  XOR U57907 ( .A(n40827), .B(n40828), .Z(n41312) );
  XOR U57908 ( .A(n41310), .B(n41312), .Z(n41314) );
  XOR U57909 ( .A(n41313), .B(n41314), .Z(n40820) );
  XOR U57910 ( .A(n40818), .B(n40820), .Z(n40823) );
  XOR U57911 ( .A(n40821), .B(n40823), .Z(n40814) );
  XOR U57912 ( .A(n40812), .B(n40814), .Z(n40816) );
  XOR U57913 ( .A(n40815), .B(n40816), .Z(n41328) );
  XOR U57914 ( .A(n41326), .B(n41328), .Z(n41331) );
  XOR U57915 ( .A(n41329), .B(n41331), .Z(n41334) );
  XOR U57916 ( .A(n41332), .B(n41334), .Z(n41336) );
  XOR U57917 ( .A(n41335), .B(n41336), .Z(n40810) );
  XOR U57918 ( .A(n40809), .B(n40810), .Z(n40805) );
  XOR U57919 ( .A(n40803), .B(n40805), .Z(n40807) );
  XOR U57920 ( .A(n40806), .B(n40807), .Z(n40798) );
  XOR U57921 ( .A(n40797), .B(n40798), .Z(n40801) );
  XOR U57922 ( .A(n40800), .B(n40801), .Z(n40793) );
  XOR U57923 ( .A(n40791), .B(n40793), .Z(n40796) );
  XOR U57924 ( .A(n40794), .B(n40796), .Z(n40786) );
  XOR U57925 ( .A(n40785), .B(n40786), .Z(n40790) );
  XOR U57926 ( .A(n40788), .B(n40790), .Z(n40780) );
  XOR U57927 ( .A(n40779), .B(n40780), .Z(n40783) );
  XOR U57928 ( .A(n40782), .B(n40783), .Z(n41345) );
  XOR U57929 ( .A(n41344), .B(n41345), .Z(n41349) );
  XOR U57930 ( .A(n41347), .B(n41349), .Z(n40775) );
  XOR U57931 ( .A(n40773), .B(n40775), .Z(n40778) );
  XOR U57932 ( .A(n40776), .B(n40778), .Z(n40768) );
  XOR U57933 ( .A(n40766), .B(n40768), .Z(n40771) );
  XOR U57934 ( .A(n40769), .B(n40771), .Z(n40764) );
  XOR U57935 ( .A(n40763), .B(n40764), .Z(n40758) );
  XOR U57936 ( .A(n40757), .B(n40758), .Z(n40762) );
  XOR U57937 ( .A(n40760), .B(n40762), .Z(n41351) );
  XOR U57938 ( .A(n41350), .B(n41351), .Z(n41354) );
  XOR U57939 ( .A(n41353), .B(n41354), .Z(n40755) );
  XOR U57940 ( .A(n40754), .B(n40755), .Z(n40750) );
  XOR U57941 ( .A(n40748), .B(n40750), .Z(n40753) );
  XOR U57942 ( .A(n40751), .B(n40753), .Z(n40743) );
  XOR U57943 ( .A(n40742), .B(n40743), .Z(n40746) );
  XOR U57944 ( .A(n40745), .B(n40746), .Z(n40738) );
  XOR U57945 ( .A(n40736), .B(n40738), .Z(n40741) );
  XOR U57946 ( .A(n40739), .B(n40741), .Z(n41361) );
  XOR U57947 ( .A(n41359), .B(n41361), .Z(n41363) );
  XOR U57948 ( .A(n41362), .B(n41363), .Z(n40734) );
  XOR U57949 ( .A(n40733), .B(n40734), .Z(n40728) );
  XOR U57950 ( .A(n40727), .B(n40728), .Z(n40732) );
  XOR U57951 ( .A(n40730), .B(n40732), .Z(n40725) );
  XOR U57952 ( .A(n40723), .B(n40725), .Z(n41368) );
  XOR U57953 ( .A(n41367), .B(n41368), .Z(n41372) );
  XOR U57954 ( .A(n41370), .B(n41372), .Z(n40719) );
  XOR U57955 ( .A(n40717), .B(n40719), .Z(n40722) );
  XOR U57956 ( .A(n40720), .B(n40722), .Z(n40716) );
  XOR U57957 ( .A(n40714), .B(n40716), .Z(n41384) );
  XOR U57958 ( .A(n41382), .B(n41384), .Z(n40712) );
  XOR U57959 ( .A(n40711), .B(n40712), .Z(n41399) );
  XOR U57960 ( .A(n41398), .B(n41399), .Z(n40709) );
  XOR U57961 ( .A(n40707), .B(n40709), .Z(n41397) );
  XOR U57962 ( .A(n41395), .B(n41397), .Z(n41407) );
  XOR U57963 ( .A(n41406), .B(n41407), .Z(n41410) );
  XOR U57964 ( .A(n41409), .B(n41410), .Z(n40703) );
  XOR U57965 ( .A(n40701), .B(n40703), .Z(n40706) );
  XOR U57966 ( .A(n40704), .B(n40706), .Z(n41414) );
  XOR U57967 ( .A(n41413), .B(n41414), .Z(n41418) );
  XOR U57968 ( .A(n41416), .B(n41418), .Z(n40697) );
  XOR U57969 ( .A(n40695), .B(n40697), .Z(n40700) );
  XOR U57970 ( .A(n40698), .B(n40700), .Z(n40693) );
  XOR U57971 ( .A(n40692), .B(n40693), .Z(n41422) );
  XOR U57972 ( .A(n41420), .B(n41422), .Z(n41424) );
  XOR U57973 ( .A(n41423), .B(n41424), .Z(n40690) );
  XOR U57974 ( .A(n40689), .B(n40690), .Z(n41431) );
  XOR U57975 ( .A(n41429), .B(n41431), .Z(n40688) );
  XOR U57976 ( .A(n40686), .B(n40688), .Z(n40682) );
  XOR U57977 ( .A(n40681), .B(n40682), .Z(n40683) );
  XOR U57978 ( .A(n40684), .B(n40683), .Z(n41439) );
  XOR U57979 ( .A(n41438), .B(n41439), .Z(n41443) );
  XOR U57980 ( .A(n41441), .B(n41443), .Z(n41444) );
  XOR U57981 ( .A(n41445), .B(n41444), .Z(n41446) );
  XOR U57982 ( .A(n41447), .B(n41446), .Z(n40676) );
  XOR U57983 ( .A(n40675), .B(n40676), .Z(n40680) );
  XOR U57984 ( .A(n40678), .B(n40680), .Z(n40670) );
  XOR U57985 ( .A(n40671), .B(n40670), .Z(n40672) );
  XOR U57986 ( .A(n40673), .B(n40672), .Z(n40669) );
  XOR U57987 ( .A(n40667), .B(n40669), .Z(n41454) );
  XOR U57988 ( .A(n41453), .B(n41454), .Z(n40665) );
  XOR U57989 ( .A(n40666), .B(n40665), .Z(n41459) );
  XOR U57990 ( .A(n41461), .B(n41459), .Z(n41463) );
  XOR U57991 ( .A(n41462), .B(n41463), .Z(n40663) );
  XOR U57992 ( .A(n40662), .B(n40663), .Z(n41469) );
  XOR U57993 ( .A(n41468), .B(n41469), .Z(n40659) );
  XOR U57994 ( .A(n40660), .B(n40659), .Z(n41477) );
  XOR U57995 ( .A(n41475), .B(n41477), .Z(n40657) );
  XOR U57996 ( .A(n40656), .B(n40657), .Z(n41487) );
  XOR U57997 ( .A(n41486), .B(n41487), .Z(n41488) );
  XOR U57998 ( .A(n41489), .B(n41488), .Z(n40651) );
  XOR U57999 ( .A(n40650), .B(n40651), .Z(n40654) );
  XOR U58000 ( .A(n40653), .B(n40654), .Z(n41505) );
  XOR U58001 ( .A(n41503), .B(n41505), .Z(n41507) );
  XOR U58002 ( .A(n41506), .B(n41507), .Z(n40645) );
  XOR U58003 ( .A(n40644), .B(n40645), .Z(n40648) );
  XOR U58004 ( .A(n40647), .B(n40648), .Z(n41510) );
  XOR U58005 ( .A(n41509), .B(n41510), .Z(n41513) );
  XOR U58006 ( .A(n41512), .B(n41513), .Z(n40640) );
  XOR U58007 ( .A(n40638), .B(n40640), .Z(n40643) );
  XOR U58008 ( .A(n40641), .B(n40643), .Z(n40632) );
  XOR U58009 ( .A(n40633), .B(n40632), .Z(n40634) );
  XOR U58010 ( .A(n40635), .B(n40634), .Z(n40630) );
  XOR U58011 ( .A(n40628), .B(n40630), .Z(n40624) );
  XOR U58012 ( .A(n40622), .B(n40624), .Z(n40626) );
  XOR U58013 ( .A(n40625), .B(n40626), .Z(n41518) );
  XOR U58014 ( .A(n41517), .B(n41518), .Z(n41522) );
  XOR U58015 ( .A(n41520), .B(n41522), .Z(n40618) );
  XOR U58016 ( .A(n40616), .B(n40618), .Z(n40620) );
  XOR U58017 ( .A(n40619), .B(n40620), .Z(n40614) );
  XOR U58018 ( .A(n40612), .B(n40614), .Z(n41525) );
  XOR U58019 ( .A(n41523), .B(n41525), .Z(n41528) );
  XOR U58020 ( .A(n41526), .B(n41528), .Z(n40607) );
  XOR U58021 ( .A(n40608), .B(n40607), .Z(n40609) );
  XOR U58022 ( .A(n40610), .B(n40609), .Z(n41532) );
  IV U58023 ( .A(n41532), .Z(n41530) );
  XOR U58024 ( .A(n41533), .B(n41530), .Z(n51317) );
  XOR U58025 ( .A(n51315), .B(n51317), .Z(n41538) );
  XOR U58026 ( .A(n41536), .B(n41538), .Z(n41539) );
  XOR U58027 ( .A(n41540), .B(n41539), .Z(n40601) );
  IV U58028 ( .A(n40601), .Z(n40604) );
  XOR U58029 ( .A(n40602), .B(n40604), .Z(n56529) );
  XOR U58030 ( .A(n56527), .B(n56529), .Z(n40596) );
  XOR U58031 ( .A(n40595), .B(n40596), .Z(n40600) );
  XOR U58032 ( .A(n40598), .B(n40600), .Z(n41544) );
  XOR U58033 ( .A(n41542), .B(n41544), .Z(n41546) );
  XOR U58034 ( .A(n41545), .B(n41546), .Z(n40593) );
  XOR U58035 ( .A(n40592), .B(n40593), .Z(n40587) );
  XOR U58036 ( .A(n40586), .B(n40587), .Z(n40591) );
  XOR U58037 ( .A(n40589), .B(n40591), .Z(n40584) );
  XOR U58038 ( .A(n40582), .B(n40584), .Z(n41551) );
  XOR U58039 ( .A(n41550), .B(n41551), .Z(n41555) );
  XOR U58040 ( .A(n41553), .B(n41555), .Z(n40576) );
  XOR U58041 ( .A(n40575), .B(n40576), .Z(n40579) );
  XOR U58042 ( .A(n40578), .B(n40579), .Z(n41558) );
  XOR U58043 ( .A(n41557), .B(n41558), .Z(n41561) );
  XOR U58044 ( .A(n41560), .B(n41561), .Z(n40571) );
  XOR U58045 ( .A(n40569), .B(n40571), .Z(n40574) );
  XOR U58046 ( .A(n40572), .B(n40574), .Z(n41564) );
  XOR U58047 ( .A(n41563), .B(n41564), .Z(n41567) );
  XOR U58048 ( .A(n41566), .B(n41567), .Z(n40567) );
  XOR U58049 ( .A(n40566), .B(n40567), .Z(n41571) );
  XOR U58050 ( .A(n41570), .B(n41571), .Z(n41574) );
  XOR U58051 ( .A(n41573), .B(n41574), .Z(n40565) );
  XOR U58052 ( .A(n40563), .B(n40565), .Z(n41580) );
  XOR U58053 ( .A(n41578), .B(n41580), .Z(n41583) );
  XOR U58054 ( .A(n41581), .B(n41583), .Z(n41586) );
  XOR U58055 ( .A(n41585), .B(n41586), .Z(n41590) );
  XOR U58056 ( .A(n41588), .B(n41590), .Z(n52158) );
  IV U58057 ( .A(n52158), .Z(n40559) );
  XOR U58058 ( .A(x[273]), .B(y[273]), .Z(n52159) );
  IV U58059 ( .A(x[274]), .Z(n38631) );
  XOR U58060 ( .A(n38631), .B(y[274]), .Z(n52161) );
  XOR U58061 ( .A(n52159), .B(n52161), .Z(n38632) );
  XOR U58062 ( .A(n40559), .B(n38632), .Z(n41593) );
  XOR U58063 ( .A(n41591), .B(n41593), .Z(n41595) );
  XOR U58064 ( .A(n41594), .B(n41595), .Z(n41600) );
  XOR U58065 ( .A(n41598), .B(n41600), .Z(n41603) );
  XOR U58066 ( .A(n41601), .B(n41603), .Z(n41606) );
  XOR U58067 ( .A(n41605), .B(n41606), .Z(n41610) );
  XOR U58068 ( .A(n41608), .B(n41610), .Z(n40556) );
  XOR U58069 ( .A(n40555), .B(n40556), .Z(n41617) );
  XOR U58070 ( .A(n41616), .B(n41617), .Z(n41620) );
  XOR U58071 ( .A(n41619), .B(n41620), .Z(n41623) );
  XOR U58072 ( .A(n41622), .B(n41623), .Z(n41626) );
  XOR U58073 ( .A(n41625), .B(n41626), .Z(n40550) );
  XOR U58074 ( .A(n40549), .B(n40550), .Z(n40554) );
  XOR U58075 ( .A(n40552), .B(n40554), .Z(n40545) );
  XOR U58076 ( .A(n40543), .B(n40545), .Z(n40547) );
  XOR U58077 ( .A(n40546), .B(n40547), .Z(n41630) );
  XOR U58078 ( .A(n41629), .B(n41630), .Z(n41633) );
  XOR U58079 ( .A(n41632), .B(n41633), .Z(n40537) );
  XOR U58080 ( .A(n40538), .B(n40537), .Z(n40542) );
  XOR U58081 ( .A(n40540), .B(n40542), .Z(n40533) );
  XOR U58082 ( .A(n40531), .B(n40533), .Z(n40535) );
  XOR U58083 ( .A(n40534), .B(n40535), .Z(n40526) );
  XOR U58084 ( .A(n40525), .B(n40526), .Z(n40530) );
  XOR U58085 ( .A(n40528), .B(n40530), .Z(n40523) );
  XOR U58086 ( .A(n40521), .B(n40523), .Z(n41636) );
  XOR U58087 ( .A(n41635), .B(n41636), .Z(n41640) );
  XOR U58088 ( .A(n41638), .B(n41640), .Z(n40517) );
  XOR U58089 ( .A(n40515), .B(n40517), .Z(n40519) );
  XOR U58090 ( .A(n40518), .B(n40519), .Z(n40513) );
  XOR U58091 ( .A(n40514), .B(n40513), .Z(n41641) );
  XOR U58092 ( .A(n41642), .B(n41641), .Z(n41645) );
  XOR U58093 ( .A(n41644), .B(n41645), .Z(n41657) );
  XOR U58094 ( .A(n41656), .B(n41657), .Z(n41651) );
  XOR U58095 ( .A(n41649), .B(n41651), .Z(n41654) );
  XOR U58096 ( .A(n41653), .B(n41654), .Z(n41666) );
  XOR U58097 ( .A(n41664), .B(n41666), .Z(n41668) );
  XOR U58098 ( .A(n41667), .B(n41668), .Z(n41672) );
  XOR U58099 ( .A(n41671), .B(n41672), .Z(n41675) );
  XOR U58100 ( .A(n41674), .B(n41675), .Z(n41680) );
  XOR U58101 ( .A(n41678), .B(n41680), .Z(n41683) );
  XOR U58102 ( .A(n41681), .B(n41683), .Z(n41686) );
  XOR U58103 ( .A(n41685), .B(n41686), .Z(n41687) );
  XOR U58104 ( .A(n41688), .B(n41687), .Z(n41692) );
  XOR U58105 ( .A(n41690), .B(n41692), .Z(n41695) );
  XOR U58106 ( .A(n41693), .B(n41695), .Z(n40508) );
  XOR U58107 ( .A(n40507), .B(n40508), .Z(n40511) );
  XOR U58108 ( .A(n40510), .B(n40511), .Z(n40503) );
  XOR U58109 ( .A(n40501), .B(n40503), .Z(n40506) );
  XOR U58110 ( .A(n40504), .B(n40506), .Z(n40496) );
  XOR U58111 ( .A(n40495), .B(n40496), .Z(n40500) );
  XOR U58112 ( .A(n40498), .B(n40500), .Z(n41700) );
  XOR U58113 ( .A(n41698), .B(n41700), .Z(n41702) );
  XOR U58114 ( .A(n41701), .B(n41702), .Z(n41715) );
  XOR U58115 ( .A(n41716), .B(n41715), .Z(n41717) );
  XOR U58116 ( .A(n41718), .B(n41717), .Z(n41723) );
  XOR U58117 ( .A(n41721), .B(n41723), .Z(n41726) );
  XOR U58118 ( .A(n41724), .B(n41726), .Z(n41729) );
  XOR U58119 ( .A(n41728), .B(n41729), .Z(n41733) );
  XOR U58120 ( .A(n41731), .B(n41733), .Z(n40490) );
  XOR U58121 ( .A(n40489), .B(n40490), .Z(n40494) );
  XOR U58122 ( .A(n40492), .B(n40494), .Z(n40483) );
  XOR U58123 ( .A(n40482), .B(n40483), .Z(n40486) );
  XOR U58124 ( .A(n40485), .B(n40486), .Z(n57401) );
  XOR U58125 ( .A(n57399), .B(n57401), .Z(n41737) );
  XOR U58126 ( .A(n41738), .B(n41737), .Z(n41743) );
  XOR U58127 ( .A(n41741), .B(n41743), .Z(n41746) );
  XOR U58128 ( .A(n41744), .B(n41746), .Z(n40478) );
  XOR U58129 ( .A(n40476), .B(n40478), .Z(n40481) );
  XOR U58130 ( .A(n40479), .B(n40481), .Z(n41749) );
  XOR U58131 ( .A(n41747), .B(n41749), .Z(n41751) );
  XOR U58132 ( .A(n41750), .B(n41751), .Z(n40471) );
  XOR U58133 ( .A(n40470), .B(n40471), .Z(n40475) );
  XOR U58134 ( .A(n40473), .B(n40475), .Z(n41756) );
  XOR U58135 ( .A(n41754), .B(n41756), .Z(n41759) );
  XOR U58136 ( .A(n41757), .B(n41759), .Z(n40466) );
  XOR U58137 ( .A(n40465), .B(n40466), .Z(n40467) );
  XOR U58138 ( .A(n40468), .B(n40467), .Z(n41762) );
  XOR U58139 ( .A(n41761), .B(n41762), .Z(n41763) );
  XOR U58140 ( .A(n41764), .B(n41763), .Z(n40462) );
  XOR U58141 ( .A(n40461), .B(n40462), .Z(n40457) );
  XOR U58142 ( .A(n40456), .B(n40457), .Z(n40460) );
  XOR U58143 ( .A(n40459), .B(n40460), .Z(n40450) );
  XOR U58144 ( .A(n40451), .B(n40450), .Z(n40455) );
  XOR U58145 ( .A(n40453), .B(n40455), .Z(n40446) );
  XOR U58146 ( .A(n40445), .B(n40446), .Z(n40448) );
  XOR U58147 ( .A(n40449), .B(n40448), .Z(n41769) );
  XOR U58148 ( .A(n41771), .B(n41769), .Z(n41774) );
  XOR U58149 ( .A(n41772), .B(n41774), .Z(n40442) );
  XOR U58150 ( .A(n40440), .B(n40442), .Z(n40443) );
  XOR U58151 ( .A(n40444), .B(n40443), .Z(n41777) );
  XOR U58152 ( .A(n41778), .B(n41777), .Z(n41782) );
  XOR U58153 ( .A(n41780), .B(n41782), .Z(n41786) );
  XOR U58154 ( .A(n41784), .B(n41786), .Z(n41788) );
  XOR U58155 ( .A(n41787), .B(n41788), .Z(n41793) );
  XOR U58156 ( .A(n41791), .B(n41793), .Z(n41795) );
  XOR U58157 ( .A(n41794), .B(n41795), .Z(n40435) );
  XOR U58158 ( .A(n40433), .B(n40435), .Z(n40437) );
  XOR U58159 ( .A(n40436), .B(n40437), .Z(n40429) );
  XOR U58160 ( .A(n40427), .B(n40429), .Z(n40431) );
  XOR U58161 ( .A(n40430), .B(n40431), .Z(n40426) );
  XOR U58162 ( .A(n40424), .B(n40426), .Z(n40418) );
  XOR U58163 ( .A(n40417), .B(n40418), .Z(n40421) );
  XOR U58164 ( .A(n40420), .B(n40421), .Z(n40412) );
  XOR U58165 ( .A(n40414), .B(n40412), .Z(n46827) );
  XOR U58166 ( .A(n46826), .B(n46827), .Z(n40407) );
  XOR U58167 ( .A(n40405), .B(n40407), .Z(n40410) );
  XOR U58168 ( .A(n40408), .B(n40410), .Z(n40400) );
  XOR U58169 ( .A(n40399), .B(n40400), .Z(n40404) );
  XOR U58170 ( .A(n40402), .B(n40404), .Z(n41802) );
  XOR U58171 ( .A(n41801), .B(n41802), .Z(n41805) );
  XOR U58172 ( .A(n41804), .B(n41805), .Z(n40395) );
  XOR U58173 ( .A(n40393), .B(n40395), .Z(n40397) );
  XOR U58174 ( .A(n40396), .B(n40397), .Z(n40392) );
  XOR U58175 ( .A(n40390), .B(n40392), .Z(n41811) );
  XOR U58176 ( .A(n41809), .B(n41811), .Z(n41814) );
  XOR U58177 ( .A(n41812), .B(n41814), .Z(n40389) );
  XOR U58178 ( .A(n40387), .B(n40389), .Z(n40382) );
  XOR U58179 ( .A(n40381), .B(n40382), .Z(n40385) );
  XOR U58180 ( .A(n40384), .B(n40385), .Z(n40377) );
  XOR U58181 ( .A(n40375), .B(n40377), .Z(n40380) );
  XOR U58182 ( .A(n40378), .B(n40380), .Z(n41819) );
  XOR U58183 ( .A(n41818), .B(n41819), .Z(n41823) );
  XOR U58184 ( .A(n41821), .B(n41823), .Z(n40371) );
  XOR U58185 ( .A(n40369), .B(n40371), .Z(n40374) );
  XOR U58186 ( .A(n40372), .B(n40374), .Z(n40364) );
  XOR U58187 ( .A(n40363), .B(n40364), .Z(n40367) );
  XOR U58188 ( .A(n40366), .B(n40367), .Z(n40359) );
  XOR U58189 ( .A(n40357), .B(n40359), .Z(n40362) );
  XOR U58190 ( .A(n40360), .B(n40362), .Z(n41833) );
  XOR U58191 ( .A(n41832), .B(n41833), .Z(n40354) );
  XOR U58192 ( .A(n40353), .B(n40354), .Z(n41831) );
  XOR U58193 ( .A(n41829), .B(n41831), .Z(n40351) );
  XOR U58194 ( .A(n40349), .B(n40351), .Z(n41845) );
  XOR U58195 ( .A(n41844), .B(n41845), .Z(n41848) );
  XOR U58196 ( .A(n41847), .B(n41848), .Z(n40345) );
  XOR U58197 ( .A(n40343), .B(n40345), .Z(n40348) );
  XOR U58198 ( .A(n40346), .B(n40348), .Z(n40338) );
  XOR U58199 ( .A(n40337), .B(n40338), .Z(n40342) );
  XOR U58200 ( .A(n40340), .B(n40342), .Z(n40333) );
  XOR U58201 ( .A(n40331), .B(n40333), .Z(n40336) );
  XOR U58202 ( .A(n40334), .B(n40336), .Z(n40329) );
  XOR U58203 ( .A(n40328), .B(n40329), .Z(n40323) );
  XOR U58204 ( .A(n40322), .B(n40323), .Z(n40327) );
  XOR U58205 ( .A(n40325), .B(n40327), .Z(n40319) );
  XOR U58206 ( .A(n40318), .B(n40319), .Z(n41853) );
  XOR U58207 ( .A(n41852), .B(n41853), .Z(n41857) );
  XOR U58208 ( .A(n41855), .B(n41857), .Z(n41861) );
  XOR U58209 ( .A(n41859), .B(n41861), .Z(n41864) );
  XOR U58210 ( .A(n41862), .B(n41864), .Z(n41866) );
  XOR U58211 ( .A(n41865), .B(n41866), .Z(n41869) );
  XOR U58212 ( .A(n41868), .B(n41869), .Z(n40313) );
  XOR U58213 ( .A(n40312), .B(n40313), .Z(n40316) );
  XOR U58214 ( .A(n40315), .B(n40316), .Z(n41874) );
  XOR U58215 ( .A(n41873), .B(n41874), .Z(n41878) );
  XOR U58216 ( .A(n41876), .B(n41878), .Z(n41882) );
  XOR U58217 ( .A(n41880), .B(n41882), .Z(n41884) );
  XOR U58218 ( .A(n41883), .B(n41884), .Z(n41888) );
  XOR U58219 ( .A(n41887), .B(n41888), .Z(n41891) );
  XOR U58220 ( .A(n41890), .B(n41891), .Z(n40308) );
  XOR U58221 ( .A(n40306), .B(n40308), .Z(n40310) );
  XOR U58222 ( .A(n40309), .B(n40310), .Z(n40301) );
  XOR U58223 ( .A(n40300), .B(n40301), .Z(n40305) );
  XOR U58224 ( .A(n40303), .B(n40305), .Z(n57589) );
  XOR U58225 ( .A(x[437]), .B(y[437]), .Z(n57588) );
  IV U58226 ( .A(n57588), .Z(n40296) );
  IV U58227 ( .A(x[438]), .Z(n38633) );
  XOR U58228 ( .A(n38633), .B(y[438]), .Z(n57591) );
  XOR U58229 ( .A(n40296), .B(n57591), .Z(n38634) );
  XOR U58230 ( .A(n57589), .B(n38634), .Z(n41896) );
  XOR U58231 ( .A(n41894), .B(n41896), .Z(n41899) );
  XOR U58232 ( .A(n41897), .B(n41899), .Z(n40291) );
  XOR U58233 ( .A(n40290), .B(n40291), .Z(n40294) );
  XOR U58234 ( .A(n40293), .B(n40294), .Z(n41903) );
  XOR U58235 ( .A(n41901), .B(n41903), .Z(n41906) );
  XOR U58236 ( .A(n41904), .B(n41906), .Z(n40288) );
  XOR U58237 ( .A(n40287), .B(n40288), .Z(n40282) );
  XOR U58238 ( .A(n40281), .B(n40282), .Z(n40286) );
  XOR U58239 ( .A(n40284), .B(n40286), .Z(n40279) );
  XOR U58240 ( .A(n40277), .B(n40279), .Z(n41911) );
  XOR U58241 ( .A(n41910), .B(n41911), .Z(n41914) );
  XOR U58242 ( .A(n41913), .B(n41914), .Z(n41918) );
  XOR U58243 ( .A(n41917), .B(n41918), .Z(n41922) );
  XOR U58244 ( .A(n41920), .B(n41922), .Z(n41926) );
  XOR U58245 ( .A(n41924), .B(n41926), .Z(n41928) );
  XOR U58246 ( .A(n41927), .B(n41928), .Z(n40275) );
  XOR U58247 ( .A(n40274), .B(n40275), .Z(n41935) );
  XOR U58248 ( .A(n41934), .B(n41935), .Z(n40273) );
  XOR U58249 ( .A(n40271), .B(n40273), .Z(n41942) );
  XOR U58250 ( .A(n41940), .B(n41942), .Z(n41944) );
  XOR U58251 ( .A(n41943), .B(n41944), .Z(n41949) );
  XOR U58252 ( .A(n41947), .B(n41949), .Z(n41952) );
  XOR U58253 ( .A(n41950), .B(n41952), .Z(n41955) );
  XOR U58254 ( .A(n41953), .B(n41955), .Z(n41957) );
  XOR U58255 ( .A(n41956), .B(n41957), .Z(n40265) );
  XOR U58256 ( .A(n40264), .B(n40265), .Z(n40268) );
  XOR U58257 ( .A(n40267), .B(n40268), .Z(n41962) );
  XOR U58258 ( .A(n41960), .B(n41962), .Z(n41964) );
  XOR U58259 ( .A(n41963), .B(n41964), .Z(n41968) );
  XOR U58260 ( .A(n41967), .B(n41968), .Z(n41971) );
  XOR U58261 ( .A(n41970), .B(n41971), .Z(n41975) );
  XOR U58262 ( .A(n41974), .B(n41975), .Z(n41978) );
  XOR U58263 ( .A(n41977), .B(n41978), .Z(n40259) );
  XOR U58264 ( .A(n40258), .B(n40259), .Z(n40263) );
  XOR U58265 ( .A(n40261), .B(n40263), .Z(n40256) );
  XOR U58266 ( .A(n40254), .B(n40256), .Z(n41982) );
  XOR U58267 ( .A(n41981), .B(n41982), .Z(n41986) );
  XOR U58268 ( .A(n41984), .B(n41986), .Z(n41990) );
  XOR U58269 ( .A(n41988), .B(n41990), .Z(n41993) );
  XOR U58270 ( .A(n41991), .B(n41993), .Z(n40252) );
  XOR U58271 ( .A(n40251), .B(n40252), .Z(n41995) );
  XOR U58272 ( .A(n41994), .B(n41995), .Z(n41999) );
  XOR U58273 ( .A(n41997), .B(n41999), .Z(n42004) );
  XOR U58274 ( .A(n42002), .B(n42004), .Z(n42006) );
  XOR U58275 ( .A(n42005), .B(n42006), .Z(n40249) );
  XOR U58276 ( .A(n40248), .B(n40249), .Z(n40244) );
  XOR U58277 ( .A(n40242), .B(n40244), .Z(n40247) );
  XOR U58278 ( .A(n40245), .B(n40247), .Z(n42017) );
  XOR U58279 ( .A(n42015), .B(n42017), .Z(n42020) );
  XOR U58280 ( .A(n42018), .B(n42020), .Z(n42023) );
  XOR U58281 ( .A(n42022), .B(n42023), .Z(n42026) );
  XOR U58282 ( .A(n42025), .B(n42026), .Z(n40238) );
  XOR U58283 ( .A(n40236), .B(n40238), .Z(n40241) );
  XOR U58284 ( .A(n40239), .B(n40241), .Z(n42034) );
  XOR U58285 ( .A(n42032), .B(n42034), .Z(n40234) );
  XOR U58286 ( .A(n40233), .B(n40234), .Z(n42044) );
  XOR U58287 ( .A(n42043), .B(n42044), .Z(n42048) );
  XOR U58288 ( .A(n42046), .B(n42048), .Z(n40232) );
  XOR U58289 ( .A(n40230), .B(n40232), .Z(n42054) );
  XOR U58290 ( .A(n42052), .B(n42054), .Z(n40228) );
  XOR U58291 ( .A(n40227), .B(n40228), .Z(n40223) );
  XOR U58292 ( .A(n40221), .B(n40223), .Z(n40226) );
  XOR U58293 ( .A(n40224), .B(n40226), .Z(n42061) );
  XOR U58294 ( .A(n42059), .B(n42061), .Z(n42063) );
  XOR U58295 ( .A(n42062), .B(n42063), .Z(n40219) );
  XOR U58296 ( .A(n40218), .B(n40219), .Z(n40214) );
  XOR U58297 ( .A(n40212), .B(n40214), .Z(n40216) );
  XOR U58298 ( .A(n40215), .B(n40216), .Z(n42069) );
  XOR U58299 ( .A(n42068), .B(n42069), .Z(n42073) );
  XOR U58300 ( .A(n42071), .B(n42073), .Z(n42076) );
  XOR U58301 ( .A(n42075), .B(n42076), .Z(n42080) );
  XOR U58302 ( .A(n42078), .B(n42080), .Z(n40210) );
  XOR U58303 ( .A(n40209), .B(n40210), .Z(n42084) );
  XOR U58304 ( .A(n42083), .B(n42084), .Z(n42088) );
  XOR U58305 ( .A(n42086), .B(n42088), .Z(n42092) );
  XOR U58306 ( .A(n42090), .B(n42092), .Z(n42095) );
  XOR U58307 ( .A(n42093), .B(n42095), .Z(n40207) );
  XOR U58308 ( .A(n40206), .B(n40207), .Z(n40201) );
  XOR U58309 ( .A(n40199), .B(n40201), .Z(n40204) );
  XOR U58310 ( .A(n40202), .B(n40204), .Z(n40195) );
  XOR U58311 ( .A(n40194), .B(n40195), .Z(n40197) );
  XOR U58312 ( .A(n40198), .B(n40197), .Z(n40191) );
  XOR U58313 ( .A(n40192), .B(n40191), .Z(n42099) );
  XOR U58314 ( .A(n42097), .B(n42099), .Z(n42101) );
  XOR U58315 ( .A(n42100), .B(n42101), .Z(n42107) );
  XOR U58316 ( .A(n42105), .B(n42107), .Z(n42110) );
  XOR U58317 ( .A(n42108), .B(n42110), .Z(n40190) );
  XOR U58318 ( .A(n40188), .B(n40190), .Z(n42119) );
  XOR U58319 ( .A(n42118), .B(n42119), .Z(n40186) );
  XOR U58320 ( .A(n40185), .B(n40186), .Z(n42133) );
  XOR U58321 ( .A(n42131), .B(n42133), .Z(n40184) );
  XOR U58322 ( .A(n40182), .B(n40184), .Z(n40177) );
  XOR U58323 ( .A(n40176), .B(n40177), .Z(n40181) );
  XOR U58324 ( .A(n40179), .B(n40181), .Z(n42143) );
  XOR U58325 ( .A(n42142), .B(n42143), .Z(n42144) );
  XOR U58326 ( .A(n42145), .B(n42144), .Z(n40174) );
  XOR U58327 ( .A(n40173), .B(n40174), .Z(n40168) );
  XOR U58328 ( .A(n40167), .B(n40168), .Z(n40172) );
  XOR U58329 ( .A(n40170), .B(n40172), .Z(n40163) );
  XOR U58330 ( .A(n40161), .B(n40163), .Z(n40165) );
  XOR U58331 ( .A(n40164), .B(n40165), .Z(n40160) );
  XOR U58332 ( .A(n40158), .B(n40160), .Z(n42155) );
  XOR U58333 ( .A(n42153), .B(n42155), .Z(n40156) );
  XOR U58334 ( .A(n40155), .B(n40156), .Z(n42162) );
  XOR U58335 ( .A(n42161), .B(n42162), .Z(n40153) );
  XOR U58336 ( .A(n40152), .B(n40153), .Z(n40148) );
  XOR U58337 ( .A(n40147), .B(n40148), .Z(n40149) );
  XOR U58338 ( .A(n40151), .B(n40149), .Z(n40143) );
  XOR U58339 ( .A(n40141), .B(n40143), .Z(n40146) );
  XOR U58340 ( .A(n40144), .B(n40146), .Z(n42176) );
  XOR U58341 ( .A(n42175), .B(n42176), .Z(n42180) );
  XOR U58342 ( .A(n42178), .B(n42180), .Z(n42184) );
  XOR U58343 ( .A(n42182), .B(n42184), .Z(n42187) );
  XOR U58344 ( .A(n42185), .B(n42187), .Z(n40136) );
  XOR U58345 ( .A(n40135), .B(n40136), .Z(n40139) );
  XOR U58346 ( .A(n40138), .B(n40139), .Z(n42192) );
  XOR U58347 ( .A(n42190), .B(n42192), .Z(n42195) );
  XOR U58348 ( .A(n42193), .B(n42195), .Z(n42197) );
  XOR U58349 ( .A(n42196), .B(n42197), .Z(n42198) );
  XOR U58350 ( .A(n42199), .B(n42198), .Z(n40133) );
  XOR U58351 ( .A(n40132), .B(n40133), .Z(n40127) );
  XOR U58352 ( .A(n40125), .B(n40127), .Z(n40130) );
  XOR U58353 ( .A(n40128), .B(n40130), .Z(n40120) );
  XOR U58354 ( .A(n40119), .B(n40120), .Z(n40123) );
  XOR U58355 ( .A(n40122), .B(n40123), .Z(n42205) );
  XOR U58356 ( .A(n42203), .B(n42205), .Z(n42208) );
  XOR U58357 ( .A(n42206), .B(n42208), .Z(n40118) );
  XOR U58358 ( .A(n40116), .B(n40118), .Z(n40112) );
  XOR U58359 ( .A(n40110), .B(n40112), .Z(n40114) );
  XOR U58360 ( .A(n40113), .B(n40114), .Z(n40105) );
  XOR U58361 ( .A(n40106), .B(n40105), .Z(n40107) );
  XOR U58362 ( .A(n40109), .B(n40107), .Z(n40101) );
  XOR U58363 ( .A(n40099), .B(n40101), .Z(n40104) );
  XOR U58364 ( .A(n40102), .B(n40104), .Z(n42215) );
  XOR U58365 ( .A(n42213), .B(n42215), .Z(n42218) );
  XOR U58366 ( .A(n42216), .B(n42218), .Z(n40097) );
  XOR U58367 ( .A(n40096), .B(n40097), .Z(n42223) );
  XOR U58368 ( .A(n42222), .B(n42223), .Z(n40095) );
  XOR U58369 ( .A(n40093), .B(n40095), .Z(n40091) );
  XOR U58370 ( .A(n40090), .B(n40091), .Z(n40085) );
  XOR U58371 ( .A(n40086), .B(n40085), .Z(n45509) );
  XOR U58372 ( .A(n45507), .B(n45509), .Z(n40082) );
  XOR U58373 ( .A(n40081), .B(n40082), .Z(n42235) );
  XOR U58374 ( .A(n42233), .B(n42235), .Z(n40079) );
  XOR U58375 ( .A(n40078), .B(n40079), .Z(n40074) );
  XOR U58376 ( .A(n40072), .B(n40074), .Z(n40076) );
  XOR U58377 ( .A(n40075), .B(n40076), .Z(n40070) );
  XOR U58378 ( .A(n40069), .B(n40070), .Z(n42242) );
  XOR U58379 ( .A(n42240), .B(n42242), .Z(n42245) );
  XOR U58380 ( .A(n42243), .B(n42245), .Z(n42248) );
  XOR U58381 ( .A(n42247), .B(n42248), .Z(n42252) );
  XOR U58382 ( .A(n42250), .B(n42252), .Z(n40067) );
  XOR U58383 ( .A(n40066), .B(n40067), .Z(n42256) );
  XOR U58384 ( .A(n42254), .B(n42256), .Z(n42258) );
  XOR U58385 ( .A(n42257), .B(n42258), .Z(n40064) );
  XOR U58386 ( .A(n40063), .B(n40064), .Z(n42266) );
  XOR U58387 ( .A(n42265), .B(n42266), .Z(n40060) );
  XOR U58388 ( .A(n40059), .B(n40060), .Z(n42264) );
  XOR U58389 ( .A(n42262), .B(n42264), .Z(n42276) );
  XOR U58390 ( .A(n42275), .B(n42276), .Z(n42279) );
  XOR U58391 ( .A(n42278), .B(n42279), .Z(n42282) );
  XOR U58392 ( .A(n42281), .B(n42282), .Z(n42286) );
  XOR U58393 ( .A(n42284), .B(n42286), .Z(n40058) );
  XOR U58394 ( .A(n40056), .B(n40058), .Z(n42290) );
  XOR U58395 ( .A(n42289), .B(n42290), .Z(n42294) );
  XOR U58396 ( .A(n42292), .B(n42294), .Z(n42298) );
  XOR U58397 ( .A(n42296), .B(n42298), .Z(n42300) );
  XOR U58398 ( .A(n42299), .B(n42300), .Z(n40054) );
  XOR U58399 ( .A(n40053), .B(n40054), .Z(n42304) );
  XOR U58400 ( .A(n42303), .B(n42304), .Z(n42308) );
  XOR U58401 ( .A(n42306), .B(n42308), .Z(n42311) );
  XOR U58402 ( .A(n42310), .B(n42311), .Z(n42315) );
  XOR U58403 ( .A(n42313), .B(n42315), .Z(n40052) );
  XOR U58404 ( .A(n40050), .B(n40052), .Z(n42319) );
  XOR U58405 ( .A(n42317), .B(n42319), .Z(n42322) );
  XOR U58406 ( .A(n42320), .B(n42322), .Z(n42326) );
  XOR U58407 ( .A(n42324), .B(n42326), .Z(n42329) );
  XOR U58408 ( .A(n42327), .B(n42329), .Z(n42332) );
  XOR U58409 ( .A(n42331), .B(n42332), .Z(n42335) );
  XOR U58410 ( .A(n42334), .B(n42335), .Z(n42340) );
  XOR U58411 ( .A(n42338), .B(n42340), .Z(n42343) );
  XOR U58412 ( .A(n42341), .B(n42343), .Z(n40046) );
  XOR U58413 ( .A(n40044), .B(n40046), .Z(n40049) );
  XOR U58414 ( .A(n40047), .B(n40049), .Z(n40039) );
  XOR U58415 ( .A(n40038), .B(n40039), .Z(n40042) );
  XOR U58416 ( .A(n40041), .B(n40042), .Z(n40037) );
  XOR U58417 ( .A(n40035), .B(n40037), .Z(n40031) );
  XOR U58418 ( .A(n40029), .B(n40031), .Z(n40033) );
  XOR U58419 ( .A(n40032), .B(n40033), .Z(n42365) );
  XOR U58420 ( .A(n42363), .B(n42365), .Z(n42368) );
  XOR U58421 ( .A(n42366), .B(n42368), .Z(n40027) );
  XOR U58422 ( .A(n40026), .B(n40027), .Z(n42371) );
  XOR U58423 ( .A(n42370), .B(n42371), .Z(n42375) );
  XOR U58424 ( .A(n42373), .B(n42375), .Z(n40021) );
  XOR U58425 ( .A(n40020), .B(n40021), .Z(n40025) );
  XOR U58426 ( .A(n40023), .B(n40025), .Z(n40019) );
  XOR U58427 ( .A(n40017), .B(n40019), .Z(n40013) );
  XOR U58428 ( .A(n40011), .B(n40013), .Z(n40016) );
  XOR U58429 ( .A(n40014), .B(n40016), .Z(n40009) );
  XOR U58430 ( .A(n40007), .B(n40009), .Z(n42379) );
  XOR U58431 ( .A(n42378), .B(n42379), .Z(n42382) );
  XOR U58432 ( .A(n42381), .B(n42382), .Z(n40002) );
  XOR U58433 ( .A(n40001), .B(n40002), .Z(n40005) );
  XOR U58434 ( .A(n40004), .B(n40005), .Z(n42386) );
  XOR U58435 ( .A(n42385), .B(n42386), .Z(n42390) );
  XOR U58436 ( .A(n42388), .B(n42390), .Z(n42393) );
  XOR U58437 ( .A(n42392), .B(n42393), .Z(n42397) );
  XOR U58438 ( .A(n42395), .B(n42397), .Z(n39997) );
  XOR U58439 ( .A(n39995), .B(n39997), .Z(n40000) );
  XOR U58440 ( .A(n39998), .B(n40000), .Z(n39992) );
  XOR U58441 ( .A(n39991), .B(n39992), .Z(n39986) );
  XOR U58442 ( .A(n39985), .B(n39986), .Z(n39990) );
  XOR U58443 ( .A(n39988), .B(n39990), .Z(n39984) );
  XOR U58444 ( .A(n39982), .B(n39984), .Z(n42403) );
  XOR U58445 ( .A(n42401), .B(n42403), .Z(n42406) );
  XOR U58446 ( .A(n42404), .B(n42406), .Z(n42410) );
  XOR U58447 ( .A(n42408), .B(n42410), .Z(n42412) );
  XOR U58448 ( .A(n42411), .B(n42412), .Z(n42415) );
  XOR U58449 ( .A(n42414), .B(n42415), .Z(n42418) );
  XOR U58450 ( .A(n42417), .B(n42418), .Z(n42423) );
  XOR U58451 ( .A(n42421), .B(n42423), .Z(n42426) );
  XOR U58452 ( .A(n42424), .B(n42426), .Z(n39978) );
  XOR U58453 ( .A(n39976), .B(n39978), .Z(n39981) );
  XOR U58454 ( .A(n39979), .B(n39981), .Z(n39971) );
  XOR U58455 ( .A(n39970), .B(n39971), .Z(n39975) );
  XOR U58456 ( .A(n39973), .B(n39975), .Z(n42432) );
  XOR U58457 ( .A(n42430), .B(n42432), .Z(n42434) );
  XOR U58458 ( .A(n42433), .B(n42434), .Z(n42438) );
  XOR U58459 ( .A(n42437), .B(n42438), .Z(n42442) );
  XOR U58460 ( .A(n42440), .B(n42442), .Z(n39966) );
  XOR U58461 ( .A(n39964), .B(n39966), .Z(n39969) );
  XOR U58462 ( .A(n39967), .B(n39969), .Z(n39959) );
  XOR U58463 ( .A(n39958), .B(n39959), .Z(n39962) );
  XOR U58464 ( .A(n39961), .B(n39962), .Z(n39954) );
  XOR U58465 ( .A(n39952), .B(n39954), .Z(n39956) );
  XOR U58466 ( .A(n39955), .B(n39956), .Z(n39948) );
  XOR U58467 ( .A(n39946), .B(n39948), .Z(n39951) );
  XOR U58468 ( .A(n39949), .B(n39951), .Z(n39942) );
  XOR U58469 ( .A(n39940), .B(n39942), .Z(n39945) );
  XOR U58470 ( .A(n39943), .B(n39945), .Z(n42449) );
  XOR U58471 ( .A(n42448), .B(n42449), .Z(n42452) );
  XOR U58472 ( .A(n42451), .B(n42452), .Z(n39936) );
  XOR U58473 ( .A(n39934), .B(n39936), .Z(n39939) );
  XOR U58474 ( .A(n39937), .B(n39939), .Z(n39930) );
  XOR U58475 ( .A(n39928), .B(n39930), .Z(n39933) );
  XOR U58476 ( .A(n39931), .B(n39933), .Z(n42457) );
  XOR U58477 ( .A(n42456), .B(n42457), .Z(n42460) );
  XOR U58478 ( .A(n42459), .B(n42460), .Z(n42465) );
  XOR U58479 ( .A(n42464), .B(n42465), .Z(n42469) );
  XOR U58480 ( .A(n42467), .B(n42469), .Z(n42473) );
  XOR U58481 ( .A(n42471), .B(n42473), .Z(n42476) );
  XOR U58482 ( .A(n42474), .B(n42476), .Z(n39926) );
  XOR U58483 ( .A(n39925), .B(n39926), .Z(n39920) );
  XOR U58484 ( .A(n39919), .B(n39920), .Z(n39924) );
  XOR U58485 ( .A(n39922), .B(n39924), .Z(n42480) );
  XOR U58486 ( .A(n42478), .B(n42480), .Z(n42482) );
  XOR U58487 ( .A(n42481), .B(n42482), .Z(n39917) );
  XOR U58488 ( .A(n39916), .B(n39917), .Z(n39912) );
  XOR U58489 ( .A(n39910), .B(n39912), .Z(n39914) );
  XOR U58490 ( .A(n39913), .B(n39914), .Z(n39905) );
  XOR U58491 ( .A(n39904), .B(n39905), .Z(n39908) );
  XOR U58492 ( .A(n39907), .B(n39908), .Z(n39899) );
  XOR U58493 ( .A(n39898), .B(n39899), .Z(n39902) );
  XOR U58494 ( .A(n39901), .B(n39902), .Z(n42487) );
  XOR U58495 ( .A(n42486), .B(n42487), .Z(n42491) );
  XOR U58496 ( .A(n42489), .B(n42491), .Z(n39894) );
  XOR U58497 ( .A(n39892), .B(n39894), .Z(n39896) );
  XOR U58498 ( .A(n39895), .B(n39896), .Z(n42495) );
  XOR U58499 ( .A(n42493), .B(n42495), .Z(n42498) );
  XOR U58500 ( .A(n42496), .B(n42498), .Z(n42502) );
  XOR U58501 ( .A(n42500), .B(n42502), .Z(n42505) );
  XOR U58502 ( .A(n42503), .B(n42505), .Z(n42508) );
  XOR U58503 ( .A(n42507), .B(n42508), .Z(n42511) );
  XOR U58504 ( .A(n42510), .B(n42511), .Z(n42516) );
  XOR U58505 ( .A(n42514), .B(n42516), .Z(n42519) );
  XOR U58506 ( .A(n42517), .B(n42519), .Z(n42521) );
  XOR U58507 ( .A(n42520), .B(n42521), .Z(n42525) );
  XOR U58508 ( .A(n42523), .B(n42525), .Z(n39888) );
  XOR U58509 ( .A(n39886), .B(n39888), .Z(n39891) );
  XOR U58510 ( .A(n39889), .B(n39891), .Z(n42527) );
  XOR U58511 ( .A(n42526), .B(n42527), .Z(n42531) );
  XOR U58512 ( .A(n42529), .B(n42531), .Z(n39885) );
  XOR U58513 ( .A(n39883), .B(n39885), .Z(n39878) );
  XOR U58514 ( .A(n39876), .B(n39878), .Z(n39880) );
  XOR U58515 ( .A(n39879), .B(n39880), .Z(n39875) );
  XOR U58516 ( .A(n39873), .B(n39875), .Z(n42536) );
  XOR U58517 ( .A(n42534), .B(n42536), .Z(n42538) );
  XOR U58518 ( .A(n42537), .B(n42538), .Z(n42542) );
  XOR U58519 ( .A(n42541), .B(n42542), .Z(n42545) );
  XOR U58520 ( .A(n42544), .B(n42545), .Z(n42549) );
  XOR U58521 ( .A(n42548), .B(n42549), .Z(n42552) );
  XOR U58522 ( .A(n42551), .B(n42552), .Z(n39869) );
  XOR U58523 ( .A(n39867), .B(n39869), .Z(n39872) );
  XOR U58524 ( .A(n39870), .B(n39872), .Z(n42556) );
  XOR U58525 ( .A(n42554), .B(n42556), .Z(n42558) );
  XOR U58526 ( .A(n42557), .B(n42558), .Z(n42564) );
  XOR U58527 ( .A(n42563), .B(n42564), .Z(n39865) );
  XOR U58528 ( .A(n39864), .B(n39865), .Z(n42577) );
  XOR U58529 ( .A(n42575), .B(n42577), .Z(n39862) );
  XOR U58530 ( .A(n39861), .B(n39862), .Z(n45259) );
  IV U58531 ( .A(n45259), .Z(n42587) );
  XOR U58532 ( .A(n45258), .B(n42587), .Z(n42588) );
  XOR U58533 ( .A(n42589), .B(n42588), .Z(n39860) );
  XOR U58534 ( .A(n39858), .B(n39860), .Z(n42594) );
  XOR U58535 ( .A(n42593), .B(n42594), .Z(n42597) );
  XOR U58536 ( .A(n42596), .B(n42597), .Z(n42602) );
  XOR U58537 ( .A(n42600), .B(n42602), .Z(n42604) );
  XOR U58538 ( .A(n42603), .B(n42604), .Z(n42608) );
  XOR U58539 ( .A(n42606), .B(n42608), .Z(n42611) );
  XOR U58540 ( .A(n42609), .B(n42611), .Z(n39855) );
  XOR U58541 ( .A(n39853), .B(n39855), .Z(n39856) );
  XOR U58542 ( .A(n39857), .B(n39856), .Z(n42613) );
  XOR U58543 ( .A(n42614), .B(n42613), .Z(n42616) );
  XOR U58544 ( .A(n42617), .B(n42616), .Z(n42618) );
  XOR U58545 ( .A(n42620), .B(n42618), .Z(n42623) );
  XOR U58546 ( .A(n42621), .B(n42623), .Z(n42625) );
  XOR U58547 ( .A(n42624), .B(n42625), .Z(n42628) );
  XOR U58548 ( .A(n42627), .B(n42628), .Z(n39847) );
  XOR U58549 ( .A(n39849), .B(n39847), .Z(n39852) );
  XOR U58550 ( .A(n39850), .B(n39852), .Z(n39843) );
  XOR U58551 ( .A(n39841), .B(n39843), .Z(n39845) );
  XOR U58552 ( .A(n39844), .B(n39845), .Z(n39839) );
  XOR U58553 ( .A(n39837), .B(n39839), .Z(n39833) );
  XOR U58554 ( .A(n39831), .B(n39833), .Z(n39835) );
  XOR U58555 ( .A(n39834), .B(n39835), .Z(n39826) );
  XOR U58556 ( .A(n39825), .B(n39826), .Z(n39830) );
  XOR U58557 ( .A(n39828), .B(n39830), .Z(n39821) );
  XOR U58558 ( .A(n39819), .B(n39821), .Z(n39824) );
  XOR U58559 ( .A(n39822), .B(n39824), .Z(n42634) );
  XOR U58560 ( .A(n42633), .B(n42634), .Z(n42637) );
  XOR U58561 ( .A(n42636), .B(n42637), .Z(n47481) );
  XOR U58562 ( .A(n47479), .B(n47481), .Z(n42642) );
  XOR U58563 ( .A(n42643), .B(n42642), .Z(n39815) );
  XOR U58564 ( .A(n39813), .B(n39815), .Z(n39817) );
  XOR U58565 ( .A(n39816), .B(n39817), .Z(n42649) );
  XOR U58566 ( .A(n42647), .B(n42649), .Z(n42652) );
  XOR U58567 ( .A(n42650), .B(n42652), .Z(n42655) );
  XOR U58568 ( .A(n42654), .B(n42655), .Z(n42658) );
  XOR U58569 ( .A(n42657), .B(n42658), .Z(n39809) );
  XOR U58570 ( .A(n39807), .B(n39809), .Z(n39812) );
  XOR U58571 ( .A(n39810), .B(n39812), .Z(n39802) );
  XOR U58572 ( .A(n39803), .B(n39802), .Z(n39804) );
  XOR U58573 ( .A(n39805), .B(n39804), .Z(n42662) );
  XOR U58574 ( .A(n42661), .B(n42662), .Z(n42663) );
  XOR U58575 ( .A(n42664), .B(n42663), .Z(n39796) );
  XOR U58576 ( .A(n39797), .B(n39796), .Z(n39798) );
  XOR U58577 ( .A(n39800), .B(n39798), .Z(n42667) );
  XOR U58578 ( .A(n42666), .B(n42667), .Z(n42668) );
  XOR U58579 ( .A(n42669), .B(n42668), .Z(n39792) );
  XOR U58580 ( .A(n39791), .B(n39792), .Z(n39793) );
  XOR U58581 ( .A(n39794), .B(n39793), .Z(n42674) );
  XOR U58582 ( .A(n42672), .B(n42674), .Z(n42677) );
  XOR U58583 ( .A(n42675), .B(n42677), .Z(n42681) );
  XOR U58584 ( .A(n42682), .B(n42681), .Z(n39788) );
  XOR U58585 ( .A(n39790), .B(n39788), .Z(n42692) );
  XOR U58586 ( .A(n42690), .B(n42692), .Z(n42694) );
  XOR U58587 ( .A(n42693), .B(n42694), .Z(n42697) );
  XOR U58588 ( .A(n42698), .B(n42697), .Z(n42699) );
  XOR U58589 ( .A(n42700), .B(n42699), .Z(n39786) );
  XOR U58590 ( .A(n39785), .B(n39786), .Z(n42706) );
  XOR U58591 ( .A(n42704), .B(n42706), .Z(n42707) );
  XOR U58592 ( .A(n42708), .B(n42707), .Z(n39782) );
  XOR U58593 ( .A(n39784), .B(n39782), .Z(n39777) );
  XOR U58594 ( .A(n39775), .B(n39777), .Z(n39779) );
  XOR U58595 ( .A(n39778), .B(n39779), .Z(n39774) );
  XOR U58596 ( .A(n39773), .B(n39774), .Z(n42712) );
  XOR U58597 ( .A(n42713), .B(n42712), .Z(n42716) );
  XOR U58598 ( .A(n42715), .B(n42716), .Z(n42722) );
  XOR U58599 ( .A(n42720), .B(n42722), .Z(n42724) );
  XOR U58600 ( .A(n42723), .B(n42724), .Z(n42726) );
  XOR U58601 ( .A(n42727), .B(n42726), .Z(n42730) );
  XOR U58602 ( .A(n42729), .B(n42730), .Z(n42735) );
  XOR U58603 ( .A(n42733), .B(n42735), .Z(n42737) );
  XOR U58604 ( .A(n42736), .B(n42737), .Z(n42739) );
  XOR U58605 ( .A(n42740), .B(n42739), .Z(n42744) );
  XOR U58606 ( .A(n42742), .B(n42744), .Z(n39770) );
  XOR U58607 ( .A(n39768), .B(n39770), .Z(n39771) );
  XOR U58608 ( .A(n39772), .B(n39771), .Z(n39765) );
  XOR U58609 ( .A(n39767), .B(n39765), .Z(n39761) );
  XOR U58610 ( .A(n39759), .B(n39761), .Z(n39764) );
  XOR U58611 ( .A(n39762), .B(n39764), .Z(n39755) );
  XOR U58612 ( .A(n39754), .B(n39755), .Z(n39756) );
  XOR U58613 ( .A(n39757), .B(n39756), .Z(n39752) );
  XOR U58614 ( .A(n39751), .B(n39752), .Z(n39747) );
  XOR U58615 ( .A(n39745), .B(n39747), .Z(n39749) );
  XOR U58616 ( .A(n39748), .B(n39749), .Z(n39740) );
  XOR U58617 ( .A(n39739), .B(n39740), .Z(n39744) );
  XOR U58618 ( .A(n39742), .B(n39744), .Z(n39735) );
  XOR U58619 ( .A(n39733), .B(n39735), .Z(n39737) );
  XOR U58620 ( .A(n39736), .B(n39737), .Z(n42755) );
  XOR U58621 ( .A(n42753), .B(n42755), .Z(n42758) );
  XOR U58622 ( .A(n42756), .B(n42758), .Z(n39727) );
  XOR U58623 ( .A(n39726), .B(n39727), .Z(n39730) );
  XOR U58624 ( .A(n39729), .B(n39730), .Z(n39724) );
  XOR U58625 ( .A(n39723), .B(n39724), .Z(n47587) );
  XOR U58626 ( .A(n47586), .B(n47587), .Z(n42761) );
  XOR U58627 ( .A(n47599), .B(n42761), .Z(n42767) );
  XOR U58628 ( .A(n42765), .B(n42767), .Z(n42769) );
  XOR U58629 ( .A(n42768), .B(n42769), .Z(n42774) );
  XOR U58630 ( .A(n42772), .B(n42774), .Z(n42777) );
  XOR U58631 ( .A(n42775), .B(n42777), .Z(n42780) );
  XOR U58632 ( .A(n42779), .B(n42780), .Z(n42784) );
  XOR U58633 ( .A(n42782), .B(n42784), .Z(n39719) );
  XOR U58634 ( .A(n39717), .B(n39719), .Z(n39721) );
  XOR U58635 ( .A(n39720), .B(n39721), .Z(n42787) );
  XOR U58636 ( .A(n42786), .B(n42787), .Z(n42791) );
  XOR U58637 ( .A(n42789), .B(n42791), .Z(n39716) );
  XOR U58638 ( .A(n39714), .B(n39716), .Z(n42798) );
  XOR U58639 ( .A(n42796), .B(n42798), .Z(n39712) );
  XOR U58640 ( .A(n39711), .B(n39712), .Z(n42803) );
  XOR U58641 ( .A(n42802), .B(n42803), .Z(n42807) );
  XOR U58642 ( .A(n42805), .B(n42807), .Z(n39707) );
  XOR U58643 ( .A(n39705), .B(n39707), .Z(n39709) );
  XOR U58644 ( .A(n39708), .B(n39709), .Z(n39703) );
  XOR U58645 ( .A(n39702), .B(n39703), .Z(n42812) );
  XOR U58646 ( .A(n42810), .B(n42812), .Z(n42815) );
  XOR U58647 ( .A(n42813), .B(n42815), .Z(n42819) );
  XOR U58648 ( .A(n42817), .B(n42819), .Z(n42822) );
  XOR U58649 ( .A(n42820), .B(n42822), .Z(n42824) );
  XOR U58650 ( .A(n42823), .B(n42824), .Z(n42827) );
  XOR U58651 ( .A(n42826), .B(n42827), .Z(n42832) );
  XOR U58652 ( .A(n42830), .B(n42832), .Z(n42835) );
  XOR U58653 ( .A(n42833), .B(n42835), .Z(n42838) );
  XOR U58654 ( .A(n42837), .B(n42838), .Z(n42842) );
  XOR U58655 ( .A(n42840), .B(n42842), .Z(n39697) );
  XOR U58656 ( .A(n39696), .B(n39697), .Z(n39700) );
  XOR U58657 ( .A(n39699), .B(n39700), .Z(n42846) );
  XOR U58658 ( .A(n42845), .B(n42846), .Z(n55410) );
  XOR U58659 ( .A(n55409), .B(n55410), .Z(n42851) );
  XOR U58660 ( .A(n42850), .B(n42851), .Z(n42855) );
  XOR U58661 ( .A(n42853), .B(n42855), .Z(n39692) );
  XOR U58662 ( .A(n39690), .B(n39692), .Z(n39695) );
  XOR U58663 ( .A(n39693), .B(n39695), .Z(n42859) );
  XOR U58664 ( .A(n42858), .B(n42859), .Z(n42862) );
  XOR U58665 ( .A(n42861), .B(n42862), .Z(n42867) );
  XOR U58666 ( .A(n42865), .B(n42867), .Z(n42870) );
  XOR U58667 ( .A(n42868), .B(n42870), .Z(n42872) );
  XOR U58668 ( .A(n42871), .B(n42872), .Z(n42876) );
  XOR U58669 ( .A(n42874), .B(n42876), .Z(n39685) );
  XOR U58670 ( .A(n39684), .B(n39685), .Z(n39689) );
  XOR U58671 ( .A(n39687), .B(n39689), .Z(n42879) );
  XOR U58672 ( .A(n42878), .B(n42879), .Z(n42882) );
  XOR U58673 ( .A(n42881), .B(n42882), .Z(n39680) );
  XOR U58674 ( .A(n39678), .B(n39680), .Z(n39683) );
  XOR U58675 ( .A(n39681), .B(n39683), .Z(n39676) );
  XOR U58676 ( .A(n39675), .B(n39676), .Z(n42888) );
  XOR U58677 ( .A(n42886), .B(n42888), .Z(n42891) );
  XOR U58678 ( .A(n42889), .B(n42891), .Z(n42905) );
  XOR U58679 ( .A(n42903), .B(n42905), .Z(n42907) );
  XOR U58680 ( .A(n42906), .B(n42907), .Z(n42910) );
  XOR U58681 ( .A(n42909), .B(n42910), .Z(n42914) );
  XOR U58682 ( .A(n42912), .B(n42914), .Z(n42918) );
  XOR U58683 ( .A(n42916), .B(n42918), .Z(n42920) );
  XOR U58684 ( .A(n42919), .B(n42920), .Z(n42925) );
  XOR U58685 ( .A(n42923), .B(n42925), .Z(n42927) );
  XOR U58686 ( .A(n42926), .B(n42927), .Z(n42932) );
  XOR U58687 ( .A(n42930), .B(n42932), .Z(n42934) );
  XOR U58688 ( .A(n42933), .B(n42934), .Z(n42938) );
  XOR U58689 ( .A(n42937), .B(n42938), .Z(n42942) );
  XOR U58690 ( .A(n42940), .B(n42942), .Z(n39673) );
  XOR U58691 ( .A(n39672), .B(n39673), .Z(n42948) );
  XOR U58692 ( .A(n42946), .B(n42948), .Z(n39671) );
  XOR U58693 ( .A(n39669), .B(n39671), .Z(n42958) );
  XOR U58694 ( .A(n42956), .B(n42958), .Z(n39668) );
  XOR U58695 ( .A(n39666), .B(n39668), .Z(n39664) );
  XOR U58696 ( .A(n39662), .B(n39664), .Z(n42970) );
  XOR U58697 ( .A(n42968), .B(n42970), .Z(n42972) );
  XOR U58698 ( .A(n42971), .B(n42972), .Z(n39657) );
  XOR U58699 ( .A(n39656), .B(n39657), .Z(n39661) );
  XOR U58700 ( .A(n39659), .B(n39661), .Z(n42980) );
  XOR U58701 ( .A(n42978), .B(n42980), .Z(n39653) );
  XOR U58702 ( .A(n39652), .B(n39653), .Z(n42977) );
  XOR U58703 ( .A(n42975), .B(n42977), .Z(n42988) );
  XOR U58704 ( .A(n42986), .B(n42988), .Z(n42995) );
  XOR U58705 ( .A(n42993), .B(n42995), .Z(n39649) );
  XOR U58706 ( .A(n39648), .B(n39649), .Z(n42991) );
  XOR U58707 ( .A(n42990), .B(n42991), .Z(n43003) );
  XOR U58708 ( .A(n43001), .B(n43003), .Z(n43006) );
  XOR U58709 ( .A(n43004), .B(n43006), .Z(n39644) );
  XOR U58710 ( .A(n39642), .B(n39644), .Z(n39647) );
  XOR U58711 ( .A(n39645), .B(n39647), .Z(n43009) );
  XOR U58712 ( .A(n43008), .B(n43009), .Z(n43013) );
  XOR U58713 ( .A(n43011), .B(n43013), .Z(n39640) );
  XOR U58714 ( .A(n39638), .B(n39640), .Z(n43016) );
  XOR U58715 ( .A(n43015), .B(n43016), .Z(n43019) );
  XOR U58716 ( .A(n43018), .B(n43019), .Z(n39634) );
  XOR U58717 ( .A(n39632), .B(n39634), .Z(n39636) );
  XOR U58718 ( .A(n39635), .B(n39636), .Z(n39628) );
  XOR U58719 ( .A(n39626), .B(n39628), .Z(n39630) );
  XOR U58720 ( .A(n39629), .B(n39630), .Z(n43023) );
  XOR U58721 ( .A(n43022), .B(n43023), .Z(n43027) );
  XOR U58722 ( .A(n43025), .B(n43027), .Z(n39624) );
  XOR U58723 ( .A(n39623), .B(n39624), .Z(n39619) );
  XOR U58724 ( .A(n39617), .B(n39619), .Z(n39621) );
  XOR U58725 ( .A(n39620), .B(n39621), .Z(n39612) );
  XOR U58726 ( .A(n39611), .B(n39612), .Z(n39616) );
  XOR U58727 ( .A(n39614), .B(n39616), .Z(n39609) );
  XOR U58728 ( .A(n39607), .B(n39609), .Z(n43035) );
  XOR U58729 ( .A(n43033), .B(n43035), .Z(n39605) );
  XOR U58730 ( .A(n39604), .B(n39605), .Z(n39602) );
  XOR U58731 ( .A(n39601), .B(n39602), .Z(n43046) );
  XOR U58732 ( .A(n43045), .B(n43046), .Z(n43050) );
  XOR U58733 ( .A(n43048), .B(n43050), .Z(n39600) );
  XOR U58734 ( .A(n39598), .B(n39600), .Z(n39594) );
  XOR U58735 ( .A(n39592), .B(n39594), .Z(n39597) );
  XOR U58736 ( .A(n39595), .B(n39597), .Z(n43056) );
  XOR U58737 ( .A(n43054), .B(n43056), .Z(n43058) );
  XOR U58738 ( .A(n43057), .B(n43058), .Z(n39590) );
  XOR U58739 ( .A(n39589), .B(n39590), .Z(n39585) );
  XOR U58740 ( .A(n39583), .B(n39585), .Z(n39588) );
  XOR U58741 ( .A(n39586), .B(n39588), .Z(n39578) );
  XOR U58742 ( .A(n39577), .B(n39578), .Z(n39582) );
  XOR U58743 ( .A(n39580), .B(n39582), .Z(n39576) );
  XOR U58744 ( .A(n39574), .B(n39576), .Z(n39570) );
  XOR U58745 ( .A(n39568), .B(n39570), .Z(n39572) );
  XOR U58746 ( .A(n39571), .B(n39572), .Z(n39562) );
  XOR U58747 ( .A(n39561), .B(n39562), .Z(n39566) );
  XOR U58748 ( .A(n39564), .B(n39566), .Z(n39557) );
  XOR U58749 ( .A(n39555), .B(n39557), .Z(n39559) );
  XOR U58750 ( .A(n39558), .B(n39559), .Z(n39553) );
  XOR U58751 ( .A(n39552), .B(n39553), .Z(n43070) );
  XOR U58752 ( .A(n43068), .B(n43070), .Z(n43072) );
  XOR U58753 ( .A(n43071), .B(n43072), .Z(n43076) );
  XOR U58754 ( .A(n43078), .B(n43076), .Z(n45062) );
  XOR U58755 ( .A(n43079), .B(n45062), .Z(n43085) );
  XOR U58756 ( .A(n43083), .B(n43085), .Z(n43088) );
  XOR U58757 ( .A(n43086), .B(n43088), .Z(n39547) );
  XOR U58758 ( .A(n39546), .B(n39547), .Z(n39551) );
  XOR U58759 ( .A(n39549), .B(n39551), .Z(n39541) );
  XOR U58760 ( .A(n39539), .B(n39541), .Z(n39544) );
  XOR U58761 ( .A(n39542), .B(n39544), .Z(n39537) );
  XOR U58762 ( .A(n39536), .B(n39537), .Z(n43094) );
  XOR U58763 ( .A(n43093), .B(n43094), .Z(n39535) );
  XOR U58764 ( .A(n39533), .B(n39535), .Z(n39532) );
  XOR U58765 ( .A(n39530), .B(n39532), .Z(n39525) );
  XOR U58766 ( .A(n39524), .B(n39525), .Z(n39529) );
  XOR U58767 ( .A(n39527), .B(n39529), .Z(n43107) );
  XOR U58768 ( .A(n43105), .B(n43107), .Z(n43110) );
  XOR U58769 ( .A(n43108), .B(n43110), .Z(n39520) );
  XOR U58770 ( .A(n39518), .B(n39520), .Z(n39523) );
  XOR U58771 ( .A(n39521), .B(n39523), .Z(n43115) );
  XOR U58772 ( .A(n43114), .B(n43115), .Z(n43119) );
  XOR U58773 ( .A(n43117), .B(n43119), .Z(n43123) );
  XOR U58774 ( .A(n43121), .B(n43123), .Z(n43125) );
  XOR U58775 ( .A(n43124), .B(n43125), .Z(n43129) );
  XOR U58776 ( .A(n43128), .B(n43129), .Z(n43132) );
  XOR U58777 ( .A(n43131), .B(n43132), .Z(n43137) );
  XOR U58778 ( .A(n43135), .B(n43137), .Z(n43140) );
  XOR U58779 ( .A(n43138), .B(n43140), .Z(n43143) );
  XOR U58780 ( .A(n43142), .B(n43143), .Z(n43147) );
  XOR U58781 ( .A(n43145), .B(n43147), .Z(n39517) );
  XOR U58782 ( .A(n39515), .B(n39517), .Z(n39511) );
  XOR U58783 ( .A(n39509), .B(n39511), .Z(n39513) );
  XOR U58784 ( .A(n39512), .B(n39513), .Z(n39504) );
  XOR U58785 ( .A(n39503), .B(n39504), .Z(n39508) );
  XOR U58786 ( .A(n39506), .B(n39508), .Z(n39495) );
  XOR U58787 ( .A(n39494), .B(n39495), .Z(n39499) );
  XOR U58788 ( .A(n39497), .B(n39499), .Z(n39502) );
  XOR U58789 ( .A(n39500), .B(n39502), .Z(n39490) );
  XOR U58790 ( .A(n39488), .B(n39490), .Z(n39492) );
  XOR U58791 ( .A(n39491), .B(n39492), .Z(n43157) );
  XOR U58792 ( .A(n43156), .B(n43157), .Z(n43160) );
  XOR U58793 ( .A(n43159), .B(n43160), .Z(n39487) );
  XOR U58794 ( .A(n39485), .B(n39487), .Z(n39480) );
  XOR U58795 ( .A(n39479), .B(n39480), .Z(n39483) );
  XOR U58796 ( .A(n39482), .B(n39483), .Z(n43167) );
  XOR U58797 ( .A(n43165), .B(n43167), .Z(n43170) );
  XOR U58798 ( .A(n43168), .B(n43170), .Z(n39478) );
  XOR U58799 ( .A(n39476), .B(n39478), .Z(n39470) );
  XOR U58800 ( .A(n39469), .B(n39470), .Z(n39474) );
  XOR U58801 ( .A(n39472), .B(n39474), .Z(n39465) );
  XOR U58802 ( .A(n39463), .B(n39465), .Z(n39468) );
  XOR U58803 ( .A(n39466), .B(n39468), .Z(n39461) );
  XOR U58804 ( .A(n39460), .B(n39461), .Z(n39455) );
  XOR U58805 ( .A(n39454), .B(n39455), .Z(n39459) );
  XOR U58806 ( .A(n39457), .B(n39459), .Z(n39450) );
  XOR U58807 ( .A(n39448), .B(n39450), .Z(n39452) );
  XOR U58808 ( .A(n39451), .B(n39452), .Z(n39447) );
  XOR U58809 ( .A(n39445), .B(n39447), .Z(n39441) );
  XOR U58810 ( .A(n39439), .B(n39441), .Z(n39444) );
  XOR U58811 ( .A(n39442), .B(n39444), .Z(n39434) );
  XOR U58812 ( .A(n39433), .B(n39434), .Z(n39438) );
  XOR U58813 ( .A(n39436), .B(n39438), .Z(n39428) );
  XOR U58814 ( .A(n39427), .B(n39428), .Z(n39432) );
  XOR U58815 ( .A(n39430), .B(n39432), .Z(n43176) );
  XOR U58816 ( .A(n43175), .B(n43176), .Z(n43180) );
  XOR U58817 ( .A(n43178), .B(n43180), .Z(n39426) );
  XOR U58818 ( .A(n39424), .B(n39426), .Z(n43186) );
  XOR U58819 ( .A(n43185), .B(n43186), .Z(n39421) );
  XOR U58820 ( .A(n39420), .B(n39421), .Z(n43184) );
  XOR U58821 ( .A(n43182), .B(n43184), .Z(n39416) );
  XOR U58822 ( .A(n39414), .B(n39416), .Z(n39419) );
  XOR U58823 ( .A(n39417), .B(n39419), .Z(n43195) );
  XOR U58824 ( .A(n43194), .B(n43195), .Z(n43199) );
  XOR U58825 ( .A(n43197), .B(n43199), .Z(n39409) );
  XOR U58826 ( .A(n39408), .B(n39409), .Z(n39413) );
  XOR U58827 ( .A(n39411), .B(n39413), .Z(n39403) );
  XOR U58828 ( .A(n39402), .B(n39403), .Z(n39407) );
  XOR U58829 ( .A(n39405), .B(n39407), .Z(n43202) );
  XOR U58830 ( .A(n43201), .B(n43202), .Z(n43205) );
  XOR U58831 ( .A(n43204), .B(n43205), .Z(n39398) );
  XOR U58832 ( .A(n39396), .B(n39398), .Z(n39401) );
  XOR U58833 ( .A(n39399), .B(n39401), .Z(n39391) );
  XOR U58834 ( .A(n39390), .B(n39391), .Z(n39395) );
  XOR U58835 ( .A(n39393), .B(n39395), .Z(n39385) );
  XOR U58836 ( .A(n39384), .B(n39385), .Z(n39389) );
  XOR U58837 ( .A(n39387), .B(n39389), .Z(n39380) );
  XOR U58838 ( .A(n39378), .B(n39380), .Z(n39383) );
  XOR U58839 ( .A(n39381), .B(n39383), .Z(n43210) );
  XOR U58840 ( .A(n43209), .B(n43210), .Z(n43214) );
  XOR U58841 ( .A(n43212), .B(n43214), .Z(n39374) );
  XOR U58842 ( .A(n39372), .B(n39374), .Z(n39377) );
  XOR U58843 ( .A(n39375), .B(n39377), .Z(n43217) );
  XOR U58844 ( .A(n43216), .B(n43217), .Z(n43221) );
  XOR U58845 ( .A(n43219), .B(n43221), .Z(n39367) );
  XOR U58846 ( .A(n39366), .B(n39367), .Z(n39371) );
  XOR U58847 ( .A(n39369), .B(n39371), .Z(n43224) );
  XOR U58848 ( .A(n43222), .B(n43224), .Z(n43227) );
  XOR U58849 ( .A(n43225), .B(n43227), .Z(n39360) );
  XOR U58850 ( .A(n39359), .B(n39360), .Z(n39363) );
  XOR U58851 ( .A(n39362), .B(n39363), .Z(n44955) );
  IV U58852 ( .A(n44955), .Z(n43230) );
  XOR U58853 ( .A(x[1059]), .B(y[1059]), .Z(n44956) );
  IV U58854 ( .A(n44956), .Z(n43229) );
  XOR U58855 ( .A(x[1060]), .B(y[1060]), .Z(n43231) );
  XOR U58856 ( .A(n43229), .B(n43231), .Z(n38635) );
  XOR U58857 ( .A(n43230), .B(n38635), .Z(n39357) );
  XOR U58858 ( .A(n39356), .B(n39357), .Z(n43237) );
  XOR U58859 ( .A(n43235), .B(n43237), .Z(n43240) );
  XOR U58860 ( .A(n43238), .B(n43240), .Z(n39352) );
  XOR U58861 ( .A(n39350), .B(n39352), .Z(n39355) );
  XOR U58862 ( .A(n39353), .B(n39355), .Z(n39346) );
  XOR U58863 ( .A(n39344), .B(n39346), .Z(n39348) );
  XOR U58864 ( .A(n39347), .B(n39348), .Z(n43244) );
  XOR U58865 ( .A(n43243), .B(n43244), .Z(n43248) );
  XOR U58866 ( .A(n43246), .B(n43248), .Z(n43254) );
  XOR U58867 ( .A(n43253), .B(n43254), .Z(n39341) );
  XOR U58868 ( .A(n39340), .B(n39341), .Z(n43252) );
  XOR U58869 ( .A(n43250), .B(n43252), .Z(n39336) );
  XOR U58870 ( .A(n39334), .B(n39336), .Z(n39339) );
  XOR U58871 ( .A(n39337), .B(n39339), .Z(n43262) );
  XOR U58872 ( .A(n43263), .B(n43262), .Z(n43264) );
  XOR U58873 ( .A(n43265), .B(n43264), .Z(n39333) );
  XOR U58874 ( .A(n39331), .B(n39333), .Z(n39327) );
  XOR U58875 ( .A(n39325), .B(n39327), .Z(n39329) );
  XOR U58876 ( .A(n39328), .B(n39329), .Z(n43270) );
  XOR U58877 ( .A(n43269), .B(n43270), .Z(n43274) );
  XOR U58878 ( .A(n43272), .B(n43274), .Z(n39320) );
  XOR U58879 ( .A(n39319), .B(n39320), .Z(n39323) );
  XOR U58880 ( .A(n39322), .B(n39323), .Z(n39317) );
  XOR U58881 ( .A(n39315), .B(n39317), .Z(n43278) );
  XOR U58882 ( .A(n43277), .B(n43278), .Z(n43282) );
  XOR U58883 ( .A(n43280), .B(n43282), .Z(n43284) );
  XOR U58884 ( .A(n43285), .B(n43284), .Z(n43286) );
  XOR U58885 ( .A(n43287), .B(n43286), .Z(n43291) );
  XOR U58886 ( .A(n43289), .B(n43291), .Z(n43294) );
  XOR U58887 ( .A(n43292), .B(n43294), .Z(n43298) );
  XOR U58888 ( .A(n43296), .B(n43298), .Z(n43301) );
  XOR U58889 ( .A(n43299), .B(n43301), .Z(n43304) );
  XOR U58890 ( .A(n43303), .B(n43304), .Z(n43308) );
  XOR U58891 ( .A(n43306), .B(n43308), .Z(n43312) );
  XOR U58892 ( .A(n43310), .B(n43312), .Z(n43315) );
  XOR U58893 ( .A(n43313), .B(n43315), .Z(n44902) );
  XOR U58894 ( .A(x[1097]), .B(y[1097]), .Z(n44903) );
  IV U58895 ( .A(n44903), .Z(n43316) );
  IV U58896 ( .A(x[1098]), .Z(n38636) );
  XOR U58897 ( .A(n38636), .B(y[1098]), .Z(n44905) );
  XOR U58898 ( .A(n43316), .B(n44905), .Z(n38637) );
  XOR U58899 ( .A(n44902), .B(n38637), .Z(n39313) );
  XOR U58900 ( .A(n39312), .B(n39313), .Z(n43325) );
  XOR U58901 ( .A(n43323), .B(n43325), .Z(n39311) );
  XOR U58902 ( .A(n39309), .B(n39311), .Z(n43331) );
  XOR U58903 ( .A(n43329), .B(n43331), .Z(n43333) );
  XOR U58904 ( .A(n43332), .B(n43333), .Z(n43337) );
  XOR U58905 ( .A(n43336), .B(n43337), .Z(n43340) );
  XOR U58906 ( .A(n43339), .B(n43340), .Z(n43345) );
  XOR U58907 ( .A(n43343), .B(n43345), .Z(n43347) );
  XOR U58908 ( .A(n43346), .B(n43347), .Z(n43352) );
  XOR U58909 ( .A(n43350), .B(n43352), .Z(n43355) );
  XOR U58910 ( .A(n43353), .B(n43355), .Z(n43358) );
  XOR U58911 ( .A(n43357), .B(n43358), .Z(n43361) );
  XOR U58912 ( .A(n43360), .B(n43361), .Z(n39307) );
  XOR U58913 ( .A(n39306), .B(n39307), .Z(n43383) );
  XOR U58914 ( .A(n43381), .B(n43383), .Z(n39305) );
  XOR U58915 ( .A(n39303), .B(n39305), .Z(n39298) );
  XOR U58916 ( .A(n39297), .B(n39298), .Z(n39302) );
  XOR U58917 ( .A(n39300), .B(n39302), .Z(n39293) );
  XOR U58918 ( .A(n39291), .B(n39293), .Z(n39295) );
  XOR U58919 ( .A(n39294), .B(n39295), .Z(n39288) );
  XOR U58920 ( .A(n39287), .B(n39288), .Z(n43394) );
  XOR U58921 ( .A(n43392), .B(n43394), .Z(n43397) );
  XOR U58922 ( .A(n43395), .B(n43397), .Z(n39285) );
  XOR U58923 ( .A(n39284), .B(n39285), .Z(n43403) );
  XOR U58924 ( .A(n43401), .B(n43403), .Z(n39283) );
  XOR U58925 ( .A(n39281), .B(n39283), .Z(n43411) );
  XOR U58926 ( .A(n43409), .B(n43411), .Z(n43413) );
  XOR U58927 ( .A(n43412), .B(n43413), .Z(n39278) );
  XOR U58928 ( .A(n39280), .B(n39278), .Z(n43417) );
  XOR U58929 ( .A(n43415), .B(n43417), .Z(n43420) );
  XOR U58930 ( .A(n43418), .B(n43420), .Z(n39273) );
  XOR U58931 ( .A(n39272), .B(n39273), .Z(n39276) );
  XOR U58932 ( .A(n39275), .B(n39276), .Z(n39267) );
  XOR U58933 ( .A(n39265), .B(n39267), .Z(n39269) );
  XOR U58934 ( .A(n39268), .B(n39269), .Z(n43424) );
  XOR U58935 ( .A(n43422), .B(n43424), .Z(n43426) );
  XOR U58936 ( .A(n43425), .B(n43426), .Z(n43430) );
  XOR U58937 ( .A(n43429), .B(n43430), .Z(n43434) );
  XOR U58938 ( .A(n43432), .B(n43434), .Z(n39264) );
  XOR U58939 ( .A(n39262), .B(n39264), .Z(n39257) );
  XOR U58940 ( .A(n39258), .B(n39257), .Z(n39259) );
  XOR U58941 ( .A(n39260), .B(n39259), .Z(n39253) );
  XOR U58942 ( .A(n39251), .B(n39253), .Z(n39255) );
  XOR U58943 ( .A(n39254), .B(n39255), .Z(n43439) );
  XOR U58944 ( .A(n43438), .B(n43439), .Z(n43442) );
  XOR U58945 ( .A(n43441), .B(n43442), .Z(n39250) );
  XOR U58946 ( .A(n39248), .B(n39250), .Z(n39244) );
  XOR U58947 ( .A(n39242), .B(n39244), .Z(n39246) );
  XOR U58948 ( .A(n39245), .B(n39246), .Z(n43453) );
  XOR U58949 ( .A(n43451), .B(n43453), .Z(n43455) );
  XOR U58950 ( .A(n43454), .B(n43455), .Z(n39241) );
  XOR U58951 ( .A(n39239), .B(n39241), .Z(n43459) );
  XOR U58952 ( .A(n43460), .B(n43459), .Z(n39236) );
  XOR U58953 ( .A(n39238), .B(n39236), .Z(n43468) );
  XOR U58954 ( .A(n43466), .B(n43468), .Z(n43470) );
  XOR U58955 ( .A(n43469), .B(n43470), .Z(n39231) );
  XOR U58956 ( .A(n39230), .B(n39231), .Z(n39235) );
  XOR U58957 ( .A(n39233), .B(n39235), .Z(n43473) );
  XOR U58958 ( .A(n43472), .B(n43473), .Z(n43477) );
  XOR U58959 ( .A(n43475), .B(n43477), .Z(n39229) );
  XOR U58960 ( .A(n39227), .B(n39229), .Z(n43482) );
  XOR U58961 ( .A(n43480), .B(n43482), .Z(n39225) );
  XOR U58962 ( .A(n39224), .B(n39225), .Z(n43487) );
  XOR U58963 ( .A(n43486), .B(n43487), .Z(n43490) );
  XOR U58964 ( .A(n43489), .B(n43490), .Z(n43495) );
  XOR U58965 ( .A(n43497), .B(n43495), .Z(n43499) );
  XOR U58966 ( .A(n43498), .B(n43499), .Z(n43493) );
  XOR U58967 ( .A(n43492), .B(n43493), .Z(n43509) );
  XOR U58968 ( .A(n43507), .B(n43509), .Z(n43512) );
  XOR U58969 ( .A(n43510), .B(n43512), .Z(n43515) );
  XOR U58970 ( .A(n43514), .B(n43515), .Z(n43519) );
  XOR U58971 ( .A(n43517), .B(n43519), .Z(n39220) );
  XOR U58972 ( .A(n39218), .B(n39220), .Z(n39223) );
  XOR U58973 ( .A(n39221), .B(n39223), .Z(n43522) );
  XOR U58974 ( .A(n43520), .B(n43522), .Z(n43524) );
  XOR U58975 ( .A(n43523), .B(n43524), .Z(n39216) );
  XOR U58976 ( .A(n39217), .B(n39216), .Z(n39210) );
  XOR U58977 ( .A(n39211), .B(n39210), .Z(n39214) );
  XOR U58978 ( .A(n39213), .B(n39214), .Z(n39206) );
  XOR U58979 ( .A(n39204), .B(n39206), .Z(n39208) );
  XOR U58980 ( .A(n39207), .B(n39208), .Z(n39203) );
  XOR U58981 ( .A(n39201), .B(n39203), .Z(n39197) );
  XOR U58982 ( .A(n39195), .B(n39197), .Z(n39199) );
  XOR U58983 ( .A(n39198), .B(n39199), .Z(n39190) );
  XOR U58984 ( .A(n39189), .B(n39190), .Z(n39194) );
  XOR U58985 ( .A(n39192), .B(n39194), .Z(n64082) );
  IV U58986 ( .A(n64082), .Z(n39185) );
  XOR U58987 ( .A(x[1185]), .B(y[1185]), .Z(n64081) );
  XOR U58988 ( .A(x[1186]), .B(y[1186]), .Z(n39186) );
  XOR U58989 ( .A(n64081), .B(n39186), .Z(n38638) );
  XOR U58990 ( .A(n39185), .B(n38638), .Z(n43530) );
  XOR U58991 ( .A(x[1187]), .B(y[1187]), .Z(n53577) );
  IV U58992 ( .A(x[1188]), .Z(n38639) );
  XOR U58993 ( .A(n38639), .B(y[1188]), .Z(n53580) );
  XOR U58994 ( .A(n53577), .B(n53580), .Z(n38640) );
  XOR U58995 ( .A(n43530), .B(n38640), .Z(n39179) );
  XOR U58996 ( .A(n39178), .B(n39179), .Z(n39183) );
  XOR U58997 ( .A(n39181), .B(n39183), .Z(n43536) );
  XOR U58998 ( .A(n43534), .B(n43536), .Z(n43538) );
  XOR U58999 ( .A(n43537), .B(n43538), .Z(n43543) );
  XOR U59000 ( .A(n43541), .B(n43543), .Z(n43546) );
  XOR U59001 ( .A(n43544), .B(n43546), .Z(n43549) );
  XOR U59002 ( .A(n43548), .B(n43549), .Z(n43552) );
  XOR U59003 ( .A(n43551), .B(n43552), .Z(n43557) );
  XOR U59004 ( .A(n43555), .B(n43557), .Z(n43560) );
  XOR U59005 ( .A(n43558), .B(n43560), .Z(n39176) );
  XOR U59006 ( .A(n39175), .B(n39176), .Z(n43564) );
  XOR U59007 ( .A(n43563), .B(n43564), .Z(n43568) );
  XOR U59008 ( .A(n43566), .B(n43568), .Z(n43572) );
  XOR U59009 ( .A(n43570), .B(n43572), .Z(n43574) );
  XOR U59010 ( .A(n43573), .B(n43574), .Z(n43578) );
  XOR U59011 ( .A(n43577), .B(n43578), .Z(n43581) );
  XOR U59012 ( .A(n43580), .B(n43581), .Z(n39172) );
  XOR U59013 ( .A(n39174), .B(n39172), .Z(n43586) );
  XOR U59014 ( .A(n43585), .B(n43586), .Z(n39171) );
  XOR U59015 ( .A(n39169), .B(n39171), .Z(n43595) );
  XOR U59016 ( .A(n43593), .B(n43595), .Z(n39168) );
  XOR U59017 ( .A(n39166), .B(n39168), .Z(n43605) );
  XOR U59018 ( .A(n43604), .B(n43605), .Z(n43609) );
  XOR U59019 ( .A(n43607), .B(n43609), .Z(n43612) );
  XOR U59020 ( .A(n43611), .B(n43612), .Z(n43616) );
  XOR U59021 ( .A(n43614), .B(n43616), .Z(n39164) );
  XOR U59022 ( .A(n39163), .B(n39164), .Z(n43620) );
  XOR U59023 ( .A(n43619), .B(n43620), .Z(n43623) );
  XOR U59024 ( .A(n43622), .B(n43623), .Z(n39160) );
  XOR U59025 ( .A(n39162), .B(n39160), .Z(n43629) );
  XOR U59026 ( .A(n43627), .B(n43629), .Z(n39159) );
  XOR U59027 ( .A(n39157), .B(n39159), .Z(n43636) );
  XOR U59028 ( .A(n43635), .B(n43636), .Z(n43640) );
  XOR U59029 ( .A(n43638), .B(n43640), .Z(n39153) );
  XOR U59030 ( .A(n39151), .B(n39153), .Z(n39156) );
  XOR U59031 ( .A(n39154), .B(n39156), .Z(n43646) );
  XOR U59032 ( .A(n43645), .B(n43646), .Z(n39149) );
  XOR U59033 ( .A(n39148), .B(n39149), .Z(n43657) );
  XOR U59034 ( .A(n43655), .B(n43657), .Z(n43660) );
  XOR U59035 ( .A(n43658), .B(n43660), .Z(n43663) );
  XOR U59036 ( .A(n43662), .B(n43663), .Z(n43664) );
  XOR U59037 ( .A(n43665), .B(n43664), .Z(n43668) );
  XOR U59038 ( .A(n43667), .B(n43668), .Z(n43671) );
  XOR U59039 ( .A(n43670), .B(n43671), .Z(n39144) );
  XOR U59040 ( .A(n39142), .B(n39144), .Z(n39147) );
  XOR U59041 ( .A(n39145), .B(n39147), .Z(n43675) );
  XOR U59042 ( .A(n43674), .B(n43675), .Z(n43679) );
  XOR U59043 ( .A(n43677), .B(n43679), .Z(n39137) );
  XOR U59044 ( .A(n39135), .B(n39137), .Z(n39140) );
  XOR U59045 ( .A(n39138), .B(n39140), .Z(n43682) );
  XOR U59046 ( .A(n43681), .B(n43682), .Z(n43685) );
  XOR U59047 ( .A(n43684), .B(n43685), .Z(n43689) );
  XOR U59048 ( .A(n43688), .B(n43689), .Z(n43690) );
  XOR U59049 ( .A(n43691), .B(n43690), .Z(n43694) );
  XOR U59050 ( .A(n43693), .B(n43694), .Z(n43698) );
  XOR U59051 ( .A(n43696), .B(n43698), .Z(n39131) );
  XOR U59052 ( .A(n39129), .B(n39131), .Z(n39134) );
  XOR U59053 ( .A(n39132), .B(n39134), .Z(n39127) );
  XOR U59054 ( .A(n39126), .B(n39127), .Z(n43700) );
  XOR U59055 ( .A(n43699), .B(n43700), .Z(n43704) );
  XOR U59056 ( .A(n43702), .B(n43704), .Z(n39124) );
  XOR U59057 ( .A(n39123), .B(n39124), .Z(n39116) );
  IV U59058 ( .A(n39116), .Z(n39118) );
  XOR U59059 ( .A(n39117), .B(n39118), .Z(n49652) );
  XOR U59060 ( .A(n39120), .B(n49652), .Z(n43708) );
  XOR U59061 ( .A(n43706), .B(n43708), .Z(n43710) );
  XOR U59062 ( .A(n43709), .B(n43710), .Z(n39114) );
  XOR U59063 ( .A(n39113), .B(n39114), .Z(n43715) );
  XOR U59064 ( .A(n43714), .B(n43715), .Z(n43719) );
  XOR U59065 ( .A(n43717), .B(n43719), .Z(n39108) );
  XOR U59066 ( .A(n39107), .B(n39108), .Z(n39111) );
  XOR U59067 ( .A(n39110), .B(n39111), .Z(n39103) );
  XOR U59068 ( .A(n39101), .B(n39103), .Z(n39106) );
  XOR U59069 ( .A(n39104), .B(n39106), .Z(n43724) );
  XOR U59070 ( .A(n43722), .B(n43724), .Z(n43726) );
  XOR U59071 ( .A(n43725), .B(n43726), .Z(n39096) );
  XOR U59072 ( .A(n39095), .B(n39096), .Z(n39100) );
  XOR U59073 ( .A(n39098), .B(n39100), .Z(n39091) );
  XOR U59074 ( .A(n39089), .B(n39091), .Z(n39093) );
  XOR U59075 ( .A(n39092), .B(n39093), .Z(n39087) );
  XOR U59076 ( .A(n39086), .B(n39087), .Z(n39082) );
  XOR U59077 ( .A(n39080), .B(n39082), .Z(n39084) );
  XOR U59078 ( .A(n39083), .B(n39084), .Z(n39075) );
  XOR U59079 ( .A(n39074), .B(n39075), .Z(n39079) );
  XOR U59080 ( .A(n39077), .B(n39079), .Z(n39070) );
  XOR U59081 ( .A(n39068), .B(n39070), .Z(n39073) );
  XOR U59082 ( .A(n39071), .B(n39073), .Z(n43732) );
  XOR U59083 ( .A(n43731), .B(n43732), .Z(n43736) );
  XOR U59084 ( .A(n43734), .B(n43736), .Z(n43740) );
  XOR U59085 ( .A(n43738), .B(n43740), .Z(n43743) );
  XOR U59086 ( .A(n43741), .B(n43743), .Z(n43746) );
  XOR U59087 ( .A(n43745), .B(n43746), .Z(n43749) );
  XOR U59088 ( .A(n43748), .B(n43749), .Z(n43756) );
  XOR U59089 ( .A(n43754), .B(n43756), .Z(n39066) );
  XOR U59090 ( .A(n39065), .B(n39066), .Z(n44683) );
  XOR U59091 ( .A(x[1283]), .B(y[1283]), .Z(n44684) );
  IV U59092 ( .A(n44684), .Z(n39061) );
  IV U59093 ( .A(x[1284]), .Z(n38641) );
  XOR U59094 ( .A(n38641), .B(y[1284]), .Z(n44686) );
  XOR U59095 ( .A(n39061), .B(n44686), .Z(n38642) );
  XOR U59096 ( .A(n44683), .B(n38642), .Z(n39056) );
  XOR U59097 ( .A(n39054), .B(n39056), .Z(n39059) );
  XOR U59098 ( .A(n39057), .B(n39059), .Z(n39049) );
  XOR U59099 ( .A(n39048), .B(n39049), .Z(n39053) );
  XOR U59100 ( .A(n39051), .B(n39053), .Z(n43769) );
  XOR U59101 ( .A(n43767), .B(n43769), .Z(n43772) );
  XOR U59102 ( .A(n43770), .B(n43772), .Z(n39047) );
  XOR U59103 ( .A(n39045), .B(n39047), .Z(n39041) );
  XOR U59104 ( .A(n39039), .B(n39041), .Z(n39044) );
  XOR U59105 ( .A(n39042), .B(n39044), .Z(n39034) );
  XOR U59106 ( .A(n39033), .B(n39034), .Z(n39037) );
  XOR U59107 ( .A(n39036), .B(n39037), .Z(n39032) );
  XOR U59108 ( .A(n39030), .B(n39032), .Z(n39027) );
  XOR U59109 ( .A(n39025), .B(n39027), .Z(n39028) );
  XOR U59110 ( .A(n39029), .B(n39028), .Z(n39018) );
  XOR U59111 ( .A(n39020), .B(n39018), .Z(n39023) );
  XOR U59112 ( .A(n39021), .B(n39023), .Z(n39013) );
  XOR U59113 ( .A(n39012), .B(n39013), .Z(n39016) );
  XOR U59114 ( .A(n39015), .B(n39016), .Z(n39007) );
  XOR U59115 ( .A(n39006), .B(n39007), .Z(n39010) );
  XOR U59116 ( .A(n39009), .B(n39010), .Z(n39002) );
  XOR U59117 ( .A(n39000), .B(n39002), .Z(n39005) );
  XOR U59118 ( .A(n39003), .B(n39005), .Z(n38998) );
  XOR U59119 ( .A(n38997), .B(n38998), .Z(n43777) );
  IV U59120 ( .A(n43777), .Z(n43779) );
  XOR U59121 ( .A(n43776), .B(n43779), .Z(n48591) );
  XOR U59122 ( .A(n43780), .B(n48591), .Z(n43785) );
  XOR U59123 ( .A(n43784), .B(n43785), .Z(n43788) );
  XOR U59124 ( .A(n43787), .B(n43788), .Z(n38996) );
  XOR U59125 ( .A(n38994), .B(n38996), .Z(n48600) );
  XOR U59126 ( .A(n48598), .B(n48600), .Z(n44667) );
  XOR U59127 ( .A(n44665), .B(n44667), .Z(n38993) );
  XOR U59128 ( .A(n38991), .B(n38993), .Z(n43797) );
  XOR U59129 ( .A(n43795), .B(n43797), .Z(n43800) );
  XOR U59130 ( .A(n43798), .B(n43800), .Z(n43803) );
  XOR U59131 ( .A(n43802), .B(n43803), .Z(n43806) );
  XOR U59132 ( .A(n43805), .B(n43806), .Z(n43810) );
  XOR U59133 ( .A(n43808), .B(n43810), .Z(n43812) );
  XOR U59134 ( .A(n43811), .B(n43812), .Z(n38986) );
  XOR U59135 ( .A(n38985), .B(n38986), .Z(n38989) );
  XOR U59136 ( .A(n38988), .B(n38989), .Z(n43816) );
  XOR U59137 ( .A(n43815), .B(n43816), .Z(n43819) );
  XOR U59138 ( .A(n43818), .B(n43819), .Z(n38981) );
  XOR U59139 ( .A(n38979), .B(n38981), .Z(n38983) );
  XOR U59140 ( .A(n38982), .B(n38983), .Z(n38977) );
  XOR U59141 ( .A(n38976), .B(n38977), .Z(n43825) );
  XOR U59142 ( .A(n43823), .B(n43825), .Z(n43827) );
  XOR U59143 ( .A(n43826), .B(n43827), .Z(n43833) );
  XOR U59144 ( .A(n43831), .B(n43833), .Z(n43836) );
  XOR U59145 ( .A(n43834), .B(n43836), .Z(n38975) );
  XOR U59146 ( .A(n38973), .B(n38975), .Z(n43844) );
  XOR U59147 ( .A(n43842), .B(n43844), .Z(n43846) );
  XOR U59148 ( .A(n43845), .B(n43846), .Z(n43851) );
  XOR U59149 ( .A(n43849), .B(n43851), .Z(n43854) );
  XOR U59150 ( .A(n43852), .B(n43854), .Z(n38972) );
  XOR U59151 ( .A(n38970), .B(n38972), .Z(n38965) );
  XOR U59152 ( .A(n38964), .B(n38965), .Z(n38969) );
  XOR U59153 ( .A(n38967), .B(n38969), .Z(n38959) );
  XOR U59154 ( .A(n38958), .B(n38959), .Z(n38963) );
  XOR U59155 ( .A(n38961), .B(n38963), .Z(n38953) );
  XOR U59156 ( .A(n38952), .B(n38953), .Z(n38957) );
  XOR U59157 ( .A(n38955), .B(n38957), .Z(n38948) );
  XOR U59158 ( .A(n38946), .B(n38948), .Z(n38950) );
  XOR U59159 ( .A(n38949), .B(n38950), .Z(n44631) );
  IV U59160 ( .A(n44631), .Z(n43860) );
  XOR U59161 ( .A(x[1347]), .B(y[1347]), .Z(n44630) );
  IV U59162 ( .A(x[1348]), .Z(n38643) );
  XOR U59163 ( .A(n38643), .B(y[1348]), .Z(n44633) );
  XOR U59164 ( .A(n44630), .B(n44633), .Z(n38644) );
  XOR U59165 ( .A(n43860), .B(n38644), .Z(n43865) );
  XOR U59166 ( .A(n43864), .B(n43865), .Z(n43869) );
  XOR U59167 ( .A(n43867), .B(n43869), .Z(n43873) );
  XOR U59168 ( .A(n43871), .B(n43873), .Z(n43876) );
  XOR U59169 ( .A(n43874), .B(n43876), .Z(n43879) );
  XOR U59170 ( .A(n43878), .B(n43879), .Z(n43882) );
  XOR U59171 ( .A(n43881), .B(n43882), .Z(n43886) );
  XOR U59172 ( .A(n43885), .B(n43886), .Z(n43890) );
  XOR U59173 ( .A(n43888), .B(n43890), .Z(n38942) );
  XOR U59174 ( .A(n38940), .B(n38942), .Z(n38945) );
  XOR U59175 ( .A(n38943), .B(n38945), .Z(n43893) );
  XOR U59176 ( .A(n43892), .B(n43893), .Z(n43896) );
  XOR U59177 ( .A(n43895), .B(n43896), .Z(n38936) );
  XOR U59178 ( .A(n38934), .B(n38936), .Z(n38939) );
  XOR U59179 ( .A(n38937), .B(n38939), .Z(n38929) );
  XOR U59180 ( .A(n38928), .B(n38929), .Z(n38933) );
  XOR U59181 ( .A(n38931), .B(n38933), .Z(n43907) );
  XOR U59182 ( .A(n43905), .B(n43907), .Z(n38927) );
  XOR U59183 ( .A(n38925), .B(n38927), .Z(n43903) );
  XOR U59184 ( .A(n43904), .B(n43903), .Z(n38919) );
  XOR U59185 ( .A(n38921), .B(n38919), .Z(n38924) );
  XOR U59186 ( .A(n38922), .B(n38924), .Z(n38918) );
  XOR U59187 ( .A(n38916), .B(n38918), .Z(n43919) );
  XOR U59188 ( .A(n43918), .B(n43919), .Z(n43923) );
  XOR U59189 ( .A(n43921), .B(n43923), .Z(n43928) );
  XOR U59190 ( .A(n43926), .B(n43928), .Z(n43930) );
  XOR U59191 ( .A(n43929), .B(n43930), .Z(n43934) );
  XOR U59192 ( .A(n43933), .B(n43934), .Z(n43937) );
  XOR U59193 ( .A(n43936), .B(n43937), .Z(n38911) );
  XOR U59194 ( .A(n38912), .B(n38911), .Z(n48766) );
  XOR U59195 ( .A(n48765), .B(n48766), .Z(n38904) );
  XOR U59196 ( .A(n38906), .B(n38904), .Z(n59206) );
  XOR U59197 ( .A(n59205), .B(n59206), .Z(n38898) );
  XOR U59198 ( .A(n38897), .B(n38898), .Z(n38902) );
  XOR U59199 ( .A(n38900), .B(n38902), .Z(n43943) );
  XOR U59200 ( .A(n43941), .B(n43943), .Z(n43945) );
  XOR U59201 ( .A(n43944), .B(n43945), .Z(n43950) );
  XOR U59202 ( .A(n43949), .B(n43950), .Z(n48790) );
  XOR U59203 ( .A(n48789), .B(n48790), .Z(n43956) );
  XOR U59204 ( .A(n43955), .B(n43956), .Z(n43959) );
  XOR U59205 ( .A(n43958), .B(n43959), .Z(n38895) );
  XOR U59206 ( .A(n38893), .B(n38895), .Z(n43963) );
  XOR U59207 ( .A(n43961), .B(n43963), .Z(n43965) );
  XOR U59208 ( .A(n43964), .B(n43965), .Z(n43969) );
  XOR U59209 ( .A(n43968), .B(n43969), .Z(n43973) );
  XOR U59210 ( .A(n43971), .B(n43973), .Z(n43976) );
  XOR U59211 ( .A(n43974), .B(n43976), .Z(n43978) );
  XOR U59212 ( .A(n43977), .B(n43978), .Z(n43983) );
  XOR U59213 ( .A(n43981), .B(n43983), .Z(n43986) );
  XOR U59214 ( .A(n43984), .B(n43986), .Z(n43989) );
  XOR U59215 ( .A(n43988), .B(n43989), .Z(n43992) );
  XOR U59216 ( .A(n43991), .B(n43992), .Z(n43998) );
  XOR U59217 ( .A(n43997), .B(n43998), .Z(n38892) );
  XOR U59218 ( .A(n38890), .B(n38892), .Z(n44009) );
  XOR U59219 ( .A(n44008), .B(n44009), .Z(n44012) );
  XOR U59220 ( .A(n44011), .B(n44012), .Z(n44017) );
  XOR U59221 ( .A(n44015), .B(n44017), .Z(n44020) );
  XOR U59222 ( .A(n44018), .B(n44020), .Z(n44023) );
  XOR U59223 ( .A(n44021), .B(n44023), .Z(n44025) );
  XOR U59224 ( .A(n44024), .B(n44025), .Z(n38886) );
  XOR U59225 ( .A(n38884), .B(n38886), .Z(n38889) );
  XOR U59226 ( .A(n38887), .B(n38889), .Z(n38882) );
  XOR U59227 ( .A(n38881), .B(n38882), .Z(n48815) );
  IV U59228 ( .A(n48815), .Z(n44028) );
  XOR U59229 ( .A(n48814), .B(n44028), .Z(n48828) );
  XOR U59230 ( .A(n48827), .B(n48828), .Z(n44034) );
  XOR U59231 ( .A(n44032), .B(n44034), .Z(n44037) );
  XOR U59232 ( .A(n44035), .B(n44037), .Z(n38877) );
  XOR U59233 ( .A(n38875), .B(n38877), .Z(n38880) );
  XOR U59234 ( .A(n38878), .B(n38880), .Z(n44042) );
  XOR U59235 ( .A(n44041), .B(n44042), .Z(n48839) );
  XOR U59236 ( .A(n48838), .B(n48839), .Z(n44049) );
  XOR U59237 ( .A(n44047), .B(n44049), .Z(n44051) );
  XOR U59238 ( .A(n44050), .B(n44051), .Z(n38874) );
  XOR U59239 ( .A(n38872), .B(n38874), .Z(n44059) );
  XOR U59240 ( .A(n44057), .B(n44059), .Z(n38870) );
  XOR U59241 ( .A(n38869), .B(n38870), .Z(n38865) );
  XOR U59242 ( .A(n38863), .B(n38865), .Z(n38868) );
  XOR U59243 ( .A(n38866), .B(n38868), .Z(n38859) );
  XOR U59244 ( .A(n38857), .B(n38859), .Z(n38861) );
  XOR U59245 ( .A(n38860), .B(n38861), .Z(n38853) );
  XOR U59246 ( .A(n38851), .B(n38853), .Z(n38856) );
  XOR U59247 ( .A(n38854), .B(n38856), .Z(n44066) );
  XOR U59248 ( .A(n44065), .B(n44066), .Z(n44069) );
  XOR U59249 ( .A(n44068), .B(n44069), .Z(n38849) );
  XOR U59250 ( .A(n38848), .B(n38849), .Z(n38844) );
  XOR U59251 ( .A(n38842), .B(n38844), .Z(n38847) );
  XOR U59252 ( .A(n38845), .B(n38847), .Z(n38836) );
  XOR U59253 ( .A(n38838), .B(n38836), .Z(n64516) );
  XOR U59254 ( .A(n38839), .B(n64516), .Z(n38834) );
  XOR U59255 ( .A(n38832), .B(n38834), .Z(n38828) );
  XOR U59256 ( .A(n38826), .B(n38828), .Z(n38831) );
  XOR U59257 ( .A(n38829), .B(n38831), .Z(n38821) );
  XOR U59258 ( .A(n38820), .B(n38821), .Z(n38824) );
  XOR U59259 ( .A(n38823), .B(n38824), .Z(n44079) );
  XOR U59260 ( .A(n44078), .B(n44079), .Z(n38818) );
  XOR U59261 ( .A(n38817), .B(n38818), .Z(n44077) );
  XOR U59262 ( .A(n44075), .B(n44077), .Z(n44088) );
  XOR U59263 ( .A(n44086), .B(n44088), .Z(n44091) );
  XOR U59264 ( .A(n44089), .B(n44091), .Z(n44094) );
  XOR U59265 ( .A(n44093), .B(n44094), .Z(n44097) );
  XOR U59266 ( .A(n44096), .B(n44097), .Z(n38816) );
  XOR U59267 ( .A(n38814), .B(n38816), .Z(n38810) );
  XOR U59268 ( .A(n38808), .B(n38810), .Z(n38812) );
  XOR U59269 ( .A(n38811), .B(n38812), .Z(n44112) );
  XOR U59270 ( .A(n44110), .B(n44112), .Z(n44115) );
  XOR U59271 ( .A(n44113), .B(n44115), .Z(n38804) );
  XOR U59272 ( .A(n38802), .B(n38804), .Z(n38806) );
  XOR U59273 ( .A(n38805), .B(n38806), .Z(n44118) );
  XOR U59274 ( .A(n44117), .B(n44118), .Z(n44122) );
  XOR U59275 ( .A(n44120), .B(n44122), .Z(n38801) );
  XOR U59276 ( .A(n38799), .B(n38801), .Z(n38793) );
  XOR U59277 ( .A(n38792), .B(n38793), .Z(n38797) );
  XOR U59278 ( .A(n38795), .B(n38797), .Z(n44126) );
  XOR U59279 ( .A(n44124), .B(n44126), .Z(n44129) );
  XOR U59280 ( .A(n44127), .B(n44129), .Z(n38788) );
  XOR U59281 ( .A(n38786), .B(n38788), .Z(n38791) );
  XOR U59282 ( .A(n38789), .B(n38791), .Z(n44132) );
  XOR U59283 ( .A(n44130), .B(n44132), .Z(n44135) );
  XOR U59284 ( .A(n44133), .B(n44135), .Z(n38785) );
  XOR U59285 ( .A(n38783), .B(n38785), .Z(n38779) );
  XOR U59286 ( .A(n38777), .B(n38779), .Z(n38782) );
  XOR U59287 ( .A(n38780), .B(n38782), .Z(n38773) );
  XOR U59288 ( .A(n38771), .B(n38773), .Z(n38775) );
  XOR U59289 ( .A(n38774), .B(n38775), .Z(n38770) );
  XOR U59290 ( .A(n38768), .B(n38770), .Z(n44141) );
  XOR U59291 ( .A(n44140), .B(n44141), .Z(n38766) );
  XOR U59292 ( .A(n38765), .B(n38766), .Z(n44148) );
  XOR U59293 ( .A(n44147), .B(n44148), .Z(n44152) );
  XOR U59294 ( .A(n44150), .B(n44152), .Z(n44155) );
  XOR U59295 ( .A(n44154), .B(n44155), .Z(n44159) );
  XOR U59296 ( .A(n44157), .B(n44159), .Z(n38764) );
  XOR U59297 ( .A(n38762), .B(n38764), .Z(n44163) );
  XOR U59298 ( .A(n44161), .B(n44163), .Z(n44165) );
  XOR U59299 ( .A(n44164), .B(n44165), .Z(n38761) );
  XOR U59300 ( .A(n38759), .B(n38761), .Z(n44179) );
  XOR U59301 ( .A(n44178), .B(n44179), .Z(n44183) );
  XOR U59302 ( .A(n44181), .B(n44183), .Z(n44187) );
  XOR U59303 ( .A(n44185), .B(n44187), .Z(n44190) );
  XOR U59304 ( .A(n44188), .B(n44190), .Z(n38757) );
  XOR U59305 ( .A(n38756), .B(n38757), .Z(n44193) );
  XOR U59306 ( .A(n44192), .B(n44193), .Z(n44196) );
  XOR U59307 ( .A(n44195), .B(n44196), .Z(n44201) );
  XOR U59308 ( .A(n44199), .B(n44201), .Z(n44204) );
  XOR U59309 ( .A(n44202), .B(n44204), .Z(n38755) );
  XOR U59310 ( .A(n38753), .B(n38755), .Z(n44207) );
  XOR U59311 ( .A(n44206), .B(n44207), .Z(n44211) );
  XOR U59312 ( .A(n44209), .B(n44211), .Z(n44214) );
  XOR U59313 ( .A(n44213), .B(n44214), .Z(n44217) );
  XOR U59314 ( .A(n44216), .B(n44217), .Z(n44221) );
  XOR U59315 ( .A(n44219), .B(n44221), .Z(n44223) );
  XOR U59316 ( .A(n44222), .B(n44223), .Z(n38748) );
  XOR U59317 ( .A(n38747), .B(n38748), .Z(n38752) );
  XOR U59318 ( .A(n38750), .B(n38752), .Z(n44227) );
  XOR U59319 ( .A(n44225), .B(n44227), .Z(n44230) );
  XOR U59320 ( .A(n44228), .B(n44230), .Z(n38742) );
  XOR U59321 ( .A(n38741), .B(n38742), .Z(n38746) );
  XOR U59322 ( .A(n38744), .B(n38746), .Z(n38739) );
  XOR U59323 ( .A(n38738), .B(n38739), .Z(n44236) );
  XOR U59324 ( .A(n44234), .B(n44236), .Z(n44461) );
  XOR U59325 ( .A(n44459), .B(n44461), .Z(n44244) );
  XOR U59326 ( .A(n44245), .B(n44244), .Z(n38734) );
  XOR U59327 ( .A(n38732), .B(n38734), .Z(n38737) );
  XOR U59328 ( .A(n38735), .B(n38737), .Z(n38730) );
  XOR U59329 ( .A(n38728), .B(n38730), .Z(n44250) );
  XOR U59330 ( .A(n44248), .B(n44250), .Z(n44252) );
  XOR U59331 ( .A(n44251), .B(n44252), .Z(n44264) );
  XOR U59332 ( .A(n44263), .B(n44264), .Z(n44257) );
  XOR U59333 ( .A(n44256), .B(n44257), .Z(n44261) );
  XOR U59334 ( .A(n44260), .B(n44261), .Z(n38727) );
  XOR U59335 ( .A(n38725), .B(n38727), .Z(n44274) );
  XOR U59336 ( .A(n44273), .B(n44274), .Z(n38722) );
  XOR U59337 ( .A(n38724), .B(n38722), .Z(n44281) );
  XOR U59338 ( .A(n44280), .B(n44281), .Z(n44282) );
  XOR U59339 ( .A(n44283), .B(n44282), .Z(n38718) );
  XOR U59340 ( .A(n38716), .B(n38718), .Z(n38720) );
  XOR U59341 ( .A(n38719), .B(n38720), .Z(n38712) );
  XOR U59342 ( .A(n38710), .B(n38712), .Z(n38715) );
  XOR U59343 ( .A(n38713), .B(n38715), .Z(n44288) );
  XOR U59344 ( .A(n44287), .B(n44288), .Z(n44291) );
  XOR U59345 ( .A(n44290), .B(n44291), .Z(n38705) );
  XOR U59346 ( .A(n38704), .B(n38705), .Z(n38709) );
  XOR U59347 ( .A(n38707), .B(n38709), .Z(n38700) );
  XOR U59348 ( .A(n38698), .B(n38700), .Z(n38702) );
  XOR U59349 ( .A(n38701), .B(n38702), .Z(n38693) );
  XOR U59350 ( .A(n38692), .B(n38693), .Z(n38697) );
  XOR U59351 ( .A(n38695), .B(n38697), .Z(n44296) );
  XOR U59352 ( .A(n44294), .B(n44296), .Z(n44298) );
  XOR U59353 ( .A(n44297), .B(n44298), .Z(n44302) );
  XOR U59354 ( .A(n44301), .B(n44302), .Z(n44306) );
  XOR U59355 ( .A(n44304), .B(n44306), .Z(n44309) );
  XOR U59356 ( .A(n44308), .B(n44309), .Z(n44313) );
  XOR U59357 ( .A(n44311), .B(n44313), .Z(n38688) );
  XOR U59358 ( .A(n38687), .B(n38688), .Z(n38689) );
  XOR U59359 ( .A(n38691), .B(n38689), .Z(n44318) );
  XOR U59360 ( .A(n44316), .B(n44318), .Z(n44320) );
  XOR U59361 ( .A(n44319), .B(n44320), .Z(n38685) );
  XOR U59362 ( .A(n38684), .B(n38685), .Z(n38680) );
  XOR U59363 ( .A(n38678), .B(n38680), .Z(n38683) );
  XOR U59364 ( .A(n38681), .B(n38683), .Z(n44327) );
  XOR U59365 ( .A(n44325), .B(n44327), .Z(n44330) );
  XOR U59366 ( .A(n44328), .B(n44330), .Z(n44332) );
  XOR U59367 ( .A(n44333), .B(n44332), .Z(n44334) );
  XOR U59368 ( .A(n44335), .B(n44334), .Z(n38673) );
  XOR U59369 ( .A(n38672), .B(n38673), .Z(n38677) );
  XOR U59370 ( .A(n38675), .B(n38677), .Z(n38667) );
  XOR U59371 ( .A(n38668), .B(n38667), .Z(n38669) );
  XOR U59372 ( .A(n38670), .B(n38669), .Z(n44339) );
  XOR U59373 ( .A(n44338), .B(n44339), .Z(n44343) );
  XOR U59374 ( .A(n44341), .B(n44343), .Z(n38662) );
  XOR U59375 ( .A(n38663), .B(n38662), .Z(n38664) );
  XOR U59376 ( .A(n38665), .B(n38664), .Z(n44348) );
  XOR U59377 ( .A(n44347), .B(n44348), .Z(n44351) );
  XOR U59378 ( .A(n44350), .B(n44351), .Z(n38661) );
  XOR U59379 ( .A(n38660), .B(n38661), .Z(n38653) );
  XOR U59380 ( .A(n38654), .B(n38653), .Z(n38657) );
  XOR U59381 ( .A(n38656), .B(n38657), .Z(n38649) );
  XOR U59382 ( .A(n38648), .B(n38649), .Z(n38652) );
  XOR U59383 ( .A(n38651), .B(n38652), .Z(n44354) );
  XOR U59384 ( .A(n44355), .B(n44354), .Z(n44359) );
  XOR U59385 ( .A(n44357), .B(n44359), .Z(n38646) );
  XOR U59386 ( .A(n38645), .B(n38646), .Z(n44361) );
  XOR U59387 ( .A(n44362), .B(n44361), .Z(n44363) );
  XOR U59388 ( .A(n44365), .B(n44363), .Z(n44369) );
  XOR U59389 ( .A(n44367), .B(n44369), .Z(n44371) );
  XOR U59390 ( .A(n44370), .B(n44371), .Z(n44374) );
  XOR U59391 ( .A(n44375), .B(n44374), .Z(n44376) );
  XOR U59392 ( .A(n44378), .B(n44376), .Z(n44385) );
  XOR U59393 ( .A(n44384), .B(n44385), .Z(n44381) );
  XOR U59394 ( .A(n44380), .B(n44381), .Z(n49125) );
  XOR U59395 ( .A(n49126), .B(n49125), .Z(n54244) );
  XOR U59396 ( .A(n54246), .B(n54244), .Z(n54254) );
  XOR U59397 ( .A(n54253), .B(n54254), .Z(n59562) );
  XOR U59398 ( .A(n59561), .B(n59562), .Z(n59564) );
  XOR U59399 ( .A(n59565), .B(n59564), .Z(n59579) );
  XOR U59400 ( .A(n59581), .B(n59579), .Z(n59605) );
  XOR U59401 ( .A(n59604), .B(n59605), .Z(n59618) );
  XOR U59402 ( .A(n59617), .B(n59618), .Z(n59625) );
  XOR U59403 ( .A(n59626), .B(n59625), .Z(n59647) );
  XOR U59404 ( .A(n59649), .B(n59647), .Z(n64843) );
  XOR U59405 ( .A(n64842), .B(n64843), .Z(n64860) );
  XOR U59406 ( .A(n64859), .B(n64860), .Z(n70019) );
  XOR U59407 ( .A(n70018), .B(n70019), .Z(n75321) );
  XOR U59408 ( .A(n75320), .B(n75321), .Z(n80656) );
  XOR U59409 ( .A(n80655), .B(n80656), .Z(n86365) );
  XOR U59410 ( .A(n86364), .B(n86365), .Z(n86393) );
  XOR U59411 ( .A(n86392), .B(n86393), .Z(n92123) );
  XOR U59412 ( .A(n92122), .B(n92123), .Z(n92148) );
  XOR U59413 ( .A(n92147), .B(n92148), .Z(n92158) );
  XOR U59414 ( .A(n92157), .B(n92158), .Z(n92185) );
  XOR U59415 ( .A(n92184), .B(n92185), .Z(n92218) );
  XOR U59416 ( .A(n92217), .B(n92218), .Z(n92271) );
  XOR U59417 ( .A(n92272), .B(n92271), .Z(o[0]) );
  IV U59418 ( .A(n38645), .Z(n38647) );
  NOR U59419 ( .A(n38647), .B(n38646), .Z(n49107) );
  IV U59420 ( .A(n38648), .Z(n38650) );
  NOR U59421 ( .A(n38650), .B(n38649), .Z(n54207) );
  NOR U59422 ( .A(n38652), .B(n38651), .Z(n54211) );
  NOR U59423 ( .A(n54207), .B(n54211), .Z(n49101) );
  IV U59424 ( .A(n38653), .Z(n38655) );
  NOR U59425 ( .A(n38655), .B(n38654), .Z(n49142) );
  IV U59426 ( .A(n38656), .Z(n38658) );
  NOR U59427 ( .A(n38658), .B(n38657), .Z(n54204) );
  NOR U59428 ( .A(n49142), .B(n54204), .Z(n38659) );
  IV U59429 ( .A(n38659), .Z(n49097) );
  NOR U59430 ( .A(n38661), .B(n38660), .Z(n49096) );
  IV U59431 ( .A(n49096), .Z(n49151) );
  NOR U59432 ( .A(n38663), .B(n38662), .Z(n44416) );
  IV U59433 ( .A(n38664), .Z(n38666) );
  NOR U59434 ( .A(n38666), .B(n38665), .Z(n44403) );
  NOR U59435 ( .A(n44416), .B(n44403), .Z(n44345) );
  NOR U59436 ( .A(n38668), .B(n38667), .Z(n59500) );
  IV U59437 ( .A(n38669), .Z(n38671) );
  NOR U59438 ( .A(n38671), .B(n38670), .Z(n54293) );
  NOR U59439 ( .A(n59500), .B(n54293), .Z(n44422) );
  IV U59440 ( .A(n38672), .Z(n38674) );
  NOR U59441 ( .A(n38674), .B(n38673), .Z(n49171) );
  IV U59442 ( .A(n38675), .Z(n38676) );
  NOR U59443 ( .A(n38677), .B(n38676), .Z(n49167) );
  NOR U59444 ( .A(n49171), .B(n49167), .Z(n44421) );
  IV U59445 ( .A(n38678), .Z(n38679) );
  NOR U59446 ( .A(n38680), .B(n38679), .Z(n44427) );
  IV U59447 ( .A(n38681), .Z(n38682) );
  NOR U59448 ( .A(n38683), .B(n38682), .Z(n49081) );
  NOR U59449 ( .A(n44427), .B(n49081), .Z(n44324) );
  IV U59450 ( .A(n38684), .Z(n38686) );
  NOR U59451 ( .A(n38686), .B(n38685), .Z(n44429) );
  NOR U59452 ( .A(n38688), .B(n38687), .Z(n49068) );
  IV U59453 ( .A(n38689), .Z(n38690) );
  NOR U59454 ( .A(n38691), .B(n38690), .Z(n49070) );
  NOR U59455 ( .A(n49068), .B(n49070), .Z(n44315) );
  IV U59456 ( .A(n38692), .Z(n38694) );
  NOR U59457 ( .A(n38694), .B(n38693), .Z(n49207) );
  IV U59458 ( .A(n38695), .Z(n38696) );
  NOR U59459 ( .A(n38697), .B(n38696), .Z(n49202) );
  NOR U59460 ( .A(n49207), .B(n49202), .Z(n44442) );
  IV U59461 ( .A(n38698), .Z(n38699) );
  NOR U59462 ( .A(n38700), .B(n38699), .Z(n49216) );
  IV U59463 ( .A(n38701), .Z(n38703) );
  NOR U59464 ( .A(n38703), .B(n38702), .Z(n49210) );
  NOR U59465 ( .A(n49216), .B(n49210), .Z(n44446) );
  IV U59466 ( .A(n38704), .Z(n38706) );
  NOR U59467 ( .A(n38706), .B(n38705), .Z(n54330) );
  IV U59468 ( .A(n38707), .Z(n38708) );
  NOR U59469 ( .A(n38709), .B(n38708), .Z(n54322) );
  NOR U59470 ( .A(n54330), .B(n54322), .Z(n49054) );
  IV U59471 ( .A(n38710), .Z(n38711) );
  NOR U59472 ( .A(n38712), .B(n38711), .Z(n49049) );
  IV U59473 ( .A(n38713), .Z(n38714) );
  NOR U59474 ( .A(n38715), .B(n38714), .Z(n49045) );
  NOR U59475 ( .A(n49049), .B(n49045), .Z(n44286) );
  IV U59476 ( .A(n38716), .Z(n38717) );
  NOR U59477 ( .A(n38718), .B(n38717), .Z(n54179) );
  IV U59478 ( .A(n38719), .Z(n38721) );
  NOR U59479 ( .A(n38721), .B(n38720), .Z(n49226) );
  NOR U59480 ( .A(n54179), .B(n49226), .Z(n49040) );
  IV U59481 ( .A(n38722), .Z(n38723) );
  NOR U59482 ( .A(n38724), .B(n38723), .Z(n44278) );
  IV U59483 ( .A(n44278), .Z(n44272) );
  IV U59484 ( .A(n38725), .Z(n38726) );
  NOR U59485 ( .A(n38727), .B(n38726), .Z(n44447) );
  IV U59486 ( .A(n38728), .Z(n38729) );
  NOR U59487 ( .A(n38730), .B(n38729), .Z(n38731) );
  IV U59488 ( .A(n38731), .Z(n49015) );
  IV U59489 ( .A(n38732), .Z(n38733) );
  NOR U59490 ( .A(n38734), .B(n38733), .Z(n49247) );
  IV U59491 ( .A(n38735), .Z(n38736) );
  NOR U59492 ( .A(n38737), .B(n38736), .Z(n49242) );
  NOR U59493 ( .A(n49247), .B(n49242), .Z(n49013) );
  IV U59494 ( .A(n38738), .Z(n38740) );
  NOR U59495 ( .A(n38740), .B(n38739), .Z(n49005) );
  IV U59496 ( .A(n38741), .Z(n38743) );
  NOR U59497 ( .A(n38743), .B(n38742), .Z(n48994) );
  IV U59498 ( .A(n38744), .Z(n38745) );
  NOR U59499 ( .A(n38746), .B(n38745), .Z(n49008) );
  NOR U59500 ( .A(n48994), .B(n49008), .Z(n44232) );
  IV U59501 ( .A(n38747), .Z(n38749) );
  NOR U59502 ( .A(n38749), .B(n38748), .Z(n54395) );
  IV U59503 ( .A(n38750), .Z(n38751) );
  NOR U59504 ( .A(n38752), .B(n38751), .Z(n54387) );
  NOR U59505 ( .A(n54395), .B(n54387), .Z(n48991) );
  IV U59506 ( .A(n38753), .Z(n38754) );
  NOR U59507 ( .A(n38755), .B(n38754), .Z(n44476) );
  IV U59508 ( .A(n38756), .Z(n38758) );
  NOR U59509 ( .A(n38758), .B(n38757), .Z(n48966) );
  IV U59510 ( .A(n38759), .Z(n38760) );
  NOR U59511 ( .A(n38761), .B(n38760), .Z(n48954) );
  IV U59512 ( .A(n38762), .Z(n38763) );
  NOR U59513 ( .A(n38764), .B(n38763), .Z(n48949) );
  IV U59514 ( .A(n38765), .Z(n38767) );
  NOR U59515 ( .A(n38767), .B(n38766), .Z(n44145) );
  IV U59516 ( .A(n44145), .Z(n44139) );
  IV U59517 ( .A(n38768), .Z(n38769) );
  NOR U59518 ( .A(n38770), .B(n38769), .Z(n48944) );
  IV U59519 ( .A(n38771), .Z(n38772) );
  NOR U59520 ( .A(n38773), .B(n38772), .Z(n54445) );
  IV U59521 ( .A(n38774), .Z(n38776) );
  NOR U59522 ( .A(n38776), .B(n38775), .Z(n54438) );
  NOR U59523 ( .A(n54445), .B(n54438), .Z(n48943) );
  IV U59524 ( .A(n38777), .Z(n38778) );
  NOR U59525 ( .A(n38779), .B(n38778), .Z(n48933) );
  IV U59526 ( .A(n38780), .Z(n38781) );
  NOR U59527 ( .A(n38782), .B(n38781), .Z(n44501) );
  NOR U59528 ( .A(n48933), .B(n44501), .Z(n44137) );
  IV U59529 ( .A(n38783), .Z(n38784) );
  NOR U59530 ( .A(n38785), .B(n38784), .Z(n48931) );
  IV U59531 ( .A(n38786), .Z(n38787) );
  NOR U59532 ( .A(n38788), .B(n38787), .Z(n49306) );
  IV U59533 ( .A(n38789), .Z(n38790) );
  NOR U59534 ( .A(n38791), .B(n38790), .Z(n49301) );
  NOR U59535 ( .A(n49306), .B(n49301), .Z(n48923) );
  IV U59536 ( .A(n38792), .Z(n38794) );
  NOR U59537 ( .A(n38794), .B(n38793), .Z(n49313) );
  IV U59538 ( .A(n38795), .Z(n38796) );
  NOR U59539 ( .A(n38797), .B(n38796), .Z(n38798) );
  NOR U59540 ( .A(n49313), .B(n38798), .Z(n44512) );
  IV U59541 ( .A(n38799), .Z(n38800) );
  NOR U59542 ( .A(n38801), .B(n38800), .Z(n44509) );
  IV U59543 ( .A(n38802), .Z(n38803) );
  NOR U59544 ( .A(n38804), .B(n38803), .Z(n48899) );
  IV U59545 ( .A(n38805), .Z(n38807) );
  NOR U59546 ( .A(n38807), .B(n38806), .Z(n48903) );
  NOR U59547 ( .A(n48899), .B(n48903), .Z(n44116) );
  IV U59548 ( .A(n38808), .Z(n38809) );
  NOR U59549 ( .A(n38810), .B(n38809), .Z(n44104) );
  IV U59550 ( .A(n38811), .Z(n38813) );
  NOR U59551 ( .A(n38813), .B(n38812), .Z(n44106) );
  IV U59552 ( .A(n38814), .Z(n38815) );
  NOR U59553 ( .A(n38816), .B(n38815), .Z(n48892) );
  IV U59554 ( .A(n38817), .Z(n38819) );
  NOR U59555 ( .A(n38819), .B(n38818), .Z(n44522) );
  IV U59556 ( .A(n44522), .Z(n44081) );
  IV U59557 ( .A(n38820), .Z(n38822) );
  NOR U59558 ( .A(n38822), .B(n38821), .Z(n54045) );
  IV U59559 ( .A(n38823), .Z(n38825) );
  NOR U59560 ( .A(n38825), .B(n38824), .Z(n54052) );
  NOR U59561 ( .A(n54045), .B(n54052), .Z(n44527) );
  IV U59562 ( .A(n38826), .Z(n38827) );
  NOR U59563 ( .A(n38828), .B(n38827), .Z(n48884) );
  IV U59564 ( .A(n38829), .Z(n38830) );
  NOR U59565 ( .A(n38831), .B(n38830), .Z(n44533) );
  NOR U59566 ( .A(n48884), .B(n44533), .Z(n44074) );
  IV U59567 ( .A(n38832), .Z(n38833) );
  NOR U59568 ( .A(n38834), .B(n38833), .Z(n48881) );
  IV U59569 ( .A(n38838), .Z(n38835) );
  NOR U59570 ( .A(n38835), .B(n38836), .Z(n59823) );
  IV U59571 ( .A(n38836), .Z(n38837) );
  NOR U59572 ( .A(n38838), .B(n38837), .Z(n38840) );
  IV U59573 ( .A(n38839), .Z(n64515) );
  NOR U59574 ( .A(n38840), .B(n64515), .Z(n38841) );
  NOR U59575 ( .A(n59823), .B(n38841), .Z(n48880) );
  IV U59576 ( .A(n38842), .Z(n38843) );
  NOR U59577 ( .A(n38844), .B(n38843), .Z(n44539) );
  IV U59578 ( .A(n38845), .Z(n38846) );
  NOR U59579 ( .A(n38847), .B(n38846), .Z(n44536) );
  NOR U59580 ( .A(n44539), .B(n44536), .Z(n44073) );
  IV U59581 ( .A(n38848), .Z(n38850) );
  NOR U59582 ( .A(n38850), .B(n38849), .Z(n44542) );
  IV U59583 ( .A(n38851), .Z(n38852) );
  NOR U59584 ( .A(n38853), .B(n38852), .Z(n48862) );
  IV U59585 ( .A(n38854), .Z(n38855) );
  NOR U59586 ( .A(n38856), .B(n38855), .Z(n48867) );
  NOR U59587 ( .A(n48862), .B(n48867), .Z(n44064) );
  IV U59588 ( .A(n38857), .Z(n38858) );
  NOR U59589 ( .A(n38859), .B(n38858), .Z(n59839) );
  IV U59590 ( .A(n38860), .Z(n38862) );
  NOR U59591 ( .A(n38862), .B(n38861), .Z(n64502) );
  NOR U59592 ( .A(n59839), .B(n64502), .Z(n54529) );
  IV U59593 ( .A(n38863), .Z(n38864) );
  NOR U59594 ( .A(n38865), .B(n38864), .Z(n44549) );
  IV U59595 ( .A(n38866), .Z(n38867) );
  NOR U59596 ( .A(n38868), .B(n38867), .Z(n44545) );
  NOR U59597 ( .A(n44549), .B(n44545), .Z(n44063) );
  IV U59598 ( .A(n38869), .Z(n38871) );
  NOR U59599 ( .A(n38871), .B(n38870), .Z(n44061) );
  IV U59600 ( .A(n44061), .Z(n44056) );
  IV U59601 ( .A(n38872), .Z(n38873) );
  NOR U59602 ( .A(n38874), .B(n38873), .Z(n48854) );
  IV U59603 ( .A(n38875), .Z(n38876) );
  NOR U59604 ( .A(n38877), .B(n38876), .Z(n54565) );
  IV U59605 ( .A(n38878), .Z(n38879) );
  NOR U59606 ( .A(n38880), .B(n38879), .Z(n54557) );
  NOR U59607 ( .A(n54565), .B(n54557), .Z(n54018) );
  IV U59608 ( .A(n54018), .Z(n44039) );
  IV U59609 ( .A(n38881), .Z(n38883) );
  NOR U59610 ( .A(n38883), .B(n38882), .Z(n48820) );
  IV U59611 ( .A(n38884), .Z(n38885) );
  NOR U59612 ( .A(n38886), .B(n38885), .Z(n49402) );
  IV U59613 ( .A(n38887), .Z(n38888) );
  NOR U59614 ( .A(n38889), .B(n38888), .Z(n53990) );
  NOR U59615 ( .A(n49402), .B(n53990), .Z(n48819) );
  IV U59616 ( .A(n38890), .Z(n38891) );
  NOR U59617 ( .A(n38892), .B(n38891), .Z(n44005) );
  IV U59618 ( .A(n44005), .Z(n43996) );
  IV U59619 ( .A(n38893), .Z(n38894) );
  NOR U59620 ( .A(n38895), .B(n38894), .Z(n38896) );
  IV U59621 ( .A(n38896), .Z(n48798) );
  IV U59622 ( .A(n38897), .Z(n38899) );
  NOR U59623 ( .A(n38899), .B(n38898), .Z(n49454) );
  IV U59624 ( .A(n38900), .Z(n38901) );
  NOR U59625 ( .A(n38902), .B(n38901), .Z(n49450) );
  NOR U59626 ( .A(n49454), .B(n49450), .Z(n48775) );
  NOR U59627 ( .A(n38903), .B(n38904), .Z(n38908) );
  IV U59628 ( .A(n38904), .Z(n38905) );
  NOR U59629 ( .A(n38906), .B(n38905), .Z(n59197) );
  NOR U59630 ( .A(n59205), .B(n59197), .Z(n38907) );
  NOR U59631 ( .A(n38908), .B(n38907), .Z(n44594) );
  IV U59632 ( .A(n38912), .Z(n38909) );
  NOR U59633 ( .A(n38911), .B(n38909), .Z(n44595) );
  NOR U59634 ( .A(n44595), .B(n38910), .Z(n38915) );
  IV U59635 ( .A(n38911), .Z(n38913) );
  NOR U59636 ( .A(n38913), .B(n38912), .Z(n38914) );
  NOR U59637 ( .A(n38915), .B(n38914), .Z(n43940) );
  IV U59638 ( .A(n38916), .Z(n38917) );
  NOR U59639 ( .A(n38918), .B(n38917), .Z(n44608) );
  IV U59640 ( .A(n38919), .Z(n38920) );
  NOR U59641 ( .A(n38921), .B(n38920), .Z(n49482) );
  IV U59642 ( .A(n38922), .Z(n38923) );
  NOR U59643 ( .A(n38924), .B(n38923), .Z(n53921) );
  NOR U59644 ( .A(n49482), .B(n53921), .Z(n44607) );
  IV U59645 ( .A(n38925), .Z(n38926) );
  NOR U59646 ( .A(n38927), .B(n38926), .Z(n43912) );
  IV U59647 ( .A(n43912), .Z(n43902) );
  IV U59648 ( .A(n38928), .Z(n38930) );
  NOR U59649 ( .A(n38930), .B(n38929), .Z(n48741) );
  IV U59650 ( .A(n38931), .Z(n38932) );
  NOR U59651 ( .A(n38933), .B(n38932), .Z(n48725) );
  NOR U59652 ( .A(n48741), .B(n48725), .Z(n43900) );
  IV U59653 ( .A(n38934), .Z(n38935) );
  NOR U59654 ( .A(n38936), .B(n38935), .Z(n48729) );
  IV U59655 ( .A(n38937), .Z(n38938) );
  NOR U59656 ( .A(n38939), .B(n38938), .Z(n48738) );
  NOR U59657 ( .A(n48729), .B(n48738), .Z(n43899) );
  IV U59658 ( .A(n38940), .Z(n38941) );
  NOR U59659 ( .A(n38942), .B(n38941), .Z(n59158) );
  IV U59660 ( .A(n38943), .Z(n38944) );
  NOR U59661 ( .A(n38945), .B(n38944), .Z(n54624) );
  NOR U59662 ( .A(n59158), .B(n54624), .Z(n48716) );
  IV U59663 ( .A(n38946), .Z(n38947) );
  NOR U59664 ( .A(n38948), .B(n38947), .Z(n44638) );
  IV U59665 ( .A(n38949), .Z(n38951) );
  NOR U59666 ( .A(n38951), .B(n38950), .Z(n44623) );
  NOR U59667 ( .A(n44638), .B(n44623), .Z(n43858) );
  IV U59668 ( .A(n38952), .Z(n38954) );
  NOR U59669 ( .A(n38954), .B(n38953), .Z(n53885) );
  IV U59670 ( .A(n38955), .Z(n38956) );
  NOR U59671 ( .A(n38957), .B(n38956), .Z(n53891) );
  NOR U59672 ( .A(n53885), .B(n53891), .Z(n44637) );
  IV U59673 ( .A(n38958), .Z(n38960) );
  NOR U59674 ( .A(n38960), .B(n38959), .Z(n48678) );
  IV U59675 ( .A(n38961), .Z(n38962) );
  NOR U59676 ( .A(n38963), .B(n38962), .Z(n48675) );
  NOR U59677 ( .A(n48678), .B(n48675), .Z(n43857) );
  IV U59678 ( .A(n38964), .Z(n38966) );
  NOR U59679 ( .A(n38966), .B(n38965), .Z(n49536) );
  IV U59680 ( .A(n38967), .Z(n38968) );
  NOR U59681 ( .A(n38969), .B(n38968), .Z(n49532) );
  NOR U59682 ( .A(n49536), .B(n49532), .Z(n44645) );
  IV U59683 ( .A(n38970), .Z(n38971) );
  NOR U59684 ( .A(n38972), .B(n38971), .Z(n44642) );
  IV U59685 ( .A(n38973), .Z(n38974) );
  NOR U59686 ( .A(n38975), .B(n38974), .Z(n43838) );
  IV U59687 ( .A(n38976), .Z(n38978) );
  NOR U59688 ( .A(n38978), .B(n38977), .Z(n48639) );
  IV U59689 ( .A(n38979), .Z(n38980) );
  NOR U59690 ( .A(n38981), .B(n38980), .Z(n48634) );
  IV U59691 ( .A(n38982), .Z(n38984) );
  NOR U59692 ( .A(n38984), .B(n38983), .Z(n48642) );
  NOR U59693 ( .A(n48634), .B(n48642), .Z(n43822) );
  IV U59694 ( .A(n38985), .Z(n38987) );
  NOR U59695 ( .A(n38987), .B(n38986), .Z(n53861) );
  IV U59696 ( .A(n38988), .Z(n38990) );
  NOR U59697 ( .A(n38990), .B(n38989), .Z(n53868) );
  NOR U59698 ( .A(n53861), .B(n53868), .Z(n48626) );
  IV U59699 ( .A(n38991), .Z(n38992) );
  NOR U59700 ( .A(n38993), .B(n38992), .Z(n44662) );
  IV U59701 ( .A(n38994), .Z(n38995) );
  NOR U59702 ( .A(n38996), .B(n38995), .Z(n48596) );
  IV U59703 ( .A(n38997), .Z(n38999) );
  NOR U59704 ( .A(n38999), .B(n38998), .Z(n48587) );
  IV U59705 ( .A(n39000), .Z(n39001) );
  NOR U59706 ( .A(n39002), .B(n39001), .Z(n59076) );
  IV U59707 ( .A(n39003), .Z(n39004) );
  NOR U59708 ( .A(n39005), .B(n39004), .Z(n54721) );
  NOR U59709 ( .A(n59076), .B(n54721), .Z(n48580) );
  IV U59710 ( .A(n39006), .Z(n39008) );
  NOR U59711 ( .A(n39008), .B(n39007), .Z(n49585) );
  IV U59712 ( .A(n39009), .Z(n39011) );
  NOR U59713 ( .A(n39011), .B(n39010), .Z(n49579) );
  NOR U59714 ( .A(n49585), .B(n49579), .Z(n44675) );
  IV U59715 ( .A(n39012), .Z(n39014) );
  NOR U59716 ( .A(n39014), .B(n39013), .Z(n49592) );
  IV U59717 ( .A(n39015), .Z(n39017) );
  NOR U59718 ( .A(n39017), .B(n39016), .Z(n49588) );
  NOR U59719 ( .A(n49592), .B(n49588), .Z(n48572) );
  IV U59720 ( .A(n39018), .Z(n39019) );
  NOR U59721 ( .A(n39020), .B(n39019), .Z(n53819) );
  IV U59722 ( .A(n39021), .Z(n39022) );
  NOR U59723 ( .A(n39023), .B(n39022), .Z(n39024) );
  NOR U59724 ( .A(n53819), .B(n39024), .Z(n48570) );
  IV U59725 ( .A(n39025), .Z(n39026) );
  NOR U59726 ( .A(n39027), .B(n39026), .Z(n44676) );
  NOR U59727 ( .A(n39029), .B(n39028), .Z(n48567) );
  NOR U59728 ( .A(n44676), .B(n48567), .Z(n43774) );
  IV U59729 ( .A(n39030), .Z(n39031) );
  NOR U59730 ( .A(n39032), .B(n39031), .Z(n44680) );
  IV U59731 ( .A(n39033), .Z(n39035) );
  NOR U59732 ( .A(n39035), .B(n39034), .Z(n60044) );
  IV U59733 ( .A(n39036), .Z(n39038) );
  NOR U59734 ( .A(n39038), .B(n39037), .Z(n60036) );
  NOR U59735 ( .A(n60044), .B(n60036), .Z(n44679) );
  IV U59736 ( .A(n39039), .Z(n39040) );
  NOR U59737 ( .A(n39041), .B(n39040), .Z(n48558) );
  IV U59738 ( .A(n39042), .Z(n39043) );
  NOR U59739 ( .A(n39044), .B(n39043), .Z(n48554) );
  NOR U59740 ( .A(n48558), .B(n48554), .Z(n43773) );
  IV U59741 ( .A(n39045), .Z(n39046) );
  NOR U59742 ( .A(n39047), .B(n39046), .Z(n48561) );
  IV U59743 ( .A(n39048), .Z(n39050) );
  NOR U59744 ( .A(n39050), .B(n39049), .Z(n48546) );
  IV U59745 ( .A(n39051), .Z(n39052) );
  NOR U59746 ( .A(n39053), .B(n39052), .Z(n48544) );
  NOR U59747 ( .A(n48546), .B(n48544), .Z(n43766) );
  IV U59748 ( .A(n39054), .Z(n39055) );
  NOR U59749 ( .A(n39056), .B(n39055), .Z(n48537) );
  IV U59750 ( .A(n39057), .Z(n39058) );
  NOR U59751 ( .A(n39059), .B(n39058), .Z(n48539) );
  NOR U59752 ( .A(n48537), .B(n48539), .Z(n39060) );
  IV U59753 ( .A(n39060), .Z(n43765) );
  NOR U59754 ( .A(n39061), .B(n44683), .Z(n44691) );
  IV U59755 ( .A(n44683), .Z(n39062) );
  NOR U59756 ( .A(n44684), .B(n39062), .Z(n39063) );
  NOR U59757 ( .A(n39063), .B(n44686), .Z(n39064) );
  NOR U59758 ( .A(n44691), .B(n39064), .Z(n43764) );
  IV U59759 ( .A(n39065), .Z(n39067) );
  NOR U59760 ( .A(n39067), .B(n39066), .Z(n43762) );
  IV U59761 ( .A(n43762), .Z(n43753) );
  IV U59762 ( .A(n39068), .Z(n39069) );
  NOR U59763 ( .A(n39070), .B(n39069), .Z(n48512) );
  IV U59764 ( .A(n39071), .Z(n39072) );
  NOR U59765 ( .A(n39073), .B(n39072), .Z(n44702) );
  NOR U59766 ( .A(n48512), .B(n44702), .Z(n43730) );
  IV U59767 ( .A(n39074), .Z(n39076) );
  NOR U59768 ( .A(n39076), .B(n39075), .Z(n59018) );
  IV U59769 ( .A(n39077), .Z(n39078) );
  NOR U59770 ( .A(n39079), .B(n39078), .Z(n54776) );
  NOR U59771 ( .A(n59018), .B(n54776), .Z(n48511) );
  IV U59772 ( .A(n39080), .Z(n39081) );
  NOR U59773 ( .A(n39082), .B(n39081), .Z(n48496) );
  IV U59774 ( .A(n39083), .Z(n39085) );
  NOR U59775 ( .A(n39085), .B(n39084), .Z(n48500) );
  NOR U59776 ( .A(n48496), .B(n48500), .Z(n43729) );
  IV U59777 ( .A(n39086), .Z(n39088) );
  NOR U59778 ( .A(n39088), .B(n39087), .Z(n48485) );
  IV U59779 ( .A(n39089), .Z(n39090) );
  NOR U59780 ( .A(n39091), .B(n39090), .Z(n44705) );
  IV U59781 ( .A(n39092), .Z(n39094) );
  NOR U59782 ( .A(n39094), .B(n39093), .Z(n48489) );
  NOR U59783 ( .A(n44705), .B(n48489), .Z(n49625) );
  IV U59784 ( .A(n39095), .Z(n39097) );
  NOR U59785 ( .A(n39097), .B(n39096), .Z(n44709) );
  IV U59786 ( .A(n39098), .Z(n39099) );
  NOR U59787 ( .A(n39100), .B(n39099), .Z(n44707) );
  NOR U59788 ( .A(n44709), .B(n44707), .Z(n43728) );
  IV U59789 ( .A(n39101), .Z(n39102) );
  NOR U59790 ( .A(n39103), .B(n39102), .Z(n54797) );
  IV U59791 ( .A(n39104), .Z(n39105) );
  NOR U59792 ( .A(n39106), .B(n39105), .Z(n54789) );
  NOR U59793 ( .A(n54797), .B(n54789), .Z(n48478) );
  IV U59794 ( .A(n39107), .Z(n39109) );
  NOR U59795 ( .A(n39109), .B(n39108), .Z(n44714) );
  IV U59796 ( .A(n39110), .Z(n39112) );
  NOR U59797 ( .A(n39112), .B(n39111), .Z(n48472) );
  NOR U59798 ( .A(n44714), .B(n48472), .Z(n43721) );
  IV U59799 ( .A(n39113), .Z(n39115) );
  NOR U59800 ( .A(n39115), .B(n39114), .Z(n44722) );
  NOR U59801 ( .A(n39117), .B(n39116), .Z(n53730) );
  NOR U59802 ( .A(n39119), .B(n39118), .Z(n39121) );
  IV U59803 ( .A(n39120), .Z(n49653) );
  NOR U59804 ( .A(n39121), .B(n49653), .Z(n39122) );
  NOR U59805 ( .A(n53730), .B(n39122), .Z(n44727) );
  IV U59806 ( .A(n39123), .Z(n39125) );
  NOR U59807 ( .A(n39125), .B(n39124), .Z(n44733) );
  IV U59808 ( .A(n39126), .Z(n39128) );
  NOR U59809 ( .A(n39128), .B(n39127), .Z(n44738) );
  IV U59810 ( .A(n39129), .Z(n39130) );
  NOR U59811 ( .A(n39131), .B(n39130), .Z(n60138) );
  IV U59812 ( .A(n39132), .Z(n39133) );
  NOR U59813 ( .A(n39134), .B(n39133), .Z(n60143) );
  NOR U59814 ( .A(n60138), .B(n60143), .Z(n53716) );
  IV U59815 ( .A(n39135), .Z(n39136) );
  NOR U59816 ( .A(n39137), .B(n39136), .Z(n48454) );
  IV U59817 ( .A(n39138), .Z(n39139) );
  NOR U59818 ( .A(n39140), .B(n39139), .Z(n48458) );
  NOR U59819 ( .A(n48454), .B(n48458), .Z(n39141) );
  IV U59820 ( .A(n39141), .Z(n43680) );
  IV U59821 ( .A(n39142), .Z(n39143) );
  NOR U59822 ( .A(n39144), .B(n39143), .Z(n54828) );
  IV U59823 ( .A(n39145), .Z(n39146) );
  NOR U59824 ( .A(n39147), .B(n39146), .Z(n54820) );
  NOR U59825 ( .A(n54828), .B(n54820), .Z(n48450) );
  IV U59826 ( .A(n39148), .Z(n39150) );
  NOR U59827 ( .A(n39150), .B(n39149), .Z(n43653) );
  IV U59828 ( .A(n43653), .Z(n43644) );
  IV U59829 ( .A(n39151), .Z(n39152) );
  NOR U59830 ( .A(n39153), .B(n39152), .Z(n49686) );
  IV U59831 ( .A(n39154), .Z(n39155) );
  NOR U59832 ( .A(n39156), .B(n39155), .Z(n44754) );
  NOR U59833 ( .A(n49686), .B(n44754), .Z(n43642) );
  IV U59834 ( .A(n39157), .Z(n39158) );
  NOR U59835 ( .A(n39159), .B(n39158), .Z(n43633) );
  IV U59836 ( .A(n43633), .Z(n43626) );
  IV U59837 ( .A(n39160), .Z(n39161) );
  NOR U59838 ( .A(n39162), .B(n39161), .Z(n48424) );
  IV U59839 ( .A(n39163), .Z(n39165) );
  NOR U59840 ( .A(n39165), .B(n39164), .Z(n48412) );
  IV U59841 ( .A(n39166), .Z(n39167) );
  NOR U59842 ( .A(n39168), .B(n39167), .Z(n43602) );
  IV U59843 ( .A(n43602), .Z(n43592) );
  IV U59844 ( .A(n39169), .Z(n39170) );
  NOR U59845 ( .A(n39171), .B(n39170), .Z(n43589) );
  IV U59846 ( .A(n43589), .Z(n43584) );
  IV U59847 ( .A(n39172), .Z(n39173) );
  NOR U59848 ( .A(n39174), .B(n39173), .Z(n44781) );
  IV U59849 ( .A(n39175), .Z(n39177) );
  NOR U59850 ( .A(n39177), .B(n39176), .Z(n44796) );
  IV U59851 ( .A(n39178), .Z(n39180) );
  NOR U59852 ( .A(n39180), .B(n39179), .Z(n44827) );
  IV U59853 ( .A(n39181), .Z(n39182) );
  NOR U59854 ( .A(n39183), .B(n39182), .Z(n44825) );
  NOR U59855 ( .A(n44827), .B(n44825), .Z(n43533) );
  IV U59856 ( .A(n64081), .Z(n39184) );
  NOR U59857 ( .A(n64082), .B(n39184), .Z(n64100) );
  NOR U59858 ( .A(n39185), .B(n64081), .Z(n39187) );
  IV U59859 ( .A(n39186), .Z(n64084) );
  NOR U59860 ( .A(n39187), .B(n64084), .Z(n39188) );
  NOR U59861 ( .A(n64100), .B(n39188), .Z(n44830) );
  IV U59862 ( .A(n39189), .Z(n39191) );
  NOR U59863 ( .A(n39191), .B(n39190), .Z(n53573) );
  IV U59864 ( .A(n39192), .Z(n39193) );
  NOR U59865 ( .A(n39194), .B(n39193), .Z(n49720) );
  NOR U59866 ( .A(n53573), .B(n49720), .Z(n48395) );
  IV U59867 ( .A(n39195), .Z(n39196) );
  NOR U59868 ( .A(n39197), .B(n39196), .Z(n48384) );
  IV U59869 ( .A(n39198), .Z(n39200) );
  NOR U59870 ( .A(n39200), .B(n39199), .Z(n48396) );
  NOR U59871 ( .A(n48384), .B(n48396), .Z(n43528) );
  IV U59872 ( .A(n39201), .Z(n39202) );
  NOR U59873 ( .A(n39203), .B(n39202), .Z(n48388) );
  IV U59874 ( .A(n39204), .Z(n39205) );
  NOR U59875 ( .A(n39206), .B(n39205), .Z(n54928) );
  IV U59876 ( .A(n39207), .Z(n39209) );
  NOR U59877 ( .A(n39209), .B(n39208), .Z(n54923) );
  NOR U59878 ( .A(n54928), .B(n54923), .Z(n48387) );
  IV U59879 ( .A(n39210), .Z(n39212) );
  NOR U59880 ( .A(n39212), .B(n39211), .Z(n44837) );
  IV U59881 ( .A(n39213), .Z(n39215) );
  NOR U59882 ( .A(n39215), .B(n39214), .Z(n44834) );
  NOR U59883 ( .A(n44837), .B(n44834), .Z(n43527) );
  NOR U59884 ( .A(n39217), .B(n39216), .Z(n48377) );
  IV U59885 ( .A(n39218), .Z(n39219) );
  NOR U59886 ( .A(n39220), .B(n39219), .Z(n60259) );
  IV U59887 ( .A(n39221), .Z(n39222) );
  NOR U59888 ( .A(n39223), .B(n39222), .Z(n60251) );
  NOR U59889 ( .A(n60259), .B(n60251), .Z(n48372) );
  IV U59890 ( .A(n39224), .Z(n39226) );
  NOR U59891 ( .A(n39226), .B(n39225), .Z(n43484) );
  IV U59892 ( .A(n43484), .Z(n43479) );
  IV U59893 ( .A(n39227), .Z(n39228) );
  NOR U59894 ( .A(n39229), .B(n39228), .Z(n48339) );
  IV U59895 ( .A(n39230), .Z(n39232) );
  NOR U59896 ( .A(n39232), .B(n39231), .Z(n49758) );
  IV U59897 ( .A(n39233), .Z(n39234) );
  NOR U59898 ( .A(n39235), .B(n39234), .Z(n49754) );
  NOR U59899 ( .A(n49758), .B(n49754), .Z(n48331) );
  IV U59900 ( .A(n39236), .Z(n39237) );
  NOR U59901 ( .A(n39238), .B(n39237), .Z(n43464) );
  IV U59902 ( .A(n43464), .Z(n43458) );
  IV U59903 ( .A(n39239), .Z(n39240) );
  NOR U59904 ( .A(n39241), .B(n39240), .Z(n43461) );
  IV U59905 ( .A(n43461), .Z(n48324) );
  IV U59906 ( .A(n39242), .Z(n39243) );
  NOR U59907 ( .A(n39244), .B(n39243), .Z(n44843) );
  IV U59908 ( .A(n39245), .Z(n39247) );
  NOR U59909 ( .A(n39247), .B(n39246), .Z(n44846) );
  NOR U59910 ( .A(n44843), .B(n44846), .Z(n43450) );
  IV U59911 ( .A(n39248), .Z(n39249) );
  NOR U59912 ( .A(n39250), .B(n39249), .Z(n43446) );
  IV U59913 ( .A(n39251), .Z(n39252) );
  NOR U59914 ( .A(n39253), .B(n39252), .Z(n48304) );
  IV U59915 ( .A(n39254), .Z(n39256) );
  NOR U59916 ( .A(n39256), .B(n39255), .Z(n48310) );
  NOR U59917 ( .A(n48304), .B(n48310), .Z(n43437) );
  NOR U59918 ( .A(n39258), .B(n39257), .Z(n44853) );
  IV U59919 ( .A(n39259), .Z(n39261) );
  NOR U59920 ( .A(n39261), .B(n39260), .Z(n48306) );
  NOR U59921 ( .A(n44853), .B(n48306), .Z(n43436) );
  IV U59922 ( .A(n39262), .Z(n39263) );
  NOR U59923 ( .A(n39264), .B(n39263), .Z(n44851) );
  IV U59924 ( .A(n39265), .Z(n39266) );
  NOR U59925 ( .A(n39267), .B(n39266), .Z(n49808) );
  IV U59926 ( .A(n39268), .Z(n39270) );
  NOR U59927 ( .A(n39270), .B(n39269), .Z(n49802) );
  NOR U59928 ( .A(n49808), .B(n49802), .Z(n39271) );
  IV U59929 ( .A(n39271), .Z(n48285) );
  IV U59930 ( .A(n39272), .Z(n39274) );
  NOR U59931 ( .A(n39274), .B(n39273), .Z(n49816) );
  IV U59932 ( .A(n39275), .Z(n39277) );
  NOR U59933 ( .A(n39277), .B(n39276), .Z(n49811) );
  NOR U59934 ( .A(n49816), .B(n49811), .Z(n48283) );
  IV U59935 ( .A(n39278), .Z(n39279) );
  NOR U59936 ( .A(n39280), .B(n39279), .Z(n48266) );
  IV U59937 ( .A(n39281), .Z(n39282) );
  NOR U59938 ( .A(n39283), .B(n39282), .Z(n43407) );
  IV U59939 ( .A(n43407), .Z(n43400) );
  IV U59940 ( .A(n39284), .Z(n39286) );
  NOR U59941 ( .A(n39286), .B(n39285), .Z(n48258) );
  IV U59942 ( .A(n39287), .Z(n39289) );
  NOR U59943 ( .A(n39289), .B(n39288), .Z(n39290) );
  IV U59944 ( .A(n39290), .Z(n44865) );
  IV U59945 ( .A(n39291), .Z(n39292) );
  NOR U59946 ( .A(n39293), .B(n39292), .Z(n53448) );
  IV U59947 ( .A(n39294), .Z(n39296) );
  NOR U59948 ( .A(n39296), .B(n39295), .Z(n53441) );
  NOR U59949 ( .A(n53448), .B(n53441), .Z(n44870) );
  IV U59950 ( .A(n39297), .Z(n39299) );
  NOR U59951 ( .A(n39299), .B(n39298), .Z(n58733) );
  IV U59952 ( .A(n39300), .Z(n39301) );
  NOR U59953 ( .A(n39302), .B(n39301), .Z(n58740) );
  NOR U59954 ( .A(n58733), .B(n58740), .Z(n49834) );
  IV U59955 ( .A(n39303), .Z(n39304) );
  NOR U59956 ( .A(n39305), .B(n39304), .Z(n43385) );
  IV U59957 ( .A(n39306), .Z(n39308) );
  NOR U59958 ( .A(n39308), .B(n39307), .Z(n44872) );
  IV U59959 ( .A(n39309), .Z(n39310) );
  NOR U59960 ( .A(n39311), .B(n39310), .Z(n43327) );
  IV U59961 ( .A(n43327), .Z(n43322) );
  IV U59962 ( .A(n39312), .Z(n39314) );
  NOR U59963 ( .A(n39314), .B(n39313), .Z(n44892) );
  IV U59964 ( .A(n39315), .Z(n39316) );
  NOR U59965 ( .A(n39317), .B(n39316), .Z(n39318) );
  IV U59966 ( .A(n39318), .Z(n48226) );
  IV U59967 ( .A(n39319), .Z(n39321) );
  NOR U59968 ( .A(n39321), .B(n39320), .Z(n48212) );
  IV U59969 ( .A(n39322), .Z(n39324) );
  NOR U59970 ( .A(n39324), .B(n39323), .Z(n48222) );
  NOR U59971 ( .A(n48212), .B(n48222), .Z(n43276) );
  IV U59972 ( .A(n39325), .Z(n39326) );
  NOR U59973 ( .A(n39327), .B(n39326), .Z(n44935) );
  IV U59974 ( .A(n39328), .Z(n39330) );
  NOR U59975 ( .A(n39330), .B(n39329), .Z(n44930) );
  NOR U59976 ( .A(n44935), .B(n44930), .Z(n43268) );
  IV U59977 ( .A(n39331), .Z(n39332) );
  NOR U59978 ( .A(n39333), .B(n39332), .Z(n44933) );
  IV U59979 ( .A(n39334), .Z(n39335) );
  NOR U59980 ( .A(n39336), .B(n39335), .Z(n48202) );
  IV U59981 ( .A(n39337), .Z(n39338) );
  NOR U59982 ( .A(n39339), .B(n39338), .Z(n44938) );
  NOR U59983 ( .A(n48202), .B(n44938), .Z(n43261) );
  IV U59984 ( .A(n39340), .Z(n39342) );
  NOR U59985 ( .A(n39342), .B(n39341), .Z(n39343) );
  IV U59986 ( .A(n39343), .Z(n43256) );
  IV U59987 ( .A(n39344), .Z(n39345) );
  NOR U59988 ( .A(n39346), .B(n39345), .Z(n48185) );
  IV U59989 ( .A(n39347), .Z(n39349) );
  NOR U59990 ( .A(n39349), .B(n39348), .Z(n48183) );
  NOR U59991 ( .A(n48185), .B(n48183), .Z(n43242) );
  IV U59992 ( .A(n39350), .Z(n39351) );
  NOR U59993 ( .A(n39352), .B(n39351), .Z(n49928) );
  IV U59994 ( .A(n39353), .Z(n39354) );
  NOR U59995 ( .A(n39355), .B(n39354), .Z(n53365) );
  NOR U59996 ( .A(n49928), .B(n53365), .Z(n44951) );
  IV U59997 ( .A(n39356), .Z(n39358) );
  NOR U59998 ( .A(n39358), .B(n39357), .Z(n48178) );
  IV U59999 ( .A(n39359), .Z(n39361) );
  NOR U60000 ( .A(n39361), .B(n39360), .Z(n48160) );
  IV U60001 ( .A(n39362), .Z(n39364) );
  NOR U60002 ( .A(n39364), .B(n39363), .Z(n48158) );
  NOR U60003 ( .A(n48160), .B(n48158), .Z(n39365) );
  IV U60004 ( .A(n39365), .Z(n43228) );
  IV U60005 ( .A(n39366), .Z(n39368) );
  NOR U60006 ( .A(n39368), .B(n39367), .Z(n49946) );
  IV U60007 ( .A(n39369), .Z(n39370) );
  NOR U60008 ( .A(n39371), .B(n39370), .Z(n49941) );
  NOR U60009 ( .A(n49946), .B(n49941), .Z(n48149) );
  IV U60010 ( .A(n39372), .Z(n39373) );
  NOR U60011 ( .A(n39374), .B(n39373), .Z(n44966) );
  IV U60012 ( .A(n39375), .Z(n39376) );
  NOR U60013 ( .A(n39377), .B(n39376), .Z(n44964) );
  NOR U60014 ( .A(n44966), .B(n44964), .Z(n43215) );
  IV U60015 ( .A(n39378), .Z(n39379) );
  NOR U60016 ( .A(n39380), .B(n39379), .Z(n53323) );
  IV U60017 ( .A(n39381), .Z(n39382) );
  NOR U60018 ( .A(n39383), .B(n39382), .Z(n53330) );
  NOR U60019 ( .A(n53323), .B(n53330), .Z(n48145) );
  IV U60020 ( .A(n39384), .Z(n39386) );
  NOR U60021 ( .A(n39386), .B(n39385), .Z(n48132) );
  IV U60022 ( .A(n39387), .Z(n39388) );
  NOR U60023 ( .A(n39389), .B(n39388), .Z(n48136) );
  NOR U60024 ( .A(n48132), .B(n48136), .Z(n44970) );
  IV U60025 ( .A(n39390), .Z(n39392) );
  NOR U60026 ( .A(n39392), .B(n39391), .Z(n44973) );
  IV U60027 ( .A(n39393), .Z(n39394) );
  NOR U60028 ( .A(n39395), .B(n39394), .Z(n44971) );
  NOR U60029 ( .A(n44973), .B(n44971), .Z(n43208) );
  IV U60030 ( .A(n39396), .Z(n39397) );
  NOR U60031 ( .A(n39398), .B(n39397), .Z(n58576) );
  IV U60032 ( .A(n39399), .Z(n39400) );
  NOR U60033 ( .A(n39401), .B(n39400), .Z(n58586) );
  NOR U60034 ( .A(n58576), .B(n58586), .Z(n44977) );
  IV U60035 ( .A(n39402), .Z(n39404) );
  NOR U60036 ( .A(n39404), .B(n39403), .Z(n53319) );
  IV U60037 ( .A(n39405), .Z(n39406) );
  NOR U60038 ( .A(n39407), .B(n39406), .Z(n49968) );
  NOR U60039 ( .A(n53319), .B(n49968), .Z(n44978) );
  IV U60040 ( .A(n39408), .Z(n39410) );
  NOR U60041 ( .A(n39410), .B(n39409), .Z(n44985) );
  IV U60042 ( .A(n39411), .Z(n39412) );
  NOR U60043 ( .A(n39413), .B(n39412), .Z(n48111) );
  NOR U60044 ( .A(n44985), .B(n48111), .Z(n43200) );
  IV U60045 ( .A(n39414), .Z(n39415) );
  NOR U60046 ( .A(n39416), .B(n39415), .Z(n44989) );
  IV U60047 ( .A(n39417), .Z(n39418) );
  NOR U60048 ( .A(n39419), .B(n39418), .Z(n44992) );
  NOR U60049 ( .A(n44989), .B(n44992), .Z(n43193) );
  IV U60050 ( .A(n39420), .Z(n39422) );
  NOR U60051 ( .A(n39422), .B(n39421), .Z(n39423) );
  IV U60052 ( .A(n39423), .Z(n43188) );
  IV U60053 ( .A(n39424), .Z(n39425) );
  NOR U60054 ( .A(n39426), .B(n39425), .Z(n48102) );
  IV U60055 ( .A(n39427), .Z(n39429) );
  NOR U60056 ( .A(n39429), .B(n39428), .Z(n45004) );
  IV U60057 ( .A(n39430), .Z(n39431) );
  NOR U60058 ( .A(n39432), .B(n39431), .Z(n48098) );
  NOR U60059 ( .A(n45004), .B(n48098), .Z(n43174) );
  IV U60060 ( .A(n39433), .Z(n39435) );
  NOR U60061 ( .A(n39435), .B(n39434), .Z(n53303) );
  IV U60062 ( .A(n39436), .Z(n39437) );
  NOR U60063 ( .A(n39438), .B(n39437), .Z(n50004) );
  NOR U60064 ( .A(n53303), .B(n50004), .Z(n45008) );
  IV U60065 ( .A(n39439), .Z(n39440) );
  NOR U60066 ( .A(n39441), .B(n39440), .Z(n48081) );
  IV U60067 ( .A(n39442), .Z(n39443) );
  NOR U60068 ( .A(n39444), .B(n39443), .Z(n45009) );
  NOR U60069 ( .A(n48081), .B(n45009), .Z(n43173) );
  IV U60070 ( .A(n39445), .Z(n39446) );
  NOR U60071 ( .A(n39447), .B(n39446), .Z(n48079) );
  IV U60072 ( .A(n39448), .Z(n39449) );
  NOR U60073 ( .A(n39450), .B(n39449), .Z(n55162) );
  IV U60074 ( .A(n39451), .Z(n39453) );
  NOR U60075 ( .A(n39453), .B(n39452), .Z(n55154) );
  NOR U60076 ( .A(n55162), .B(n55154), .Z(n48087) );
  IV U60077 ( .A(n39454), .Z(n39456) );
  NOR U60078 ( .A(n39456), .B(n39455), .Z(n45013) );
  IV U60079 ( .A(n39457), .Z(n39458) );
  NOR U60080 ( .A(n39459), .B(n39458), .Z(n48076) );
  NOR U60081 ( .A(n45013), .B(n48076), .Z(n43172) );
  IV U60082 ( .A(n39460), .Z(n39462) );
  NOR U60083 ( .A(n39462), .B(n39461), .Z(n48056) );
  IV U60084 ( .A(n39463), .Z(n39464) );
  NOR U60085 ( .A(n39465), .B(n39464), .Z(n48050) );
  IV U60086 ( .A(n39466), .Z(n39467) );
  NOR U60087 ( .A(n39468), .B(n39467), .Z(n55173) );
  NOR U60088 ( .A(n48050), .B(n55173), .Z(n48063) );
  IV U60089 ( .A(n39469), .Z(n39471) );
  NOR U60090 ( .A(n39471), .B(n39470), .Z(n50015) );
  IV U60091 ( .A(n39472), .Z(n39473) );
  NOR U60092 ( .A(n39474), .B(n39473), .Z(n39475) );
  NOR U60093 ( .A(n50015), .B(n39475), .Z(n45016) );
  IV U60094 ( .A(n39476), .Z(n39477) );
  NOR U60095 ( .A(n39478), .B(n39477), .Z(n48041) );
  IV U60096 ( .A(n39479), .Z(n39481) );
  NOR U60097 ( .A(n39481), .B(n39480), .Z(n48019) );
  IV U60098 ( .A(n39482), .Z(n39484) );
  NOR U60099 ( .A(n39484), .B(n39483), .Z(n45017) );
  NOR U60100 ( .A(n48019), .B(n45017), .Z(n43164) );
  IV U60101 ( .A(n39485), .Z(n39486) );
  NOR U60102 ( .A(n39487), .B(n39486), .Z(n48021) );
  IV U60103 ( .A(n39488), .Z(n39489) );
  NOR U60104 ( .A(n39490), .B(n39489), .Z(n47997) );
  IV U60105 ( .A(n39491), .Z(n39493) );
  NOR U60106 ( .A(n39493), .B(n39492), .Z(n47993) );
  NOR U60107 ( .A(n47997), .B(n47993), .Z(n43155) );
  IV U60108 ( .A(n39494), .Z(n39496) );
  NOR U60109 ( .A(n39496), .B(n39495), .Z(n47978) );
  IV U60110 ( .A(n39497), .Z(n39498) );
  NOR U60111 ( .A(n39499), .B(n39498), .Z(n45022) );
  IV U60112 ( .A(n39500), .Z(n39501) );
  NOR U60113 ( .A(n39502), .B(n39501), .Z(n47977) );
  NOR U60114 ( .A(n45022), .B(n47977), .Z(n43150) );
  IV U60115 ( .A(n39503), .Z(n39505) );
  NOR U60116 ( .A(n39505), .B(n39504), .Z(n55203) );
  IV U60117 ( .A(n39506), .Z(n39507) );
  NOR U60118 ( .A(n39508), .B(n39507), .Z(n58499) );
  NOR U60119 ( .A(n55203), .B(n58499), .Z(n47971) );
  IV U60120 ( .A(n39509), .Z(n39510) );
  NOR U60121 ( .A(n39511), .B(n39510), .Z(n45025) );
  IV U60122 ( .A(n39512), .Z(n39514) );
  NOR U60123 ( .A(n39514), .B(n39513), .Z(n47972) );
  NOR U60124 ( .A(n45025), .B(n47972), .Z(n43149) );
  IV U60125 ( .A(n39515), .Z(n39516) );
  NOR U60126 ( .A(n39517), .B(n39516), .Z(n45030) );
  IV U60127 ( .A(n39518), .Z(n39519) );
  NOR U60128 ( .A(n39520), .B(n39519), .Z(n47945) );
  IV U60129 ( .A(n39521), .Z(n39522) );
  NOR U60130 ( .A(n39523), .B(n39522), .Z(n47943) );
  NOR U60131 ( .A(n47945), .B(n47943), .Z(n43113) );
  IV U60132 ( .A(n39524), .Z(n39526) );
  NOR U60133 ( .A(n39526), .B(n39525), .Z(n47925) );
  IV U60134 ( .A(n39527), .Z(n39528) );
  NOR U60135 ( .A(n39529), .B(n39528), .Z(n47933) );
  NOR U60136 ( .A(n47925), .B(n47933), .Z(n43104) );
  IV U60137 ( .A(n39530), .Z(n39531) );
  NOR U60138 ( .A(n39532), .B(n39531), .Z(n43099) );
  IV U60139 ( .A(n39533), .Z(n39534) );
  NOR U60140 ( .A(n39535), .B(n39534), .Z(n43097) );
  IV U60141 ( .A(n43097), .Z(n43092) );
  IV U60142 ( .A(n39536), .Z(n39538) );
  NOR U60143 ( .A(n39538), .B(n39537), .Z(n47916) );
  IV U60144 ( .A(n39539), .Z(n39540) );
  NOR U60145 ( .A(n39541), .B(n39540), .Z(n53234) );
  IV U60146 ( .A(n39542), .Z(n39543) );
  NOR U60147 ( .A(n39544), .B(n39543), .Z(n39545) );
  NOR U60148 ( .A(n53234), .B(n39545), .Z(n45054) );
  IV U60149 ( .A(n39546), .Z(n39548) );
  NOR U60150 ( .A(n39548), .B(n39547), .Z(n45058) );
  IV U60151 ( .A(n39549), .Z(n39550) );
  NOR U60152 ( .A(n39551), .B(n39550), .Z(n45055) );
  NOR U60153 ( .A(n45058), .B(n45055), .Z(n43090) );
  IV U60154 ( .A(n39552), .Z(n39554) );
  NOR U60155 ( .A(n39554), .B(n39553), .Z(n43064) );
  IV U60156 ( .A(n39555), .Z(n39556) );
  NOR U60157 ( .A(n39557), .B(n39556), .Z(n45068) );
  IV U60158 ( .A(n39558), .Z(n39560) );
  NOR U60159 ( .A(n39560), .B(n39559), .Z(n45066) );
  NOR U60160 ( .A(n45068), .B(n45066), .Z(n43063) );
  IV U60161 ( .A(n39561), .Z(n39563) );
  NOR U60162 ( .A(n39563), .B(n39562), .Z(n58391) );
  IV U60163 ( .A(n39564), .Z(n39565) );
  NOR U60164 ( .A(n39566), .B(n39565), .Z(n39567) );
  NOR U60165 ( .A(n58391), .B(n39567), .Z(n45072) );
  IV U60166 ( .A(n39568), .Z(n39569) );
  NOR U60167 ( .A(n39570), .B(n39569), .Z(n45076) );
  IV U60168 ( .A(n39571), .Z(n39573) );
  NOR U60169 ( .A(n39573), .B(n39572), .Z(n45073) );
  NOR U60170 ( .A(n45076), .B(n45073), .Z(n43062) );
  IV U60171 ( .A(n39574), .Z(n39575) );
  NOR U60172 ( .A(n39576), .B(n39575), .Z(n45078) );
  IV U60173 ( .A(n39577), .Z(n39579) );
  NOR U60174 ( .A(n39579), .B(n39578), .Z(n50087) );
  IV U60175 ( .A(n39580), .Z(n39581) );
  NOR U60176 ( .A(n39582), .B(n39581), .Z(n53216) );
  NOR U60177 ( .A(n50087), .B(n53216), .Z(n47883) );
  IV U60178 ( .A(n39583), .Z(n39584) );
  NOR U60179 ( .A(n39585), .B(n39584), .Z(n45081) );
  IV U60180 ( .A(n39586), .Z(n39587) );
  NOR U60181 ( .A(n39588), .B(n39587), .Z(n47884) );
  NOR U60182 ( .A(n45081), .B(n47884), .Z(n43061) );
  IV U60183 ( .A(n39589), .Z(n39591) );
  NOR U60184 ( .A(n39591), .B(n39590), .Z(n45083) );
  IV U60185 ( .A(n39592), .Z(n39593) );
  NOR U60186 ( .A(n39594), .B(n39593), .Z(n47867) );
  IV U60187 ( .A(n39595), .Z(n39596) );
  NOR U60188 ( .A(n39597), .B(n39596), .Z(n47874) );
  NOR U60189 ( .A(n47867), .B(n47874), .Z(n43053) );
  IV U60190 ( .A(n39598), .Z(n39599) );
  NOR U60191 ( .A(n39600), .B(n39599), .Z(n47865) );
  IV U60192 ( .A(n39601), .Z(n39603) );
  NOR U60193 ( .A(n39603), .B(n39602), .Z(n47855) );
  IV U60194 ( .A(n39604), .Z(n39606) );
  NOR U60195 ( .A(n39606), .B(n39605), .Z(n43039) );
  IV U60196 ( .A(n43039), .Z(n43032) );
  IV U60197 ( .A(n39607), .Z(n39608) );
  NOR U60198 ( .A(n39609), .B(n39608), .Z(n39610) );
  IV U60199 ( .A(n39610), .Z(n47848) );
  IV U60200 ( .A(n39611), .Z(n39613) );
  NOR U60201 ( .A(n39613), .B(n39612), .Z(n47837) );
  IV U60202 ( .A(n39614), .Z(n39615) );
  NOR U60203 ( .A(n39616), .B(n39615), .Z(n47844) );
  NOR U60204 ( .A(n47837), .B(n47844), .Z(n43030) );
  IV U60205 ( .A(n39617), .Z(n39618) );
  NOR U60206 ( .A(n39619), .B(n39618), .Z(n47819) );
  IV U60207 ( .A(n39620), .Z(n39622) );
  NOR U60208 ( .A(n39622), .B(n39621), .Z(n47839) );
  NOR U60209 ( .A(n47819), .B(n47839), .Z(n43029) );
  IV U60210 ( .A(n39623), .Z(n39625) );
  NOR U60211 ( .A(n39625), .B(n39624), .Z(n47817) );
  IV U60212 ( .A(n39626), .Z(n39627) );
  NOR U60213 ( .A(n39628), .B(n39627), .Z(n50108) );
  IV U60214 ( .A(n39629), .Z(n39631) );
  NOR U60215 ( .A(n39631), .B(n39630), .Z(n50104) );
  NOR U60216 ( .A(n50108), .B(n50104), .Z(n45088) );
  IV U60217 ( .A(n39632), .Z(n39633) );
  NOR U60218 ( .A(n39634), .B(n39633), .Z(n55318) );
  IV U60219 ( .A(n39635), .Z(n39637) );
  NOR U60220 ( .A(n39637), .B(n39636), .Z(n55310) );
  NOR U60221 ( .A(n55318), .B(n55310), .Z(n45089) );
  IV U60222 ( .A(n39638), .Z(n39639) );
  NOR U60223 ( .A(n39640), .B(n39639), .Z(n39641) );
  IV U60224 ( .A(n39641), .Z(n47805) );
  IV U60225 ( .A(n39642), .Z(n39643) );
  NOR U60226 ( .A(n39644), .B(n39643), .Z(n47797) );
  IV U60227 ( .A(n39645), .Z(n39646) );
  NOR U60228 ( .A(n39647), .B(n39646), .Z(n47795) );
  NOR U60229 ( .A(n47797), .B(n47795), .Z(n43007) );
  IV U60230 ( .A(n39648), .Z(n39650) );
  NOR U60231 ( .A(n39650), .B(n39649), .Z(n39651) );
  IV U60232 ( .A(n39651), .Z(n42996) );
  IV U60233 ( .A(n39652), .Z(n39654) );
  NOR U60234 ( .A(n39654), .B(n39653), .Z(n39655) );
  IV U60235 ( .A(n39655), .Z(n42981) );
  IV U60236 ( .A(n39656), .Z(n39658) );
  NOR U60237 ( .A(n39658), .B(n39657), .Z(n55337) );
  IV U60238 ( .A(n39659), .Z(n39660) );
  NOR U60239 ( .A(n39661), .B(n39660), .Z(n58317) );
  NOR U60240 ( .A(n55337), .B(n58317), .Z(n45113) );
  IV U60241 ( .A(n39662), .Z(n39663) );
  NOR U60242 ( .A(n39664), .B(n39663), .Z(n39665) );
  IV U60243 ( .A(n39665), .Z(n47775) );
  IV U60244 ( .A(n39666), .Z(n39667) );
  NOR U60245 ( .A(n39668), .B(n39667), .Z(n42963) );
  IV U60246 ( .A(n42963), .Z(n42955) );
  IV U60247 ( .A(n39669), .Z(n39670) );
  NOR U60248 ( .A(n39671), .B(n39670), .Z(n42952) );
  IV U60249 ( .A(n42952), .Z(n42945) );
  IV U60250 ( .A(n39672), .Z(n39674) );
  NOR U60251 ( .A(n39674), .B(n39673), .Z(n42949) );
  IV U60252 ( .A(n42949), .Z(n45119) );
  IV U60253 ( .A(n39675), .Z(n39677) );
  NOR U60254 ( .A(n39677), .B(n39676), .Z(n47739) );
  IV U60255 ( .A(n39678), .Z(n39679) );
  NOR U60256 ( .A(n39680), .B(n39679), .Z(n47733) );
  IV U60257 ( .A(n39681), .Z(n39682) );
  NOR U60258 ( .A(n39683), .B(n39682), .Z(n47727) );
  NOR U60259 ( .A(n47733), .B(n47727), .Z(n42885) );
  IV U60260 ( .A(n39684), .Z(n39686) );
  NOR U60261 ( .A(n39686), .B(n39685), .Z(n47716) );
  IV U60262 ( .A(n39687), .Z(n39688) );
  NOR U60263 ( .A(n39689), .B(n39688), .Z(n45141) );
  NOR U60264 ( .A(n47716), .B(n45141), .Z(n42877) );
  IV U60265 ( .A(n39690), .Z(n39691) );
  NOR U60266 ( .A(n39692), .B(n39691), .Z(n45153) );
  IV U60267 ( .A(n39693), .Z(n39694) );
  NOR U60268 ( .A(n39695), .B(n39694), .Z(n47710) );
  NOR U60269 ( .A(n45153), .B(n47710), .Z(n42857) );
  IV U60270 ( .A(n39696), .Z(n39698) );
  NOR U60271 ( .A(n39698), .B(n39697), .Z(n50193) );
  IV U60272 ( .A(n39699), .Z(n39701) );
  NOR U60273 ( .A(n39701), .B(n39700), .Z(n50186) );
  NOR U60274 ( .A(n50193), .B(n50186), .Z(n47690) );
  IV U60275 ( .A(n39702), .Z(n39704) );
  NOR U60276 ( .A(n39704), .B(n39703), .Z(n47651) );
  IV U60277 ( .A(n39705), .Z(n39706) );
  NOR U60278 ( .A(n39707), .B(n39706), .Z(n58231) );
  IV U60279 ( .A(n39708), .Z(n39710) );
  NOR U60280 ( .A(n39710), .B(n39709), .Z(n55442) );
  NOR U60281 ( .A(n58231), .B(n55442), .Z(n50221) );
  IV U60282 ( .A(n50221), .Z(n42809) );
  IV U60283 ( .A(n39711), .Z(n39713) );
  NOR U60284 ( .A(n39713), .B(n39712), .Z(n42800) );
  IV U60285 ( .A(n42800), .Z(n42795) );
  IV U60286 ( .A(n39714), .Z(n39715) );
  NOR U60287 ( .A(n39716), .B(n39715), .Z(n45161) );
  IV U60288 ( .A(n39717), .Z(n39718) );
  NOR U60289 ( .A(n39719), .B(n39718), .Z(n45168) );
  IV U60290 ( .A(n39720), .Z(n39722) );
  NOR U60291 ( .A(n39722), .B(n39721), .Z(n47636) );
  NOR U60292 ( .A(n45168), .B(n47636), .Z(n42785) );
  IV U60293 ( .A(n39723), .Z(n39725) );
  NOR U60294 ( .A(n39725), .B(n39724), .Z(n47592) );
  IV U60295 ( .A(n39726), .Z(n39728) );
  NOR U60296 ( .A(n39728), .B(n39727), .Z(n47566) );
  IV U60297 ( .A(n39729), .Z(n39731) );
  NOR U60298 ( .A(n39731), .B(n39730), .Z(n45175) );
  NOR U60299 ( .A(n47566), .B(n45175), .Z(n39732) );
  IV U60300 ( .A(n39732), .Z(n42760) );
  IV U60301 ( .A(n39733), .Z(n39734) );
  NOR U60302 ( .A(n39735), .B(n39734), .Z(n50264) );
  IV U60303 ( .A(n39736), .Z(n39738) );
  NOR U60304 ( .A(n39738), .B(n39737), .Z(n50259) );
  NOR U60305 ( .A(n50264), .B(n50259), .Z(n47561) );
  IV U60306 ( .A(n39739), .Z(n39741) );
  NOR U60307 ( .A(n39741), .B(n39740), .Z(n52984) );
  IV U60308 ( .A(n39742), .Z(n39743) );
  NOR U60309 ( .A(n39744), .B(n39743), .Z(n52993) );
  NOR U60310 ( .A(n52984), .B(n52993), .Z(n45178) );
  IV U60311 ( .A(n39745), .Z(n39746) );
  NOR U60312 ( .A(n39747), .B(n39746), .Z(n45184) );
  IV U60313 ( .A(n39748), .Z(n39750) );
  NOR U60314 ( .A(n39750), .B(n39749), .Z(n45179) );
  NOR U60315 ( .A(n45184), .B(n45179), .Z(n42752) );
  IV U60316 ( .A(n39751), .Z(n39753) );
  NOR U60317 ( .A(n39753), .B(n39752), .Z(n45182) );
  NOR U60318 ( .A(n39755), .B(n39754), .Z(n50283) );
  IV U60319 ( .A(n39756), .Z(n39758) );
  NOR U60320 ( .A(n39758), .B(n39757), .Z(n50279) );
  NOR U60321 ( .A(n50283), .B(n50279), .Z(n45187) );
  IV U60322 ( .A(n39759), .Z(n39760) );
  NOR U60323 ( .A(n39761), .B(n39760), .Z(n45193) );
  IV U60324 ( .A(n39762), .Z(n39763) );
  NOR U60325 ( .A(n39764), .B(n39763), .Z(n45188) );
  NOR U60326 ( .A(n45193), .B(n45188), .Z(n42750) );
  IV U60327 ( .A(n39765), .Z(n39766) );
  NOR U60328 ( .A(n39767), .B(n39766), .Z(n42746) );
  IV U60329 ( .A(n39768), .Z(n39769) );
  NOR U60330 ( .A(n39770), .B(n39769), .Z(n47550) );
  NOR U60331 ( .A(n39772), .B(n39771), .Z(n47546) );
  NOR U60332 ( .A(n47550), .B(n47546), .Z(n42745) );
  NOR U60333 ( .A(n39774), .B(n39773), .Z(n45214) );
  IV U60334 ( .A(n39775), .Z(n39776) );
  NOR U60335 ( .A(n39777), .B(n39776), .Z(n47535) );
  IV U60336 ( .A(n39778), .Z(n39780) );
  NOR U60337 ( .A(n39780), .B(n39779), .Z(n45217) );
  NOR U60338 ( .A(n47535), .B(n45217), .Z(n39781) );
  IV U60339 ( .A(n39781), .Z(n42711) );
  IV U60340 ( .A(n39782), .Z(n39783) );
  NOR U60341 ( .A(n39784), .B(n39783), .Z(n47533) );
  IV U60342 ( .A(n39785), .Z(n39787) );
  NOR U60343 ( .A(n39787), .B(n39786), .Z(n47525) );
  IV U60344 ( .A(n39788), .Z(n39789) );
  NOR U60345 ( .A(n39790), .B(n39789), .Z(n42688) );
  IV U60346 ( .A(n42688), .Z(n42680) );
  NOR U60347 ( .A(n39792), .B(n39791), .Z(n50356) );
  IV U60348 ( .A(n39793), .Z(n39795) );
  NOR U60349 ( .A(n39795), .B(n39794), .Z(n50351) );
  NOR U60350 ( .A(n50356), .B(n50351), .Z(n45238) );
  NOR U60351 ( .A(n39797), .B(n39796), .Z(n50370) );
  IV U60352 ( .A(n39798), .Z(n39799) );
  NOR U60353 ( .A(n39800), .B(n39799), .Z(n39801) );
  NOR U60354 ( .A(n50370), .B(n39801), .Z(n45241) );
  NOR U60355 ( .A(n39803), .B(n39802), .Z(n50389) );
  IV U60356 ( .A(n39804), .Z(n39806) );
  NOR U60357 ( .A(n39806), .B(n39805), .Z(n50384) );
  NOR U60358 ( .A(n50389), .B(n50384), .Z(n47508) );
  IV U60359 ( .A(n39807), .Z(n39808) );
  NOR U60360 ( .A(n39809), .B(n39808), .Z(n52945) );
  IV U60361 ( .A(n39810), .Z(n39811) );
  NOR U60362 ( .A(n39812), .B(n39811), .Z(n50392) );
  NOR U60363 ( .A(n52945), .B(n50392), .Z(n45244) );
  IV U60364 ( .A(n39813), .Z(n39814) );
  NOR U60365 ( .A(n39815), .B(n39814), .Z(n47490) );
  IV U60366 ( .A(n39816), .Z(n39818) );
  NOR U60367 ( .A(n39818), .B(n39817), .Z(n47492) );
  NOR U60368 ( .A(n47490), .B(n47492), .Z(n42646) );
  IV U60369 ( .A(n39819), .Z(n39820) );
  NOR U60370 ( .A(n39821), .B(n39820), .Z(n47465) );
  IV U60371 ( .A(n39822), .Z(n39823) );
  NOR U60372 ( .A(n39824), .B(n39823), .Z(n47457) );
  NOR U60373 ( .A(n47465), .B(n47457), .Z(n42632) );
  IV U60374 ( .A(n39825), .Z(n39827) );
  NOR U60375 ( .A(n39827), .B(n39826), .Z(n52913) );
  IV U60376 ( .A(n39828), .Z(n39829) );
  NOR U60377 ( .A(n39830), .B(n39829), .Z(n52920) );
  NOR U60378 ( .A(n52913), .B(n52920), .Z(n47450) );
  IV U60379 ( .A(n39831), .Z(n39832) );
  NOR U60380 ( .A(n39833), .B(n39832), .Z(n47442) );
  IV U60381 ( .A(n39834), .Z(n39836) );
  NOR U60382 ( .A(n39836), .B(n39835), .Z(n47451) );
  NOR U60383 ( .A(n47442), .B(n47451), .Z(n42630) );
  IV U60384 ( .A(n39837), .Z(n39838) );
  NOR U60385 ( .A(n39839), .B(n39838), .Z(n39840) );
  IV U60386 ( .A(n39840), .Z(n47446) );
  IV U60387 ( .A(n39841), .Z(n39842) );
  NOR U60388 ( .A(n39843), .B(n39842), .Z(n55580) );
  IV U60389 ( .A(n39844), .Z(n39846) );
  NOR U60390 ( .A(n39846), .B(n39845), .Z(n58070) );
  NOR U60391 ( .A(n55580), .B(n58070), .Z(n50412) );
  IV U60392 ( .A(n39847), .Z(n39848) );
  NOR U60393 ( .A(n39849), .B(n39848), .Z(n50417) );
  IV U60394 ( .A(n39850), .Z(n39851) );
  NOR U60395 ( .A(n39852), .B(n39851), .Z(n50413) );
  NOR U60396 ( .A(n50417), .B(n50413), .Z(n47433) );
  IV U60397 ( .A(n39853), .Z(n39854) );
  NOR U60398 ( .A(n39855), .B(n39854), .Z(n50436) );
  NOR U60399 ( .A(n39857), .B(n39856), .Z(n50430) );
  NOR U60400 ( .A(n50436), .B(n50430), .Z(n47420) );
  IV U60401 ( .A(n39858), .Z(n39859) );
  NOR U60402 ( .A(n39860), .B(n39859), .Z(n47408) );
  IV U60403 ( .A(n39861), .Z(n39863) );
  NOR U60404 ( .A(n39863), .B(n39862), .Z(n42584) );
  IV U60405 ( .A(n42584), .Z(n42574) );
  IV U60406 ( .A(n39864), .Z(n39866) );
  NOR U60407 ( .A(n39866), .B(n39865), .Z(n42571) );
  IV U60408 ( .A(n42571), .Z(n42562) );
  IV U60409 ( .A(n39867), .Z(n39868) );
  NOR U60410 ( .A(n39869), .B(n39868), .Z(n50468) );
  IV U60411 ( .A(n39870), .Z(n39871) );
  NOR U60412 ( .A(n39872), .B(n39871), .Z(n50463) );
  NOR U60413 ( .A(n50468), .B(n50463), .Z(n47399) );
  IV U60414 ( .A(n39873), .Z(n39874) );
  NOR U60415 ( .A(n39875), .B(n39874), .Z(n45278) );
  IV U60416 ( .A(n39876), .Z(n39877) );
  NOR U60417 ( .A(n39878), .B(n39877), .Z(n47382) );
  IV U60418 ( .A(n39879), .Z(n39881) );
  NOR U60419 ( .A(n39881), .B(n39880), .Z(n45280) );
  NOR U60420 ( .A(n47382), .B(n45280), .Z(n39882) );
  IV U60421 ( .A(n39882), .Z(n42533) );
  IV U60422 ( .A(n39883), .Z(n39884) );
  NOR U60423 ( .A(n39885), .B(n39884), .Z(n47378) );
  IV U60424 ( .A(n39886), .Z(n39887) );
  NOR U60425 ( .A(n39888), .B(n39887), .Z(n50499) );
  IV U60426 ( .A(n39889), .Z(n39890) );
  NOR U60427 ( .A(n39891), .B(n39890), .Z(n50495) );
  NOR U60428 ( .A(n50499), .B(n50495), .Z(n45286) );
  IV U60429 ( .A(n39892), .Z(n39893) );
  NOR U60430 ( .A(n39894), .B(n39893), .Z(n47356) );
  IV U60431 ( .A(n39895), .Z(n39897) );
  NOR U60432 ( .A(n39897), .B(n39896), .Z(n45309) );
  NOR U60433 ( .A(n47356), .B(n45309), .Z(n42492) );
  IV U60434 ( .A(n39898), .Z(n39900) );
  NOR U60435 ( .A(n39900), .B(n39899), .Z(n52808) );
  IV U60436 ( .A(n39901), .Z(n39903) );
  NOR U60437 ( .A(n39903), .B(n39902), .Z(n52818) );
  NOR U60438 ( .A(n52808), .B(n52818), .Z(n45313) );
  IV U60439 ( .A(n39904), .Z(n39906) );
  NOR U60440 ( .A(n39906), .B(n39905), .Z(n50534) );
  IV U60441 ( .A(n39907), .Z(n39909) );
  NOR U60442 ( .A(n39909), .B(n39908), .Z(n52813) );
  NOR U60443 ( .A(n50534), .B(n52813), .Z(n45312) );
  IV U60444 ( .A(n39910), .Z(n39911) );
  NOR U60445 ( .A(n39912), .B(n39911), .Z(n45320) );
  IV U60446 ( .A(n39913), .Z(n39915) );
  NOR U60447 ( .A(n39915), .B(n39914), .Z(n45315) );
  NOR U60448 ( .A(n45320), .B(n45315), .Z(n42485) );
  IV U60449 ( .A(n39916), .Z(n39918) );
  NOR U60450 ( .A(n39918), .B(n39917), .Z(n45318) );
  IV U60451 ( .A(n39919), .Z(n39921) );
  NOR U60452 ( .A(n39921), .B(n39920), .Z(n52802) );
  IV U60453 ( .A(n39922), .Z(n39923) );
  NOR U60454 ( .A(n39924), .B(n39923), .Z(n50549) );
  NOR U60455 ( .A(n52802), .B(n50549), .Z(n45323) );
  IV U60456 ( .A(n39925), .Z(n39927) );
  NOR U60457 ( .A(n39927), .B(n39926), .Z(n47339) );
  IV U60458 ( .A(n39928), .Z(n39929) );
  NOR U60459 ( .A(n39930), .B(n39929), .Z(n50571) );
  IV U60460 ( .A(n39931), .Z(n39932) );
  NOR U60461 ( .A(n39933), .B(n39932), .Z(n50566) );
  NOR U60462 ( .A(n50571), .B(n50566), .Z(n45339) );
  IV U60463 ( .A(n39934), .Z(n39935) );
  NOR U60464 ( .A(n39936), .B(n39935), .Z(n47319) );
  IV U60465 ( .A(n39937), .Z(n39938) );
  NOR U60466 ( .A(n39939), .B(n39938), .Z(n45340) );
  NOR U60467 ( .A(n47319), .B(n45340), .Z(n42455) );
  IV U60468 ( .A(n39940), .Z(n39941) );
  NOR U60469 ( .A(n39942), .B(n39941), .Z(n45347) );
  IV U60470 ( .A(n39943), .Z(n39944) );
  NOR U60471 ( .A(n39945), .B(n39944), .Z(n45345) );
  NOR U60472 ( .A(n45347), .B(n45345), .Z(n42447) );
  IV U60473 ( .A(n39946), .Z(n39947) );
  NOR U60474 ( .A(n39948), .B(n39947), .Z(n47308) );
  IV U60475 ( .A(n39949), .Z(n39950) );
  NOR U60476 ( .A(n39951), .B(n39950), .Z(n47305) );
  NOR U60477 ( .A(n47308), .B(n47305), .Z(n42446) );
  IV U60478 ( .A(n39952), .Z(n39953) );
  NOR U60479 ( .A(n39954), .B(n39953), .Z(n47298) );
  IV U60480 ( .A(n39955), .Z(n39957) );
  NOR U60481 ( .A(n39957), .B(n39956), .Z(n45350) );
  NOR U60482 ( .A(n47298), .B(n45350), .Z(n42445) );
  IV U60483 ( .A(n39958), .Z(n39960) );
  NOR U60484 ( .A(n39960), .B(n39959), .Z(n45356) );
  IV U60485 ( .A(n39961), .Z(n39963) );
  NOR U60486 ( .A(n39963), .B(n39962), .Z(n45353) );
  NOR U60487 ( .A(n45356), .B(n45353), .Z(n42444) );
  IV U60488 ( .A(n39964), .Z(n39965) );
  NOR U60489 ( .A(n39966), .B(n39965), .Z(n52756) );
  IV U60490 ( .A(n39967), .Z(n39968) );
  NOR U60491 ( .A(n39969), .B(n39968), .Z(n52762) );
  NOR U60492 ( .A(n52756), .B(n52762), .Z(n45360) );
  IV U60493 ( .A(n39970), .Z(n39972) );
  NOR U60494 ( .A(n39972), .B(n39971), .Z(n47273) );
  IV U60495 ( .A(n39973), .Z(n39974) );
  NOR U60496 ( .A(n39975), .B(n39974), .Z(n47274) );
  NOR U60497 ( .A(n47273), .B(n47274), .Z(n42429) );
  IV U60498 ( .A(n39976), .Z(n39977) );
  NOR U60499 ( .A(n39978), .B(n39977), .Z(n45371) );
  IV U60500 ( .A(n39979), .Z(n39980) );
  NOR U60501 ( .A(n39981), .B(n39980), .Z(n45369) );
  NOR U60502 ( .A(n45371), .B(n45369), .Z(n42428) );
  IV U60503 ( .A(n39982), .Z(n39983) );
  NOR U60504 ( .A(n39984), .B(n39983), .Z(n45386) );
  IV U60505 ( .A(n39985), .Z(n39987) );
  NOR U60506 ( .A(n39987), .B(n39986), .Z(n47258) );
  IV U60507 ( .A(n39988), .Z(n39989) );
  NOR U60508 ( .A(n39990), .B(n39989), .Z(n45389) );
  NOR U60509 ( .A(n47258), .B(n45389), .Z(n42399) );
  IV U60510 ( .A(n39991), .Z(n39993) );
  NOR U60511 ( .A(n39993), .B(n39992), .Z(n39994) );
  IV U60512 ( .A(n39994), .Z(n47255) );
  IV U60513 ( .A(n39995), .Z(n39996) );
  NOR U60514 ( .A(n39997), .B(n39996), .Z(n55788) );
  IV U60515 ( .A(n39998), .Z(n39999) );
  NOR U60516 ( .A(n40000), .B(n39999), .Z(n55781) );
  NOR U60517 ( .A(n55788), .B(n55781), .Z(n52717) );
  IV U60518 ( .A(n40001), .Z(n40003) );
  NOR U60519 ( .A(n40003), .B(n40002), .Z(n45405) );
  IV U60520 ( .A(n40004), .Z(n40006) );
  NOR U60521 ( .A(n40006), .B(n40005), .Z(n45402) );
  NOR U60522 ( .A(n45405), .B(n45402), .Z(n42384) );
  IV U60523 ( .A(n40007), .Z(n40008) );
  NOR U60524 ( .A(n40009), .B(n40008), .Z(n40010) );
  IV U60525 ( .A(n40010), .Z(n47247) );
  IV U60526 ( .A(n40011), .Z(n40012) );
  NOR U60527 ( .A(n40013), .B(n40012), .Z(n45411) );
  IV U60528 ( .A(n40014), .Z(n40015) );
  NOR U60529 ( .A(n40016), .B(n40015), .Z(n47242) );
  NOR U60530 ( .A(n45411), .B(n47242), .Z(n42377) );
  IV U60531 ( .A(n40017), .Z(n40018) );
  NOR U60532 ( .A(n40019), .B(n40018), .Z(n45416) );
  IV U60533 ( .A(n40020), .Z(n40022) );
  NOR U60534 ( .A(n40022), .B(n40021), .Z(n50629) );
  IV U60535 ( .A(n40023), .Z(n40024) );
  NOR U60536 ( .A(n40025), .B(n40024), .Z(n50625) );
  NOR U60537 ( .A(n50629), .B(n50625), .Z(n45415) );
  IV U60538 ( .A(n40026), .Z(n40028) );
  NOR U60539 ( .A(n40028), .B(n40027), .Z(n47236) );
  IV U60540 ( .A(n40029), .Z(n40030) );
  NOR U60541 ( .A(n40031), .B(n40030), .Z(n42357) );
  IV U60542 ( .A(n40032), .Z(n40034) );
  NOR U60543 ( .A(n40034), .B(n40033), .Z(n42353) );
  IV U60544 ( .A(n40035), .Z(n40036) );
  NOR U60545 ( .A(n40037), .B(n40036), .Z(n42347) );
  IV U60546 ( .A(n40038), .Z(n40040) );
  NOR U60547 ( .A(n40040), .B(n40039), .Z(n45424) );
  IV U60548 ( .A(n40041), .Z(n40043) );
  NOR U60549 ( .A(n40043), .B(n40042), .Z(n45426) );
  NOR U60550 ( .A(n45424), .B(n45426), .Z(n42346) );
  IV U60551 ( .A(n40044), .Z(n40045) );
  NOR U60552 ( .A(n40046), .B(n40045), .Z(n63046) );
  IV U60553 ( .A(n40047), .Z(n40048) );
  NOR U60554 ( .A(n40049), .B(n40048), .Z(n63060) );
  NOR U60555 ( .A(n63046), .B(n63060), .Z(n45429) );
  IV U60556 ( .A(n40050), .Z(n40051) );
  NOR U60557 ( .A(n40052), .B(n40051), .Z(n45451) );
  IV U60558 ( .A(n40053), .Z(n40055) );
  NOR U60559 ( .A(n40055), .B(n40054), .Z(n47193) );
  IV U60560 ( .A(n40056), .Z(n40057) );
  NOR U60561 ( .A(n40058), .B(n40057), .Z(n47179) );
  IV U60562 ( .A(n40059), .Z(n40061) );
  NOR U60563 ( .A(n40061), .B(n40060), .Z(n40062) );
  IV U60564 ( .A(n40062), .Z(n42270) );
  IV U60565 ( .A(n40063), .Z(n40065) );
  NOR U60566 ( .A(n40065), .B(n40064), .Z(n45470) );
  IV U60567 ( .A(n40066), .Z(n40068) );
  NOR U60568 ( .A(n40068), .B(n40067), .Z(n45483) );
  IV U60569 ( .A(n40069), .Z(n40071) );
  NOR U60570 ( .A(n40071), .B(n40070), .Z(n45494) );
  IV U60571 ( .A(n40072), .Z(n40073) );
  NOR U60572 ( .A(n40074), .B(n40073), .Z(n47162) );
  IV U60573 ( .A(n40075), .Z(n40077) );
  NOR U60574 ( .A(n40077), .B(n40076), .Z(n45497) );
  NOR U60575 ( .A(n47162), .B(n45497), .Z(n42239) );
  IV U60576 ( .A(n40078), .Z(n40080) );
  NOR U60577 ( .A(n40080), .B(n40079), .Z(n42237) );
  IV U60578 ( .A(n42237), .Z(n42232) );
  IV U60579 ( .A(n40081), .Z(n40083) );
  NOR U60580 ( .A(n40083), .B(n40082), .Z(n45503) );
  IV U60581 ( .A(n40086), .Z(n40084) );
  NOR U60582 ( .A(n40085), .B(n40084), .Z(n45513) );
  NOR U60583 ( .A(n45513), .B(n45507), .Z(n40089) );
  IV U60584 ( .A(n40085), .Z(n40087) );
  NOR U60585 ( .A(n40087), .B(n40086), .Z(n40088) );
  NOR U60586 ( .A(n40089), .B(n40088), .Z(n42230) );
  IV U60587 ( .A(n40090), .Z(n40092) );
  NOR U60588 ( .A(n40092), .B(n40091), .Z(n47156) );
  IV U60589 ( .A(n40093), .Z(n40094) );
  NOR U60590 ( .A(n40095), .B(n40094), .Z(n42227) );
  IV U60591 ( .A(n42227), .Z(n42221) );
  IV U60592 ( .A(n40096), .Z(n40098) );
  NOR U60593 ( .A(n40098), .B(n40097), .Z(n47152) );
  IV U60594 ( .A(n40099), .Z(n40100) );
  NOR U60595 ( .A(n40101), .B(n40100), .Z(n52596) );
  IV U60596 ( .A(n40102), .Z(n40103) );
  NOR U60597 ( .A(n40104), .B(n40103), .Z(n52603) );
  NOR U60598 ( .A(n52596), .B(n52603), .Z(n47144) );
  NOR U60599 ( .A(n40106), .B(n40105), .Z(n45520) );
  IV U60600 ( .A(n40107), .Z(n40108) );
  NOR U60601 ( .A(n40109), .B(n40108), .Z(n45518) );
  NOR U60602 ( .A(n45520), .B(n45518), .Z(n42212) );
  IV U60603 ( .A(n40110), .Z(n40111) );
  NOR U60604 ( .A(n40112), .B(n40111), .Z(n45527) );
  IV U60605 ( .A(n40113), .Z(n40115) );
  NOR U60606 ( .A(n40115), .B(n40114), .Z(n45523) );
  NOR U60607 ( .A(n45527), .B(n45523), .Z(n42211) );
  IV U60608 ( .A(n40116), .Z(n40117) );
  NOR U60609 ( .A(n40118), .B(n40117), .Z(n45529) );
  IV U60610 ( .A(n40119), .Z(n40121) );
  NOR U60611 ( .A(n40121), .B(n40120), .Z(n50756) );
  IV U60612 ( .A(n40122), .Z(n40124) );
  NOR U60613 ( .A(n40124), .B(n40123), .Z(n50752) );
  NOR U60614 ( .A(n50756), .B(n50752), .Z(n45535) );
  IV U60615 ( .A(n40125), .Z(n40126) );
  NOR U60616 ( .A(n40127), .B(n40126), .Z(n50763) );
  IV U60617 ( .A(n40128), .Z(n40129) );
  NOR U60618 ( .A(n40130), .B(n40129), .Z(n40131) );
  NOR U60619 ( .A(n50763), .B(n40131), .Z(n45541) );
  IV U60620 ( .A(n40132), .Z(n40134) );
  NOR U60621 ( .A(n40134), .B(n40133), .Z(n47134) );
  IV U60622 ( .A(n40135), .Z(n40137) );
  NOR U60623 ( .A(n40137), .B(n40136), .Z(n50790) );
  IV U60624 ( .A(n40138), .Z(n40140) );
  NOR U60625 ( .A(n40140), .B(n40139), .Z(n50785) );
  NOR U60626 ( .A(n50790), .B(n50785), .Z(n45547) );
  IV U60627 ( .A(n40141), .Z(n40142) );
  NOR U60628 ( .A(n40143), .B(n40142), .Z(n47126) );
  IV U60629 ( .A(n40144), .Z(n40145) );
  NOR U60630 ( .A(n40146), .B(n40145), .Z(n47120) );
  NOR U60631 ( .A(n47126), .B(n47120), .Z(n42174) );
  NOR U60632 ( .A(n40148), .B(n40147), .Z(n47106) );
  IV U60633 ( .A(n40149), .Z(n40150) );
  NOR U60634 ( .A(n40151), .B(n40150), .Z(n47110) );
  NOR U60635 ( .A(n47106), .B(n47110), .Z(n42173) );
  IV U60636 ( .A(n40152), .Z(n40154) );
  NOR U60637 ( .A(n40154), .B(n40153), .Z(n42171) );
  IV U60638 ( .A(n42171), .Z(n42160) );
  IV U60639 ( .A(n40155), .Z(n40157) );
  NOR U60640 ( .A(n40157), .B(n40156), .Z(n42157) );
  IV U60641 ( .A(n42157), .Z(n42152) );
  IV U60642 ( .A(n40158), .Z(n40159) );
  NOR U60643 ( .A(n40160), .B(n40159), .Z(n45557) );
  IV U60644 ( .A(n40161), .Z(n40162) );
  NOR U60645 ( .A(n40163), .B(n40162), .Z(n45565) );
  IV U60646 ( .A(n40164), .Z(n40166) );
  NOR U60647 ( .A(n40166), .B(n40165), .Z(n45563) );
  NOR U60648 ( .A(n45565), .B(n45563), .Z(n42150) );
  IV U60649 ( .A(n40167), .Z(n40169) );
  NOR U60650 ( .A(n40169), .B(n40168), .Z(n45571) );
  IV U60651 ( .A(n40170), .Z(n40171) );
  NOR U60652 ( .A(n40172), .B(n40171), .Z(n45568) );
  NOR U60653 ( .A(n45571), .B(n45568), .Z(n42149) );
  IV U60654 ( .A(n40173), .Z(n40175) );
  NOR U60655 ( .A(n40175), .B(n40174), .Z(n45573) );
  IV U60656 ( .A(n40176), .Z(n40178) );
  NOR U60657 ( .A(n40178), .B(n40177), .Z(n52547) );
  IV U60658 ( .A(n40179), .Z(n40180) );
  NOR U60659 ( .A(n40181), .B(n40180), .Z(n50816) );
  NOR U60660 ( .A(n52547), .B(n50816), .Z(n47098) );
  IV U60661 ( .A(n40182), .Z(n40183) );
  NOR U60662 ( .A(n40184), .B(n40183), .Z(n42140) );
  IV U60663 ( .A(n42140), .Z(n42130) );
  IV U60664 ( .A(n40185), .Z(n40187) );
  NOR U60665 ( .A(n40187), .B(n40186), .Z(n42127) );
  IV U60666 ( .A(n42127), .Z(n42117) );
  IV U60667 ( .A(n40188), .Z(n40189) );
  NOR U60668 ( .A(n40190), .B(n40189), .Z(n42112) );
  IV U60669 ( .A(n40191), .Z(n40193) );
  NOR U60670 ( .A(n40193), .B(n40192), .Z(n47088) );
  IV U60671 ( .A(n40194), .Z(n40196) );
  NOR U60672 ( .A(n40196), .B(n40195), .Z(n50847) );
  NOR U60673 ( .A(n40198), .B(n40197), .Z(n50841) );
  NOR U60674 ( .A(n50847), .B(n50841), .Z(n47087) );
  IV U60675 ( .A(n40199), .Z(n40200) );
  NOR U60676 ( .A(n40201), .B(n40200), .Z(n50852) );
  IV U60677 ( .A(n40202), .Z(n40203) );
  NOR U60678 ( .A(n40204), .B(n40203), .Z(n40205) );
  NOR U60679 ( .A(n50852), .B(n40205), .Z(n45592) );
  IV U60680 ( .A(n40206), .Z(n40208) );
  NOR U60681 ( .A(n40208), .B(n40207), .Z(n47077) );
  IV U60682 ( .A(n40209), .Z(n40211) );
  NOR U60683 ( .A(n40211), .B(n40210), .Z(n47065) );
  IV U60684 ( .A(n40212), .Z(n40213) );
  NOR U60685 ( .A(n40214), .B(n40213), .Z(n47045) );
  IV U60686 ( .A(n40215), .Z(n40217) );
  NOR U60687 ( .A(n40217), .B(n40216), .Z(n45603) );
  NOR U60688 ( .A(n47045), .B(n45603), .Z(n42067) );
  IV U60689 ( .A(n40218), .Z(n40220) );
  NOR U60690 ( .A(n40220), .B(n40219), .Z(n47040) );
  IV U60691 ( .A(n40221), .Z(n40222) );
  NOR U60692 ( .A(n40223), .B(n40222), .Z(n50874) );
  IV U60693 ( .A(n40224), .Z(n40225) );
  NOR U60694 ( .A(n40226), .B(n40225), .Z(n52505) );
  NOR U60695 ( .A(n50874), .B(n52505), .Z(n45613) );
  IV U60696 ( .A(n40227), .Z(n40229) );
  NOR U60697 ( .A(n40229), .B(n40228), .Z(n42057) );
  IV U60698 ( .A(n42057), .Z(n42051) );
  IV U60699 ( .A(n40230), .Z(n40231) );
  NOR U60700 ( .A(n40232), .B(n40231), .Z(n45615) );
  IV U60701 ( .A(n40233), .Z(n40235) );
  NOR U60702 ( .A(n40235), .B(n40234), .Z(n42041) );
  IV U60703 ( .A(n42041), .Z(n42031) );
  IV U60704 ( .A(n40236), .Z(n40237) );
  NOR U60705 ( .A(n40238), .B(n40237), .Z(n47027) );
  IV U60706 ( .A(n40239), .Z(n40240) );
  NOR U60707 ( .A(n40241), .B(n40240), .Z(n47025) );
  NOR U60708 ( .A(n47027), .B(n47025), .Z(n42029) );
  IV U60709 ( .A(n40242), .Z(n40243) );
  NOR U60710 ( .A(n40244), .B(n40243), .Z(n47015) );
  IV U60711 ( .A(n40245), .Z(n40246) );
  NOR U60712 ( .A(n40247), .B(n40246), .Z(n45634) );
  NOR U60713 ( .A(n47015), .B(n45634), .Z(n42014) );
  IV U60714 ( .A(n40248), .Z(n40250) );
  NOR U60715 ( .A(n40250), .B(n40249), .Z(n42010) );
  IV U60716 ( .A(n40251), .Z(n40253) );
  NOR U60717 ( .A(n40253), .B(n40252), .Z(n45640) );
  IV U60718 ( .A(n40254), .Z(n40255) );
  NOR U60719 ( .A(n40256), .B(n40255), .Z(n40257) );
  IV U60720 ( .A(n40257), .Z(n45648) );
  IV U60721 ( .A(n40258), .Z(n40260) );
  NOR U60722 ( .A(n40260), .B(n40259), .Z(n56104) );
  IV U60723 ( .A(n40261), .Z(n40262) );
  NOR U60724 ( .A(n40263), .B(n40262), .Z(n56096) );
  NOR U60725 ( .A(n56104), .B(n56096), .Z(n45653) );
  IV U60726 ( .A(n40264), .Z(n40266) );
  NOR U60727 ( .A(n40266), .B(n40265), .Z(n57649) );
  IV U60728 ( .A(n40267), .Z(n40269) );
  NOR U60729 ( .A(n40269), .B(n40268), .Z(n40270) );
  NOR U60730 ( .A(n57649), .B(n40270), .Z(n45664) );
  IV U60731 ( .A(n40271), .Z(n40272) );
  NOR U60732 ( .A(n40273), .B(n40272), .Z(n41938) );
  IV U60733 ( .A(n41938), .Z(n41933) );
  IV U60734 ( .A(n40274), .Z(n40276) );
  NOR U60735 ( .A(n40276), .B(n40275), .Z(n45681) );
  IV U60736 ( .A(n40277), .Z(n40278) );
  NOR U60737 ( .A(n40279), .B(n40278), .Z(n40280) );
  IV U60738 ( .A(n40280), .Z(n45698) );
  IV U60739 ( .A(n40281), .Z(n40283) );
  NOR U60740 ( .A(n40283), .B(n40282), .Z(n46972) );
  IV U60741 ( .A(n40284), .Z(n40285) );
  NOR U60742 ( .A(n40286), .B(n40285), .Z(n45700) );
  NOR U60743 ( .A(n46972), .B(n45700), .Z(n41909) );
  IV U60744 ( .A(n40287), .Z(n40289) );
  NOR U60745 ( .A(n40289), .B(n40288), .Z(n46965) );
  IV U60746 ( .A(n40290), .Z(n40292) );
  NOR U60747 ( .A(n40292), .B(n40291), .Z(n46960) );
  IV U60748 ( .A(n40293), .Z(n40295) );
  NOR U60749 ( .A(n40295), .B(n40294), .Z(n45705) );
  NOR U60750 ( .A(n46960), .B(n45705), .Z(n41900) );
  NOR U60751 ( .A(n57589), .B(n40296), .Z(n57579) );
  IV U60752 ( .A(n57589), .Z(n40297) );
  NOR U60753 ( .A(n40297), .B(n57588), .Z(n40298) );
  NOR U60754 ( .A(n40298), .B(n57591), .Z(n40299) );
  NOR U60755 ( .A(n57579), .B(n40299), .Z(n50990) );
  IV U60756 ( .A(n40300), .Z(n40302) );
  NOR U60757 ( .A(n40302), .B(n40301), .Z(n50996) );
  IV U60758 ( .A(n40303), .Z(n40304) );
  NOR U60759 ( .A(n40305), .B(n40304), .Z(n50991) );
  NOR U60760 ( .A(n50996), .B(n50991), .Z(n46954) );
  IV U60761 ( .A(n40306), .Z(n40307) );
  NOR U60762 ( .A(n40308), .B(n40307), .Z(n45708) );
  IV U60763 ( .A(n40309), .Z(n40311) );
  NOR U60764 ( .A(n40311), .B(n40310), .Z(n46950) );
  NOR U60765 ( .A(n45708), .B(n46950), .Z(n41893) );
  IV U60766 ( .A(n40312), .Z(n40314) );
  NOR U60767 ( .A(n40314), .B(n40313), .Z(n46930) );
  IV U60768 ( .A(n40315), .Z(n40317) );
  NOR U60769 ( .A(n40317), .B(n40316), .Z(n45714) );
  NOR U60770 ( .A(n46930), .B(n45714), .Z(n41872) );
  IV U60771 ( .A(n40318), .Z(n40320) );
  NOR U60772 ( .A(n40320), .B(n40319), .Z(n40321) );
  IV U60773 ( .A(n40321), .Z(n45726) );
  IV U60774 ( .A(n40322), .Z(n40324) );
  NOR U60775 ( .A(n40324), .B(n40323), .Z(n56196) );
  IV U60776 ( .A(n40325), .Z(n40326) );
  NOR U60777 ( .A(n40327), .B(n40326), .Z(n56190) );
  NOR U60778 ( .A(n56196), .B(n56190), .Z(n45724) );
  IV U60779 ( .A(n40328), .Z(n40330) );
  NOR U60780 ( .A(n40330), .B(n40329), .Z(n45727) );
  IV U60781 ( .A(n40331), .Z(n40332) );
  NOR U60782 ( .A(n40333), .B(n40332), .Z(n51011) );
  IV U60783 ( .A(n40334), .Z(n40335) );
  NOR U60784 ( .A(n40336), .B(n40335), .Z(n52390) );
  NOR U60785 ( .A(n51011), .B(n52390), .Z(n46915) );
  IV U60786 ( .A(n40337), .Z(n40339) );
  NOR U60787 ( .A(n40339), .B(n40338), .Z(n51020) );
  IV U60788 ( .A(n40340), .Z(n40341) );
  NOR U60789 ( .A(n40342), .B(n40341), .Z(n51016) );
  NOR U60790 ( .A(n51020), .B(n51016), .Z(n46913) );
  IV U60791 ( .A(n40343), .Z(n40344) );
  NOR U60792 ( .A(n40345), .B(n40344), .Z(n45733) );
  IV U60793 ( .A(n40346), .Z(n40347) );
  NOR U60794 ( .A(n40348), .B(n40347), .Z(n45731) );
  NOR U60795 ( .A(n45733), .B(n45731), .Z(n41851) );
  IV U60796 ( .A(n40349), .Z(n40350) );
  NOR U60797 ( .A(n40351), .B(n40350), .Z(n40352) );
  IV U60798 ( .A(n40352), .Z(n45740) );
  IV U60799 ( .A(n40353), .Z(n40355) );
  NOR U60800 ( .A(n40355), .B(n40354), .Z(n40356) );
  IV U60801 ( .A(n40356), .Z(n41840) );
  IV U60802 ( .A(n40357), .Z(n40358) );
  NOR U60803 ( .A(n40359), .B(n40358), .Z(n45741) );
  IV U60804 ( .A(n40360), .Z(n40361) );
  NOR U60805 ( .A(n40362), .B(n40361), .Z(n46872) );
  NOR U60806 ( .A(n45741), .B(n46872), .Z(n41827) );
  IV U60807 ( .A(n40363), .Z(n40365) );
  NOR U60808 ( .A(n40365), .B(n40364), .Z(n45745) );
  IV U60809 ( .A(n40366), .Z(n40368) );
  NOR U60810 ( .A(n40368), .B(n40367), .Z(n46877) );
  NOR U60811 ( .A(n45745), .B(n46877), .Z(n41825) );
  IV U60812 ( .A(n40369), .Z(n40370) );
  NOR U60813 ( .A(n40371), .B(n40370), .Z(n52376) );
  IV U60814 ( .A(n40372), .Z(n40373) );
  NOR U60815 ( .A(n40374), .B(n40373), .Z(n52381) );
  NOR U60816 ( .A(n52376), .B(n52381), .Z(n45744) );
  IV U60817 ( .A(n40375), .Z(n40376) );
  NOR U60818 ( .A(n40377), .B(n40376), .Z(n46850) );
  IV U60819 ( .A(n40378), .Z(n40379) );
  NOR U60820 ( .A(n40380), .B(n40379), .Z(n45751) );
  NOR U60821 ( .A(n46850), .B(n45751), .Z(n41817) );
  IV U60822 ( .A(n40381), .Z(n40383) );
  NOR U60823 ( .A(n40383), .B(n40382), .Z(n46861) );
  IV U60824 ( .A(n40384), .Z(n40386) );
  NOR U60825 ( .A(n40386), .B(n40385), .Z(n46854) );
  NOR U60826 ( .A(n46861), .B(n46854), .Z(n41816) );
  IV U60827 ( .A(n40387), .Z(n40388) );
  NOR U60828 ( .A(n40389), .B(n40388), .Z(n45757) );
  IV U60829 ( .A(n40390), .Z(n40391) );
  NOR U60830 ( .A(n40392), .B(n40391), .Z(n46845) );
  IV U60831 ( .A(n40393), .Z(n40394) );
  NOR U60832 ( .A(n40395), .B(n40394), .Z(n45760) );
  IV U60833 ( .A(n40396), .Z(n40398) );
  NOR U60834 ( .A(n40398), .B(n40397), .Z(n46840) );
  NOR U60835 ( .A(n45760), .B(n46840), .Z(n41808) );
  IV U60836 ( .A(n40399), .Z(n40401) );
  NOR U60837 ( .A(n40401), .B(n40400), .Z(n51068) );
  IV U60838 ( .A(n40402), .Z(n40403) );
  NOR U60839 ( .A(n40404), .B(n40403), .Z(n52353) );
  NOR U60840 ( .A(n51068), .B(n52353), .Z(n46835) );
  IV U60841 ( .A(n40405), .Z(n40406) );
  NOR U60842 ( .A(n40407), .B(n40406), .Z(n51073) );
  IV U60843 ( .A(n40408), .Z(n40409) );
  NOR U60844 ( .A(n40410), .B(n40409), .Z(n52345) );
  NOR U60845 ( .A(n51073), .B(n52345), .Z(n46833) );
  IV U60846 ( .A(n40414), .Z(n40411) );
  NOR U60847 ( .A(n40411), .B(n40412), .Z(n46820) );
  NOR U60848 ( .A(n46826), .B(n46820), .Z(n40416) );
  IV U60849 ( .A(n40412), .Z(n40413) );
  NOR U60850 ( .A(n40414), .B(n40413), .Z(n40415) );
  NOR U60851 ( .A(n40416), .B(n40415), .Z(n41800) );
  IV U60852 ( .A(n40417), .Z(n40419) );
  NOR U60853 ( .A(n40419), .B(n40418), .Z(n46812) );
  IV U60854 ( .A(n40420), .Z(n40422) );
  NOR U60855 ( .A(n40422), .B(n40421), .Z(n46807) );
  NOR U60856 ( .A(n46812), .B(n46807), .Z(n40423) );
  IV U60857 ( .A(n40423), .Z(n41799) );
  IV U60858 ( .A(n40424), .Z(n40425) );
  NOR U60859 ( .A(n40426), .B(n40425), .Z(n46796) );
  IV U60860 ( .A(n40427), .Z(n40428) );
  NOR U60861 ( .A(n40429), .B(n40428), .Z(n46801) );
  IV U60862 ( .A(n40430), .Z(n40432) );
  NOR U60863 ( .A(n40432), .B(n40431), .Z(n46799) );
  NOR U60864 ( .A(n46801), .B(n46799), .Z(n41797) );
  IV U60865 ( .A(n40433), .Z(n40434) );
  NOR U60866 ( .A(n40435), .B(n40434), .Z(n52334) );
  IV U60867 ( .A(n40436), .Z(n40438) );
  NOR U60868 ( .A(n40438), .B(n40437), .Z(n51089) );
  NOR U60869 ( .A(n52334), .B(n51089), .Z(n40439) );
  IV U60870 ( .A(n40439), .Z(n46792) );
  IV U60871 ( .A(n40440), .Z(n40441) );
  NOR U60872 ( .A(n40442), .B(n40441), .Z(n45785) );
  NOR U60873 ( .A(n40444), .B(n40443), .Z(n45783) );
  NOR U60874 ( .A(n45785), .B(n45783), .Z(n41776) );
  IV U60875 ( .A(n40445), .Z(n40447) );
  NOR U60876 ( .A(n40447), .B(n40446), .Z(n45798) );
  NOR U60877 ( .A(n40449), .B(n40448), .Z(n52318) );
  NOR U60878 ( .A(n45798), .B(n52318), .Z(n41768) );
  IV U60879 ( .A(n40450), .Z(n40452) );
  NOR U60880 ( .A(n40452), .B(n40451), .Z(n45801) );
  IV U60881 ( .A(n40453), .Z(n40454) );
  NOR U60882 ( .A(n40455), .B(n40454), .Z(n45796) );
  NOR U60883 ( .A(n45801), .B(n45796), .Z(n41767) );
  IV U60884 ( .A(n40456), .Z(n40458) );
  NOR U60885 ( .A(n40458), .B(n40457), .Z(n46772) );
  NOR U60886 ( .A(n40460), .B(n40459), .Z(n46782) );
  NOR U60887 ( .A(n46772), .B(n46782), .Z(n41766) );
  IV U60888 ( .A(n40461), .Z(n40463) );
  NOR U60889 ( .A(n40463), .B(n40462), .Z(n40464) );
  IV U60890 ( .A(n40464), .Z(n46777) );
  NOR U60891 ( .A(n40466), .B(n40465), .Z(n45808) );
  IV U60892 ( .A(n40467), .Z(n40469) );
  NOR U60893 ( .A(n40469), .B(n40468), .Z(n45804) );
  NOR U60894 ( .A(n45808), .B(n45804), .Z(n41760) );
  IV U60895 ( .A(n40470), .Z(n40472) );
  NOR U60896 ( .A(n40472), .B(n40471), .Z(n46759) );
  IV U60897 ( .A(n40473), .Z(n40474) );
  NOR U60898 ( .A(n40475), .B(n40474), .Z(n45812) );
  NOR U60899 ( .A(n46759), .B(n45812), .Z(n41753) );
  IV U60900 ( .A(n40476), .Z(n40477) );
  NOR U60901 ( .A(n40478), .B(n40477), .Z(n52280) );
  IV U60902 ( .A(n40479), .Z(n40480) );
  NOR U60903 ( .A(n40481), .B(n40480), .Z(n51126) );
  NOR U60904 ( .A(n52280), .B(n51126), .Z(n57429) );
  IV U60905 ( .A(n40482), .Z(n40484) );
  NOR U60906 ( .A(n40484), .B(n40483), .Z(n52269) );
  IV U60907 ( .A(n40485), .Z(n40487) );
  NOR U60908 ( .A(n40487), .B(n40486), .Z(n40488) );
  NOR U60909 ( .A(n52269), .B(n40488), .Z(n46742) );
  IV U60910 ( .A(n40489), .Z(n40491) );
  NOR U60911 ( .A(n40491), .B(n40490), .Z(n52271) );
  IV U60912 ( .A(n40492), .Z(n40493) );
  NOR U60913 ( .A(n40494), .B(n40493), .Z(n46746) );
  NOR U60914 ( .A(n52271), .B(n46746), .Z(n41735) );
  IV U60915 ( .A(n40495), .Z(n40497) );
  NOR U60916 ( .A(n40497), .B(n40496), .Z(n41711) );
  IV U60917 ( .A(n40498), .Z(n40499) );
  NOR U60918 ( .A(n40500), .B(n40499), .Z(n46727) );
  NOR U60919 ( .A(n41711), .B(n46727), .Z(n41697) );
  IV U60920 ( .A(n40501), .Z(n40502) );
  NOR U60921 ( .A(n40503), .B(n40502), .Z(n56367) );
  IV U60922 ( .A(n40504), .Z(n40505) );
  NOR U60923 ( .A(n40506), .B(n40505), .Z(n56356) );
  NOR U60924 ( .A(n56367), .B(n56356), .Z(n45830) );
  IV U60925 ( .A(n40507), .Z(n40509) );
  NOR U60926 ( .A(n40509), .B(n40508), .Z(n45834) );
  IV U60927 ( .A(n40510), .Z(n40512) );
  NOR U60928 ( .A(n40512), .B(n40511), .Z(n46717) );
  NOR U60929 ( .A(n45834), .B(n46717), .Z(n41696) );
  NOR U60930 ( .A(n40514), .B(n40513), .Z(n45859) );
  IV U60931 ( .A(n40515), .Z(n40516) );
  NOR U60932 ( .A(n40517), .B(n40516), .Z(n52212) );
  IV U60933 ( .A(n40518), .Z(n40520) );
  NOR U60934 ( .A(n40520), .B(n40519), .Z(n52220) );
  NOR U60935 ( .A(n52212), .B(n52220), .Z(n45858) );
  IV U60936 ( .A(n40521), .Z(n40522) );
  NOR U60937 ( .A(n40523), .B(n40522), .Z(n40524) );
  IV U60938 ( .A(n40524), .Z(n46688) );
  IV U60939 ( .A(n40525), .Z(n40527) );
  NOR U60940 ( .A(n40527), .B(n40526), .Z(n56413) );
  IV U60941 ( .A(n40528), .Z(n40529) );
  NOR U60942 ( .A(n40530), .B(n40529), .Z(n56405) );
  NOR U60943 ( .A(n56413), .B(n56405), .Z(n52206) );
  IV U60944 ( .A(n40531), .Z(n40532) );
  NOR U60945 ( .A(n40533), .B(n40532), .Z(n51208) );
  IV U60946 ( .A(n40534), .Z(n40536) );
  NOR U60947 ( .A(n40536), .B(n40535), .Z(n51202) );
  NOR U60948 ( .A(n51208), .B(n51202), .Z(n45864) );
  IV U60949 ( .A(n40537), .Z(n40539) );
  NOR U60950 ( .A(n40539), .B(n40538), .Z(n45867) );
  IV U60951 ( .A(n40540), .Z(n40541) );
  NOR U60952 ( .A(n40542), .B(n40541), .Z(n45871) );
  NOR U60953 ( .A(n45867), .B(n45871), .Z(n41634) );
  IV U60954 ( .A(n40543), .Z(n40544) );
  NOR U60955 ( .A(n40545), .B(n40544), .Z(n51225) );
  IV U60956 ( .A(n40546), .Z(n40548) );
  NOR U60957 ( .A(n40548), .B(n40547), .Z(n51220) );
  NOR U60958 ( .A(n51225), .B(n51220), .Z(n46681) );
  IV U60959 ( .A(n40549), .Z(n40551) );
  NOR U60960 ( .A(n40551), .B(n40550), .Z(n52199) );
  IV U60961 ( .A(n40552), .Z(n40553) );
  NOR U60962 ( .A(n40554), .B(n40553), .Z(n51228) );
  NOR U60963 ( .A(n52199), .B(n51228), .Z(n46680) );
  IV U60964 ( .A(n40555), .Z(n40557) );
  NOR U60965 ( .A(n40557), .B(n40556), .Z(n41612) );
  IV U60966 ( .A(n52159), .Z(n40558) );
  NOR U60967 ( .A(n40558), .B(n52158), .Z(n52171) );
  NOR U60968 ( .A(n52159), .B(n40559), .Z(n40560) );
  NOR U60969 ( .A(n40560), .B(n52161), .Z(n40561) );
  NOR U60970 ( .A(n52171), .B(n40561), .Z(n40562) );
  IV U60971 ( .A(n40562), .Z(n45902) );
  IV U60972 ( .A(n40563), .Z(n40564) );
  NOR U60973 ( .A(n40565), .B(n40564), .Z(n45905) );
  IV U60974 ( .A(n40566), .Z(n40568) );
  NOR U60975 ( .A(n40568), .B(n40567), .Z(n45912) );
  IV U60976 ( .A(n40569), .Z(n40570) );
  NOR U60977 ( .A(n40571), .B(n40570), .Z(n56493) );
  IV U60978 ( .A(n40572), .Z(n40573) );
  NOR U60979 ( .A(n40574), .B(n40573), .Z(n56485) );
  NOR U60980 ( .A(n56493), .B(n56485), .Z(n45917) );
  IV U60981 ( .A(n40575), .Z(n40577) );
  NOR U60982 ( .A(n40577), .B(n40576), .Z(n51283) );
  IV U60983 ( .A(n40578), .Z(n40580) );
  NOR U60984 ( .A(n40580), .B(n40579), .Z(n40581) );
  NOR U60985 ( .A(n51283), .B(n40581), .Z(n45919) );
  IV U60986 ( .A(n40582), .Z(n40583) );
  NOR U60987 ( .A(n40584), .B(n40583), .Z(n40585) );
  IV U60988 ( .A(n40585), .Z(n45926) );
  IV U60989 ( .A(n40586), .Z(n40588) );
  NOR U60990 ( .A(n40588), .B(n40587), .Z(n45931) );
  IV U60991 ( .A(n40589), .Z(n40590) );
  NOR U60992 ( .A(n40591), .B(n40590), .Z(n45928) );
  NOR U60993 ( .A(n45931), .B(n45928), .Z(n41549) );
  IV U60994 ( .A(n40592), .Z(n40594) );
  NOR U60995 ( .A(n40594), .B(n40593), .Z(n46634) );
  IV U60996 ( .A(n40595), .Z(n40597) );
  NOR U60997 ( .A(n40597), .B(n40596), .Z(n51302) );
  IV U60998 ( .A(n40598), .Z(n40599) );
  NOR U60999 ( .A(n40600), .B(n40599), .Z(n51298) );
  NOR U61000 ( .A(n51302), .B(n51298), .Z(n46626) );
  NOR U61001 ( .A(n40601), .B(n40602), .Z(n40606) );
  IV U61002 ( .A(n40602), .Z(n40603) );
  NOR U61003 ( .A(n40604), .B(n40603), .Z(n56539) );
  NOR U61004 ( .A(n56539), .B(n56527), .Z(n40605) );
  NOR U61005 ( .A(n40606), .B(n40605), .Z(n45933) );
  NOR U61006 ( .A(n40608), .B(n40607), .Z(n52123) );
  IV U61007 ( .A(n40609), .Z(n40611) );
  NOR U61008 ( .A(n40611), .B(n40610), .Z(n51331) );
  NOR U61009 ( .A(n52123), .B(n51331), .Z(n45935) );
  IV U61010 ( .A(n45935), .Z(n51320) );
  IV U61011 ( .A(n40612), .Z(n40613) );
  NOR U61012 ( .A(n40614), .B(n40613), .Z(n40615) );
  IV U61013 ( .A(n40615), .Z(n46599) );
  IV U61014 ( .A(n40616), .Z(n40617) );
  NOR U61015 ( .A(n40618), .B(n40617), .Z(n57290) );
  IV U61016 ( .A(n40619), .Z(n40621) );
  NOR U61017 ( .A(n40621), .B(n40620), .Z(n56571) );
  NOR U61018 ( .A(n57290), .B(n56571), .Z(n46606) );
  IV U61019 ( .A(n40622), .Z(n40623) );
  NOR U61020 ( .A(n40624), .B(n40623), .Z(n45939) );
  IV U61021 ( .A(n40625), .Z(n40627) );
  NOR U61022 ( .A(n40627), .B(n40626), .Z(n46594) );
  NOR U61023 ( .A(n45939), .B(n46594), .Z(n41516) );
  IV U61024 ( .A(n40628), .Z(n40629) );
  NOR U61025 ( .A(n40630), .B(n40629), .Z(n40631) );
  IV U61026 ( .A(n40631), .Z(n45944) );
  NOR U61027 ( .A(n40633), .B(n40632), .Z(n62315) );
  IV U61028 ( .A(n40634), .Z(n40636) );
  NOR U61029 ( .A(n40636), .B(n40635), .Z(n40637) );
  NOR U61030 ( .A(n62315), .B(n40637), .Z(n45942) );
  IV U61031 ( .A(n40638), .Z(n40639) );
  NOR U61032 ( .A(n40640), .B(n40639), .Z(n46574) );
  IV U61033 ( .A(n40641), .Z(n40642) );
  NOR U61034 ( .A(n40643), .B(n40642), .Z(n45946) );
  NOR U61035 ( .A(n46574), .B(n45946), .Z(n41515) );
  IV U61036 ( .A(n40644), .Z(n40646) );
  NOR U61037 ( .A(n40646), .B(n40645), .Z(n56602) );
  IV U61038 ( .A(n40647), .Z(n40649) );
  NOR U61039 ( .A(n40649), .B(n40648), .Z(n56592) );
  NOR U61040 ( .A(n56602), .B(n56592), .Z(n45951) );
  IV U61041 ( .A(n40650), .Z(n40652) );
  NOR U61042 ( .A(n40652), .B(n40651), .Z(n45957) );
  IV U61043 ( .A(n40653), .Z(n40655) );
  NOR U61044 ( .A(n40655), .B(n40654), .Z(n45954) );
  NOR U61045 ( .A(n45957), .B(n45954), .Z(n41502) );
  IV U61046 ( .A(n40656), .Z(n40658) );
  NOR U61047 ( .A(n40658), .B(n40657), .Z(n41484) );
  IV U61048 ( .A(n41484), .Z(n41474) );
  IV U61049 ( .A(n40659), .Z(n40661) );
  NOR U61050 ( .A(n40661), .B(n40660), .Z(n41471) );
  IV U61051 ( .A(n41471), .Z(n41467) );
  IV U61052 ( .A(n40662), .Z(n40664) );
  NOR U61053 ( .A(n40664), .B(n40663), .Z(n45964) );
  NOR U61054 ( .A(n40666), .B(n40665), .Z(n41457) );
  IV U61055 ( .A(n41457), .Z(n41452) );
  IV U61056 ( .A(n40667), .Z(n40668) );
  NOR U61057 ( .A(n40669), .B(n40668), .Z(n45977) );
  NOR U61058 ( .A(n40671), .B(n40670), .Z(n56647) );
  IV U61059 ( .A(n40672), .Z(n40674) );
  NOR U61060 ( .A(n40674), .B(n40673), .Z(n56639) );
  NOR U61061 ( .A(n56647), .B(n56639), .Z(n51367) );
  IV U61062 ( .A(n40675), .Z(n40677) );
  NOR U61063 ( .A(n40677), .B(n40676), .Z(n45982) );
  IV U61064 ( .A(n40678), .Z(n40679) );
  NOR U61065 ( .A(n40680), .B(n40679), .Z(n46560) );
  NOR U61066 ( .A(n45982), .B(n46560), .Z(n41450) );
  NOR U61067 ( .A(n40682), .B(n40681), .Z(n45995) );
  IV U61068 ( .A(n40683), .Z(n40685) );
  NOR U61069 ( .A(n40685), .B(n40684), .Z(n45991) );
  NOR U61070 ( .A(n45995), .B(n45991), .Z(n41437) );
  IV U61071 ( .A(n40686), .Z(n40687) );
  NOR U61072 ( .A(n40688), .B(n40687), .Z(n41435) );
  IV U61073 ( .A(n41435), .Z(n41428) );
  IV U61074 ( .A(n40689), .Z(n40691) );
  NOR U61075 ( .A(n40691), .B(n40690), .Z(n45998) );
  IV U61076 ( .A(n40692), .Z(n40694) );
  NOR U61077 ( .A(n40694), .B(n40693), .Z(n51395) );
  IV U61078 ( .A(n40695), .Z(n40696) );
  NOR U61079 ( .A(n40697), .B(n40696), .Z(n56670) );
  IV U61080 ( .A(n40698), .Z(n40699) );
  NOR U61081 ( .A(n40700), .B(n40699), .Z(n56662) );
  NOR U61082 ( .A(n56670), .B(n56662), .Z(n46009) );
  IV U61083 ( .A(n40701), .Z(n40702) );
  NOR U61084 ( .A(n40703), .B(n40702), .Z(n52027) );
  IV U61085 ( .A(n40704), .Z(n40705) );
  NOR U61086 ( .A(n40706), .B(n40705), .Z(n52018) );
  NOR U61087 ( .A(n52027), .B(n52018), .Z(n46551) );
  IV U61088 ( .A(n46551), .Z(n41412) );
  IV U61089 ( .A(n40707), .Z(n40708) );
  NOR U61090 ( .A(n40709), .B(n40708), .Z(n40710) );
  IV U61091 ( .A(n40710), .Z(n41401) );
  IV U61092 ( .A(n40711), .Z(n40713) );
  NOR U61093 ( .A(n40713), .B(n40712), .Z(n41392) );
  IV U61094 ( .A(n41392), .Z(n41381) );
  IV U61095 ( .A(n40714), .Z(n40715) );
  NOR U61096 ( .A(n40716), .B(n40715), .Z(n41376) );
  IV U61097 ( .A(n40717), .Z(n40718) );
  NOR U61098 ( .A(n40719), .B(n40718), .Z(n46527) );
  IV U61099 ( .A(n40720), .Z(n40721) );
  NOR U61100 ( .A(n40722), .B(n40721), .Z(n46019) );
  NOR U61101 ( .A(n46527), .B(n46019), .Z(n41375) );
  IV U61102 ( .A(n40723), .Z(n40724) );
  NOR U61103 ( .A(n40725), .B(n40724), .Z(n40726) );
  IV U61104 ( .A(n40726), .Z(n46022) );
  IV U61105 ( .A(n40727), .Z(n40729) );
  NOR U61106 ( .A(n40729), .B(n40728), .Z(n46519) );
  IV U61107 ( .A(n40730), .Z(n40731) );
  NOR U61108 ( .A(n40732), .B(n40731), .Z(n46025) );
  NOR U61109 ( .A(n46519), .B(n46025), .Z(n41366) );
  IV U61110 ( .A(n40733), .Z(n40735) );
  NOR U61111 ( .A(n40735), .B(n40734), .Z(n46028) );
  IV U61112 ( .A(n40736), .Z(n40737) );
  NOR U61113 ( .A(n40738), .B(n40737), .Z(n46036) );
  IV U61114 ( .A(n40739), .Z(n40740) );
  NOR U61115 ( .A(n40741), .B(n40740), .Z(n46034) );
  NOR U61116 ( .A(n46036), .B(n46034), .Z(n41358) );
  IV U61117 ( .A(n40742), .Z(n40744) );
  NOR U61118 ( .A(n40744), .B(n40743), .Z(n46040) );
  IV U61119 ( .A(n40745), .Z(n40747) );
  NOR U61120 ( .A(n40747), .B(n40746), .Z(n46503) );
  NOR U61121 ( .A(n46040), .B(n46503), .Z(n41357) );
  IV U61122 ( .A(n40748), .Z(n40749) );
  NOR U61123 ( .A(n40750), .B(n40749), .Z(n46493) );
  IV U61124 ( .A(n40751), .Z(n40752) );
  NOR U61125 ( .A(n40753), .B(n40752), .Z(n46487) );
  NOR U61126 ( .A(n46493), .B(n46487), .Z(n41356) );
  IV U61127 ( .A(n40754), .Z(n40756) );
  NOR U61128 ( .A(n40756), .B(n40755), .Z(n46491) );
  IV U61129 ( .A(n40757), .Z(n40759) );
  NOR U61130 ( .A(n40759), .B(n40758), .Z(n51453) );
  IV U61131 ( .A(n40760), .Z(n40761) );
  NOR U61132 ( .A(n40762), .B(n40761), .Z(n51448) );
  NOR U61133 ( .A(n51453), .B(n51448), .Z(n46486) );
  IV U61134 ( .A(n40763), .Z(n40765) );
  NOR U61135 ( .A(n40765), .B(n40764), .Z(n46478) );
  IV U61136 ( .A(n40766), .Z(n40767) );
  NOR U61137 ( .A(n40768), .B(n40767), .Z(n51976) );
  IV U61138 ( .A(n40769), .Z(n40770) );
  NOR U61139 ( .A(n40771), .B(n40770), .Z(n40772) );
  NOR U61140 ( .A(n51976), .B(n40772), .Z(n46477) );
  IV U61141 ( .A(n40773), .Z(n40774) );
  NOR U61142 ( .A(n40775), .B(n40774), .Z(n51468) );
  IV U61143 ( .A(n40776), .Z(n40777) );
  NOR U61144 ( .A(n40778), .B(n40777), .Z(n51463) );
  NOR U61145 ( .A(n51468), .B(n51463), .Z(n46473) );
  IV U61146 ( .A(n40779), .Z(n40781) );
  NOR U61147 ( .A(n40781), .B(n40780), .Z(n46045) );
  IV U61148 ( .A(n40782), .Z(n40784) );
  NOR U61149 ( .A(n40784), .B(n40783), .Z(n46047) );
  NOR U61150 ( .A(n46045), .B(n46047), .Z(n41343) );
  IV U61151 ( .A(n40785), .Z(n40787) );
  NOR U61152 ( .A(n40787), .B(n40786), .Z(n46050) );
  IV U61153 ( .A(n40788), .Z(n40789) );
  NOR U61154 ( .A(n40790), .B(n40789), .Z(n46043) );
  NOR U61155 ( .A(n46050), .B(n46043), .Z(n41342) );
  IV U61156 ( .A(n40791), .Z(n40792) );
  NOR U61157 ( .A(n40793), .B(n40792), .Z(n46055) );
  IV U61158 ( .A(n40794), .Z(n40795) );
  NOR U61159 ( .A(n40796), .B(n40795), .Z(n46053) );
  NOR U61160 ( .A(n46055), .B(n46053), .Z(n41341) );
  IV U61161 ( .A(n40797), .Z(n40799) );
  NOR U61162 ( .A(n40799), .B(n40798), .Z(n46458) );
  IV U61163 ( .A(n40800), .Z(n40802) );
  NOR U61164 ( .A(n40802), .B(n40801), .Z(n46452) );
  NOR U61165 ( .A(n46458), .B(n46452), .Z(n46060) );
  IV U61166 ( .A(n40803), .Z(n40804) );
  NOR U61167 ( .A(n40805), .B(n40804), .Z(n46064) );
  IV U61168 ( .A(n40806), .Z(n40808) );
  NOR U61169 ( .A(n40808), .B(n40807), .Z(n46061) );
  NOR U61170 ( .A(n46064), .B(n46061), .Z(n41340) );
  IV U61171 ( .A(n40809), .Z(n40811) );
  NOR U61172 ( .A(n40811), .B(n40810), .Z(n46445) );
  IV U61173 ( .A(n40812), .Z(n40813) );
  NOR U61174 ( .A(n40814), .B(n40813), .Z(n41323) );
  IV U61175 ( .A(n40815), .Z(n40817) );
  NOR U61176 ( .A(n40817), .B(n40816), .Z(n41319) );
  IV U61177 ( .A(n40818), .Z(n40819) );
  NOR U61178 ( .A(n40820), .B(n40819), .Z(n46431) );
  IV U61179 ( .A(n40821), .Z(n40822) );
  NOR U61180 ( .A(n40823), .B(n40822), .Z(n46433) );
  NOR U61181 ( .A(n46431), .B(n46433), .Z(n41316) );
  IV U61182 ( .A(n40824), .Z(n40825) );
  NOR U61183 ( .A(n40826), .B(n40825), .Z(n51508) );
  IV U61184 ( .A(n40827), .Z(n40829) );
  NOR U61185 ( .A(n40829), .B(n40828), .Z(n51499) );
  NOR U61186 ( .A(n51508), .B(n51499), .Z(n46075) );
  IV U61187 ( .A(n40830), .Z(n40831) );
  NOR U61188 ( .A(n40832), .B(n40831), .Z(n46410) );
  IV U61189 ( .A(n40833), .Z(n40834) );
  NOR U61190 ( .A(n40835), .B(n40834), .Z(n41287) );
  IV U61191 ( .A(n41287), .Z(n41282) );
  IV U61192 ( .A(n40836), .Z(n40838) );
  NOR U61193 ( .A(n40838), .B(n40837), .Z(n46076) );
  IV U61194 ( .A(n40839), .Z(n40840) );
  NOR U61195 ( .A(n40841), .B(n40840), .Z(n46082) );
  IV U61196 ( .A(n40842), .Z(n40844) );
  NOR U61197 ( .A(n40844), .B(n40843), .Z(n46381) );
  NOR U61198 ( .A(n46082), .B(n46381), .Z(n41280) );
  IV U61199 ( .A(n40845), .Z(n40846) );
  NOR U61200 ( .A(n40847), .B(n40846), .Z(n46389) );
  IV U61201 ( .A(n40848), .Z(n40850) );
  NOR U61202 ( .A(n40850), .B(n40849), .Z(n46384) );
  NOR U61203 ( .A(n46389), .B(n46384), .Z(n41279) );
  IV U61204 ( .A(n40851), .Z(n40853) );
  NOR U61205 ( .A(n40853), .B(n40852), .Z(n46387) );
  IV U61206 ( .A(n40854), .Z(n40855) );
  NOR U61207 ( .A(n40856), .B(n40855), .Z(n46089) );
  IV U61208 ( .A(n40857), .Z(n40859) );
  NOR U61209 ( .A(n40859), .B(n40858), .Z(n46087) );
  NOR U61210 ( .A(n46089), .B(n46087), .Z(n41271) );
  IV U61211 ( .A(n40860), .Z(n40862) );
  NOR U61212 ( .A(n40862), .B(n40861), .Z(n51532) );
  IV U61213 ( .A(n40863), .Z(n40865) );
  NOR U61214 ( .A(n40865), .B(n40864), .Z(n51527) );
  NOR U61215 ( .A(n51532), .B(n51527), .Z(n46374) );
  IV U61216 ( .A(n46374), .Z(n41270) );
  IV U61217 ( .A(n40866), .Z(n40867) );
  NOR U61218 ( .A(n40868), .B(n40867), .Z(n46369) );
  IV U61219 ( .A(n40869), .Z(n40870) );
  NOR U61220 ( .A(n40871), .B(n40870), .Z(n46375) );
  NOR U61221 ( .A(n46369), .B(n46375), .Z(n41269) );
  IV U61222 ( .A(n40872), .Z(n40874) );
  NOR U61223 ( .A(n40874), .B(n40873), .Z(n46371) );
  IV U61224 ( .A(n40875), .Z(n40876) );
  NOR U61225 ( .A(n40877), .B(n40876), .Z(n46093) );
  NOR U61226 ( .A(n46371), .B(n46093), .Z(n41268) );
  IV U61227 ( .A(n40878), .Z(n40880) );
  NOR U61228 ( .A(n40880), .B(n40879), .Z(n46355) );
  IV U61229 ( .A(n40881), .Z(n40883) );
  NOR U61230 ( .A(n40883), .B(n40882), .Z(n46353) );
  NOR U61231 ( .A(n46355), .B(n46353), .Z(n41260) );
  IV U61232 ( .A(n40884), .Z(n40886) );
  NOR U61233 ( .A(n40886), .B(n40885), .Z(n46343) );
  IV U61234 ( .A(n40887), .Z(n40888) );
  NOR U61235 ( .A(n40889), .B(n40888), .Z(n46348) );
  NOR U61236 ( .A(n46343), .B(n46348), .Z(n41259) );
  IV U61237 ( .A(n40890), .Z(n40891) );
  NOR U61238 ( .A(n40892), .B(n40891), .Z(n51842) );
  IV U61239 ( .A(n40893), .Z(n40895) );
  NOR U61240 ( .A(n40895), .B(n40894), .Z(n51837) );
  NOR U61241 ( .A(n51842), .B(n51837), .Z(n46326) );
  IV U61242 ( .A(n40896), .Z(n40897) );
  NOR U61243 ( .A(n40898), .B(n40897), .Z(n51835) );
  IV U61244 ( .A(n40899), .Z(n40901) );
  NOR U61245 ( .A(n40901), .B(n40900), .Z(n40902) );
  NOR U61246 ( .A(n51835), .B(n40902), .Z(n46100) );
  IV U61247 ( .A(n40903), .Z(n40905) );
  NOR U61248 ( .A(n40905), .B(n40904), .Z(n46106) );
  IV U61249 ( .A(n40906), .Z(n40907) );
  NOR U61250 ( .A(n40908), .B(n40907), .Z(n46104) );
  NOR U61251 ( .A(n46106), .B(n46104), .Z(n41231) );
  IV U61252 ( .A(n40909), .Z(n40910) );
  NOR U61253 ( .A(n40911), .B(n40910), .Z(n46113) );
  IV U61254 ( .A(n40912), .Z(n40914) );
  NOR U61255 ( .A(n40914), .B(n40913), .Z(n46110) );
  NOR U61256 ( .A(n46113), .B(n46110), .Z(n41229) );
  IV U61257 ( .A(n40915), .Z(n40916) );
  NOR U61258 ( .A(n40917), .B(n40916), .Z(n46314) );
  IV U61259 ( .A(n40918), .Z(n40919) );
  NOR U61260 ( .A(n40920), .B(n40919), .Z(n46287) );
  IV U61261 ( .A(n40921), .Z(n40922) );
  NOR U61262 ( .A(n40923), .B(n40922), .Z(n46274) );
  IV U61263 ( .A(n40924), .Z(n40925) );
  NOR U61264 ( .A(n40926), .B(n40925), .Z(n51764) );
  IV U61265 ( .A(n40927), .Z(n40929) );
  NOR U61266 ( .A(n40929), .B(n40928), .Z(n51614) );
  NOR U61267 ( .A(n51764), .B(n51614), .Z(n46262) );
  IV U61268 ( .A(n40930), .Z(n40931) );
  NOR U61269 ( .A(n40932), .B(n40931), .Z(n40933) );
  IV U61270 ( .A(n40933), .Z(n41164) );
  IV U61271 ( .A(n40934), .Z(n40936) );
  NOR U61272 ( .A(n40936), .B(n40935), .Z(n46131) );
  IV U61273 ( .A(n40937), .Z(n40938) );
  NOR U61274 ( .A(n40939), .B(n40938), .Z(n51618) );
  IV U61275 ( .A(n40940), .Z(n40942) );
  NOR U61276 ( .A(n40942), .B(n40941), .Z(n51760) );
  NOR U61277 ( .A(n51618), .B(n51760), .Z(n40943) );
  IV U61278 ( .A(n40943), .Z(n46135) );
  IV U61279 ( .A(n40944), .Z(n40945) );
  NOR U61280 ( .A(n40946), .B(n40945), .Z(n56888) );
  IV U61281 ( .A(n40947), .Z(n40949) );
  NOR U61282 ( .A(n40949), .B(n40948), .Z(n56879) );
  NOR U61283 ( .A(n56888), .B(n56879), .Z(n51755) );
  IV U61284 ( .A(n40950), .Z(n40951) );
  NOR U61285 ( .A(n40952), .B(n40951), .Z(n51628) );
  IV U61286 ( .A(n40953), .Z(n40954) );
  NOR U61287 ( .A(n40955), .B(n40954), .Z(n51623) );
  NOR U61288 ( .A(n51628), .B(n51623), .Z(n46138) );
  IV U61289 ( .A(n40956), .Z(n40958) );
  NOR U61290 ( .A(n40958), .B(n40957), .Z(n40959) );
  IV U61291 ( .A(n40959), .Z(n46251) );
  IV U61292 ( .A(n40960), .Z(n40961) );
  NOR U61293 ( .A(n40962), .B(n40961), .Z(n46148) );
  IV U61294 ( .A(n40963), .Z(n40965) );
  NOR U61295 ( .A(n40965), .B(n40964), .Z(n46243) );
  NOR U61296 ( .A(n46148), .B(n46243), .Z(n41141) );
  IV U61297 ( .A(n40966), .Z(n40968) );
  NOR U61298 ( .A(n40968), .B(n40967), .Z(n51735) );
  IV U61299 ( .A(n40969), .Z(n40970) );
  NOR U61300 ( .A(n40971), .B(n40970), .Z(n40972) );
  NOR U61301 ( .A(n51735), .B(n40972), .Z(n46233) );
  IV U61302 ( .A(n40973), .Z(n40974) );
  NOR U61303 ( .A(n40975), .B(n40974), .Z(n41139) );
  IV U61304 ( .A(n41139), .Z(n41129) );
  IV U61305 ( .A(n40976), .Z(n40978) );
  NOR U61306 ( .A(n40978), .B(n40977), .Z(n41126) );
  IV U61307 ( .A(n41126), .Z(n41116) );
  IV U61308 ( .A(n40979), .Z(n40980) );
  NOR U61309 ( .A(n40981), .B(n40980), .Z(n41113) );
  IV U61310 ( .A(n41113), .Z(n41108) );
  IV U61311 ( .A(n40982), .Z(n40983) );
  NOR U61312 ( .A(n40984), .B(n40983), .Z(n46226) );
  IV U61313 ( .A(n40985), .Z(n40987) );
  NOR U61314 ( .A(n40987), .B(n40986), .Z(n46152) );
  IV U61315 ( .A(n40988), .Z(n40990) );
  NOR U61316 ( .A(n40990), .B(n40989), .Z(n46224) );
  NOR U61317 ( .A(n46152), .B(n46224), .Z(n40991) );
  IV U61318 ( .A(n40991), .Z(n41106) );
  IV U61319 ( .A(n40992), .Z(n40993) );
  NOR U61320 ( .A(n40994), .B(n40993), .Z(n46159) );
  IV U61321 ( .A(n40995), .Z(n40997) );
  NOR U61322 ( .A(n40997), .B(n40996), .Z(n46154) );
  NOR U61323 ( .A(n46159), .B(n46154), .Z(n41105) );
  IV U61324 ( .A(n40998), .Z(n40999) );
  NOR U61325 ( .A(n41000), .B(n40999), .Z(n41103) );
  IV U61326 ( .A(n41103), .Z(n41093) );
  IV U61327 ( .A(n41001), .Z(n41002) );
  NOR U61328 ( .A(n41003), .B(n41002), .Z(n41090) );
  IV U61329 ( .A(n41090), .Z(n41079) );
  IV U61330 ( .A(n41004), .Z(n41005) );
  NOR U61331 ( .A(n41006), .B(n41005), .Z(n51673) );
  IV U61332 ( .A(n41007), .Z(n41008) );
  NOR U61333 ( .A(n41009), .B(n41008), .Z(n51680) );
  NOR U61334 ( .A(n51673), .B(n51680), .Z(n46169) );
  IV U61335 ( .A(n41010), .Z(n41011) );
  NOR U61336 ( .A(n41012), .B(n41011), .Z(n41069) );
  IV U61337 ( .A(n41069), .Z(n41063) );
  IV U61338 ( .A(n41013), .Z(n41014) );
  NOR U61339 ( .A(n41015), .B(n41014), .Z(n46207) );
  IV U61340 ( .A(n41016), .Z(n41017) );
  NOR U61341 ( .A(n41018), .B(n41017), .Z(n46196) );
  IV U61342 ( .A(n41019), .Z(n41020) );
  NOR U61343 ( .A(n41021), .B(n41020), .Z(n46212) );
  NOR U61344 ( .A(n46196), .B(n46212), .Z(n41061) );
  IV U61345 ( .A(n41022), .Z(n41023) );
  NOR U61346 ( .A(n41024), .B(n41023), .Z(n46173) );
  IV U61347 ( .A(n41025), .Z(n41026) );
  NOR U61348 ( .A(n41027), .B(n41026), .Z(n46199) );
  NOR U61349 ( .A(n46173), .B(n46199), .Z(n41060) );
  NOR U61350 ( .A(n41029), .B(n41028), .Z(n41033) );
  NOR U61351 ( .A(n41031), .B(n41030), .Z(n41032) );
  NOR U61352 ( .A(n41033), .B(n41032), .Z(n41034) );
  IV U61353 ( .A(n41034), .Z(n46185) );
  IV U61354 ( .A(n41035), .Z(n41037) );
  NOR U61355 ( .A(n41037), .B(n41036), .Z(n41046) );
  IV U61356 ( .A(n41038), .Z(n41040) );
  NOR U61357 ( .A(n41040), .B(n41039), .Z(n41041) );
  IV U61358 ( .A(n41041), .Z(n46179) );
  IV U61359 ( .A(n41042), .Z(n41043) );
  NOR U61360 ( .A(n41044), .B(n41043), .Z(n46178) );
  XOR U61361 ( .A(n46179), .B(n46178), .Z(n41045) );
  NOR U61362 ( .A(n41046), .B(n41045), .Z(n41052) );
  IV U61363 ( .A(n41046), .Z(n46177) );
  IV U61364 ( .A(n41047), .Z(n41049) );
  NOR U61365 ( .A(n41049), .B(n41048), .Z(n46175) );
  XOR U61366 ( .A(n46177), .B(n46175), .Z(n41050) );
  NOR U61367 ( .A(n46178), .B(n41050), .Z(n41051) );
  NOR U61368 ( .A(n41052), .B(n41051), .Z(n46187) );
  IV U61369 ( .A(n41053), .Z(n41055) );
  NOR U61370 ( .A(n41055), .B(n41054), .Z(n41059) );
  NOR U61371 ( .A(n41057), .B(n41056), .Z(n41058) );
  NOR U61372 ( .A(n41059), .B(n41058), .Z(n46188) );
  XOR U61373 ( .A(n46187), .B(n46188), .Z(n46184) );
  XOR U61374 ( .A(n46185), .B(n46184), .Z(n46201) );
  XOR U61375 ( .A(n41060), .B(n46201), .Z(n46195) );
  XOR U61376 ( .A(n41061), .B(n46195), .Z(n46208) );
  XOR U61377 ( .A(n46207), .B(n46208), .Z(n41062) );
  NOR U61378 ( .A(n41063), .B(n41062), .Z(n51670) );
  IV U61379 ( .A(n41064), .Z(n41065) );
  NOR U61380 ( .A(n41066), .B(n41065), .Z(n46171) );
  NOR U61381 ( .A(n46207), .B(n46171), .Z(n41067) );
  XOR U61382 ( .A(n41067), .B(n46208), .Z(n41068) );
  NOR U61383 ( .A(n41069), .B(n41068), .Z(n41070) );
  NOR U61384 ( .A(n51670), .B(n41070), .Z(n46168) );
  XOR U61385 ( .A(n46169), .B(n46168), .Z(n46166) );
  IV U61386 ( .A(n41071), .Z(n41073) );
  NOR U61387 ( .A(n41073), .B(n41072), .Z(n41080) );
  IV U61388 ( .A(n41074), .Z(n41075) );
  NOR U61389 ( .A(n41076), .B(n41075), .Z(n46164) );
  NOR U61390 ( .A(n41080), .B(n46164), .Z(n41077) );
  XOR U61391 ( .A(n46166), .B(n41077), .Z(n41087) );
  IV U61392 ( .A(n41087), .Z(n41078) );
  NOR U61393 ( .A(n41079), .B(n41078), .Z(n51660) );
  IV U61394 ( .A(n41080), .Z(n46167) );
  XOR U61395 ( .A(n46167), .B(n46166), .Z(n41081) );
  NOR U61396 ( .A(n46164), .B(n41081), .Z(n41086) );
  IV U61397 ( .A(n41082), .Z(n41083) );
  NOR U61398 ( .A(n41084), .B(n41083), .Z(n41088) );
  IV U61399 ( .A(n41088), .Z(n41085) );
  NOR U61400 ( .A(n41086), .B(n41085), .Z(n51657) );
  NOR U61401 ( .A(n41088), .B(n41087), .Z(n41089) );
  NOR U61402 ( .A(n51657), .B(n41089), .Z(n41099) );
  NOR U61403 ( .A(n41090), .B(n41099), .Z(n41091) );
  NOR U61404 ( .A(n51660), .B(n41091), .Z(n41097) );
  IV U61405 ( .A(n41097), .Z(n41092) );
  NOR U61406 ( .A(n41093), .B(n41092), .Z(n46163) );
  IV U61407 ( .A(n41094), .Z(n41095) );
  NOR U61408 ( .A(n41096), .B(n41095), .Z(n41098) );
  NOR U61409 ( .A(n41098), .B(n41097), .Z(n41102) );
  IV U61410 ( .A(n41098), .Z(n41101) );
  IV U61411 ( .A(n41099), .Z(n41100) );
  NOR U61412 ( .A(n41101), .B(n41100), .Z(n51655) );
  NOR U61413 ( .A(n41102), .B(n51655), .Z(n46160) );
  NOR U61414 ( .A(n41103), .B(n46160), .Z(n41104) );
  NOR U61415 ( .A(n46163), .B(n41104), .Z(n46155) );
  XOR U61416 ( .A(n41105), .B(n46155), .Z(n51719) );
  XOR U61417 ( .A(n41106), .B(n51719), .Z(n46227) );
  XOR U61418 ( .A(n46226), .B(n46227), .Z(n41107) );
  NOR U61419 ( .A(n41108), .B(n41107), .Z(n51723) );
  IV U61420 ( .A(n41109), .Z(n41110) );
  NOR U61421 ( .A(n41111), .B(n41110), .Z(n46150) );
  NOR U61422 ( .A(n46226), .B(n46150), .Z(n41112) );
  XOR U61423 ( .A(n41112), .B(n46227), .Z(n41120) );
  NOR U61424 ( .A(n41113), .B(n41120), .Z(n41114) );
  NOR U61425 ( .A(n51723), .B(n41114), .Z(n41123) );
  IV U61426 ( .A(n41123), .Z(n41115) );
  NOR U61427 ( .A(n41116), .B(n41115), .Z(n51642) );
  IV U61428 ( .A(n41117), .Z(n41119) );
  NOR U61429 ( .A(n41119), .B(n41118), .Z(n41124) );
  IV U61430 ( .A(n41124), .Z(n41122) );
  IV U61431 ( .A(n41120), .Z(n41121) );
  NOR U61432 ( .A(n41122), .B(n41121), .Z(n51645) );
  NOR U61433 ( .A(n41124), .B(n41123), .Z(n41125) );
  NOR U61434 ( .A(n51645), .B(n41125), .Z(n41133) );
  NOR U61435 ( .A(n41126), .B(n41133), .Z(n41127) );
  NOR U61436 ( .A(n51642), .B(n41127), .Z(n41136) );
  IV U61437 ( .A(n41136), .Z(n41128) );
  NOR U61438 ( .A(n41129), .B(n41128), .Z(n51731) );
  IV U61439 ( .A(n41130), .Z(n41131) );
  NOR U61440 ( .A(n41132), .B(n41131), .Z(n41137) );
  IV U61441 ( .A(n41137), .Z(n41135) );
  IV U61442 ( .A(n41133), .Z(n41134) );
  NOR U61443 ( .A(n41135), .B(n41134), .Z(n51728) );
  NOR U61444 ( .A(n41137), .B(n41136), .Z(n41138) );
  NOR U61445 ( .A(n51728), .B(n41138), .Z(n51736) );
  NOR U61446 ( .A(n41139), .B(n51736), .Z(n41140) );
  NOR U61447 ( .A(n51731), .B(n41140), .Z(n46231) );
  XOR U61448 ( .A(n46233), .B(n46231), .Z(n46244) );
  XOR U61449 ( .A(n41141), .B(n46244), .Z(n46239) );
  XOR U61450 ( .A(n46251), .B(n46239), .Z(n46257) );
  IV U61451 ( .A(n41142), .Z(n41144) );
  NOR U61452 ( .A(n41144), .B(n41143), .Z(n46238) );
  IV U61453 ( .A(n41145), .Z(n41146) );
  NOR U61454 ( .A(n41147), .B(n41146), .Z(n46256) );
  NOR U61455 ( .A(n46238), .B(n46256), .Z(n41148) );
  XOR U61456 ( .A(n46257), .B(n41148), .Z(n46139) );
  IV U61457 ( .A(n41149), .Z(n41150) );
  NOR U61458 ( .A(n41151), .B(n41150), .Z(n46140) );
  IV U61459 ( .A(n41152), .Z(n41154) );
  NOR U61460 ( .A(n41154), .B(n41153), .Z(n46142) );
  NOR U61461 ( .A(n46140), .B(n46142), .Z(n41155) );
  XOR U61462 ( .A(n46139), .B(n41155), .Z(n51624) );
  XOR U61463 ( .A(n46138), .B(n51624), .Z(n51749) );
  XOR U61464 ( .A(n51755), .B(n51749), .Z(n51619) );
  XOR U61465 ( .A(n46135), .B(n51619), .Z(n46133) );
  XOR U61466 ( .A(n46131), .B(n46133), .Z(n41156) );
  NOR U61467 ( .A(n41164), .B(n41156), .Z(n51771) );
  IV U61468 ( .A(n41157), .Z(n41158) );
  NOR U61469 ( .A(n41159), .B(n41158), .Z(n46125) );
  IV U61470 ( .A(n41160), .Z(n41161) );
  NOR U61471 ( .A(n41162), .B(n41161), .Z(n46129) );
  NOR U61472 ( .A(n46131), .B(n46129), .Z(n41163) );
  XOR U61473 ( .A(n46133), .B(n41163), .Z(n46126) );
  XOR U61474 ( .A(n46125), .B(n46126), .Z(n41166) );
  NOR U61475 ( .A(n46126), .B(n41164), .Z(n41165) );
  NOR U61476 ( .A(n41166), .B(n41165), .Z(n41167) );
  NOR U61477 ( .A(n51771), .B(n41167), .Z(n46261) );
  XOR U61478 ( .A(n46262), .B(n46261), .Z(n46270) );
  IV U61479 ( .A(n41168), .Z(n41170) );
  NOR U61480 ( .A(n41170), .B(n41169), .Z(n46263) );
  IV U61481 ( .A(n41171), .Z(n41172) );
  NOR U61482 ( .A(n41173), .B(n41172), .Z(n46269) );
  NOR U61483 ( .A(n46263), .B(n46269), .Z(n41174) );
  XOR U61484 ( .A(n46270), .B(n41174), .Z(n46267) );
  IV U61485 ( .A(n41175), .Z(n41176) );
  NOR U61486 ( .A(n41177), .B(n41176), .Z(n51787) );
  IV U61487 ( .A(n41178), .Z(n41180) );
  NOR U61488 ( .A(n41180), .B(n41179), .Z(n51795) );
  NOR U61489 ( .A(n51787), .B(n51795), .Z(n46268) );
  XOR U61490 ( .A(n46267), .B(n46268), .Z(n46277) );
  XOR U61491 ( .A(n46274), .B(n46277), .Z(n46284) );
  IV U61492 ( .A(n41181), .Z(n41182) );
  NOR U61493 ( .A(n41183), .B(n41182), .Z(n46276) );
  IV U61494 ( .A(n41184), .Z(n41185) );
  NOR U61495 ( .A(n41186), .B(n41185), .Z(n46283) );
  NOR U61496 ( .A(n46276), .B(n46283), .Z(n41187) );
  XOR U61497 ( .A(n46284), .B(n41187), .Z(n46280) );
  IV U61498 ( .A(n41188), .Z(n41190) );
  NOR U61499 ( .A(n41190), .B(n41189), .Z(n46281) );
  IV U61500 ( .A(n41191), .Z(n41193) );
  NOR U61501 ( .A(n41193), .B(n41192), .Z(n46290) );
  NOR U61502 ( .A(n46281), .B(n46290), .Z(n41194) );
  XOR U61503 ( .A(n46280), .B(n41194), .Z(n46288) );
  XOR U61504 ( .A(n46287), .B(n46288), .Z(n46122) );
  IV U61505 ( .A(n41195), .Z(n41197) );
  NOR U61506 ( .A(n41197), .B(n41196), .Z(n46121) );
  IV U61507 ( .A(n41198), .Z(n41200) );
  NOR U61508 ( .A(n41200), .B(n41199), .Z(n46119) );
  NOR U61509 ( .A(n46121), .B(n46119), .Z(n41201) );
  XOR U61510 ( .A(n46122), .B(n41201), .Z(n46299) );
  IV U61511 ( .A(n41202), .Z(n41203) );
  NOR U61512 ( .A(n41204), .B(n41203), .Z(n46300) );
  IV U61513 ( .A(n41205), .Z(n41206) );
  NOR U61514 ( .A(n41207), .B(n41206), .Z(n46304) );
  NOR U61515 ( .A(n46300), .B(n46304), .Z(n41208) );
  XOR U61516 ( .A(n46299), .B(n41208), .Z(n46296) );
  IV U61517 ( .A(n41209), .Z(n41211) );
  NOR U61518 ( .A(n41211), .B(n41210), .Z(n46295) );
  IV U61519 ( .A(n41212), .Z(n41214) );
  NOR U61520 ( .A(n41214), .B(n41213), .Z(n46117) );
  NOR U61521 ( .A(n46295), .B(n46117), .Z(n41215) );
  XOR U61522 ( .A(n46296), .B(n41215), .Z(n51577) );
  IV U61523 ( .A(n51577), .Z(n51590) );
  IV U61524 ( .A(n41216), .Z(n41217) );
  NOR U61525 ( .A(n41218), .B(n41217), .Z(n51593) );
  IV U61526 ( .A(n41219), .Z(n41220) );
  NOR U61527 ( .A(n41221), .B(n41220), .Z(n51589) );
  NOR U61528 ( .A(n51593), .B(n51589), .Z(n46116) );
  IV U61529 ( .A(n46116), .Z(n51576) );
  XOR U61530 ( .A(n51590), .B(n51576), .Z(n46312) );
  IV U61531 ( .A(n46312), .Z(n41228) );
  IV U61532 ( .A(n41222), .Z(n41223) );
  NOR U61533 ( .A(n41224), .B(n41223), .Z(n51586) );
  IV U61534 ( .A(n41225), .Z(n41227) );
  NOR U61535 ( .A(n41227), .B(n41226), .Z(n51575) );
  NOR U61536 ( .A(n51586), .B(n51575), .Z(n46313) );
  XOR U61537 ( .A(n41228), .B(n46313), .Z(n46315) );
  XOR U61538 ( .A(n46314), .B(n46315), .Z(n46111) );
  XOR U61539 ( .A(n41229), .B(n46111), .Z(n41230) );
  IV U61540 ( .A(n41230), .Z(n46108) );
  XOR U61541 ( .A(n41231), .B(n46108), .Z(n46322) );
  IV U61542 ( .A(n41232), .Z(n41234) );
  NOR U61543 ( .A(n41234), .B(n41233), .Z(n46101) );
  IV U61544 ( .A(n41235), .Z(n41237) );
  NOR U61545 ( .A(n41237), .B(n41236), .Z(n46321) );
  NOR U61546 ( .A(n46101), .B(n46321), .Z(n41238) );
  XOR U61547 ( .A(n46322), .B(n41238), .Z(n51826) );
  XOR U61548 ( .A(n46100), .B(n51826), .Z(n46328) );
  XOR U61549 ( .A(n46326), .B(n46328), .Z(n51557) );
  IV U61550 ( .A(n41239), .Z(n41241) );
  NOR U61551 ( .A(n41241), .B(n41240), .Z(n46325) );
  IV U61552 ( .A(n41242), .Z(n41244) );
  NOR U61553 ( .A(n41244), .B(n41243), .Z(n46339) );
  NOR U61554 ( .A(n46325), .B(n46339), .Z(n41245) );
  XOR U61555 ( .A(n51557), .B(n41245), .Z(n46333) );
  IV U61556 ( .A(n41246), .Z(n41248) );
  NOR U61557 ( .A(n41248), .B(n41247), .Z(n46336) );
  IV U61558 ( .A(n41249), .Z(n41251) );
  NOR U61559 ( .A(n41251), .B(n41250), .Z(n46334) );
  NOR U61560 ( .A(n46336), .B(n46334), .Z(n41252) );
  XOR U61561 ( .A(n46333), .B(n41252), .Z(n51861) );
  IV U61562 ( .A(n41253), .Z(n41254) );
  NOR U61563 ( .A(n41255), .B(n41254), .Z(n57062) );
  IV U61564 ( .A(n41256), .Z(n41257) );
  NOR U61565 ( .A(n41258), .B(n41257), .Z(n57070) );
  NOR U61566 ( .A(n57062), .B(n57070), .Z(n51863) );
  XOR U61567 ( .A(n51861), .B(n51863), .Z(n46344) );
  XOR U61568 ( .A(n41259), .B(n46344), .Z(n46357) );
  XOR U61569 ( .A(n41260), .B(n46357), .Z(n46098) );
  IV U61570 ( .A(n41261), .Z(n41262) );
  NOR U61571 ( .A(n41263), .B(n41262), .Z(n46097) );
  IV U61572 ( .A(n41264), .Z(n41265) );
  NOR U61573 ( .A(n41266), .B(n41265), .Z(n46361) );
  NOR U61574 ( .A(n46097), .B(n46361), .Z(n41267) );
  XOR U61575 ( .A(n46098), .B(n41267), .Z(n46370) );
  XOR U61576 ( .A(n41268), .B(n46370), .Z(n46376) );
  XOR U61577 ( .A(n41269), .B(n46376), .Z(n51529) );
  XOR U61578 ( .A(n41270), .B(n51529), .Z(n46090) );
  XOR U61579 ( .A(n41271), .B(n46090), .Z(n46085) );
  IV U61580 ( .A(n41272), .Z(n41274) );
  NOR U61581 ( .A(n41274), .B(n41273), .Z(n51893) );
  IV U61582 ( .A(n41275), .Z(n41276) );
  NOR U61583 ( .A(n41277), .B(n41276), .Z(n41278) );
  NOR U61584 ( .A(n51893), .B(n41278), .Z(n46086) );
  XOR U61585 ( .A(n46085), .B(n46086), .Z(n46390) );
  XOR U61586 ( .A(n46387), .B(n46390), .Z(n46385) );
  XOR U61587 ( .A(n41279), .B(n46385), .Z(n46081) );
  XOR U61588 ( .A(n41280), .B(n46081), .Z(n46079) );
  XOR U61589 ( .A(n46076), .B(n46079), .Z(n41281) );
  NOR U61590 ( .A(n41282), .B(n41281), .Z(n51908) );
  IV U61591 ( .A(n41283), .Z(n41284) );
  NOR U61592 ( .A(n41285), .B(n41284), .Z(n46078) );
  NOR U61593 ( .A(n46076), .B(n46078), .Z(n41286) );
  XOR U61594 ( .A(n41286), .B(n46079), .Z(n46402) );
  NOR U61595 ( .A(n41287), .B(n46402), .Z(n41288) );
  NOR U61596 ( .A(n51908), .B(n41288), .Z(n46406) );
  IV U61597 ( .A(n41289), .Z(n41290) );
  NOR U61598 ( .A(n41291), .B(n41290), .Z(n46401) );
  IV U61599 ( .A(n41292), .Z(n41293) );
  NOR U61600 ( .A(n41294), .B(n41293), .Z(n46405) );
  NOR U61601 ( .A(n46401), .B(n46405), .Z(n41295) );
  XOR U61602 ( .A(n46406), .B(n41295), .Z(n46414) );
  XOR U61603 ( .A(n46410), .B(n46414), .Z(n46421) );
  IV U61604 ( .A(n41296), .Z(n41297) );
  NOR U61605 ( .A(n41298), .B(n41297), .Z(n46412) );
  IV U61606 ( .A(n41299), .Z(n41301) );
  NOR U61607 ( .A(n41301), .B(n41300), .Z(n46420) );
  NOR U61608 ( .A(n46412), .B(n46420), .Z(n41302) );
  XOR U61609 ( .A(n46421), .B(n41302), .Z(n46417) );
  IV U61610 ( .A(n41303), .Z(n41304) );
  NOR U61611 ( .A(n41305), .B(n41304), .Z(n46418) );
  IV U61612 ( .A(n41306), .Z(n41307) );
  NOR U61613 ( .A(n41308), .B(n41307), .Z(n46424) );
  NOR U61614 ( .A(n46418), .B(n46424), .Z(n41309) );
  XOR U61615 ( .A(n46417), .B(n41309), .Z(n51501) );
  XOR U61616 ( .A(n46075), .B(n51501), .Z(n46429) );
  IV U61617 ( .A(n41310), .Z(n41311) );
  NOR U61618 ( .A(n41312), .B(n41311), .Z(n51496) );
  IV U61619 ( .A(n41313), .Z(n41315) );
  NOR U61620 ( .A(n41315), .B(n41314), .Z(n51492) );
  NOR U61621 ( .A(n51496), .B(n51492), .Z(n46430) );
  XOR U61622 ( .A(n46429), .B(n46430), .Z(n46434) );
  XOR U61623 ( .A(n41316), .B(n46434), .Z(n41320) );
  NOR U61624 ( .A(n41319), .B(n41320), .Z(n41317) );
  IV U61625 ( .A(n41317), .Z(n41318) );
  NOR U61626 ( .A(n41323), .B(n41318), .Z(n51946) );
  IV U61627 ( .A(n41319), .Z(n41322) );
  IV U61628 ( .A(n41320), .Z(n41321) );
  NOR U61629 ( .A(n41322), .B(n41321), .Z(n51939) );
  IV U61630 ( .A(n41323), .Z(n41325) );
  XOR U61631 ( .A(n46431), .B(n46434), .Z(n41324) );
  NOR U61632 ( .A(n41325), .B(n41324), .Z(n51485) );
  NOR U61633 ( .A(n51939), .B(n51485), .Z(n46440) );
  IV U61634 ( .A(n46440), .Z(n51942) );
  NOR U61635 ( .A(n51946), .B(n51942), .Z(n46068) );
  IV U61636 ( .A(n41326), .Z(n41327) );
  NOR U61637 ( .A(n41328), .B(n41327), .Z(n51941) );
  IV U61638 ( .A(n41329), .Z(n41330) );
  NOR U61639 ( .A(n41331), .B(n41330), .Z(n51949) );
  NOR U61640 ( .A(n51941), .B(n51949), .Z(n46070) );
  XOR U61641 ( .A(n46068), .B(n46070), .Z(n46072) );
  IV U61642 ( .A(n46072), .Z(n41339) );
  IV U61643 ( .A(n41332), .Z(n41333) );
  NOR U61644 ( .A(n41334), .B(n41333), .Z(n46071) );
  IV U61645 ( .A(n41335), .Z(n41337) );
  NOR U61646 ( .A(n41337), .B(n41336), .Z(n46066) );
  NOR U61647 ( .A(n46071), .B(n46066), .Z(n41338) );
  XOR U61648 ( .A(n41339), .B(n41338), .Z(n46447) );
  XOR U61649 ( .A(n46445), .B(n46447), .Z(n46062) );
  XOR U61650 ( .A(n41340), .B(n46062), .Z(n46059) );
  XOR U61651 ( .A(n46060), .B(n46059), .Z(n46056) );
  XOR U61652 ( .A(n41341), .B(n46056), .Z(n46042) );
  XOR U61653 ( .A(n41342), .B(n46042), .Z(n46048) );
  XOR U61654 ( .A(n41343), .B(n46048), .Z(n46471) );
  IV U61655 ( .A(n41344), .Z(n41346) );
  NOR U61656 ( .A(n41346), .B(n41345), .Z(n56737) );
  IV U61657 ( .A(n41347), .Z(n41348) );
  NOR U61658 ( .A(n41349), .B(n41348), .Z(n57154) );
  NOR U61659 ( .A(n56737), .B(n57154), .Z(n46472) );
  XOR U61660 ( .A(n46471), .B(n46472), .Z(n51465) );
  XOR U61661 ( .A(n46473), .B(n51465), .Z(n46476) );
  XOR U61662 ( .A(n46477), .B(n46476), .Z(n46479) );
  XOR U61663 ( .A(n46478), .B(n46479), .Z(n51450) );
  XOR U61664 ( .A(n46486), .B(n51450), .Z(n46482) );
  IV U61665 ( .A(n41350), .Z(n41352) );
  NOR U61666 ( .A(n41352), .B(n41351), .Z(n51981) );
  IV U61667 ( .A(n41353), .Z(n41355) );
  NOR U61668 ( .A(n41355), .B(n41354), .Z(n51989) );
  NOR U61669 ( .A(n51981), .B(n51989), .Z(n46483) );
  XOR U61670 ( .A(n46482), .B(n46483), .Z(n46494) );
  XOR U61671 ( .A(n46491), .B(n46494), .Z(n46488) );
  XOR U61672 ( .A(n41356), .B(n46488), .Z(n46039) );
  XOR U61673 ( .A(n41357), .B(n46039), .Z(n46037) );
  XOR U61674 ( .A(n41358), .B(n46037), .Z(n46509) );
  IV U61675 ( .A(n41359), .Z(n41360) );
  NOR U61676 ( .A(n41361), .B(n41360), .Z(n46030) );
  IV U61677 ( .A(n41362), .Z(n41364) );
  NOR U61678 ( .A(n41364), .B(n41363), .Z(n46508) );
  NOR U61679 ( .A(n46030), .B(n46508), .Z(n41365) );
  XOR U61680 ( .A(n46509), .B(n41365), .Z(n46521) );
  XOR U61681 ( .A(n46028), .B(n46521), .Z(n46026) );
  XOR U61682 ( .A(n41366), .B(n46026), .Z(n46021) );
  XOR U61683 ( .A(n46022), .B(n46021), .Z(n46023) );
  IV U61684 ( .A(n46023), .Z(n41374) );
  IV U61685 ( .A(n41367), .Z(n41369) );
  NOR U61686 ( .A(n41369), .B(n41368), .Z(n51419) );
  IV U61687 ( .A(n41370), .Z(n41371) );
  NOR U61688 ( .A(n41372), .B(n41371), .Z(n41373) );
  NOR U61689 ( .A(n51419), .B(n41373), .Z(n46024) );
  XOR U61690 ( .A(n41374), .B(n46024), .Z(n46528) );
  XOR U61691 ( .A(n41375), .B(n46528), .Z(n41385) );
  NOR U61692 ( .A(n41376), .B(n41385), .Z(n41379) );
  IV U61693 ( .A(n41376), .Z(n41378) );
  XOR U61694 ( .A(n46527), .B(n46528), .Z(n41377) );
  NOR U61695 ( .A(n41378), .B(n41377), .Z(n46526) );
  NOR U61696 ( .A(n41379), .B(n46526), .Z(n41388) );
  IV U61697 ( .A(n41388), .Z(n41380) );
  NOR U61698 ( .A(n41381), .B(n41380), .Z(n56684) );
  IV U61699 ( .A(n41382), .Z(n41383) );
  NOR U61700 ( .A(n41384), .B(n41383), .Z(n41389) );
  IV U61701 ( .A(n41389), .Z(n41387) );
  IV U61702 ( .A(n41385), .Z(n41386) );
  NOR U61703 ( .A(n41387), .B(n41386), .Z(n46533) );
  NOR U61704 ( .A(n41389), .B(n41388), .Z(n41390) );
  NOR U61705 ( .A(n46533), .B(n41390), .Z(n41391) );
  NOR U61706 ( .A(n41392), .B(n41391), .Z(n41393) );
  NOR U61707 ( .A(n56684), .B(n41393), .Z(n41394) );
  IV U61708 ( .A(n41394), .Z(n46537) );
  NOR U61709 ( .A(n41401), .B(n46537), .Z(n46541) );
  IV U61710 ( .A(n41395), .Z(n41396) );
  NOR U61711 ( .A(n41397), .B(n41396), .Z(n46016) );
  IV U61712 ( .A(n41398), .Z(n41400) );
  NOR U61713 ( .A(n41400), .B(n41399), .Z(n46536) );
  XOR U61714 ( .A(n46536), .B(n46537), .Z(n46017) );
  IV U61715 ( .A(n46017), .Z(n41402) );
  XOR U61716 ( .A(n46016), .B(n41402), .Z(n41404) );
  NOR U61717 ( .A(n41402), .B(n41401), .Z(n41403) );
  NOR U61718 ( .A(n41404), .B(n41403), .Z(n41405) );
  NOR U61719 ( .A(n46541), .B(n41405), .Z(n46544) );
  IV U61720 ( .A(n41406), .Z(n41408) );
  NOR U61721 ( .A(n41408), .B(n41407), .Z(n52007) );
  IV U61722 ( .A(n41409), .Z(n41411) );
  NOR U61723 ( .A(n41411), .B(n41410), .Z(n51405) );
  NOR U61724 ( .A(n52007), .B(n51405), .Z(n46545) );
  XOR U61725 ( .A(n46544), .B(n46545), .Z(n52024) );
  XOR U61726 ( .A(n41412), .B(n52024), .Z(n46553) );
  IV U61727 ( .A(n41413), .Z(n41415) );
  NOR U61728 ( .A(n41415), .B(n41414), .Z(n46552) );
  IV U61729 ( .A(n41416), .Z(n41417) );
  NOR U61730 ( .A(n41418), .B(n41417), .Z(n46014) );
  NOR U61731 ( .A(n46552), .B(n46014), .Z(n41419) );
  XOR U61732 ( .A(n46553), .B(n41419), .Z(n46008) );
  XOR U61733 ( .A(n46009), .B(n46008), .Z(n51396) );
  XOR U61734 ( .A(n51395), .B(n51396), .Z(n46001) );
  IV U61735 ( .A(n41420), .Z(n41421) );
  NOR U61736 ( .A(n41422), .B(n41421), .Z(n46011) );
  IV U61737 ( .A(n41423), .Z(n41425) );
  NOR U61738 ( .A(n41425), .B(n41424), .Z(n46000) );
  NOR U61739 ( .A(n46011), .B(n46000), .Z(n41426) );
  XOR U61740 ( .A(n46001), .B(n41426), .Z(n41433) );
  IV U61741 ( .A(n41433), .Z(n46005) );
  XOR U61742 ( .A(n45998), .B(n46005), .Z(n41427) );
  NOR U61743 ( .A(n41428), .B(n41427), .Z(n51384) );
  IV U61744 ( .A(n41429), .Z(n41430) );
  NOR U61745 ( .A(n41431), .B(n41430), .Z(n46003) );
  NOR U61746 ( .A(n45998), .B(n46003), .Z(n41432) );
  XOR U61747 ( .A(n41433), .B(n41432), .Z(n45996) );
  IV U61748 ( .A(n45996), .Z(n41434) );
  NOR U61749 ( .A(n41435), .B(n41434), .Z(n41436) );
  NOR U61750 ( .A(n51384), .B(n41436), .Z(n45992) );
  XOR U61751 ( .A(n41437), .B(n45992), .Z(n51381) );
  IV U61752 ( .A(n41438), .Z(n41440) );
  NOR U61753 ( .A(n41440), .B(n41439), .Z(n52052) );
  IV U61754 ( .A(n41441), .Z(n41442) );
  NOR U61755 ( .A(n41443), .B(n41442), .Z(n51380) );
  NOR U61756 ( .A(n52052), .B(n51380), .Z(n45987) );
  XOR U61757 ( .A(n51381), .B(n45987), .Z(n45984) );
  NOR U61758 ( .A(n41445), .B(n41444), .Z(n45983) );
  IV U61759 ( .A(n41446), .Z(n41448) );
  NOR U61760 ( .A(n41448), .B(n41447), .Z(n45980) );
  NOR U61761 ( .A(n45983), .B(n45980), .Z(n41449) );
  XOR U61762 ( .A(n45984), .B(n41449), .Z(n46561) );
  XOR U61763 ( .A(n41450), .B(n46561), .Z(n46563) );
  XOR U61764 ( .A(n51367), .B(n46563), .Z(n45978) );
  XOR U61765 ( .A(n45977), .B(n45978), .Z(n41451) );
  NOR U61766 ( .A(n41452), .B(n41451), .Z(n56636) );
  IV U61767 ( .A(n41453), .Z(n41455) );
  NOR U61768 ( .A(n41455), .B(n41454), .Z(n45975) );
  NOR U61769 ( .A(n45977), .B(n45975), .Z(n41456) );
  XOR U61770 ( .A(n41456), .B(n45978), .Z(n45972) );
  NOR U61771 ( .A(n41457), .B(n45972), .Z(n41458) );
  NOR U61772 ( .A(n56636), .B(n41458), .Z(n45968) );
  IV U61773 ( .A(n41459), .Z(n41460) );
  NOR U61774 ( .A(n41461), .B(n41460), .Z(n45971) );
  IV U61775 ( .A(n41462), .Z(n41464) );
  NOR U61776 ( .A(n41464), .B(n41463), .Z(n45967) );
  NOR U61777 ( .A(n45971), .B(n45967), .Z(n41465) );
  XOR U61778 ( .A(n45968), .B(n41465), .Z(n45966) );
  XOR U61779 ( .A(n45964), .B(n45966), .Z(n41466) );
  NOR U61780 ( .A(n41467), .B(n41466), .Z(n52070) );
  NOR U61781 ( .A(n41469), .B(n41468), .Z(n45961) );
  NOR U61782 ( .A(n45964), .B(n45961), .Z(n41470) );
  XOR U61783 ( .A(n45966), .B(n41470), .Z(n41478) );
  NOR U61784 ( .A(n41471), .B(n41478), .Z(n41472) );
  NOR U61785 ( .A(n52070), .B(n41472), .Z(n41481) );
  IV U61786 ( .A(n41481), .Z(n41473) );
  NOR U61787 ( .A(n41474), .B(n41473), .Z(n51350) );
  IV U61788 ( .A(n41475), .Z(n41476) );
  NOR U61789 ( .A(n41477), .B(n41476), .Z(n41482) );
  IV U61790 ( .A(n41482), .Z(n41480) );
  IV U61791 ( .A(n41478), .Z(n41479) );
  NOR U61792 ( .A(n41480), .B(n41479), .Z(n51352) );
  NOR U61793 ( .A(n41482), .B(n41481), .Z(n41483) );
  NOR U61794 ( .A(n51352), .B(n41483), .Z(n41498) );
  NOR U61795 ( .A(n41484), .B(n41498), .Z(n41485) );
  NOR U61796 ( .A(n51350), .B(n41485), .Z(n41494) );
  NOR U61797 ( .A(n41487), .B(n41486), .Z(n41497) );
  IV U61798 ( .A(n41488), .Z(n41490) );
  NOR U61799 ( .A(n41490), .B(n41489), .Z(n41493) );
  NOR U61800 ( .A(n41497), .B(n41493), .Z(n41491) );
  IV U61801 ( .A(n41491), .Z(n41492) );
  NOR U61802 ( .A(n41494), .B(n41492), .Z(n41501) );
  IV U61803 ( .A(n41493), .Z(n41496) );
  IV U61804 ( .A(n41494), .Z(n41495) );
  NOR U61805 ( .A(n41496), .B(n41495), .Z(n56609) );
  IV U61806 ( .A(n41497), .Z(n41500) );
  IV U61807 ( .A(n41498), .Z(n41499) );
  NOR U61808 ( .A(n41500), .B(n41499), .Z(n56618) );
  NOR U61809 ( .A(n56609), .B(n56618), .Z(n52081) );
  IV U61810 ( .A(n52081), .Z(n45960) );
  NOR U61811 ( .A(n41501), .B(n45960), .Z(n45955) );
  XOR U61812 ( .A(n41502), .B(n45955), .Z(n52085) );
  IV U61813 ( .A(n41503), .Z(n41504) );
  NOR U61814 ( .A(n41505), .B(n41504), .Z(n52083) );
  IV U61815 ( .A(n41506), .Z(n41508) );
  NOR U61816 ( .A(n41508), .B(n41507), .Z(n52096) );
  NOR U61817 ( .A(n52083), .B(n52096), .Z(n45953) );
  XOR U61818 ( .A(n52085), .B(n45953), .Z(n45950) );
  XOR U61819 ( .A(n45951), .B(n45950), .Z(n46580) );
  IV U61820 ( .A(n41509), .Z(n41511) );
  NOR U61821 ( .A(n41511), .B(n41510), .Z(n46577) );
  IV U61822 ( .A(n41512), .Z(n41514) );
  NOR U61823 ( .A(n41514), .B(n41513), .Z(n46584) );
  NOR U61824 ( .A(n46577), .B(n46584), .Z(n46581) );
  XOR U61825 ( .A(n46580), .B(n46581), .Z(n45947) );
  XOR U61826 ( .A(n41515), .B(n45947), .Z(n62313) );
  XOR U61827 ( .A(n45942), .B(n62313), .Z(n45940) );
  XOR U61828 ( .A(n45944), .B(n45940), .Z(n46595) );
  XOR U61829 ( .A(n41516), .B(n46595), .Z(n46607) );
  IV U61830 ( .A(n41517), .Z(n41519) );
  NOR U61831 ( .A(n41519), .B(n41518), .Z(n52109) );
  IV U61832 ( .A(n41520), .Z(n41521) );
  NOR U61833 ( .A(n41522), .B(n41521), .Z(n52114) );
  NOR U61834 ( .A(n52109), .B(n52114), .Z(n46608) );
  XOR U61835 ( .A(n46607), .B(n46608), .Z(n46605) );
  XOR U61836 ( .A(n46606), .B(n46605), .Z(n46598) );
  XOR U61837 ( .A(n46599), .B(n46598), .Z(n45937) );
  IV U61838 ( .A(n41523), .Z(n41524) );
  NOR U61839 ( .A(n41525), .B(n41524), .Z(n46600) );
  IV U61840 ( .A(n41526), .Z(n41527) );
  NOR U61841 ( .A(n41528), .B(n41527), .Z(n45936) );
  NOR U61842 ( .A(n46600), .B(n45936), .Z(n41529) );
  XOR U61843 ( .A(n45937), .B(n41529), .Z(n51319) );
  IV U61844 ( .A(n51319), .Z(n51332) );
  XOR U61845 ( .A(n51320), .B(n51332), .Z(n46620) );
  NOR U61846 ( .A(n41531), .B(n41530), .Z(n41535) );
  NOR U61847 ( .A(n41533), .B(n41532), .Z(n51328) );
  NOR U61848 ( .A(n51328), .B(n51315), .Z(n41534) );
  NOR U61849 ( .A(n41535), .B(n41534), .Z(n46618) );
  XOR U61850 ( .A(n46620), .B(n46618), .Z(n51308) );
  IV U61851 ( .A(n51308), .Z(n41541) );
  IV U61852 ( .A(n41536), .Z(n41537) );
  NOR U61853 ( .A(n41538), .B(n41537), .Z(n51312) );
  NOR U61854 ( .A(n41540), .B(n41539), .Z(n51307) );
  NOR U61855 ( .A(n51312), .B(n51307), .Z(n46621) );
  XOR U61856 ( .A(n41541), .B(n46621), .Z(n56540) );
  XOR U61857 ( .A(n45933), .B(n56540), .Z(n51299) );
  XOR U61858 ( .A(n46626), .B(n51299), .Z(n46630) );
  IV U61859 ( .A(n41542), .Z(n41543) );
  NOR U61860 ( .A(n41544), .B(n41543), .Z(n46627) );
  IV U61861 ( .A(n41545), .Z(n41547) );
  NOR U61862 ( .A(n41547), .B(n41546), .Z(n46640) );
  NOR U61863 ( .A(n46627), .B(n46640), .Z(n41548) );
  XOR U61864 ( .A(n46630), .B(n41548), .Z(n46635) );
  XOR U61865 ( .A(n46634), .B(n46635), .Z(n45929) );
  XOR U61866 ( .A(n41549), .B(n45929), .Z(n45923) );
  XOR U61867 ( .A(n45926), .B(n45923), .Z(n45921) );
  IV U61868 ( .A(n41550), .Z(n41552) );
  NOR U61869 ( .A(n41552), .B(n41551), .Z(n45924) );
  IV U61870 ( .A(n41553), .Z(n41554) );
  NOR U61871 ( .A(n41555), .B(n41554), .Z(n45920) );
  NOR U61872 ( .A(n45924), .B(n45920), .Z(n41556) );
  XOR U61873 ( .A(n45921), .B(n41556), .Z(n45918) );
  XOR U61874 ( .A(n45919), .B(n45918), .Z(n51270) );
  IV U61875 ( .A(n41557), .Z(n41559) );
  NOR U61876 ( .A(n41559), .B(n41558), .Z(n51273) );
  IV U61877 ( .A(n41560), .Z(n41562) );
  NOR U61878 ( .A(n41562), .B(n41561), .Z(n51268) );
  NOR U61879 ( .A(n51273), .B(n51268), .Z(n46653) );
  XOR U61880 ( .A(n51270), .B(n46653), .Z(n45916) );
  XOR U61881 ( .A(n45917), .B(n45916), .Z(n51262) );
  IV U61882 ( .A(n41563), .Z(n41565) );
  NOR U61883 ( .A(n41565), .B(n41564), .Z(n51265) );
  IV U61884 ( .A(n41566), .Z(n41568) );
  NOR U61885 ( .A(n41568), .B(n41567), .Z(n51259) );
  NOR U61886 ( .A(n51265), .B(n51259), .Z(n45915) );
  XOR U61887 ( .A(n51262), .B(n45915), .Z(n41569) );
  IV U61888 ( .A(n41569), .Z(n45913) );
  XOR U61889 ( .A(n45912), .B(n45913), .Z(n45907) );
  IV U61890 ( .A(n41570), .Z(n41572) );
  NOR U61891 ( .A(n41572), .B(n41571), .Z(n45910) );
  IV U61892 ( .A(n41573), .Z(n41575) );
  NOR U61893 ( .A(n41575), .B(n41574), .Z(n52154) );
  NOR U61894 ( .A(n45910), .B(n52154), .Z(n41576) );
  XOR U61895 ( .A(n45907), .B(n41576), .Z(n41577) );
  IV U61896 ( .A(n41577), .Z(n46671) );
  XOR U61897 ( .A(n45905), .B(n46671), .Z(n46667) );
  IV U61898 ( .A(n41578), .Z(n41579) );
  NOR U61899 ( .A(n41580), .B(n41579), .Z(n46669) );
  IV U61900 ( .A(n41581), .Z(n41582) );
  NOR U61901 ( .A(n41583), .B(n41582), .Z(n46666) );
  NOR U61902 ( .A(n46669), .B(n46666), .Z(n41584) );
  XOR U61903 ( .A(n46667), .B(n41584), .Z(n45901) );
  IV U61904 ( .A(n45901), .Z(n56462) );
  IV U61905 ( .A(n41585), .Z(n41587) );
  NOR U61906 ( .A(n41587), .B(n41586), .Z(n56457) );
  IV U61907 ( .A(n41588), .Z(n41589) );
  NOR U61908 ( .A(n41590), .B(n41589), .Z(n56465) );
  NOR U61909 ( .A(n56457), .B(n56465), .Z(n51251) );
  IV U61910 ( .A(n51251), .Z(n45900) );
  XOR U61911 ( .A(n56462), .B(n45900), .Z(n52164) );
  XOR U61912 ( .A(n45902), .B(n52164), .Z(n45899) );
  IV U61913 ( .A(n41591), .Z(n41592) );
  NOR U61914 ( .A(n41593), .B(n41592), .Z(n45897) );
  IV U61915 ( .A(n41594), .Z(n41596) );
  NOR U61916 ( .A(n41596), .B(n41595), .Z(n45895) );
  NOR U61917 ( .A(n45897), .B(n45895), .Z(n41597) );
  XOR U61918 ( .A(n45899), .B(n41597), .Z(n45882) );
  IV U61919 ( .A(n41598), .Z(n41599) );
  NOR U61920 ( .A(n41600), .B(n41599), .Z(n45892) );
  IV U61921 ( .A(n41601), .Z(n41602) );
  NOR U61922 ( .A(n41603), .B(n41602), .Z(n45881) );
  NOR U61923 ( .A(n45892), .B(n45881), .Z(n41604) );
  XOR U61924 ( .A(n45882), .B(n41604), .Z(n45889) );
  IV U61925 ( .A(n41605), .Z(n41607) );
  NOR U61926 ( .A(n41607), .B(n41606), .Z(n45885) );
  IV U61927 ( .A(n41608), .Z(n41609) );
  NOR U61928 ( .A(n41610), .B(n41609), .Z(n45887) );
  NOR U61929 ( .A(n45885), .B(n45887), .Z(n41611) );
  XOR U61930 ( .A(n45889), .B(n41611), .Z(n52182) );
  NOR U61931 ( .A(n41612), .B(n52182), .Z(n41615) );
  IV U61932 ( .A(n41612), .Z(n41614) );
  XOR U61933 ( .A(n45885), .B(n45889), .Z(n41613) );
  NOR U61934 ( .A(n41614), .B(n41613), .Z(n52185) );
  NOR U61935 ( .A(n41615), .B(n52185), .Z(n45878) );
  IV U61936 ( .A(n41616), .Z(n41618) );
  NOR U61937 ( .A(n41618), .B(n41617), .Z(n52183) );
  IV U61938 ( .A(n41619), .Z(n41621) );
  NOR U61939 ( .A(n41621), .B(n41620), .Z(n51232) );
  NOR U61940 ( .A(n52183), .B(n51232), .Z(n45879) );
  XOR U61941 ( .A(n45878), .B(n45879), .Z(n46677) );
  IV U61942 ( .A(n41622), .Z(n41624) );
  NOR U61943 ( .A(n41624), .B(n41623), .Z(n46676) );
  IV U61944 ( .A(n41625), .Z(n41627) );
  NOR U61945 ( .A(n41627), .B(n41626), .Z(n45876) );
  NOR U61946 ( .A(n46676), .B(n45876), .Z(n41628) );
  XOR U61947 ( .A(n46677), .B(n41628), .Z(n46679) );
  XOR U61948 ( .A(n46680), .B(n46679), .Z(n51222) );
  XOR U61949 ( .A(n46681), .B(n51222), .Z(n45869) );
  IV U61950 ( .A(n41629), .Z(n41631) );
  NOR U61951 ( .A(n41631), .B(n41630), .Z(n57345) );
  NOR U61952 ( .A(n41633), .B(n41632), .Z(n56425) );
  NOR U61953 ( .A(n57345), .B(n56425), .Z(n45870) );
  XOR U61954 ( .A(n45869), .B(n45870), .Z(n45872) );
  XOR U61955 ( .A(n41634), .B(n45872), .Z(n45863) );
  XOR U61956 ( .A(n45864), .B(n45863), .Z(n52204) );
  XOR U61957 ( .A(n52206), .B(n52204), .Z(n46686) );
  XOR U61958 ( .A(n46688), .B(n46686), .Z(n51196) );
  IV U61959 ( .A(n41635), .Z(n41637) );
  NOR U61960 ( .A(n41637), .B(n41636), .Z(n51194) );
  IV U61961 ( .A(n41638), .Z(n41639) );
  NOR U61962 ( .A(n41640), .B(n41639), .Z(n52209) );
  NOR U61963 ( .A(n51194), .B(n52209), .Z(n46689) );
  XOR U61964 ( .A(n51196), .B(n46689), .Z(n45857) );
  XOR U61965 ( .A(n45858), .B(n45857), .Z(n45860) );
  XOR U61966 ( .A(n45859), .B(n45860), .Z(n46697) );
  IV U61967 ( .A(n41641), .Z(n41643) );
  NOR U61968 ( .A(n41643), .B(n41642), .Z(n45854) );
  IV U61969 ( .A(n41644), .Z(n41646) );
  NOR U61970 ( .A(n41646), .B(n41645), .Z(n46696) );
  NOR U61971 ( .A(n45854), .B(n46696), .Z(n41647) );
  XOR U61972 ( .A(n46697), .B(n41647), .Z(n41648) );
  IV U61973 ( .A(n41648), .Z(n46695) );
  IV U61974 ( .A(n41649), .Z(n41650) );
  NOR U61975 ( .A(n41651), .B(n41650), .Z(n41652) );
  IV U61976 ( .A(n41652), .Z(n41659) );
  NOR U61977 ( .A(n46695), .B(n41659), .Z(n51190) );
  IV U61978 ( .A(n41653), .Z(n41655) );
  NOR U61979 ( .A(n41655), .B(n41654), .Z(n45850) );
  IV U61980 ( .A(n41656), .Z(n41658) );
  NOR U61981 ( .A(n41658), .B(n41657), .Z(n46693) );
  XOR U61982 ( .A(n46693), .B(n46695), .Z(n45851) );
  IV U61983 ( .A(n45851), .Z(n41660) );
  XOR U61984 ( .A(n45850), .B(n41660), .Z(n41662) );
  NOR U61985 ( .A(n41660), .B(n41659), .Z(n41661) );
  NOR U61986 ( .A(n41662), .B(n41661), .Z(n41663) );
  NOR U61987 ( .A(n51190), .B(n41663), .Z(n45848) );
  IV U61988 ( .A(n41664), .Z(n41665) );
  NOR U61989 ( .A(n41666), .B(n41665), .Z(n45847) );
  IV U61990 ( .A(n41667), .Z(n41669) );
  NOR U61991 ( .A(n41669), .B(n41668), .Z(n46701) );
  NOR U61992 ( .A(n45847), .B(n46701), .Z(n41670) );
  XOR U61993 ( .A(n45848), .B(n41670), .Z(n45846) );
  IV U61994 ( .A(n41671), .Z(n41673) );
  NOR U61995 ( .A(n41673), .B(n41672), .Z(n45844) );
  IV U61996 ( .A(n41674), .Z(n41676) );
  NOR U61997 ( .A(n41676), .B(n41675), .Z(n45842) );
  NOR U61998 ( .A(n45844), .B(n45842), .Z(n41677) );
  XOR U61999 ( .A(n45846), .B(n41677), .Z(n45840) );
  IV U62000 ( .A(n41678), .Z(n41679) );
  NOR U62001 ( .A(n41680), .B(n41679), .Z(n45839) );
  IV U62002 ( .A(n41681), .Z(n41682) );
  NOR U62003 ( .A(n41683), .B(n41682), .Z(n46711) );
  NOR U62004 ( .A(n45839), .B(n46711), .Z(n41684) );
  XOR U62005 ( .A(n45840), .B(n41684), .Z(n51170) );
  NOR U62006 ( .A(n41686), .B(n41685), .Z(n51169) );
  IV U62007 ( .A(n41687), .Z(n41689) );
  NOR U62008 ( .A(n41689), .B(n41688), .Z(n52233) );
  NOR U62009 ( .A(n51169), .B(n52233), .Z(n45838) );
  IV U62010 ( .A(n45838), .Z(n51157) );
  XOR U62011 ( .A(n51170), .B(n51157), .Z(n45832) );
  IV U62012 ( .A(n41690), .Z(n41691) );
  NOR U62013 ( .A(n41692), .B(n41691), .Z(n51166) );
  IV U62014 ( .A(n41693), .Z(n41694) );
  NOR U62015 ( .A(n41695), .B(n41694), .Z(n51156) );
  NOR U62016 ( .A(n51166), .B(n51156), .Z(n45833) );
  XOR U62017 ( .A(n45832), .B(n45833), .Z(n45835) );
  XOR U62018 ( .A(n41696), .B(n45835), .Z(n56361) );
  XOR U62019 ( .A(n45830), .B(n56361), .Z(n46715) );
  XOR U62020 ( .A(n41697), .B(n46715), .Z(n41708) );
  IV U62021 ( .A(n41708), .Z(n41706) );
  IV U62022 ( .A(n41698), .Z(n41699) );
  NOR U62023 ( .A(n41700), .B(n41699), .Z(n41710) );
  IV U62024 ( .A(n41701), .Z(n41703) );
  NOR U62025 ( .A(n41703), .B(n41702), .Z(n41707) );
  NOR U62026 ( .A(n41710), .B(n41707), .Z(n41704) );
  IV U62027 ( .A(n41704), .Z(n41705) );
  NOR U62028 ( .A(n41706), .B(n41705), .Z(n41714) );
  IV U62029 ( .A(n41707), .Z(n41709) );
  NOR U62030 ( .A(n41709), .B(n41708), .Z(n56343) );
  IV U62031 ( .A(n41710), .Z(n41713) );
  IV U62032 ( .A(n41711), .Z(n46716) );
  XOR U62033 ( .A(n46716), .B(n46715), .Z(n41712) );
  NOR U62034 ( .A(n41713), .B(n41712), .Z(n56348) );
  NOR U62035 ( .A(n56343), .B(n56348), .Z(n52250) );
  IV U62036 ( .A(n52250), .Z(n46730) );
  NOR U62037 ( .A(n41714), .B(n46730), .Z(n45822) );
  NOR U62038 ( .A(n41716), .B(n41715), .Z(n45827) );
  IV U62039 ( .A(n41717), .Z(n41719) );
  NOR U62040 ( .A(n41719), .B(n41718), .Z(n51155) );
  NOR U62041 ( .A(n45827), .B(n51155), .Z(n41720) );
  XOR U62042 ( .A(n45822), .B(n41720), .Z(n46735) );
  IV U62043 ( .A(n41721), .Z(n41722) );
  NOR U62044 ( .A(n41723), .B(n41722), .Z(n45824) );
  IV U62045 ( .A(n41724), .Z(n41725) );
  NOR U62046 ( .A(n41726), .B(n41725), .Z(n46733) );
  NOR U62047 ( .A(n45824), .B(n46733), .Z(n41727) );
  XOR U62048 ( .A(n46735), .B(n41727), .Z(n45819) );
  IV U62049 ( .A(n41728), .Z(n41730) );
  NOR U62050 ( .A(n41730), .B(n41729), .Z(n46736) );
  IV U62051 ( .A(n41731), .Z(n41732) );
  NOR U62052 ( .A(n41733), .B(n41732), .Z(n45818) );
  NOR U62053 ( .A(n46736), .B(n45818), .Z(n41734) );
  XOR U62054 ( .A(n45819), .B(n41734), .Z(n52270) );
  XOR U62055 ( .A(n41735), .B(n52270), .Z(n46740) );
  XOR U62056 ( .A(n46742), .B(n46740), .Z(n57411) );
  IV U62057 ( .A(n57401), .Z(n41736) );
  NOR U62058 ( .A(n41736), .B(n57399), .Z(n41740) );
  NOR U62059 ( .A(n41738), .B(n41737), .Z(n41739) );
  NOR U62060 ( .A(n41740), .B(n41739), .Z(n46755) );
  XOR U62061 ( .A(n57411), .B(n46755), .Z(n51138) );
  IV U62062 ( .A(n51138), .Z(n51128) );
  IV U62063 ( .A(n41741), .Z(n41742) );
  NOR U62064 ( .A(n41743), .B(n41742), .Z(n51141) );
  IV U62065 ( .A(n41744), .Z(n41745) );
  NOR U62066 ( .A(n41746), .B(n41745), .Z(n51137) );
  NOR U62067 ( .A(n51141), .B(n51137), .Z(n46757) );
  IV U62068 ( .A(n46757), .Z(n51127) );
  XOR U62069 ( .A(n51128), .B(n51127), .Z(n57431) );
  XOR U62070 ( .A(n57429), .B(n57431), .Z(n46764) );
  IV U62071 ( .A(n41747), .Z(n41748) );
  NOR U62072 ( .A(n41749), .B(n41748), .Z(n57428) );
  IV U62073 ( .A(n41750), .Z(n41752) );
  NOR U62074 ( .A(n41752), .B(n41751), .Z(n57444) );
  NOR U62075 ( .A(n57428), .B(n57444), .Z(n46765) );
  XOR U62076 ( .A(n46764), .B(n46765), .Z(n45813) );
  XOR U62077 ( .A(n41753), .B(n45813), .Z(n52288) );
  IV U62078 ( .A(n41754), .Z(n41755) );
  NOR U62079 ( .A(n41756), .B(n41755), .Z(n52286) );
  IV U62080 ( .A(n41757), .Z(n41758) );
  NOR U62081 ( .A(n41759), .B(n41758), .Z(n52292) );
  NOR U62082 ( .A(n52286), .B(n52292), .Z(n45807) );
  XOR U62083 ( .A(n52288), .B(n45807), .Z(n45805) );
  XOR U62084 ( .A(n41760), .B(n45805), .Z(n66968) );
  NOR U62085 ( .A(n41762), .B(n41761), .Z(n66964) );
  IV U62086 ( .A(n41763), .Z(n41765) );
  NOR U62087 ( .A(n41765), .B(n41764), .Z(n68014) );
  NOR U62088 ( .A(n66964), .B(n68014), .Z(n46775) );
  XOR U62089 ( .A(n66968), .B(n46775), .Z(n46773) );
  XOR U62090 ( .A(n46777), .B(n46773), .Z(n46783) );
  XOR U62091 ( .A(n41766), .B(n46783), .Z(n45795) );
  XOR U62092 ( .A(n41767), .B(n45795), .Z(n45799) );
  XOR U62093 ( .A(n41768), .B(n45799), .Z(n45780) );
  IV U62094 ( .A(n41769), .Z(n41770) );
  NOR U62095 ( .A(n41771), .B(n41770), .Z(n45791) );
  IV U62096 ( .A(n41772), .Z(n41773) );
  NOR U62097 ( .A(n41774), .B(n41773), .Z(n45781) );
  NOR U62098 ( .A(n45791), .B(n45781), .Z(n41775) );
  XOR U62099 ( .A(n45780), .B(n41775), .Z(n45786) );
  XOR U62100 ( .A(n41776), .B(n45786), .Z(n45770) );
  IV U62101 ( .A(n41777), .Z(n41779) );
  NOR U62102 ( .A(n41779), .B(n41778), .Z(n45777) );
  IV U62103 ( .A(n41780), .Z(n41781) );
  NOR U62104 ( .A(n41782), .B(n41781), .Z(n45769) );
  NOR U62105 ( .A(n45777), .B(n45769), .Z(n41783) );
  XOR U62106 ( .A(n45770), .B(n41783), .Z(n45775) );
  IV U62107 ( .A(n41784), .Z(n41785) );
  NOR U62108 ( .A(n41786), .B(n41785), .Z(n45767) );
  IV U62109 ( .A(n41787), .Z(n41789) );
  NOR U62110 ( .A(n41789), .B(n41788), .Z(n45773) );
  NOR U62111 ( .A(n45767), .B(n45773), .Z(n41790) );
  XOR U62112 ( .A(n45775), .B(n41790), .Z(n52329) );
  IV U62113 ( .A(n41791), .Z(n41792) );
  NOR U62114 ( .A(n41793), .B(n41792), .Z(n52328) );
  IV U62115 ( .A(n41794), .Z(n41796) );
  NOR U62116 ( .A(n41796), .B(n41795), .Z(n52337) );
  NOR U62117 ( .A(n52328), .B(n52337), .Z(n46790) );
  XOR U62118 ( .A(n52329), .B(n46790), .Z(n51090) );
  XOR U62119 ( .A(n46792), .B(n51090), .Z(n46803) );
  XOR U62120 ( .A(n41797), .B(n46803), .Z(n41798) );
  IV U62121 ( .A(n41798), .Z(n46813) );
  XOR U62122 ( .A(n46796), .B(n46813), .Z(n46808) );
  XOR U62123 ( .A(n41799), .B(n46808), .Z(n46831) );
  XOR U62124 ( .A(n41800), .B(n46831), .Z(n51075) );
  XOR U62125 ( .A(n46833), .B(n51075), .Z(n46834) );
  XOR U62126 ( .A(n46835), .B(n46834), .Z(n45765) );
  IV U62127 ( .A(n41801), .Z(n41803) );
  NOR U62128 ( .A(n41803), .B(n41802), .Z(n45764) );
  IV U62129 ( .A(n41804), .Z(n41806) );
  NOR U62130 ( .A(n41806), .B(n41805), .Z(n51062) );
  NOR U62131 ( .A(n45764), .B(n51062), .Z(n41807) );
  XOR U62132 ( .A(n45765), .B(n41807), .Z(n46841) );
  XOR U62133 ( .A(n41808), .B(n46841), .Z(n52366) );
  XOR U62134 ( .A(n46845), .B(n52366), .Z(n51054) );
  IV U62135 ( .A(n51054), .Z(n41815) );
  IV U62136 ( .A(n41809), .Z(n41810) );
  NOR U62137 ( .A(n41811), .B(n41810), .Z(n52364) );
  IV U62138 ( .A(n41812), .Z(n41813) );
  NOR U62139 ( .A(n41814), .B(n41813), .Z(n51053) );
  NOR U62140 ( .A(n52364), .B(n51053), .Z(n46847) );
  XOR U62141 ( .A(n41815), .B(n46847), .Z(n46862) );
  XOR U62142 ( .A(n45757), .B(n46862), .Z(n46855) );
  XOR U62143 ( .A(n41816), .B(n46855), .Z(n45750) );
  XOR U62144 ( .A(n41817), .B(n45750), .Z(n45754) );
  IV U62145 ( .A(n41818), .Z(n41820) );
  NOR U62146 ( .A(n41820), .B(n41819), .Z(n45748) );
  IV U62147 ( .A(n41821), .Z(n41822) );
  NOR U62148 ( .A(n41823), .B(n41822), .Z(n45753) );
  NOR U62149 ( .A(n45748), .B(n45753), .Z(n41824) );
  XOR U62150 ( .A(n45754), .B(n41824), .Z(n45743) );
  XOR U62151 ( .A(n45744), .B(n45743), .Z(n46878) );
  XOR U62152 ( .A(n41825), .B(n46878), .Z(n41826) );
  IV U62153 ( .A(n41826), .Z(n46874) );
  XOR U62154 ( .A(n41827), .B(n46874), .Z(n41837) );
  IV U62155 ( .A(n41837), .Z(n41828) );
  NOR U62156 ( .A(n41840), .B(n41828), .Z(n46897) );
  IV U62157 ( .A(n41829), .Z(n41830) );
  NOR U62158 ( .A(n41831), .B(n41830), .Z(n46901) );
  IV U62159 ( .A(n41832), .Z(n41834) );
  NOR U62160 ( .A(n41834), .B(n41833), .Z(n41838) );
  IV U62161 ( .A(n41838), .Z(n41836) );
  XOR U62162 ( .A(n45741), .B(n46874), .Z(n41835) );
  NOR U62163 ( .A(n41836), .B(n41835), .Z(n46893) );
  NOR U62164 ( .A(n41838), .B(n41837), .Z(n41839) );
  NOR U62165 ( .A(n46893), .B(n41839), .Z(n46902) );
  XOR U62166 ( .A(n46901), .B(n46902), .Z(n41842) );
  NOR U62167 ( .A(n46902), .B(n41840), .Z(n41841) );
  NOR U62168 ( .A(n41842), .B(n41841), .Z(n41843) );
  NOR U62169 ( .A(n46897), .B(n41843), .Z(n45739) );
  XOR U62170 ( .A(n45740), .B(n45739), .Z(n45737) );
  IV U62171 ( .A(n41844), .Z(n41846) );
  NOR U62172 ( .A(n41846), .B(n41845), .Z(n46908) );
  IV U62173 ( .A(n41847), .Z(n41849) );
  NOR U62174 ( .A(n41849), .B(n41848), .Z(n45736) );
  NOR U62175 ( .A(n46908), .B(n45736), .Z(n41850) );
  XOR U62176 ( .A(n45737), .B(n41850), .Z(n45730) );
  XOR U62177 ( .A(n41851), .B(n45730), .Z(n51017) );
  XOR U62178 ( .A(n46913), .B(n51017), .Z(n46914) );
  XOR U62179 ( .A(n46915), .B(n46914), .Z(n45728) );
  XOR U62180 ( .A(n45727), .B(n45728), .Z(n56193) );
  XOR U62181 ( .A(n45724), .B(n56193), .Z(n45721) );
  XOR U62182 ( .A(n45726), .B(n45721), .Z(n45718) );
  IV U62183 ( .A(n41852), .Z(n41854) );
  NOR U62184 ( .A(n41854), .B(n41853), .Z(n45720) );
  IV U62185 ( .A(n41855), .Z(n41856) );
  NOR U62186 ( .A(n41857), .B(n41856), .Z(n45717) );
  NOR U62187 ( .A(n45720), .B(n45717), .Z(n41858) );
  XOR U62188 ( .A(n45718), .B(n41858), .Z(n46921) );
  IV U62189 ( .A(n41859), .Z(n41860) );
  NOR U62190 ( .A(n41861), .B(n41860), .Z(n52411) );
  IV U62191 ( .A(n41862), .Z(n41863) );
  NOR U62192 ( .A(n41864), .B(n41863), .Z(n52407) );
  NOR U62193 ( .A(n52411), .B(n52407), .Z(n46922) );
  XOR U62194 ( .A(n46921), .B(n46922), .Z(n46928) );
  IV U62195 ( .A(n41865), .Z(n41867) );
  NOR U62196 ( .A(n41867), .B(n41866), .Z(n46923) );
  IV U62197 ( .A(n41868), .Z(n41870) );
  NOR U62198 ( .A(n41870), .B(n41869), .Z(n46927) );
  NOR U62199 ( .A(n46923), .B(n46927), .Z(n41871) );
  XOR U62200 ( .A(n46928), .B(n41871), .Z(n45715) );
  XOR U62201 ( .A(n41872), .B(n45715), .Z(n46939) );
  IV U62202 ( .A(n41873), .Z(n41875) );
  NOR U62203 ( .A(n41875), .B(n41874), .Z(n46933) );
  IV U62204 ( .A(n41876), .Z(n41877) );
  NOR U62205 ( .A(n41878), .B(n41877), .Z(n46938) );
  NOR U62206 ( .A(n46933), .B(n46938), .Z(n41879) );
  XOR U62207 ( .A(n46939), .B(n41879), .Z(n45711) );
  IV U62208 ( .A(n41880), .Z(n41881) );
  NOR U62209 ( .A(n41882), .B(n41881), .Z(n46935) );
  IV U62210 ( .A(n41883), .Z(n41885) );
  NOR U62211 ( .A(n41885), .B(n41884), .Z(n45712) );
  NOR U62212 ( .A(n46935), .B(n45712), .Z(n41886) );
  XOR U62213 ( .A(n45711), .B(n41886), .Z(n56149) );
  IV U62214 ( .A(n41887), .Z(n41889) );
  NOR U62215 ( .A(n41889), .B(n41888), .Z(n56155) );
  IV U62216 ( .A(n41890), .Z(n41892) );
  NOR U62217 ( .A(n41892), .B(n41891), .Z(n56144) );
  NOR U62218 ( .A(n56155), .B(n56144), .Z(n46944) );
  XOR U62219 ( .A(n56149), .B(n46944), .Z(n45709) );
  XOR U62220 ( .A(n41893), .B(n45709), .Z(n50993) );
  XOR U62221 ( .A(n46954), .B(n50993), .Z(n46955) );
  XOR U62222 ( .A(n50990), .B(n46955), .Z(n50980) );
  IV U62223 ( .A(n41894), .Z(n41895) );
  NOR U62224 ( .A(n41896), .B(n41895), .Z(n50984) );
  IV U62225 ( .A(n41897), .Z(n41898) );
  NOR U62226 ( .A(n41899), .B(n41898), .Z(n50979) );
  NOR U62227 ( .A(n50984), .B(n50979), .Z(n46959) );
  XOR U62228 ( .A(n50980), .B(n46959), .Z(n45706) );
  XOR U62229 ( .A(n41900), .B(n45706), .Z(n46968) );
  IV U62230 ( .A(n46968), .Z(n41908) );
  IV U62231 ( .A(n41901), .Z(n41902) );
  NOR U62232 ( .A(n41903), .B(n41902), .Z(n45703) );
  IV U62233 ( .A(n41904), .Z(n41905) );
  NOR U62234 ( .A(n41906), .B(n41905), .Z(n46967) );
  NOR U62235 ( .A(n45703), .B(n46967), .Z(n41907) );
  XOR U62236 ( .A(n41908), .B(n41907), .Z(n46974) );
  XOR U62237 ( .A(n46965), .B(n46974), .Z(n45701) );
  XOR U62238 ( .A(n41909), .B(n45701), .Z(n45694) );
  XOR U62239 ( .A(n45698), .B(n45694), .Z(n45692) );
  IV U62240 ( .A(n41910), .Z(n41912) );
  NOR U62241 ( .A(n41912), .B(n41911), .Z(n45695) );
  IV U62242 ( .A(n41913), .Z(n41915) );
  NOR U62243 ( .A(n41915), .B(n41914), .Z(n45691) );
  NOR U62244 ( .A(n45695), .B(n45691), .Z(n41916) );
  XOR U62245 ( .A(n45692), .B(n41916), .Z(n45688) );
  IV U62246 ( .A(n41917), .Z(n41919) );
  NOR U62247 ( .A(n41919), .B(n41918), .Z(n45689) );
  IV U62248 ( .A(n41920), .Z(n41921) );
  NOR U62249 ( .A(n41922), .B(n41921), .Z(n46979) );
  NOR U62250 ( .A(n45689), .B(n46979), .Z(n41923) );
  XOR U62251 ( .A(n45688), .B(n41923), .Z(n46977) );
  IV U62252 ( .A(n46977), .Z(n41931) );
  IV U62253 ( .A(n41924), .Z(n41925) );
  NOR U62254 ( .A(n41926), .B(n41925), .Z(n46976) );
  IV U62255 ( .A(n41927), .Z(n41929) );
  NOR U62256 ( .A(n41929), .B(n41928), .Z(n45686) );
  NOR U62257 ( .A(n46976), .B(n45686), .Z(n41930) );
  XOR U62258 ( .A(n41931), .B(n41930), .Z(n45684) );
  XOR U62259 ( .A(n45681), .B(n45684), .Z(n41932) );
  NOR U62260 ( .A(n41933), .B(n41932), .Z(n52454) );
  IV U62261 ( .A(n41934), .Z(n41936) );
  NOR U62262 ( .A(n41936), .B(n41935), .Z(n45683) );
  NOR U62263 ( .A(n45681), .B(n45683), .Z(n41937) );
  XOR U62264 ( .A(n41937), .B(n45684), .Z(n45678) );
  NOR U62265 ( .A(n41938), .B(n45678), .Z(n41939) );
  NOR U62266 ( .A(n52454), .B(n41939), .Z(n45674) );
  IV U62267 ( .A(n41940), .Z(n41941) );
  NOR U62268 ( .A(n41942), .B(n41941), .Z(n45677) );
  IV U62269 ( .A(n41943), .Z(n41945) );
  NOR U62270 ( .A(n41945), .B(n41944), .Z(n45673) );
  NOR U62271 ( .A(n45677), .B(n45673), .Z(n41946) );
  XOR U62272 ( .A(n45674), .B(n41946), .Z(n56123) );
  IV U62273 ( .A(n41947), .Z(n41948) );
  NOR U62274 ( .A(n41949), .B(n41948), .Z(n56119) );
  IV U62275 ( .A(n41950), .Z(n41951) );
  NOR U62276 ( .A(n41952), .B(n41951), .Z(n57635) );
  NOR U62277 ( .A(n56119), .B(n57635), .Z(n45672) );
  XOR U62278 ( .A(n56123), .B(n45672), .Z(n57650) );
  IV U62279 ( .A(n41953), .Z(n41954) );
  NOR U62280 ( .A(n41955), .B(n41954), .Z(n45668) );
  IV U62281 ( .A(n41956), .Z(n41958) );
  NOR U62282 ( .A(n41958), .B(n41957), .Z(n45669) );
  NOR U62283 ( .A(n45668), .B(n45669), .Z(n41959) );
  XOR U62284 ( .A(n57650), .B(n41959), .Z(n45663) );
  XOR U62285 ( .A(n45664), .B(n45663), .Z(n45666) );
  IV U62286 ( .A(n41960), .Z(n41961) );
  NOR U62287 ( .A(n41962), .B(n41961), .Z(n45665) );
  IV U62288 ( .A(n41963), .Z(n41965) );
  NOR U62289 ( .A(n41965), .B(n41964), .Z(n46994) );
  NOR U62290 ( .A(n45665), .B(n46994), .Z(n41966) );
  XOR U62291 ( .A(n45666), .B(n41966), .Z(n46992) );
  IV U62292 ( .A(n41967), .Z(n41969) );
  NOR U62293 ( .A(n41969), .B(n41968), .Z(n46990) );
  IV U62294 ( .A(n41970), .Z(n41972) );
  NOR U62295 ( .A(n41972), .B(n41971), .Z(n45661) );
  NOR U62296 ( .A(n46990), .B(n45661), .Z(n41973) );
  XOR U62297 ( .A(n46992), .B(n41973), .Z(n45655) );
  IV U62298 ( .A(n41974), .Z(n41976) );
  NOR U62299 ( .A(n41976), .B(n41975), .Z(n45654) );
  IV U62300 ( .A(n41977), .Z(n41979) );
  NOR U62301 ( .A(n41979), .B(n41978), .Z(n45657) );
  NOR U62302 ( .A(n45654), .B(n45657), .Z(n41980) );
  XOR U62303 ( .A(n45655), .B(n41980), .Z(n56101) );
  XOR U62304 ( .A(n45653), .B(n56101), .Z(n45647) );
  XOR U62305 ( .A(n45648), .B(n45647), .Z(n45645) );
  IV U62306 ( .A(n41981), .Z(n41983) );
  NOR U62307 ( .A(n41983), .B(n41982), .Z(n45649) );
  IV U62308 ( .A(n41984), .Z(n41985) );
  NOR U62309 ( .A(n41986), .B(n41985), .Z(n45644) );
  NOR U62310 ( .A(n45649), .B(n45644), .Z(n41987) );
  XOR U62311 ( .A(n45645), .B(n41987), .Z(n45639) );
  IV U62312 ( .A(n41988), .Z(n41989) );
  NOR U62313 ( .A(n41990), .B(n41989), .Z(n56082) );
  IV U62314 ( .A(n41991), .Z(n41992) );
  NOR U62315 ( .A(n41993), .B(n41992), .Z(n57668) );
  NOR U62316 ( .A(n56082), .B(n57668), .Z(n50927) );
  XOR U62317 ( .A(n45639), .B(n50927), .Z(n45641) );
  XOR U62318 ( .A(n45640), .B(n45641), .Z(n47007) );
  IV U62319 ( .A(n41994), .Z(n41996) );
  NOR U62320 ( .A(n41996), .B(n41995), .Z(n45637) );
  IV U62321 ( .A(n41997), .Z(n41998) );
  NOR U62322 ( .A(n41999), .B(n41998), .Z(n47006) );
  NOR U62323 ( .A(n45637), .B(n47006), .Z(n42000) );
  XOR U62324 ( .A(n47007), .B(n42000), .Z(n42001) );
  IV U62325 ( .A(n42001), .Z(n47013) );
  IV U62326 ( .A(n42002), .Z(n42003) );
  NOR U62327 ( .A(n42004), .B(n42003), .Z(n47011) );
  IV U62328 ( .A(n42005), .Z(n42007) );
  NOR U62329 ( .A(n42007), .B(n42006), .Z(n47009) );
  NOR U62330 ( .A(n47011), .B(n47009), .Z(n42008) );
  XOR U62331 ( .A(n47013), .B(n42008), .Z(n42009) );
  NOR U62332 ( .A(n42010), .B(n42009), .Z(n42013) );
  IV U62333 ( .A(n42010), .Z(n42012) );
  XOR U62334 ( .A(n47011), .B(n47013), .Z(n42011) );
  NOR U62335 ( .A(n42012), .B(n42011), .Z(n52491) );
  NOR U62336 ( .A(n42013), .B(n52491), .Z(n45635) );
  XOR U62337 ( .A(n42014), .B(n45635), .Z(n45631) );
  IV U62338 ( .A(n42015), .Z(n42016) );
  NOR U62339 ( .A(n42017), .B(n42016), .Z(n45630) );
  IV U62340 ( .A(n42018), .Z(n42019) );
  NOR U62341 ( .A(n42020), .B(n42019), .Z(n45625) );
  NOR U62342 ( .A(n45630), .B(n45625), .Z(n42021) );
  XOR U62343 ( .A(n45631), .B(n42021), .Z(n47022) );
  IV U62344 ( .A(n42022), .Z(n42024) );
  NOR U62345 ( .A(n42024), .B(n42023), .Z(n45627) );
  IV U62346 ( .A(n42025), .Z(n42027) );
  NOR U62347 ( .A(n42027), .B(n42026), .Z(n47021) );
  NOR U62348 ( .A(n45627), .B(n47021), .Z(n42028) );
  XOR U62349 ( .A(n47022), .B(n42028), .Z(n47029) );
  XOR U62350 ( .A(n42029), .B(n47029), .Z(n42037) );
  IV U62351 ( .A(n42037), .Z(n42030) );
  NOR U62352 ( .A(n42031), .B(n42030), .Z(n50891) );
  IV U62353 ( .A(n42032), .Z(n42033) );
  NOR U62354 ( .A(n42034), .B(n42033), .Z(n42038) );
  IV U62355 ( .A(n42038), .Z(n42036) );
  XOR U62356 ( .A(n47027), .B(n47029), .Z(n42035) );
  NOR U62357 ( .A(n42036), .B(n42035), .Z(n50889) );
  NOR U62358 ( .A(n42038), .B(n42037), .Z(n42039) );
  NOR U62359 ( .A(n50889), .B(n42039), .Z(n42040) );
  NOR U62360 ( .A(n42041), .B(n42040), .Z(n42042) );
  NOR U62361 ( .A(n50891), .B(n42042), .Z(n45620) );
  IV U62362 ( .A(n42043), .Z(n42045) );
  NOR U62363 ( .A(n42045), .B(n42044), .Z(n47032) );
  IV U62364 ( .A(n42046), .Z(n42047) );
  NOR U62365 ( .A(n42048), .B(n42047), .Z(n42049) );
  NOR U62366 ( .A(n47032), .B(n42049), .Z(n45621) );
  XOR U62367 ( .A(n45620), .B(n45621), .Z(n45618) );
  XOR U62368 ( .A(n45615), .B(n45618), .Z(n42050) );
  NOR U62369 ( .A(n42051), .B(n42050), .Z(n50879) );
  IV U62370 ( .A(n42052), .Z(n42053) );
  NOR U62371 ( .A(n42054), .B(n42053), .Z(n45617) );
  NOR U62372 ( .A(n45615), .B(n45617), .Z(n42055) );
  XOR U62373 ( .A(n45618), .B(n42055), .Z(n42056) );
  NOR U62374 ( .A(n42057), .B(n42056), .Z(n42058) );
  NOR U62375 ( .A(n50879), .B(n42058), .Z(n45612) );
  XOR U62376 ( .A(n45613), .B(n45612), .Z(n45609) );
  IV U62377 ( .A(n45609), .Z(n42066) );
  IV U62378 ( .A(n42059), .Z(n42060) );
  NOR U62379 ( .A(n42061), .B(n42060), .Z(n45608) );
  IV U62380 ( .A(n42062), .Z(n42064) );
  NOR U62381 ( .A(n42064), .B(n42063), .Z(n45606) );
  NOR U62382 ( .A(n45608), .B(n45606), .Z(n42065) );
  XOR U62383 ( .A(n42066), .B(n42065), .Z(n47046) );
  XOR U62384 ( .A(n47040), .B(n47046), .Z(n45604) );
  XOR U62385 ( .A(n42067), .B(n45604), .Z(n47055) );
  IV U62386 ( .A(n42068), .Z(n42070) );
  NOR U62387 ( .A(n42070), .B(n42069), .Z(n47056) );
  IV U62388 ( .A(n42071), .Z(n42072) );
  NOR U62389 ( .A(n42073), .B(n42072), .Z(n47060) );
  NOR U62390 ( .A(n47056), .B(n47060), .Z(n42074) );
  XOR U62391 ( .A(n47055), .B(n42074), .Z(n47068) );
  IV U62392 ( .A(n42075), .Z(n42077) );
  NOR U62393 ( .A(n42077), .B(n42076), .Z(n47052) );
  IV U62394 ( .A(n42078), .Z(n42079) );
  NOR U62395 ( .A(n42080), .B(n42079), .Z(n47067) );
  NOR U62396 ( .A(n47052), .B(n47067), .Z(n42081) );
  XOR U62397 ( .A(n47068), .B(n42081), .Z(n42082) );
  IV U62398 ( .A(n42082), .Z(n47074) );
  XOR U62399 ( .A(n47065), .B(n47074), .Z(n45601) );
  IV U62400 ( .A(n42083), .Z(n42085) );
  NOR U62401 ( .A(n42085), .B(n42084), .Z(n47072) );
  IV U62402 ( .A(n42086), .Z(n42087) );
  NOR U62403 ( .A(n42088), .B(n42087), .Z(n45600) );
  NOR U62404 ( .A(n47072), .B(n45600), .Z(n42089) );
  XOR U62405 ( .A(n45601), .B(n42089), .Z(n45593) );
  IV U62406 ( .A(n42090), .Z(n42091) );
  NOR U62407 ( .A(n42092), .B(n42091), .Z(n45597) );
  IV U62408 ( .A(n42093), .Z(n42094) );
  NOR U62409 ( .A(n42095), .B(n42094), .Z(n45594) );
  NOR U62410 ( .A(n45597), .B(n45594), .Z(n42096) );
  XOR U62411 ( .A(n45593), .B(n42096), .Z(n47079) );
  XOR U62412 ( .A(n47077), .B(n47079), .Z(n45591) );
  XOR U62413 ( .A(n45592), .B(n45591), .Z(n47086) );
  XOR U62414 ( .A(n47087), .B(n47086), .Z(n47093) );
  XOR U62415 ( .A(n47088), .B(n47093), .Z(n45589) );
  IV U62416 ( .A(n45589), .Z(n42104) );
  IV U62417 ( .A(n42097), .Z(n42098) );
  NOR U62418 ( .A(n42099), .B(n42098), .Z(n47092) );
  IV U62419 ( .A(n42100), .Z(n42102) );
  NOR U62420 ( .A(n42102), .B(n42101), .Z(n45588) );
  NOR U62421 ( .A(n47092), .B(n45588), .Z(n42103) );
  XOR U62422 ( .A(n42104), .B(n42103), .Z(n45587) );
  IV U62423 ( .A(n42105), .Z(n42106) );
  NOR U62424 ( .A(n42107), .B(n42106), .Z(n45583) );
  IV U62425 ( .A(n42108), .Z(n42109) );
  NOR U62426 ( .A(n42110), .B(n42109), .Z(n45585) );
  NOR U62427 ( .A(n45583), .B(n45585), .Z(n42111) );
  XOR U62428 ( .A(n45587), .B(n42111), .Z(n42123) );
  NOR U62429 ( .A(n42112), .B(n42123), .Z(n42115) );
  IV U62430 ( .A(n42112), .Z(n42114) );
  XOR U62431 ( .A(n45583), .B(n45587), .Z(n42113) );
  NOR U62432 ( .A(n42114), .B(n42113), .Z(n50822) );
  NOR U62433 ( .A(n42115), .B(n50822), .Z(n42121) );
  IV U62434 ( .A(n42121), .Z(n42116) );
  NOR U62435 ( .A(n42117), .B(n42116), .Z(n52538) );
  IV U62436 ( .A(n42118), .Z(n42120) );
  NOR U62437 ( .A(n42120), .B(n42119), .Z(n42122) );
  NOR U62438 ( .A(n42122), .B(n42121), .Z(n42126) );
  IV U62439 ( .A(n42122), .Z(n42125) );
  IV U62440 ( .A(n42123), .Z(n42124) );
  NOR U62441 ( .A(n42125), .B(n42124), .Z(n52535) );
  NOR U62442 ( .A(n42126), .B(n52535), .Z(n42134) );
  NOR U62443 ( .A(n42127), .B(n42134), .Z(n42128) );
  NOR U62444 ( .A(n52538), .B(n42128), .Z(n42137) );
  IV U62445 ( .A(n42137), .Z(n42129) );
  NOR U62446 ( .A(n42130), .B(n42129), .Z(n52550) );
  IV U62447 ( .A(n42131), .Z(n42132) );
  NOR U62448 ( .A(n42133), .B(n42132), .Z(n42138) );
  IV U62449 ( .A(n42138), .Z(n42136) );
  IV U62450 ( .A(n42134), .Z(n42135) );
  NOR U62451 ( .A(n42136), .B(n42135), .Z(n52542) );
  NOR U62452 ( .A(n42138), .B(n42137), .Z(n42139) );
  NOR U62453 ( .A(n52542), .B(n42139), .Z(n52548) );
  NOR U62454 ( .A(n42140), .B(n52548), .Z(n42141) );
  NOR U62455 ( .A(n52550), .B(n42141), .Z(n47097) );
  XOR U62456 ( .A(n47098), .B(n47097), .Z(n45581) );
  NOR U62457 ( .A(n42143), .B(n42142), .Z(n45580) );
  IV U62458 ( .A(n42144), .Z(n42146) );
  NOR U62459 ( .A(n42146), .B(n42145), .Z(n45576) );
  NOR U62460 ( .A(n45580), .B(n45576), .Z(n42147) );
  XOR U62461 ( .A(n45581), .B(n42147), .Z(n42148) );
  IV U62462 ( .A(n42148), .Z(n45574) );
  XOR U62463 ( .A(n45573), .B(n45574), .Z(n45569) );
  XOR U62464 ( .A(n42149), .B(n45569), .Z(n45562) );
  XOR U62465 ( .A(n42150), .B(n45562), .Z(n45560) );
  XOR U62466 ( .A(n45557), .B(n45560), .Z(n42151) );
  NOR U62467 ( .A(n42152), .B(n42151), .Z(n52568) );
  IV U62468 ( .A(n42153), .Z(n42154) );
  NOR U62469 ( .A(n42155), .B(n42154), .Z(n45559) );
  NOR U62470 ( .A(n45557), .B(n45559), .Z(n42156) );
  XOR U62471 ( .A(n42156), .B(n45560), .Z(n42164) );
  NOR U62472 ( .A(n42157), .B(n42164), .Z(n42158) );
  NOR U62473 ( .A(n52568), .B(n42158), .Z(n42167) );
  IV U62474 ( .A(n42167), .Z(n42159) );
  NOR U62475 ( .A(n42160), .B(n42159), .Z(n52576) );
  IV U62476 ( .A(n42161), .Z(n42163) );
  NOR U62477 ( .A(n42163), .B(n42162), .Z(n42168) );
  IV U62478 ( .A(n42168), .Z(n42166) );
  IV U62479 ( .A(n42164), .Z(n42165) );
  NOR U62480 ( .A(n42166), .B(n42165), .Z(n45556) );
  NOR U62481 ( .A(n42168), .B(n42167), .Z(n42169) );
  NOR U62482 ( .A(n45556), .B(n42169), .Z(n42170) );
  NOR U62483 ( .A(n42171), .B(n42170), .Z(n42172) );
  NOR U62484 ( .A(n52576), .B(n42172), .Z(n47107) );
  XOR U62485 ( .A(n42173), .B(n47107), .Z(n47125) );
  XOR U62486 ( .A(n42174), .B(n47125), .Z(n47115) );
  IV U62487 ( .A(n42175), .Z(n42177) );
  NOR U62488 ( .A(n42177), .B(n42176), .Z(n47124) );
  IV U62489 ( .A(n42178), .Z(n42179) );
  NOR U62490 ( .A(n42180), .B(n42179), .Z(n47114) );
  NOR U62491 ( .A(n47124), .B(n47114), .Z(n42181) );
  XOR U62492 ( .A(n47115), .B(n42181), .Z(n45552) );
  IV U62493 ( .A(n42182), .Z(n42183) );
  NOR U62494 ( .A(n42184), .B(n42183), .Z(n45550) );
  IV U62495 ( .A(n42185), .Z(n42186) );
  NOR U62496 ( .A(n42187), .B(n42186), .Z(n45548) );
  NOR U62497 ( .A(n45550), .B(n45548), .Z(n42188) );
  XOR U62498 ( .A(n45552), .B(n42188), .Z(n42189) );
  IV U62499 ( .A(n42189), .Z(n50787) );
  XOR U62500 ( .A(n45547), .B(n50787), .Z(n45543) );
  IV U62501 ( .A(n45543), .Z(n50782) );
  IV U62502 ( .A(n42190), .Z(n42191) );
  NOR U62503 ( .A(n42192), .B(n42191), .Z(n57766) );
  IV U62504 ( .A(n42193), .Z(n42194) );
  NOR U62505 ( .A(n42195), .B(n42194), .Z(n57772) );
  NOR U62506 ( .A(n57766), .B(n57772), .Z(n50784) );
  IV U62507 ( .A(n50784), .Z(n45542) );
  XOR U62508 ( .A(n50782), .B(n45542), .Z(n47137) );
  NOR U62509 ( .A(n42197), .B(n42196), .Z(n45544) );
  IV U62510 ( .A(n42198), .Z(n42200) );
  NOR U62511 ( .A(n42200), .B(n42199), .Z(n47136) );
  NOR U62512 ( .A(n45544), .B(n47136), .Z(n42201) );
  XOR U62513 ( .A(n47137), .B(n42201), .Z(n42202) );
  IV U62514 ( .A(n42202), .Z(n50765) );
  XOR U62515 ( .A(n47134), .B(n50765), .Z(n45540) );
  XOR U62516 ( .A(n45541), .B(n45540), .Z(n45534) );
  XOR U62517 ( .A(n45535), .B(n45534), .Z(n45537) );
  IV U62518 ( .A(n45537), .Z(n42210) );
  IV U62519 ( .A(n42203), .Z(n42204) );
  NOR U62520 ( .A(n42205), .B(n42204), .Z(n45536) );
  IV U62521 ( .A(n42206), .Z(n42207) );
  NOR U62522 ( .A(n42208), .B(n42207), .Z(n45532) );
  NOR U62523 ( .A(n45536), .B(n45532), .Z(n42209) );
  XOR U62524 ( .A(n42210), .B(n42209), .Z(n45531) );
  XOR U62525 ( .A(n45529), .B(n45531), .Z(n45524) );
  XOR U62526 ( .A(n42211), .B(n45524), .Z(n45517) );
  XOR U62527 ( .A(n42212), .B(n45517), .Z(n52598) );
  XOR U62528 ( .A(n47144), .B(n52598), .Z(n47146) );
  IV U62529 ( .A(n42213), .Z(n42214) );
  NOR U62530 ( .A(n42215), .B(n42214), .Z(n47145) );
  IV U62531 ( .A(n42216), .Z(n42217) );
  NOR U62532 ( .A(n42218), .B(n42217), .Z(n52616) );
  NOR U62533 ( .A(n47145), .B(n52616), .Z(n42219) );
  XOR U62534 ( .A(n47146), .B(n42219), .Z(n47153) );
  XOR U62535 ( .A(n47152), .B(n47153), .Z(n42220) );
  NOR U62536 ( .A(n42221), .B(n42220), .Z(n55913) );
  IV U62537 ( .A(n42222), .Z(n42224) );
  NOR U62538 ( .A(n42224), .B(n42223), .Z(n45515) );
  NOR U62539 ( .A(n47152), .B(n45515), .Z(n42225) );
  XOR U62540 ( .A(n42225), .B(n47153), .Z(n42226) );
  NOR U62541 ( .A(n42227), .B(n42226), .Z(n42228) );
  NOR U62542 ( .A(n55913), .B(n42228), .Z(n42229) );
  IV U62543 ( .A(n42229), .Z(n47157) );
  XOR U62544 ( .A(n47156), .B(n47157), .Z(n45511) );
  XOR U62545 ( .A(n42230), .B(n45511), .Z(n45504) );
  XOR U62546 ( .A(n45503), .B(n45504), .Z(n42231) );
  NOR U62547 ( .A(n42232), .B(n42231), .Z(n50720) );
  IV U62548 ( .A(n42233), .Z(n42234) );
  NOR U62549 ( .A(n42235), .B(n42234), .Z(n45501) );
  NOR U62550 ( .A(n45503), .B(n45501), .Z(n42236) );
  XOR U62551 ( .A(n42236), .B(n45504), .Z(n47163) );
  NOR U62552 ( .A(n42237), .B(n47163), .Z(n42238) );
  NOR U62553 ( .A(n50720), .B(n42238), .Z(n45498) );
  XOR U62554 ( .A(n42239), .B(n45498), .Z(n45496) );
  XOR U62555 ( .A(n45494), .B(n45496), .Z(n45489) );
  IV U62556 ( .A(n42240), .Z(n42241) );
  NOR U62557 ( .A(n42242), .B(n42241), .Z(n45492) );
  IV U62558 ( .A(n42243), .Z(n42244) );
  NOR U62559 ( .A(n42245), .B(n42244), .Z(n45488) );
  NOR U62560 ( .A(n45492), .B(n45488), .Z(n42246) );
  XOR U62561 ( .A(n45489), .B(n42246), .Z(n45480) );
  IV U62562 ( .A(n42247), .Z(n42249) );
  NOR U62563 ( .A(n42249), .B(n42248), .Z(n45486) );
  IV U62564 ( .A(n42250), .Z(n42251) );
  NOR U62565 ( .A(n42252), .B(n42251), .Z(n45481) );
  NOR U62566 ( .A(n45486), .B(n45481), .Z(n42253) );
  XOR U62567 ( .A(n45480), .B(n42253), .Z(n45484) );
  XOR U62568 ( .A(n45483), .B(n45484), .Z(n45473) );
  IV U62569 ( .A(n42254), .Z(n42255) );
  NOR U62570 ( .A(n42256), .B(n42255), .Z(n45477) );
  IV U62571 ( .A(n42257), .Z(n42259) );
  NOR U62572 ( .A(n42259), .B(n42258), .Z(n45472) );
  NOR U62573 ( .A(n45477), .B(n45472), .Z(n42260) );
  XOR U62574 ( .A(n45473), .B(n42260), .Z(n42269) );
  IV U62575 ( .A(n42269), .Z(n47171) );
  XOR U62576 ( .A(n45470), .B(n47171), .Z(n42261) );
  NOR U62577 ( .A(n42270), .B(n42261), .Z(n47168) );
  IV U62578 ( .A(n42262), .Z(n42263) );
  NOR U62579 ( .A(n42264), .B(n42263), .Z(n45467) );
  IV U62580 ( .A(n42265), .Z(n42267) );
  NOR U62581 ( .A(n42267), .B(n42266), .Z(n47169) );
  NOR U62582 ( .A(n45470), .B(n47169), .Z(n42268) );
  XOR U62583 ( .A(n42269), .B(n42268), .Z(n45468) );
  IV U62584 ( .A(n45468), .Z(n42271) );
  XOR U62585 ( .A(n45467), .B(n42271), .Z(n42273) );
  NOR U62586 ( .A(n42271), .B(n42270), .Z(n42272) );
  NOR U62587 ( .A(n42273), .B(n42272), .Z(n42274) );
  NOR U62588 ( .A(n47168), .B(n42274), .Z(n45463) );
  IV U62589 ( .A(n42275), .Z(n42277) );
  NOR U62590 ( .A(n42277), .B(n42276), .Z(n55866) );
  IV U62591 ( .A(n42278), .Z(n42280) );
  NOR U62592 ( .A(n42280), .B(n42279), .Z(n55858) );
  NOR U62593 ( .A(n55866), .B(n55858), .Z(n45464) );
  XOR U62594 ( .A(n45463), .B(n45464), .Z(n47182) );
  IV U62595 ( .A(n42281), .Z(n42283) );
  NOR U62596 ( .A(n42283), .B(n42282), .Z(n45465) );
  IV U62597 ( .A(n42284), .Z(n42285) );
  NOR U62598 ( .A(n42286), .B(n42285), .Z(n47181) );
  NOR U62599 ( .A(n45465), .B(n47181), .Z(n42287) );
  XOR U62600 ( .A(n47182), .B(n42287), .Z(n42288) );
  IV U62601 ( .A(n42288), .Z(n47188) );
  XOR U62602 ( .A(n47179), .B(n47188), .Z(n45461) );
  IV U62603 ( .A(n42289), .Z(n42291) );
  NOR U62604 ( .A(n42291), .B(n42290), .Z(n47186) );
  IV U62605 ( .A(n42292), .Z(n42293) );
  NOR U62606 ( .A(n42294), .B(n42293), .Z(n45460) );
  NOR U62607 ( .A(n47186), .B(n45460), .Z(n42295) );
  XOR U62608 ( .A(n45461), .B(n42295), .Z(n47189) );
  IV U62609 ( .A(n42296), .Z(n42297) );
  NOR U62610 ( .A(n42298), .B(n42297), .Z(n47195) );
  IV U62611 ( .A(n42299), .Z(n42301) );
  NOR U62612 ( .A(n42301), .B(n42300), .Z(n47190) );
  NOR U62613 ( .A(n47195), .B(n47190), .Z(n42302) );
  XOR U62614 ( .A(n47189), .B(n42302), .Z(n47205) );
  XOR U62615 ( .A(n47193), .B(n47205), .Z(n47208) );
  IV U62616 ( .A(n42303), .Z(n42305) );
  NOR U62617 ( .A(n42305), .B(n42304), .Z(n47204) );
  IV U62618 ( .A(n42306), .Z(n42307) );
  NOR U62619 ( .A(n42308), .B(n42307), .Z(n47207) );
  NOR U62620 ( .A(n47204), .B(n47207), .Z(n42309) );
  XOR U62621 ( .A(n47208), .B(n42309), .Z(n45454) );
  IV U62622 ( .A(n42310), .Z(n42312) );
  NOR U62623 ( .A(n42312), .B(n42311), .Z(n45457) );
  IV U62624 ( .A(n42313), .Z(n42314) );
  NOR U62625 ( .A(n42315), .B(n42314), .Z(n45455) );
  NOR U62626 ( .A(n45457), .B(n45455), .Z(n42316) );
  XOR U62627 ( .A(n45454), .B(n42316), .Z(n45452) );
  XOR U62628 ( .A(n45451), .B(n45452), .Z(n47214) );
  IV U62629 ( .A(n42317), .Z(n42318) );
  NOR U62630 ( .A(n42319), .B(n42318), .Z(n45449) );
  IV U62631 ( .A(n42320), .Z(n42321) );
  NOR U62632 ( .A(n42322), .B(n42321), .Z(n47213) );
  NOR U62633 ( .A(n45449), .B(n47213), .Z(n42323) );
  XOR U62634 ( .A(n47214), .B(n42323), .Z(n45439) );
  IV U62635 ( .A(n42324), .Z(n42325) );
  NOR U62636 ( .A(n42326), .B(n42325), .Z(n47210) );
  IV U62637 ( .A(n42327), .Z(n42328) );
  NOR U62638 ( .A(n42329), .B(n42328), .Z(n45440) );
  NOR U62639 ( .A(n47210), .B(n45440), .Z(n42330) );
  XOR U62640 ( .A(n45439), .B(n42330), .Z(n45445) );
  IV U62641 ( .A(n42331), .Z(n42333) );
  NOR U62642 ( .A(n42333), .B(n42332), .Z(n45444) );
  IV U62643 ( .A(n42334), .Z(n42336) );
  NOR U62644 ( .A(n42336), .B(n42335), .Z(n45442) );
  NOR U62645 ( .A(n45444), .B(n45442), .Z(n42337) );
  XOR U62646 ( .A(n45445), .B(n42337), .Z(n45433) );
  IV U62647 ( .A(n42338), .Z(n42339) );
  NOR U62648 ( .A(n42340), .B(n42339), .Z(n45436) );
  IV U62649 ( .A(n42341), .Z(n42342) );
  NOR U62650 ( .A(n42343), .B(n42342), .Z(n45432) );
  NOR U62651 ( .A(n45436), .B(n45432), .Z(n42344) );
  XOR U62652 ( .A(n45433), .B(n42344), .Z(n63048) );
  XOR U62653 ( .A(n45429), .B(n63048), .Z(n42345) );
  IV U62654 ( .A(n42345), .Z(n45427) );
  XOR U62655 ( .A(n42346), .B(n45427), .Z(n42358) );
  NOR U62656 ( .A(n42347), .B(n42358), .Z(n42350) );
  IV U62657 ( .A(n42347), .Z(n42349) );
  XOR U62658 ( .A(n45424), .B(n45427), .Z(n42348) );
  NOR U62659 ( .A(n42349), .B(n42348), .Z(n50644) );
  NOR U62660 ( .A(n42350), .B(n50644), .Z(n42354) );
  NOR U62661 ( .A(n42353), .B(n42354), .Z(n42351) );
  IV U62662 ( .A(n42351), .Z(n42352) );
  NOR U62663 ( .A(n42357), .B(n42352), .Z(n42362) );
  IV U62664 ( .A(n42353), .Z(n42356) );
  IV U62665 ( .A(n42354), .Z(n42355) );
  NOR U62666 ( .A(n42356), .B(n42355), .Z(n50642) );
  IV U62667 ( .A(n42357), .Z(n42360) );
  IV U62668 ( .A(n42358), .Z(n42359) );
  NOR U62669 ( .A(n42360), .B(n42359), .Z(n50647) );
  NOR U62670 ( .A(n50642), .B(n50647), .Z(n42361) );
  IV U62671 ( .A(n42361), .Z(n45423) );
  NOR U62672 ( .A(n42362), .B(n45423), .Z(n47222) );
  IV U62673 ( .A(n42363), .Z(n42364) );
  NOR U62674 ( .A(n42365), .B(n42364), .Z(n47226) );
  IV U62675 ( .A(n42366), .Z(n42367) );
  NOR U62676 ( .A(n42368), .B(n42367), .Z(n47221) );
  NOR U62677 ( .A(n47226), .B(n47221), .Z(n42369) );
  XOR U62678 ( .A(n47222), .B(n42369), .Z(n47240) );
  XOR U62679 ( .A(n47236), .B(n47240), .Z(n45421) );
  IV U62680 ( .A(n42370), .Z(n42372) );
  NOR U62681 ( .A(n42372), .B(n42371), .Z(n47238) );
  IV U62682 ( .A(n42373), .Z(n42374) );
  NOR U62683 ( .A(n42375), .B(n42374), .Z(n45420) );
  NOR U62684 ( .A(n47238), .B(n45420), .Z(n42376) );
  XOR U62685 ( .A(n45421), .B(n42376), .Z(n45414) );
  XOR U62686 ( .A(n45415), .B(n45414), .Z(n45417) );
  XOR U62687 ( .A(n45416), .B(n45417), .Z(n47243) );
  XOR U62688 ( .A(n42377), .B(n47243), .Z(n47246) );
  XOR U62689 ( .A(n47247), .B(n47246), .Z(n50620) );
  IV U62690 ( .A(n42378), .Z(n42380) );
  NOR U62691 ( .A(n42380), .B(n42379), .Z(n50617) );
  IV U62692 ( .A(n42381), .Z(n42383) );
  NOR U62693 ( .A(n42383), .B(n42382), .Z(n52704) );
  NOR U62694 ( .A(n50617), .B(n52704), .Z(n47249) );
  XOR U62695 ( .A(n50620), .B(n47249), .Z(n45406) );
  XOR U62696 ( .A(n42384), .B(n45406), .Z(n45400) );
  IV U62697 ( .A(n42385), .Z(n42387) );
  NOR U62698 ( .A(n42387), .B(n42386), .Z(n45404) );
  IV U62699 ( .A(n42388), .Z(n42389) );
  NOR U62700 ( .A(n42390), .B(n42389), .Z(n45399) );
  NOR U62701 ( .A(n45404), .B(n45399), .Z(n42391) );
  XOR U62702 ( .A(n45400), .B(n42391), .Z(n45392) );
  IV U62703 ( .A(n42392), .Z(n42394) );
  NOR U62704 ( .A(n42394), .B(n42393), .Z(n45396) );
  IV U62705 ( .A(n42395), .Z(n42396) );
  NOR U62706 ( .A(n42397), .B(n42396), .Z(n45393) );
  NOR U62707 ( .A(n45396), .B(n45393), .Z(n42398) );
  XOR U62708 ( .A(n45392), .B(n42398), .Z(n52715) );
  XOR U62709 ( .A(n52717), .B(n52715), .Z(n47254) );
  XOR U62710 ( .A(n47255), .B(n47254), .Z(n45390) );
  XOR U62711 ( .A(n42399), .B(n45390), .Z(n42400) );
  IV U62712 ( .A(n42400), .Z(n45388) );
  XOR U62713 ( .A(n45386), .B(n45388), .Z(n47263) );
  IV U62714 ( .A(n42401), .Z(n42402) );
  NOR U62715 ( .A(n42403), .B(n42402), .Z(n45383) );
  IV U62716 ( .A(n42404), .Z(n42405) );
  NOR U62717 ( .A(n42406), .B(n42405), .Z(n47262) );
  NOR U62718 ( .A(n45383), .B(n47262), .Z(n42407) );
  XOR U62719 ( .A(n47263), .B(n42407), .Z(n47265) );
  IV U62720 ( .A(n42408), .Z(n42409) );
  NOR U62721 ( .A(n42410), .B(n42409), .Z(n55766) );
  IV U62722 ( .A(n42411), .Z(n42413) );
  NOR U62723 ( .A(n42413), .B(n42412), .Z(n55761) );
  NOR U62724 ( .A(n55766), .B(n55761), .Z(n52730) );
  XOR U62725 ( .A(n47265), .B(n52730), .Z(n47267) );
  IV U62726 ( .A(n42414), .Z(n42416) );
  NOR U62727 ( .A(n42416), .B(n42415), .Z(n47266) );
  IV U62728 ( .A(n42417), .Z(n42419) );
  NOR U62729 ( .A(n42419), .B(n42418), .Z(n45381) );
  NOR U62730 ( .A(n47266), .B(n45381), .Z(n42420) );
  XOR U62731 ( .A(n47267), .B(n42420), .Z(n45374) );
  IV U62732 ( .A(n42421), .Z(n42422) );
  NOR U62733 ( .A(n42423), .B(n42422), .Z(n45378) );
  IV U62734 ( .A(n42424), .Z(n42425) );
  NOR U62735 ( .A(n42426), .B(n42425), .Z(n52737) );
  NOR U62736 ( .A(n45378), .B(n52737), .Z(n42427) );
  XOR U62737 ( .A(n45374), .B(n42427), .Z(n45373) );
  XOR U62738 ( .A(n42428), .B(n45373), .Z(n47284) );
  XOR U62739 ( .A(n42429), .B(n47284), .Z(n47279) );
  IV U62740 ( .A(n42430), .Z(n42431) );
  NOR U62741 ( .A(n42432), .B(n42431), .Z(n47283) );
  IV U62742 ( .A(n42433), .Z(n42435) );
  NOR U62743 ( .A(n42435), .B(n42434), .Z(n47278) );
  NOR U62744 ( .A(n47283), .B(n47278), .Z(n42436) );
  XOR U62745 ( .A(n47279), .B(n42436), .Z(n45361) );
  IV U62746 ( .A(n42437), .Z(n42439) );
  NOR U62747 ( .A(n42439), .B(n42438), .Z(n45365) );
  IV U62748 ( .A(n42440), .Z(n42441) );
  NOR U62749 ( .A(n42442), .B(n42441), .Z(n45362) );
  NOR U62750 ( .A(n45365), .B(n45362), .Z(n42443) );
  XOR U62751 ( .A(n45361), .B(n42443), .Z(n52758) );
  XOR U62752 ( .A(n45360), .B(n52758), .Z(n45354) );
  XOR U62753 ( .A(n42444), .B(n45354), .Z(n47297) );
  XOR U62754 ( .A(n42445), .B(n47297), .Z(n47306) );
  XOR U62755 ( .A(n42446), .B(n47306), .Z(n45349) );
  XOR U62756 ( .A(n42447), .B(n45349), .Z(n45343) );
  IV U62757 ( .A(n42448), .Z(n42450) );
  NOR U62758 ( .A(n42450), .B(n42449), .Z(n45342) );
  IV U62759 ( .A(n42451), .Z(n42453) );
  NOR U62760 ( .A(n42453), .B(n42452), .Z(n47322) );
  NOR U62761 ( .A(n45342), .B(n47322), .Z(n42454) );
  XOR U62762 ( .A(n45343), .B(n42454), .Z(n47321) );
  XOR U62763 ( .A(n42455), .B(n47321), .Z(n45338) );
  XOR U62764 ( .A(n45339), .B(n45338), .Z(n47334) );
  IV U62765 ( .A(n47334), .Z(n42463) );
  IV U62766 ( .A(n42456), .Z(n42458) );
  NOR U62767 ( .A(n42458), .B(n42457), .Z(n45336) );
  IV U62768 ( .A(n42459), .Z(n42461) );
  NOR U62769 ( .A(n42461), .B(n42460), .Z(n47333) );
  NOR U62770 ( .A(n45336), .B(n47333), .Z(n42462) );
  XOR U62771 ( .A(n42463), .B(n42462), .Z(n45335) );
  IV U62772 ( .A(n42464), .Z(n42466) );
  NOR U62773 ( .A(n42466), .B(n42465), .Z(n45333) );
  IV U62774 ( .A(n42467), .Z(n42468) );
  NOR U62775 ( .A(n42469), .B(n42468), .Z(n45331) );
  NOR U62776 ( .A(n45333), .B(n45331), .Z(n42470) );
  XOR U62777 ( .A(n45335), .B(n42470), .Z(n47343) );
  IV U62778 ( .A(n42471), .Z(n42472) );
  NOR U62779 ( .A(n42473), .B(n42472), .Z(n45328) );
  IV U62780 ( .A(n42474), .Z(n42475) );
  NOR U62781 ( .A(n42476), .B(n42475), .Z(n47342) );
  NOR U62782 ( .A(n45328), .B(n47342), .Z(n42477) );
  XOR U62783 ( .A(n47343), .B(n42477), .Z(n47341) );
  XOR U62784 ( .A(n47339), .B(n47341), .Z(n50550) );
  XOR U62785 ( .A(n45323), .B(n50550), .Z(n45325) );
  IV U62786 ( .A(n42478), .Z(n42479) );
  NOR U62787 ( .A(n42480), .B(n42479), .Z(n45324) );
  IV U62788 ( .A(n42481), .Z(n42483) );
  NOR U62789 ( .A(n42483), .B(n42482), .Z(n47347) );
  NOR U62790 ( .A(n45324), .B(n47347), .Z(n42484) );
  XOR U62791 ( .A(n45325), .B(n42484), .Z(n45322) );
  XOR U62792 ( .A(n45318), .B(n45322), .Z(n45316) );
  XOR U62793 ( .A(n42485), .B(n45316), .Z(n45311) );
  XOR U62794 ( .A(n45312), .B(n45311), .Z(n52809) );
  XOR U62795 ( .A(n45313), .B(n52809), .Z(n47355) );
  IV U62796 ( .A(n42486), .Z(n42488) );
  NOR U62797 ( .A(n42488), .B(n42487), .Z(n57986) );
  IV U62798 ( .A(n42489), .Z(n42490) );
  NOR U62799 ( .A(n42491), .B(n42490), .Z(n55680) );
  NOR U62800 ( .A(n57986), .B(n55680), .Z(n50533) );
  XOR U62801 ( .A(n47355), .B(n50533), .Z(n47357) );
  XOR U62802 ( .A(n42492), .B(n47357), .Z(n45302) );
  IV U62803 ( .A(n42493), .Z(n42494) );
  NOR U62804 ( .A(n42495), .B(n42494), .Z(n45305) );
  IV U62805 ( .A(n42496), .Z(n42497) );
  NOR U62806 ( .A(n42498), .B(n42497), .Z(n45301) );
  NOR U62807 ( .A(n45305), .B(n45301), .Z(n42499) );
  XOR U62808 ( .A(n45302), .B(n42499), .Z(n47368) );
  IV U62809 ( .A(n42500), .Z(n42501) );
  NOR U62810 ( .A(n42502), .B(n42501), .Z(n47362) );
  IV U62811 ( .A(n42503), .Z(n42504) );
  NOR U62812 ( .A(n42505), .B(n42504), .Z(n47366) );
  NOR U62813 ( .A(n47362), .B(n47366), .Z(n42506) );
  XOR U62814 ( .A(n47368), .B(n42506), .Z(n45295) );
  IV U62815 ( .A(n42507), .Z(n42509) );
  NOR U62816 ( .A(n42509), .B(n42508), .Z(n45298) );
  IV U62817 ( .A(n42510), .Z(n42512) );
  NOR U62818 ( .A(n42512), .B(n42511), .Z(n45294) );
  NOR U62819 ( .A(n45298), .B(n45294), .Z(n42513) );
  XOR U62820 ( .A(n45295), .B(n42513), .Z(n50511) );
  IV U62821 ( .A(n42514), .Z(n42515) );
  NOR U62822 ( .A(n42516), .B(n42515), .Z(n50508) );
  IV U62823 ( .A(n42517), .Z(n42518) );
  NOR U62824 ( .A(n42519), .B(n42518), .Z(n52832) );
  NOR U62825 ( .A(n50508), .B(n52832), .Z(n45293) );
  XOR U62826 ( .A(n50511), .B(n45293), .Z(n45291) );
  IV U62827 ( .A(n42520), .Z(n42522) );
  NOR U62828 ( .A(n42522), .B(n42521), .Z(n52829) );
  IV U62829 ( .A(n42523), .Z(n42524) );
  NOR U62830 ( .A(n42525), .B(n42524), .Z(n50502) );
  NOR U62831 ( .A(n52829), .B(n50502), .Z(n45292) );
  XOR U62832 ( .A(n45291), .B(n45292), .Z(n50496) );
  XOR U62833 ( .A(n45286), .B(n50496), .Z(n45284) );
  IV U62834 ( .A(n42526), .Z(n42528) );
  NOR U62835 ( .A(n42528), .B(n42527), .Z(n45287) );
  IV U62836 ( .A(n42529), .Z(n42530) );
  NOR U62837 ( .A(n42531), .B(n42530), .Z(n45283) );
  NOR U62838 ( .A(n45287), .B(n45283), .Z(n42532) );
  XOR U62839 ( .A(n45284), .B(n42532), .Z(n47383) );
  XOR U62840 ( .A(n47378), .B(n47383), .Z(n45281) );
  XOR U62841 ( .A(n42533), .B(n45281), .Z(n47392) );
  XOR U62842 ( .A(n45278), .B(n47392), .Z(n45276) );
  IV U62843 ( .A(n42534), .Z(n42535) );
  NOR U62844 ( .A(n42536), .B(n42535), .Z(n47390) );
  IV U62845 ( .A(n42537), .Z(n42539) );
  NOR U62846 ( .A(n42539), .B(n42538), .Z(n45275) );
  NOR U62847 ( .A(n47390), .B(n45275), .Z(n42540) );
  XOR U62848 ( .A(n45276), .B(n42540), .Z(n45271) );
  IV U62849 ( .A(n42541), .Z(n42543) );
  NOR U62850 ( .A(n42543), .B(n42542), .Z(n47393) );
  IV U62851 ( .A(n42544), .Z(n42546) );
  NOR U62852 ( .A(n42546), .B(n42545), .Z(n45272) );
  NOR U62853 ( .A(n47393), .B(n45272), .Z(n42547) );
  XOR U62854 ( .A(n45271), .B(n42547), .Z(n50471) );
  IV U62855 ( .A(n42548), .Z(n42550) );
  NOR U62856 ( .A(n42550), .B(n42549), .Z(n55643) );
  IV U62857 ( .A(n42551), .Z(n42553) );
  NOR U62858 ( .A(n42553), .B(n42552), .Z(n55638) );
  NOR U62859 ( .A(n55643), .B(n55638), .Z(n50473) );
  XOR U62860 ( .A(n50471), .B(n50473), .Z(n47398) );
  XOR U62861 ( .A(n47399), .B(n47398), .Z(n47401) );
  IV U62862 ( .A(n42554), .Z(n42555) );
  NOR U62863 ( .A(n42556), .B(n42555), .Z(n47400) );
  IV U62864 ( .A(n42557), .Z(n42559) );
  NOR U62865 ( .A(n42559), .B(n42558), .Z(n45269) );
  NOR U62866 ( .A(n47400), .B(n45269), .Z(n42560) );
  XOR U62867 ( .A(n47401), .B(n42560), .Z(n42568) );
  IV U62868 ( .A(n42568), .Z(n42561) );
  NOR U62869 ( .A(n42562), .B(n42561), .Z(n50458) );
  IV U62870 ( .A(n42563), .Z(n42565) );
  NOR U62871 ( .A(n42565), .B(n42564), .Z(n42569) );
  IV U62872 ( .A(n42569), .Z(n42567) );
  XOR U62873 ( .A(n47400), .B(n47401), .Z(n42566) );
  NOR U62874 ( .A(n42567), .B(n42566), .Z(n52863) );
  NOR U62875 ( .A(n42569), .B(n42568), .Z(n42570) );
  NOR U62876 ( .A(n52863), .B(n42570), .Z(n42580) );
  NOR U62877 ( .A(n42571), .B(n42580), .Z(n42572) );
  NOR U62878 ( .A(n50458), .B(n42572), .Z(n42578) );
  IV U62879 ( .A(n42578), .Z(n42573) );
  NOR U62880 ( .A(n42574), .B(n42573), .Z(n50450) );
  IV U62881 ( .A(n42575), .Z(n42576) );
  NOR U62882 ( .A(n42577), .B(n42576), .Z(n42579) );
  NOR U62883 ( .A(n42579), .B(n42578), .Z(n42583) );
  IV U62884 ( .A(n42579), .Z(n42582) );
  IV U62885 ( .A(n42580), .Z(n42581) );
  NOR U62886 ( .A(n42582), .B(n42581), .Z(n50455) );
  NOR U62887 ( .A(n42583), .B(n50455), .Z(n45260) );
  NOR U62888 ( .A(n42584), .B(n45260), .Z(n42585) );
  NOR U62889 ( .A(n50450), .B(n42585), .Z(n45263) );
  NOR U62890 ( .A(n42587), .B(n42586), .Z(n42591) );
  NOR U62891 ( .A(n42589), .B(n42588), .Z(n42590) );
  NOR U62892 ( .A(n42591), .B(n42590), .Z(n42592) );
  IV U62893 ( .A(n42592), .Z(n45264) );
  XOR U62894 ( .A(n45263), .B(n45264), .Z(n47411) );
  XOR U62895 ( .A(n47408), .B(n47411), .Z(n47415) );
  IV U62896 ( .A(n42593), .Z(n42595) );
  NOR U62897 ( .A(n42595), .B(n42594), .Z(n47410) );
  IV U62898 ( .A(n42596), .Z(n42598) );
  NOR U62899 ( .A(n42598), .B(n42597), .Z(n47414) );
  NOR U62900 ( .A(n47410), .B(n47414), .Z(n42599) );
  XOR U62901 ( .A(n47415), .B(n42599), .Z(n45253) );
  IV U62902 ( .A(n42600), .Z(n42601) );
  NOR U62903 ( .A(n42602), .B(n42601), .Z(n50443) );
  IV U62904 ( .A(n42603), .Z(n42605) );
  NOR U62905 ( .A(n42605), .B(n42604), .Z(n52891) );
  NOR U62906 ( .A(n50443), .B(n52891), .Z(n45254) );
  XOR U62907 ( .A(n45253), .B(n45254), .Z(n45256) );
  IV U62908 ( .A(n42606), .Z(n42607) );
  NOR U62909 ( .A(n42608), .B(n42607), .Z(n45255) );
  IV U62910 ( .A(n42609), .Z(n42610) );
  NOR U62911 ( .A(n42611), .B(n42610), .Z(n45251) );
  NOR U62912 ( .A(n45255), .B(n45251), .Z(n42612) );
  XOR U62913 ( .A(n45256), .B(n42612), .Z(n47422) );
  XOR U62914 ( .A(n47420), .B(n47422), .Z(n50427) );
  IV U62915 ( .A(n42613), .Z(n42615) );
  NOR U62916 ( .A(n42615), .B(n42614), .Z(n47419) );
  NOR U62917 ( .A(n42617), .B(n42616), .Z(n47428) );
  NOR U62918 ( .A(n47419), .B(n47428), .Z(n50429) );
  XOR U62919 ( .A(n50427), .B(n50429), .Z(n47427) );
  IV U62920 ( .A(n42618), .Z(n42619) );
  NOR U62921 ( .A(n42620), .B(n42619), .Z(n55604) );
  IV U62922 ( .A(n42621), .Z(n42622) );
  NOR U62923 ( .A(n42623), .B(n42622), .Z(n55599) );
  NOR U62924 ( .A(n55604), .B(n55599), .Z(n50425) );
  XOR U62925 ( .A(n47427), .B(n50425), .Z(n47437) );
  IV U62926 ( .A(n42624), .Z(n42626) );
  NOR U62927 ( .A(n42626), .B(n42625), .Z(n47434) );
  NOR U62928 ( .A(n42628), .B(n42627), .Z(n47436) );
  NOR U62929 ( .A(n47434), .B(n47436), .Z(n42629) );
  XOR U62930 ( .A(n47437), .B(n42629), .Z(n47432) );
  XOR U62931 ( .A(n47433), .B(n47432), .Z(n50410) );
  XOR U62932 ( .A(n50412), .B(n50410), .Z(n47443) );
  XOR U62933 ( .A(n47446), .B(n47443), .Z(n47452) );
  XOR U62934 ( .A(n42630), .B(n47452), .Z(n42631) );
  IV U62935 ( .A(n42631), .Z(n52916) );
  XOR U62936 ( .A(n47450), .B(n52916), .Z(n47463) );
  XOR U62937 ( .A(n42632), .B(n47463), .Z(n47477) );
  IV U62938 ( .A(n42633), .Z(n42635) );
  NOR U62939 ( .A(n42635), .B(n42634), .Z(n47456) );
  IV U62940 ( .A(n42636), .Z(n42638) );
  NOR U62941 ( .A(n42638), .B(n42637), .Z(n47476) );
  NOR U62942 ( .A(n47456), .B(n47476), .Z(n42639) );
  XOR U62943 ( .A(n47477), .B(n42639), .Z(n42640) );
  IV U62944 ( .A(n42640), .Z(n47484) );
  IV U62945 ( .A(n47481), .Z(n42641) );
  NOR U62946 ( .A(n42641), .B(n47479), .Z(n42645) );
  NOR U62947 ( .A(n42643), .B(n42642), .Z(n42644) );
  NOR U62948 ( .A(n42645), .B(n42644), .Z(n47474) );
  XOR U62949 ( .A(n47484), .B(n47474), .Z(n47493) );
  XOR U62950 ( .A(n42646), .B(n47493), .Z(n47488) );
  IV U62951 ( .A(n42647), .Z(n42648) );
  NOR U62952 ( .A(n42649), .B(n42648), .Z(n47487) );
  IV U62953 ( .A(n42650), .Z(n42651) );
  NOR U62954 ( .A(n42652), .B(n42651), .Z(n47497) );
  NOR U62955 ( .A(n47487), .B(n47497), .Z(n42653) );
  XOR U62956 ( .A(n47488), .B(n42653), .Z(n45250) );
  IV U62957 ( .A(n42654), .Z(n42656) );
  NOR U62958 ( .A(n42656), .B(n42655), .Z(n45248) );
  IV U62959 ( .A(n42657), .Z(n42659) );
  NOR U62960 ( .A(n42659), .B(n42658), .Z(n45245) );
  NOR U62961 ( .A(n45248), .B(n45245), .Z(n42660) );
  XOR U62962 ( .A(n45250), .B(n42660), .Z(n45243) );
  XOR U62963 ( .A(n45244), .B(n45243), .Z(n50386) );
  XOR U62964 ( .A(n47508), .B(n50386), .Z(n47509) );
  NOR U62965 ( .A(n42662), .B(n42661), .Z(n50381) );
  IV U62966 ( .A(n42663), .Z(n42665) );
  NOR U62967 ( .A(n42665), .B(n42664), .Z(n50376) );
  NOR U62968 ( .A(n50381), .B(n50376), .Z(n47510) );
  XOR U62969 ( .A(n47509), .B(n47510), .Z(n50371) );
  XOR U62970 ( .A(n45241), .B(n50371), .Z(n45236) );
  NOR U62971 ( .A(n42667), .B(n42666), .Z(n50364) );
  IV U62972 ( .A(n42668), .Z(n42670) );
  NOR U62973 ( .A(n42670), .B(n42669), .Z(n50359) );
  NOR U62974 ( .A(n50364), .B(n50359), .Z(n45237) );
  XOR U62975 ( .A(n45236), .B(n45237), .Z(n50353) );
  XOR U62976 ( .A(n45238), .B(n50353), .Z(n42671) );
  IV U62977 ( .A(n42671), .Z(n47516) );
  IV U62978 ( .A(n42672), .Z(n42673) );
  NOR U62979 ( .A(n42674), .B(n42673), .Z(n45233) );
  IV U62980 ( .A(n42675), .Z(n42676) );
  NOR U62981 ( .A(n42677), .B(n42676), .Z(n47515) );
  NOR U62982 ( .A(n45233), .B(n47515), .Z(n42678) );
  XOR U62983 ( .A(n47516), .B(n42678), .Z(n42685) );
  IV U62984 ( .A(n42685), .Z(n42679) );
  NOR U62985 ( .A(n42680), .B(n42679), .Z(n52955) );
  NOR U62986 ( .A(n42682), .B(n42681), .Z(n42686) );
  IV U62987 ( .A(n42686), .Z(n42684) );
  XOR U62988 ( .A(n45233), .B(n47516), .Z(n42683) );
  NOR U62989 ( .A(n42684), .B(n42683), .Z(n52951) );
  NOR U62990 ( .A(n42686), .B(n42685), .Z(n42687) );
  NOR U62991 ( .A(n52951), .B(n42687), .Z(n45230) );
  NOR U62992 ( .A(n42688), .B(n45230), .Z(n42689) );
  NOR U62993 ( .A(n52955), .B(n42689), .Z(n45225) );
  IV U62994 ( .A(n42690), .Z(n42691) );
  NOR U62995 ( .A(n42692), .B(n42691), .Z(n45229) );
  IV U62996 ( .A(n42693), .Z(n42695) );
  NOR U62997 ( .A(n42695), .B(n42694), .Z(n45224) );
  NOR U62998 ( .A(n45229), .B(n45224), .Z(n42696) );
  XOR U62999 ( .A(n45225), .B(n42696), .Z(n50339) );
  NOR U63000 ( .A(n42698), .B(n42697), .Z(n50337) );
  IV U63001 ( .A(n42699), .Z(n42701) );
  NOR U63002 ( .A(n42701), .B(n42700), .Z(n42702) );
  NOR U63003 ( .A(n50337), .B(n42702), .Z(n45223) );
  XOR U63004 ( .A(n50339), .B(n45223), .Z(n42703) );
  IV U63005 ( .A(n42703), .Z(n47526) );
  XOR U63006 ( .A(n47525), .B(n47526), .Z(n45221) );
  IV U63007 ( .A(n45221), .Z(n42710) );
  IV U63008 ( .A(n42704), .Z(n42705) );
  NOR U63009 ( .A(n42706), .B(n42705), .Z(n47522) );
  NOR U63010 ( .A(n42708), .B(n42707), .Z(n45220) );
  NOR U63011 ( .A(n47522), .B(n45220), .Z(n42709) );
  XOR U63012 ( .A(n42710), .B(n42709), .Z(n47537) );
  XOR U63013 ( .A(n47533), .B(n47537), .Z(n45218) );
  XOR U63014 ( .A(n42711), .B(n45218), .Z(n45216) );
  XOR U63015 ( .A(n45214), .B(n45216), .Z(n45210) );
  IV U63016 ( .A(n45210), .Z(n42719) );
  IV U63017 ( .A(n42712), .Z(n42714) );
  NOR U63018 ( .A(n42714), .B(n42713), .Z(n45212) );
  IV U63019 ( .A(n42715), .Z(n42717) );
  NOR U63020 ( .A(n42717), .B(n42716), .Z(n45209) );
  NOR U63021 ( .A(n45212), .B(n45209), .Z(n42718) );
  XOR U63022 ( .A(n42719), .B(n42718), .Z(n45207) );
  IV U63023 ( .A(n42720), .Z(n42721) );
  NOR U63024 ( .A(n42722), .B(n42721), .Z(n45203) );
  NOR U63025 ( .A(n42724), .B(n42723), .Z(n45205) );
  NOR U63026 ( .A(n45203), .B(n45205), .Z(n42725) );
  XOR U63027 ( .A(n45207), .B(n42725), .Z(n45198) );
  IV U63028 ( .A(n42726), .Z(n42728) );
  NOR U63029 ( .A(n42728), .B(n42727), .Z(n45200) );
  IV U63030 ( .A(n42729), .Z(n42731) );
  NOR U63031 ( .A(n42731), .B(n42730), .Z(n45197) );
  NOR U63032 ( .A(n45200), .B(n45197), .Z(n42732) );
  XOR U63033 ( .A(n45198), .B(n42732), .Z(n47545) );
  IV U63034 ( .A(n42733), .Z(n42734) );
  NOR U63035 ( .A(n42735), .B(n42734), .Z(n47541) );
  NOR U63036 ( .A(n42737), .B(n42736), .Z(n47543) );
  NOR U63037 ( .A(n47541), .B(n47543), .Z(n42738) );
  XOR U63038 ( .A(n47545), .B(n42738), .Z(n47548) );
  IV U63039 ( .A(n42739), .Z(n42741) );
  NOR U63040 ( .A(n42741), .B(n42740), .Z(n52974) );
  IV U63041 ( .A(n42742), .Z(n42743) );
  NOR U63042 ( .A(n42744), .B(n42743), .Z(n50294) );
  NOR U63043 ( .A(n52974), .B(n50294), .Z(n47549) );
  XOR U63044 ( .A(n47548), .B(n47549), .Z(n47551) );
  XOR U63045 ( .A(n42745), .B(n47551), .Z(n45194) );
  NOR U63046 ( .A(n42746), .B(n45194), .Z(n42749) );
  IV U63047 ( .A(n42746), .Z(n42748) );
  XOR U63048 ( .A(n47550), .B(n47551), .Z(n42747) );
  NOR U63049 ( .A(n42748), .B(n42747), .Z(n52977) );
  NOR U63050 ( .A(n42749), .B(n52977), .Z(n45189) );
  XOR U63051 ( .A(n42750), .B(n45189), .Z(n50280) );
  XOR U63052 ( .A(n45187), .B(n50280), .Z(n42751) );
  IV U63053 ( .A(n42751), .Z(n45185) );
  XOR U63054 ( .A(n45182), .B(n45185), .Z(n45180) );
  XOR U63055 ( .A(n42752), .B(n45180), .Z(n45177) );
  XOR U63056 ( .A(n45178), .B(n45177), .Z(n50261) );
  XOR U63057 ( .A(n47561), .B(n50261), .Z(n47572) );
  IV U63058 ( .A(n42753), .Z(n42754) );
  NOR U63059 ( .A(n42755), .B(n42754), .Z(n47574) );
  IV U63060 ( .A(n42756), .Z(n42757) );
  NOR U63061 ( .A(n42758), .B(n42757), .Z(n47571) );
  NOR U63062 ( .A(n47574), .B(n47571), .Z(n42759) );
  XOR U63063 ( .A(n47572), .B(n42759), .Z(n47567) );
  XOR U63064 ( .A(n42760), .B(n47567), .Z(n47594) );
  XOR U63065 ( .A(n47592), .B(n47594), .Z(n47606) );
  IV U63066 ( .A(n47587), .Z(n47600) );
  NOR U63067 ( .A(n47600), .B(n47586), .Z(n42763) );
  NOR U63068 ( .A(n47599), .B(n42761), .Z(n42762) );
  NOR U63069 ( .A(n42763), .B(n42762), .Z(n42764) );
  XOR U63070 ( .A(n47606), .B(n42764), .Z(n47614) );
  IV U63071 ( .A(n42765), .Z(n42766) );
  NOR U63072 ( .A(n42767), .B(n42766), .Z(n47611) );
  IV U63073 ( .A(n42768), .Z(n42770) );
  NOR U63074 ( .A(n42770), .B(n42769), .Z(n47613) );
  NOR U63075 ( .A(n47611), .B(n47613), .Z(n42771) );
  XOR U63076 ( .A(n47614), .B(n42771), .Z(n45172) );
  IV U63077 ( .A(n42772), .Z(n42773) );
  NOR U63078 ( .A(n42774), .B(n42773), .Z(n47607) );
  IV U63079 ( .A(n42775), .Z(n42776) );
  NOR U63080 ( .A(n42777), .B(n42776), .Z(n45173) );
  NOR U63081 ( .A(n47607), .B(n45173), .Z(n42778) );
  XOR U63082 ( .A(n45172), .B(n42778), .Z(n47628) );
  IV U63083 ( .A(n42779), .Z(n42781) );
  NOR U63084 ( .A(n42781), .B(n42780), .Z(n47626) );
  IV U63085 ( .A(n42782), .Z(n42783) );
  NOR U63086 ( .A(n42784), .B(n42783), .Z(n47621) );
  NOR U63087 ( .A(n47626), .B(n47621), .Z(n45171) );
  XOR U63088 ( .A(n47628), .B(n45171), .Z(n45169) );
  XOR U63089 ( .A(n42785), .B(n45169), .Z(n47640) );
  IV U63090 ( .A(n42786), .Z(n42788) );
  NOR U63091 ( .A(n42788), .B(n42787), .Z(n47639) );
  IV U63092 ( .A(n42789), .Z(n42790) );
  NOR U63093 ( .A(n42791), .B(n42790), .Z(n45166) );
  NOR U63094 ( .A(n47639), .B(n45166), .Z(n42792) );
  XOR U63095 ( .A(n47640), .B(n42792), .Z(n42793) );
  IV U63096 ( .A(n42793), .Z(n45165) );
  XOR U63097 ( .A(n45161), .B(n45165), .Z(n42794) );
  NOR U63098 ( .A(n42795), .B(n42794), .Z(n45160) );
  IV U63099 ( .A(n42796), .Z(n42797) );
  NOR U63100 ( .A(n42798), .B(n42797), .Z(n45163) );
  NOR U63101 ( .A(n45161), .B(n45163), .Z(n42799) );
  XOR U63102 ( .A(n45165), .B(n42799), .Z(n47646) );
  NOR U63103 ( .A(n42800), .B(n47646), .Z(n42801) );
  NOR U63104 ( .A(n45160), .B(n42801), .Z(n45157) );
  IV U63105 ( .A(n42802), .Z(n42804) );
  NOR U63106 ( .A(n42804), .B(n42803), .Z(n47645) );
  IV U63107 ( .A(n42805), .Z(n42806) );
  NOR U63108 ( .A(n42807), .B(n42806), .Z(n45156) );
  NOR U63109 ( .A(n47645), .B(n45156), .Z(n42808) );
  XOR U63110 ( .A(n45157), .B(n42808), .Z(n50219) );
  XOR U63111 ( .A(n42809), .B(n50219), .Z(n47652) );
  XOR U63112 ( .A(n47651), .B(n47652), .Z(n47659) );
  IV U63113 ( .A(n42810), .Z(n42811) );
  NOR U63114 ( .A(n42812), .B(n42811), .Z(n47649) );
  IV U63115 ( .A(n42813), .Z(n42814) );
  NOR U63116 ( .A(n42815), .B(n42814), .Z(n47658) );
  NOR U63117 ( .A(n47649), .B(n47658), .Z(n42816) );
  XOR U63118 ( .A(n47659), .B(n42816), .Z(n47663) );
  IV U63119 ( .A(n42817), .Z(n42818) );
  NOR U63120 ( .A(n42819), .B(n42818), .Z(n58239) );
  IV U63121 ( .A(n42820), .Z(n42821) );
  NOR U63122 ( .A(n42822), .B(n42821), .Z(n55428) );
  NOR U63123 ( .A(n58239), .B(n55428), .Z(n47664) );
  XOR U63124 ( .A(n47663), .B(n47664), .Z(n47674) );
  IV U63125 ( .A(n42823), .Z(n42825) );
  NOR U63126 ( .A(n42825), .B(n42824), .Z(n47675) );
  IV U63127 ( .A(n42826), .Z(n42828) );
  NOR U63128 ( .A(n42828), .B(n42827), .Z(n47671) );
  NOR U63129 ( .A(n47675), .B(n47671), .Z(n42829) );
  XOR U63130 ( .A(n47674), .B(n42829), .Z(n47682) );
  IV U63131 ( .A(n42830), .Z(n42831) );
  NOR U63132 ( .A(n42832), .B(n42831), .Z(n47673) );
  IV U63133 ( .A(n42833), .Z(n42834) );
  NOR U63134 ( .A(n42835), .B(n42834), .Z(n47681) );
  NOR U63135 ( .A(n47673), .B(n47681), .Z(n42836) );
  XOR U63136 ( .A(n47682), .B(n42836), .Z(n47688) );
  IV U63137 ( .A(n42837), .Z(n42839) );
  NOR U63138 ( .A(n42839), .B(n42838), .Z(n47679) );
  IV U63139 ( .A(n42840), .Z(n42841) );
  NOR U63140 ( .A(n42842), .B(n42841), .Z(n47686) );
  NOR U63141 ( .A(n47679), .B(n47686), .Z(n42843) );
  XOR U63142 ( .A(n47688), .B(n42843), .Z(n47689) );
  XOR U63143 ( .A(n47690), .B(n47689), .Z(n55417) );
  IV U63144 ( .A(n42846), .Z(n42844) );
  NOR U63145 ( .A(n42845), .B(n42844), .Z(n42849) );
  IV U63146 ( .A(n42845), .Z(n42847) );
  NOR U63147 ( .A(n42847), .B(n42846), .Z(n58261) );
  NOR U63148 ( .A(n55409), .B(n58261), .Z(n42848) );
  NOR U63149 ( .A(n42849), .B(n42848), .Z(n47691) );
  XOR U63150 ( .A(n55417), .B(n47691), .Z(n47699) );
  IV U63151 ( .A(n42850), .Z(n42852) );
  NOR U63152 ( .A(n42852), .B(n42851), .Z(n47698) );
  IV U63153 ( .A(n42853), .Z(n42854) );
  NOR U63154 ( .A(n42855), .B(n42854), .Z(n47696) );
  NOR U63155 ( .A(n47698), .B(n47696), .Z(n42856) );
  XOR U63156 ( .A(n47699), .B(n42856), .Z(n45150) );
  XOR U63157 ( .A(n42857), .B(n45150), .Z(n45147) );
  IV U63158 ( .A(n42858), .Z(n42860) );
  NOR U63159 ( .A(n42860), .B(n42859), .Z(n45149) );
  IV U63160 ( .A(n42861), .Z(n42863) );
  NOR U63161 ( .A(n42863), .B(n42862), .Z(n45146) );
  NOR U63162 ( .A(n45149), .B(n45146), .Z(n42864) );
  XOR U63163 ( .A(n45147), .B(n42864), .Z(n45144) );
  IV U63164 ( .A(n42865), .Z(n42866) );
  NOR U63165 ( .A(n42867), .B(n42866), .Z(n50174) );
  IV U63166 ( .A(n42868), .Z(n42869) );
  NOR U63167 ( .A(n42870), .B(n42869), .Z(n50164) );
  NOR U63168 ( .A(n50174), .B(n50164), .Z(n45145) );
  XOR U63169 ( .A(n45144), .B(n45145), .Z(n50161) );
  IV U63170 ( .A(n42871), .Z(n42873) );
  NOR U63171 ( .A(n42873), .B(n42872), .Z(n50168) );
  IV U63172 ( .A(n42874), .Z(n42875) );
  NOR U63173 ( .A(n42876), .B(n42875), .Z(n50159) );
  NOR U63174 ( .A(n50168), .B(n50159), .Z(n47715) );
  XOR U63175 ( .A(n50161), .B(n47715), .Z(n45142) );
  XOR U63176 ( .A(n42877), .B(n45142), .Z(n47731) );
  IV U63177 ( .A(n42878), .Z(n42880) );
  NOR U63178 ( .A(n42880), .B(n42879), .Z(n47721) );
  IV U63179 ( .A(n42881), .Z(n42883) );
  NOR U63180 ( .A(n42883), .B(n42882), .Z(n47730) );
  NOR U63181 ( .A(n47721), .B(n47730), .Z(n42884) );
  XOR U63182 ( .A(n47731), .B(n42884), .Z(n47728) );
  XOR U63183 ( .A(n42885), .B(n47728), .Z(n47740) );
  XOR U63184 ( .A(n47739), .B(n47740), .Z(n42896) );
  IV U63185 ( .A(n42896), .Z(n42894) );
  IV U63186 ( .A(n42886), .Z(n42887) );
  NOR U63187 ( .A(n42888), .B(n42887), .Z(n42898) );
  IV U63188 ( .A(n42889), .Z(n42890) );
  NOR U63189 ( .A(n42891), .B(n42890), .Z(n42895) );
  NOR U63190 ( .A(n42898), .B(n42895), .Z(n42892) );
  IV U63191 ( .A(n42892), .Z(n42893) );
  NOR U63192 ( .A(n42894), .B(n42893), .Z(n42902) );
  IV U63193 ( .A(n42895), .Z(n42897) );
  NOR U63194 ( .A(n42897), .B(n42896), .Z(n45140) );
  IV U63195 ( .A(n42898), .Z(n42899) );
  NOR U63196 ( .A(n42899), .B(n47740), .Z(n53049) );
  NOR U63197 ( .A(n45140), .B(n53049), .Z(n42900) );
  IV U63198 ( .A(n42900), .Z(n42901) );
  NOR U63199 ( .A(n42902), .B(n42901), .Z(n47753) );
  IV U63200 ( .A(n42903), .Z(n42904) );
  NOR U63201 ( .A(n42905), .B(n42904), .Z(n58302) );
  IV U63202 ( .A(n42906), .Z(n42908) );
  NOR U63203 ( .A(n42908), .B(n42907), .Z(n58297) );
  NOR U63204 ( .A(n58302), .B(n58297), .Z(n50158) );
  XOR U63205 ( .A(n47753), .B(n50158), .Z(n47759) );
  IV U63206 ( .A(n42909), .Z(n42911) );
  NOR U63207 ( .A(n42911), .B(n42910), .Z(n47754) );
  IV U63208 ( .A(n42912), .Z(n42913) );
  NOR U63209 ( .A(n42914), .B(n42913), .Z(n47758) );
  NOR U63210 ( .A(n47754), .B(n47758), .Z(n42915) );
  XOR U63211 ( .A(n47759), .B(n42915), .Z(n45134) );
  IV U63212 ( .A(n42916), .Z(n42917) );
  NOR U63213 ( .A(n42918), .B(n42917), .Z(n45137) );
  IV U63214 ( .A(n42919), .Z(n42921) );
  NOR U63215 ( .A(n42921), .B(n42920), .Z(n45135) );
  NOR U63216 ( .A(n45137), .B(n45135), .Z(n42922) );
  XOR U63217 ( .A(n45134), .B(n42922), .Z(n47765) );
  IV U63218 ( .A(n42923), .Z(n42924) );
  NOR U63219 ( .A(n42925), .B(n42924), .Z(n45132) );
  IV U63220 ( .A(n42926), .Z(n42928) );
  NOR U63221 ( .A(n42928), .B(n42927), .Z(n53075) );
  NOR U63222 ( .A(n45132), .B(n53075), .Z(n42929) );
  XOR U63223 ( .A(n47765), .B(n42929), .Z(n45127) );
  IV U63224 ( .A(n42930), .Z(n42931) );
  NOR U63225 ( .A(n42932), .B(n42931), .Z(n47762) );
  IV U63226 ( .A(n42933), .Z(n42935) );
  NOR U63227 ( .A(n42935), .B(n42934), .Z(n45130) );
  NOR U63228 ( .A(n47762), .B(n45130), .Z(n42936) );
  XOR U63229 ( .A(n45127), .B(n42936), .Z(n45124) );
  IV U63230 ( .A(n42937), .Z(n42939) );
  NOR U63231 ( .A(n42939), .B(n42938), .Z(n45126) );
  IV U63232 ( .A(n42940), .Z(n42941) );
  NOR U63233 ( .A(n42942), .B(n42941), .Z(n45123) );
  NOR U63234 ( .A(n45126), .B(n45123), .Z(n42943) );
  XOR U63235 ( .A(n45124), .B(n42943), .Z(n45118) );
  XOR U63236 ( .A(n45119), .B(n45118), .Z(n42944) );
  NOR U63237 ( .A(n42945), .B(n42944), .Z(n45117) );
  IV U63238 ( .A(n42946), .Z(n42947) );
  NOR U63239 ( .A(n42948), .B(n42947), .Z(n45120) );
  NOR U63240 ( .A(n42949), .B(n45120), .Z(n42950) );
  XOR U63241 ( .A(n45118), .B(n42950), .Z(n42959) );
  IV U63242 ( .A(n42959), .Z(n42951) );
  NOR U63243 ( .A(n42952), .B(n42951), .Z(n42953) );
  NOR U63244 ( .A(n45117), .B(n42953), .Z(n42966) );
  IV U63245 ( .A(n42966), .Z(n42954) );
  NOR U63246 ( .A(n42955), .B(n42954), .Z(n53093) );
  IV U63247 ( .A(n42956), .Z(n42957) );
  NOR U63248 ( .A(n42958), .B(n42957), .Z(n42962) );
  IV U63249 ( .A(n42962), .Z(n42960) );
  NOR U63250 ( .A(n42960), .B(n42959), .Z(n53089) );
  NOR U63251 ( .A(n53093), .B(n53089), .Z(n42961) );
  IV U63252 ( .A(n42961), .Z(n47780) );
  NOR U63253 ( .A(n42963), .B(n42962), .Z(n42964) );
  IV U63254 ( .A(n42964), .Z(n42965) );
  NOR U63255 ( .A(n42966), .B(n42965), .Z(n42967) );
  NOR U63256 ( .A(n47780), .B(n42967), .Z(n47774) );
  XOR U63257 ( .A(n47775), .B(n47774), .Z(n47770) );
  IV U63258 ( .A(n42968), .Z(n42969) );
  NOR U63259 ( .A(n42970), .B(n42969), .Z(n47776) );
  IV U63260 ( .A(n42971), .Z(n42973) );
  NOR U63261 ( .A(n42973), .B(n42972), .Z(n47769) );
  NOR U63262 ( .A(n47776), .B(n47769), .Z(n42974) );
  XOR U63263 ( .A(n47770), .B(n42974), .Z(n45112) );
  XOR U63264 ( .A(n45113), .B(n45112), .Z(n45115) );
  NOR U63265 ( .A(n42981), .B(n45115), .Z(n50124) );
  IV U63266 ( .A(n42975), .Z(n42976) );
  NOR U63267 ( .A(n42977), .B(n42976), .Z(n45109) );
  IV U63268 ( .A(n42978), .Z(n42979) );
  NOR U63269 ( .A(n42980), .B(n42979), .Z(n45114) );
  XOR U63270 ( .A(n45114), .B(n45115), .Z(n45110) );
  IV U63271 ( .A(n45110), .Z(n42982) );
  XOR U63272 ( .A(n45109), .B(n42982), .Z(n42984) );
  NOR U63273 ( .A(n42982), .B(n42981), .Z(n42983) );
  NOR U63274 ( .A(n42984), .B(n42983), .Z(n42985) );
  NOR U63275 ( .A(n50124), .B(n42985), .Z(n45106) );
  IV U63276 ( .A(n42986), .Z(n42987) );
  NOR U63277 ( .A(n42988), .B(n42987), .Z(n42989) );
  IV U63278 ( .A(n42989), .Z(n45108) );
  XOR U63279 ( .A(n45106), .B(n45108), .Z(n45103) );
  NOR U63280 ( .A(n42996), .B(n45103), .Z(n50113) );
  IV U63281 ( .A(n42990), .Z(n42992) );
  NOR U63282 ( .A(n42992), .B(n42991), .Z(n47788) );
  IV U63283 ( .A(n42993), .Z(n42994) );
  NOR U63284 ( .A(n42995), .B(n42994), .Z(n45102) );
  XOR U63285 ( .A(n45102), .B(n45103), .Z(n47789) );
  IV U63286 ( .A(n47789), .Z(n42997) );
  XOR U63287 ( .A(n47788), .B(n42997), .Z(n42999) );
  NOR U63288 ( .A(n42997), .B(n42996), .Z(n42998) );
  NOR U63289 ( .A(n42999), .B(n42998), .Z(n43000) );
  NOR U63290 ( .A(n50113), .B(n43000), .Z(n47791) );
  IV U63291 ( .A(n43001), .Z(n43002) );
  NOR U63292 ( .A(n43003), .B(n43002), .Z(n53111) );
  IV U63293 ( .A(n43004), .Z(n43005) );
  NOR U63294 ( .A(n43006), .B(n43005), .Z(n53119) );
  NOR U63295 ( .A(n53111), .B(n53119), .Z(n47792) );
  XOR U63296 ( .A(n47791), .B(n47792), .Z(n47798) );
  XOR U63297 ( .A(n43007), .B(n47798), .Z(n45095) );
  IV U63298 ( .A(n43008), .Z(n43010) );
  NOR U63299 ( .A(n43010), .B(n43009), .Z(n45098) );
  IV U63300 ( .A(n43011), .Z(n43012) );
  NOR U63301 ( .A(n43013), .B(n43012), .Z(n45094) );
  NOR U63302 ( .A(n45098), .B(n45094), .Z(n43014) );
  XOR U63303 ( .A(n45095), .B(n43014), .Z(n47806) );
  XOR U63304 ( .A(n47805), .B(n47806), .Z(n45091) );
  IV U63305 ( .A(n43015), .Z(n43017) );
  NOR U63306 ( .A(n43017), .B(n43016), .Z(n47802) );
  IV U63307 ( .A(n43018), .Z(n43020) );
  NOR U63308 ( .A(n43020), .B(n43019), .Z(n45090) );
  NOR U63309 ( .A(n47802), .B(n45090), .Z(n43021) );
  XOR U63310 ( .A(n45091), .B(n43021), .Z(n55315) );
  XOR U63311 ( .A(n45089), .B(n55315), .Z(n45087) );
  XOR U63312 ( .A(n45088), .B(n45087), .Z(n47824) );
  IV U63313 ( .A(n47824), .Z(n43028) );
  IV U63314 ( .A(n43022), .Z(n43024) );
  NOR U63315 ( .A(n43024), .B(n43023), .Z(n55304) );
  IV U63316 ( .A(n43025), .Z(n43026) );
  NOR U63317 ( .A(n43027), .B(n43026), .Z(n55296) );
  NOR U63318 ( .A(n55304), .B(n55296), .Z(n47825) );
  XOR U63319 ( .A(n43028), .B(n47825), .Z(n47820) );
  XOR U63320 ( .A(n47817), .B(n47820), .Z(n47840) );
  XOR U63321 ( .A(n43029), .B(n47840), .Z(n47836) );
  XOR U63322 ( .A(n43030), .B(n47836), .Z(n47847) );
  XOR U63323 ( .A(n47848), .B(n47847), .Z(n43042) );
  IV U63324 ( .A(n43042), .Z(n43031) );
  NOR U63325 ( .A(n43032), .B(n43031), .Z(n53171) );
  IV U63326 ( .A(n43033), .Z(n43034) );
  NOR U63327 ( .A(n43035), .B(n43034), .Z(n43038) );
  IV U63328 ( .A(n43038), .Z(n43036) );
  NOR U63329 ( .A(n43036), .B(n47847), .Z(n53164) );
  NOR U63330 ( .A(n53171), .B(n53164), .Z(n43037) );
  IV U63331 ( .A(n43037), .Z(n47849) );
  NOR U63332 ( .A(n43039), .B(n43038), .Z(n43040) );
  IV U63333 ( .A(n43040), .Z(n43041) );
  NOR U63334 ( .A(n43042), .B(n43041), .Z(n43043) );
  NOR U63335 ( .A(n47849), .B(n43043), .Z(n43044) );
  IV U63336 ( .A(n43044), .Z(n47856) );
  XOR U63337 ( .A(n47855), .B(n47856), .Z(n47862) );
  IV U63338 ( .A(n47862), .Z(n43052) );
  IV U63339 ( .A(n43045), .Z(n43047) );
  NOR U63340 ( .A(n43047), .B(n43046), .Z(n47852) );
  IV U63341 ( .A(n43048), .Z(n43049) );
  NOR U63342 ( .A(n43050), .B(n43049), .Z(n47861) );
  NOR U63343 ( .A(n47852), .B(n47861), .Z(n43051) );
  XOR U63344 ( .A(n43052), .B(n43051), .Z(n47869) );
  XOR U63345 ( .A(n47865), .B(n47869), .Z(n47875) );
  XOR U63346 ( .A(n43053), .B(n47875), .Z(n47871) );
  IV U63347 ( .A(n43054), .Z(n43055) );
  NOR U63348 ( .A(n43056), .B(n43055), .Z(n47872) );
  IV U63349 ( .A(n43057), .Z(n43059) );
  NOR U63350 ( .A(n43059), .B(n43058), .Z(n47878) );
  NOR U63351 ( .A(n47872), .B(n47878), .Z(n43060) );
  XOR U63352 ( .A(n47871), .B(n43060), .Z(n45084) );
  XOR U63353 ( .A(n45083), .B(n45084), .Z(n47885) );
  XOR U63354 ( .A(n43061), .B(n47885), .Z(n47882) );
  XOR U63355 ( .A(n47883), .B(n47882), .Z(n45079) );
  XOR U63356 ( .A(n45078), .B(n45079), .Z(n45074) );
  XOR U63357 ( .A(n43062), .B(n45074), .Z(n45071) );
  XOR U63358 ( .A(n45072), .B(n45071), .Z(n45069) );
  XOR U63359 ( .A(n43063), .B(n45069), .Z(n47895) );
  NOR U63360 ( .A(n43064), .B(n47895), .Z(n43067) );
  IV U63361 ( .A(n43064), .Z(n43066) );
  XOR U63362 ( .A(n45068), .B(n45069), .Z(n43065) );
  NOR U63363 ( .A(n43066), .B(n43065), .Z(n50071) );
  NOR U63364 ( .A(n43067), .B(n50071), .Z(n47900) );
  IV U63365 ( .A(n43068), .Z(n43069) );
  NOR U63366 ( .A(n43070), .B(n43069), .Z(n47894) );
  IV U63367 ( .A(n43071), .Z(n43073) );
  NOR U63368 ( .A(n43073), .B(n43072), .Z(n47899) );
  NOR U63369 ( .A(n47894), .B(n47899), .Z(n43074) );
  XOR U63370 ( .A(n47900), .B(n43074), .Z(n47905) );
  IV U63371 ( .A(n43078), .Z(n43075) );
  NOR U63372 ( .A(n43075), .B(n43076), .Z(n47903) );
  IV U63373 ( .A(n43076), .Z(n43077) );
  NOR U63374 ( .A(n43078), .B(n43077), .Z(n43080) );
  IV U63375 ( .A(n43079), .Z(n45063) );
  NOR U63376 ( .A(n43080), .B(n45063), .Z(n43081) );
  NOR U63377 ( .A(n47903), .B(n43081), .Z(n43082) );
  XOR U63378 ( .A(n47905), .B(n43082), .Z(n47908) );
  IV U63379 ( .A(n43083), .Z(n43084) );
  NOR U63380 ( .A(n43085), .B(n43084), .Z(n45059) );
  IV U63381 ( .A(n43086), .Z(n43087) );
  NOR U63382 ( .A(n43088), .B(n43087), .Z(n47910) );
  NOR U63383 ( .A(n45059), .B(n47910), .Z(n43089) );
  XOR U63384 ( .A(n47908), .B(n43089), .Z(n45056) );
  XOR U63385 ( .A(n43090), .B(n45056), .Z(n45053) );
  XOR U63386 ( .A(n45054), .B(n45053), .Z(n47919) );
  XOR U63387 ( .A(n47916), .B(n47919), .Z(n43091) );
  NOR U63388 ( .A(n43092), .B(n43091), .Z(n47923) );
  IV U63389 ( .A(n43093), .Z(n43095) );
  NOR U63390 ( .A(n43095), .B(n43094), .Z(n47918) );
  NOR U63391 ( .A(n47916), .B(n47918), .Z(n43096) );
  XOR U63392 ( .A(n43096), .B(n47919), .Z(n43100) );
  NOR U63393 ( .A(n43097), .B(n43100), .Z(n43098) );
  NOR U63394 ( .A(n47923), .B(n43098), .Z(n47926) );
  NOR U63395 ( .A(n43099), .B(n47926), .Z(n43103) );
  IV U63396 ( .A(n43099), .Z(n43102) );
  IV U63397 ( .A(n43100), .Z(n43101) );
  NOR U63398 ( .A(n43102), .B(n43101), .Z(n50050) );
  NOR U63399 ( .A(n43103), .B(n50050), .Z(n47934) );
  XOR U63400 ( .A(n43104), .B(n47934), .Z(n47932) );
  IV U63401 ( .A(n43105), .Z(n43106) );
  NOR U63402 ( .A(n43107), .B(n43106), .Z(n47930) );
  IV U63403 ( .A(n43108), .Z(n43109) );
  NOR U63404 ( .A(n43110), .B(n43109), .Z(n45051) );
  NOR U63405 ( .A(n47930), .B(n45051), .Z(n43111) );
  XOR U63406 ( .A(n47932), .B(n43111), .Z(n43112) );
  IV U63407 ( .A(n43112), .Z(n47946) );
  XOR U63408 ( .A(n43113), .B(n47946), .Z(n45044) );
  IV U63409 ( .A(n43114), .Z(n43116) );
  NOR U63410 ( .A(n43116), .B(n43115), .Z(n45047) );
  IV U63411 ( .A(n43117), .Z(n43118) );
  NOR U63412 ( .A(n43119), .B(n43118), .Z(n45043) );
  NOR U63413 ( .A(n45047), .B(n45043), .Z(n43120) );
  XOR U63414 ( .A(n45044), .B(n43120), .Z(n47956) );
  IV U63415 ( .A(n43121), .Z(n43122) );
  NOR U63416 ( .A(n43123), .B(n43122), .Z(n47950) );
  IV U63417 ( .A(n43124), .Z(n43126) );
  NOR U63418 ( .A(n43126), .B(n43125), .Z(n47954) );
  NOR U63419 ( .A(n47950), .B(n47954), .Z(n43127) );
  XOR U63420 ( .A(n47956), .B(n43127), .Z(n45037) );
  IV U63421 ( .A(n43128), .Z(n43130) );
  NOR U63422 ( .A(n43130), .B(n43129), .Z(n45040) );
  IV U63423 ( .A(n43131), .Z(n43133) );
  NOR U63424 ( .A(n43133), .B(n43132), .Z(n45036) );
  NOR U63425 ( .A(n45040), .B(n45036), .Z(n43134) );
  XOR U63426 ( .A(n45037), .B(n43134), .Z(n47967) );
  IV U63427 ( .A(n43135), .Z(n43136) );
  NOR U63428 ( .A(n43137), .B(n43136), .Z(n47965) );
  IV U63429 ( .A(n43138), .Z(n43139) );
  NOR U63430 ( .A(n43140), .B(n43139), .Z(n47962) );
  NOR U63431 ( .A(n47965), .B(n47962), .Z(n43141) );
  XOR U63432 ( .A(n47967), .B(n43141), .Z(n45028) );
  IV U63433 ( .A(n43142), .Z(n43144) );
  NOR U63434 ( .A(n43144), .B(n43143), .Z(n45033) );
  IV U63435 ( .A(n43145), .Z(n43146) );
  NOR U63436 ( .A(n43147), .B(n43146), .Z(n45027) );
  NOR U63437 ( .A(n45033), .B(n45027), .Z(n43148) );
  XOR U63438 ( .A(n45028), .B(n43148), .Z(n45031) );
  XOR U63439 ( .A(n45030), .B(n45031), .Z(n47973) );
  XOR U63440 ( .A(n43149), .B(n47973), .Z(n47970) );
  XOR U63441 ( .A(n47971), .B(n47970), .Z(n47981) );
  XOR U63442 ( .A(n43150), .B(n47981), .Z(n43151) );
  NOR U63443 ( .A(n47978), .B(n43151), .Z(n43154) );
  IV U63444 ( .A(n47978), .Z(n47982) );
  XOR U63445 ( .A(n47977), .B(n47981), .Z(n43152) );
  NOR U63446 ( .A(n47982), .B(n43152), .Z(n43153) );
  NOR U63447 ( .A(n43154), .B(n43153), .Z(n47992) );
  XOR U63448 ( .A(n43155), .B(n47992), .Z(n48010) );
  IV U63449 ( .A(n48010), .Z(n43163) );
  IV U63450 ( .A(n43156), .Z(n43158) );
  NOR U63451 ( .A(n43158), .B(n43157), .Z(n48009) );
  IV U63452 ( .A(n43159), .Z(n43161) );
  NOR U63453 ( .A(n43161), .B(n43160), .Z(n45020) );
  NOR U63454 ( .A(n48009), .B(n45020), .Z(n43162) );
  XOR U63455 ( .A(n43163), .B(n43162), .Z(n48022) );
  XOR U63456 ( .A(n48021), .B(n48022), .Z(n45018) );
  XOR U63457 ( .A(n43164), .B(n45018), .Z(n48034) );
  IV U63458 ( .A(n43165), .Z(n43166) );
  NOR U63459 ( .A(n43167), .B(n43166), .Z(n48035) );
  IV U63460 ( .A(n43168), .Z(n43169) );
  NOR U63461 ( .A(n43170), .B(n43169), .Z(n48037) );
  NOR U63462 ( .A(n48035), .B(n48037), .Z(n43171) );
  XOR U63463 ( .A(n48034), .B(n43171), .Z(n55188) );
  XOR U63464 ( .A(n48041), .B(n55188), .Z(n45015) );
  XOR U63465 ( .A(n45016), .B(n45015), .Z(n48051) );
  XOR U63466 ( .A(n48063), .B(n48051), .Z(n48057) );
  XOR U63467 ( .A(n48056), .B(n48057), .Z(n48077) );
  XOR U63468 ( .A(n43172), .B(n48077), .Z(n48086) );
  XOR U63469 ( .A(n48087), .B(n48086), .Z(n48082) );
  XOR U63470 ( .A(n48079), .B(n48082), .Z(n45010) );
  XOR U63471 ( .A(n43173), .B(n45010), .Z(n45007) );
  XOR U63472 ( .A(n45008), .B(n45007), .Z(n48099) );
  XOR U63473 ( .A(n43174), .B(n48099), .Z(n48095) );
  IV U63474 ( .A(n43175), .Z(n43177) );
  NOR U63475 ( .A(n43177), .B(n43176), .Z(n48096) );
  IV U63476 ( .A(n43178), .Z(n43179) );
  NOR U63477 ( .A(n43180), .B(n43179), .Z(n48105) );
  NOR U63478 ( .A(n48096), .B(n48105), .Z(n43181) );
  XOR U63479 ( .A(n48095), .B(n43181), .Z(n48103) );
  XOR U63480 ( .A(n48102), .B(n48103), .Z(n45001) );
  NOR U63481 ( .A(n43188), .B(n45001), .Z(n58536) );
  IV U63482 ( .A(n43182), .Z(n43183) );
  NOR U63483 ( .A(n43184), .B(n43183), .Z(n44997) );
  IV U63484 ( .A(n43185), .Z(n43187) );
  NOR U63485 ( .A(n43187), .B(n43186), .Z(n45000) );
  XOR U63486 ( .A(n45000), .B(n45001), .Z(n44998) );
  IV U63487 ( .A(n44998), .Z(n43189) );
  XOR U63488 ( .A(n44997), .B(n43189), .Z(n43191) );
  NOR U63489 ( .A(n43189), .B(n43188), .Z(n43190) );
  NOR U63490 ( .A(n43191), .B(n43190), .Z(n43192) );
  NOR U63491 ( .A(n58536), .B(n43192), .Z(n44990) );
  XOR U63492 ( .A(n43193), .B(n44990), .Z(n49979) );
  IV U63493 ( .A(n43194), .Z(n43196) );
  NOR U63494 ( .A(n43196), .B(n43195), .Z(n49983) );
  IV U63495 ( .A(n43197), .Z(n43198) );
  NOR U63496 ( .A(n43199), .B(n43198), .Z(n49978) );
  NOR U63497 ( .A(n49983), .B(n49978), .Z(n44988) );
  XOR U63498 ( .A(n49979), .B(n44988), .Z(n44986) );
  XOR U63499 ( .A(n43200), .B(n44986), .Z(n49969) );
  IV U63500 ( .A(n49969), .Z(n44980) );
  XOR U63501 ( .A(n44978), .B(n44980), .Z(n48116) );
  IV U63502 ( .A(n43201), .Z(n43203) );
  NOR U63503 ( .A(n43203), .B(n43202), .Z(n44981) );
  IV U63504 ( .A(n43204), .Z(n43206) );
  NOR U63505 ( .A(n43206), .B(n43205), .Z(n48115) );
  NOR U63506 ( .A(n44981), .B(n48115), .Z(n43207) );
  XOR U63507 ( .A(n48116), .B(n43207), .Z(n44976) );
  XOR U63508 ( .A(n44977), .B(n44976), .Z(n44974) );
  XOR U63509 ( .A(n43208), .B(n44974), .Z(n44969) );
  XOR U63510 ( .A(n44970), .B(n44969), .Z(n53325) );
  XOR U63511 ( .A(n48145), .B(n53325), .Z(n48143) );
  IV U63512 ( .A(n43209), .Z(n43211) );
  NOR U63513 ( .A(n43211), .B(n43210), .Z(n49956) );
  IV U63514 ( .A(n43212), .Z(n43213) );
  NOR U63515 ( .A(n43214), .B(n43213), .Z(n49951) );
  NOR U63516 ( .A(n49956), .B(n49951), .Z(n48144) );
  XOR U63517 ( .A(n48143), .B(n48144), .Z(n44967) );
  XOR U63518 ( .A(n43215), .B(n44967), .Z(n48147) );
  IV U63519 ( .A(n43216), .Z(n43218) );
  NOR U63520 ( .A(n43218), .B(n43217), .Z(n53337) );
  IV U63521 ( .A(n43219), .Z(n43220) );
  NOR U63522 ( .A(n43221), .B(n43220), .Z(n53343) );
  NOR U63523 ( .A(n53337), .B(n53343), .Z(n48148) );
  XOR U63524 ( .A(n48147), .B(n48148), .Z(n49943) );
  XOR U63525 ( .A(n48149), .B(n49943), .Z(n44962) );
  IV U63526 ( .A(n43222), .Z(n43223) );
  NOR U63527 ( .A(n43224), .B(n43223), .Z(n58614) );
  IV U63528 ( .A(n43225), .Z(n43226) );
  NOR U63529 ( .A(n43227), .B(n43226), .Z(n55081) );
  NOR U63530 ( .A(n58614), .B(n55081), .Z(n44963) );
  XOR U63531 ( .A(n44962), .B(n44963), .Z(n48161) );
  XOR U63532 ( .A(n43228), .B(n48161), .Z(n44960) );
  NOR U63533 ( .A(n43229), .B(n44955), .Z(n48153) );
  NOR U63534 ( .A(n44956), .B(n43230), .Z(n43232) );
  IV U63535 ( .A(n43231), .Z(n44958) );
  NOR U63536 ( .A(n43232), .B(n44958), .Z(n43233) );
  NOR U63537 ( .A(n48153), .B(n43233), .Z(n43234) );
  XOR U63538 ( .A(n44960), .B(n43234), .Z(n48177) );
  IV U63539 ( .A(n48177), .Z(n48176) );
  XOR U63540 ( .A(n48178), .B(n48176), .Z(n44953) );
  IV U63541 ( .A(n43235), .Z(n43236) );
  NOR U63542 ( .A(n43237), .B(n43236), .Z(n48179) );
  IV U63543 ( .A(n43238), .Z(n43239) );
  NOR U63544 ( .A(n43240), .B(n43239), .Z(n44952) );
  NOR U63545 ( .A(n48179), .B(n44952), .Z(n43241) );
  XOR U63546 ( .A(n44953), .B(n43241), .Z(n44950) );
  XOR U63547 ( .A(n44951), .B(n44950), .Z(n48186) );
  XOR U63548 ( .A(n43242), .B(n48186), .Z(n44947) );
  IV U63549 ( .A(n43243), .Z(n43245) );
  NOR U63550 ( .A(n43245), .B(n43244), .Z(n44946) );
  IV U63551 ( .A(n43246), .Z(n43247) );
  NOR U63552 ( .A(n43248), .B(n43247), .Z(n48194) );
  NOR U63553 ( .A(n44946), .B(n48194), .Z(n43249) );
  XOR U63554 ( .A(n44947), .B(n43249), .Z(n44944) );
  NOR U63555 ( .A(n43256), .B(n44944), .Z(n53376) );
  IV U63556 ( .A(n43250), .Z(n43251) );
  NOR U63557 ( .A(n43252), .B(n43251), .Z(n48199) );
  IV U63558 ( .A(n43253), .Z(n43255) );
  NOR U63559 ( .A(n43255), .B(n43254), .Z(n44943) );
  XOR U63560 ( .A(n44943), .B(n44944), .Z(n48200) );
  IV U63561 ( .A(n48200), .Z(n43257) );
  XOR U63562 ( .A(n48199), .B(n43257), .Z(n43259) );
  NOR U63563 ( .A(n43257), .B(n43256), .Z(n43258) );
  NOR U63564 ( .A(n43259), .B(n43258), .Z(n43260) );
  NOR U63565 ( .A(n53376), .B(n43260), .Z(n44939) );
  XOR U63566 ( .A(n43261), .B(n44939), .Z(n49906) );
  IV U63567 ( .A(n49906), .Z(n43267) );
  NOR U63568 ( .A(n43263), .B(n43262), .Z(n49909) );
  IV U63569 ( .A(n43264), .Z(n43266) );
  NOR U63570 ( .A(n43266), .B(n43265), .Z(n49904) );
  NOR U63571 ( .A(n49909), .B(n49904), .Z(n44941) );
  XOR U63572 ( .A(n43267), .B(n44941), .Z(n44936) );
  XOR U63573 ( .A(n44933), .B(n44936), .Z(n44931) );
  XOR U63574 ( .A(n43268), .B(n44931), .Z(n48208) );
  IV U63575 ( .A(n43269), .Z(n43271) );
  NOR U63576 ( .A(n43271), .B(n43270), .Z(n48214) );
  IV U63577 ( .A(n43272), .Z(n43273) );
  NOR U63578 ( .A(n43274), .B(n43273), .Z(n48209) );
  NOR U63579 ( .A(n48214), .B(n48209), .Z(n43275) );
  XOR U63580 ( .A(n48208), .B(n43275), .Z(n48223) );
  XOR U63581 ( .A(n43276), .B(n48223), .Z(n48225) );
  XOR U63582 ( .A(n48226), .B(n48225), .Z(n44928) );
  IV U63583 ( .A(n43277), .Z(n43279) );
  NOR U63584 ( .A(n43279), .B(n43278), .Z(n48228) );
  IV U63585 ( .A(n43280), .Z(n43281) );
  NOR U63586 ( .A(n43282), .B(n43281), .Z(n44927) );
  NOR U63587 ( .A(n48228), .B(n44927), .Z(n43283) );
  XOR U63588 ( .A(n44928), .B(n43283), .Z(n44923) );
  IV U63589 ( .A(n44923), .Z(n55042) );
  NOR U63590 ( .A(n43285), .B(n43284), .Z(n55037) );
  IV U63591 ( .A(n43286), .Z(n43288) );
  NOR U63592 ( .A(n43288), .B(n43287), .Z(n58679) );
  NOR U63593 ( .A(n55037), .B(n58679), .Z(n53389) );
  IV U63594 ( .A(n53389), .Z(n44922) );
  XOR U63595 ( .A(n55042), .B(n44922), .Z(n49877) );
  IV U63596 ( .A(n43289), .Z(n43290) );
  NOR U63597 ( .A(n43291), .B(n43290), .Z(n49875) );
  IV U63598 ( .A(n43292), .Z(n43293) );
  NOR U63599 ( .A(n43294), .B(n43293), .Z(n53396) );
  NOR U63600 ( .A(n49875), .B(n53396), .Z(n43295) );
  IV U63601 ( .A(n43295), .Z(n44924) );
  XOR U63602 ( .A(n49877), .B(n44924), .Z(n44921) );
  IV U63603 ( .A(n43296), .Z(n43297) );
  NOR U63604 ( .A(n43298), .B(n43297), .Z(n44919) );
  IV U63605 ( .A(n43299), .Z(n43300) );
  NOR U63606 ( .A(n43301), .B(n43300), .Z(n44917) );
  NOR U63607 ( .A(n44919), .B(n44917), .Z(n43302) );
  XOR U63608 ( .A(n44921), .B(n43302), .Z(n44911) );
  IV U63609 ( .A(n43303), .Z(n43305) );
  NOR U63610 ( .A(n43305), .B(n43304), .Z(n44914) );
  IV U63611 ( .A(n43306), .Z(n43307) );
  NOR U63612 ( .A(n43308), .B(n43307), .Z(n44910) );
  NOR U63613 ( .A(n44914), .B(n44910), .Z(n43309) );
  XOR U63614 ( .A(n44911), .B(n43309), .Z(n49867) );
  IV U63615 ( .A(n43310), .Z(n43311) );
  NOR U63616 ( .A(n43312), .B(n43311), .Z(n49870) );
  IV U63617 ( .A(n43313), .Z(n43314) );
  NOR U63618 ( .A(n43315), .B(n43314), .Z(n49865) );
  NOR U63619 ( .A(n49870), .B(n49865), .Z(n44897) );
  XOR U63620 ( .A(n49867), .B(n44897), .Z(n44899) );
  NOR U63621 ( .A(n43316), .B(n44902), .Z(n44898) );
  IV U63622 ( .A(n44902), .Z(n43317) );
  NOR U63623 ( .A(n44903), .B(n43317), .Z(n43318) );
  NOR U63624 ( .A(n43318), .B(n44905), .Z(n43319) );
  NOR U63625 ( .A(n44898), .B(n43319), .Z(n43320) );
  XOR U63626 ( .A(n44899), .B(n43320), .Z(n44896) );
  XOR U63627 ( .A(n44892), .B(n44896), .Z(n43321) );
  NOR U63628 ( .A(n43322), .B(n43321), .Z(n49851) );
  IV U63629 ( .A(n43323), .Z(n43324) );
  NOR U63630 ( .A(n43325), .B(n43324), .Z(n44894) );
  NOR U63631 ( .A(n44892), .B(n44894), .Z(n43326) );
  XOR U63632 ( .A(n44896), .B(n43326), .Z(n44889) );
  NOR U63633 ( .A(n43327), .B(n44889), .Z(n43328) );
  NOR U63634 ( .A(n49851), .B(n43328), .Z(n48241) );
  IV U63635 ( .A(n43329), .Z(n43330) );
  NOR U63636 ( .A(n43331), .B(n43330), .Z(n44888) );
  IV U63637 ( .A(n43332), .Z(n43334) );
  NOR U63638 ( .A(n43334), .B(n43333), .Z(n48240) );
  NOR U63639 ( .A(n44888), .B(n48240), .Z(n43335) );
  XOR U63640 ( .A(n48241), .B(n43335), .Z(n48239) );
  IV U63641 ( .A(n43336), .Z(n43338) );
  NOR U63642 ( .A(n43338), .B(n43337), .Z(n48237) );
  IV U63643 ( .A(n43339), .Z(n43341) );
  NOR U63644 ( .A(n43341), .B(n43340), .Z(n44886) );
  NOR U63645 ( .A(n48237), .B(n44886), .Z(n43342) );
  XOR U63646 ( .A(n48239), .B(n43342), .Z(n44880) );
  IV U63647 ( .A(n43343), .Z(n43344) );
  NOR U63648 ( .A(n43345), .B(n43344), .Z(n44882) );
  IV U63649 ( .A(n43346), .Z(n43348) );
  NOR U63650 ( .A(n43348), .B(n43347), .Z(n44879) );
  NOR U63651 ( .A(n44882), .B(n44879), .Z(n43349) );
  XOR U63652 ( .A(n44880), .B(n43349), .Z(n44878) );
  IV U63653 ( .A(n43350), .Z(n43351) );
  NOR U63654 ( .A(n43352), .B(n43351), .Z(n43371) );
  IV U63655 ( .A(n43353), .Z(n43354) );
  NOR U63656 ( .A(n43355), .B(n43354), .Z(n43370) );
  NOR U63657 ( .A(n43371), .B(n43370), .Z(n43356) );
  XOR U63658 ( .A(n44878), .B(n43356), .Z(n43366) );
  IV U63659 ( .A(n43357), .Z(n43359) );
  NOR U63660 ( .A(n43359), .B(n43358), .Z(n43369) );
  IV U63661 ( .A(n43360), .Z(n43362) );
  NOR U63662 ( .A(n43362), .B(n43361), .Z(n43365) );
  NOR U63663 ( .A(n43369), .B(n43365), .Z(n43363) );
  IV U63664 ( .A(n43363), .Z(n43364) );
  NOR U63665 ( .A(n43366), .B(n43364), .Z(n43377) );
  IV U63666 ( .A(n43365), .Z(n43368) );
  IV U63667 ( .A(n43366), .Z(n43367) );
  NOR U63668 ( .A(n43368), .B(n43367), .Z(n48249) );
  IV U63669 ( .A(n43369), .Z(n43375) );
  IV U63670 ( .A(n43371), .Z(n44877) );
  XOR U63671 ( .A(n44878), .B(n44877), .Z(n43373) );
  IV U63672 ( .A(n43370), .Z(n44876) );
  NOR U63673 ( .A(n43371), .B(n44876), .Z(n43372) );
  NOR U63674 ( .A(n43373), .B(n43372), .Z(n43374) );
  NOR U63675 ( .A(n43375), .B(n43374), .Z(n48251) );
  NOR U63676 ( .A(n48249), .B(n48251), .Z(n43376) );
  IV U63677 ( .A(n43376), .Z(n48248) );
  NOR U63678 ( .A(n43377), .B(n48248), .Z(n43378) );
  IV U63679 ( .A(n43378), .Z(n44873) );
  XOR U63680 ( .A(n44872), .B(n44873), .Z(n43386) );
  IV U63681 ( .A(n43386), .Z(n43379) );
  NOR U63682 ( .A(n43385), .B(n43379), .Z(n43380) );
  IV U63683 ( .A(n43380), .Z(n43384) );
  IV U63684 ( .A(n43381), .Z(n43382) );
  NOR U63685 ( .A(n43383), .B(n43382), .Z(n43388) );
  NOR U63686 ( .A(n43384), .B(n43388), .Z(n43391) );
  IV U63687 ( .A(n43385), .Z(n43387) );
  NOR U63688 ( .A(n43387), .B(n43386), .Z(n53435) );
  IV U63689 ( .A(n43388), .Z(n43389) );
  NOR U63690 ( .A(n43389), .B(n44873), .Z(n53421) );
  NOR U63691 ( .A(n53435), .B(n53421), .Z(n43390) );
  IV U63692 ( .A(n43390), .Z(n48256) );
  NOR U63693 ( .A(n43391), .B(n48256), .Z(n44869) );
  XOR U63694 ( .A(n49834), .B(n44869), .Z(n53445) );
  XOR U63695 ( .A(n44870), .B(n53445), .Z(n44864) );
  XOR U63696 ( .A(n44865), .B(n44864), .Z(n48262) );
  IV U63697 ( .A(n43392), .Z(n43393) );
  NOR U63698 ( .A(n43394), .B(n43393), .Z(n44866) );
  IV U63699 ( .A(n43395), .Z(n43396) );
  NOR U63700 ( .A(n43397), .B(n43396), .Z(n48261) );
  NOR U63701 ( .A(n44866), .B(n48261), .Z(n43398) );
  XOR U63702 ( .A(n48262), .B(n43398), .Z(n43405) );
  IV U63703 ( .A(n43405), .Z(n48260) );
  XOR U63704 ( .A(n48258), .B(n48260), .Z(n43399) );
  NOR U63705 ( .A(n43400), .B(n43399), .Z(n54984) );
  IV U63706 ( .A(n43401), .Z(n43402) );
  NOR U63707 ( .A(n43403), .B(n43402), .Z(n44861) );
  NOR U63708 ( .A(n48258), .B(n44861), .Z(n43404) );
  XOR U63709 ( .A(n43405), .B(n43404), .Z(n44859) );
  IV U63710 ( .A(n44859), .Z(n43406) );
  NOR U63711 ( .A(n43407), .B(n43406), .Z(n43408) );
  NOR U63712 ( .A(n54984), .B(n43408), .Z(n48269) );
  IV U63713 ( .A(n43409), .Z(n43410) );
  NOR U63714 ( .A(n43411), .B(n43410), .Z(n44858) );
  NOR U63715 ( .A(n43413), .B(n43412), .Z(n48268) );
  NOR U63716 ( .A(n44858), .B(n48268), .Z(n43414) );
  XOR U63717 ( .A(n48269), .B(n43414), .Z(n48277) );
  XOR U63718 ( .A(n48266), .B(n48277), .Z(n48281) );
  IV U63719 ( .A(n43415), .Z(n43416) );
  NOR U63720 ( .A(n43417), .B(n43416), .Z(n48275) );
  IV U63721 ( .A(n43418), .Z(n43419) );
  NOR U63722 ( .A(n43420), .B(n43419), .Z(n48280) );
  NOR U63723 ( .A(n48275), .B(n48280), .Z(n43421) );
  XOR U63724 ( .A(n48281), .B(n43421), .Z(n49812) );
  XOR U63725 ( .A(n48283), .B(n49812), .Z(n49804) );
  XOR U63726 ( .A(n48285), .B(n49804), .Z(n48292) );
  IV U63727 ( .A(n43422), .Z(n43423) );
  NOR U63728 ( .A(n43424), .B(n43423), .Z(n48293) );
  IV U63729 ( .A(n43425), .Z(n43427) );
  NOR U63730 ( .A(n43427), .B(n43426), .Z(n48289) );
  NOR U63731 ( .A(n48293), .B(n48289), .Z(n43428) );
  XOR U63732 ( .A(n48292), .B(n43428), .Z(n48299) );
  IV U63733 ( .A(n43429), .Z(n43431) );
  NOR U63734 ( .A(n43431), .B(n43430), .Z(n48291) );
  IV U63735 ( .A(n43432), .Z(n43433) );
  NOR U63736 ( .A(n43434), .B(n43433), .Z(n48298) );
  NOR U63737 ( .A(n48291), .B(n48298), .Z(n43435) );
  XOR U63738 ( .A(n48299), .B(n43435), .Z(n44855) );
  XOR U63739 ( .A(n44851), .B(n44855), .Z(n48307) );
  XOR U63740 ( .A(n43436), .B(n48307), .Z(n48303) );
  XOR U63741 ( .A(n43437), .B(n48303), .Z(n48314) );
  IV U63742 ( .A(n43438), .Z(n43440) );
  NOR U63743 ( .A(n43440), .B(n43439), .Z(n48313) );
  IV U63744 ( .A(n43441), .Z(n43443) );
  NOR U63745 ( .A(n43443), .B(n43442), .Z(n44849) );
  NOR U63746 ( .A(n48313), .B(n44849), .Z(n43444) );
  XOR U63747 ( .A(n48314), .B(n43444), .Z(n43445) );
  NOR U63748 ( .A(n43446), .B(n43445), .Z(n43449) );
  IV U63749 ( .A(n43446), .Z(n43448) );
  XOR U63750 ( .A(n48313), .B(n48314), .Z(n43447) );
  NOR U63751 ( .A(n43448), .B(n43447), .Z(n49773) );
  NOR U63752 ( .A(n43449), .B(n49773), .Z(n44844) );
  XOR U63753 ( .A(n43450), .B(n44844), .Z(n49763) );
  IV U63754 ( .A(n43451), .Z(n43452) );
  NOR U63755 ( .A(n43453), .B(n43452), .Z(n49766) );
  IV U63756 ( .A(n43454), .Z(n43456) );
  NOR U63757 ( .A(n43456), .B(n43455), .Z(n49761) );
  NOR U63758 ( .A(n49766), .B(n49761), .Z(n48322) );
  XOR U63759 ( .A(n49763), .B(n48322), .Z(n48320) );
  XOR U63760 ( .A(n48324), .B(n48320), .Z(n43457) );
  NOR U63761 ( .A(n43458), .B(n43457), .Z(n53493) );
  NOR U63762 ( .A(n43460), .B(n43459), .Z(n48319) );
  NOR U63763 ( .A(n43461), .B(n48319), .Z(n43462) );
  XOR U63764 ( .A(n43462), .B(n48320), .Z(n53502) );
  IV U63765 ( .A(n53502), .Z(n43463) );
  NOR U63766 ( .A(n43464), .B(n43463), .Z(n43465) );
  NOR U63767 ( .A(n53493), .B(n43465), .Z(n48329) );
  IV U63768 ( .A(n43466), .Z(n43467) );
  NOR U63769 ( .A(n43468), .B(n43467), .Z(n53500) );
  IV U63770 ( .A(n43469), .Z(n43471) );
  NOR U63771 ( .A(n43471), .B(n43470), .Z(n53506) );
  NOR U63772 ( .A(n53500), .B(n53506), .Z(n48330) );
  XOR U63773 ( .A(n48329), .B(n48330), .Z(n49755) );
  XOR U63774 ( .A(n48331), .B(n49755), .Z(n48337) );
  IV U63775 ( .A(n43472), .Z(n43474) );
  NOR U63776 ( .A(n43474), .B(n43473), .Z(n49750) );
  IV U63777 ( .A(n43475), .Z(n43476) );
  NOR U63778 ( .A(n43477), .B(n43476), .Z(n53516) );
  NOR U63779 ( .A(n49750), .B(n53516), .Z(n48338) );
  XOR U63780 ( .A(n48337), .B(n48338), .Z(n48340) );
  XOR U63781 ( .A(n48339), .B(n48340), .Z(n43478) );
  NOR U63782 ( .A(n43479), .B(n43478), .Z(n53519) );
  IV U63783 ( .A(n43480), .Z(n43481) );
  NOR U63784 ( .A(n43482), .B(n43481), .Z(n48335) );
  NOR U63785 ( .A(n48339), .B(n48335), .Z(n43483) );
  XOR U63786 ( .A(n43483), .B(n48340), .Z(n48347) );
  NOR U63787 ( .A(n43484), .B(n48347), .Z(n43485) );
  NOR U63788 ( .A(n53519), .B(n43485), .Z(n44840) );
  IV U63789 ( .A(n43486), .Z(n43488) );
  NOR U63790 ( .A(n43488), .B(n43487), .Z(n48346) );
  NOR U63791 ( .A(n43490), .B(n43489), .Z(n44839) );
  NOR U63792 ( .A(n48346), .B(n44839), .Z(n43491) );
  XOR U63793 ( .A(n44840), .B(n43491), .Z(n48356) );
  IV U63794 ( .A(n43492), .Z(n43494) );
  NOR U63795 ( .A(n43494), .B(n43493), .Z(n43503) );
  IV U63796 ( .A(n43503), .Z(n48353) );
  IV U63797 ( .A(n43495), .Z(n43496) );
  NOR U63798 ( .A(n43497), .B(n43496), .Z(n48351) );
  IV U63799 ( .A(n48351), .Z(n48350) );
  NOR U63800 ( .A(n48353), .B(n48350), .Z(n43505) );
  IV U63801 ( .A(n43498), .Z(n43500) );
  NOR U63802 ( .A(n43500), .B(n43499), .Z(n48354) );
  NOR U63803 ( .A(n48351), .B(n48354), .Z(n43501) );
  IV U63804 ( .A(n43501), .Z(n43502) );
  NOR U63805 ( .A(n43503), .B(n43502), .Z(n43504) );
  NOR U63806 ( .A(n43505), .B(n43504), .Z(n43506) );
  XOR U63807 ( .A(n48356), .B(n43506), .Z(n48368) );
  IV U63808 ( .A(n43507), .Z(n43508) );
  NOR U63809 ( .A(n43509), .B(n43508), .Z(n48364) );
  IV U63810 ( .A(n43510), .Z(n43511) );
  NOR U63811 ( .A(n43512), .B(n43511), .Z(n48366) );
  NOR U63812 ( .A(n48364), .B(n48366), .Z(n43513) );
  XOR U63813 ( .A(n48368), .B(n43513), .Z(n48361) );
  IV U63814 ( .A(n43514), .Z(n43516) );
  NOR U63815 ( .A(n43516), .B(n43515), .Z(n54944) );
  IV U63816 ( .A(n43517), .Z(n43518) );
  NOR U63817 ( .A(n43519), .B(n43518), .Z(n54938) );
  NOR U63818 ( .A(n54944), .B(n54938), .Z(n48362) );
  XOR U63819 ( .A(n48361), .B(n48362), .Z(n60256) );
  XOR U63820 ( .A(n48372), .B(n60256), .Z(n48374) );
  IV U63821 ( .A(n43520), .Z(n43521) );
  NOR U63822 ( .A(n43522), .B(n43521), .Z(n48373) );
  IV U63823 ( .A(n43523), .Z(n43525) );
  NOR U63824 ( .A(n43525), .B(n43524), .Z(n48380) );
  NOR U63825 ( .A(n48373), .B(n48380), .Z(n43526) );
  XOR U63826 ( .A(n48374), .B(n43526), .Z(n48379) );
  XOR U63827 ( .A(n48377), .B(n48379), .Z(n44835) );
  XOR U63828 ( .A(n43527), .B(n44835), .Z(n48386) );
  XOR U63829 ( .A(n48387), .B(n48386), .Z(n48389) );
  XOR U63830 ( .A(n48388), .B(n48389), .Z(n48397) );
  XOR U63831 ( .A(n43528), .B(n48397), .Z(n48394) );
  XOR U63832 ( .A(n48395), .B(n48394), .Z(n64089) );
  XOR U63833 ( .A(n44830), .B(n64089), .Z(n44831) );
  IV U63834 ( .A(n43530), .Z(n53578) );
  IV U63835 ( .A(n53577), .Z(n43529) );
  NOR U63836 ( .A(n53578), .B(n43529), .Z(n53589) );
  NOR U63837 ( .A(n43530), .B(n53577), .Z(n43531) );
  NOR U63838 ( .A(n43531), .B(n53580), .Z(n43532) );
  NOR U63839 ( .A(n53589), .B(n43532), .Z(n44832) );
  XOR U63840 ( .A(n44831), .B(n44832), .Z(n44828) );
  XOR U63841 ( .A(n43533), .B(n44828), .Z(n44819) );
  IV U63842 ( .A(n43534), .Z(n43535) );
  NOR U63843 ( .A(n43536), .B(n43535), .Z(n44822) );
  IV U63844 ( .A(n43537), .Z(n43539) );
  NOR U63845 ( .A(n43539), .B(n43538), .Z(n44818) );
  NOR U63846 ( .A(n44822), .B(n44818), .Z(n43540) );
  XOR U63847 ( .A(n44819), .B(n43540), .Z(n44817) );
  IV U63848 ( .A(n43541), .Z(n43542) );
  NOR U63849 ( .A(n43543), .B(n43542), .Z(n44815) );
  IV U63850 ( .A(n43544), .Z(n43545) );
  NOR U63851 ( .A(n43546), .B(n43545), .Z(n44813) );
  NOR U63852 ( .A(n44815), .B(n44813), .Z(n43547) );
  XOR U63853 ( .A(n44817), .B(n43547), .Z(n44809) );
  IV U63854 ( .A(n43548), .Z(n43550) );
  NOR U63855 ( .A(n43550), .B(n43549), .Z(n44805) );
  IV U63856 ( .A(n43551), .Z(n43553) );
  NOR U63857 ( .A(n43553), .B(n43552), .Z(n44808) );
  NOR U63858 ( .A(n44805), .B(n44808), .Z(n43554) );
  XOR U63859 ( .A(n44809), .B(n43554), .Z(n44802) );
  IV U63860 ( .A(n43555), .Z(n43556) );
  NOR U63861 ( .A(n43557), .B(n43556), .Z(n44804) );
  IV U63862 ( .A(n43558), .Z(n43559) );
  NOR U63863 ( .A(n43560), .B(n43559), .Z(n44801) );
  NOR U63864 ( .A(n44804), .B(n44801), .Z(n43561) );
  XOR U63865 ( .A(n44802), .B(n43561), .Z(n43562) );
  IV U63866 ( .A(n43562), .Z(n44800) );
  XOR U63867 ( .A(n44796), .B(n44800), .Z(n44794) );
  IV U63868 ( .A(n43563), .Z(n43565) );
  NOR U63869 ( .A(n43565), .B(n43564), .Z(n44798) );
  IV U63870 ( .A(n43566), .Z(n43567) );
  NOR U63871 ( .A(n43568), .B(n43567), .Z(n44793) );
  NOR U63872 ( .A(n44798), .B(n44793), .Z(n43569) );
  XOR U63873 ( .A(n44794), .B(n43569), .Z(n44784) );
  IV U63874 ( .A(n43570), .Z(n43571) );
  NOR U63875 ( .A(n43572), .B(n43571), .Z(n44790) );
  IV U63876 ( .A(n43573), .Z(n43575) );
  NOR U63877 ( .A(n43575), .B(n43574), .Z(n44785) );
  NOR U63878 ( .A(n44790), .B(n44785), .Z(n43576) );
  XOR U63879 ( .A(n44784), .B(n43576), .Z(n49705) );
  IV U63880 ( .A(n49705), .Z(n43582) );
  IV U63881 ( .A(n43577), .Z(n43579) );
  NOR U63882 ( .A(n43579), .B(n43578), .Z(n53637) );
  NOR U63883 ( .A(n43581), .B(n43580), .Z(n49704) );
  NOR U63884 ( .A(n53637), .B(n49704), .Z(n44787) );
  XOR U63885 ( .A(n43582), .B(n44787), .Z(n44782) );
  XOR U63886 ( .A(n44781), .B(n44782), .Z(n43583) );
  NOR U63887 ( .A(n43584), .B(n43583), .Z(n53641) );
  IV U63888 ( .A(n43585), .Z(n43587) );
  NOR U63889 ( .A(n43587), .B(n43586), .Z(n44779) );
  NOR U63890 ( .A(n44781), .B(n44779), .Z(n43588) );
  XOR U63891 ( .A(n43588), .B(n44782), .Z(n43598) );
  NOR U63892 ( .A(n43589), .B(n43598), .Z(n43590) );
  NOR U63893 ( .A(n53641), .B(n43590), .Z(n43596) );
  IV U63894 ( .A(n43596), .Z(n43591) );
  NOR U63895 ( .A(n43592), .B(n43591), .Z(n53648) );
  IV U63896 ( .A(n43593), .Z(n43594) );
  NOR U63897 ( .A(n43595), .B(n43594), .Z(n43597) );
  NOR U63898 ( .A(n43597), .B(n43596), .Z(n43601) );
  IV U63899 ( .A(n43597), .Z(n43600) );
  IV U63900 ( .A(n43598), .Z(n43599) );
  NOR U63901 ( .A(n43600), .B(n43599), .Z(n53644) );
  NOR U63902 ( .A(n43601), .B(n53644), .Z(n44775) );
  NOR U63903 ( .A(n43602), .B(n44775), .Z(n43603) );
  NOR U63904 ( .A(n53648), .B(n43603), .Z(n44771) );
  IV U63905 ( .A(n43604), .Z(n43606) );
  NOR U63906 ( .A(n43606), .B(n43605), .Z(n44774) );
  IV U63907 ( .A(n43607), .Z(n43608) );
  NOR U63908 ( .A(n43609), .B(n43608), .Z(n44770) );
  NOR U63909 ( .A(n44774), .B(n44770), .Z(n43610) );
  XOR U63910 ( .A(n44771), .B(n43610), .Z(n48418) );
  IV U63911 ( .A(n43611), .Z(n43613) );
  NOR U63912 ( .A(n43613), .B(n43612), .Z(n48416) );
  IV U63913 ( .A(n43614), .Z(n43615) );
  NOR U63914 ( .A(n43616), .B(n43615), .Z(n48414) );
  NOR U63915 ( .A(n48416), .B(n48414), .Z(n43617) );
  XOR U63916 ( .A(n48418), .B(n43617), .Z(n43618) );
  IV U63917 ( .A(n43618), .Z(n48422) );
  XOR U63918 ( .A(n48412), .B(n48422), .Z(n44768) );
  IV U63919 ( .A(n43619), .Z(n43621) );
  NOR U63920 ( .A(n43621), .B(n43620), .Z(n48421) );
  NOR U63921 ( .A(n43623), .B(n43622), .Z(n44767) );
  NOR U63922 ( .A(n48421), .B(n44767), .Z(n43624) );
  XOR U63923 ( .A(n44768), .B(n43624), .Z(n43631) );
  IV U63924 ( .A(n43631), .Z(n48428) );
  XOR U63925 ( .A(n48424), .B(n48428), .Z(n43625) );
  NOR U63926 ( .A(n43626), .B(n43625), .Z(n49687) );
  IV U63927 ( .A(n43627), .Z(n43628) );
  NOR U63928 ( .A(n43629), .B(n43628), .Z(n48426) );
  NOR U63929 ( .A(n48424), .B(n48426), .Z(n43630) );
  XOR U63930 ( .A(n43631), .B(n43630), .Z(n44765) );
  IV U63931 ( .A(n44765), .Z(n43632) );
  NOR U63932 ( .A(n43633), .B(n43632), .Z(n43634) );
  NOR U63933 ( .A(n49687), .B(n43634), .Z(n44760) );
  IV U63934 ( .A(n43635), .Z(n43637) );
  NOR U63935 ( .A(n43637), .B(n43636), .Z(n44764) );
  IV U63936 ( .A(n43638), .Z(n43639) );
  NOR U63937 ( .A(n43640), .B(n43639), .Z(n44759) );
  NOR U63938 ( .A(n44764), .B(n44759), .Z(n43641) );
  XOR U63939 ( .A(n44760), .B(n43641), .Z(n44757) );
  XOR U63940 ( .A(n43642), .B(n44757), .Z(n43648) );
  IV U63941 ( .A(n43648), .Z(n43643) );
  NOR U63942 ( .A(n43644), .B(n43643), .Z(n53669) );
  IV U63943 ( .A(n43645), .Z(n43647) );
  NOR U63944 ( .A(n43647), .B(n43646), .Z(n43649) );
  NOR U63945 ( .A(n43649), .B(n43648), .Z(n43652) );
  IV U63946 ( .A(n43649), .Z(n43651) );
  XOR U63947 ( .A(n49686), .B(n44757), .Z(n43650) );
  NOR U63948 ( .A(n43651), .B(n43650), .Z(n49680) );
  NOR U63949 ( .A(n43652), .B(n49680), .Z(n44751) );
  NOR U63950 ( .A(n43653), .B(n44751), .Z(n43654) );
  NOR U63951 ( .A(n53669), .B(n43654), .Z(n48438) );
  IV U63952 ( .A(n43655), .Z(n43656) );
  NOR U63953 ( .A(n43657), .B(n43656), .Z(n44750) );
  IV U63954 ( .A(n43658), .Z(n43659) );
  NOR U63955 ( .A(n43660), .B(n43659), .Z(n48437) );
  NOR U63956 ( .A(n44750), .B(n48437), .Z(n43661) );
  XOR U63957 ( .A(n48438), .B(n43661), .Z(n54834) );
  NOR U63958 ( .A(n43663), .B(n43662), .Z(n54839) );
  IV U63959 ( .A(n43664), .Z(n43666) );
  NOR U63960 ( .A(n43666), .B(n43665), .Z(n54831) );
  NOR U63961 ( .A(n54839), .B(n54831), .Z(n48441) );
  XOR U63962 ( .A(n54834), .B(n48441), .Z(n48443) );
  IV U63963 ( .A(n43667), .Z(n43669) );
  NOR U63964 ( .A(n43669), .B(n43668), .Z(n48442) );
  IV U63965 ( .A(n43670), .Z(n43672) );
  NOR U63966 ( .A(n43672), .B(n43671), .Z(n48447) );
  NOR U63967 ( .A(n48442), .B(n48447), .Z(n43673) );
  XOR U63968 ( .A(n48443), .B(n43673), .Z(n54825) );
  XOR U63969 ( .A(n48450), .B(n54825), .Z(n48452) );
  IV U63970 ( .A(n43674), .Z(n43676) );
  NOR U63971 ( .A(n43676), .B(n43675), .Z(n53679) );
  IV U63972 ( .A(n43677), .Z(n43678) );
  NOR U63973 ( .A(n43679), .B(n43678), .Z(n53684) );
  NOR U63974 ( .A(n53679), .B(n53684), .Z(n48453) );
  XOR U63975 ( .A(n48452), .B(n48453), .Z(n48459) );
  XOR U63976 ( .A(n43680), .B(n48459), .Z(n48465) );
  IV U63977 ( .A(n43681), .Z(n43683) );
  NOR U63978 ( .A(n43683), .B(n43682), .Z(n48461) );
  IV U63979 ( .A(n43684), .Z(n43686) );
  NOR U63980 ( .A(n43686), .B(n43685), .Z(n48464) );
  NOR U63981 ( .A(n48461), .B(n48464), .Z(n43687) );
  XOR U63982 ( .A(n48465), .B(n43687), .Z(n44748) );
  NOR U63983 ( .A(n43689), .B(n43688), .Z(n53694) );
  IV U63984 ( .A(n43690), .Z(n43692) );
  NOR U63985 ( .A(n43692), .B(n43691), .Z(n49664) );
  NOR U63986 ( .A(n53694), .B(n49664), .Z(n44749) );
  XOR U63987 ( .A(n44748), .B(n44749), .Z(n49660) );
  IV U63988 ( .A(n43693), .Z(n43695) );
  NOR U63989 ( .A(n43695), .B(n43694), .Z(n49668) );
  IV U63990 ( .A(n43696), .Z(n43697) );
  NOR U63991 ( .A(n43698), .B(n43697), .Z(n49659) );
  NOR U63992 ( .A(n49668), .B(n49659), .Z(n44744) );
  XOR U63993 ( .A(n49660), .B(n44744), .Z(n44745) );
  XOR U63994 ( .A(n53716), .B(n44745), .Z(n44741) );
  XOR U63995 ( .A(n44738), .B(n44741), .Z(n44736) );
  IV U63996 ( .A(n43699), .Z(n43701) );
  NOR U63997 ( .A(n43701), .B(n43700), .Z(n44740) );
  IV U63998 ( .A(n43702), .Z(n43703) );
  NOR U63999 ( .A(n43704), .B(n43703), .Z(n44735) );
  NOR U64000 ( .A(n44740), .B(n44735), .Z(n43705) );
  XOR U64001 ( .A(n44736), .B(n43705), .Z(n44732) );
  XOR U64002 ( .A(n44733), .B(n44732), .Z(n44729) );
  XOR U64003 ( .A(n44727), .B(n44729), .Z(n53737) );
  IV U64004 ( .A(n53737), .Z(n43713) );
  IV U64005 ( .A(n43706), .Z(n43707) );
  NOR U64006 ( .A(n43708), .B(n43707), .Z(n53739) );
  IV U64007 ( .A(n43709), .Z(n43711) );
  NOR U64008 ( .A(n43711), .B(n43710), .Z(n44725) );
  NOR U64009 ( .A(n53739), .B(n44725), .Z(n43712) );
  XOR U64010 ( .A(n43713), .B(n43712), .Z(n44724) );
  XOR U64011 ( .A(n44722), .B(n44724), .Z(n44717) );
  IV U64012 ( .A(n43714), .Z(n43716) );
  NOR U64013 ( .A(n43716), .B(n43715), .Z(n44719) );
  IV U64014 ( .A(n43717), .Z(n43718) );
  NOR U64015 ( .A(n43719), .B(n43718), .Z(n44716) );
  NOR U64016 ( .A(n44719), .B(n44716), .Z(n43720) );
  XOR U64017 ( .A(n44717), .B(n43720), .Z(n44713) );
  XOR U64018 ( .A(n43721), .B(n44713), .Z(n54794) );
  XOR U64019 ( .A(n48478), .B(n54794), .Z(n48479) );
  IV U64020 ( .A(n43722), .Z(n43723) );
  NOR U64021 ( .A(n43724), .B(n43723), .Z(n49636) );
  IV U64022 ( .A(n43725), .Z(n43727) );
  NOR U64023 ( .A(n43727), .B(n43726), .Z(n49632) );
  NOR U64024 ( .A(n49636), .B(n49632), .Z(n48480) );
  XOR U64025 ( .A(n48479), .B(n48480), .Z(n44710) );
  XOR U64026 ( .A(n43728), .B(n44710), .Z(n44704) );
  XOR U64027 ( .A(n49625), .B(n44704), .Z(n48497) );
  XOR U64028 ( .A(n48485), .B(n48497), .Z(n48501) );
  XOR U64029 ( .A(n43729), .B(n48501), .Z(n48510) );
  XOR U64030 ( .A(n48511), .B(n48510), .Z(n48513) );
  XOR U64031 ( .A(n43730), .B(n48513), .Z(n48521) );
  IV U64032 ( .A(n43731), .Z(n43733) );
  NOR U64033 ( .A(n43733), .B(n43732), .Z(n48525) );
  IV U64034 ( .A(n43734), .Z(n43735) );
  NOR U64035 ( .A(n43736), .B(n43735), .Z(n48520) );
  NOR U64036 ( .A(n48525), .B(n48520), .Z(n43737) );
  XOR U64037 ( .A(n48521), .B(n43737), .Z(n53758) );
  IV U64038 ( .A(n53758), .Z(n43744) );
  IV U64039 ( .A(n43738), .Z(n43739) );
  NOR U64040 ( .A(n43740), .B(n43739), .Z(n53761) );
  IV U64041 ( .A(n43741), .Z(n43742) );
  NOR U64042 ( .A(n43743), .B(n43742), .Z(n53756) );
  NOR U64043 ( .A(n53761), .B(n53756), .Z(n44697) );
  XOR U64044 ( .A(n43744), .B(n44697), .Z(n44699) );
  IV U64045 ( .A(n43745), .Z(n43747) );
  NOR U64046 ( .A(n43747), .B(n43746), .Z(n44698) );
  IV U64047 ( .A(n43748), .Z(n43750) );
  NOR U64048 ( .A(n43750), .B(n43749), .Z(n44695) );
  NOR U64049 ( .A(n44698), .B(n44695), .Z(n43751) );
  XOR U64050 ( .A(n44699), .B(n43751), .Z(n43759) );
  IV U64051 ( .A(n43759), .Z(n43752) );
  NOR U64052 ( .A(n43753), .B(n43752), .Z(n53777) );
  IV U64053 ( .A(n43754), .Z(n43755) );
  NOR U64054 ( .A(n43756), .B(n43755), .Z(n43760) );
  IV U64055 ( .A(n43760), .Z(n43758) );
  XOR U64056 ( .A(n44698), .B(n44699), .Z(n43757) );
  NOR U64057 ( .A(n43758), .B(n43757), .Z(n53769) );
  NOR U64058 ( .A(n43760), .B(n43759), .Z(n43761) );
  NOR U64059 ( .A(n53769), .B(n43761), .Z(n44692) );
  NOR U64060 ( .A(n43762), .B(n44692), .Z(n43763) );
  NOR U64061 ( .A(n53777), .B(n43763), .Z(n44688) );
  XOR U64062 ( .A(n43764), .B(n44688), .Z(n48541) );
  XOR U64063 ( .A(n43765), .B(n48541), .Z(n48547) );
  XOR U64064 ( .A(n43766), .B(n48547), .Z(n48542) );
  IV U64065 ( .A(n43767), .Z(n43768) );
  NOR U64066 ( .A(n43769), .B(n43768), .Z(n49604) );
  IV U64067 ( .A(n43770), .Z(n43771) );
  NOR U64068 ( .A(n43772), .B(n43771), .Z(n53798) );
  NOR U64069 ( .A(n49604), .B(n53798), .Z(n48543) );
  XOR U64070 ( .A(n48542), .B(n48543), .Z(n48562) );
  XOR U64071 ( .A(n48561), .B(n48562), .Z(n48555) );
  XOR U64072 ( .A(n43773), .B(n48555), .Z(n44678) );
  XOR U64073 ( .A(n44679), .B(n44678), .Z(n44681) );
  XOR U64074 ( .A(n44680), .B(n44681), .Z(n48568) );
  XOR U64075 ( .A(n43774), .B(n48568), .Z(n43775) );
  IV U64076 ( .A(n43775), .Z(n53821) );
  XOR U64077 ( .A(n48570), .B(n53821), .Z(n48571) );
  XOR U64078 ( .A(n48572), .B(n48571), .Z(n49580) );
  XOR U64079 ( .A(n44675), .B(n49580), .Z(n48579) );
  XOR U64080 ( .A(n48580), .B(n48579), .Z(n48588) );
  XOR U64081 ( .A(n48587), .B(n48588), .Z(n48593) );
  NOR U64082 ( .A(n43777), .B(n43776), .Z(n48575) );
  NOR U64083 ( .A(n43779), .B(n43778), .Z(n43781) );
  IV U64084 ( .A(n43780), .Z(n48590) );
  NOR U64085 ( .A(n43781), .B(n48590), .Z(n43782) );
  NOR U64086 ( .A(n48575), .B(n43782), .Z(n43783) );
  XOR U64087 ( .A(n48593), .B(n43783), .Z(n44670) );
  IV U64088 ( .A(n43784), .Z(n43786) );
  NOR U64089 ( .A(n43786), .B(n43785), .Z(n54713) );
  IV U64090 ( .A(n43787), .Z(n43789) );
  NOR U64091 ( .A(n43789), .B(n43788), .Z(n44671) );
  NOR U64092 ( .A(n54713), .B(n44671), .Z(n43790) );
  XOR U64093 ( .A(n44670), .B(n43790), .Z(n48602) );
  XOR U64094 ( .A(n48596), .B(n48602), .Z(n44666) );
  IV U64095 ( .A(n48600), .Z(n43791) );
  NOR U64096 ( .A(n43791), .B(n48598), .Z(n43793) );
  NOR U64097 ( .A(n44665), .B(n44667), .Z(n43792) );
  NOR U64098 ( .A(n43793), .B(n43792), .Z(n43794) );
  XOR U64099 ( .A(n44666), .B(n43794), .Z(n44663) );
  XOR U64100 ( .A(n44662), .B(n44663), .Z(n44657) );
  IV U64101 ( .A(n43795), .Z(n43796) );
  NOR U64102 ( .A(n43797), .B(n43796), .Z(n44660) );
  IV U64103 ( .A(n43798), .Z(n43799) );
  NOR U64104 ( .A(n43800), .B(n43799), .Z(n44656) );
  NOR U64105 ( .A(n44660), .B(n44656), .Z(n43801) );
  XOR U64106 ( .A(n44657), .B(n43801), .Z(n48609) );
  IV U64107 ( .A(n43802), .Z(n43804) );
  NOR U64108 ( .A(n43804), .B(n43803), .Z(n48608) );
  IV U64109 ( .A(n43805), .Z(n43807) );
  NOR U64110 ( .A(n43807), .B(n43806), .Z(n48612) );
  NOR U64111 ( .A(n48608), .B(n48612), .Z(n48615) );
  XOR U64112 ( .A(n48609), .B(n48615), .Z(n44654) );
  IV U64113 ( .A(n43808), .Z(n43809) );
  NOR U64114 ( .A(n43810), .B(n43809), .Z(n44653) );
  IV U64115 ( .A(n43811), .Z(n43813) );
  NOR U64116 ( .A(n43813), .B(n43812), .Z(n44651) );
  NOR U64117 ( .A(n44653), .B(n44651), .Z(n43814) );
  XOR U64118 ( .A(n44654), .B(n43814), .Z(n48625) );
  XOR U64119 ( .A(n48626), .B(n48625), .Z(n48628) );
  IV U64120 ( .A(n43815), .Z(n43817) );
  NOR U64121 ( .A(n43817), .B(n43816), .Z(n48627) );
  IV U64122 ( .A(n43818), .Z(n43820) );
  NOR U64123 ( .A(n43820), .B(n43819), .Z(n44649) );
  NOR U64124 ( .A(n48627), .B(n44649), .Z(n43821) );
  XOR U64125 ( .A(n48628), .B(n43821), .Z(n48635) );
  XOR U64126 ( .A(n43822), .B(n48635), .Z(n48641) );
  XOR U64127 ( .A(n48639), .B(n48641), .Z(n48652) );
  IV U64128 ( .A(n48652), .Z(n43830) );
  IV U64129 ( .A(n43823), .Z(n43824) );
  NOR U64130 ( .A(n43825), .B(n43824), .Z(n44647) );
  IV U64131 ( .A(n43826), .Z(n43828) );
  NOR U64132 ( .A(n43828), .B(n43827), .Z(n48651) );
  NOR U64133 ( .A(n44647), .B(n48651), .Z(n43829) );
  XOR U64134 ( .A(n43830), .B(n43829), .Z(n48657) );
  IV U64135 ( .A(n43831), .Z(n43832) );
  NOR U64136 ( .A(n43833), .B(n43832), .Z(n48649) );
  IV U64137 ( .A(n43834), .Z(n43835) );
  NOR U64138 ( .A(n43836), .B(n43835), .Z(n48655) );
  NOR U64139 ( .A(n48649), .B(n48655), .Z(n43837) );
  XOR U64140 ( .A(n48657), .B(n43837), .Z(n48659) );
  NOR U64141 ( .A(n43838), .B(n48659), .Z(n43841) );
  IV U64142 ( .A(n43838), .Z(n43840) );
  XOR U64143 ( .A(n48649), .B(n48657), .Z(n43839) );
  NOR U64144 ( .A(n43840), .B(n43839), .Z(n54655) );
  NOR U64145 ( .A(n43841), .B(n54655), .Z(n48667) );
  IV U64146 ( .A(n43842), .Z(n43843) );
  NOR U64147 ( .A(n43844), .B(n43843), .Z(n48658) );
  IV U64148 ( .A(n43845), .Z(n43847) );
  NOR U64149 ( .A(n43847), .B(n43846), .Z(n48666) );
  NOR U64150 ( .A(n48658), .B(n48666), .Z(n43848) );
  XOR U64151 ( .A(n48667), .B(n43848), .Z(n48673) );
  IV U64152 ( .A(n43849), .Z(n43850) );
  NOR U64153 ( .A(n43851), .B(n43850), .Z(n48664) );
  IV U64154 ( .A(n43852), .Z(n43853) );
  NOR U64155 ( .A(n43854), .B(n43853), .Z(n48671) );
  NOR U64156 ( .A(n48664), .B(n48671), .Z(n43855) );
  XOR U64157 ( .A(n48673), .B(n43855), .Z(n43856) );
  IV U64158 ( .A(n43856), .Z(n44643) );
  XOR U64159 ( .A(n44642), .B(n44643), .Z(n49533) );
  XOR U64160 ( .A(n44645), .B(n49533), .Z(n48676) );
  XOR U64161 ( .A(n43857), .B(n48676), .Z(n53888) );
  XOR U64162 ( .A(n44637), .B(n53888), .Z(n44624) );
  XOR U64163 ( .A(n43858), .B(n44624), .Z(n44635) );
  IV U64164 ( .A(n44630), .Z(n43859) );
  NOR U64165 ( .A(n44631), .B(n43859), .Z(n44626) );
  NOR U64166 ( .A(n43860), .B(n44630), .Z(n43861) );
  NOR U64167 ( .A(n43861), .B(n44633), .Z(n43862) );
  NOR U64168 ( .A(n44626), .B(n43862), .Z(n43863) );
  XOR U64169 ( .A(n44635), .B(n43863), .Z(n48686) );
  IV U64170 ( .A(n43864), .Z(n43866) );
  NOR U64171 ( .A(n43866), .B(n43865), .Z(n48689) );
  IV U64172 ( .A(n43867), .Z(n43868) );
  NOR U64173 ( .A(n43869), .B(n43868), .Z(n48687) );
  NOR U64174 ( .A(n48689), .B(n48687), .Z(n43870) );
  XOR U64175 ( .A(n48686), .B(n43870), .Z(n48703) );
  IV U64176 ( .A(n43871), .Z(n43872) );
  NOR U64177 ( .A(n43873), .B(n43872), .Z(n44621) );
  IV U64178 ( .A(n43874), .Z(n43875) );
  NOR U64179 ( .A(n43876), .B(n43875), .Z(n48702) );
  NOR U64180 ( .A(n44621), .B(n48702), .Z(n43877) );
  XOR U64181 ( .A(n48703), .B(n43877), .Z(n44617) );
  IV U64182 ( .A(n43878), .Z(n43880) );
  NOR U64183 ( .A(n43880), .B(n43879), .Z(n53910) );
  IV U64184 ( .A(n43881), .Z(n43883) );
  NOR U64185 ( .A(n43883), .B(n43882), .Z(n44618) );
  NOR U64186 ( .A(n53910), .B(n44618), .Z(n43884) );
  XOR U64187 ( .A(n44617), .B(n43884), .Z(n44615) );
  IV U64188 ( .A(n43885), .Z(n43887) );
  NOR U64189 ( .A(n43887), .B(n43886), .Z(n53908) );
  IV U64190 ( .A(n43888), .Z(n43889) );
  NOR U64191 ( .A(n43890), .B(n43889), .Z(n43891) );
  NOR U64192 ( .A(n53908), .B(n43891), .Z(n44616) );
  XOR U64193 ( .A(n44615), .B(n44616), .Z(n48712) );
  XOR U64194 ( .A(n48716), .B(n48712), .Z(n48723) );
  IV U64195 ( .A(n43892), .Z(n43894) );
  NOR U64196 ( .A(n43894), .B(n43893), .Z(n44613) );
  IV U64197 ( .A(n43895), .Z(n43897) );
  NOR U64198 ( .A(n43897), .B(n43896), .Z(n48722) );
  NOR U64199 ( .A(n44613), .B(n48722), .Z(n43898) );
  XOR U64200 ( .A(n48723), .B(n43898), .Z(n48730) );
  XOR U64201 ( .A(n43899), .B(n48730), .Z(n48743) );
  XOR U64202 ( .A(n43900), .B(n48743), .Z(n43901) );
  IV U64203 ( .A(n43901), .Z(n48748) );
  NOR U64204 ( .A(n43902), .B(n48748), .Z(n49489) );
  NOR U64205 ( .A(n43904), .B(n43903), .Z(n43913) );
  IV U64206 ( .A(n43913), .Z(n43910) );
  IV U64207 ( .A(n43905), .Z(n43906) );
  NOR U64208 ( .A(n43907), .B(n43906), .Z(n43908) );
  IV U64209 ( .A(n43908), .Z(n48749) );
  XOR U64210 ( .A(n48749), .B(n48748), .Z(n43916) );
  IV U64211 ( .A(n43916), .Z(n43909) );
  NOR U64212 ( .A(n43910), .B(n43909), .Z(n49487) );
  NOR U64213 ( .A(n49489), .B(n49487), .Z(n43911) );
  IV U64214 ( .A(n43911), .Z(n48750) );
  NOR U64215 ( .A(n43913), .B(n43912), .Z(n43914) );
  IV U64216 ( .A(n43914), .Z(n43915) );
  NOR U64217 ( .A(n43916), .B(n43915), .Z(n43917) );
  NOR U64218 ( .A(n48750), .B(n43917), .Z(n44606) );
  XOR U64219 ( .A(n44607), .B(n44606), .Z(n44609) );
  XOR U64220 ( .A(n44608), .B(n44609), .Z(n48756) );
  IV U64221 ( .A(n48756), .Z(n43925) );
  IV U64222 ( .A(n43918), .Z(n43920) );
  NOR U64223 ( .A(n43920), .B(n43919), .Z(n44604) );
  IV U64224 ( .A(n43921), .Z(n43922) );
  NOR U64225 ( .A(n43923), .B(n43922), .Z(n48755) );
  NOR U64226 ( .A(n44604), .B(n48755), .Z(n43924) );
  XOR U64227 ( .A(n43925), .B(n43924), .Z(n48762) );
  IV U64228 ( .A(n43926), .Z(n43927) );
  NOR U64229 ( .A(n43928), .B(n43927), .Z(n48753) );
  IV U64230 ( .A(n43929), .Z(n43931) );
  NOR U64231 ( .A(n43931), .B(n43930), .Z(n48760) );
  NOR U64232 ( .A(n48753), .B(n48760), .Z(n43932) );
  XOR U64233 ( .A(n48762), .B(n43932), .Z(n44598) );
  IV U64234 ( .A(n43933), .Z(n43935) );
  NOR U64235 ( .A(n43935), .B(n43934), .Z(n44597) );
  IV U64236 ( .A(n43936), .Z(n43938) );
  NOR U64237 ( .A(n43938), .B(n43937), .Z(n44600) );
  NOR U64238 ( .A(n44597), .B(n44600), .Z(n43939) );
  XOR U64239 ( .A(n44598), .B(n43939), .Z(n48768) );
  XOR U64240 ( .A(n43940), .B(n48768), .Z(n49458) );
  XOR U64241 ( .A(n44594), .B(n49458), .Z(n49451) );
  XOR U64242 ( .A(n48775), .B(n49451), .Z(n48772) );
  IV U64243 ( .A(n43941), .Z(n43942) );
  NOR U64244 ( .A(n43943), .B(n43942), .Z(n48776) );
  IV U64245 ( .A(n43944), .Z(n43946) );
  NOR U64246 ( .A(n43946), .B(n43945), .Z(n48771) );
  NOR U64247 ( .A(n48776), .B(n48771), .Z(n43947) );
  XOR U64248 ( .A(n48772), .B(n43947), .Z(n48794) );
  IV U64249 ( .A(n43950), .Z(n43948) );
  NOR U64250 ( .A(n43949), .B(n43948), .Z(n43953) );
  IV U64251 ( .A(n43949), .Z(n43951) );
  NOR U64252 ( .A(n43951), .B(n43950), .Z(n48782) );
  NOR U64253 ( .A(n48789), .B(n48782), .Z(n43952) );
  NOR U64254 ( .A(n43953), .B(n43952), .Z(n43954) );
  XOR U64255 ( .A(n48794), .B(n43954), .Z(n49440) );
  IV U64256 ( .A(n43955), .Z(n43957) );
  NOR U64257 ( .A(n43957), .B(n43956), .Z(n49443) );
  IV U64258 ( .A(n43958), .Z(n43960) );
  NOR U64259 ( .A(n43960), .B(n43959), .Z(n49438) );
  NOR U64260 ( .A(n49443), .B(n49438), .Z(n48796) );
  XOR U64261 ( .A(n49440), .B(n48796), .Z(n48797) );
  XOR U64262 ( .A(n48798), .B(n48797), .Z(n44592) );
  IV U64263 ( .A(n43961), .Z(n43962) );
  NOR U64264 ( .A(n43963), .B(n43962), .Z(n48801) );
  IV U64265 ( .A(n43964), .Z(n43966) );
  NOR U64266 ( .A(n43966), .B(n43965), .Z(n44591) );
  NOR U64267 ( .A(n48801), .B(n44591), .Z(n43967) );
  XOR U64268 ( .A(n44592), .B(n43967), .Z(n44586) );
  IV U64269 ( .A(n43968), .Z(n43970) );
  NOR U64270 ( .A(n43970), .B(n43969), .Z(n49427) );
  IV U64271 ( .A(n43971), .Z(n43972) );
  NOR U64272 ( .A(n43973), .B(n43972), .Z(n49422) );
  NOR U64273 ( .A(n49427), .B(n49422), .Z(n44587) );
  XOR U64274 ( .A(n44586), .B(n44587), .Z(n48806) );
  IV U64275 ( .A(n43974), .Z(n43975) );
  NOR U64276 ( .A(n43976), .B(n43975), .Z(n44588) );
  IV U64277 ( .A(n43977), .Z(n43979) );
  NOR U64278 ( .A(n43979), .B(n43978), .Z(n48805) );
  NOR U64279 ( .A(n44588), .B(n48805), .Z(n43980) );
  XOR U64280 ( .A(n48806), .B(n43980), .Z(n44575) );
  IV U64281 ( .A(n43981), .Z(n43982) );
  NOR U64282 ( .A(n43983), .B(n43982), .Z(n44576) );
  IV U64283 ( .A(n43984), .Z(n43985) );
  NOR U64284 ( .A(n43986), .B(n43985), .Z(n44581) );
  NOR U64285 ( .A(n44576), .B(n44581), .Z(n43987) );
  XOR U64286 ( .A(n44575), .B(n43987), .Z(n44579) );
  IV U64287 ( .A(n43988), .Z(n43990) );
  NOR U64288 ( .A(n43990), .B(n43989), .Z(n44578) );
  IV U64289 ( .A(n43991), .Z(n43993) );
  NOR U64290 ( .A(n43993), .B(n43992), .Z(n44573) );
  NOR U64291 ( .A(n44578), .B(n44573), .Z(n43994) );
  XOR U64292 ( .A(n44579), .B(n43994), .Z(n44002) );
  IV U64293 ( .A(n44002), .Z(n43995) );
  NOR U64294 ( .A(n43996), .B(n43995), .Z(n49411) );
  IV U64295 ( .A(n43997), .Z(n43999) );
  NOR U64296 ( .A(n43999), .B(n43998), .Z(n44003) );
  IV U64297 ( .A(n44003), .Z(n44001) );
  XOR U64298 ( .A(n44578), .B(n44579), .Z(n44000) );
  NOR U64299 ( .A(n44001), .B(n44000), .Z(n53956) );
  NOR U64300 ( .A(n44003), .B(n44002), .Z(n44004) );
  NOR U64301 ( .A(n53956), .B(n44004), .Z(n44568) );
  NOR U64302 ( .A(n44005), .B(n44568), .Z(n44006) );
  NOR U64303 ( .A(n49411), .B(n44006), .Z(n44007) );
  IV U64304 ( .A(n44007), .Z(n44565) );
  IV U64305 ( .A(n44008), .Z(n44010) );
  NOR U64306 ( .A(n44010), .B(n44009), .Z(n44567) );
  IV U64307 ( .A(n44011), .Z(n44013) );
  NOR U64308 ( .A(n44013), .B(n44012), .Z(n44564) );
  NOR U64309 ( .A(n44567), .B(n44564), .Z(n44014) );
  XOR U64310 ( .A(n44565), .B(n44014), .Z(n53972) );
  IV U64311 ( .A(n44015), .Z(n44016) );
  NOR U64312 ( .A(n44017), .B(n44016), .Z(n53965) );
  IV U64313 ( .A(n44018), .Z(n44019) );
  NOR U64314 ( .A(n44020), .B(n44019), .Z(n49407) );
  NOR U64315 ( .A(n53965), .B(n49407), .Z(n53970) );
  XOR U64316 ( .A(n53972), .B(n53970), .Z(n44561) );
  IV U64317 ( .A(n44021), .Z(n44022) );
  NOR U64318 ( .A(n44023), .B(n44022), .Z(n53980) );
  IV U64319 ( .A(n44024), .Z(n44026) );
  NOR U64320 ( .A(n44026), .B(n44025), .Z(n53969) );
  NOR U64321 ( .A(n53980), .B(n53969), .Z(n44562) );
  XOR U64322 ( .A(n44561), .B(n44562), .Z(n48818) );
  XOR U64323 ( .A(n48819), .B(n48818), .Z(n48821) );
  XOR U64324 ( .A(n48820), .B(n48821), .Z(n48832) );
  NOR U64325 ( .A(n44028), .B(n44027), .Z(n44030) );
  NOR U64326 ( .A(n48827), .B(n48828), .Z(n44029) );
  NOR U64327 ( .A(n44030), .B(n44029), .Z(n44031) );
  XOR U64328 ( .A(n48832), .B(n44031), .Z(n44558) );
  IV U64329 ( .A(n44558), .Z(n54007) );
  IV U64330 ( .A(n44032), .Z(n44033) );
  NOR U64331 ( .A(n44034), .B(n44033), .Z(n54011) );
  IV U64332 ( .A(n44035), .Z(n44036) );
  NOR U64333 ( .A(n44037), .B(n44036), .Z(n54008) );
  NOR U64334 ( .A(n54011), .B(n54008), .Z(n44038) );
  XOR U64335 ( .A(n54007), .B(n44038), .Z(n44553) );
  XOR U64336 ( .A(n44039), .B(n44553), .Z(n48842) );
  IV U64337 ( .A(n44042), .Z(n44040) );
  NOR U64338 ( .A(n44041), .B(n44040), .Z(n44045) );
  IV U64339 ( .A(n44041), .Z(n44043) );
  NOR U64340 ( .A(n44043), .B(n44042), .Z(n44554) );
  NOR U64341 ( .A(n48838), .B(n44554), .Z(n44044) );
  NOR U64342 ( .A(n44045), .B(n44044), .Z(n44046) );
  XOR U64343 ( .A(n48842), .B(n44046), .Z(n48852) );
  IV U64344 ( .A(n44047), .Z(n44048) );
  NOR U64345 ( .A(n44049), .B(n44048), .Z(n48834) );
  IV U64346 ( .A(n44050), .Z(n44052) );
  NOR U64347 ( .A(n44052), .B(n44051), .Z(n48851) );
  NOR U64348 ( .A(n48834), .B(n48851), .Z(n44053) );
  XOR U64349 ( .A(n48852), .B(n44053), .Z(n44054) );
  IV U64350 ( .A(n44054), .Z(n48858) );
  XOR U64351 ( .A(n48854), .B(n48858), .Z(n44055) );
  NOR U64352 ( .A(n44056), .B(n44055), .Z(n54028) );
  IV U64353 ( .A(n44057), .Z(n44058) );
  NOR U64354 ( .A(n44059), .B(n44058), .Z(n48856) );
  NOR U64355 ( .A(n48854), .B(n48856), .Z(n44060) );
  XOR U64356 ( .A(n48858), .B(n44060), .Z(n44550) );
  NOR U64357 ( .A(n44061), .B(n44550), .Z(n44062) );
  NOR U64358 ( .A(n54028), .B(n44062), .Z(n44546) );
  XOR U64359 ( .A(n44063), .B(n44546), .Z(n54527) );
  XOR U64360 ( .A(n54529), .B(n54527), .Z(n48863) );
  XOR U64361 ( .A(n44064), .B(n48863), .Z(n48875) );
  IV U64362 ( .A(n48875), .Z(n44072) );
  IV U64363 ( .A(n44065), .Z(n44067) );
  NOR U64364 ( .A(n44067), .B(n44066), .Z(n48870) );
  IV U64365 ( .A(n44068), .Z(n44070) );
  NOR U64366 ( .A(n44070), .B(n44069), .Z(n48873) );
  NOR U64367 ( .A(n48870), .B(n48873), .Z(n44071) );
  XOR U64368 ( .A(n44072), .B(n44071), .Z(n44543) );
  XOR U64369 ( .A(n44542), .B(n44543), .Z(n44537) );
  XOR U64370 ( .A(n44073), .B(n44537), .Z(n48879) );
  XOR U64371 ( .A(n48880), .B(n48879), .Z(n48885) );
  XOR U64372 ( .A(n48881), .B(n48885), .Z(n44534) );
  XOR U64373 ( .A(n44074), .B(n44534), .Z(n44526) );
  XOR U64374 ( .A(n44527), .B(n44526), .Z(n44529) );
  NOR U64375 ( .A(n44081), .B(n44529), .Z(n49361) );
  IV U64376 ( .A(n44075), .Z(n44076) );
  NOR U64377 ( .A(n44077), .B(n44076), .Z(n49352) );
  IV U64378 ( .A(n44078), .Z(n44080) );
  NOR U64379 ( .A(n44080), .B(n44079), .Z(n44528) );
  XOR U64380 ( .A(n44528), .B(n44529), .Z(n49353) );
  IV U64381 ( .A(n49353), .Z(n44519) );
  XOR U64382 ( .A(n49352), .B(n44519), .Z(n44083) );
  NOR U64383 ( .A(n44519), .B(n44081), .Z(n44082) );
  NOR U64384 ( .A(n44083), .B(n44082), .Z(n44084) );
  NOR U64385 ( .A(n49361), .B(n44084), .Z(n44085) );
  IV U64386 ( .A(n44085), .Z(n49349) );
  IV U64387 ( .A(n44086), .Z(n44087) );
  NOR U64388 ( .A(n44088), .B(n44087), .Z(n49358) );
  IV U64389 ( .A(n44089), .Z(n44090) );
  NOR U64390 ( .A(n44091), .B(n44090), .Z(n49348) );
  NOR U64391 ( .A(n49358), .B(n49348), .Z(n44092) );
  IV U64392 ( .A(n44092), .Z(n44523) );
  XOR U64393 ( .A(n49349), .B(n44523), .Z(n48891) );
  IV U64394 ( .A(n44093), .Z(n44095) );
  NOR U64395 ( .A(n44095), .B(n44094), .Z(n44517) );
  IV U64396 ( .A(n44096), .Z(n44098) );
  NOR U64397 ( .A(n44098), .B(n44097), .Z(n48889) );
  NOR U64398 ( .A(n44517), .B(n48889), .Z(n44099) );
  XOR U64399 ( .A(n48891), .B(n44099), .Z(n44100) );
  IV U64400 ( .A(n44100), .Z(n48893) );
  XOR U64401 ( .A(n48892), .B(n48893), .Z(n44107) );
  IV U64402 ( .A(n44107), .Z(n44101) );
  NOR U64403 ( .A(n44106), .B(n44101), .Z(n44102) );
  IV U64404 ( .A(n44102), .Z(n44103) );
  NOR U64405 ( .A(n44104), .B(n44103), .Z(n49333) );
  IV U64406 ( .A(n44104), .Z(n44105) );
  NOR U64407 ( .A(n44105), .B(n48893), .Z(n49337) );
  IV U64408 ( .A(n44106), .Z(n44108) );
  NOR U64409 ( .A(n44108), .B(n44107), .Z(n54059) );
  NOR U64410 ( .A(n49337), .B(n54059), .Z(n44109) );
  IV U64411 ( .A(n44109), .Z(n49330) );
  NOR U64412 ( .A(n49333), .B(n49330), .Z(n48896) );
  IV U64413 ( .A(n44110), .Z(n44111) );
  NOR U64414 ( .A(n44112), .B(n44111), .Z(n54062) );
  IV U64415 ( .A(n44113), .Z(n44114) );
  NOR U64416 ( .A(n44115), .B(n44114), .Z(n49329) );
  NOR U64417 ( .A(n54062), .B(n49329), .Z(n48898) );
  XOR U64418 ( .A(n48896), .B(n48898), .Z(n48904) );
  XOR U64419 ( .A(n44116), .B(n48904), .Z(n44514) );
  IV U64420 ( .A(n44117), .Z(n44119) );
  NOR U64421 ( .A(n44119), .B(n44118), .Z(n48906) );
  IV U64422 ( .A(n44120), .Z(n44121) );
  NOR U64423 ( .A(n44122), .B(n44121), .Z(n44513) );
  NOR U64424 ( .A(n48906), .B(n44513), .Z(n44123) );
  XOR U64425 ( .A(n44514), .B(n44123), .Z(n49315) );
  XOR U64426 ( .A(n44509), .B(n49315), .Z(n44511) );
  XOR U64427 ( .A(n44512), .B(n44511), .Z(n44507) );
  IV U64428 ( .A(n44124), .Z(n44125) );
  NOR U64429 ( .A(n44126), .B(n44125), .Z(n48917) );
  IV U64430 ( .A(n44127), .Z(n44128) );
  NOR U64431 ( .A(n44129), .B(n44128), .Z(n48913) );
  NOR U64432 ( .A(n48917), .B(n48913), .Z(n44508) );
  XOR U64433 ( .A(n44507), .B(n44508), .Z(n49303) );
  XOR U64434 ( .A(n48923), .B(n49303), .Z(n44505) );
  IV U64435 ( .A(n44130), .Z(n44131) );
  NOR U64436 ( .A(n44132), .B(n44131), .Z(n48924) );
  IV U64437 ( .A(n44133), .Z(n44134) );
  NOR U64438 ( .A(n44135), .B(n44134), .Z(n44504) );
  NOR U64439 ( .A(n48924), .B(n44504), .Z(n44136) );
  XOR U64440 ( .A(n44505), .B(n44136), .Z(n48934) );
  XOR U64441 ( .A(n48931), .B(n48934), .Z(n44502) );
  XOR U64442 ( .A(n44137), .B(n44502), .Z(n48942) );
  XOR U64443 ( .A(n48943), .B(n48942), .Z(n48945) );
  XOR U64444 ( .A(n48944), .B(n48945), .Z(n44138) );
  NOR U64445 ( .A(n44139), .B(n44138), .Z(n54091) );
  IV U64446 ( .A(n44140), .Z(n44142) );
  NOR U64447 ( .A(n44142), .B(n44141), .Z(n44499) );
  NOR U64448 ( .A(n48944), .B(n44499), .Z(n44143) );
  XOR U64449 ( .A(n44143), .B(n48945), .Z(n44144) );
  NOR U64450 ( .A(n44145), .B(n44144), .Z(n44146) );
  NOR U64451 ( .A(n54091), .B(n44146), .Z(n44493) );
  IV U64452 ( .A(n44147), .Z(n44149) );
  NOR U64453 ( .A(n44149), .B(n44148), .Z(n44496) );
  IV U64454 ( .A(n44150), .Z(n44151) );
  NOR U64455 ( .A(n44152), .B(n44151), .Z(n44492) );
  NOR U64456 ( .A(n44496), .B(n44492), .Z(n44153) );
  XOR U64457 ( .A(n44493), .B(n44153), .Z(n49286) );
  IV U64458 ( .A(n44154), .Z(n44156) );
  NOR U64459 ( .A(n44156), .B(n44155), .Z(n59761) );
  IV U64460 ( .A(n44157), .Z(n44158) );
  NOR U64461 ( .A(n44159), .B(n44158), .Z(n59748) );
  NOR U64462 ( .A(n59761), .B(n59748), .Z(n49288) );
  XOR U64463 ( .A(n49286), .B(n49288), .Z(n44160) );
  IV U64464 ( .A(n44160), .Z(n48950) );
  XOR U64465 ( .A(n48949), .B(n48950), .Z(n44173) );
  IV U64466 ( .A(n44173), .Z(n44169) );
  IV U64467 ( .A(n44161), .Z(n44162) );
  NOR U64468 ( .A(n44163), .B(n44162), .Z(n44170) );
  IV U64469 ( .A(n44164), .Z(n44166) );
  NOR U64470 ( .A(n44166), .B(n44165), .Z(n44172) );
  NOR U64471 ( .A(n44170), .B(n44172), .Z(n44167) );
  IV U64472 ( .A(n44167), .Z(n44168) );
  NOR U64473 ( .A(n44169), .B(n44168), .Z(n44176) );
  IV U64474 ( .A(n44170), .Z(n44171) );
  NOR U64475 ( .A(n44171), .B(n48950), .Z(n54096) );
  IV U64476 ( .A(n44172), .Z(n44174) );
  NOR U64477 ( .A(n44174), .B(n44173), .Z(n54104) );
  NOR U64478 ( .A(n54096), .B(n54104), .Z(n44175) );
  IV U64479 ( .A(n44175), .Z(n48956) );
  NOR U64480 ( .A(n44176), .B(n48956), .Z(n44177) );
  IV U64481 ( .A(n44177), .Z(n48959) );
  XOR U64482 ( .A(n48954), .B(n48959), .Z(n44490) );
  IV U64483 ( .A(n44178), .Z(n44180) );
  NOR U64484 ( .A(n44180), .B(n44179), .Z(n48958) );
  IV U64485 ( .A(n44181), .Z(n44182) );
  NOR U64486 ( .A(n44183), .B(n44182), .Z(n44489) );
  NOR U64487 ( .A(n48958), .B(n44489), .Z(n44184) );
  XOR U64488 ( .A(n44490), .B(n44184), .Z(n44485) );
  IV U64489 ( .A(n44185), .Z(n44186) );
  NOR U64490 ( .A(n44187), .B(n44186), .Z(n44486) );
  IV U64491 ( .A(n44188), .Z(n44189) );
  NOR U64492 ( .A(n44190), .B(n44189), .Z(n48963) );
  NOR U64493 ( .A(n44486), .B(n48963), .Z(n44191) );
  XOR U64494 ( .A(n44485), .B(n44191), .Z(n48967) );
  XOR U64495 ( .A(n48966), .B(n48967), .Z(n48973) );
  IV U64496 ( .A(n44192), .Z(n44194) );
  NOR U64497 ( .A(n44194), .B(n44193), .Z(n48961) );
  IV U64498 ( .A(n44195), .Z(n44197) );
  NOR U64499 ( .A(n44197), .B(n44196), .Z(n48972) );
  NOR U64500 ( .A(n48961), .B(n48972), .Z(n44198) );
  XOR U64501 ( .A(n48973), .B(n44198), .Z(n44478) );
  IV U64502 ( .A(n44199), .Z(n44200) );
  NOR U64503 ( .A(n44201), .B(n44200), .Z(n44479) );
  IV U64504 ( .A(n44202), .Z(n44203) );
  NOR U64505 ( .A(n44204), .B(n44203), .Z(n44481) );
  NOR U64506 ( .A(n44479), .B(n44481), .Z(n44205) );
  XOR U64507 ( .A(n44478), .B(n44205), .Z(n48978) );
  XOR U64508 ( .A(n44476), .B(n48978), .Z(n44474) );
  IV U64509 ( .A(n44206), .Z(n44208) );
  NOR U64510 ( .A(n44208), .B(n44207), .Z(n48977) );
  IV U64511 ( .A(n44209), .Z(n44210) );
  NOR U64512 ( .A(n44211), .B(n44210), .Z(n44473) );
  NOR U64513 ( .A(n48977), .B(n44473), .Z(n44212) );
  XOR U64514 ( .A(n44474), .B(n44212), .Z(n44471) );
  IV U64515 ( .A(n44213), .Z(n44215) );
  NOR U64516 ( .A(n44215), .B(n44214), .Z(n49272) );
  IV U64517 ( .A(n44216), .Z(n44218) );
  NOR U64518 ( .A(n44218), .B(n44217), .Z(n49263) );
  NOR U64519 ( .A(n49272), .B(n49263), .Z(n44472) );
  XOR U64520 ( .A(n44471), .B(n44472), .Z(n49269) );
  IV U64521 ( .A(n44219), .Z(n44220) );
  NOR U64522 ( .A(n44221), .B(n44220), .Z(n49267) );
  IV U64523 ( .A(n44222), .Z(n44224) );
  NOR U64524 ( .A(n44224), .B(n44223), .Z(n54142) );
  NOR U64525 ( .A(n49267), .B(n54142), .Z(n48989) );
  XOR U64526 ( .A(n49269), .B(n48989), .Z(n48990) );
  XOR U64527 ( .A(n48991), .B(n48990), .Z(n49000) );
  IV U64528 ( .A(n44225), .Z(n44226) );
  NOR U64529 ( .A(n44227), .B(n44226), .Z(n48997) );
  IV U64530 ( .A(n44228), .Z(n44229) );
  NOR U64531 ( .A(n44230), .B(n44229), .Z(n48999) );
  NOR U64532 ( .A(n48997), .B(n48999), .Z(n44231) );
  XOR U64533 ( .A(n49000), .B(n44231), .Z(n48995) );
  XOR U64534 ( .A(n44232), .B(n48995), .Z(n49007) );
  IV U64535 ( .A(n49007), .Z(n44233) );
  NOR U64536 ( .A(n49005), .B(n44233), .Z(n44238) );
  IV U64537 ( .A(n44234), .Z(n44235) );
  NOR U64538 ( .A(n44236), .B(n44235), .Z(n44240) );
  IV U64539 ( .A(n44240), .Z(n44237) );
  NOR U64540 ( .A(n44238), .B(n44237), .Z(n44470) );
  XOR U64541 ( .A(n49005), .B(n49007), .Z(n44468) );
  IV U64542 ( .A(n44468), .Z(n44239) );
  NOR U64543 ( .A(n44240), .B(n44239), .Z(n44241) );
  NOR U64544 ( .A(n44470), .B(n44241), .Z(n44242) );
  IV U64545 ( .A(n44242), .Z(n44464) );
  IV U64546 ( .A(n44461), .Z(n44243) );
  NOR U64547 ( .A(n44243), .B(n44459), .Z(n44247) );
  NOR U64548 ( .A(n44245), .B(n44244), .Z(n44246) );
  NOR U64549 ( .A(n44247), .B(n44246), .Z(n44462) );
  XOR U64550 ( .A(n44464), .B(n44462), .Z(n49244) );
  XOR U64551 ( .A(n49013), .B(n49244), .Z(n49014) );
  XOR U64552 ( .A(n49015), .B(n49014), .Z(n44456) );
  IV U64553 ( .A(n44248), .Z(n44249) );
  NOR U64554 ( .A(n44250), .B(n44249), .Z(n49018) );
  IV U64555 ( .A(n44251), .Z(n44253) );
  NOR U64556 ( .A(n44253), .B(n44252), .Z(n44455) );
  NOR U64557 ( .A(n49018), .B(n44455), .Z(n44254) );
  XOR U64558 ( .A(n44456), .B(n44254), .Z(n44255) );
  IV U64559 ( .A(n44255), .Z(n44454) );
  IV U64560 ( .A(n44256), .Z(n44258) );
  NOR U64561 ( .A(n44258), .B(n44257), .Z(n44259) );
  IV U64562 ( .A(n44259), .Z(n44266) );
  NOR U64563 ( .A(n44454), .B(n44266), .Z(n54162) );
  IV U64564 ( .A(n44260), .Z(n44262) );
  NOR U64565 ( .A(n44262), .B(n44261), .Z(n49024) );
  IV U64566 ( .A(n44263), .Z(n44265) );
  NOR U64567 ( .A(n44265), .B(n44264), .Z(n44452) );
  XOR U64568 ( .A(n44452), .B(n44454), .Z(n49025) );
  IV U64569 ( .A(n49025), .Z(n44267) );
  XOR U64570 ( .A(n49024), .B(n44267), .Z(n44269) );
  NOR U64571 ( .A(n44267), .B(n44266), .Z(n44268) );
  NOR U64572 ( .A(n44269), .B(n44268), .Z(n44270) );
  NOR U64573 ( .A(n54162), .B(n44270), .Z(n44275) );
  IV U64574 ( .A(n44275), .Z(n44450) );
  XOR U64575 ( .A(n44447), .B(n44450), .Z(n44271) );
  NOR U64576 ( .A(n44272), .B(n44271), .Z(n49231) );
  NOR U64577 ( .A(n44274), .B(n44273), .Z(n44449) );
  NOR U64578 ( .A(n44447), .B(n44449), .Z(n44276) );
  XOR U64579 ( .A(n44276), .B(n44275), .Z(n49033) );
  IV U64580 ( .A(n49033), .Z(n44277) );
  NOR U64581 ( .A(n44278), .B(n44277), .Z(n44279) );
  NOR U64582 ( .A(n49231), .B(n44279), .Z(n49036) );
  NOR U64583 ( .A(n44281), .B(n44280), .Z(n49032) );
  IV U64584 ( .A(n44282), .Z(n44284) );
  NOR U64585 ( .A(n44284), .B(n44283), .Z(n49035) );
  NOR U64586 ( .A(n49032), .B(n49035), .Z(n44285) );
  XOR U64587 ( .A(n49036), .B(n44285), .Z(n49228) );
  XOR U64588 ( .A(n49040), .B(n49228), .Z(n49041) );
  XOR U64589 ( .A(n44286), .B(n49041), .Z(n49056) );
  IV U64590 ( .A(n44287), .Z(n44289) );
  NOR U64591 ( .A(n44289), .B(n44288), .Z(n49047) );
  IV U64592 ( .A(n44290), .Z(n44292) );
  NOR U64593 ( .A(n44292), .B(n44291), .Z(n49055) );
  NOR U64594 ( .A(n49047), .B(n49055), .Z(n44293) );
  XOR U64595 ( .A(n49056), .B(n44293), .Z(n49053) );
  XOR U64596 ( .A(n49054), .B(n49053), .Z(n49213) );
  XOR U64597 ( .A(n44446), .B(n49213), .Z(n44441) );
  XOR U64598 ( .A(n44442), .B(n44441), .Z(n49061) );
  IV U64599 ( .A(n44294), .Z(n44295) );
  NOR U64600 ( .A(n44296), .B(n44295), .Z(n44443) );
  IV U64601 ( .A(n44297), .Z(n44299) );
  NOR U64602 ( .A(n44299), .B(n44298), .Z(n49060) );
  NOR U64603 ( .A(n44443), .B(n49060), .Z(n44300) );
  XOR U64604 ( .A(n49061), .B(n44300), .Z(n44435) );
  IV U64605 ( .A(n44301), .Z(n44303) );
  NOR U64606 ( .A(n44303), .B(n44302), .Z(n44438) );
  IV U64607 ( .A(n44304), .Z(n44305) );
  NOR U64608 ( .A(n44306), .B(n44305), .Z(n44436) );
  NOR U64609 ( .A(n44438), .B(n44436), .Z(n44307) );
  XOR U64610 ( .A(n44435), .B(n44307), .Z(n69931) );
  IV U64611 ( .A(n44308), .Z(n44310) );
  NOR U64612 ( .A(n44310), .B(n44309), .Z(n69930) );
  IV U64613 ( .A(n44311), .Z(n44312) );
  NOR U64614 ( .A(n44313), .B(n44312), .Z(n44314) );
  NOR U64615 ( .A(n69930), .B(n44314), .Z(n44432) );
  XOR U64616 ( .A(n69931), .B(n44432), .Z(n49067) );
  XOR U64617 ( .A(n44315), .B(n49067), .Z(n44425) );
  IV U64618 ( .A(n44316), .Z(n44317) );
  NOR U64619 ( .A(n44318), .B(n44317), .Z(n49071) );
  IV U64620 ( .A(n44319), .Z(n44321) );
  NOR U64621 ( .A(n44321), .B(n44320), .Z(n44424) );
  NOR U64622 ( .A(n49071), .B(n44424), .Z(n44322) );
  XOR U64623 ( .A(n44425), .B(n44322), .Z(n44323) );
  IV U64624 ( .A(n44323), .Z(n44431) );
  XOR U64625 ( .A(n44429), .B(n44431), .Z(n49082) );
  XOR U64626 ( .A(n44324), .B(n49082), .Z(n49078) );
  IV U64627 ( .A(n44325), .Z(n44326) );
  NOR U64628 ( .A(n44327), .B(n44326), .Z(n49079) );
  IV U64629 ( .A(n44328), .Z(n44329) );
  NOR U64630 ( .A(n44330), .B(n44329), .Z(n49086) );
  NOR U64631 ( .A(n49079), .B(n49086), .Z(n44331) );
  XOR U64632 ( .A(n49078), .B(n44331), .Z(n49091) );
  NOR U64633 ( .A(n44333), .B(n44332), .Z(n49084) );
  IV U64634 ( .A(n44334), .Z(n44336) );
  NOR U64635 ( .A(n44336), .B(n44335), .Z(n49090) );
  NOR U64636 ( .A(n49084), .B(n49090), .Z(n44337) );
  XOR U64637 ( .A(n49091), .B(n44337), .Z(n44420) );
  XOR U64638 ( .A(n44421), .B(n44420), .Z(n54298) );
  XOR U64639 ( .A(n44422), .B(n54298), .Z(n44410) );
  IV U64640 ( .A(n44338), .Z(n44340) );
  NOR U64641 ( .A(n44340), .B(n44339), .Z(n44409) );
  IV U64642 ( .A(n44341), .Z(n44342) );
  NOR U64643 ( .A(n44343), .B(n44342), .Z(n44412) );
  NOR U64644 ( .A(n44409), .B(n44412), .Z(n44344) );
  XOR U64645 ( .A(n44410), .B(n44344), .Z(n44417) );
  XOR U64646 ( .A(n44345), .B(n44417), .Z(n44346) );
  IV U64647 ( .A(n44346), .Z(n44406) );
  IV U64648 ( .A(n44347), .Z(n44349) );
  NOR U64649 ( .A(n44349), .B(n44348), .Z(n44405) );
  IV U64650 ( .A(n44350), .Z(n44352) );
  NOR U64651 ( .A(n44352), .B(n44351), .Z(n44401) );
  NOR U64652 ( .A(n44405), .B(n44401), .Z(n44353) );
  XOR U64653 ( .A(n44406), .B(n44353), .Z(n49150) );
  XOR U64654 ( .A(n49151), .B(n49150), .Z(n49143) );
  XOR U64655 ( .A(n49097), .B(n49143), .Z(n54208) );
  XOR U64656 ( .A(n49101), .B(n54208), .Z(n49103) );
  IV U64657 ( .A(n44354), .Z(n44356) );
  NOR U64658 ( .A(n44356), .B(n44355), .Z(n49110) );
  IV U64659 ( .A(n44357), .Z(n44358) );
  NOR U64660 ( .A(n44359), .B(n44358), .Z(n49102) );
  NOR U64661 ( .A(n49110), .B(n49102), .Z(n44360) );
  XOR U64662 ( .A(n49103), .B(n44360), .Z(n49109) );
  XOR U64663 ( .A(n49107), .B(n49109), .Z(n44398) );
  NOR U64664 ( .A(n44362), .B(n44361), .Z(n44399) );
  IV U64665 ( .A(n44363), .Z(n44364) );
  NOR U64666 ( .A(n44365), .B(n44364), .Z(n44396) );
  NOR U64667 ( .A(n44399), .B(n44396), .Z(n44366) );
  XOR U64668 ( .A(n44398), .B(n44366), .Z(n44392) );
  IV U64669 ( .A(n44367), .Z(n44368) );
  NOR U64670 ( .A(n44369), .B(n44368), .Z(n49116) );
  IV U64671 ( .A(n44370), .Z(n44372) );
  NOR U64672 ( .A(n44372), .B(n44371), .Z(n49114) );
  NOR U64673 ( .A(n49116), .B(n49114), .Z(n44373) );
  XOR U64674 ( .A(n44392), .B(n44373), .Z(n44391) );
  NOR U64675 ( .A(n44375), .B(n44374), .Z(n44393) );
  IV U64676 ( .A(n44376), .Z(n44377) );
  NOR U64677 ( .A(n44378), .B(n44377), .Z(n44389) );
  NOR U64678 ( .A(n44393), .B(n44389), .Z(n44379) );
  XOR U64679 ( .A(n44391), .B(n44379), .Z(n49124) );
  IV U64680 ( .A(n49124), .Z(n44388) );
  IV U64681 ( .A(n44380), .Z(n44382) );
  NOR U64682 ( .A(n44382), .B(n44381), .Z(n49121) );
  IV U64683 ( .A(n49121), .Z(n44383) );
  NOR U64684 ( .A(n44388), .B(n44383), .Z(n49133) );
  IV U64685 ( .A(n44384), .Z(n44386) );
  NOR U64686 ( .A(n44386), .B(n44385), .Z(n49122) );
  IV U64687 ( .A(n49122), .Z(n44387) );
  NOR U64688 ( .A(n44388), .B(n44387), .Z(n49130) );
  IV U64689 ( .A(n44389), .Z(n44390) );
  NOR U64690 ( .A(n44391), .B(n44390), .Z(n54240) );
  IV U64691 ( .A(n44392), .Z(n49118) );
  XOR U64692 ( .A(n49118), .B(n49116), .Z(n44395) );
  IV U64693 ( .A(n44393), .Z(n44394) );
  NOR U64694 ( .A(n44395), .B(n44394), .Z(n54236) );
  IV U64695 ( .A(n44396), .Z(n44397) );
  NOR U64696 ( .A(n44398), .B(n44397), .Z(n49136) );
  IV U64697 ( .A(n44399), .Z(n44400) );
  NOR U64698 ( .A(n49109), .B(n44400), .Z(n54225) );
  IV U64699 ( .A(n44401), .Z(n44402) );
  NOR U64700 ( .A(n44402), .B(n44406), .Z(n49147) );
  IV U64701 ( .A(n44403), .Z(n44404) );
  NOR U64702 ( .A(n44404), .B(n44417), .Z(n54285) );
  IV U64703 ( .A(n44405), .Z(n44407) );
  NOR U64704 ( .A(n44407), .B(n44406), .Z(n49156) );
  NOR U64705 ( .A(n54285), .B(n49156), .Z(n44408) );
  IV U64706 ( .A(n44408), .Z(n49095) );
  IV U64707 ( .A(n44409), .Z(n44411) );
  IV U64708 ( .A(n44410), .Z(n44413) );
  NOR U64709 ( .A(n44411), .B(n44413), .Z(n49163) );
  IV U64710 ( .A(n44412), .Z(n44414) );
  NOR U64711 ( .A(n44414), .B(n44413), .Z(n49161) );
  NOR U64712 ( .A(n49163), .B(n49161), .Z(n44415) );
  IV U64713 ( .A(n44415), .Z(n44419) );
  IV U64714 ( .A(n44416), .Z(n44418) );
  NOR U64715 ( .A(n44418), .B(n44417), .Z(n59503) );
  NOR U64716 ( .A(n44419), .B(n59503), .Z(n49094) );
  IV U64717 ( .A(n44420), .Z(n49168) );
  NOR U64718 ( .A(n49168), .B(n44421), .Z(n44423) );
  NOR U64719 ( .A(n44422), .B(n54298), .Z(n49165) );
  NOR U64720 ( .A(n44423), .B(n49165), .Z(n49093) );
  IV U64721 ( .A(n44424), .Z(n44426) );
  NOR U64722 ( .A(n44426), .B(n44425), .Z(n54194) );
  IV U64723 ( .A(n44427), .Z(n44428) );
  NOR U64724 ( .A(n44431), .B(n44428), .Z(n54197) );
  NOR U64725 ( .A(n54194), .B(n54197), .Z(n49076) );
  IV U64726 ( .A(n44429), .Z(n44430) );
  NOR U64727 ( .A(n44431), .B(n44430), .Z(n54192) );
  NOR U64728 ( .A(n44432), .B(n69931), .Z(n54308) );
  IV U64729 ( .A(n49068), .Z(n44433) );
  IV U64730 ( .A(n49067), .Z(n59457) );
  NOR U64731 ( .A(n44433), .B(n59457), .Z(n44434) );
  NOR U64732 ( .A(n54308), .B(n44434), .Z(n49188) );
  IV U64733 ( .A(n44435), .Z(n44440) );
  IV U64734 ( .A(n44436), .Z(n44437) );
  NOR U64735 ( .A(n44440), .B(n44437), .Z(n49193) );
  IV U64736 ( .A(n44438), .Z(n44439) );
  NOR U64737 ( .A(n44440), .B(n44439), .Z(n49195) );
  NOR U64738 ( .A(n49193), .B(n49195), .Z(n49065) );
  IV U64739 ( .A(n44441), .Z(n49204) );
  NOR U64740 ( .A(n44442), .B(n49204), .Z(n44445) );
  IV U64741 ( .A(n44443), .Z(n44444) );
  NOR U64742 ( .A(n44444), .B(n49061), .Z(n49199) );
  NOR U64743 ( .A(n44445), .B(n49199), .Z(n49064) );
  NOR U64744 ( .A(n44446), .B(n49213), .Z(n49059) );
  IV U64745 ( .A(n44447), .Z(n44448) );
  NOR U64746 ( .A(n44448), .B(n44450), .Z(n65000) );
  IV U64747 ( .A(n44449), .Z(n44451) );
  NOR U64748 ( .A(n44451), .B(n44450), .Z(n69903) );
  NOR U64749 ( .A(n65000), .B(n69903), .Z(n49021) );
  IV U64750 ( .A(n44452), .Z(n44453) );
  NOR U64751 ( .A(n44454), .B(n44453), .Z(n54166) );
  IV U64752 ( .A(n44455), .Z(n44457) );
  NOR U64753 ( .A(n44457), .B(n44456), .Z(n44458) );
  IV U64754 ( .A(n44458), .Z(n54164) );
  IV U64755 ( .A(n44459), .Z(n44460) );
  NOR U64756 ( .A(n44461), .B(n44460), .Z(n44467) );
  IV U64757 ( .A(n44462), .Z(n44463) );
  NOR U64758 ( .A(n44464), .B(n44463), .Z(n44465) );
  IV U64759 ( .A(n44465), .Z(n44466) );
  NOR U64760 ( .A(n44467), .B(n44466), .Z(n49250) );
  IV U64761 ( .A(n44467), .Z(n44469) );
  NOR U64762 ( .A(n44469), .B(n44468), .Z(n49252) );
  NOR U64763 ( .A(n49250), .B(n49252), .Z(n49012) );
  IV U64764 ( .A(n44470), .Z(n49259) );
  IV U64765 ( .A(n44471), .Z(n49264) );
  NOR U64766 ( .A(n49264), .B(n44472), .Z(n48988) );
  IV U64767 ( .A(n44473), .Z(n44475) );
  NOR U64768 ( .A(n44475), .B(n44474), .Z(n48982) );
  IV U64769 ( .A(n44476), .Z(n44477) );
  NOR U64770 ( .A(n44477), .B(n48978), .Z(n49275) );
  IV U64771 ( .A(n44478), .Z(n44483) );
  IV U64772 ( .A(n44479), .Z(n44480) );
  NOR U64773 ( .A(n44483), .B(n44480), .Z(n48983) );
  IV U64774 ( .A(n44481), .Z(n44482) );
  NOR U64775 ( .A(n44483), .B(n44482), .Z(n49280) );
  XOR U64776 ( .A(n48983), .B(n49280), .Z(n44484) );
  NOR U64777 ( .A(n49275), .B(n44484), .Z(n48976) );
  IV U64778 ( .A(n44485), .Z(n48965) );
  IV U64779 ( .A(n44486), .Z(n44487) );
  NOR U64780 ( .A(n48965), .B(n44487), .Z(n44488) );
  IV U64781 ( .A(n44488), .Z(n54121) );
  IV U64782 ( .A(n44489), .Z(n44491) );
  NOR U64783 ( .A(n44491), .B(n44490), .Z(n54111) );
  IV U64784 ( .A(n44492), .Z(n44494) );
  IV U64785 ( .A(n44493), .Z(n44497) );
  NOR U64786 ( .A(n44494), .B(n44497), .Z(n44495) );
  IV U64787 ( .A(n44495), .Z(n49289) );
  IV U64788 ( .A(n44496), .Z(n44498) );
  NOR U64789 ( .A(n44498), .B(n44497), .Z(n49291) );
  NOR U64790 ( .A(n54091), .B(n49291), .Z(n48948) );
  IV U64791 ( .A(n44499), .Z(n44500) );
  NOR U64792 ( .A(n44500), .B(n48945), .Z(n54088) );
  IV U64793 ( .A(n44501), .Z(n44503) );
  NOR U64794 ( .A(n44503), .B(n44502), .Z(n48940) );
  IV U64795 ( .A(n48940), .Z(n48930) );
  IV U64796 ( .A(n44504), .Z(n44506) );
  IV U64797 ( .A(n44505), .Z(n48925) );
  NOR U64798 ( .A(n44506), .B(n48925), .Z(n54079) );
  IV U64799 ( .A(n44507), .Z(n48914) );
  NOR U64800 ( .A(n44508), .B(n48914), .Z(n48912) );
  IV U64801 ( .A(n44509), .Z(n44510) );
  NOR U64802 ( .A(n49315), .B(n44510), .Z(n54069) );
  NOR U64803 ( .A(n44512), .B(n44511), .Z(n49309) );
  NOR U64804 ( .A(n54069), .B(n49309), .Z(n48910) );
  IV U64805 ( .A(n44513), .Z(n44515) );
  IV U64806 ( .A(n44514), .Z(n48907) );
  NOR U64807 ( .A(n44515), .B(n48907), .Z(n44516) );
  IV U64808 ( .A(n44516), .Z(n54067) );
  IV U64809 ( .A(n44517), .Z(n44518) );
  NOR U64810 ( .A(n48891), .B(n44518), .Z(n49345) );
  NOR U64811 ( .A(n49352), .B(n44519), .Z(n44520) );
  IV U64812 ( .A(n44520), .Z(n44521) );
  NOR U64813 ( .A(n44522), .B(n44521), .Z(n44525) );
  NOR U64814 ( .A(n49349), .B(n44523), .Z(n44524) );
  NOR U64815 ( .A(n44525), .B(n44524), .Z(n48888) );
  IV U64816 ( .A(n44526), .Z(n54047) );
  NOR U64817 ( .A(n54047), .B(n44527), .Z(n44531) );
  IV U64818 ( .A(n44528), .Z(n44530) );
  NOR U64819 ( .A(n44530), .B(n44529), .Z(n49363) );
  NOR U64820 ( .A(n44531), .B(n49363), .Z(n44532) );
  IV U64821 ( .A(n44532), .Z(n48887) );
  IV U64822 ( .A(n44533), .Z(n44535) );
  NOR U64823 ( .A(n44535), .B(n44534), .Z(n54043) );
  IV U64824 ( .A(n44536), .Z(n44538) );
  NOR U64825 ( .A(n44538), .B(n44537), .Z(n48877) );
  IV U64826 ( .A(n44539), .Z(n44540) );
  NOR U64827 ( .A(n44540), .B(n44543), .Z(n44541) );
  IV U64828 ( .A(n44541), .Z(n49373) );
  IV U64829 ( .A(n44542), .Z(n44544) );
  NOR U64830 ( .A(n44544), .B(n44543), .Z(n49369) );
  IV U64831 ( .A(n44545), .Z(n44548) );
  IV U64832 ( .A(n44546), .Z(n44547) );
  NOR U64833 ( .A(n44548), .B(n44547), .Z(n49388) );
  IV U64834 ( .A(n44549), .Z(n44552) );
  IV U64835 ( .A(n44550), .Z(n44551) );
  NOR U64836 ( .A(n44552), .B(n44551), .Z(n54031) );
  NOR U64837 ( .A(n54018), .B(n44553), .Z(n44556) );
  IV U64838 ( .A(n44554), .Z(n44555) );
  NOR U64839 ( .A(n44555), .B(n48842), .Z(n54020) );
  NOR U64840 ( .A(n44556), .B(n54020), .Z(n48833) );
  IV U64841 ( .A(n54008), .Z(n44557) );
  NOR U64842 ( .A(n44557), .B(n44558), .Z(n54005) );
  IV U64843 ( .A(n54011), .Z(n44559) );
  NOR U64844 ( .A(n44559), .B(n44558), .Z(n54002) );
  NOR U64845 ( .A(n54005), .B(n54002), .Z(n44560) );
  IV U64846 ( .A(n44560), .Z(n54013) );
  IV U64847 ( .A(n53972), .Z(n49408) );
  NOR U64848 ( .A(n49408), .B(n53970), .Z(n53974) );
  NOR U64849 ( .A(n44562), .B(n44561), .Z(n44563) );
  NOR U64850 ( .A(n53974), .B(n44563), .Z(n48813) );
  IV U64851 ( .A(n44564), .Z(n44566) );
  NOR U64852 ( .A(n44566), .B(n44565), .Z(n53949) );
  IV U64853 ( .A(n44567), .Z(n44570) );
  IV U64854 ( .A(n44568), .Z(n44569) );
  NOR U64855 ( .A(n44570), .B(n44569), .Z(n53948) );
  NOR U64856 ( .A(n53956), .B(n49411), .Z(n65163) );
  IV U64857 ( .A(n65163), .Z(n44571) );
  NOR U64858 ( .A(n53948), .B(n44571), .Z(n44572) );
  IV U64859 ( .A(n44572), .Z(n48812) );
  IV U64860 ( .A(n44573), .Z(n44574) );
  NOR U64861 ( .A(n44574), .B(n44579), .Z(n49414) );
  IV U64862 ( .A(n44575), .Z(n44583) );
  IV U64863 ( .A(n44576), .Z(n44577) );
  NOR U64864 ( .A(n44583), .B(n44577), .Z(n53943) );
  NOR U64865 ( .A(n49414), .B(n53943), .Z(n44585) );
  IV U64866 ( .A(n44578), .Z(n44580) );
  NOR U64867 ( .A(n44580), .B(n44579), .Z(n49416) );
  IV U64868 ( .A(n44581), .Z(n44582) );
  NOR U64869 ( .A(n44583), .B(n44582), .Z(n53945) );
  NOR U64870 ( .A(n49416), .B(n53945), .Z(n44584) );
  XOR U64871 ( .A(n44585), .B(n44584), .Z(n48811) );
  IV U64872 ( .A(n44586), .Z(n49424) );
  NOR U64873 ( .A(n49424), .B(n44587), .Z(n44590) );
  IV U64874 ( .A(n44588), .Z(n44589) );
  NOR U64875 ( .A(n44589), .B(n48806), .Z(n49419) );
  NOR U64876 ( .A(n44590), .B(n49419), .Z(n48810) );
  IV U64877 ( .A(n44591), .Z(n44593) );
  NOR U64878 ( .A(n44593), .B(n44592), .Z(n49432) );
  IV U64879 ( .A(n44594), .Z(n49460) );
  NOR U64880 ( .A(n49460), .B(n49458), .Z(n48770) );
  IV U64881 ( .A(n44595), .Z(n44596) );
  NOR U64882 ( .A(n44596), .B(n48768), .Z(n49461) );
  IV U64883 ( .A(n44597), .Z(n44599) );
  IV U64884 ( .A(n44598), .Z(n44601) );
  NOR U64885 ( .A(n44599), .B(n44601), .Z(n49469) );
  IV U64886 ( .A(n44600), .Z(n44602) );
  NOR U64887 ( .A(n44602), .B(n44601), .Z(n49466) );
  XOR U64888 ( .A(n49469), .B(n49466), .Z(n44603) );
  NOR U64889 ( .A(n49461), .B(n44603), .Z(n48763) );
  IV U64890 ( .A(n44604), .Z(n44605) );
  NOR U64891 ( .A(n44605), .B(n44609), .Z(n53924) );
  IV U64892 ( .A(n44606), .Z(n49484) );
  NOR U64893 ( .A(n44607), .B(n49484), .Z(n44611) );
  IV U64894 ( .A(n44608), .Z(n44610) );
  NOR U64895 ( .A(n44610), .B(n44609), .Z(n49479) );
  NOR U64896 ( .A(n44611), .B(n49479), .Z(n44612) );
  IV U64897 ( .A(n44612), .Z(n48752) );
  IV U64898 ( .A(n44613), .Z(n44614) );
  NOR U64899 ( .A(n44614), .B(n48723), .Z(n48720) );
  IV U64900 ( .A(n48720), .Z(n48711) );
  NOR U64901 ( .A(n44616), .B(n44615), .Z(n48706) );
  IV U64902 ( .A(n44617), .Z(n53909) );
  IV U64903 ( .A(n44618), .Z(n44619) );
  NOR U64904 ( .A(n53909), .B(n44619), .Z(n53905) );
  IV U64905 ( .A(n53910), .Z(n44620) );
  NOR U64906 ( .A(n53909), .B(n44620), .Z(n49509) );
  NOR U64907 ( .A(n53905), .B(n49509), .Z(n48705) );
  IV U64908 ( .A(n44621), .Z(n44622) );
  NOR U64909 ( .A(n44622), .B(n48703), .Z(n48699) );
  IV U64910 ( .A(n48699), .Z(n48685) );
  IV U64911 ( .A(n44623), .Z(n44625) );
  IV U64912 ( .A(n44624), .Z(n44639) );
  NOR U64913 ( .A(n44625), .B(n44639), .Z(n49522) );
  IV U64914 ( .A(n44626), .Z(n44628) );
  XOR U64915 ( .A(n44638), .B(n44639), .Z(n44627) );
  NOR U64916 ( .A(n44628), .B(n44627), .Z(n49519) );
  NOR U64917 ( .A(n49522), .B(n49519), .Z(n44629) );
  IV U64918 ( .A(n44629), .Z(n48692) );
  XOR U64919 ( .A(n44631), .B(n44630), .Z(n44632) );
  NOR U64920 ( .A(n44633), .B(n44632), .Z(n44634) );
  IV U64921 ( .A(n44634), .Z(n44636) );
  NOR U64922 ( .A(n44636), .B(n44635), .Z(n49517) );
  NOR U64923 ( .A(n48692), .B(n49517), .Z(n48684) );
  NOR U64924 ( .A(n44637), .B(n53888), .Z(n44641) );
  IV U64925 ( .A(n44638), .Z(n44640) );
  NOR U64926 ( .A(n44640), .B(n44639), .Z(n49529) );
  NOR U64927 ( .A(n44641), .B(n49529), .Z(n49523) );
  IV U64928 ( .A(n44642), .Z(n44644) );
  NOR U64929 ( .A(n44644), .B(n44643), .Z(n49541) );
  NOR U64930 ( .A(n44645), .B(n49533), .Z(n44646) );
  NOR U64931 ( .A(n49541), .B(n44646), .Z(n48674) );
  IV U64932 ( .A(n44647), .Z(n44648) );
  NOR U64933 ( .A(n48641), .B(n44648), .Z(n48647) );
  IV U64934 ( .A(n48647), .Z(n48633) );
  IV U64935 ( .A(n44649), .Z(n44650) );
  NOR U64936 ( .A(n44650), .B(n48628), .Z(n48637) );
  IV U64937 ( .A(n48637), .Z(n49562) );
  IV U64938 ( .A(n44651), .Z(n44652) );
  NOR U64939 ( .A(n44652), .B(n44654), .Z(n53858) );
  IV U64940 ( .A(n44653), .Z(n44655) );
  NOR U64941 ( .A(n44655), .B(n44654), .Z(n48622) );
  IV U64942 ( .A(n48622), .Z(n48607) );
  IV U64943 ( .A(n44656), .Z(n44658) );
  NOR U64944 ( .A(n44658), .B(n44657), .Z(n44659) );
  IV U64945 ( .A(n44659), .Z(n53856) );
  IV U64946 ( .A(n44660), .Z(n44661) );
  NOR U64947 ( .A(n44661), .B(n44663), .Z(n53851) );
  IV U64948 ( .A(n44662), .Z(n44664) );
  NOR U64949 ( .A(n44664), .B(n44663), .Z(n53848) );
  IV U64950 ( .A(n44665), .Z(n44669) );
  NOR U64951 ( .A(n44667), .B(n44666), .Z(n44668) );
  IV U64952 ( .A(n44668), .Z(n54707) );
  NOR U64953 ( .A(n44669), .B(n54707), .Z(n49569) );
  IV U64954 ( .A(n44670), .Z(n44674) );
  IV U64955 ( .A(n44671), .Z(n44672) );
  NOR U64956 ( .A(n44674), .B(n44672), .Z(n53843) );
  IV U64957 ( .A(n54713), .Z(n44673) );
  NOR U64958 ( .A(n44674), .B(n44673), .Z(n53840) );
  NOR U64959 ( .A(n44675), .B(n49580), .Z(n48581) );
  IV U64960 ( .A(n44676), .Z(n44677) );
  NOR U64961 ( .A(n44677), .B(n44681), .Z(n53811) );
  IV U64962 ( .A(n44678), .Z(n60041) );
  NOR U64963 ( .A(n60041), .B(n44679), .Z(n59065) );
  IV U64964 ( .A(n44680), .Z(n44682) );
  NOR U64965 ( .A(n44682), .B(n44681), .Z(n49599) );
  NOR U64966 ( .A(n59065), .B(n49599), .Z(n48566) );
  XOR U64967 ( .A(n44684), .B(n44683), .Z(n44685) );
  NOR U64968 ( .A(n44686), .B(n44685), .Z(n44687) );
  IV U64969 ( .A(n44687), .Z(n44690) );
  IV U64970 ( .A(n44688), .Z(n44689) );
  NOR U64971 ( .A(n44690), .B(n44689), .Z(n53774) );
  IV U64972 ( .A(n44691), .Z(n44694) );
  IV U64973 ( .A(n44692), .Z(n44693) );
  NOR U64974 ( .A(n44694), .B(n44693), .Z(n49612) );
  IV U64975 ( .A(n44695), .Z(n44696) );
  NOR U64976 ( .A(n44696), .B(n44699), .Z(n53766) );
  NOR U64977 ( .A(n53758), .B(n44697), .Z(n44701) );
  IV U64978 ( .A(n44698), .Z(n44700) );
  NOR U64979 ( .A(n44700), .B(n44699), .Z(n49616) );
  NOR U64980 ( .A(n44701), .B(n49616), .Z(n48536) );
  IV U64981 ( .A(n44702), .Z(n44703) );
  NOR U64982 ( .A(n44703), .B(n48513), .Z(n48518) );
  IV U64983 ( .A(n48518), .Z(n48509) );
  IV U64984 ( .A(n44704), .Z(n49626) );
  IV U64985 ( .A(n44705), .Z(n44706) );
  NOR U64986 ( .A(n49626), .B(n44706), .Z(n59012) );
  IV U64987 ( .A(n44707), .Z(n44708) );
  NOR U64988 ( .A(n44708), .B(n44710), .Z(n49629) );
  NOR U64989 ( .A(n59012), .B(n49629), .Z(n48491) );
  IV U64990 ( .A(n44709), .Z(n44711) );
  NOR U64991 ( .A(n44711), .B(n44710), .Z(n44712) );
  IV U64992 ( .A(n44712), .Z(n49631) );
  IV U64993 ( .A(n44713), .Z(n48474) );
  IV U64994 ( .A(n44714), .Z(n44715) );
  NOR U64995 ( .A(n48474), .B(n44715), .Z(n49642) );
  IV U64996 ( .A(n44716), .Z(n44718) );
  NOR U64997 ( .A(n44718), .B(n44717), .Z(n49646) );
  NOR U64998 ( .A(n49642), .B(n49646), .Z(n48477) );
  IV U64999 ( .A(n44719), .Z(n44720) );
  NOR U65000 ( .A(n44724), .B(n44720), .Z(n44721) );
  IV U65001 ( .A(n44721), .Z(n49648) );
  IV U65002 ( .A(n44722), .Z(n44723) );
  NOR U65003 ( .A(n44724), .B(n44723), .Z(n49650) );
  IV U65004 ( .A(n44725), .Z(n75822) );
  NOR U65005 ( .A(n75822), .B(n53737), .Z(n53741) );
  NOR U65006 ( .A(n49650), .B(n53741), .Z(n48471) );
  IV U65007 ( .A(n44729), .Z(n49655) );
  NOR U65008 ( .A(n44727), .B(n49655), .Z(n44726) );
  NOR U65009 ( .A(n53739), .B(n44726), .Z(n44731) );
  IV U65010 ( .A(n44727), .Z(n44728) );
  NOR U65011 ( .A(n44729), .B(n44728), .Z(n44730) );
  NOR U65012 ( .A(n44731), .B(n44730), .Z(n48470) );
  IV U65013 ( .A(n44732), .Z(n53732) );
  IV U65014 ( .A(n44733), .Z(n44734) );
  NOR U65015 ( .A(n53732), .B(n44734), .Z(n53727) );
  IV U65016 ( .A(n44735), .Z(n44737) );
  NOR U65017 ( .A(n44737), .B(n44736), .Z(n53724) );
  IV U65018 ( .A(n44738), .Z(n44739) );
  NOR U65019 ( .A(n44739), .B(n44741), .Z(n53717) );
  IV U65020 ( .A(n44740), .Z(n44742) );
  NOR U65021 ( .A(n44742), .B(n44741), .Z(n53720) );
  XOR U65022 ( .A(n53717), .B(n53720), .Z(n44743) );
  NOR U65023 ( .A(n53724), .B(n44743), .Z(n48469) );
  NOR U65024 ( .A(n44744), .B(n49660), .Z(n44747) );
  IV U65025 ( .A(n44745), .Z(n53713) );
  NOR U65026 ( .A(n53716), .B(n53713), .Z(n44746) );
  NOR U65027 ( .A(n44747), .B(n44746), .Z(n48468) );
  IV U65028 ( .A(n44748), .Z(n49665) );
  NOR U65029 ( .A(n49665), .B(n44749), .Z(n48467) );
  IV U65030 ( .A(n44750), .Z(n44753) );
  IV U65031 ( .A(n44751), .Z(n44752) );
  NOR U65032 ( .A(n44753), .B(n44752), .Z(n53672) );
  IV U65033 ( .A(n44754), .Z(n44755) );
  NOR U65034 ( .A(n44757), .B(n44755), .Z(n44758) );
  IV U65035 ( .A(n49686), .Z(n44756) );
  NOR U65036 ( .A(n44757), .B(n44756), .Z(n53665) );
  NOR U65037 ( .A(n44758), .B(n53665), .Z(n49683) );
  IV U65038 ( .A(n44759), .Z(n44762) );
  IV U65039 ( .A(n44760), .Z(n44761) );
  NOR U65040 ( .A(n44762), .B(n44761), .Z(n44763) );
  IV U65041 ( .A(n44763), .Z(n53662) );
  IV U65042 ( .A(n44764), .Z(n44766) );
  NOR U65043 ( .A(n44766), .B(n44765), .Z(n48432) );
  IV U65044 ( .A(n44767), .Z(n44769) );
  NOR U65045 ( .A(n44769), .B(n44768), .Z(n49693) );
  IV U65046 ( .A(n44770), .Z(n44773) );
  IV U65047 ( .A(n44771), .Z(n44772) );
  NOR U65048 ( .A(n44773), .B(n44772), .Z(n48410) );
  IV U65049 ( .A(n44774), .Z(n44777) );
  IV U65050 ( .A(n44775), .Z(n44776) );
  NOR U65051 ( .A(n44777), .B(n44776), .Z(n44778) );
  IV U65052 ( .A(n44778), .Z(n53652) );
  IV U65053 ( .A(n44779), .Z(n44780) );
  NOR U65054 ( .A(n44780), .B(n44782), .Z(n49699) );
  IV U65055 ( .A(n44781), .Z(n44783) );
  NOR U65056 ( .A(n44783), .B(n44782), .Z(n49701) );
  NOR U65057 ( .A(n49699), .B(n49701), .Z(n48407) );
  IV U65058 ( .A(n44784), .Z(n44792) );
  IV U65059 ( .A(n44785), .Z(n44786) );
  NOR U65060 ( .A(n44792), .B(n44786), .Z(n53622) );
  NOR U65061 ( .A(n44787), .B(n49705), .Z(n44788) );
  NOR U65062 ( .A(n53622), .B(n44788), .Z(n44789) );
  IV U65063 ( .A(n44789), .Z(n48406) );
  IV U65064 ( .A(n44790), .Z(n44791) );
  NOR U65065 ( .A(n44792), .B(n44791), .Z(n53627) );
  IV U65066 ( .A(n44793), .Z(n44795) );
  NOR U65067 ( .A(n44795), .B(n44794), .Z(n53629) );
  NOR U65068 ( .A(n53627), .B(n53629), .Z(n48405) );
  IV U65069 ( .A(n44796), .Z(n44797) );
  NOR U65070 ( .A(n44800), .B(n44797), .Z(n53618) );
  IV U65071 ( .A(n44798), .Z(n44799) );
  NOR U65072 ( .A(n44800), .B(n44799), .Z(n49708) );
  NOR U65073 ( .A(n53618), .B(n49708), .Z(n48404) );
  IV U65074 ( .A(n44801), .Z(n44803) );
  NOR U65075 ( .A(n44803), .B(n44802), .Z(n53615) );
  IV U65076 ( .A(n44804), .Z(n44807) );
  IV U65077 ( .A(n44805), .Z(n44812) );
  XOR U65078 ( .A(n44812), .B(n44809), .Z(n44806) );
  NOR U65079 ( .A(n44807), .B(n44806), .Z(n53612) );
  IV U65080 ( .A(n44808), .Z(n44810) );
  IV U65081 ( .A(n44809), .Z(n44811) );
  NOR U65082 ( .A(n44810), .B(n44811), .Z(n53608) );
  NOR U65083 ( .A(n44812), .B(n44811), .Z(n53605) );
  IV U65084 ( .A(n44813), .Z(n44814) );
  NOR U65085 ( .A(n44817), .B(n44814), .Z(n53599) );
  NOR U65086 ( .A(n53605), .B(n53599), .Z(n48403) );
  IV U65087 ( .A(n44815), .Z(n44816) );
  NOR U65088 ( .A(n44817), .B(n44816), .Z(n53601) );
  IV U65089 ( .A(n44818), .Z(n44821) );
  IV U65090 ( .A(n44819), .Z(n44820) );
  NOR U65091 ( .A(n44821), .B(n44820), .Z(n49710) );
  NOR U65092 ( .A(n53601), .B(n49710), .Z(n48402) );
  IV U65093 ( .A(n44822), .Z(n44824) );
  XOR U65094 ( .A(n44827), .B(n44828), .Z(n44823) );
  NOR U65095 ( .A(n44824), .B(n44823), .Z(n49715) );
  IV U65096 ( .A(n44825), .Z(n44826) );
  NOR U65097 ( .A(n44826), .B(n44828), .Z(n49712) );
  IV U65098 ( .A(n44827), .Z(n44829) );
  NOR U65099 ( .A(n44829), .B(n44828), .Z(n53586) );
  NOR U65100 ( .A(n44830), .B(n64089), .Z(n49718) );
  IV U65101 ( .A(n44831), .Z(n53582) );
  NOR U65102 ( .A(n44832), .B(n53582), .Z(n44833) );
  NOR U65103 ( .A(n49718), .B(n44833), .Z(n54918) );
  IV U65104 ( .A(n54918), .Z(n48401) );
  IV U65105 ( .A(n44834), .Z(n44836) );
  NOR U65106 ( .A(n44836), .B(n44835), .Z(n53551) );
  IV U65107 ( .A(n44837), .Z(n44838) );
  NOR U65108 ( .A(n48379), .B(n44838), .Z(n49726) );
  IV U65109 ( .A(n44839), .Z(n44842) );
  IV U65110 ( .A(n44840), .Z(n44841) );
  NOR U65111 ( .A(n44842), .B(n44841), .Z(n53531) );
  IV U65112 ( .A(n44843), .Z(n44845) );
  IV U65113 ( .A(n44844), .Z(n44847) );
  NOR U65114 ( .A(n44845), .B(n44847), .Z(n49771) );
  NOR U65115 ( .A(n49773), .B(n49771), .Z(n48318) );
  IV U65116 ( .A(n44846), .Z(n44848) );
  NOR U65117 ( .A(n44848), .B(n44847), .Z(n49769) );
  IV U65118 ( .A(n44849), .Z(n44850) );
  NOR U65119 ( .A(n44850), .B(n48314), .Z(n49776) );
  IV U65120 ( .A(n44851), .Z(n44852) );
  NOR U65121 ( .A(n44855), .B(n44852), .Z(n49794) );
  IV U65122 ( .A(n44853), .Z(n44854) );
  NOR U65123 ( .A(n44855), .B(n44854), .Z(n49788) );
  NOR U65124 ( .A(n49794), .B(n49788), .Z(n44856) );
  IV U65125 ( .A(n44856), .Z(n48302) );
  IV U65126 ( .A(n48293), .Z(n44857) );
  NOR U65127 ( .A(n48292), .B(n44857), .Z(n49800) );
  IV U65128 ( .A(n44858), .Z(n44860) );
  NOR U65129 ( .A(n44860), .B(n44859), .Z(n53462) );
  IV U65130 ( .A(n44861), .Z(n44862) );
  NOR U65131 ( .A(n48260), .B(n44862), .Z(n49824) );
  XOR U65132 ( .A(n54984), .B(n49824), .Z(n44863) );
  NOR U65133 ( .A(n53462), .B(n44863), .Z(n48265) );
  IV U65134 ( .A(n44864), .Z(n44867) );
  NOR U65135 ( .A(n44865), .B(n44867), .Z(n60332) );
  IV U65136 ( .A(n44866), .Z(n44868) );
  NOR U65137 ( .A(n44868), .B(n44867), .Z(n63977) );
  NOR U65138 ( .A(n60332), .B(n63977), .Z(n53455) );
  IV U65139 ( .A(n44869), .Z(n49832) );
  NOR U65140 ( .A(n49834), .B(n49832), .Z(n44871) );
  NOR U65141 ( .A(n44870), .B(n53445), .Z(n49830) );
  NOR U65142 ( .A(n44871), .B(n49830), .Z(n48257) );
  IV U65143 ( .A(n44872), .Z(n44874) );
  NOR U65144 ( .A(n44874), .B(n44873), .Z(n44875) );
  IV U65145 ( .A(n44875), .Z(n53420) );
  NOR U65146 ( .A(n44878), .B(n44876), .Z(n53414) );
  NOR U65147 ( .A(n44878), .B(n44877), .Z(n53411) );
  IV U65148 ( .A(n44879), .Z(n44881) );
  IV U65149 ( .A(n44880), .Z(n44883) );
  NOR U65150 ( .A(n44881), .B(n44883), .Z(n49836) );
  IV U65151 ( .A(n44882), .Z(n44884) );
  NOR U65152 ( .A(n44884), .B(n44883), .Z(n49837) );
  XOR U65153 ( .A(n49836), .B(n49837), .Z(n44885) );
  NOR U65154 ( .A(n53411), .B(n44885), .Z(n48245) );
  IV U65155 ( .A(n44886), .Z(n44887) );
  NOR U65156 ( .A(n48239), .B(n44887), .Z(n49840) );
  IV U65157 ( .A(n44888), .Z(n44891) );
  IV U65158 ( .A(n44889), .Z(n44890) );
  NOR U65159 ( .A(n44891), .B(n44890), .Z(n49846) );
  NOR U65160 ( .A(n49851), .B(n49846), .Z(n48236) );
  IV U65161 ( .A(n44892), .Z(n44893) );
  NOR U65162 ( .A(n44896), .B(n44893), .Z(n49856) );
  IV U65163 ( .A(n44894), .Z(n44895) );
  NOR U65164 ( .A(n44896), .B(n44895), .Z(n49854) );
  NOR U65165 ( .A(n49856), .B(n49854), .Z(n48234) );
  NOR U65166 ( .A(n49867), .B(n44897), .Z(n44901) );
  IV U65167 ( .A(n44898), .Z(n44900) );
  IV U65168 ( .A(n44899), .Z(n44907) );
  NOR U65169 ( .A(n44900), .B(n44907), .Z(n49860) );
  NOR U65170 ( .A(n44901), .B(n49860), .Z(n48233) );
  XOR U65171 ( .A(n44903), .B(n44902), .Z(n44904) );
  NOR U65172 ( .A(n44905), .B(n44904), .Z(n44906) );
  IV U65173 ( .A(n44906), .Z(n44908) );
  NOR U65174 ( .A(n44908), .B(n44907), .Z(n44909) );
  IV U65175 ( .A(n44909), .Z(n49859) );
  IV U65176 ( .A(n44910), .Z(n44913) );
  IV U65177 ( .A(n44911), .Z(n44912) );
  NOR U65178 ( .A(n44913), .B(n44912), .Z(n49863) );
  IV U65179 ( .A(n44914), .Z(n44916) );
  XOR U65180 ( .A(n44919), .B(n44921), .Z(n44915) );
  NOR U65181 ( .A(n44916), .B(n44915), .Z(n53403) );
  IV U65182 ( .A(n44917), .Z(n44918) );
  NOR U65183 ( .A(n44921), .B(n44918), .Z(n53400) );
  IV U65184 ( .A(n44919), .Z(n44920) );
  NOR U65185 ( .A(n44921), .B(n44920), .Z(n53393) );
  NOR U65186 ( .A(n44923), .B(n44922), .Z(n44926) );
  NOR U65187 ( .A(n49877), .B(n44924), .Z(n44925) );
  NOR U65188 ( .A(n44926), .B(n44925), .Z(n48231) );
  IV U65189 ( .A(n44927), .Z(n44929) );
  NOR U65190 ( .A(n44929), .B(n44928), .Z(n49880) );
  IV U65191 ( .A(n44930), .Z(n44932) );
  NOR U65192 ( .A(n44932), .B(n44931), .Z(n49897) );
  IV U65193 ( .A(n44933), .Z(n44934) );
  NOR U65194 ( .A(n44934), .B(n44936), .Z(n49902) );
  IV U65195 ( .A(n44935), .Z(n44937) );
  NOR U65196 ( .A(n44937), .B(n44936), .Z(n53381) );
  NOR U65197 ( .A(n49902), .B(n53381), .Z(n48207) );
  IV U65198 ( .A(n44938), .Z(n44940) );
  IV U65199 ( .A(n44939), .Z(n48203) );
  NOR U65200 ( .A(n44940), .B(n48203), .Z(n49912) );
  NOR U65201 ( .A(n44941), .B(n49906), .Z(n44942) );
  NOR U65202 ( .A(n49912), .B(n44942), .Z(n48206) );
  IV U65203 ( .A(n44943), .Z(n44945) );
  NOR U65204 ( .A(n44945), .B(n44944), .Z(n53369) );
  NOR U65205 ( .A(n53369), .B(n53376), .Z(n48198) );
  IV U65206 ( .A(n44946), .Z(n44948) );
  IV U65207 ( .A(n44947), .Z(n48195) );
  NOR U65208 ( .A(n44948), .B(n48195), .Z(n44949) );
  IV U65209 ( .A(n44949), .Z(n48190) );
  IV U65210 ( .A(n44950), .Z(n49929) );
  NOR U65211 ( .A(n49929), .B(n44951), .Z(n48188) );
  IV U65212 ( .A(n44952), .Z(n44954) );
  NOR U65213 ( .A(n44954), .B(n44953), .Z(n49932) );
  XOR U65214 ( .A(n44956), .B(n44955), .Z(n44957) );
  NOR U65215 ( .A(n44958), .B(n44957), .Z(n44959) );
  IV U65216 ( .A(n44959), .Z(n44961) );
  NOR U65217 ( .A(n44961), .B(n44960), .Z(n48171) );
  IV U65218 ( .A(n44962), .Z(n55086) );
  NOR U65219 ( .A(n44963), .B(n55086), .Z(n49939) );
  IV U65220 ( .A(n44964), .Z(n44965) );
  NOR U65221 ( .A(n44965), .B(n44967), .Z(n53334) );
  IV U65222 ( .A(n44966), .Z(n44968) );
  NOR U65223 ( .A(n44968), .B(n44967), .Z(n49949) );
  IV U65224 ( .A(n44969), .Z(n48133) );
  NOR U65225 ( .A(n48133), .B(n44970), .Z(n48131) );
  IV U65226 ( .A(n44971), .Z(n44972) );
  NOR U65227 ( .A(n44972), .B(n44974), .Z(n49960) );
  IV U65228 ( .A(n44973), .Z(n44975) );
  NOR U65229 ( .A(n44975), .B(n44974), .Z(n48125) );
  IV U65230 ( .A(n44976), .Z(n58581) );
  NOR U65231 ( .A(n58581), .B(n44977), .Z(n48122) );
  IV U65232 ( .A(n48122), .Z(n48114) );
  NOR U65233 ( .A(n49969), .B(n44978), .Z(n49967) );
  IV U65234 ( .A(n44978), .Z(n44979) );
  NOR U65235 ( .A(n44980), .B(n44979), .Z(n44983) );
  IV U65236 ( .A(n44981), .Z(n44982) );
  NOR U65237 ( .A(n44983), .B(n44982), .Z(n44984) );
  NOR U65238 ( .A(n49967), .B(n44984), .Z(n49964) );
  IV U65239 ( .A(n44985), .Z(n44987) );
  IV U65240 ( .A(n44986), .Z(n48112) );
  NOR U65241 ( .A(n44987), .B(n48112), .Z(n49972) );
  NOR U65242 ( .A(n44988), .B(n49979), .Z(n44996) );
  IV U65243 ( .A(n44989), .Z(n44991) );
  IV U65244 ( .A(n44990), .Z(n44993) );
  NOR U65245 ( .A(n44991), .B(n44993), .Z(n49990) );
  IV U65246 ( .A(n44992), .Z(n44994) );
  NOR U65247 ( .A(n44994), .B(n44993), .Z(n49988) );
  XOR U65248 ( .A(n49990), .B(n49988), .Z(n44995) );
  NOR U65249 ( .A(n44996), .B(n44995), .Z(n48109) );
  IV U65250 ( .A(n44997), .Z(n44999) );
  NOR U65251 ( .A(n44999), .B(n44998), .Z(n49993) );
  IV U65252 ( .A(n45000), .Z(n45002) );
  NOR U65253 ( .A(n45002), .B(n45001), .Z(n58543) );
  NOR U65254 ( .A(n58543), .B(n58536), .Z(n45003) );
  IV U65255 ( .A(n45003), .Z(n53310) );
  IV U65256 ( .A(n45004), .Z(n45005) );
  NOR U65257 ( .A(n45005), .B(n48099), .Z(n45006) );
  IV U65258 ( .A(n45006), .Z(n50000) );
  IV U65259 ( .A(n45007), .Z(n50005) );
  NOR U65260 ( .A(n50005), .B(n45008), .Z(n45012) );
  IV U65261 ( .A(n45009), .Z(n45011) );
  NOR U65262 ( .A(n45011), .B(n45010), .Z(n53299) );
  NOR U65263 ( .A(n45012), .B(n53299), .Z(n48094) );
  IV U65264 ( .A(n45013), .Z(n45014) );
  NOR U65265 ( .A(n45014), .B(n48057), .Z(n48072) );
  NOR U65266 ( .A(n45016), .B(n45015), .Z(n48048) );
  IV U65267 ( .A(n48048), .Z(n48040) );
  IV U65268 ( .A(n45017), .Z(n45019) );
  NOR U65269 ( .A(n45019), .B(n45018), .Z(n53279) );
  IV U65270 ( .A(n45020), .Z(n45021) );
  NOR U65271 ( .A(n45021), .B(n48010), .Z(n48017) );
  IV U65272 ( .A(n48017), .Z(n48008) );
  IV U65273 ( .A(n45022), .Z(n45023) );
  NOR U65274 ( .A(n45023), .B(n47981), .Z(n45024) );
  IV U65275 ( .A(n45024), .Z(n47988) );
  IV U65276 ( .A(n45025), .Z(n45026) );
  NOR U65277 ( .A(n45026), .B(n45031), .Z(n53265) );
  IV U65278 ( .A(n45027), .Z(n45029) );
  IV U65279 ( .A(n45028), .Z(n45034) );
  NOR U65280 ( .A(n45029), .B(n45034), .Z(n58484) );
  IV U65281 ( .A(n45030), .Z(n45032) );
  NOR U65282 ( .A(n45032), .B(n45031), .Z(n58490) );
  NOR U65283 ( .A(n58484), .B(n58490), .Z(n53262) );
  IV U65284 ( .A(n45033), .Z(n45035) );
  NOR U65285 ( .A(n45035), .B(n45034), .Z(n47968) );
  IV U65286 ( .A(n47968), .Z(n47961) );
  IV U65287 ( .A(n45036), .Z(n45038) );
  IV U65288 ( .A(n45037), .Z(n45041) );
  NOR U65289 ( .A(n45038), .B(n45041), .Z(n45039) );
  IV U65290 ( .A(n45039), .Z(n58482) );
  IV U65291 ( .A(n45040), .Z(n45042) );
  NOR U65292 ( .A(n45042), .B(n45041), .Z(n47959) );
  IV U65293 ( .A(n47959), .Z(n47949) );
  IV U65294 ( .A(n45043), .Z(n45046) );
  IV U65295 ( .A(n45044), .Z(n45045) );
  NOR U65296 ( .A(n45046), .B(n45045), .Z(n53256) );
  IV U65297 ( .A(n45047), .Z(n45049) );
  XOR U65298 ( .A(n47945), .B(n47946), .Z(n45048) );
  NOR U65299 ( .A(n45049), .B(n45048), .Z(n45050) );
  IV U65300 ( .A(n45050), .Z(n53251) );
  IV U65301 ( .A(n45051), .Z(n45052) );
  NOR U65302 ( .A(n47932), .B(n45052), .Z(n47939) );
  IV U65303 ( .A(n47923), .Z(n47915) );
  IV U65304 ( .A(n45053), .Z(n53235) );
  NOR U65305 ( .A(n45054), .B(n53235), .Z(n50055) );
  IV U65306 ( .A(n45055), .Z(n45057) );
  NOR U65307 ( .A(n45057), .B(n45056), .Z(n53230) );
  IV U65308 ( .A(n45058), .Z(n45061) );
  IV U65309 ( .A(n45059), .Z(n47909) );
  XOR U65310 ( .A(n47909), .B(n47908), .Z(n45060) );
  NOR U65311 ( .A(n45061), .B(n45060), .Z(n53227) );
  NOR U65312 ( .A(n45063), .B(n45062), .Z(n45064) );
  IV U65313 ( .A(n45064), .Z(n45065) );
  NOR U65314 ( .A(n47905), .B(n45065), .Z(n50060) );
  IV U65315 ( .A(n45066), .Z(n45067) );
  NOR U65316 ( .A(n45067), .B(n45069), .Z(n50076) );
  NOR U65317 ( .A(n50076), .B(n50071), .Z(n47893) );
  IV U65318 ( .A(n45068), .Z(n45070) );
  NOR U65319 ( .A(n45070), .B(n45069), .Z(n50073) );
  IV U65320 ( .A(n45071), .Z(n58393) );
  NOR U65321 ( .A(n58393), .B(n45072), .Z(n50079) );
  IV U65322 ( .A(n45073), .Z(n45075) );
  NOR U65323 ( .A(n45075), .B(n45074), .Z(n50084) );
  NOR U65324 ( .A(n50079), .B(n50084), .Z(n47890) );
  IV U65325 ( .A(n45076), .Z(n45077) );
  NOR U65326 ( .A(n45077), .B(n45079), .Z(n50081) );
  IV U65327 ( .A(n45078), .Z(n45080) );
  NOR U65328 ( .A(n45080), .B(n45079), .Z(n53213) );
  IV U65329 ( .A(n45081), .Z(n45082) );
  NOR U65330 ( .A(n45082), .B(n45084), .Z(n50093) );
  IV U65331 ( .A(n45083), .Z(n45085) );
  NOR U65332 ( .A(n45085), .B(n45084), .Z(n53196) );
  IV U65333 ( .A(n45088), .Z(n45086) );
  NOR U65334 ( .A(n45087), .B(n45086), .Z(n47815) );
  IV U65335 ( .A(n45087), .Z(n50105) );
  NOR U65336 ( .A(n45088), .B(n50105), .Z(n47826) );
  NOR U65337 ( .A(n55315), .B(n45089), .Z(n53149) );
  IV U65338 ( .A(n45090), .Z(n45093) );
  IV U65339 ( .A(n45091), .Z(n45092) );
  NOR U65340 ( .A(n45093), .B(n45092), .Z(n47810) );
  IV U65341 ( .A(n47810), .Z(n47801) );
  IV U65342 ( .A(n45094), .Z(n45097) );
  IV U65343 ( .A(n45095), .Z(n45096) );
  NOR U65344 ( .A(n45097), .B(n45096), .Z(n53140) );
  IV U65345 ( .A(n45098), .Z(n45100) );
  XOR U65346 ( .A(n47797), .B(n47798), .Z(n45099) );
  NOR U65347 ( .A(n45100), .B(n45099), .Z(n45101) );
  IV U65348 ( .A(n45101), .Z(n53138) );
  IV U65349 ( .A(n45102), .Z(n45104) );
  NOR U65350 ( .A(n45104), .B(n45103), .Z(n50116) );
  NOR U65351 ( .A(n50116), .B(n50113), .Z(n45105) );
  IV U65352 ( .A(n45105), .Z(n47787) );
  IV U65353 ( .A(n45106), .Z(n45107) );
  NOR U65354 ( .A(n45108), .B(n45107), .Z(n50121) );
  IV U65355 ( .A(n45109), .Z(n45111) );
  NOR U65356 ( .A(n45111), .B(n45110), .Z(n50118) );
  IV U65357 ( .A(n45112), .Z(n55339) );
  NOR U65358 ( .A(n55339), .B(n45113), .Z(n53097) );
  IV U65359 ( .A(n45114), .Z(n45116) );
  NOR U65360 ( .A(n45116), .B(n45115), .Z(n50127) );
  NOR U65361 ( .A(n53097), .B(n50127), .Z(n47785) );
  IV U65362 ( .A(n45117), .Z(n53088) );
  IV U65363 ( .A(n45118), .Z(n45122) );
  NOR U65364 ( .A(n45122), .B(n45119), .Z(n50137) );
  IV U65365 ( .A(n45120), .Z(n45121) );
  NOR U65366 ( .A(n45122), .B(n45121), .Z(n50134) );
  NOR U65367 ( .A(n50137), .B(n50134), .Z(n47768) );
  IV U65368 ( .A(n45123), .Z(n45125) );
  NOR U65369 ( .A(n45125), .B(n45124), .Z(n53080) );
  IV U65370 ( .A(n45126), .Z(n45129) );
  IV U65371 ( .A(n45127), .Z(n47764) );
  XOR U65372 ( .A(n47762), .B(n47764), .Z(n45128) );
  NOR U65373 ( .A(n45129), .B(n45128), .Z(n50140) );
  IV U65374 ( .A(n45130), .Z(n45131) );
  NOR U65375 ( .A(n47764), .B(n45131), .Z(n53067) );
  IV U65376 ( .A(n45132), .Z(n45133) );
  NOR U65377 ( .A(n45133), .B(n47765), .Z(n50146) );
  IV U65378 ( .A(n45134), .Z(n45139) );
  IV U65379 ( .A(n45135), .Z(n45136) );
  NOR U65380 ( .A(n45139), .B(n45136), .Z(n50148) );
  NOR U65381 ( .A(n50146), .B(n50148), .Z(n47761) );
  IV U65382 ( .A(n45137), .Z(n45138) );
  NOR U65383 ( .A(n45139), .B(n45138), .Z(n53055) );
  IV U65384 ( .A(n45140), .Z(n47749) );
  IV U65385 ( .A(n45141), .Z(n45143) );
  IV U65386 ( .A(n45142), .Z(n47717) );
  NOR U65387 ( .A(n45143), .B(n47717), .Z(n53033) );
  IV U65388 ( .A(n53033), .Z(n47723) );
  IV U65389 ( .A(n45144), .Z(n50165) );
  NOR U65390 ( .A(n50165), .B(n45145), .Z(n47714) );
  IV U65391 ( .A(n45146), .Z(n45148) );
  NOR U65392 ( .A(n45148), .B(n45147), .Z(n50171) );
  IV U65393 ( .A(n45149), .Z(n45152) );
  IV U65394 ( .A(n45150), .Z(n47711) );
  XOR U65395 ( .A(n45153), .B(n47711), .Z(n45151) );
  NOR U65396 ( .A(n45152), .B(n45151), .Z(n50180) );
  IV U65397 ( .A(n45153), .Z(n45154) );
  NOR U65398 ( .A(n45154), .B(n47711), .Z(n47708) );
  IV U65399 ( .A(n47708), .Z(n47695) );
  IV U65400 ( .A(n47675), .Z(n45155) );
  NOR U65401 ( .A(n45155), .B(n47674), .Z(n47668) );
  IV U65402 ( .A(n47668), .Z(n47662) );
  IV U65403 ( .A(n45156), .Z(n45159) );
  IV U65404 ( .A(n45157), .Z(n45158) );
  NOR U65405 ( .A(n45159), .B(n45158), .Z(n50222) );
  IV U65406 ( .A(n45160), .Z(n50229) );
  IV U65407 ( .A(n45161), .Z(n45162) );
  NOR U65408 ( .A(n45165), .B(n45162), .Z(n50233) );
  IV U65409 ( .A(n45163), .Z(n45164) );
  NOR U65410 ( .A(n45165), .B(n45164), .Z(n50225) );
  NOR U65411 ( .A(n50233), .B(n50225), .Z(n47644) );
  IV U65412 ( .A(n45166), .Z(n45167) );
  NOR U65413 ( .A(n45167), .B(n47640), .Z(n50230) );
  IV U65414 ( .A(n45168), .Z(n45170) );
  IV U65415 ( .A(n45169), .Z(n47637) );
  NOR U65416 ( .A(n45170), .B(n47637), .Z(n58219) );
  NOR U65417 ( .A(n45171), .B(n47628), .Z(n47620) );
  IV U65418 ( .A(n45172), .Z(n47609) );
  IV U65419 ( .A(n45173), .Z(n45174) );
  NOR U65420 ( .A(n47609), .B(n45174), .Z(n50240) );
  IV U65421 ( .A(n45175), .Z(n45176) );
  NOR U65422 ( .A(n45176), .B(n47567), .Z(n58182) );
  IV U65423 ( .A(n45177), .Z(n52990) );
  NOR U65424 ( .A(n52990), .B(n45178), .Z(n50268) );
  IV U65425 ( .A(n45179), .Z(n45181) );
  NOR U65426 ( .A(n45181), .B(n45180), .Z(n50270) );
  NOR U65427 ( .A(n50268), .B(n50270), .Z(n47560) );
  IV U65428 ( .A(n45182), .Z(n45183) );
  NOR U65429 ( .A(n45183), .B(n45185), .Z(n50276) );
  IV U65430 ( .A(n45184), .Z(n45186) );
  NOR U65431 ( .A(n45186), .B(n45185), .Z(n50274) );
  NOR U65432 ( .A(n50276), .B(n50274), .Z(n47559) );
  NOR U65433 ( .A(n50280), .B(n45187), .Z(n45192) );
  IV U65434 ( .A(n45188), .Z(n45191) );
  IV U65435 ( .A(n45189), .Z(n45190) );
  NOR U65436 ( .A(n45191), .B(n45190), .Z(n50286) );
  NOR U65437 ( .A(n45192), .B(n50286), .Z(n47558) );
  IV U65438 ( .A(n45193), .Z(n45196) );
  IV U65439 ( .A(n45194), .Z(n45195) );
  NOR U65440 ( .A(n45196), .B(n45195), .Z(n52980) );
  IV U65441 ( .A(n45197), .Z(n45199) );
  IV U65442 ( .A(n45198), .Z(n45201) );
  NOR U65443 ( .A(n45199), .B(n45201), .Z(n50300) );
  IV U65444 ( .A(n45200), .Z(n45202) );
  NOR U65445 ( .A(n45202), .B(n45201), .Z(n50298) );
  IV U65446 ( .A(n45203), .Z(n45204) );
  NOR U65447 ( .A(n45207), .B(n45204), .Z(n50309) );
  IV U65448 ( .A(n45205), .Z(n45206) );
  NOR U65449 ( .A(n45207), .B(n45206), .Z(n50303) );
  XOR U65450 ( .A(n50309), .B(n50303), .Z(n45208) );
  NOR U65451 ( .A(n50298), .B(n45208), .Z(n47539) );
  IV U65452 ( .A(n45209), .Z(n45211) );
  NOR U65453 ( .A(n45211), .B(n45210), .Z(n50306) );
  IV U65454 ( .A(n45212), .Z(n45213) );
  NOR U65455 ( .A(n45216), .B(n45213), .Z(n50318) );
  IV U65456 ( .A(n45214), .Z(n45215) );
  NOR U65457 ( .A(n45216), .B(n45215), .Z(n50315) );
  IV U65458 ( .A(n45217), .Z(n45219) );
  NOR U65459 ( .A(n45219), .B(n45218), .Z(n50312) );
  IV U65460 ( .A(n45220), .Z(n45222) );
  NOR U65461 ( .A(n45222), .B(n45221), .Z(n47531) );
  IV U65462 ( .A(n47531), .Z(n47521) );
  NOR U65463 ( .A(n50339), .B(n45223), .Z(n50333) );
  IV U65464 ( .A(n45224), .Z(n45227) );
  IV U65465 ( .A(n45225), .Z(n45226) );
  NOR U65466 ( .A(n45227), .B(n45226), .Z(n45228) );
  IV U65467 ( .A(n45228), .Z(n50343) );
  IV U65468 ( .A(n45229), .Z(n45232) );
  IV U65469 ( .A(n45230), .Z(n45231) );
  NOR U65470 ( .A(n45232), .B(n45231), .Z(n52958) );
  IV U65471 ( .A(n45233), .Z(n45234) );
  NOR U65472 ( .A(n45234), .B(n47516), .Z(n45235) );
  IV U65473 ( .A(n45235), .Z(n50347) );
  IV U65474 ( .A(n45236), .Z(n50361) );
  NOR U65475 ( .A(n45237), .B(n50361), .Z(n45240) );
  NOR U65476 ( .A(n45238), .B(n50353), .Z(n45239) );
  NOR U65477 ( .A(n45240), .B(n45239), .Z(n47514) );
  NOR U65478 ( .A(n45241), .B(n50371), .Z(n45242) );
  IV U65479 ( .A(n45242), .Z(n50367) );
  IV U65480 ( .A(n45243), .Z(n50394) );
  NOR U65481 ( .A(n45244), .B(n50394), .Z(n47507) );
  IV U65482 ( .A(n45245), .Z(n45246) );
  NOR U65483 ( .A(n45250), .B(n45246), .Z(n45247) );
  IV U65484 ( .A(n45247), .Z(n52942) );
  IV U65485 ( .A(n45248), .Z(n45249) );
  NOR U65486 ( .A(n45250), .B(n45249), .Z(n47502) );
  IV U65487 ( .A(n45251), .Z(n45252) );
  NOR U65488 ( .A(n45252), .B(n45256), .Z(n50439) );
  IV U65489 ( .A(n45253), .Z(n50444) );
  NOR U65490 ( .A(n50444), .B(n45254), .Z(n50431) );
  IV U65491 ( .A(n45255), .Z(n45257) );
  NOR U65492 ( .A(n45257), .B(n45256), .Z(n52888) );
  NOR U65493 ( .A(n50431), .B(n52888), .Z(n47417) );
  NOR U65494 ( .A(n45259), .B(n45258), .Z(n45268) );
  IV U65495 ( .A(n45268), .Z(n45262) );
  IV U65496 ( .A(n45260), .Z(n45261) );
  NOR U65497 ( .A(n45262), .B(n45261), .Z(n50453) );
  IV U65498 ( .A(n45263), .Z(n45265) );
  NOR U65499 ( .A(n45265), .B(n45264), .Z(n45266) );
  IV U65500 ( .A(n45266), .Z(n45267) );
  NOR U65501 ( .A(n45268), .B(n45267), .Z(n52868) );
  NOR U65502 ( .A(n50453), .B(n52868), .Z(n47407) );
  IV U65503 ( .A(n45269), .Z(n45270) );
  NOR U65504 ( .A(n45270), .B(n47401), .Z(n52860) );
  NOR U65505 ( .A(n50473), .B(n50471), .Z(n45274) );
  IV U65506 ( .A(n45271), .Z(n47395) );
  IV U65507 ( .A(n45272), .Z(n45273) );
  NOR U65508 ( .A(n47395), .B(n45273), .Z(n50474) );
  NOR U65509 ( .A(n45274), .B(n50474), .Z(n47397) );
  IV U65510 ( .A(n45275), .Z(n45277) );
  NOR U65511 ( .A(n45277), .B(n45276), .Z(n50479) );
  IV U65512 ( .A(n45278), .Z(n45279) );
  NOR U65513 ( .A(n47392), .B(n45279), .Z(n50482) );
  IV U65514 ( .A(n45280), .Z(n45282) );
  NOR U65515 ( .A(n45282), .B(n45281), .Z(n47387) );
  IV U65516 ( .A(n47387), .Z(n47377) );
  IV U65517 ( .A(n45283), .Z(n45285) );
  IV U65518 ( .A(n45284), .Z(n45288) );
  NOR U65519 ( .A(n45285), .B(n45288), .Z(n50489) );
  NOR U65520 ( .A(n45286), .B(n50496), .Z(n45290) );
  IV U65521 ( .A(n45287), .Z(n45289) );
  NOR U65522 ( .A(n45289), .B(n45288), .Z(n50492) );
  NOR U65523 ( .A(n45290), .B(n50492), .Z(n47375) );
  IV U65524 ( .A(n45291), .Z(n50503) );
  NOR U65525 ( .A(n45292), .B(n50503), .Z(n47374) );
  NOR U65526 ( .A(n50511), .B(n45293), .Z(n45297) );
  IV U65527 ( .A(n45294), .Z(n45296) );
  IV U65528 ( .A(n45295), .Z(n45299) );
  NOR U65529 ( .A(n45296), .B(n45299), .Z(n50515) );
  NOR U65530 ( .A(n45297), .B(n50515), .Z(n47373) );
  IV U65531 ( .A(n45298), .Z(n45300) );
  NOR U65532 ( .A(n45300), .B(n45299), .Z(n47371) );
  IV U65533 ( .A(n47371), .Z(n47361) );
  IV U65534 ( .A(n45301), .Z(n45304) );
  IV U65535 ( .A(n45302), .Z(n45303) );
  NOR U65536 ( .A(n45304), .B(n45303), .Z(n52824) );
  IV U65537 ( .A(n45305), .Z(n45307) );
  XOR U65538 ( .A(n47356), .B(n47357), .Z(n45306) );
  NOR U65539 ( .A(n45307), .B(n45306), .Z(n45308) );
  IV U65540 ( .A(n45308), .Z(n52823) );
  IV U65541 ( .A(n45309), .Z(n45310) );
  NOR U65542 ( .A(n45310), .B(n47357), .Z(n50522) );
  IV U65543 ( .A(n45311), .Z(n50535) );
  NOR U65544 ( .A(n45312), .B(n50535), .Z(n50529) );
  NOR U65545 ( .A(n45313), .B(n52809), .Z(n45314) );
  NOR U65546 ( .A(n50529), .B(n45314), .Z(n47354) );
  IV U65547 ( .A(n45315), .Z(n45317) );
  NOR U65548 ( .A(n45317), .B(n45316), .Z(n50538) );
  IV U65549 ( .A(n45318), .Z(n45319) );
  NOR U65550 ( .A(n45322), .B(n45319), .Z(n50544) );
  IV U65551 ( .A(n45320), .Z(n45321) );
  NOR U65552 ( .A(n45322), .B(n45321), .Z(n50542) );
  NOR U65553 ( .A(n50544), .B(n50542), .Z(n47353) );
  NOR U65554 ( .A(n45323), .B(n50550), .Z(n45327) );
  IV U65555 ( .A(n45324), .Z(n45326) );
  IV U65556 ( .A(n45325), .Z(n47348) );
  NOR U65557 ( .A(n45326), .B(n47348), .Z(n52805) );
  NOR U65558 ( .A(n45327), .B(n52805), .Z(n47352) );
  IV U65559 ( .A(n45328), .Z(n45330) );
  XOR U65560 ( .A(n45333), .B(n45335), .Z(n45329) );
  NOR U65561 ( .A(n45330), .B(n45329), .Z(n50558) );
  IV U65562 ( .A(n45331), .Z(n45332) );
  NOR U65563 ( .A(n45335), .B(n45332), .Z(n50561) );
  IV U65564 ( .A(n45333), .Z(n45334) );
  NOR U65565 ( .A(n45335), .B(n45334), .Z(n52796) );
  NOR U65566 ( .A(n50561), .B(n52796), .Z(n47338) );
  IV U65567 ( .A(n45336), .Z(n45337) );
  NOR U65568 ( .A(n45337), .B(n47334), .Z(n50563) );
  IV U65569 ( .A(n45338), .Z(n50568) );
  NOR U65570 ( .A(n45339), .B(n50568), .Z(n47328) );
  IV U65571 ( .A(n45340), .Z(n45341) );
  NOR U65572 ( .A(n47321), .B(n45341), .Z(n52790) );
  IV U65573 ( .A(n45342), .Z(n45344) );
  IV U65574 ( .A(n45343), .Z(n47323) );
  NOR U65575 ( .A(n45344), .B(n47323), .Z(n47315) );
  IV U65576 ( .A(n45345), .Z(n45346) );
  NOR U65577 ( .A(n45349), .B(n45346), .Z(n52778) );
  IV U65578 ( .A(n45347), .Z(n45348) );
  NOR U65579 ( .A(n45349), .B(n45348), .Z(n47312) );
  IV U65580 ( .A(n47312), .Z(n47304) );
  IV U65581 ( .A(n45350), .Z(n57932) );
  NOR U65582 ( .A(n47297), .B(n57932), .Z(n47296) );
  IV U65583 ( .A(n47298), .Z(n45351) );
  NOR U65584 ( .A(n47297), .B(n45351), .Z(n45352) );
  IV U65585 ( .A(n45352), .Z(n52769) );
  IV U65586 ( .A(n45353), .Z(n45355) );
  IV U65587 ( .A(n45354), .Z(n45357) );
  NOR U65588 ( .A(n45355), .B(n45357), .Z(n52765) );
  IV U65589 ( .A(n45356), .Z(n45358) );
  NOR U65590 ( .A(n45358), .B(n45357), .Z(n45359) );
  IV U65591 ( .A(n45359), .Z(n50577) );
  NOR U65592 ( .A(n45360), .B(n52758), .Z(n45364) );
  IV U65593 ( .A(n45361), .Z(n45367) );
  IV U65594 ( .A(n45362), .Z(n45363) );
  NOR U65595 ( .A(n45367), .B(n45363), .Z(n52753) );
  NOR U65596 ( .A(n45364), .B(n52753), .Z(n47294) );
  IV U65597 ( .A(n45365), .Z(n45366) );
  NOR U65598 ( .A(n45367), .B(n45366), .Z(n45368) );
  IV U65599 ( .A(n45368), .Z(n52751) );
  IV U65600 ( .A(n45369), .Z(n45370) );
  NOR U65601 ( .A(n45373), .B(n45370), .Z(n52738) );
  IV U65602 ( .A(n45371), .Z(n45372) );
  NOR U65603 ( .A(n45373), .B(n45372), .Z(n45377) );
  IV U65604 ( .A(n52737), .Z(n45376) );
  IV U65605 ( .A(n45374), .Z(n45375) );
  NOR U65606 ( .A(n45376), .B(n45375), .Z(n50579) );
  NOR U65607 ( .A(n45377), .B(n50579), .Z(n52734) );
  IV U65608 ( .A(n45378), .Z(n45380) );
  XOR U65609 ( .A(n47266), .B(n47267), .Z(n45379) );
  NOR U65610 ( .A(n45380), .B(n45379), .Z(n50585) );
  IV U65611 ( .A(n45381), .Z(n45382) );
  NOR U65612 ( .A(n45382), .B(n47267), .Z(n50582) );
  IV U65613 ( .A(n45383), .Z(n45384) );
  NOR U65614 ( .A(n45388), .B(n45384), .Z(n45385) );
  IV U65615 ( .A(n45385), .Z(n52723) );
  IV U65616 ( .A(n45386), .Z(n45387) );
  NOR U65617 ( .A(n45388), .B(n45387), .Z(n50591) );
  IV U65618 ( .A(n45389), .Z(n45391) );
  NOR U65619 ( .A(n45391), .B(n45390), .Z(n50594) );
  NOR U65620 ( .A(n50591), .B(n50594), .Z(n47261) );
  IV U65621 ( .A(n45392), .Z(n45398) );
  IV U65622 ( .A(n45393), .Z(n45394) );
  NOR U65623 ( .A(n45398), .B(n45394), .Z(n45395) );
  IV U65624 ( .A(n45395), .Z(n50607) );
  IV U65625 ( .A(n45396), .Z(n45397) );
  NOR U65626 ( .A(n45398), .B(n45397), .Z(n50604) );
  IV U65627 ( .A(n45399), .Z(n45401) );
  NOR U65628 ( .A(n45401), .B(n45400), .Z(n50609) );
  IV U65629 ( .A(n45402), .Z(n45403) );
  IV U65630 ( .A(n45406), .Z(n45409) );
  NOR U65631 ( .A(n45403), .B(n45409), .Z(n50614) );
  IV U65632 ( .A(n45404), .Z(n45408) );
  IV U65633 ( .A(n45405), .Z(n45410) );
  XOR U65634 ( .A(n45410), .B(n45406), .Z(n45407) );
  NOR U65635 ( .A(n45408), .B(n45407), .Z(n50612) );
  NOR U65636 ( .A(n50614), .B(n50612), .Z(n47252) );
  NOR U65637 ( .A(n45410), .B(n45409), .Z(n52701) );
  IV U65638 ( .A(n45411), .Z(n45412) );
  NOR U65639 ( .A(n45412), .B(n45417), .Z(n45413) );
  IV U65640 ( .A(n45413), .Z(n52693) );
  IV U65641 ( .A(n45414), .Z(n50631) );
  NOR U65642 ( .A(n50631), .B(n45415), .Z(n45419) );
  IV U65643 ( .A(n45416), .Z(n45418) );
  NOR U65644 ( .A(n45418), .B(n45417), .Z(n50623) );
  NOR U65645 ( .A(n45419), .B(n50623), .Z(n47241) );
  IV U65646 ( .A(n45420), .Z(n45422) );
  NOR U65647 ( .A(n45422), .B(n45421), .Z(n50637) );
  NOR U65648 ( .A(n45423), .B(n50644), .Z(n47220) );
  IV U65649 ( .A(n45424), .Z(n45425) );
  NOR U65650 ( .A(n45425), .B(n45427), .Z(n52684) );
  IV U65651 ( .A(n45426), .Z(n45428) );
  NOR U65652 ( .A(n45428), .B(n45427), .Z(n52682) );
  NOR U65653 ( .A(n45429), .B(n63048), .Z(n52680) );
  NOR U65654 ( .A(n52682), .B(n52680), .Z(n45430) );
  IV U65655 ( .A(n45430), .Z(n45431) );
  NOR U65656 ( .A(n52684), .B(n45431), .Z(n47218) );
  IV U65657 ( .A(n45432), .Z(n45435) );
  IV U65658 ( .A(n45433), .Z(n45434) );
  NOR U65659 ( .A(n45435), .B(n45434), .Z(n50653) );
  IV U65660 ( .A(n45436), .Z(n45438) );
  XOR U65661 ( .A(n45444), .B(n45445), .Z(n45437) );
  NOR U65662 ( .A(n45438), .B(n45437), .Z(n50650) );
  IV U65663 ( .A(n45439), .Z(n47212) );
  IV U65664 ( .A(n45440), .Z(n45441) );
  NOR U65665 ( .A(n47212), .B(n45441), .Z(n50660) );
  IV U65666 ( .A(n45442), .Z(n45443) );
  NOR U65667 ( .A(n45443), .B(n45445), .Z(n50658) );
  IV U65668 ( .A(n45444), .Z(n45446) );
  NOR U65669 ( .A(n45446), .B(n45445), .Z(n50655) );
  NOR U65670 ( .A(n50658), .B(n50655), .Z(n45447) );
  IV U65671 ( .A(n45447), .Z(n45448) );
  NOR U65672 ( .A(n50660), .B(n45448), .Z(n47217) );
  IV U65673 ( .A(n45449), .Z(n45450) );
  NOR U65674 ( .A(n45450), .B(n45452), .Z(n50662) );
  IV U65675 ( .A(n45451), .Z(n45453) );
  NOR U65676 ( .A(n45453), .B(n45452), .Z(n50667) );
  IV U65677 ( .A(n45454), .Z(n45459) );
  IV U65678 ( .A(n45455), .Z(n45456) );
  NOR U65679 ( .A(n45459), .B(n45456), .Z(n52670) );
  IV U65680 ( .A(n45457), .Z(n45458) );
  NOR U65681 ( .A(n45459), .B(n45458), .Z(n52667) );
  IV U65682 ( .A(n45460), .Z(n45462) );
  NOR U65683 ( .A(n45462), .B(n45461), .Z(n50674) );
  IV U65684 ( .A(n45463), .Z(n55863) );
  NOR U65685 ( .A(n45464), .B(n55863), .Z(n50691) );
  IV U65686 ( .A(n45465), .Z(n45466) );
  NOR U65687 ( .A(n45466), .B(n47182), .Z(n50688) );
  NOR U65688 ( .A(n50691), .B(n50688), .Z(n47178) );
  IV U65689 ( .A(n45467), .Z(n45469) );
  NOR U65690 ( .A(n45469), .B(n45468), .Z(n47175) );
  IV U65691 ( .A(n47175), .Z(n47167) );
  IV U65692 ( .A(n45470), .Z(n45471) );
  NOR U65693 ( .A(n47171), .B(n45471), .Z(n50694) );
  IV U65694 ( .A(n45472), .Z(n45474) );
  NOR U65695 ( .A(n45474), .B(n45473), .Z(n45475) );
  IV U65696 ( .A(n45475), .Z(n50700) );
  IV U65697 ( .A(n45484), .Z(n45476) );
  NOR U65698 ( .A(n45483), .B(n45476), .Z(n45479) );
  IV U65699 ( .A(n45477), .Z(n45478) );
  NOR U65700 ( .A(n45479), .B(n45478), .Z(n50696) );
  IV U65701 ( .A(n45480), .Z(n50706) );
  IV U65702 ( .A(n45481), .Z(n45482) );
  NOR U65703 ( .A(n50706), .B(n45482), .Z(n61062) );
  IV U65704 ( .A(n45483), .Z(n45485) );
  NOR U65705 ( .A(n45485), .B(n45484), .Z(n61056) );
  NOR U65706 ( .A(n61062), .B(n61056), .Z(n50702) );
  IV U65707 ( .A(n45486), .Z(n45487) );
  NOR U65708 ( .A(n50706), .B(n45487), .Z(n45491) );
  IV U65709 ( .A(n45488), .Z(n45490) );
  NOR U65710 ( .A(n45490), .B(n45489), .Z(n50710) );
  NOR U65711 ( .A(n45491), .B(n50710), .Z(n50703) );
  IV U65712 ( .A(n45492), .Z(n45493) );
  NOR U65713 ( .A(n45496), .B(n45493), .Z(n50707) );
  IV U65714 ( .A(n45494), .Z(n45495) );
  NOR U65715 ( .A(n45496), .B(n45495), .Z(n50717) );
  IV U65716 ( .A(n45497), .Z(n45500) );
  IV U65717 ( .A(n45498), .Z(n45499) );
  NOR U65718 ( .A(n45500), .B(n45499), .Z(n50714) );
  IV U65719 ( .A(n45501), .Z(n45502) );
  NOR U65720 ( .A(n45502), .B(n45504), .Z(n50726) );
  IV U65721 ( .A(n45503), .Z(n45505) );
  NOR U65722 ( .A(n45505), .B(n45504), .Z(n50728) );
  XOR U65723 ( .A(n50726), .B(n50728), .Z(n45506) );
  NOR U65724 ( .A(n50720), .B(n45506), .Z(n47160) );
  IV U65725 ( .A(n45507), .Z(n45508) );
  NOR U65726 ( .A(n45509), .B(n45508), .Z(n45510) );
  IV U65727 ( .A(n45510), .Z(n45512) );
  NOR U65728 ( .A(n45512), .B(n45511), .Z(n52624) );
  IV U65729 ( .A(n45513), .Z(n45514) );
  NOR U65730 ( .A(n45514), .B(n47157), .Z(n52618) );
  IV U65731 ( .A(n45515), .Z(n45516) );
  NOR U65732 ( .A(n45516), .B(n47153), .Z(n52608) );
  IV U65733 ( .A(n45517), .Z(n45522) );
  IV U65734 ( .A(n45518), .Z(n45519) );
  NOR U65735 ( .A(n45522), .B(n45519), .Z(n52595) );
  IV U65736 ( .A(n45520), .Z(n45521) );
  NOR U65737 ( .A(n45522), .B(n45521), .Z(n50736) );
  IV U65738 ( .A(n45523), .Z(n45525) );
  NOR U65739 ( .A(n45525), .B(n45524), .Z(n50738) );
  NOR U65740 ( .A(n50736), .B(n50738), .Z(n45526) );
  IV U65741 ( .A(n45526), .Z(n47143) );
  IV U65742 ( .A(n45527), .Z(n45528) );
  NOR U65743 ( .A(n45531), .B(n45528), .Z(n50740) );
  IV U65744 ( .A(n45529), .Z(n45530) );
  NOR U65745 ( .A(n45531), .B(n45530), .Z(n50744) );
  IV U65746 ( .A(n45532), .Z(n45533) );
  NOR U65747 ( .A(n45533), .B(n45537), .Z(n50747) );
  NOR U65748 ( .A(n50744), .B(n50747), .Z(n47142) );
  IV U65749 ( .A(n45534), .Z(n50753) );
  NOR U65750 ( .A(n45535), .B(n50753), .Z(n45539) );
  IV U65751 ( .A(n45536), .Z(n45538) );
  NOR U65752 ( .A(n45538), .B(n45537), .Z(n50749) );
  NOR U65753 ( .A(n45539), .B(n50749), .Z(n47141) );
  NOR U65754 ( .A(n45541), .B(n45540), .Z(n50759) );
  NOR U65755 ( .A(n45543), .B(n45542), .Z(n45546) );
  NOR U65756 ( .A(n50784), .B(n50782), .Z(n50779) );
  NOR U65757 ( .A(n45544), .B(n50779), .Z(n45545) );
  NOR U65758 ( .A(n45546), .B(n45545), .Z(n50774) );
  NOR U65759 ( .A(n45547), .B(n50787), .Z(n45554) );
  IV U65760 ( .A(n45548), .Z(n45549) );
  NOR U65761 ( .A(n45552), .B(n45549), .Z(n50796) );
  IV U65762 ( .A(n45550), .Z(n45551) );
  NOR U65763 ( .A(n45552), .B(n45551), .Z(n50780) );
  XOR U65764 ( .A(n50796), .B(n50780), .Z(n45553) );
  NOR U65765 ( .A(n45554), .B(n45553), .Z(n47133) );
  IV U65766 ( .A(n47126), .Z(n45555) );
  NOR U65767 ( .A(n47125), .B(n45555), .Z(n52584) );
  IV U65768 ( .A(n45556), .Z(n52572) );
  IV U65769 ( .A(n45557), .Z(n45558) );
  NOR U65770 ( .A(n45558), .B(n45560), .Z(n50803) );
  IV U65771 ( .A(n45559), .Z(n45561) );
  NOR U65772 ( .A(n45561), .B(n45560), .Z(n52565) );
  NOR U65773 ( .A(n50803), .B(n52565), .Z(n47104) );
  IV U65774 ( .A(n45562), .Z(n45567) );
  IV U65775 ( .A(n45563), .Z(n45564) );
  NOR U65776 ( .A(n45567), .B(n45564), .Z(n50801) );
  IV U65777 ( .A(n45565), .Z(n45566) );
  NOR U65778 ( .A(n45567), .B(n45566), .Z(n50807) );
  IV U65779 ( .A(n45568), .Z(n45570) );
  NOR U65780 ( .A(n45570), .B(n45569), .Z(n50809) );
  NOR U65781 ( .A(n50807), .B(n50809), .Z(n47103) );
  IV U65782 ( .A(n45571), .Z(n45572) );
  NOR U65783 ( .A(n45572), .B(n45574), .Z(n50812) );
  IV U65784 ( .A(n45573), .Z(n45575) );
  NOR U65785 ( .A(n45575), .B(n45574), .Z(n50814) );
  IV U65786 ( .A(n45576), .Z(n45577) );
  NOR U65787 ( .A(n45577), .B(n45581), .Z(n52559) );
  NOR U65788 ( .A(n50814), .B(n52559), .Z(n45578) );
  IV U65789 ( .A(n45578), .Z(n45579) );
  NOR U65790 ( .A(n50812), .B(n45579), .Z(n47102) );
  IV U65791 ( .A(n45580), .Z(n45582) );
  NOR U65792 ( .A(n45582), .B(n45581), .Z(n52556) );
  IV U65793 ( .A(n45583), .Z(n45584) );
  NOR U65794 ( .A(n45587), .B(n45584), .Z(n50831) );
  IV U65795 ( .A(n45585), .Z(n45586) );
  NOR U65796 ( .A(n45587), .B(n45586), .Z(n50829) );
  NOR U65797 ( .A(n50831), .B(n50829), .Z(n47095) );
  IV U65798 ( .A(n45588), .Z(n45590) );
  NOR U65799 ( .A(n45590), .B(n45589), .Z(n50826) );
  NOR U65800 ( .A(n45592), .B(n45591), .Z(n47084) );
  IV U65801 ( .A(n47084), .Z(n47076) );
  IV U65802 ( .A(n45593), .Z(n45599) );
  IV U65803 ( .A(n45594), .Z(n45595) );
  NOR U65804 ( .A(n45599), .B(n45595), .Z(n45596) );
  IV U65805 ( .A(n45596), .Z(n52530) );
  IV U65806 ( .A(n45597), .Z(n45598) );
  NOR U65807 ( .A(n45599), .B(n45598), .Z(n50855) );
  IV U65808 ( .A(n45600), .Z(n45602) );
  NOR U65809 ( .A(n45602), .B(n45601), .Z(n52520) );
  IV U65810 ( .A(n45603), .Z(n45605) );
  NOR U65811 ( .A(n45605), .B(n45604), .Z(n47050) );
  IV U65812 ( .A(n47050), .Z(n47039) );
  IV U65813 ( .A(n45606), .Z(n45607) );
  NOR U65814 ( .A(n45607), .B(n45609), .Z(n50872) );
  IV U65815 ( .A(n45608), .Z(n45610) );
  NOR U65816 ( .A(n45610), .B(n45609), .Z(n52508) );
  NOR U65817 ( .A(n50872), .B(n52508), .Z(n45611) );
  IV U65818 ( .A(n45611), .Z(n47042) );
  IV U65819 ( .A(n45612), .Z(n50876) );
  NOR U65820 ( .A(n45613), .B(n50876), .Z(n45614) );
  NOR U65821 ( .A(n50879), .B(n45614), .Z(n47037) );
  IV U65822 ( .A(n45615), .Z(n45616) );
  NOR U65823 ( .A(n45616), .B(n45618), .Z(n62853) );
  IV U65824 ( .A(n45617), .Z(n45619) );
  NOR U65825 ( .A(n45619), .B(n45618), .Z(n62861) );
  NOR U65826 ( .A(n62853), .B(n62861), .Z(n50884) );
  IV U65827 ( .A(n50884), .Z(n45624) );
  IV U65828 ( .A(n45620), .Z(n47033) );
  NOR U65829 ( .A(n45621), .B(n47033), .Z(n45622) );
  IV U65830 ( .A(n45622), .Z(n45623) );
  NOR U65831 ( .A(n47032), .B(n45623), .Z(n50880) );
  NOR U65832 ( .A(n45624), .B(n50880), .Z(n47036) );
  IV U65833 ( .A(n45625), .Z(n45626) );
  NOR U65834 ( .A(n45626), .B(n45631), .Z(n50900) );
  IV U65835 ( .A(n45627), .Z(n45629) );
  XOR U65836 ( .A(n45630), .B(n45631), .Z(n45628) );
  NOR U65837 ( .A(n45629), .B(n45628), .Z(n50896) );
  NOR U65838 ( .A(n50900), .B(n50896), .Z(n47020) );
  IV U65839 ( .A(n45630), .Z(n45632) );
  NOR U65840 ( .A(n45632), .B(n45631), .Z(n45633) );
  IV U65841 ( .A(n45633), .Z(n50899) );
  IV U65842 ( .A(n45634), .Z(n45636) );
  IV U65843 ( .A(n45635), .Z(n47016) );
  NOR U65844 ( .A(n45636), .B(n47016), .Z(n50903) );
  IV U65845 ( .A(n45637), .Z(n45638) );
  NOR U65846 ( .A(n45638), .B(n45641), .Z(n50918) );
  IV U65847 ( .A(n45639), .Z(n50925) );
  NOR U65848 ( .A(n50925), .B(n50927), .Z(n45643) );
  IV U65849 ( .A(n45640), .Z(n45642) );
  NOR U65850 ( .A(n45642), .B(n45641), .Z(n50921) );
  NOR U65851 ( .A(n45643), .B(n50921), .Z(n47005) );
  IV U65852 ( .A(n45644), .Z(n45646) );
  NOR U65853 ( .A(n45646), .B(n45645), .Z(n50928) );
  IV U65854 ( .A(n45647), .Z(n45650) );
  NOR U65855 ( .A(n45648), .B(n45650), .Z(n52483) );
  IV U65856 ( .A(n45649), .Z(n45651) );
  NOR U65857 ( .A(n45651), .B(n45650), .Z(n50931) );
  XOR U65858 ( .A(n52483), .B(n50931), .Z(n45652) );
  NOR U65859 ( .A(n50928), .B(n45652), .Z(n47004) );
  NOR U65860 ( .A(n45653), .B(n56101), .Z(n52481) );
  IV U65861 ( .A(n45654), .Z(n45656) );
  IV U65862 ( .A(n45655), .Z(n45658) );
  NOR U65863 ( .A(n45656), .B(n45658), .Z(n52473) );
  IV U65864 ( .A(n45657), .Z(n45659) );
  NOR U65865 ( .A(n45659), .B(n45658), .Z(n52472) );
  XOR U65866 ( .A(n52473), .B(n52472), .Z(n45660) );
  NOR U65867 ( .A(n52481), .B(n45660), .Z(n47003) );
  IV U65868 ( .A(n45661), .Z(n45662) );
  NOR U65869 ( .A(n46992), .B(n45662), .Z(n47001) );
  IV U65870 ( .A(n47001), .Z(n46989) );
  NOR U65871 ( .A(n45664), .B(n45663), .Z(n50937) );
  IV U65872 ( .A(n45665), .Z(n45667) );
  IV U65873 ( .A(n45666), .Z(n46995) );
  NOR U65874 ( .A(n45667), .B(n46995), .Z(n50935) );
  NOR U65875 ( .A(n50937), .B(n50935), .Z(n46997) );
  IV U65876 ( .A(n45668), .Z(n57651) );
  IV U65877 ( .A(n57650), .Z(n45670) );
  NOR U65878 ( .A(n57651), .B(n45670), .Z(n50941) );
  IV U65879 ( .A(n45669), .Z(n45671) );
  NOR U65880 ( .A(n45671), .B(n45670), .Z(n50939) );
  NOR U65881 ( .A(n50941), .B(n50939), .Z(n46987) );
  NOR U65882 ( .A(n56123), .B(n45672), .Z(n50946) );
  IV U65883 ( .A(n45673), .Z(n45676) );
  IV U65884 ( .A(n45674), .Z(n45675) );
  NOR U65885 ( .A(n45676), .B(n45675), .Z(n50943) );
  IV U65886 ( .A(n45677), .Z(n45680) );
  IV U65887 ( .A(n45678), .Z(n45679) );
  NOR U65888 ( .A(n45680), .B(n45679), .Z(n52458) );
  NOR U65889 ( .A(n52454), .B(n52458), .Z(n46985) );
  IV U65890 ( .A(n45681), .Z(n45682) );
  NOR U65891 ( .A(n45682), .B(n45684), .Z(n52447) );
  IV U65892 ( .A(n45683), .Z(n45685) );
  NOR U65893 ( .A(n45685), .B(n45684), .Z(n52450) );
  NOR U65894 ( .A(n52447), .B(n52450), .Z(n46984) );
  IV U65895 ( .A(n45686), .Z(n45687) );
  NOR U65896 ( .A(n45687), .B(n46977), .Z(n50951) );
  IV U65897 ( .A(n45688), .Z(n46981) );
  IV U65898 ( .A(n45689), .Z(n45690) );
  NOR U65899 ( .A(n46981), .B(n45690), .Z(n50954) );
  IV U65900 ( .A(n45691), .Z(n45693) );
  NOR U65901 ( .A(n45693), .B(n45692), .Z(n50962) );
  IV U65902 ( .A(n45694), .Z(n45699) );
  IV U65903 ( .A(n45695), .Z(n45696) );
  NOR U65904 ( .A(n45699), .B(n45696), .Z(n45697) );
  IV U65905 ( .A(n45697), .Z(n57615) );
  NOR U65906 ( .A(n45699), .B(n45698), .Z(n50966) );
  IV U65907 ( .A(n45700), .Z(n45702) );
  NOR U65908 ( .A(n45702), .B(n45701), .Z(n52442) );
  NOR U65909 ( .A(n50966), .B(n52442), .Z(n46975) );
  IV U65910 ( .A(n45703), .Z(n45704) );
  NOR U65911 ( .A(n45704), .B(n46968), .Z(n50974) );
  IV U65912 ( .A(n45705), .Z(n45707) );
  IV U65913 ( .A(n45706), .Z(n46961) );
  NOR U65914 ( .A(n45707), .B(n46961), .Z(n50971) );
  IV U65915 ( .A(n45708), .Z(n45710) );
  IV U65916 ( .A(n45709), .Z(n46951) );
  NOR U65917 ( .A(n45710), .B(n46951), .Z(n46948) );
  IV U65918 ( .A(n46948), .Z(n46943) );
  IV U65919 ( .A(n45711), .Z(n46937) );
  IV U65920 ( .A(n45712), .Z(n45713) );
  NOR U65921 ( .A(n46937), .B(n45713), .Z(n51001) );
  IV U65922 ( .A(n45714), .Z(n45716) );
  IV U65923 ( .A(n45715), .Z(n46931) );
  NOR U65924 ( .A(n45716), .B(n46931), .Z(n52421) );
  IV U65925 ( .A(n45717), .Z(n45719) );
  NOR U65926 ( .A(n45719), .B(n45718), .Z(n52404) );
  IV U65927 ( .A(n45720), .Z(n45722) );
  IV U65928 ( .A(n45721), .Z(n45725) );
  NOR U65929 ( .A(n45722), .B(n45725), .Z(n45723) );
  IV U65930 ( .A(n45723), .Z(n52398) );
  NOR U65931 ( .A(n45724), .B(n56193), .Z(n52394) );
  NOR U65932 ( .A(n45726), .B(n45725), .Z(n52400) );
  NOR U65933 ( .A(n52394), .B(n52400), .Z(n46920) );
  IV U65934 ( .A(n45727), .Z(n45729) );
  NOR U65935 ( .A(n45729), .B(n45728), .Z(n52393) );
  IV U65936 ( .A(n45730), .Z(n45735) );
  IV U65937 ( .A(n45731), .Z(n45732) );
  NOR U65938 ( .A(n45735), .B(n45732), .Z(n51026) );
  IV U65939 ( .A(n45733), .Z(n45734) );
  NOR U65940 ( .A(n45735), .B(n45734), .Z(n51023) );
  IV U65941 ( .A(n45736), .Z(n45738) );
  NOR U65942 ( .A(n45738), .B(n45737), .Z(n51033) );
  NOR U65943 ( .A(n51023), .B(n51033), .Z(n46912) );
  IV U65944 ( .A(n45739), .Z(n46909) );
  NOR U65945 ( .A(n45740), .B(n46909), .Z(n46907) );
  IV U65946 ( .A(n46907), .Z(n46900) );
  IV U65947 ( .A(n45741), .Z(n45742) );
  NOR U65948 ( .A(n46874), .B(n45742), .Z(n46885) );
  IV U65949 ( .A(n46885), .Z(n46871) );
  IV U65950 ( .A(n45743), .Z(n52378) );
  NOR U65951 ( .A(n52378), .B(n45744), .Z(n45747) );
  IV U65952 ( .A(n45745), .Z(n45746) );
  NOR U65953 ( .A(n45746), .B(n46878), .Z(n51041) );
  NOR U65954 ( .A(n45747), .B(n51041), .Z(n46870) );
  IV U65955 ( .A(n45748), .Z(n45749) );
  NOR U65956 ( .A(n45749), .B(n45754), .Z(n57542) );
  IV U65957 ( .A(n45750), .Z(n46852) );
  IV U65958 ( .A(n45751), .Z(n45752) );
  NOR U65959 ( .A(n46852), .B(n45752), .Z(n57533) );
  NOR U65960 ( .A(n57542), .B(n57533), .Z(n51044) );
  IV U65961 ( .A(n51044), .Z(n45756) );
  IV U65962 ( .A(n45753), .Z(n45755) );
  NOR U65963 ( .A(n45755), .B(n45754), .Z(n52373) );
  NOR U65964 ( .A(n45756), .B(n52373), .Z(n46869) );
  IV U65965 ( .A(n45757), .Z(n45758) );
  NOR U65966 ( .A(n45758), .B(n46862), .Z(n46860) );
  IV U65967 ( .A(n51062), .Z(n45759) );
  NOR U65968 ( .A(n45759), .B(n45765), .Z(n51065) );
  IV U65969 ( .A(n45760), .Z(n45762) );
  XOR U65970 ( .A(n45764), .B(n45765), .Z(n45761) );
  NOR U65971 ( .A(n45762), .B(n45761), .Z(n45763) );
  NOR U65972 ( .A(n51065), .B(n45763), .Z(n51059) );
  IV U65973 ( .A(n45764), .Z(n45766) );
  NOR U65974 ( .A(n45766), .B(n45765), .Z(n51063) );
  IV U65975 ( .A(n45767), .Z(n45768) );
  NOR U65976 ( .A(n45775), .B(n45768), .Z(n51098) );
  IV U65977 ( .A(n45769), .Z(n45772) );
  IV U65978 ( .A(n45770), .Z(n45771) );
  NOR U65979 ( .A(n45772), .B(n45771), .Z(n51103) );
  NOR U65980 ( .A(n51098), .B(n51103), .Z(n46789) );
  IV U65981 ( .A(n45773), .Z(n45774) );
  NOR U65982 ( .A(n45775), .B(n45774), .Z(n45776) );
  IV U65983 ( .A(n45776), .Z(n51097) );
  IV U65984 ( .A(n45777), .Z(n45779) );
  XOR U65985 ( .A(n45785), .B(n45786), .Z(n45778) );
  NOR U65986 ( .A(n45779), .B(n45778), .Z(n51100) );
  IV U65987 ( .A(n45780), .Z(n45793) );
  IV U65988 ( .A(n45781), .Z(n45782) );
  NOR U65989 ( .A(n45793), .B(n45782), .Z(n52319) );
  IV U65990 ( .A(n45783), .Z(n45784) );
  NOR U65991 ( .A(n45784), .B(n45786), .Z(n51106) );
  IV U65992 ( .A(n45785), .Z(n45787) );
  NOR U65993 ( .A(n45787), .B(n45786), .Z(n52322) );
  NOR U65994 ( .A(n51106), .B(n52322), .Z(n45788) );
  IV U65995 ( .A(n45788), .Z(n45789) );
  NOR U65996 ( .A(n52319), .B(n45789), .Z(n46786) );
  IV U65997 ( .A(n52318), .Z(n45790) );
  NOR U65998 ( .A(n45790), .B(n45799), .Z(n51109) );
  IV U65999 ( .A(n45791), .Z(n45792) );
  NOR U66000 ( .A(n45793), .B(n45792), .Z(n45794) );
  NOR U66001 ( .A(n51109), .B(n45794), .Z(n52314) );
  IV U66002 ( .A(n45795), .Z(n45803) );
  IV U66003 ( .A(n45796), .Z(n45797) );
  NOR U66004 ( .A(n45803), .B(n45797), .Z(n52302) );
  IV U66005 ( .A(n45798), .Z(n45800) );
  NOR U66006 ( .A(n45800), .B(n45799), .Z(n51112) );
  NOR U66007 ( .A(n52302), .B(n51112), .Z(n46785) );
  IV U66008 ( .A(n45801), .Z(n45802) );
  NOR U66009 ( .A(n45803), .B(n45802), .Z(n52306) );
  IV U66010 ( .A(n45804), .Z(n45806) );
  IV U66011 ( .A(n45805), .Z(n45809) );
  NOR U66012 ( .A(n45806), .B(n45809), .Z(n51117) );
  NOR U66013 ( .A(n45807), .B(n52288), .Z(n45811) );
  IV U66014 ( .A(n45808), .Z(n45810) );
  NOR U66015 ( .A(n45810), .B(n45809), .Z(n51121) );
  NOR U66016 ( .A(n45811), .B(n51121), .Z(n46770) );
  IV U66017 ( .A(n45812), .Z(n45814) );
  IV U66018 ( .A(n45813), .Z(n46760) );
  NOR U66019 ( .A(n45814), .B(n46760), .Z(n45815) );
  IV U66020 ( .A(n45815), .Z(n52285) );
  IV U66021 ( .A(n57431), .Z(n45816) );
  NOR U66022 ( .A(n57429), .B(n45816), .Z(n57433) );
  IV U66023 ( .A(n52271), .Z(n45817) );
  NOR U66024 ( .A(n52270), .B(n45817), .Z(n46744) );
  IV U66025 ( .A(n45818), .Z(n45820) );
  IV U66026 ( .A(n45819), .Z(n46737) );
  NOR U66027 ( .A(n45820), .B(n46737), .Z(n45821) );
  IV U66028 ( .A(n45821), .Z(n52260) );
  IV U66029 ( .A(n51155), .Z(n45823) );
  IV U66030 ( .A(n45822), .Z(n45828) );
  NOR U66031 ( .A(n45823), .B(n45828), .Z(n52256) );
  IV U66032 ( .A(n45824), .Z(n45825) );
  NOR U66033 ( .A(n46735), .B(n45825), .Z(n45826) );
  NOR U66034 ( .A(n52256), .B(n45826), .Z(n51152) );
  IV U66035 ( .A(n45827), .Z(n45829) );
  NOR U66036 ( .A(n45829), .B(n45828), .Z(n52251) );
  NOR U66037 ( .A(n56361), .B(n45830), .Z(n45831) );
  IV U66038 ( .A(n45831), .Z(n46722) );
  NOR U66039 ( .A(n45833), .B(n45832), .Z(n45837) );
  IV U66040 ( .A(n45834), .Z(n45836) );
  IV U66041 ( .A(n45835), .Z(n46718) );
  NOR U66042 ( .A(n45836), .B(n46718), .Z(n52236) );
  NOR U66043 ( .A(n45837), .B(n52236), .Z(n46714) );
  NOR U66044 ( .A(n51170), .B(n45838), .Z(n51160) );
  IV U66045 ( .A(n45839), .Z(n45841) );
  IV U66046 ( .A(n45840), .Z(n46712) );
  NOR U66047 ( .A(n45841), .B(n46712), .Z(n51176) );
  IV U66048 ( .A(n45842), .Z(n45843) );
  NOR U66049 ( .A(n45846), .B(n45843), .Z(n51179) );
  NOR U66050 ( .A(n51176), .B(n51179), .Z(n46710) );
  IV U66051 ( .A(n45844), .Z(n45845) );
  NOR U66052 ( .A(n45846), .B(n45845), .Z(n46706) );
  IV U66053 ( .A(n45847), .Z(n45849) );
  IV U66054 ( .A(n45848), .Z(n46702) );
  NOR U66055 ( .A(n45849), .B(n46702), .Z(n51187) );
  IV U66056 ( .A(n45850), .Z(n45852) );
  NOR U66057 ( .A(n45852), .B(n45851), .Z(n51184) );
  XOR U66058 ( .A(n51190), .B(n51184), .Z(n45853) );
  NOR U66059 ( .A(n51187), .B(n45853), .Z(n46700) );
  IV U66060 ( .A(n45854), .Z(n45855) );
  NOR U66061 ( .A(n45855), .B(n45860), .Z(n45856) );
  IV U66062 ( .A(n45856), .Z(n52225) );
  IV U66063 ( .A(n45857), .Z(n52213) );
  NOR U66064 ( .A(n45858), .B(n52213), .Z(n45862) );
  IV U66065 ( .A(n45859), .Z(n45861) );
  NOR U66066 ( .A(n45861), .B(n45860), .Z(n52217) );
  NOR U66067 ( .A(n45862), .B(n52217), .Z(n46692) );
  IV U66068 ( .A(n45863), .Z(n51204) );
  NOR U66069 ( .A(n45864), .B(n51204), .Z(n45866) );
  NOR U66070 ( .A(n52206), .B(n52204), .Z(n45865) );
  NOR U66071 ( .A(n45866), .B(n45865), .Z(n46685) );
  IV U66072 ( .A(n45867), .Z(n45868) );
  NOR U66073 ( .A(n45868), .B(n45872), .Z(n51214) );
  IV U66074 ( .A(n45869), .Z(n56430) );
  NOR U66075 ( .A(n45870), .B(n56430), .Z(n51217) );
  IV U66076 ( .A(n45871), .Z(n45873) );
  NOR U66077 ( .A(n45873), .B(n45872), .Z(n51211) );
  NOR U66078 ( .A(n51217), .B(n51211), .Z(n45874) );
  IV U66079 ( .A(n45874), .Z(n45875) );
  NOR U66080 ( .A(n51214), .B(n45875), .Z(n46684) );
  IV U66081 ( .A(n45876), .Z(n45877) );
  NOR U66082 ( .A(n45877), .B(n46677), .Z(n52194) );
  IV U66083 ( .A(n45878), .Z(n51234) );
  NOR U66084 ( .A(n45879), .B(n51234), .Z(n45880) );
  NOR U66085 ( .A(n52185), .B(n45880), .Z(n46675) );
  IV U66086 ( .A(n45881), .Z(n45884) );
  IV U66087 ( .A(n45882), .Z(n45883) );
  NOR U66088 ( .A(n45884), .B(n45883), .Z(n51242) );
  IV U66089 ( .A(n45885), .Z(n45886) );
  NOR U66090 ( .A(n45889), .B(n45886), .Z(n51238) );
  IV U66091 ( .A(n45887), .Z(n45888) );
  NOR U66092 ( .A(n45889), .B(n45888), .Z(n51240) );
  NOR U66093 ( .A(n51238), .B(n51240), .Z(n45890) );
  IV U66094 ( .A(n45890), .Z(n45891) );
  NOR U66095 ( .A(n51242), .B(n45891), .Z(n46674) );
  IV U66096 ( .A(n45892), .Z(n45894) );
  XOR U66097 ( .A(n45897), .B(n45899), .Z(n45893) );
  NOR U66098 ( .A(n45894), .B(n45893), .Z(n51248) );
  IV U66099 ( .A(n45895), .Z(n45896) );
  NOR U66100 ( .A(n45899), .B(n45896), .Z(n51245) );
  IV U66101 ( .A(n45897), .Z(n45898) );
  NOR U66102 ( .A(n45899), .B(n45898), .Z(n52168) );
  NOR U66103 ( .A(n45901), .B(n45900), .Z(n45904) );
  NOR U66104 ( .A(n45902), .B(n52164), .Z(n45903) );
  NOR U66105 ( .A(n45904), .B(n45903), .Z(n46673) );
  IV U66106 ( .A(n45905), .Z(n45906) );
  NOR U66107 ( .A(n46671), .B(n45906), .Z(n45909) );
  IV U66108 ( .A(n52154), .Z(n45908) );
  NOR U66109 ( .A(n45908), .B(n45907), .Z(n51257) );
  NOR U66110 ( .A(n45909), .B(n51257), .Z(n52151) );
  IV U66111 ( .A(n45910), .Z(n45911) );
  NOR U66112 ( .A(n45911), .B(n45913), .Z(n52142) );
  IV U66113 ( .A(n45912), .Z(n45914) );
  NOR U66114 ( .A(n45914), .B(n45913), .Z(n52139) );
  NOR U66115 ( .A(n45915), .B(n51262), .Z(n46662) );
  IV U66116 ( .A(n45916), .Z(n56490) );
  NOR U66117 ( .A(n45917), .B(n56490), .Z(n46659) );
  IV U66118 ( .A(n46659), .Z(n46651) );
  IV U66119 ( .A(n45918), .Z(n51285) );
  NOR U66120 ( .A(n45919), .B(n51285), .Z(n51276) );
  IV U66121 ( .A(n45920), .Z(n45922) );
  NOR U66122 ( .A(n45922), .B(n45921), .Z(n51281) );
  NOR U66123 ( .A(n51276), .B(n51281), .Z(n46650) );
  IV U66124 ( .A(n45923), .Z(n45927) );
  IV U66125 ( .A(n45924), .Z(n45925) );
  NOR U66126 ( .A(n45927), .B(n45925), .Z(n52133) );
  NOR U66127 ( .A(n45927), .B(n45926), .Z(n52130) );
  IV U66128 ( .A(n45928), .Z(n45930) );
  NOR U66129 ( .A(n45930), .B(n45929), .Z(n51292) );
  IV U66130 ( .A(n45931), .Z(n45932) );
  NOR U66131 ( .A(n45932), .B(n46635), .Z(n51289) );
  IV U66132 ( .A(n45933), .Z(n45934) );
  NOR U66133 ( .A(n56540), .B(n45934), .Z(n51305) );
  NOR U66134 ( .A(n45935), .B(n51332), .Z(n51322) );
  IV U66135 ( .A(n45936), .Z(n45938) );
  NOR U66136 ( .A(n45938), .B(n45937), .Z(n51335) );
  IV U66137 ( .A(n45939), .Z(n45941) );
  IV U66138 ( .A(n45940), .Z(n45943) );
  NOR U66139 ( .A(n45941), .B(n45943), .Z(n51342) );
  NOR U66140 ( .A(n62313), .B(n45942), .Z(n52106) );
  NOR U66141 ( .A(n45944), .B(n45943), .Z(n51345) );
  NOR U66142 ( .A(n52106), .B(n51345), .Z(n45945) );
  IV U66143 ( .A(n45945), .Z(n46593) );
  IV U66144 ( .A(n45946), .Z(n45948) );
  IV U66145 ( .A(n45947), .Z(n46575) );
  NOR U66146 ( .A(n45948), .B(n46575), .Z(n45949) );
  IV U66147 ( .A(n45949), .Z(n56588) );
  IV U66148 ( .A(n45950), .Z(n56596) );
  NOR U66149 ( .A(n45951), .B(n56596), .Z(n45952) );
  IV U66150 ( .A(n45952), .Z(n52099) );
  NOR U66151 ( .A(n45953), .B(n52085), .Z(n46573) );
  IV U66152 ( .A(n45954), .Z(n45956) );
  IV U66153 ( .A(n45955), .Z(n45958) );
  NOR U66154 ( .A(n45956), .B(n45958), .Z(n52088) );
  IV U66155 ( .A(n45957), .Z(n45959) );
  NOR U66156 ( .A(n45959), .B(n45958), .Z(n52091) );
  NOR U66157 ( .A(n45960), .B(n52091), .Z(n46572) );
  NOR U66158 ( .A(n51350), .B(n51352), .Z(n46571) );
  IV U66159 ( .A(n45961), .Z(n45962) );
  NOR U66160 ( .A(n45966), .B(n45962), .Z(n45963) );
  IV U66161 ( .A(n45963), .Z(n51358) );
  IV U66162 ( .A(n45964), .Z(n45965) );
  NOR U66163 ( .A(n45966), .B(n45965), .Z(n56628) );
  IV U66164 ( .A(n45967), .Z(n45970) );
  IV U66165 ( .A(n45968), .Z(n45969) );
  NOR U66166 ( .A(n45970), .B(n45969), .Z(n56633) );
  NOR U66167 ( .A(n56628), .B(n56633), .Z(n52073) );
  IV U66168 ( .A(n45971), .Z(n45974) );
  IV U66169 ( .A(n45972), .Z(n45973) );
  NOR U66170 ( .A(n45974), .B(n45973), .Z(n52058) );
  NOR U66171 ( .A(n56636), .B(n52058), .Z(n46570) );
  IV U66172 ( .A(n45975), .Z(n45976) );
  NOR U66173 ( .A(n45976), .B(n45978), .Z(n46568) );
  IV U66174 ( .A(n45977), .Z(n45979) );
  NOR U66175 ( .A(n45979), .B(n45978), .Z(n51361) );
  IV U66176 ( .A(n45980), .Z(n45981) );
  IV U66177 ( .A(n45984), .Z(n45988) );
  NOR U66178 ( .A(n45981), .B(n45988), .Z(n51375) );
  IV U66179 ( .A(n45982), .Z(n45986) );
  IV U66180 ( .A(n45983), .Z(n45989) );
  XOR U66181 ( .A(n45989), .B(n45984), .Z(n45985) );
  NOR U66182 ( .A(n45986), .B(n45985), .Z(n51372) );
  NOR U66183 ( .A(n51375), .B(n51372), .Z(n46559) );
  NOR U66184 ( .A(n51381), .B(n45987), .Z(n45990) );
  NOR U66185 ( .A(n45989), .B(n45988), .Z(n51377) );
  NOR U66186 ( .A(n45990), .B(n51377), .Z(n46558) );
  IV U66187 ( .A(n45991), .Z(n45994) );
  IV U66188 ( .A(n45992), .Z(n45993) );
  NOR U66189 ( .A(n45994), .B(n45993), .Z(n52047) );
  IV U66190 ( .A(n45995), .Z(n45997) );
  NOR U66191 ( .A(n45997), .B(n45996), .Z(n52044) );
  IV U66192 ( .A(n45998), .Z(n45999) );
  NOR U66193 ( .A(n46005), .B(n45999), .Z(n52041) );
  IV U66194 ( .A(n46000), .Z(n46002) );
  NOR U66195 ( .A(n46002), .B(n46001), .Z(n51388) );
  NOR U66196 ( .A(n52041), .B(n51388), .Z(n46557) );
  IV U66197 ( .A(n46003), .Z(n46004) );
  NOR U66198 ( .A(n46005), .B(n46004), .Z(n46006) );
  IV U66199 ( .A(n46006), .Z(n51387) );
  IV U66200 ( .A(n46009), .Z(n46007) );
  NOR U66201 ( .A(n46008), .B(n46007), .Z(n46013) );
  IV U66202 ( .A(n46008), .Z(n56667) );
  NOR U66203 ( .A(n46009), .B(n56667), .Z(n51401) );
  NOR U66204 ( .A(n51395), .B(n51401), .Z(n46010) );
  IV U66205 ( .A(n46010), .Z(n51394) );
  NOR U66206 ( .A(n51394), .B(n46011), .Z(n46012) );
  NOR U66207 ( .A(n46013), .B(n46012), .Z(n51390) );
  IV U66208 ( .A(n46014), .Z(n46015) );
  NOR U66209 ( .A(n46015), .B(n46553), .Z(n51403) );
  IV U66210 ( .A(n46016), .Z(n46018) );
  NOR U66211 ( .A(n46018), .B(n46017), .Z(n52003) );
  IV U66212 ( .A(n46541), .Z(n46535) );
  IV U66213 ( .A(n46019), .Z(n46020) );
  NOR U66214 ( .A(n46020), .B(n46528), .Z(n46532) );
  IV U66215 ( .A(n46532), .Z(n46525) );
  IV U66216 ( .A(n46021), .Z(n51423) );
  NOR U66217 ( .A(n51423), .B(n46022), .Z(n51421) );
  NOR U66218 ( .A(n46024), .B(n46023), .Z(n51414) );
  NOR U66219 ( .A(n51421), .B(n51414), .Z(n46523) );
  IV U66220 ( .A(n46025), .Z(n46027) );
  NOR U66221 ( .A(n46027), .B(n46026), .Z(n51429) );
  IV U66222 ( .A(n46028), .Z(n46029) );
  NOR U66223 ( .A(n46521), .B(n46029), .Z(n46517) );
  IV U66224 ( .A(n46517), .Z(n46507) );
  IV U66225 ( .A(n46030), .Z(n46032) );
  XOR U66226 ( .A(n46036), .B(n46037), .Z(n46031) );
  NOR U66227 ( .A(n46032), .B(n46031), .Z(n46033) );
  IV U66228 ( .A(n46033), .Z(n51436) );
  IV U66229 ( .A(n46034), .Z(n46035) );
  NOR U66230 ( .A(n46035), .B(n46037), .Z(n51433) );
  IV U66231 ( .A(n46036), .Z(n46038) );
  NOR U66232 ( .A(n46038), .B(n46037), .Z(n51440) );
  IV U66233 ( .A(n46039), .Z(n46505) );
  IV U66234 ( .A(n46040), .Z(n46041) );
  NOR U66235 ( .A(n46505), .B(n46041), .Z(n46500) );
  IV U66236 ( .A(n46042), .Z(n46052) );
  IV U66237 ( .A(n46043), .Z(n46044) );
  NOR U66238 ( .A(n46052), .B(n46044), .Z(n56745) );
  IV U66239 ( .A(n46045), .Z(n46046) );
  NOR U66240 ( .A(n46046), .B(n46048), .Z(n57146) );
  NOR U66241 ( .A(n56745), .B(n57146), .Z(n46470) );
  IV U66242 ( .A(n46047), .Z(n46049) );
  NOR U66243 ( .A(n46049), .B(n46048), .Z(n57151) );
  IV U66244 ( .A(n46050), .Z(n46051) );
  NOR U66245 ( .A(n46052), .B(n46051), .Z(n56750) );
  IV U66246 ( .A(n46053), .Z(n46054) );
  NOR U66247 ( .A(n46054), .B(n46056), .Z(n51963) );
  IV U66248 ( .A(n46055), .Z(n46057) );
  NOR U66249 ( .A(n46057), .B(n46056), .Z(n51961) );
  XOR U66250 ( .A(n51963), .B(n51961), .Z(n46058) );
  NOR U66251 ( .A(n56750), .B(n46058), .Z(n46468) );
  IV U66252 ( .A(n46059), .Z(n46461) );
  NOR U66253 ( .A(n46461), .B(n46060), .Z(n46451) );
  IV U66254 ( .A(n46061), .Z(n46063) );
  NOR U66255 ( .A(n46063), .B(n46062), .Z(n46449) );
  IV U66256 ( .A(n46449), .Z(n46444) );
  IV U66257 ( .A(n46064), .Z(n46065) );
  NOR U66258 ( .A(n46447), .B(n46065), .Z(n51476) );
  IV U66259 ( .A(n46066), .Z(n46067) );
  NOR U66260 ( .A(n46067), .B(n46072), .Z(n51481) );
  IV U66261 ( .A(n46068), .Z(n46069) );
  NOR U66262 ( .A(n46070), .B(n46069), .Z(n46074) );
  IV U66263 ( .A(n46071), .Z(n46073) );
  NOR U66264 ( .A(n46073), .B(n46072), .Z(n51952) );
  NOR U66265 ( .A(n46074), .B(n51952), .Z(n46441) );
  NOR U66266 ( .A(n46075), .B(n51501), .Z(n46428) );
  IV U66267 ( .A(n46076), .Z(n46077) );
  NOR U66268 ( .A(n46077), .B(n46079), .Z(n51904) );
  IV U66269 ( .A(n46078), .Z(n46080) );
  NOR U66270 ( .A(n46080), .B(n46079), .Z(n51516) );
  NOR U66271 ( .A(n51904), .B(n51516), .Z(n46400) );
  IV U66272 ( .A(n46081), .Z(n46383) );
  IV U66273 ( .A(n46082), .Z(n46083) );
  NOR U66274 ( .A(n46383), .B(n46083), .Z(n46084) );
  IV U66275 ( .A(n46084), .Z(n46395) );
  IV U66276 ( .A(n46085), .Z(n51884) );
  NOR U66277 ( .A(n46086), .B(n51884), .Z(n51889) );
  IV U66278 ( .A(n46087), .Z(n46088) );
  NOR U66279 ( .A(n46088), .B(n46090), .Z(n51521) );
  IV U66280 ( .A(n46089), .Z(n46091) );
  NOR U66281 ( .A(n46091), .B(n46090), .Z(n46092) );
  IV U66282 ( .A(n46092), .Z(n51526) );
  IV U66283 ( .A(n46093), .Z(n46094) );
  NOR U66284 ( .A(n46370), .B(n46094), .Z(n46095) );
  IV U66285 ( .A(n46095), .Z(n51542) );
  IV U66286 ( .A(n46371), .Z(n46096) );
  NOR U66287 ( .A(n46370), .B(n46096), .Z(n46365) );
  IV U66288 ( .A(n46097), .Z(n46099) );
  IV U66289 ( .A(n46098), .Z(n46362) );
  NOR U66290 ( .A(n46099), .B(n46362), .Z(n46359) );
  IV U66291 ( .A(n46359), .Z(n46352) );
  NOR U66292 ( .A(n51826), .B(n46100), .Z(n51831) );
  IV U66293 ( .A(n46101), .Z(n46103) );
  XOR U66294 ( .A(n46106), .B(n46108), .Z(n46102) );
  NOR U66295 ( .A(n46103), .B(n46102), .Z(n51561) );
  IV U66296 ( .A(n46104), .Z(n46105) );
  NOR U66297 ( .A(n46108), .B(n46105), .Z(n51564) );
  IV U66298 ( .A(n46106), .Z(n46107) );
  NOR U66299 ( .A(n46108), .B(n46107), .Z(n51566) );
  XOR U66300 ( .A(n51564), .B(n51566), .Z(n46109) );
  NOR U66301 ( .A(n51561), .B(n46109), .Z(n46319) );
  IV U66302 ( .A(n46110), .Z(n46112) );
  NOR U66303 ( .A(n46112), .B(n46111), .Z(n51569) );
  IV U66304 ( .A(n46113), .Z(n46114) );
  NOR U66305 ( .A(n46114), .B(n46315), .Z(n46115) );
  IV U66306 ( .A(n46115), .Z(n51817) );
  NOR U66307 ( .A(n51590), .B(n46116), .Z(n51580) );
  IV U66308 ( .A(n46117), .Z(n46118) );
  NOR U66309 ( .A(n46118), .B(n46296), .Z(n51809) );
  NOR U66310 ( .A(n51580), .B(n51809), .Z(n46311) );
  IV U66311 ( .A(n46119), .Z(n46120) );
  NOR U66312 ( .A(n46120), .B(n46122), .Z(n51599) );
  IV U66313 ( .A(n46121), .Z(n46123) );
  NOR U66314 ( .A(n46123), .B(n46122), .Z(n46124) );
  IV U66315 ( .A(n46124), .Z(n51803) );
  IV U66316 ( .A(n46125), .Z(n46128) );
  IV U66317 ( .A(n46126), .Z(n46127) );
  NOR U66318 ( .A(n46128), .B(n46127), .Z(n51776) );
  IV U66319 ( .A(n46129), .Z(n46130) );
  NOR U66320 ( .A(n46133), .B(n46130), .Z(n51768) );
  IV U66321 ( .A(n46131), .Z(n46132) );
  NOR U66322 ( .A(n46133), .B(n46132), .Z(n51757) );
  IV U66323 ( .A(n51755), .Z(n46134) );
  NOR U66324 ( .A(n51749), .B(n46134), .Z(n46137) );
  NOR U66325 ( .A(n46135), .B(n51619), .Z(n46136) );
  NOR U66326 ( .A(n46137), .B(n46136), .Z(n46260) );
  NOR U66327 ( .A(n46138), .B(n51624), .Z(n46146) );
  IV U66328 ( .A(n46139), .Z(n46144) );
  IV U66329 ( .A(n46140), .Z(n46141) );
  NOR U66330 ( .A(n46144), .B(n46141), .Z(n51631) );
  IV U66331 ( .A(n46142), .Z(n46143) );
  NOR U66332 ( .A(n46144), .B(n46143), .Z(n51751) );
  XOR U66333 ( .A(n51631), .B(n51751), .Z(n46145) );
  NOR U66334 ( .A(n46146), .B(n46145), .Z(n46147) );
  IV U66335 ( .A(n46147), .Z(n46259) );
  IV U66336 ( .A(n46148), .Z(n46149) );
  NOR U66337 ( .A(n46149), .B(n46244), .Z(n46236) );
  IV U66338 ( .A(n46236), .Z(n46230) );
  IV U66339 ( .A(n46150), .Z(n46151) );
  NOR U66340 ( .A(n46151), .B(n46227), .Z(n51720) );
  IV U66341 ( .A(n46152), .Z(n46153) );
  NOR U66342 ( .A(n51719), .B(n46153), .Z(n46158) );
  IV U66343 ( .A(n46154), .Z(n46157) );
  IV U66344 ( .A(n46155), .Z(n46156) );
  NOR U66345 ( .A(n46157), .B(n46156), .Z(n51703) );
  NOR U66346 ( .A(n46158), .B(n51703), .Z(n51716) );
  IV U66347 ( .A(n46159), .Z(n46162) );
  IV U66348 ( .A(n46160), .Z(n46161) );
  NOR U66349 ( .A(n46162), .B(n46161), .Z(n51708) );
  IV U66350 ( .A(n46163), .Z(n51706) );
  IV U66351 ( .A(n46164), .Z(n46165) );
  NOR U66352 ( .A(n46165), .B(n46166), .Z(n51666) );
  NOR U66353 ( .A(n46167), .B(n46166), .Z(n51663) );
  IV U66354 ( .A(n46168), .Z(n51675) );
  NOR U66355 ( .A(n46169), .B(n51675), .Z(n46170) );
  NOR U66356 ( .A(n51670), .B(n46170), .Z(n46222) );
  IV U66357 ( .A(n46171), .Z(n46172) );
  NOR U66358 ( .A(n46172), .B(n46208), .Z(n46220) );
  IV U66359 ( .A(n46220), .Z(n46206) );
  IV U66360 ( .A(n46173), .Z(n46174) );
  NOR U66361 ( .A(n46174), .B(n46201), .Z(n46194) );
  NOR U66362 ( .A(n46178), .B(n46175), .Z(n46176) );
  NOR U66363 ( .A(n46177), .B(n46176), .Z(n46182) );
  IV U66364 ( .A(n46178), .Z(n46180) );
  NOR U66365 ( .A(n46180), .B(n46179), .Z(n46181) );
  NOR U66366 ( .A(n46182), .B(n46181), .Z(n46183) );
  IV U66367 ( .A(n46183), .Z(n51691) );
  IV U66368 ( .A(n46184), .Z(n46186) );
  NOR U66369 ( .A(n46186), .B(n46185), .Z(n46190) );
  XOR U66370 ( .A(n51691), .B(n46190), .Z(n46192) );
  NOR U66371 ( .A(n46188), .B(n46187), .Z(n51692) );
  IV U66372 ( .A(n51692), .Z(n46189) );
  NOR U66373 ( .A(n46190), .B(n46189), .Z(n46191) );
  NOR U66374 ( .A(n46192), .B(n46191), .Z(n46193) );
  XOR U66375 ( .A(n46194), .B(n46193), .Z(n46203) );
  IV U66376 ( .A(n46195), .Z(n46214) );
  IV U66377 ( .A(n46196), .Z(n46197) );
  NOR U66378 ( .A(n46214), .B(n46197), .Z(n46204) );
  IV U66379 ( .A(n46204), .Z(n46198) );
  NOR U66380 ( .A(n46203), .B(n46198), .Z(n51696) );
  IV U66381 ( .A(n46199), .Z(n46200) );
  NOR U66382 ( .A(n46201), .B(n46200), .Z(n46202) );
  XOR U66383 ( .A(n46203), .B(n46202), .Z(n46210) );
  IV U66384 ( .A(n46210), .Z(n51693) );
  NOR U66385 ( .A(n51693), .B(n46204), .Z(n46205) );
  NOR U66386 ( .A(n51696), .B(n46205), .Z(n46215) );
  IV U66387 ( .A(n46215), .Z(n51687) );
  NOR U66388 ( .A(n46206), .B(n51687), .Z(n56963) );
  IV U66389 ( .A(n46207), .Z(n46209) );
  NOR U66390 ( .A(n46209), .B(n46208), .Z(n46217) );
  IV U66391 ( .A(n46217), .Z(n46211) );
  NOR U66392 ( .A(n46211), .B(n46210), .Z(n51688) );
  IV U66393 ( .A(n46212), .Z(n46213) );
  NOR U66394 ( .A(n46214), .B(n46213), .Z(n51685) );
  XOR U66395 ( .A(n46215), .B(n51685), .Z(n46216) );
  NOR U66396 ( .A(n46217), .B(n46216), .Z(n46218) );
  NOR U66397 ( .A(n51688), .B(n46218), .Z(n46219) );
  NOR U66398 ( .A(n46220), .B(n46219), .Z(n46221) );
  NOR U66399 ( .A(n56963), .B(n46221), .Z(n51671) );
  XOR U66400 ( .A(n46222), .B(n51671), .Z(n51665) );
  XOR U66401 ( .A(n51663), .B(n51665), .Z(n51667) );
  XOR U66402 ( .A(n51666), .B(n51667), .Z(n51658) );
  XOR U66403 ( .A(n51657), .B(n51658), .Z(n51661) );
  NOR U66404 ( .A(n51660), .B(n51655), .Z(n46223) );
  XOR U66405 ( .A(n51661), .B(n46223), .Z(n51705) );
  XOR U66406 ( .A(n51706), .B(n51705), .Z(n51710) );
  XOR U66407 ( .A(n51708), .B(n51710), .Z(n51715) );
  XOR U66408 ( .A(n51716), .B(n51715), .Z(n51649) );
  IV U66409 ( .A(n46224), .Z(n46225) );
  NOR U66410 ( .A(n51719), .B(n46225), .Z(n51651) );
  IV U66411 ( .A(n46226), .Z(n46228) );
  NOR U66412 ( .A(n46228), .B(n46227), .Z(n51648) );
  NOR U66413 ( .A(n51651), .B(n51648), .Z(n46229) );
  XOR U66414 ( .A(n51649), .B(n46229), .Z(n51722) );
  XOR U66415 ( .A(n51720), .B(n51722), .Z(n51724) );
  XOR U66416 ( .A(n51723), .B(n51724), .Z(n51646) );
  XOR U66417 ( .A(n51645), .B(n51646), .Z(n51643) );
  XOR U66418 ( .A(n51642), .B(n51643), .Z(n51729) );
  XOR U66419 ( .A(n51728), .B(n51729), .Z(n51732) );
  XOR U66420 ( .A(n51731), .B(n51732), .Z(n51737) );
  NOR U66421 ( .A(n46230), .B(n51737), .Z(n56900) );
  IV U66422 ( .A(n46231), .Z(n46232) );
  NOR U66423 ( .A(n46233), .B(n46232), .Z(n51638) );
  NOR U66424 ( .A(n51731), .B(n51638), .Z(n46234) );
  XOR U66425 ( .A(n51732), .B(n46234), .Z(n46235) );
  NOR U66426 ( .A(n46236), .B(n46235), .Z(n46237) );
  NOR U66427 ( .A(n56900), .B(n46237), .Z(n46246) );
  IV U66428 ( .A(n46246), .Z(n46242) );
  IV U66429 ( .A(n46238), .Z(n46240) );
  IV U66430 ( .A(n46239), .Z(n46250) );
  NOR U66431 ( .A(n46240), .B(n46250), .Z(n46253) );
  IV U66432 ( .A(n46253), .Z(n46241) );
  NOR U66433 ( .A(n46242), .B(n46241), .Z(n56897) );
  IV U66434 ( .A(n46243), .Z(n46245) );
  NOR U66435 ( .A(n46245), .B(n46244), .Z(n46247) );
  NOR U66436 ( .A(n46247), .B(n46246), .Z(n46249) );
  IV U66437 ( .A(n46247), .Z(n46248) );
  NOR U66438 ( .A(n46248), .B(n51737), .Z(n61947) );
  NOR U66439 ( .A(n46249), .B(n61947), .Z(n51635) );
  NOR U66440 ( .A(n46251), .B(n46250), .Z(n51634) );
  XOR U66441 ( .A(n51635), .B(n51634), .Z(n46252) );
  NOR U66442 ( .A(n46253), .B(n46252), .Z(n46254) );
  NOR U66443 ( .A(n56897), .B(n46254), .Z(n46255) );
  IV U66444 ( .A(n46255), .Z(n51745) );
  IV U66445 ( .A(n46256), .Z(n46258) );
  NOR U66446 ( .A(n46258), .B(n46257), .Z(n51743) );
  XOR U66447 ( .A(n51745), .B(n51743), .Z(n51632) );
  XOR U66448 ( .A(n46259), .B(n51632), .Z(n51620) );
  XOR U66449 ( .A(n46260), .B(n51620), .Z(n51759) );
  XOR U66450 ( .A(n51757), .B(n51759), .Z(n51769) );
  XOR U66451 ( .A(n51768), .B(n51769), .Z(n51772) );
  XOR U66452 ( .A(n51771), .B(n51772), .Z(n51777) );
  XOR U66453 ( .A(n51776), .B(n51777), .Z(n51785) );
  IV U66454 ( .A(n46261), .Z(n51615) );
  NOR U66455 ( .A(n46262), .B(n51615), .Z(n46265) );
  IV U66456 ( .A(n46263), .Z(n46264) );
  NOR U66457 ( .A(n46264), .B(n46270), .Z(n51612) );
  NOR U66458 ( .A(n46265), .B(n51612), .Z(n46266) );
  XOR U66459 ( .A(n51785), .B(n46266), .Z(n51788) );
  IV U66460 ( .A(n46267), .Z(n51790) );
  NOR U66461 ( .A(n51790), .B(n46268), .Z(n46272) );
  IV U66462 ( .A(n46269), .Z(n46271) );
  NOR U66463 ( .A(n46271), .B(n46270), .Z(n51784) );
  NOR U66464 ( .A(n46272), .B(n51784), .Z(n46273) );
  XOR U66465 ( .A(n51788), .B(n46273), .Z(n51801) );
  IV U66466 ( .A(n46274), .Z(n46275) );
  NOR U66467 ( .A(n46275), .B(n46277), .Z(n51793) );
  IV U66468 ( .A(n46276), .Z(n46278) );
  NOR U66469 ( .A(n46278), .B(n46277), .Z(n51800) );
  NOR U66470 ( .A(n51793), .B(n51800), .Z(n46279) );
  XOR U66471 ( .A(n51801), .B(n46279), .Z(n51604) );
  IV U66472 ( .A(n46280), .Z(n46292) );
  IV U66473 ( .A(n46281), .Z(n46282) );
  NOR U66474 ( .A(n46292), .B(n46282), .Z(n51605) );
  IV U66475 ( .A(n46283), .Z(n46285) );
  NOR U66476 ( .A(n46285), .B(n46284), .Z(n51609) );
  NOR U66477 ( .A(n51605), .B(n51609), .Z(n46286) );
  XOR U66478 ( .A(n51604), .B(n46286), .Z(n51806) );
  IV U66479 ( .A(n46287), .Z(n46289) );
  NOR U66480 ( .A(n46289), .B(n46288), .Z(n51805) );
  IV U66481 ( .A(n46290), .Z(n46291) );
  NOR U66482 ( .A(n46292), .B(n46291), .Z(n51607) );
  NOR U66483 ( .A(n51805), .B(n51607), .Z(n46293) );
  XOR U66484 ( .A(n51806), .B(n46293), .Z(n46294) );
  IV U66485 ( .A(n46294), .Z(n51804) );
  XOR U66486 ( .A(n51803), .B(n51804), .Z(n46302) );
  IV U66487 ( .A(n46302), .Z(n51603) );
  XOR U66488 ( .A(n51599), .B(n51603), .Z(n57027) );
  IV U66489 ( .A(n46295), .Z(n46297) );
  NOR U66490 ( .A(n46297), .B(n46296), .Z(n46309) );
  IV U66491 ( .A(n46309), .Z(n46298) );
  NOR U66492 ( .A(n57027), .B(n46298), .Z(n57022) );
  IV U66493 ( .A(n46299), .Z(n46306) );
  IV U66494 ( .A(n46300), .Z(n46301) );
  NOR U66495 ( .A(n46306), .B(n46301), .Z(n51601) );
  NOR U66496 ( .A(n51599), .B(n51601), .Z(n46303) );
  XOR U66497 ( .A(n46303), .B(n46302), .Z(n51598) );
  IV U66498 ( .A(n46304), .Z(n46305) );
  NOR U66499 ( .A(n46306), .B(n46305), .Z(n46307) );
  IV U66500 ( .A(n46307), .Z(n51597) );
  XOR U66501 ( .A(n51598), .B(n51597), .Z(n46308) );
  NOR U66502 ( .A(n46309), .B(n46308), .Z(n46310) );
  NOR U66503 ( .A(n57022), .B(n46310), .Z(n51578) );
  XOR U66504 ( .A(n46311), .B(n51578), .Z(n51574) );
  NOR U66505 ( .A(n46313), .B(n46312), .Z(n46317) );
  IV U66506 ( .A(n46314), .Z(n46316) );
  NOR U66507 ( .A(n46316), .B(n46315), .Z(n51572) );
  NOR U66508 ( .A(n46317), .B(n51572), .Z(n46318) );
  XOR U66509 ( .A(n51574), .B(n46318), .Z(n51815) );
  XOR U66510 ( .A(n51817), .B(n51815), .Z(n51571) );
  XOR U66511 ( .A(n51569), .B(n51571), .Z(n51565) );
  XOR U66512 ( .A(n46319), .B(n51565), .Z(n46320) );
  IV U66513 ( .A(n46320), .Z(n51825) );
  IV U66514 ( .A(n46321), .Z(n46324) );
  IV U66515 ( .A(n46322), .Z(n46323) );
  NOR U66516 ( .A(n46324), .B(n46323), .Z(n51823) );
  XOR U66517 ( .A(n51825), .B(n51823), .Z(n51838) );
  XOR U66518 ( .A(n51831), .B(n51838), .Z(n51556) );
  IV U66519 ( .A(n46328), .Z(n51839) );
  NOR U66520 ( .A(n46326), .B(n51839), .Z(n46331) );
  IV U66521 ( .A(n46325), .Z(n51560) );
  IV U66522 ( .A(n46326), .Z(n46327) );
  NOR U66523 ( .A(n46328), .B(n46327), .Z(n46329) );
  NOR U66524 ( .A(n51560), .B(n46329), .Z(n46330) );
  NOR U66525 ( .A(n46331), .B(n46330), .Z(n46332) );
  XOR U66526 ( .A(n51556), .B(n46332), .Z(n51553) );
  IV U66527 ( .A(n46333), .Z(n46338) );
  IV U66528 ( .A(n46334), .Z(n46335) );
  NOR U66529 ( .A(n46338), .B(n46335), .Z(n51554) );
  IV U66530 ( .A(n46336), .Z(n46337) );
  NOR U66531 ( .A(n46338), .B(n46337), .Z(n51852) );
  IV U66532 ( .A(n46339), .Z(n46340) );
  NOR U66533 ( .A(n46340), .B(n51557), .Z(n51853) );
  XOR U66534 ( .A(n51852), .B(n51853), .Z(n46341) );
  NOR U66535 ( .A(n51554), .B(n46341), .Z(n46342) );
  XOR U66536 ( .A(n51553), .B(n46342), .Z(n51859) );
  NOR U66537 ( .A(n51863), .B(n51861), .Z(n46346) );
  IV U66538 ( .A(n46343), .Z(n46345) );
  IV U66539 ( .A(n46344), .Z(n46349) );
  NOR U66540 ( .A(n46345), .B(n46349), .Z(n51857) );
  NOR U66541 ( .A(n46346), .B(n51857), .Z(n46347) );
  XOR U66542 ( .A(n51859), .B(n46347), .Z(n51550) );
  IV U66543 ( .A(n46348), .Z(n46350) );
  NOR U66544 ( .A(n46350), .B(n46349), .Z(n46351) );
  IV U66545 ( .A(n46351), .Z(n51551) );
  XOR U66546 ( .A(n51550), .B(n51551), .Z(n51871) );
  NOR U66547 ( .A(n46352), .B(n51871), .Z(n61786) );
  IV U66548 ( .A(n46353), .Z(n46354) );
  NOR U66549 ( .A(n46357), .B(n46354), .Z(n51547) );
  IV U66550 ( .A(n46355), .Z(n46356) );
  NOR U66551 ( .A(n46357), .B(n46356), .Z(n51870) );
  XOR U66552 ( .A(n51870), .B(n51871), .Z(n51548) );
  XOR U66553 ( .A(n51547), .B(n51548), .Z(n46366) );
  IV U66554 ( .A(n46366), .Z(n46358) );
  NOR U66555 ( .A(n46359), .B(n46358), .Z(n46360) );
  NOR U66556 ( .A(n61786), .B(n46360), .Z(n51543) );
  IV U66557 ( .A(n46361), .Z(n46363) );
  NOR U66558 ( .A(n46363), .B(n46362), .Z(n51544) );
  XOR U66559 ( .A(n51543), .B(n51544), .Z(n46364) );
  NOR U66560 ( .A(n46365), .B(n46364), .Z(n46368) );
  IV U66561 ( .A(n46365), .Z(n46367) );
  NOR U66562 ( .A(n46367), .B(n46366), .Z(n57079) );
  NOR U66563 ( .A(n46368), .B(n57079), .Z(n51538) );
  XOR U66564 ( .A(n51542), .B(n51538), .Z(n51537) );
  IV U66565 ( .A(n46369), .Z(n46373) );
  XOR U66566 ( .A(n46371), .B(n46370), .Z(n46372) );
  NOR U66567 ( .A(n46373), .B(n46372), .Z(n51535) );
  XOR U66568 ( .A(n51537), .B(n51535), .Z(n51528) );
  NOR U66569 ( .A(n51529), .B(n46374), .Z(n46379) );
  IV U66570 ( .A(n46375), .Z(n46378) );
  IV U66571 ( .A(n46376), .Z(n46377) );
  NOR U66572 ( .A(n46378), .B(n46377), .Z(n51539) );
  NOR U66573 ( .A(n46379), .B(n51539), .Z(n46380) );
  XOR U66574 ( .A(n51528), .B(n46380), .Z(n51525) );
  XOR U66575 ( .A(n51526), .B(n51525), .Z(n51522) );
  XOR U66576 ( .A(n51521), .B(n51522), .Z(n51896) );
  XOR U66577 ( .A(n51889), .B(n51896), .Z(n46392) );
  NOR U66578 ( .A(n46395), .B(n46392), .Z(n57086) );
  IV U66579 ( .A(n46381), .Z(n46382) );
  NOR U66580 ( .A(n46383), .B(n46382), .Z(n51901) );
  IV U66581 ( .A(n46384), .Z(n46386) );
  NOR U66582 ( .A(n46386), .B(n46385), .Z(n51897) );
  IV U66583 ( .A(n46387), .Z(n46388) );
  NOR U66584 ( .A(n46388), .B(n46390), .Z(n51519) );
  IV U66585 ( .A(n46389), .Z(n46391) );
  NOR U66586 ( .A(n46391), .B(n46390), .Z(n51894) );
  NOR U66587 ( .A(n51519), .B(n51894), .Z(n46393) );
  XOR U66588 ( .A(n46393), .B(n46392), .Z(n46394) );
  IV U66589 ( .A(n46394), .Z(n51899) );
  XOR U66590 ( .A(n51897), .B(n51899), .Z(n51902) );
  IV U66591 ( .A(n51902), .Z(n46396) );
  XOR U66592 ( .A(n51901), .B(n46396), .Z(n46398) );
  NOR U66593 ( .A(n46396), .B(n46395), .Z(n46397) );
  NOR U66594 ( .A(n46398), .B(n46397), .Z(n46399) );
  NOR U66595 ( .A(n57086), .B(n46399), .Z(n51517) );
  XOR U66596 ( .A(n46400), .B(n51517), .Z(n51909) );
  XOR U66597 ( .A(n51908), .B(n51909), .Z(n51913) );
  IV U66598 ( .A(n46401), .Z(n46404) );
  IV U66599 ( .A(n46402), .Z(n46403) );
  NOR U66600 ( .A(n46404), .B(n46403), .Z(n51911) );
  XOR U66601 ( .A(n51913), .B(n51911), .Z(n51922) );
  IV U66602 ( .A(n46405), .Z(n46408) );
  IV U66603 ( .A(n46406), .Z(n46407) );
  NOR U66604 ( .A(n46408), .B(n46407), .Z(n46409) );
  IV U66605 ( .A(n46409), .Z(n51515) );
  XOR U66606 ( .A(n51922), .B(n51515), .Z(n46416) );
  IV U66607 ( .A(n46410), .Z(n46411) );
  NOR U66608 ( .A(n46414), .B(n46411), .Z(n51513) );
  IV U66609 ( .A(n46412), .Z(n46413) );
  NOR U66610 ( .A(n46414), .B(n46413), .Z(n51920) );
  NOR U66611 ( .A(n51513), .B(n51920), .Z(n46415) );
  XOR U66612 ( .A(n46416), .B(n46415), .Z(n51919) );
  IV U66613 ( .A(n46417), .Z(n46426) );
  IV U66614 ( .A(n46418), .Z(n46419) );
  NOR U66615 ( .A(n46426), .B(n46419), .Z(n51917) );
  IV U66616 ( .A(n46420), .Z(n46422) );
  NOR U66617 ( .A(n46422), .B(n46421), .Z(n51511) );
  NOR U66618 ( .A(n51917), .B(n51511), .Z(n46423) );
  XOR U66619 ( .A(n51919), .B(n46423), .Z(n51505) );
  IV U66620 ( .A(n46424), .Z(n46425) );
  NOR U66621 ( .A(n46426), .B(n46425), .Z(n46427) );
  IV U66622 ( .A(n46427), .Z(n51506) );
  XOR U66623 ( .A(n51505), .B(n51506), .Z(n51500) );
  XOR U66624 ( .A(n46428), .B(n51500), .Z(n51490) );
  IV U66625 ( .A(n46429), .Z(n51493) );
  NOR U66626 ( .A(n46430), .B(n51493), .Z(n46438) );
  IV U66627 ( .A(n46431), .Z(n46432) );
  NOR U66628 ( .A(n46432), .B(n46434), .Z(n51489) );
  IV U66629 ( .A(n46433), .Z(n46435) );
  NOR U66630 ( .A(n46435), .B(n46434), .Z(n51487) );
  NOR U66631 ( .A(n51489), .B(n51487), .Z(n46436) );
  IV U66632 ( .A(n46436), .Z(n46437) );
  NOR U66633 ( .A(n46438), .B(n46437), .Z(n46439) );
  XOR U66634 ( .A(n51490), .B(n46439), .Z(n51484) );
  XOR U66635 ( .A(n46440), .B(n51484), .Z(n51954) );
  XOR U66636 ( .A(n46441), .B(n51954), .Z(n46442) );
  IV U66637 ( .A(n46442), .Z(n51482) );
  XOR U66638 ( .A(n51481), .B(n51482), .Z(n51479) );
  XOR U66639 ( .A(n51476), .B(n51479), .Z(n46443) );
  NOR U66640 ( .A(n46444), .B(n46443), .Z(n57139) );
  IV U66641 ( .A(n46445), .Z(n46446) );
  NOR U66642 ( .A(n46447), .B(n46446), .Z(n51478) );
  NOR U66643 ( .A(n51478), .B(n51476), .Z(n46448) );
  XOR U66644 ( .A(n46448), .B(n51479), .Z(n46459) );
  NOR U66645 ( .A(n46449), .B(n46459), .Z(n46450) );
  NOR U66646 ( .A(n57139), .B(n46450), .Z(n46453) );
  NOR U66647 ( .A(n46451), .B(n46453), .Z(n46467) );
  IV U66648 ( .A(n46452), .Z(n46457) );
  IV U66649 ( .A(n46453), .Z(n46454) );
  NOR U66650 ( .A(n46461), .B(n46454), .Z(n46455) );
  IV U66651 ( .A(n46455), .Z(n46456) );
  NOR U66652 ( .A(n46457), .B(n46456), .Z(n56758) );
  IV U66653 ( .A(n46458), .Z(n46464) );
  IV U66654 ( .A(n46459), .Z(n46460) );
  NOR U66655 ( .A(n46461), .B(n46460), .Z(n46462) );
  IV U66656 ( .A(n46462), .Z(n46463) );
  NOR U66657 ( .A(n46464), .B(n46463), .Z(n57137) );
  NOR U66658 ( .A(n56758), .B(n57137), .Z(n46465) );
  IV U66659 ( .A(n46465), .Z(n46466) );
  NOR U66660 ( .A(n46467), .B(n46466), .Z(n51474) );
  XOR U66661 ( .A(n46468), .B(n51474), .Z(n57148) );
  XOR U66662 ( .A(n57151), .B(n57148), .Z(n46469) );
  XOR U66663 ( .A(n46470), .B(n46469), .Z(n51464) );
  IV U66664 ( .A(n46471), .Z(n56742) );
  NOR U66665 ( .A(n46472), .B(n56742), .Z(n51471) );
  NOR U66666 ( .A(n46473), .B(n51465), .Z(n46474) );
  NOR U66667 ( .A(n51471), .B(n46474), .Z(n46475) );
  XOR U66668 ( .A(n51464), .B(n46475), .Z(n51972) );
  IV U66669 ( .A(n51972), .Z(n46485) );
  IV U66670 ( .A(n46476), .Z(n51459) );
  NOR U66671 ( .A(n46477), .B(n51459), .Z(n46484) );
  IV U66672 ( .A(n46478), .Z(n46480) );
  NOR U66673 ( .A(n46480), .B(n46479), .Z(n51457) );
  NOR U66674 ( .A(n46484), .B(n51457), .Z(n46481) );
  XOR U66675 ( .A(n46485), .B(n46481), .Z(n51982) );
  IV U66676 ( .A(n46482), .Z(n51983) );
  IV U66677 ( .A(n46484), .Z(n51973) );
  XOR U66678 ( .A(n51973), .B(n46485), .Z(n51449) );
  IV U66679 ( .A(n46487), .Z(n46489) );
  NOR U66680 ( .A(n46489), .B(n46488), .Z(n46497) );
  IV U66681 ( .A(n46497), .Z(n46490) );
  NOR U66682 ( .A(n51988), .B(n46490), .Z(n56715) );
  IV U66683 ( .A(n46491), .Z(n46492) );
  NOR U66684 ( .A(n46492), .B(n46494), .Z(n51986) );
  XOR U66685 ( .A(n51986), .B(n51988), .Z(n51446) );
  IV U66686 ( .A(n46493), .Z(n46495) );
  NOR U66687 ( .A(n46495), .B(n46494), .Z(n51444) );
  XOR U66688 ( .A(n51446), .B(n51444), .Z(n56708) );
  IV U66689 ( .A(n56708), .Z(n46496) );
  NOR U66690 ( .A(n46497), .B(n46496), .Z(n46498) );
  NOR U66691 ( .A(n56715), .B(n46498), .Z(n46499) );
  NOR U66692 ( .A(n46500), .B(n46499), .Z(n46502) );
  IV U66693 ( .A(n46500), .Z(n46501) );
  NOR U66694 ( .A(n46501), .B(n56708), .Z(n56704) );
  NOR U66695 ( .A(n46502), .B(n56704), .Z(n51438) );
  IV U66696 ( .A(n46503), .Z(n46504) );
  NOR U66697 ( .A(n46505), .B(n46504), .Z(n46506) );
  IV U66698 ( .A(n46506), .Z(n56711) );
  XOR U66699 ( .A(n51438), .B(n56711), .Z(n51441) );
  XOR U66700 ( .A(n51440), .B(n51441), .Z(n51434) );
  XOR U66701 ( .A(n51433), .B(n51434), .Z(n51437) );
  XOR U66702 ( .A(n51436), .B(n51437), .Z(n46513) );
  IV U66703 ( .A(n46513), .Z(n57179) );
  NOR U66704 ( .A(n46507), .B(n57179), .Z(n56697) );
  IV U66705 ( .A(n46508), .Z(n46511) );
  IV U66706 ( .A(n46509), .Z(n46510) );
  NOR U66707 ( .A(n46511), .B(n46510), .Z(n46514) );
  IV U66708 ( .A(n46514), .Z(n46512) );
  NOR U66709 ( .A(n46512), .B(n51434), .Z(n57171) );
  NOR U66710 ( .A(n46514), .B(n46513), .Z(n46515) );
  NOR U66711 ( .A(n57171), .B(n46515), .Z(n46516) );
  NOR U66712 ( .A(n46517), .B(n46516), .Z(n46518) );
  NOR U66713 ( .A(n56697), .B(n46518), .Z(n51427) );
  IV U66714 ( .A(n46519), .Z(n46520) );
  NOR U66715 ( .A(n46521), .B(n46520), .Z(n46522) );
  IV U66716 ( .A(n46522), .Z(n57182) );
  XOR U66717 ( .A(n51427), .B(n57182), .Z(n51431) );
  XOR U66718 ( .A(n51429), .B(n51431), .Z(n51420) );
  XOR U66719 ( .A(n46523), .B(n51420), .Z(n46524) );
  IV U66720 ( .A(n46524), .Z(n51412) );
  NOR U66721 ( .A(n46525), .B(n51412), .Z(n51998) );
  IV U66722 ( .A(n51998), .Z(n56693) );
  IV U66723 ( .A(n46526), .Z(n51410) );
  IV U66724 ( .A(n46527), .Z(n46529) );
  NOR U66725 ( .A(n46529), .B(n46528), .Z(n46530) );
  IV U66726 ( .A(n46530), .Z(n51413) );
  XOR U66727 ( .A(n51413), .B(n51412), .Z(n46531) );
  NOR U66728 ( .A(n46532), .B(n46531), .Z(n51411) );
  IV U66729 ( .A(n46533), .Z(n46534) );
  NOR U66730 ( .A(n46534), .B(n51412), .Z(n56690) );
  IV U66731 ( .A(n46539), .Z(n56681) );
  NOR U66732 ( .A(n46535), .B(n56681), .Z(n56677) );
  IV U66733 ( .A(n46536), .Z(n46538) );
  NOR U66734 ( .A(n46538), .B(n46537), .Z(n56680) );
  NOR U66735 ( .A(n56684), .B(n56680), .Z(n51999) );
  XOR U66736 ( .A(n51999), .B(n46539), .Z(n51406) );
  IV U66737 ( .A(n51406), .Z(n46540) );
  NOR U66738 ( .A(n46541), .B(n46540), .Z(n46542) );
  NOR U66739 ( .A(n56677), .B(n46542), .Z(n46543) );
  IV U66740 ( .A(n46543), .Z(n52004) );
  XOR U66741 ( .A(n52003), .B(n52004), .Z(n52021) );
  IV U66742 ( .A(n52021), .Z(n46546) );
  IV U66743 ( .A(n46544), .Z(n51407) );
  NOR U66744 ( .A(n46545), .B(n51407), .Z(n46547) );
  NOR U66745 ( .A(n46546), .B(n46547), .Z(n46550) );
  IV U66746 ( .A(n46547), .Z(n46548) );
  NOR U66747 ( .A(n46548), .B(n51406), .Z(n46549) );
  NOR U66748 ( .A(n46550), .B(n46549), .Z(n52034) );
  NOR U66749 ( .A(n46551), .B(n52024), .Z(n52015) );
  IV U66750 ( .A(n46552), .Z(n46554) );
  NOR U66751 ( .A(n46554), .B(n46553), .Z(n52035) );
  NOR U66752 ( .A(n52015), .B(n52035), .Z(n46555) );
  XOR U66753 ( .A(n52034), .B(n46555), .Z(n56664) );
  XOR U66754 ( .A(n51403), .B(n56664), .Z(n51399) );
  XOR U66755 ( .A(n51390), .B(n51399), .Z(n52042) );
  XOR U66756 ( .A(n51387), .B(n52042), .Z(n46556) );
  XOR U66757 ( .A(n46557), .B(n46556), .Z(n51386) );
  XOR U66758 ( .A(n51384), .B(n51386), .Z(n52045) );
  XOR U66759 ( .A(n52044), .B(n52045), .Z(n52049) );
  XOR U66760 ( .A(n52047), .B(n52049), .Z(n51378) );
  XOR U66761 ( .A(n46558), .B(n51378), .Z(n51371) );
  XOR U66762 ( .A(n46559), .B(n51371), .Z(n51370) );
  IV U66763 ( .A(n51370), .Z(n46566) );
  IV U66764 ( .A(n46560), .Z(n46562) );
  NOR U66765 ( .A(n46562), .B(n46561), .Z(n51368) );
  IV U66766 ( .A(n46563), .Z(n51365) );
  NOR U66767 ( .A(n51365), .B(n51367), .Z(n46564) );
  NOR U66768 ( .A(n51368), .B(n46564), .Z(n46565) );
  XOR U66769 ( .A(n46566), .B(n46565), .Z(n51362) );
  XOR U66770 ( .A(n51361), .B(n51362), .Z(n52060) );
  IV U66771 ( .A(n52060), .Z(n46567) );
  NOR U66772 ( .A(n46568), .B(n46567), .Z(n52063) );
  IV U66773 ( .A(n46568), .Z(n46569) );
  NOR U66774 ( .A(n46569), .B(n51362), .Z(n57262) );
  NOR U66775 ( .A(n52063), .B(n57262), .Z(n51360) );
  XOR U66776 ( .A(n46570), .B(n51360), .Z(n56630) );
  XOR U66777 ( .A(n52073), .B(n56630), .Z(n51356) );
  XOR U66778 ( .A(n51358), .B(n51356), .Z(n52071) );
  XOR U66779 ( .A(n52070), .B(n52071), .Z(n51353) );
  XOR U66780 ( .A(n46571), .B(n51353), .Z(n52080) );
  XOR U66781 ( .A(n46572), .B(n52080), .Z(n52089) );
  XOR U66782 ( .A(n52088), .B(n52089), .Z(n52084) );
  XOR U66783 ( .A(n46573), .B(n52084), .Z(n56593) );
  XOR U66784 ( .A(n52099), .B(n56593), .Z(n46582) );
  IV U66785 ( .A(n46582), .Z(n56586) );
  IV U66786 ( .A(n46574), .Z(n46576) );
  NOR U66787 ( .A(n46576), .B(n46575), .Z(n46591) );
  IV U66788 ( .A(n46591), .Z(n57277) );
  NOR U66789 ( .A(n56586), .B(n57277), .Z(n52104) );
  IV U66790 ( .A(n46577), .Z(n46579) );
  NOR U66791 ( .A(n46580), .B(n56593), .Z(n46578) );
  IV U66792 ( .A(n46578), .Z(n46585) );
  NOR U66793 ( .A(n46579), .B(n46585), .Z(n56589) );
  NOR U66794 ( .A(n46581), .B(n46580), .Z(n46583) );
  NOR U66795 ( .A(n46583), .B(n46582), .Z(n46587) );
  IV U66796 ( .A(n46584), .Z(n46586) );
  NOR U66797 ( .A(n46586), .B(n46585), .Z(n51349) );
  NOR U66798 ( .A(n46587), .B(n51349), .Z(n46588) );
  IV U66799 ( .A(n46588), .Z(n46589) );
  NOR U66800 ( .A(n56589), .B(n46589), .Z(n46590) );
  NOR U66801 ( .A(n46591), .B(n46590), .Z(n46592) );
  NOR U66802 ( .A(n52104), .B(n46592), .Z(n52102) );
  XOR U66803 ( .A(n56588), .B(n52102), .Z(n51346) );
  XOR U66804 ( .A(n46593), .B(n51346), .Z(n51344) );
  XOR U66805 ( .A(n51342), .B(n51344), .Z(n52110) );
  IV U66806 ( .A(n46594), .Z(n46596) );
  NOR U66807 ( .A(n46596), .B(n46595), .Z(n51340) );
  XOR U66808 ( .A(n52110), .B(n51340), .Z(n46609) );
  NOR U66809 ( .A(n46609), .B(n46605), .Z(n46597) );
  IV U66810 ( .A(n46597), .Z(n56573) );
  NOR U66811 ( .A(n46606), .B(n56573), .Z(n56564) );
  IV U66812 ( .A(n46598), .Z(n46601) );
  NOR U66813 ( .A(n46599), .B(n46601), .Z(n52117) );
  IV U66814 ( .A(n46600), .Z(n46602) );
  NOR U66815 ( .A(n46602), .B(n46601), .Z(n51338) );
  NOR U66816 ( .A(n52117), .B(n51338), .Z(n46615) );
  IV U66817 ( .A(n46615), .Z(n46603) );
  NOR U66818 ( .A(n56564), .B(n46603), .Z(n46604) );
  IV U66819 ( .A(n46604), .Z(n46613) );
  NOR U66820 ( .A(n46606), .B(n46605), .Z(n46611) );
  IV U66821 ( .A(n46607), .Z(n52111) );
  NOR U66822 ( .A(n52111), .B(n46608), .Z(n46610) );
  XOR U66823 ( .A(n46610), .B(n46609), .Z(n52119) );
  IV U66824 ( .A(n52119), .Z(n46614) );
  NOR U66825 ( .A(n46611), .B(n46614), .Z(n46612) );
  NOR U66826 ( .A(n46613), .B(n46612), .Z(n46617) );
  NOR U66827 ( .A(n46615), .B(n46614), .Z(n46616) );
  NOR U66828 ( .A(n46617), .B(n46616), .Z(n51337) );
  XOR U66829 ( .A(n51335), .B(n51337), .Z(n51321) );
  XOR U66830 ( .A(n51322), .B(n51321), .Z(n51309) );
  IV U66831 ( .A(n51309), .Z(n46625) );
  IV U66832 ( .A(n46618), .Z(n46619) );
  NOR U66833 ( .A(n46620), .B(n46619), .Z(n46623) );
  NOR U66834 ( .A(n46621), .B(n51308), .Z(n46622) );
  NOR U66835 ( .A(n46623), .B(n46622), .Z(n46624) );
  XOR U66836 ( .A(n46625), .B(n46624), .Z(n56537) );
  XOR U66837 ( .A(n51305), .B(n56537), .Z(n51296) );
  NOR U66838 ( .A(n46626), .B(n51299), .Z(n46628) );
  IV U66839 ( .A(n46627), .Z(n46631) );
  IV U66840 ( .A(n46630), .Z(n46642) );
  NOR U66841 ( .A(n46631), .B(n46642), .Z(n51295) );
  NOR U66842 ( .A(n46628), .B(n51295), .Z(n46629) );
  XOR U66843 ( .A(n51296), .B(n46629), .Z(n46644) );
  IV U66844 ( .A(n46644), .Z(n46633) );
  XOR U66845 ( .A(n46631), .B(n46630), .Z(n46632) );
  NOR U66846 ( .A(n46633), .B(n46632), .Z(n46638) );
  IV U66847 ( .A(n46634), .Z(n46639) );
  NOR U66848 ( .A(n46639), .B(n46635), .Z(n46636) );
  IV U66849 ( .A(n46636), .Z(n46637) );
  NOR U66850 ( .A(n46638), .B(n46637), .Z(n46649) );
  IV U66851 ( .A(n46638), .Z(n46641) );
  NOR U66852 ( .A(n46639), .B(n46641), .Z(n57301) );
  IV U66853 ( .A(n46640), .Z(n46643) );
  NOR U66854 ( .A(n46643), .B(n46641), .Z(n56515) );
  NOR U66855 ( .A(n57301), .B(n56515), .Z(n52128) );
  IV U66856 ( .A(n52128), .Z(n46647) );
  NOR U66857 ( .A(n46643), .B(n46642), .Z(n46645) );
  NOR U66858 ( .A(n46645), .B(n46644), .Z(n46646) );
  NOR U66859 ( .A(n46647), .B(n46646), .Z(n46648) );
  NOR U66860 ( .A(n46649), .B(n46648), .Z(n51291) );
  XOR U66861 ( .A(n51289), .B(n51291), .Z(n51294) );
  XOR U66862 ( .A(n51292), .B(n51294), .Z(n52131) );
  XOR U66863 ( .A(n52130), .B(n52131), .Z(n52134) );
  XOR U66864 ( .A(n52133), .B(n52134), .Z(n51284) );
  XOR U66865 ( .A(n46650), .B(n51284), .Z(n46654) );
  IV U66866 ( .A(n46654), .Z(n56487) );
  NOR U66867 ( .A(n46651), .B(n56487), .Z(n52138) );
  NOR U66868 ( .A(n46662), .B(n52138), .Z(n46652) );
  IV U66869 ( .A(n46652), .Z(n46661) );
  NOR U66870 ( .A(n46653), .B(n51270), .Z(n46655) );
  NOR U66871 ( .A(n46655), .B(n46654), .Z(n46658) );
  XOR U66872 ( .A(n51281), .B(n51284), .Z(n51269) );
  IV U66873 ( .A(n46655), .Z(n46656) );
  NOR U66874 ( .A(n51269), .B(n46656), .Z(n46657) );
  NOR U66875 ( .A(n46658), .B(n46657), .Z(n51260) );
  NOR U66876 ( .A(n46659), .B(n51260), .Z(n46660) );
  NOR U66877 ( .A(n46661), .B(n46660), .Z(n46665) );
  IV U66878 ( .A(n46662), .Z(n46663) );
  NOR U66879 ( .A(n51260), .B(n46663), .Z(n46664) );
  NOR U66880 ( .A(n46665), .B(n46664), .Z(n52141) );
  XOR U66881 ( .A(n52139), .B(n52141), .Z(n52144) );
  XOR U66882 ( .A(n52142), .B(n52144), .Z(n52150) );
  XOR U66883 ( .A(n52151), .B(n52150), .Z(n51253) );
  IV U66884 ( .A(n46666), .Z(n46668) );
  NOR U66885 ( .A(n46668), .B(n46667), .Z(n51255) );
  IV U66886 ( .A(n46669), .Z(n46670) );
  NOR U66887 ( .A(n46671), .B(n46670), .Z(n52147) );
  NOR U66888 ( .A(n51255), .B(n52147), .Z(n46672) );
  XOR U66889 ( .A(n51253), .B(n46672), .Z(n52163) );
  XOR U66890 ( .A(n46673), .B(n52163), .Z(n52169) );
  XOR U66891 ( .A(n52168), .B(n52169), .Z(n51246) );
  XOR U66892 ( .A(n51245), .B(n51246), .Z(n51249) );
  XOR U66893 ( .A(n51248), .B(n51249), .Z(n51244) );
  XOR U66894 ( .A(n46674), .B(n51244), .Z(n51233) );
  XOR U66895 ( .A(n46675), .B(n51233), .Z(n52193) );
  IV U66896 ( .A(n46676), .Z(n46678) );
  NOR U66897 ( .A(n46678), .B(n46677), .Z(n52191) );
  XOR U66898 ( .A(n52193), .B(n52191), .Z(n52195) );
  XOR U66899 ( .A(n52194), .B(n52195), .Z(n51221) );
  IV U66900 ( .A(n46679), .Z(n51229) );
  NOR U66901 ( .A(n51229), .B(n46680), .Z(n51218) );
  NOR U66902 ( .A(n46681), .B(n51222), .Z(n46682) );
  NOR U66903 ( .A(n51218), .B(n46682), .Z(n46683) );
  XOR U66904 ( .A(n51221), .B(n46683), .Z(n51212) );
  XOR U66905 ( .A(n46684), .B(n51212), .Z(n52203) );
  XOR U66906 ( .A(n46685), .B(n52203), .Z(n51195) );
  IV U66907 ( .A(n46686), .Z(n46687) );
  NOR U66908 ( .A(n46688), .B(n46687), .Z(n51199) );
  NOR U66909 ( .A(n46689), .B(n51196), .Z(n46690) );
  NOR U66910 ( .A(n51199), .B(n46690), .Z(n46691) );
  XOR U66911 ( .A(n51195), .B(n46691), .Z(n52218) );
  XOR U66912 ( .A(n46692), .B(n52218), .Z(n52224) );
  XOR U66913 ( .A(n52225), .B(n52224), .Z(n57356) );
  IV U66914 ( .A(n46693), .Z(n46694) );
  NOR U66915 ( .A(n46695), .B(n46694), .Z(n51189) );
  IV U66916 ( .A(n46696), .Z(n46698) );
  NOR U66917 ( .A(n46698), .B(n46697), .Z(n52227) );
  NOR U66918 ( .A(n51189), .B(n52227), .Z(n46699) );
  XOR U66919 ( .A(n57356), .B(n46699), .Z(n46707) );
  XOR U66920 ( .A(n46700), .B(n46707), .Z(n51183) );
  IV U66921 ( .A(n46701), .Z(n46703) );
  NOR U66922 ( .A(n46703), .B(n46702), .Z(n46704) );
  IV U66923 ( .A(n46704), .Z(n51182) );
  XOR U66924 ( .A(n51183), .B(n51182), .Z(n46705) );
  NOR U66925 ( .A(n46706), .B(n46705), .Z(n46709) );
  IV U66926 ( .A(n46706), .Z(n46708) );
  IV U66927 ( .A(n46707), .Z(n51191) );
  XOR U66928 ( .A(n51190), .B(n51191), .Z(n51185) );
  XOR U66929 ( .A(n51184), .B(n51185), .Z(n57382) );
  NOR U66930 ( .A(n46708), .B(n57382), .Z(n57377) );
  NOR U66931 ( .A(n46709), .B(n57377), .Z(n51177) );
  XOR U66932 ( .A(n46710), .B(n51177), .Z(n51175) );
  IV U66933 ( .A(n46711), .Z(n46713) );
  NOR U66934 ( .A(n46713), .B(n46712), .Z(n51173) );
  XOR U66935 ( .A(n51175), .B(n51173), .Z(n51159) );
  XOR U66936 ( .A(n51160), .B(n51159), .Z(n52238) );
  XOR U66937 ( .A(n46714), .B(n52238), .Z(n46721) );
  IV U66938 ( .A(n46721), .Z(n56358) );
  NOR U66939 ( .A(n46722), .B(n56358), .Z(n52240) );
  IV U66940 ( .A(n46715), .Z(n46728) );
  NOR U66941 ( .A(n46716), .B(n46728), .Z(n52243) );
  IV U66942 ( .A(n46717), .Z(n46719) );
  NOR U66943 ( .A(n46719), .B(n46718), .Z(n46720) );
  IV U66944 ( .A(n46720), .Z(n52239) );
  XOR U66945 ( .A(n52239), .B(n46721), .Z(n52244) );
  IV U66946 ( .A(n52244), .Z(n46723) );
  XOR U66947 ( .A(n52243), .B(n46723), .Z(n46725) );
  NOR U66948 ( .A(n46723), .B(n46722), .Z(n46724) );
  NOR U66949 ( .A(n46725), .B(n46724), .Z(n46726) );
  NOR U66950 ( .A(n52240), .B(n46726), .Z(n52247) );
  IV U66951 ( .A(n46727), .Z(n46729) );
  NOR U66952 ( .A(n46729), .B(n46728), .Z(n52246) );
  NOR U66953 ( .A(n52246), .B(n46730), .Z(n46731) );
  XOR U66954 ( .A(n52247), .B(n46731), .Z(n52252) );
  XOR U66955 ( .A(n52251), .B(n52252), .Z(n52258) );
  XOR U66956 ( .A(n51152), .B(n52258), .Z(n46732) );
  IV U66957 ( .A(n46732), .Z(n52263) );
  IV U66958 ( .A(n46733), .Z(n46734) );
  NOR U66959 ( .A(n46735), .B(n46734), .Z(n52261) );
  XOR U66960 ( .A(n52263), .B(n52261), .Z(n51150) );
  IV U66961 ( .A(n46736), .Z(n46738) );
  NOR U66962 ( .A(n46738), .B(n46737), .Z(n51148) );
  XOR U66963 ( .A(n51150), .B(n51148), .Z(n52259) );
  XOR U66964 ( .A(n52260), .B(n52259), .Z(n46739) );
  NOR U66965 ( .A(n46744), .B(n46739), .Z(n46749) );
  IV U66966 ( .A(n46740), .Z(n46741) );
  NOR U66967 ( .A(n46742), .B(n46741), .Z(n46753) );
  IV U66968 ( .A(n46753), .Z(n46743) );
  NOR U66969 ( .A(n46749), .B(n46743), .Z(n51146) );
  IV U66970 ( .A(n46744), .Z(n46745) );
  NOR U66971 ( .A(n46745), .B(n51150), .Z(n62516) );
  IV U66972 ( .A(n46746), .Z(n46747) );
  NOR U66973 ( .A(n52270), .B(n46747), .Z(n46750) );
  IV U66974 ( .A(n46750), .Z(n46748) );
  NOR U66975 ( .A(n46748), .B(n51150), .Z(n61414) );
  NOR U66976 ( .A(n62516), .B(n61414), .Z(n56330) );
  IV U66977 ( .A(n56330), .Z(n52278) );
  IV U66978 ( .A(n46749), .Z(n46751) );
  NOR U66979 ( .A(n46751), .B(n46750), .Z(n46752) );
  NOR U66980 ( .A(n52278), .B(n46752), .Z(n52272) );
  NOR U66981 ( .A(n46753), .B(n52272), .Z(n46754) );
  NOR U66982 ( .A(n51146), .B(n46754), .Z(n51129) );
  IV U66983 ( .A(n46755), .Z(n46756) );
  NOR U66984 ( .A(n57411), .B(n46756), .Z(n51144) );
  NOR U66985 ( .A(n46757), .B(n51138), .Z(n51131) );
  NOR U66986 ( .A(n51144), .B(n51131), .Z(n46758) );
  XOR U66987 ( .A(n51129), .B(n46758), .Z(n57432) );
  XOR U66988 ( .A(n57433), .B(n57432), .Z(n46763) );
  IV U66989 ( .A(n46759), .Z(n46761) );
  NOR U66990 ( .A(n46761), .B(n46760), .Z(n46768) );
  IV U66991 ( .A(n46768), .Z(n46762) );
  NOR U66992 ( .A(n46763), .B(n46762), .Z(n56310) );
  NOR U66993 ( .A(n46765), .B(n46764), .Z(n51124) );
  NOR U66994 ( .A(n57433), .B(n51124), .Z(n46766) );
  XOR U66995 ( .A(n57432), .B(n46766), .Z(n46767) );
  NOR U66996 ( .A(n46768), .B(n46767), .Z(n46769) );
  NOR U66997 ( .A(n56310), .B(n46769), .Z(n52284) );
  XOR U66998 ( .A(n52285), .B(n52284), .Z(n51122) );
  XOR U66999 ( .A(n46770), .B(n51122), .Z(n46771) );
  IV U67000 ( .A(n46771), .Z(n66966) );
  XOR U67001 ( .A(n51117), .B(n66966), .Z(n52299) );
  IV U67002 ( .A(n46772), .Z(n46774) );
  IV U67003 ( .A(n46773), .Z(n46776) );
  NOR U67004 ( .A(n46774), .B(n46776), .Z(n52296) );
  NOR U67005 ( .A(n46775), .B(n66968), .Z(n51119) );
  NOR U67006 ( .A(n46777), .B(n46776), .Z(n52298) );
  NOR U67007 ( .A(n51119), .B(n52298), .Z(n46778) );
  IV U67008 ( .A(n46778), .Z(n46779) );
  NOR U67009 ( .A(n52296), .B(n46779), .Z(n46780) );
  XOR U67010 ( .A(n52299), .B(n46780), .Z(n46781) );
  IV U67011 ( .A(n46781), .Z(n52304) );
  IV U67012 ( .A(n46782), .Z(n46784) );
  NOR U67013 ( .A(n46784), .B(n46783), .Z(n51115) );
  XOR U67014 ( .A(n52304), .B(n51115), .Z(n52307) );
  XOR U67015 ( .A(n52306), .B(n52307), .Z(n51114) );
  XOR U67016 ( .A(n46785), .B(n51114), .Z(n51108) );
  XOR U67017 ( .A(n52314), .B(n51108), .Z(n52323) );
  XOR U67018 ( .A(n46786), .B(n52323), .Z(n46787) );
  IV U67019 ( .A(n46787), .Z(n51102) );
  XOR U67020 ( .A(n51100), .B(n51102), .Z(n51104) );
  XOR U67021 ( .A(n51097), .B(n51104), .Z(n46788) );
  XOR U67022 ( .A(n46789), .B(n46788), .Z(n52331) );
  IV U67023 ( .A(n46790), .Z(n46791) );
  NOR U67024 ( .A(n52329), .B(n46791), .Z(n46794) );
  NOR U67025 ( .A(n51090), .B(n46792), .Z(n46793) );
  NOR U67026 ( .A(n46794), .B(n46793), .Z(n46795) );
  XOR U67027 ( .A(n52331), .B(n46795), .Z(n51088) );
  IV U67028 ( .A(n46796), .Z(n46797) );
  NOR U67029 ( .A(n46797), .B(n46813), .Z(n46805) );
  IV U67030 ( .A(n46805), .Z(n46798) );
  NOR U67031 ( .A(n51088), .B(n46798), .Z(n57505) );
  IV U67032 ( .A(n46799), .Z(n46800) );
  NOR U67033 ( .A(n46803), .B(n46800), .Z(n51093) );
  IV U67034 ( .A(n46801), .Z(n46802) );
  NOR U67035 ( .A(n46803), .B(n46802), .Z(n51086) );
  XOR U67036 ( .A(n51086), .B(n51088), .Z(n51094) );
  XOR U67037 ( .A(n51093), .B(n51094), .Z(n46816) );
  IV U67038 ( .A(n46816), .Z(n46804) );
  NOR U67039 ( .A(n46805), .B(n46804), .Z(n46806) );
  NOR U67040 ( .A(n57505), .B(n46806), .Z(n46818) );
  IV U67041 ( .A(n46818), .Z(n46811) );
  IV U67042 ( .A(n46807), .Z(n46809) );
  NOR U67043 ( .A(n46809), .B(n46808), .Z(n46810) );
  IV U67044 ( .A(n46810), .Z(n46822) );
  NOR U67045 ( .A(n46811), .B(n46822), .Z(n56273) );
  IV U67046 ( .A(n46812), .Z(n46814) );
  NOR U67047 ( .A(n46814), .B(n46813), .Z(n46817) );
  IV U67048 ( .A(n46817), .Z(n46815) );
  NOR U67049 ( .A(n46816), .B(n46815), .Z(n61363) );
  NOR U67050 ( .A(n46818), .B(n46817), .Z(n46819) );
  NOR U67051 ( .A(n61363), .B(n46819), .Z(n51080) );
  IV U67052 ( .A(n46820), .Z(n46821) );
  NOR U67053 ( .A(n46831), .B(n46821), .Z(n51081) );
  XOR U67054 ( .A(n51080), .B(n51081), .Z(n46824) );
  NOR U67055 ( .A(n51081), .B(n46822), .Z(n46823) );
  NOR U67056 ( .A(n46824), .B(n46823), .Z(n46825) );
  NOR U67057 ( .A(n56273), .B(n46825), .Z(n51074) );
  IV U67058 ( .A(n46826), .Z(n46828) );
  NOR U67059 ( .A(n46828), .B(n46827), .Z(n46829) );
  IV U67060 ( .A(n46829), .Z(n46830) );
  NOR U67061 ( .A(n46831), .B(n46830), .Z(n46832) );
  IV U67062 ( .A(n46832), .Z(n51078) );
  XOR U67063 ( .A(n51074), .B(n51078), .Z(n51069) );
  IV U67064 ( .A(n51069), .Z(n46839) );
  NOR U67065 ( .A(n51075), .B(n46833), .Z(n46837) );
  IV U67066 ( .A(n46834), .Z(n51070) );
  NOR U67067 ( .A(n46835), .B(n51070), .Z(n46836) );
  NOR U67068 ( .A(n46837), .B(n46836), .Z(n46838) );
  XOR U67069 ( .A(n46839), .B(n46838), .Z(n51067) );
  XOR U67070 ( .A(n51063), .B(n51067), .Z(n51058) );
  XOR U67071 ( .A(n51059), .B(n51058), .Z(n52358) );
  IV U67072 ( .A(n46840), .Z(n46843) );
  IV U67073 ( .A(n46841), .Z(n46842) );
  NOR U67074 ( .A(n46843), .B(n46842), .Z(n46844) );
  IV U67075 ( .A(n46844), .Z(n52359) );
  XOR U67076 ( .A(n52358), .B(n52359), .Z(n52361) );
  IV U67077 ( .A(n46845), .Z(n46846) );
  NOR U67078 ( .A(n52366), .B(n46846), .Z(n52360) );
  NOR U67079 ( .A(n46847), .B(n51054), .Z(n46848) );
  NOR U67080 ( .A(n52360), .B(n46848), .Z(n46849) );
  XOR U67081 ( .A(n52361), .B(n46849), .Z(n46859) );
  IV U67082 ( .A(n46859), .Z(n46858) );
  XOR U67083 ( .A(n46860), .B(n46858), .Z(n57540) );
  IV U67084 ( .A(n46850), .Z(n46851) );
  NOR U67085 ( .A(n46852), .B(n46851), .Z(n46867) );
  IV U67086 ( .A(n46867), .Z(n46853) );
  NOR U67087 ( .A(n57540), .B(n46853), .Z(n57532) );
  IV U67088 ( .A(n46854), .Z(n46856) );
  NOR U67089 ( .A(n46856), .B(n46855), .Z(n51048) );
  IV U67090 ( .A(n46860), .Z(n46857) );
  NOR U67091 ( .A(n46858), .B(n46857), .Z(n57523) );
  NOR U67092 ( .A(n46860), .B(n46859), .Z(n46864) );
  IV U67093 ( .A(n46861), .Z(n46863) );
  NOR U67094 ( .A(n46863), .B(n46862), .Z(n51045) );
  XOR U67095 ( .A(n46864), .B(n51045), .Z(n46865) );
  NOR U67096 ( .A(n57523), .B(n46865), .Z(n51049) );
  XOR U67097 ( .A(n51048), .B(n51049), .Z(n46866) );
  NOR U67098 ( .A(n46867), .B(n46866), .Z(n46868) );
  NOR U67099 ( .A(n57532), .B(n46868), .Z(n51043) );
  XOR U67100 ( .A(n46869), .B(n51043), .Z(n52377) );
  XOR U67101 ( .A(n46870), .B(n52377), .Z(n46882) );
  IV U67102 ( .A(n46882), .Z(n46875) );
  NOR U67103 ( .A(n46871), .B(n46875), .Z(n56239) );
  IV U67104 ( .A(n46872), .Z(n46873) );
  NOR U67105 ( .A(n46874), .B(n46873), .Z(n46884) );
  IV U67106 ( .A(n46884), .Z(n46876) );
  NOR U67107 ( .A(n46876), .B(n46875), .Z(n56242) );
  IV U67108 ( .A(n46877), .Z(n46879) );
  NOR U67109 ( .A(n46879), .B(n46878), .Z(n46881) );
  IV U67110 ( .A(n46881), .Z(n46880) );
  NOR U67111 ( .A(n52377), .B(n46880), .Z(n56248) );
  NOR U67112 ( .A(n46882), .B(n46881), .Z(n46883) );
  NOR U67113 ( .A(n56248), .B(n46883), .Z(n46888) );
  NOR U67114 ( .A(n46885), .B(n46884), .Z(n46886) );
  IV U67115 ( .A(n46886), .Z(n46887) );
  NOR U67116 ( .A(n46888), .B(n46887), .Z(n46889) );
  NOR U67117 ( .A(n56242), .B(n46889), .Z(n46890) );
  IV U67118 ( .A(n46890), .Z(n46891) );
  NOR U67119 ( .A(n56239), .B(n46891), .Z(n51036) );
  IV U67120 ( .A(n46897), .Z(n51038) );
  NOR U67121 ( .A(n51036), .B(n51038), .Z(n46899) );
  IV U67122 ( .A(n46893), .Z(n46892) );
  NOR U67123 ( .A(n46892), .B(n46891), .Z(n56237) );
  NOR U67124 ( .A(n51036), .B(n46893), .Z(n46894) );
  NOR U67125 ( .A(n56237), .B(n46894), .Z(n46895) );
  IV U67126 ( .A(n46895), .Z(n46896) );
  NOR U67127 ( .A(n46897), .B(n46896), .Z(n46898) );
  NOR U67128 ( .A(n46899), .B(n46898), .Z(n51039) );
  NOR U67129 ( .A(n46900), .B(n51039), .Z(n56228) );
  IV U67130 ( .A(n46901), .Z(n46904) );
  IV U67131 ( .A(n46902), .Z(n46903) );
  NOR U67132 ( .A(n46904), .B(n46903), .Z(n46905) );
  IV U67133 ( .A(n46905), .Z(n51040) );
  XOR U67134 ( .A(n51040), .B(n51039), .Z(n46906) );
  NOR U67135 ( .A(n46907), .B(n46906), .Z(n51031) );
  IV U67136 ( .A(n46908), .Z(n46910) );
  NOR U67137 ( .A(n46910), .B(n46909), .Z(n51029) );
  XOR U67138 ( .A(n51031), .B(n51029), .Z(n46911) );
  NOR U67139 ( .A(n56228), .B(n46911), .Z(n51024) );
  XOR U67140 ( .A(n46912), .B(n51024), .Z(n51027) );
  XOR U67141 ( .A(n51026), .B(n51027), .Z(n51012) );
  IV U67142 ( .A(n51012), .Z(n46919) );
  NOR U67143 ( .A(n46913), .B(n51017), .Z(n46917) );
  IV U67144 ( .A(n46914), .Z(n51013) );
  NOR U67145 ( .A(n46915), .B(n51013), .Z(n46916) );
  NOR U67146 ( .A(n46917), .B(n46916), .Z(n46918) );
  XOR U67147 ( .A(n46919), .B(n46918), .Z(n56200) );
  XOR U67148 ( .A(n52393), .B(n56200), .Z(n52401) );
  XOR U67149 ( .A(n46920), .B(n52401), .Z(n52397) );
  XOR U67150 ( .A(n52398), .B(n52397), .Z(n52405) );
  XOR U67151 ( .A(n52404), .B(n52405), .Z(n52418) );
  IV U67152 ( .A(n46921), .Z(n52408) );
  NOR U67153 ( .A(n52408), .B(n46922), .Z(n46925) );
  IV U67154 ( .A(n46923), .Z(n46924) );
  NOR U67155 ( .A(n46924), .B(n46928), .Z(n52417) );
  NOR U67156 ( .A(n46925), .B(n52417), .Z(n46926) );
  XOR U67157 ( .A(n52418), .B(n46926), .Z(n51009) );
  IV U67158 ( .A(n46927), .Z(n46929) );
  NOR U67159 ( .A(n46929), .B(n46928), .Z(n56170) );
  IV U67160 ( .A(n46930), .Z(n46932) );
  NOR U67161 ( .A(n46932), .B(n46931), .Z(n56163) );
  NOR U67162 ( .A(n56170), .B(n56163), .Z(n51010) );
  XOR U67163 ( .A(n51009), .B(n51010), .Z(n52422) );
  XOR U67164 ( .A(n52421), .B(n52422), .Z(n52426) );
  IV U67165 ( .A(n46933), .Z(n46934) );
  NOR U67166 ( .A(n46934), .B(n46939), .Z(n52424) );
  XOR U67167 ( .A(n52426), .B(n52424), .Z(n51006) );
  IV U67168 ( .A(n46935), .Z(n46936) );
  NOR U67169 ( .A(n46937), .B(n46936), .Z(n51005) );
  IV U67170 ( .A(n46938), .Z(n46940) );
  NOR U67171 ( .A(n46940), .B(n46939), .Z(n51003) );
  NOR U67172 ( .A(n51005), .B(n51003), .Z(n46941) );
  XOR U67173 ( .A(n51006), .B(n46941), .Z(n46945) );
  IV U67174 ( .A(n46945), .Z(n56146) );
  XOR U67175 ( .A(n51001), .B(n56146), .Z(n46942) );
  NOR U67176 ( .A(n46943), .B(n46942), .Z(n61314) );
  NOR U67177 ( .A(n46944), .B(n56149), .Z(n50999) );
  NOR U67178 ( .A(n50999), .B(n51001), .Z(n46946) );
  XOR U67179 ( .A(n46946), .B(n46945), .Z(n50992) );
  IV U67180 ( .A(n50992), .Z(n46947) );
  NOR U67181 ( .A(n46948), .B(n46947), .Z(n46949) );
  NOR U67182 ( .A(n61314), .B(n46949), .Z(n52430) );
  IV U67183 ( .A(n46950), .Z(n46952) );
  NOR U67184 ( .A(n46952), .B(n46951), .Z(n46953) );
  IV U67185 ( .A(n46953), .Z(n52431) );
  XOR U67186 ( .A(n52430), .B(n52431), .Z(n50987) );
  NOR U67187 ( .A(n50993), .B(n46954), .Z(n46957) );
  IV U67188 ( .A(n46955), .Z(n50988) );
  NOR U67189 ( .A(n50990), .B(n50988), .Z(n46956) );
  NOR U67190 ( .A(n46957), .B(n46956), .Z(n46958) );
  XOR U67191 ( .A(n50987), .B(n46958), .Z(n50976) );
  NOR U67192 ( .A(n46959), .B(n50980), .Z(n46963) );
  IV U67193 ( .A(n46960), .Z(n46962) );
  NOR U67194 ( .A(n46962), .B(n46961), .Z(n50977) );
  NOR U67195 ( .A(n46963), .B(n50977), .Z(n46964) );
  XOR U67196 ( .A(n50976), .B(n46964), .Z(n50972) );
  XOR U67197 ( .A(n50971), .B(n50972), .Z(n52437) );
  XOR U67198 ( .A(n50974), .B(n52437), .Z(n50970) );
  IV U67199 ( .A(n50970), .Z(n46971) );
  IV U67200 ( .A(n46965), .Z(n46966) );
  NOR U67201 ( .A(n46974), .B(n46966), .Z(n52436) );
  IV U67202 ( .A(n46967), .Z(n46969) );
  NOR U67203 ( .A(n46969), .B(n46968), .Z(n50968) );
  NOR U67204 ( .A(n52436), .B(n50968), .Z(n46970) );
  XOR U67205 ( .A(n46971), .B(n46970), .Z(n52441) );
  IV U67206 ( .A(n46972), .Z(n46973) );
  NOR U67207 ( .A(n46974), .B(n46973), .Z(n52439) );
  XOR U67208 ( .A(n52441), .B(n52439), .Z(n57612) );
  XOR U67209 ( .A(n46975), .B(n57612), .Z(n50960) );
  XOR U67210 ( .A(n57615), .B(n50960), .Z(n50963) );
  XOR U67211 ( .A(n50962), .B(n50963), .Z(n50955) );
  XOR U67212 ( .A(n50954), .B(n50955), .Z(n50959) );
  IV U67213 ( .A(n50959), .Z(n46983) );
  IV U67214 ( .A(n46976), .Z(n46978) );
  NOR U67215 ( .A(n46978), .B(n46977), .Z(n50949) );
  IV U67216 ( .A(n46979), .Z(n46980) );
  NOR U67217 ( .A(n46981), .B(n46980), .Z(n50957) );
  NOR U67218 ( .A(n50949), .B(n50957), .Z(n46982) );
  XOR U67219 ( .A(n46983), .B(n46982), .Z(n50952) );
  XOR U67220 ( .A(n50951), .B(n50952), .Z(n52451) );
  XOR U67221 ( .A(n46984), .B(n52451), .Z(n52453) );
  XOR U67222 ( .A(n46985), .B(n52453), .Z(n50945) );
  XOR U67223 ( .A(n50943), .B(n50945), .Z(n56120) );
  XOR U67224 ( .A(n50946), .B(n56120), .Z(n46986) );
  XOR U67225 ( .A(n46987), .B(n46986), .Z(n50934) );
  XOR U67226 ( .A(n46997), .B(n50934), .Z(n46988) );
  NOR U67227 ( .A(n46989), .B(n46988), .Z(n57657) );
  IV U67228 ( .A(n46990), .Z(n46991) );
  NOR U67229 ( .A(n46992), .B(n46991), .Z(n46993) );
  IV U67230 ( .A(n46993), .Z(n52466) );
  IV U67231 ( .A(n46994), .Z(n46996) );
  NOR U67232 ( .A(n46996), .B(n46995), .Z(n52463) );
  IV U67233 ( .A(n46997), .Z(n46998) );
  NOR U67234 ( .A(n52463), .B(n46998), .Z(n46999) );
  XOR U67235 ( .A(n50934), .B(n46999), .Z(n52465) );
  XOR U67236 ( .A(n52466), .B(n52465), .Z(n47000) );
  NOR U67237 ( .A(n47001), .B(n47000), .Z(n47002) );
  NOR U67238 ( .A(n57657), .B(n47002), .Z(n52469) );
  XOR U67239 ( .A(n47003), .B(n52469), .Z(n52484) );
  XOR U67240 ( .A(n47004), .B(n52484), .Z(n50922) );
  XOR U67241 ( .A(n47005), .B(n50922), .Z(n50920) );
  XOR U67242 ( .A(n50918), .B(n50920), .Z(n50913) );
  IV U67243 ( .A(n47006), .Z(n47008) );
  NOR U67244 ( .A(n47008), .B(n47007), .Z(n50911) );
  XOR U67245 ( .A(n50913), .B(n50911), .Z(n50915) );
  IV U67246 ( .A(n47009), .Z(n47010) );
  NOR U67247 ( .A(n47013), .B(n47010), .Z(n50909) );
  IV U67248 ( .A(n47011), .Z(n47012) );
  NOR U67249 ( .A(n47013), .B(n47012), .Z(n50914) );
  NOR U67250 ( .A(n50909), .B(n50914), .Z(n47014) );
  XOR U67251 ( .A(n50915), .B(n47014), .Z(n50907) );
  IV U67252 ( .A(n47015), .Z(n47017) );
  NOR U67253 ( .A(n47017), .B(n47016), .Z(n50906) );
  NOR U67254 ( .A(n52491), .B(n50906), .Z(n47018) );
  XOR U67255 ( .A(n50907), .B(n47018), .Z(n50905) );
  XOR U67256 ( .A(n50903), .B(n50905), .Z(n50901) );
  XOR U67257 ( .A(n50899), .B(n50901), .Z(n47019) );
  XOR U67258 ( .A(n47020), .B(n47019), .Z(n52498) );
  IV U67259 ( .A(n47021), .Z(n47024) );
  IV U67260 ( .A(n47022), .Z(n47023) );
  NOR U67261 ( .A(n47024), .B(n47023), .Z(n52496) );
  XOR U67262 ( .A(n52498), .B(n52496), .Z(n52500) );
  IV U67263 ( .A(n52500), .Z(n47031) );
  IV U67264 ( .A(n47025), .Z(n47026) );
  NOR U67265 ( .A(n47029), .B(n47026), .Z(n50894) );
  IV U67266 ( .A(n47027), .Z(n47028) );
  NOR U67267 ( .A(n47029), .B(n47028), .Z(n52499) );
  NOR U67268 ( .A(n50894), .B(n52499), .Z(n47030) );
  XOR U67269 ( .A(n47031), .B(n47030), .Z(n50892) );
  XOR U67270 ( .A(n50889), .B(n50892), .Z(n50888) );
  IV U67271 ( .A(n47032), .Z(n47034) );
  NOR U67272 ( .A(n47034), .B(n47033), .Z(n50886) );
  NOR U67273 ( .A(n50891), .B(n50886), .Z(n47035) );
  XOR U67274 ( .A(n50888), .B(n47035), .Z(n50883) );
  XOR U67275 ( .A(n47036), .B(n50883), .Z(n50875) );
  XOR U67276 ( .A(n47037), .B(n50875), .Z(n47044) );
  IV U67277 ( .A(n47044), .Z(n52510) );
  XOR U67278 ( .A(n47042), .B(n52510), .Z(n47038) );
  NOR U67279 ( .A(n47039), .B(n47038), .Z(n57703) );
  IV U67280 ( .A(n47040), .Z(n47041) );
  NOR U67281 ( .A(n47041), .B(n47046), .Z(n50870) );
  NOR U67282 ( .A(n50870), .B(n47042), .Z(n47043) );
  XOR U67283 ( .A(n47044), .B(n47043), .Z(n52514) );
  IV U67284 ( .A(n47045), .Z(n47047) );
  NOR U67285 ( .A(n47047), .B(n47046), .Z(n47048) );
  IV U67286 ( .A(n47048), .Z(n52513) );
  XOR U67287 ( .A(n52514), .B(n52513), .Z(n47049) );
  NOR U67288 ( .A(n47050), .B(n47049), .Z(n47051) );
  NOR U67289 ( .A(n57703), .B(n47051), .Z(n47059) );
  IV U67290 ( .A(n47059), .Z(n50866) );
  IV U67291 ( .A(n47052), .Z(n47053) );
  NOR U67292 ( .A(n47053), .B(n47068), .Z(n47064) );
  IV U67293 ( .A(n47064), .Z(n47054) );
  NOR U67294 ( .A(n50866), .B(n47054), .Z(n62893) );
  IV U67295 ( .A(n47055), .Z(n47062) );
  IV U67296 ( .A(n47056), .Z(n47057) );
  NOR U67297 ( .A(n47062), .B(n47057), .Z(n47058) );
  IV U67298 ( .A(n47058), .Z(n50865) );
  XOR U67299 ( .A(n47059), .B(n50865), .Z(n50869) );
  IV U67300 ( .A(n47060), .Z(n47061) );
  NOR U67301 ( .A(n47062), .B(n47061), .Z(n50867) );
  XOR U67302 ( .A(n50869), .B(n50867), .Z(n50859) );
  IV U67303 ( .A(n50859), .Z(n47063) );
  NOR U67304 ( .A(n47064), .B(n47063), .Z(n50863) );
  NOR U67305 ( .A(n62893), .B(n50863), .Z(n47071) );
  IV U67306 ( .A(n47065), .Z(n47066) );
  NOR U67307 ( .A(n47074), .B(n47066), .Z(n50858) );
  IV U67308 ( .A(n47067), .Z(n47069) );
  NOR U67309 ( .A(n47069), .B(n47068), .Z(n50862) );
  NOR U67310 ( .A(n50858), .B(n50862), .Z(n47070) );
  XOR U67311 ( .A(n47071), .B(n47070), .Z(n52519) );
  IV U67312 ( .A(n47072), .Z(n47073) );
  NOR U67313 ( .A(n47074), .B(n47073), .Z(n52517) );
  XOR U67314 ( .A(n52519), .B(n52517), .Z(n52522) );
  XOR U67315 ( .A(n52520), .B(n52522), .Z(n50857) );
  XOR U67316 ( .A(n50855), .B(n50857), .Z(n52529) );
  XOR U67317 ( .A(n52530), .B(n52529), .Z(n47081) );
  IV U67318 ( .A(n47081), .Z(n47075) );
  NOR U67319 ( .A(n47076), .B(n47075), .Z(n50850) );
  IV U67320 ( .A(n47077), .Z(n47080) );
  NOR U67321 ( .A(n47079), .B(n50857), .Z(n47078) );
  IV U67322 ( .A(n47078), .Z(n50853) );
  NOR U67323 ( .A(n47080), .B(n50853), .Z(n56022) );
  NOR U67324 ( .A(n47080), .B(n47079), .Z(n47082) );
  NOR U67325 ( .A(n47082), .B(n47081), .Z(n47083) );
  NOR U67326 ( .A(n56022), .B(n47083), .Z(n50842) );
  NOR U67327 ( .A(n47084), .B(n50842), .Z(n47085) );
  NOR U67328 ( .A(n50850), .B(n47085), .Z(n50838) );
  IV U67329 ( .A(n47086), .Z(n50844) );
  NOR U67330 ( .A(n47087), .B(n50844), .Z(n47090) );
  IV U67331 ( .A(n47088), .Z(n47089) );
  NOR U67332 ( .A(n47089), .B(n47093), .Z(n50837) );
  NOR U67333 ( .A(n47090), .B(n50837), .Z(n47091) );
  XOR U67334 ( .A(n50838), .B(n47091), .Z(n50836) );
  IV U67335 ( .A(n47092), .Z(n47094) );
  NOR U67336 ( .A(n47094), .B(n47093), .Z(n50834) );
  XOR U67337 ( .A(n50836), .B(n50834), .Z(n50827) );
  XOR U67338 ( .A(n50826), .B(n50827), .Z(n50832) );
  XOR U67339 ( .A(n47095), .B(n50832), .Z(n47096) );
  IV U67340 ( .A(n47096), .Z(n50824) );
  XOR U67341 ( .A(n50822), .B(n50824), .Z(n52536) );
  XOR U67342 ( .A(n52535), .B(n52536), .Z(n52539) );
  XOR U67343 ( .A(n52538), .B(n52539), .Z(n52543) );
  XOR U67344 ( .A(n52542), .B(n52543), .Z(n52549) );
  IV U67345 ( .A(n47097), .Z(n50817) );
  NOR U67346 ( .A(n47098), .B(n50817), .Z(n47099) );
  NOR U67347 ( .A(n52550), .B(n47099), .Z(n47100) );
  XOR U67348 ( .A(n52549), .B(n47100), .Z(n47101) );
  IV U67349 ( .A(n47101), .Z(n52557) );
  XOR U67350 ( .A(n52556), .B(n52557), .Z(n52560) );
  XOR U67351 ( .A(n47102), .B(n52560), .Z(n50806) );
  XOR U67352 ( .A(n47103), .B(n50806), .Z(n50804) );
  XOR U67353 ( .A(n50801), .B(n50804), .Z(n52566) );
  XOR U67354 ( .A(n47104), .B(n52566), .Z(n47105) );
  IV U67355 ( .A(n47105), .Z(n52570) );
  XOR U67356 ( .A(n52568), .B(n52570), .Z(n52571) );
  XOR U67357 ( .A(n52572), .B(n52571), .Z(n52577) );
  IV U67358 ( .A(n47106), .Z(n47108) );
  IV U67359 ( .A(n47107), .Z(n47111) );
  NOR U67360 ( .A(n47108), .B(n47111), .Z(n52579) );
  NOR U67361 ( .A(n52576), .B(n52579), .Z(n47109) );
  XOR U67362 ( .A(n52577), .B(n47109), .Z(n52575) );
  IV U67363 ( .A(n47110), .Z(n47112) );
  NOR U67364 ( .A(n47112), .B(n47111), .Z(n47113) );
  IV U67365 ( .A(n47113), .Z(n52574) );
  XOR U67366 ( .A(n52575), .B(n52574), .Z(n47122) );
  IV U67367 ( .A(n47122), .Z(n52587) );
  XOR U67368 ( .A(n52584), .B(n52587), .Z(n47119) );
  IV U67369 ( .A(n47114), .Z(n47117) );
  IV U67370 ( .A(n47115), .Z(n47116) );
  NOR U67371 ( .A(n47117), .B(n47116), .Z(n47131) );
  IV U67372 ( .A(n47131), .Z(n47118) );
  NOR U67373 ( .A(n47119), .B(n47118), .Z(n55955) );
  IV U67374 ( .A(n47120), .Z(n47121) );
  NOR U67375 ( .A(n47125), .B(n47121), .Z(n52586) );
  NOR U67376 ( .A(n52586), .B(n52584), .Z(n47123) );
  XOR U67377 ( .A(n47123), .B(n47122), .Z(n50800) );
  IV U67378 ( .A(n47124), .Z(n47128) );
  XOR U67379 ( .A(n47126), .B(n47125), .Z(n47127) );
  NOR U67380 ( .A(n47128), .B(n47127), .Z(n47129) );
  IV U67381 ( .A(n47129), .Z(n50799) );
  XOR U67382 ( .A(n50800), .B(n50799), .Z(n47130) );
  NOR U67383 ( .A(n47131), .B(n47130), .Z(n47132) );
  NOR U67384 ( .A(n55955), .B(n47132), .Z(n50786) );
  XOR U67385 ( .A(n47133), .B(n50786), .Z(n50776) );
  XOR U67386 ( .A(n50774), .B(n50776), .Z(n50770) );
  IV U67387 ( .A(n50770), .Z(n47140) );
  IV U67388 ( .A(n47134), .Z(n47135) );
  NOR U67389 ( .A(n50765), .B(n47135), .Z(n50769) );
  IV U67390 ( .A(n47136), .Z(n47138) );
  NOR U67391 ( .A(n47138), .B(n47137), .Z(n50772) );
  NOR U67392 ( .A(n50769), .B(n50772), .Z(n47139) );
  XOR U67393 ( .A(n47140), .B(n47139), .Z(n50764) );
  XOR U67394 ( .A(n50759), .B(n50764), .Z(n50750) );
  XOR U67395 ( .A(n47141), .B(n50750), .Z(n50743) );
  XOR U67396 ( .A(n47142), .B(n50743), .Z(n50742) );
  XOR U67397 ( .A(n50740), .B(n50742), .Z(n57803) );
  XOR U67398 ( .A(n47143), .B(n57803), .Z(n52597) );
  XOR U67399 ( .A(n52595), .B(n52597), .Z(n50734) );
  NOR U67400 ( .A(n47144), .B(n52598), .Z(n47148) );
  IV U67401 ( .A(n47145), .Z(n47147) );
  IV U67402 ( .A(n47146), .Z(n47150) );
  NOR U67403 ( .A(n47147), .B(n47150), .Z(n50733) );
  NOR U67404 ( .A(n47148), .B(n50733), .Z(n47149) );
  XOR U67405 ( .A(n50734), .B(n47149), .Z(n52611) );
  IV U67406 ( .A(n52616), .Z(n47151) );
  NOR U67407 ( .A(n47151), .B(n47150), .Z(n50731) );
  IV U67408 ( .A(n47152), .Z(n47154) );
  NOR U67409 ( .A(n47154), .B(n47153), .Z(n47155) );
  NOR U67410 ( .A(n50731), .B(n47155), .Z(n52612) );
  XOR U67411 ( .A(n52611), .B(n52612), .Z(n52609) );
  XOR U67412 ( .A(n52608), .B(n52609), .Z(n55908) );
  IV U67413 ( .A(n47156), .Z(n47158) );
  NOR U67414 ( .A(n47158), .B(n47157), .Z(n55907) );
  NOR U67415 ( .A(n55913), .B(n55907), .Z(n52622) );
  XOR U67416 ( .A(n55908), .B(n52622), .Z(n47159) );
  IV U67417 ( .A(n47159), .Z(n52619) );
  XOR U67418 ( .A(n52618), .B(n52619), .Z(n52625) );
  XOR U67419 ( .A(n52624), .B(n52625), .Z(n50727) );
  XOR U67420 ( .A(n47160), .B(n50727), .Z(n47161) );
  IV U67421 ( .A(n47161), .Z(n50724) );
  IV U67422 ( .A(n47162), .Z(n47165) );
  IV U67423 ( .A(n47163), .Z(n47164) );
  NOR U67424 ( .A(n47165), .B(n47164), .Z(n50722) );
  XOR U67425 ( .A(n50724), .B(n50722), .Z(n50715) );
  XOR U67426 ( .A(n50714), .B(n50715), .Z(n50718) );
  XOR U67427 ( .A(n50717), .B(n50718), .Z(n50708) );
  XOR U67428 ( .A(n50707), .B(n50708), .Z(n50712) );
  XOR U67429 ( .A(n50703), .B(n50712), .Z(n50701) );
  XOR U67430 ( .A(n50702), .B(n50701), .Z(n50697) );
  XOR U67431 ( .A(n50696), .B(n50697), .Z(n50699) );
  XOR U67432 ( .A(n50700), .B(n50699), .Z(n47172) );
  IV U67433 ( .A(n47172), .Z(n52638) );
  XOR U67434 ( .A(n50694), .B(n52638), .Z(n47166) );
  NOR U67435 ( .A(n47167), .B(n47166), .Z(n55873) );
  IV U67436 ( .A(n47168), .Z(n50693) );
  IV U67437 ( .A(n47169), .Z(n47170) );
  NOR U67438 ( .A(n47171), .B(n47170), .Z(n52637) );
  NOR U67439 ( .A(n50694), .B(n52637), .Z(n47173) );
  XOR U67440 ( .A(n47173), .B(n47172), .Z(n55860) );
  XOR U67441 ( .A(n50693), .B(n55860), .Z(n47174) );
  NOR U67442 ( .A(n47175), .B(n47174), .Z(n47176) );
  NOR U67443 ( .A(n55873), .B(n47176), .Z(n47177) );
  IV U67444 ( .A(n47177), .Z(n50689) );
  XOR U67445 ( .A(n47178), .B(n50689), .Z(n47185) );
  IV U67446 ( .A(n47179), .Z(n47180) );
  NOR U67447 ( .A(n47188), .B(n47180), .Z(n50683) );
  IV U67448 ( .A(n47181), .Z(n47183) );
  NOR U67449 ( .A(n47183), .B(n47182), .Z(n50686) );
  NOR U67450 ( .A(n50683), .B(n50686), .Z(n47184) );
  XOR U67451 ( .A(n47185), .B(n47184), .Z(n50682) );
  IV U67452 ( .A(n47186), .Z(n47187) );
  NOR U67453 ( .A(n47188), .B(n47187), .Z(n50680) );
  XOR U67454 ( .A(n50682), .B(n50680), .Z(n50675) );
  XOR U67455 ( .A(n50674), .B(n50675), .Z(n50679) );
  IV U67456 ( .A(n47189), .Z(n47197) );
  IV U67457 ( .A(n47190), .Z(n47191) );
  NOR U67458 ( .A(n47197), .B(n47191), .Z(n47192) );
  IV U67459 ( .A(n47192), .Z(n47198) );
  NOR U67460 ( .A(n50679), .B(n47198), .Z(n57840) );
  IV U67461 ( .A(n47193), .Z(n47194) );
  NOR U67462 ( .A(n47194), .B(n47205), .Z(n52659) );
  IV U67463 ( .A(n47195), .Z(n47196) );
  NOR U67464 ( .A(n47197), .B(n47196), .Z(n50677) );
  XOR U67465 ( .A(n50679), .B(n50677), .Z(n52660) );
  IV U67466 ( .A(n52660), .Z(n47199) );
  XOR U67467 ( .A(n52659), .B(n47199), .Z(n47201) );
  NOR U67468 ( .A(n47199), .B(n47198), .Z(n47200) );
  NOR U67469 ( .A(n47201), .B(n47200), .Z(n47202) );
  NOR U67470 ( .A(n57840), .B(n47202), .Z(n47203) );
  IV U67471 ( .A(n47203), .Z(n50672) );
  IV U67472 ( .A(n47204), .Z(n47206) );
  NOR U67473 ( .A(n47206), .B(n47205), .Z(n50670) );
  XOR U67474 ( .A(n50672), .B(n50670), .Z(n52658) );
  IV U67475 ( .A(n47207), .Z(n47209) );
  NOR U67476 ( .A(n47209), .B(n47208), .Z(n52656) );
  XOR U67477 ( .A(n52658), .B(n52656), .Z(n52668) );
  XOR U67478 ( .A(n52667), .B(n52668), .Z(n52671) );
  XOR U67479 ( .A(n52670), .B(n52671), .Z(n50668) );
  XOR U67480 ( .A(n50667), .B(n50668), .Z(n50663) );
  XOR U67481 ( .A(n50662), .B(n50663), .Z(n55825) );
  IV U67482 ( .A(n47210), .Z(n47211) );
  NOR U67483 ( .A(n47212), .B(n47211), .Z(n52676) );
  IV U67484 ( .A(n47213), .Z(n47215) );
  NOR U67485 ( .A(n47215), .B(n47214), .Z(n50665) );
  NOR U67486 ( .A(n52676), .B(n50665), .Z(n47216) );
  XOR U67487 ( .A(n55825), .B(n47216), .Z(n50656) );
  XOR U67488 ( .A(n47217), .B(n50656), .Z(n50651) );
  XOR U67489 ( .A(n50650), .B(n50651), .Z(n63050) );
  XOR U67490 ( .A(n50653), .B(n63050), .Z(n52685) );
  XOR U67491 ( .A(n47218), .B(n52685), .Z(n47219) );
  IV U67492 ( .A(n47219), .Z(n50646) );
  XOR U67493 ( .A(n47220), .B(n50646), .Z(n47231) );
  IV U67494 ( .A(n47231), .Z(n47225) );
  IV U67495 ( .A(n47221), .Z(n47223) );
  IV U67496 ( .A(n47222), .Z(n47227) );
  NOR U67497 ( .A(n47223), .B(n47227), .Z(n47234) );
  IV U67498 ( .A(n47234), .Z(n47224) );
  NOR U67499 ( .A(n47225), .B(n47224), .Z(n50641) );
  XOR U67500 ( .A(n50644), .B(n50646), .Z(n50648) );
  IV U67501 ( .A(n47226), .Z(n47228) );
  NOR U67502 ( .A(n47228), .B(n47227), .Z(n47230) );
  IV U67503 ( .A(n47230), .Z(n47229) );
  NOR U67504 ( .A(n50648), .B(n47229), .Z(n55801) );
  NOR U67505 ( .A(n47231), .B(n47230), .Z(n47232) );
  NOR U67506 ( .A(n55801), .B(n47232), .Z(n47233) );
  NOR U67507 ( .A(n47234), .B(n47233), .Z(n47235) );
  NOR U67508 ( .A(n50641), .B(n47235), .Z(n50635) );
  IV U67509 ( .A(n47236), .Z(n47237) );
  NOR U67510 ( .A(n47240), .B(n47237), .Z(n55796) );
  IV U67511 ( .A(n47238), .Z(n47239) );
  NOR U67512 ( .A(n47240), .B(n47239), .Z(n57854) );
  NOR U67513 ( .A(n55796), .B(n57854), .Z(n50636) );
  XOR U67514 ( .A(n50635), .B(n50636), .Z(n50638) );
  XOR U67515 ( .A(n50637), .B(n50638), .Z(n50630) );
  XOR U67516 ( .A(n47241), .B(n50630), .Z(n52692) );
  XOR U67517 ( .A(n52693), .B(n52692), .Z(n52698) );
  IV U67518 ( .A(n47242), .Z(n47244) );
  NOR U67519 ( .A(n47244), .B(n47243), .Z(n47245) );
  IV U67520 ( .A(n47245), .Z(n52695) );
  XOR U67521 ( .A(n52698), .B(n52695), .Z(n50618) );
  IV U67522 ( .A(n47246), .Z(n47248) );
  NOR U67523 ( .A(n47248), .B(n47247), .Z(n52697) );
  NOR U67524 ( .A(n47249), .B(n50620), .Z(n47250) );
  NOR U67525 ( .A(n52697), .B(n47250), .Z(n47251) );
  XOR U67526 ( .A(n50618), .B(n47251), .Z(n52703) );
  XOR U67527 ( .A(n52701), .B(n52703), .Z(n50615) );
  XOR U67528 ( .A(n47252), .B(n50615), .Z(n47253) );
  IV U67529 ( .A(n47253), .Z(n50611) );
  XOR U67530 ( .A(n50609), .B(n50611), .Z(n52714) );
  XOR U67531 ( .A(n50604), .B(n52714), .Z(n50606) );
  XOR U67532 ( .A(n50607), .B(n50606), .Z(n50601) );
  NOR U67533 ( .A(n52717), .B(n52715), .Z(n47256) );
  IV U67534 ( .A(n47254), .Z(n47259) );
  NOR U67535 ( .A(n47255), .B(n47259), .Z(n50600) );
  NOR U67536 ( .A(n47256), .B(n50600), .Z(n47257) );
  XOR U67537 ( .A(n50601), .B(n47257), .Z(n50599) );
  IV U67538 ( .A(n47258), .Z(n47260) );
  NOR U67539 ( .A(n47260), .B(n47259), .Z(n50597) );
  XOR U67540 ( .A(n50599), .B(n50597), .Z(n50596) );
  XOR U67541 ( .A(n47261), .B(n50596), .Z(n52721) );
  XOR U67542 ( .A(n52723), .B(n52721), .Z(n52727) );
  IV U67543 ( .A(n47262), .Z(n47264) );
  NOR U67544 ( .A(n47264), .B(n47263), .Z(n52724) );
  XOR U67545 ( .A(n52727), .B(n52724), .Z(n50589) );
  IV U67546 ( .A(n47265), .Z(n52728) );
  NOR U67547 ( .A(n52728), .B(n52730), .Z(n47269) );
  IV U67548 ( .A(n47266), .Z(n47268) );
  NOR U67549 ( .A(n47268), .B(n47267), .Z(n50588) );
  NOR U67550 ( .A(n47269), .B(n50588), .Z(n47270) );
  XOR U67551 ( .A(n50589), .B(n47270), .Z(n47271) );
  IV U67552 ( .A(n47271), .Z(n50584) );
  XOR U67553 ( .A(n50582), .B(n50584), .Z(n50587) );
  XOR U67554 ( .A(n50585), .B(n50587), .Z(n52733) );
  XOR U67555 ( .A(n52734), .B(n52733), .Z(n47272) );
  IV U67556 ( .A(n47272), .Z(n52739) );
  XOR U67557 ( .A(n52738), .B(n52739), .Z(n52747) );
  IV U67558 ( .A(n52747), .Z(n47277) );
  IV U67559 ( .A(n47273), .Z(n47285) );
  IV U67560 ( .A(n47284), .Z(n47275) );
  NOR U67561 ( .A(n47285), .B(n47275), .Z(n52741) );
  IV U67562 ( .A(n47274), .Z(n47276) );
  NOR U67563 ( .A(n47276), .B(n47275), .Z(n52744) );
  NOR U67564 ( .A(n52741), .B(n52744), .Z(n47288) );
  XOR U67565 ( .A(n47277), .B(n47288), .Z(n47282) );
  IV U67566 ( .A(n47278), .Z(n47280) );
  NOR U67567 ( .A(n47280), .B(n47279), .Z(n47291) );
  IV U67568 ( .A(n47291), .Z(n47281) );
  NOR U67569 ( .A(n47282), .B(n47281), .Z(n55741) );
  IV U67570 ( .A(n47283), .Z(n47287) );
  XOR U67571 ( .A(n47285), .B(n47284), .Z(n47286) );
  NOR U67572 ( .A(n47287), .B(n47286), .Z(n52746) );
  IV U67573 ( .A(n47288), .Z(n47289) );
  NOR U67574 ( .A(n52746), .B(n47289), .Z(n47290) );
  XOR U67575 ( .A(n47290), .B(n52747), .Z(n47292) );
  NOR U67576 ( .A(n47292), .B(n47291), .Z(n47293) );
  NOR U67577 ( .A(n55741), .B(n47293), .Z(n52750) );
  XOR U67578 ( .A(n52751), .B(n52750), .Z(n52755) );
  XOR U67579 ( .A(n47294), .B(n52755), .Z(n50576) );
  XOR U67580 ( .A(n50577), .B(n50576), .Z(n52766) );
  XOR U67581 ( .A(n52765), .B(n52766), .Z(n52768) );
  XOR U67582 ( .A(n52769), .B(n52768), .Z(n47295) );
  NOR U67583 ( .A(n47296), .B(n47295), .Z(n52773) );
  IV U67584 ( .A(n47296), .Z(n47301) );
  XOR U67585 ( .A(n47298), .B(n47297), .Z(n47299) );
  NOR U67586 ( .A(n47299), .B(n52768), .Z(n47300) );
  IV U67587 ( .A(n47300), .Z(n55724) );
  NOR U67588 ( .A(n47301), .B(n55724), .Z(n47302) );
  NOR U67589 ( .A(n52773), .B(n47302), .Z(n47303) );
  IV U67590 ( .A(n47303), .Z(n47311) );
  NOR U67591 ( .A(n47304), .B(n47311), .Z(n55722) );
  IV U67592 ( .A(n47305), .Z(n47307) );
  IV U67593 ( .A(n47306), .Z(n47309) );
  NOR U67594 ( .A(n47307), .B(n47309), .Z(n57933) );
  IV U67595 ( .A(n47308), .Z(n55726) );
  NOR U67596 ( .A(n47309), .B(n55726), .Z(n47310) );
  XOR U67597 ( .A(n47311), .B(n47310), .Z(n57934) );
  XOR U67598 ( .A(n57933), .B(n57934), .Z(n47316) );
  IV U67599 ( .A(n47316), .Z(n52772) );
  NOR U67600 ( .A(n47312), .B(n52772), .Z(n47313) );
  NOR U67601 ( .A(n55722), .B(n47313), .Z(n52779) );
  XOR U67602 ( .A(n52778), .B(n52779), .Z(n47314) );
  NOR U67603 ( .A(n47315), .B(n47314), .Z(n47318) );
  IV U67604 ( .A(n47315), .Z(n47317) );
  NOR U67605 ( .A(n47317), .B(n47316), .Z(n52777) );
  NOR U67606 ( .A(n47318), .B(n52777), .Z(n50574) );
  IV U67607 ( .A(n47319), .Z(n47320) );
  NOR U67608 ( .A(n47321), .B(n47320), .Z(n52787) );
  IV U67609 ( .A(n47322), .Z(n47324) );
  NOR U67610 ( .A(n47324), .B(n47323), .Z(n47327) );
  NOR U67611 ( .A(n52787), .B(n47327), .Z(n47325) );
  XOR U67612 ( .A(n50574), .B(n47325), .Z(n52791) );
  XOR U67613 ( .A(n52790), .B(n52791), .Z(n47326) );
  NOR U67614 ( .A(n47328), .B(n47326), .Z(n47332) );
  IV U67615 ( .A(n47327), .Z(n50575) );
  XOR U67616 ( .A(n50574), .B(n50575), .Z(n50567) );
  IV U67617 ( .A(n50567), .Z(n47330) );
  IV U67618 ( .A(n47328), .Z(n47329) );
  NOR U67619 ( .A(n47330), .B(n47329), .Z(n47331) );
  NOR U67620 ( .A(n47332), .B(n47331), .Z(n50565) );
  XOR U67621 ( .A(n50563), .B(n50565), .Z(n52797) );
  IV U67622 ( .A(n47333), .Z(n47335) );
  NOR U67623 ( .A(n47335), .B(n47334), .Z(n47336) );
  IV U67624 ( .A(n47336), .Z(n52795) );
  XOR U67625 ( .A(n52797), .B(n52795), .Z(n47337) );
  XOR U67626 ( .A(n47338), .B(n47337), .Z(n50560) );
  XOR U67627 ( .A(n50558), .B(n50560), .Z(n50557) );
  IV U67628 ( .A(n47339), .Z(n47340) );
  NOR U67629 ( .A(n47341), .B(n47340), .Z(n50553) );
  IV U67630 ( .A(n47342), .Z(n47345) );
  IV U67631 ( .A(n47343), .Z(n47344) );
  NOR U67632 ( .A(n47345), .B(n47344), .Z(n50555) );
  NOR U67633 ( .A(n50553), .B(n50555), .Z(n47346) );
  XOR U67634 ( .A(n50557), .B(n47346), .Z(n50547) );
  IV U67635 ( .A(n47347), .Z(n47349) );
  NOR U67636 ( .A(n47349), .B(n47348), .Z(n47350) );
  IV U67637 ( .A(n47350), .Z(n50548) );
  XOR U67638 ( .A(n50547), .B(n50548), .Z(n47351) );
  XOR U67639 ( .A(n47352), .B(n47351), .Z(n50541) );
  XOR U67640 ( .A(n47353), .B(n50541), .Z(n50540) );
  XOR U67641 ( .A(n50538), .B(n50540), .Z(n52810) );
  XOR U67642 ( .A(n47354), .B(n52810), .Z(n50526) );
  IV U67643 ( .A(n47355), .Z(n50530) );
  NOR U67644 ( .A(n50533), .B(n50530), .Z(n47359) );
  IV U67645 ( .A(n47356), .Z(n47358) );
  NOR U67646 ( .A(n47358), .B(n47357), .Z(n50525) );
  NOR U67647 ( .A(n47359), .B(n50525), .Z(n47360) );
  XOR U67648 ( .A(n50526), .B(n47360), .Z(n50524) );
  XOR U67649 ( .A(n50522), .B(n50524), .Z(n52822) );
  XOR U67650 ( .A(n52823), .B(n52822), .Z(n47364) );
  IV U67651 ( .A(n47364), .Z(n55670) );
  XOR U67652 ( .A(n52824), .B(n55670), .Z(n50517) );
  NOR U67653 ( .A(n47361), .B(n50517), .Z(n57999) );
  IV U67654 ( .A(n47362), .Z(n47363) );
  NOR U67655 ( .A(n47368), .B(n47363), .Z(n50518) );
  NOR U67656 ( .A(n50518), .B(n52824), .Z(n47365) );
  XOR U67657 ( .A(n47365), .B(n47364), .Z(n50520) );
  IV U67658 ( .A(n47366), .Z(n47367) );
  NOR U67659 ( .A(n47368), .B(n47367), .Z(n47369) );
  IV U67660 ( .A(n47369), .Z(n55667) );
  XOR U67661 ( .A(n50520), .B(n55667), .Z(n47370) );
  NOR U67662 ( .A(n47371), .B(n47370), .Z(n47372) );
  NOR U67663 ( .A(n57999), .B(n47372), .Z(n50509) );
  XOR U67664 ( .A(n47373), .B(n50509), .Z(n50504) );
  XOR U67665 ( .A(n47374), .B(n50504), .Z(n50494) );
  XOR U67666 ( .A(n47375), .B(n50494), .Z(n47380) );
  IV U67667 ( .A(n47380), .Z(n50490) );
  XOR U67668 ( .A(n50489), .B(n50490), .Z(n47376) );
  NOR U67669 ( .A(n47377), .B(n47376), .Z(n55649) );
  IV U67670 ( .A(n47378), .Z(n47379) );
  NOR U67671 ( .A(n47379), .B(n47383), .Z(n50487) );
  NOR U67672 ( .A(n50489), .B(n50487), .Z(n47381) );
  XOR U67673 ( .A(n47381), .B(n47380), .Z(n50486) );
  IV U67674 ( .A(n47382), .Z(n47384) );
  NOR U67675 ( .A(n47384), .B(n47383), .Z(n47385) );
  IV U67676 ( .A(n47385), .Z(n50485) );
  XOR U67677 ( .A(n50486), .B(n50485), .Z(n47386) );
  NOR U67678 ( .A(n47387), .B(n47386), .Z(n47388) );
  NOR U67679 ( .A(n55649), .B(n47388), .Z(n47389) );
  IV U67680 ( .A(n47389), .Z(n50483) );
  XOR U67681 ( .A(n50482), .B(n50483), .Z(n52843) );
  IV U67682 ( .A(n47390), .Z(n47391) );
  NOR U67683 ( .A(n47392), .B(n47391), .Z(n52841) );
  XOR U67684 ( .A(n52843), .B(n52841), .Z(n50480) );
  XOR U67685 ( .A(n50479), .B(n50480), .Z(n50478) );
  IV U67686 ( .A(n47393), .Z(n47394) );
  NOR U67687 ( .A(n47395), .B(n47394), .Z(n50476) );
  XOR U67688 ( .A(n50478), .B(n50476), .Z(n47396) );
  XOR U67689 ( .A(n47397), .B(n47396), .Z(n50460) );
  IV U67690 ( .A(n47398), .Z(n50464) );
  NOR U67691 ( .A(n47399), .B(n50464), .Z(n47403) );
  IV U67692 ( .A(n47400), .Z(n47402) );
  NOR U67693 ( .A(n47402), .B(n47401), .Z(n50461) );
  NOR U67694 ( .A(n47403), .B(n50461), .Z(n47404) );
  XOR U67695 ( .A(n50460), .B(n47404), .Z(n52861) );
  XOR U67696 ( .A(n52860), .B(n52861), .Z(n52864) );
  NOR U67697 ( .A(n50458), .B(n52863), .Z(n47405) );
  XOR U67698 ( .A(n52864), .B(n47405), .Z(n47406) );
  IV U67699 ( .A(n47406), .Z(n50457) );
  XOR U67700 ( .A(n50455), .B(n50457), .Z(n50451) );
  XOR U67701 ( .A(n50450), .B(n50451), .Z(n52870) );
  XOR U67702 ( .A(n47407), .B(n52870), .Z(n52872) );
  IV U67703 ( .A(n47408), .Z(n47409) );
  NOR U67704 ( .A(n47409), .B(n47411), .Z(n52871) );
  IV U67705 ( .A(n47410), .Z(n47412) );
  NOR U67706 ( .A(n47412), .B(n47411), .Z(n52877) );
  NOR U67707 ( .A(n52871), .B(n52877), .Z(n47413) );
  XOR U67708 ( .A(n52872), .B(n47413), .Z(n50449) );
  IV U67709 ( .A(n47414), .Z(n47416) );
  NOR U67710 ( .A(n47416), .B(n47415), .Z(n50447) );
  XOR U67711 ( .A(n50449), .B(n50447), .Z(n52889) );
  XOR U67712 ( .A(n47417), .B(n52889), .Z(n47418) );
  IV U67713 ( .A(n47418), .Z(n50440) );
  XOR U67714 ( .A(n50439), .B(n50440), .Z(n50426) );
  IV U67715 ( .A(n47422), .Z(n50433) );
  NOR U67716 ( .A(n47420), .B(n50433), .Z(n47425) );
  IV U67717 ( .A(n47419), .Z(n55615) );
  IV U67718 ( .A(n47420), .Z(n47421) );
  NOR U67719 ( .A(n47422), .B(n47421), .Z(n47423) );
  NOR U67720 ( .A(n55615), .B(n47423), .Z(n47424) );
  NOR U67721 ( .A(n47425), .B(n47424), .Z(n47426) );
  XOR U67722 ( .A(n50426), .B(n47426), .Z(n50421) );
  IV U67723 ( .A(n47427), .Z(n50423) );
  NOR U67724 ( .A(n50423), .B(n50425), .Z(n47430) );
  IV U67725 ( .A(n47428), .Z(n55610) );
  NOR U67726 ( .A(n50427), .B(n55610), .Z(n47429) );
  NOR U67727 ( .A(n47430), .B(n47429), .Z(n47431) );
  XOR U67728 ( .A(n50421), .B(n47431), .Z(n55593) );
  IV U67729 ( .A(n47432), .Z(n50414) );
  NOR U67730 ( .A(n47433), .B(n50414), .Z(n47440) );
  IV U67731 ( .A(n47434), .Z(n47435) );
  NOR U67732 ( .A(n47435), .B(n47437), .Z(n55596) );
  IV U67733 ( .A(n47436), .Z(n47438) );
  NOR U67734 ( .A(n47438), .B(n47437), .Z(n55591) );
  NOR U67735 ( .A(n55596), .B(n55591), .Z(n50420) );
  IV U67736 ( .A(n50420), .Z(n47439) );
  NOR U67737 ( .A(n47440), .B(n47439), .Z(n47441) );
  XOR U67738 ( .A(n55593), .B(n47441), .Z(n52901) );
  IV U67739 ( .A(n52901), .Z(n52909) );
  IV U67740 ( .A(n47442), .Z(n47444) );
  IV U67741 ( .A(n47443), .Z(n47445) );
  NOR U67742 ( .A(n47444), .B(n47445), .Z(n52905) );
  NOR U67743 ( .A(n50412), .B(n50410), .Z(n47447) );
  NOR U67744 ( .A(n47446), .B(n47445), .Z(n52907) );
  NOR U67745 ( .A(n47447), .B(n52907), .Z(n52902) );
  IV U67746 ( .A(n52902), .Z(n47448) );
  NOR U67747 ( .A(n52905), .B(n47448), .Z(n47449) );
  XOR U67748 ( .A(n52909), .B(n47449), .Z(n52914) );
  NOR U67749 ( .A(n52916), .B(n47450), .Z(n47454) );
  IV U67750 ( .A(n47451), .Z(n47453) );
  NOR U67751 ( .A(n47453), .B(n47452), .Z(n52900) );
  NOR U67752 ( .A(n47454), .B(n52900), .Z(n47455) );
  XOR U67753 ( .A(n52914), .B(n47455), .Z(n52931) );
  IV U67754 ( .A(n47456), .Z(n47461) );
  XOR U67755 ( .A(n47465), .B(n47463), .Z(n47459) );
  IV U67756 ( .A(n47457), .Z(n47464) );
  NOR U67757 ( .A(n47463), .B(n47464), .Z(n47458) );
  NOR U67758 ( .A(n47459), .B(n47458), .Z(n47460) );
  NOR U67759 ( .A(n47461), .B(n47460), .Z(n47462) );
  IV U67760 ( .A(n47462), .Z(n47468) );
  NOR U67761 ( .A(n52931), .B(n47468), .Z(n55564) );
  IV U67762 ( .A(n47463), .Z(n47466) );
  NOR U67763 ( .A(n47464), .B(n47466), .Z(n52925) );
  IV U67764 ( .A(n47465), .Z(n47467) );
  NOR U67765 ( .A(n47467), .B(n47466), .Z(n52923) );
  XOR U67766 ( .A(n52923), .B(n52931), .Z(n52926) );
  IV U67767 ( .A(n52926), .Z(n47469) );
  XOR U67768 ( .A(n52925), .B(n47469), .Z(n47471) );
  NOR U67769 ( .A(n47469), .B(n47468), .Z(n47470) );
  NOR U67770 ( .A(n47471), .B(n47470), .Z(n47472) );
  NOR U67771 ( .A(n55564), .B(n47472), .Z(n47473) );
  IV U67772 ( .A(n47473), .Z(n52935) );
  IV U67773 ( .A(n47474), .Z(n47475) );
  NOR U67774 ( .A(n47484), .B(n47475), .Z(n50405) );
  IV U67775 ( .A(n47476), .Z(n47478) );
  NOR U67776 ( .A(n47478), .B(n47477), .Z(n52929) );
  IV U67777 ( .A(n47479), .Z(n47480) );
  NOR U67778 ( .A(n47481), .B(n47480), .Z(n47482) );
  IV U67779 ( .A(n47482), .Z(n47483) );
  NOR U67780 ( .A(n47484), .B(n47483), .Z(n52933) );
  NOR U67781 ( .A(n52929), .B(n52933), .Z(n47485) );
  IV U67782 ( .A(n47485), .Z(n50406) );
  NOR U67783 ( .A(n50405), .B(n50406), .Z(n47486) );
  XOR U67784 ( .A(n52935), .B(n47486), .Z(n50397) );
  IV U67785 ( .A(n47487), .Z(n47489) );
  IV U67786 ( .A(n47488), .Z(n47498) );
  NOR U67787 ( .A(n47489), .B(n47498), .Z(n50402) );
  IV U67788 ( .A(n47490), .Z(n47491) );
  NOR U67789 ( .A(n47491), .B(n47493), .Z(n47503) );
  IV U67790 ( .A(n47492), .Z(n47494) );
  NOR U67791 ( .A(n47494), .B(n47493), .Z(n50399) );
  XOR U67792 ( .A(n47503), .B(n50399), .Z(n47495) );
  NOR U67793 ( .A(n50402), .B(n47495), .Z(n47496) );
  XOR U67794 ( .A(n50397), .B(n47496), .Z(n52939) );
  IV U67795 ( .A(n47497), .Z(n47499) );
  NOR U67796 ( .A(n47499), .B(n47498), .Z(n47500) );
  IV U67797 ( .A(n47500), .Z(n52938) );
  XOR U67798 ( .A(n52939), .B(n52938), .Z(n47501) );
  NOR U67799 ( .A(n47502), .B(n47501), .Z(n47506) );
  IV U67800 ( .A(n47502), .Z(n47505) );
  IV U67801 ( .A(n47503), .Z(n50398) );
  XOR U67802 ( .A(n50398), .B(n50397), .Z(n50400) );
  XOR U67803 ( .A(n50399), .B(n50400), .Z(n47504) );
  NOR U67804 ( .A(n47505), .B(n47504), .Z(n55550) );
  NOR U67805 ( .A(n47506), .B(n55550), .Z(n50393) );
  XOR U67806 ( .A(n52942), .B(n50393), .Z(n50385) );
  XOR U67807 ( .A(n47507), .B(n50385), .Z(n50377) );
  NOR U67808 ( .A(n47508), .B(n50386), .Z(n47512) );
  IV U67809 ( .A(n47509), .Z(n50378) );
  NOR U67810 ( .A(n47510), .B(n50378), .Z(n47511) );
  NOR U67811 ( .A(n47512), .B(n47511), .Z(n47513) );
  XOR U67812 ( .A(n50377), .B(n47513), .Z(n50360) );
  XOR U67813 ( .A(n50367), .B(n50360), .Z(n50352) );
  XOR U67814 ( .A(n47514), .B(n50352), .Z(n50346) );
  XOR U67815 ( .A(n50347), .B(n50346), .Z(n50349) );
  IV U67816 ( .A(n47515), .Z(n47517) );
  NOR U67817 ( .A(n47517), .B(n47516), .Z(n50348) );
  NOR U67818 ( .A(n50348), .B(n52951), .Z(n47518) );
  XOR U67819 ( .A(n50349), .B(n47518), .Z(n47519) );
  IV U67820 ( .A(n47519), .Z(n52957) );
  XOR U67821 ( .A(n52955), .B(n52957), .Z(n52959) );
  XOR U67822 ( .A(n52958), .B(n52959), .Z(n50344) );
  XOR U67823 ( .A(n50343), .B(n50344), .Z(n47528) );
  IV U67824 ( .A(n47528), .Z(n50338) );
  XOR U67825 ( .A(n50333), .B(n50338), .Z(n47520) );
  NOR U67826 ( .A(n47521), .B(n47520), .Z(n58131) );
  IV U67827 ( .A(n47522), .Z(n47523) );
  NOR U67828 ( .A(n47523), .B(n47526), .Z(n47524) );
  IV U67829 ( .A(n47524), .Z(n50332) );
  IV U67830 ( .A(n47525), .Z(n47527) );
  NOR U67831 ( .A(n47527), .B(n47526), .Z(n50329) );
  NOR U67832 ( .A(n50333), .B(n50329), .Z(n47529) );
  XOR U67833 ( .A(n47529), .B(n47528), .Z(n50331) );
  XOR U67834 ( .A(n50332), .B(n50331), .Z(n47530) );
  NOR U67835 ( .A(n47531), .B(n47530), .Z(n47532) );
  NOR U67836 ( .A(n58131), .B(n47532), .Z(n50324) );
  IV U67837 ( .A(n47533), .Z(n47534) );
  NOR U67838 ( .A(n47537), .B(n47534), .Z(n50326) );
  IV U67839 ( .A(n47535), .Z(n47536) );
  NOR U67840 ( .A(n47537), .B(n47536), .Z(n50323) );
  NOR U67841 ( .A(n50326), .B(n50323), .Z(n47538) );
  XOR U67842 ( .A(n50324), .B(n47538), .Z(n50313) );
  XOR U67843 ( .A(n50312), .B(n50313), .Z(n50316) );
  XOR U67844 ( .A(n50315), .B(n50316), .Z(n50319) );
  XOR U67845 ( .A(n50318), .B(n50319), .Z(n50308) );
  XOR U67846 ( .A(n50306), .B(n50308), .Z(n50311) );
  XOR U67847 ( .A(n47539), .B(n50311), .Z(n47540) );
  IV U67848 ( .A(n47540), .Z(n50301) );
  XOR U67849 ( .A(n50300), .B(n50301), .Z(n52969) );
  IV U67850 ( .A(n47541), .Z(n47542) );
  NOR U67851 ( .A(n47545), .B(n47542), .Z(n52967) );
  XOR U67852 ( .A(n52969), .B(n52967), .Z(n52972) );
  IV U67853 ( .A(n47543), .Z(n47544) );
  NOR U67854 ( .A(n47545), .B(n47544), .Z(n52970) );
  XOR U67855 ( .A(n52972), .B(n52970), .Z(n50292) );
  IV U67856 ( .A(n47546), .Z(n47547) );
  NOR U67857 ( .A(n47547), .B(n47551), .Z(n50291) );
  IV U67858 ( .A(n47548), .Z(n50295) );
  NOR U67859 ( .A(n47549), .B(n50295), .Z(n47553) );
  IV U67860 ( .A(n47550), .Z(n47552) );
  NOR U67861 ( .A(n47552), .B(n47551), .Z(n50289) );
  NOR U67862 ( .A(n47553), .B(n50289), .Z(n47554) );
  IV U67863 ( .A(n47554), .Z(n47555) );
  NOR U67864 ( .A(n50291), .B(n47555), .Z(n47556) );
  XOR U67865 ( .A(n50292), .B(n47556), .Z(n47557) );
  IV U67866 ( .A(n47557), .Z(n52979) );
  XOR U67867 ( .A(n52977), .B(n52979), .Z(n52982) );
  XOR U67868 ( .A(n52980), .B(n52982), .Z(n50288) );
  XOR U67869 ( .A(n47558), .B(n50288), .Z(n50273) );
  XOR U67870 ( .A(n47559), .B(n50273), .Z(n52987) );
  XOR U67871 ( .A(n47560), .B(n52987), .Z(n47577) );
  NOR U67872 ( .A(n47561), .B(n50261), .Z(n47562) );
  NOR U67873 ( .A(n47577), .B(n47562), .Z(n47565) );
  IV U67874 ( .A(n47562), .Z(n47563) );
  XOR U67875 ( .A(n50270), .B(n52987), .Z(n50260) );
  NOR U67876 ( .A(n47563), .B(n50260), .Z(n47564) );
  NOR U67877 ( .A(n47565), .B(n47564), .Z(n47580) );
  IV U67878 ( .A(n47580), .Z(n47570) );
  IV U67879 ( .A(n47566), .Z(n47568) );
  NOR U67880 ( .A(n47568), .B(n47567), .Z(n47584) );
  IV U67881 ( .A(n47584), .Z(n47569) );
  NOR U67882 ( .A(n47570), .B(n47569), .Z(n58179) );
  IV U67883 ( .A(n47571), .Z(n47573) );
  IV U67884 ( .A(n47572), .Z(n47575) );
  NOR U67885 ( .A(n47573), .B(n47575), .Z(n50255) );
  IV U67886 ( .A(n47574), .Z(n47576) );
  NOR U67887 ( .A(n47576), .B(n47575), .Z(n47581) );
  IV U67888 ( .A(n47581), .Z(n47579) );
  IV U67889 ( .A(n47577), .Z(n47578) );
  NOR U67890 ( .A(n47579), .B(n47578), .Z(n58169) );
  NOR U67891 ( .A(n47581), .B(n47580), .Z(n47582) );
  NOR U67892 ( .A(n58169), .B(n47582), .Z(n50256) );
  XOR U67893 ( .A(n50255), .B(n50256), .Z(n47583) );
  NOR U67894 ( .A(n47584), .B(n47583), .Z(n50254) );
  NOR U67895 ( .A(n58179), .B(n50254), .Z(n47585) );
  IV U67896 ( .A(n47585), .Z(n58183) );
  XOR U67897 ( .A(n58182), .B(n58183), .Z(n47591) );
  IV U67898 ( .A(n47586), .Z(n47601) );
  NOR U67899 ( .A(n47587), .B(n47601), .Z(n47588) );
  IV U67900 ( .A(n47588), .Z(n47589) );
  NOR U67901 ( .A(n47594), .B(n47589), .Z(n47596) );
  IV U67902 ( .A(n47596), .Z(n47590) );
  NOR U67903 ( .A(n47591), .B(n47590), .Z(n58192) );
  IV U67904 ( .A(n47592), .Z(n47593) );
  NOR U67905 ( .A(n47594), .B(n47593), .Z(n55460) );
  NOR U67906 ( .A(n55460), .B(n58182), .Z(n47595) );
  XOR U67907 ( .A(n47595), .B(n58183), .Z(n50253) );
  NOR U67908 ( .A(n50253), .B(n47596), .Z(n47597) );
  NOR U67909 ( .A(n58192), .B(n47597), .Z(n47598) );
  IV U67910 ( .A(n47598), .Z(n50252) );
  IV U67911 ( .A(n47599), .Z(n47603) );
  XOR U67912 ( .A(n47601), .B(n47600), .Z(n47602) );
  NOR U67913 ( .A(n47603), .B(n47602), .Z(n47604) );
  IV U67914 ( .A(n47604), .Z(n47605) );
  NOR U67915 ( .A(n47606), .B(n47605), .Z(n50250) );
  XOR U67916 ( .A(n50252), .B(n50250), .Z(n50246) );
  IV U67917 ( .A(n47607), .Z(n47608) );
  NOR U67918 ( .A(n47609), .B(n47608), .Z(n47616) );
  IV U67919 ( .A(n47616), .Z(n47610) );
  NOR U67920 ( .A(n50246), .B(n47610), .Z(n58206) );
  IV U67921 ( .A(n47611), .Z(n47612) );
  NOR U67922 ( .A(n47612), .B(n47614), .Z(n50244) );
  XOR U67923 ( .A(n50246), .B(n50244), .Z(n50249) );
  IV U67924 ( .A(n47613), .Z(n47615) );
  NOR U67925 ( .A(n47615), .B(n47614), .Z(n50247) );
  XOR U67926 ( .A(n50249), .B(n50247), .Z(n47627) );
  IV U67927 ( .A(n47627), .Z(n47617) );
  NOR U67928 ( .A(n47617), .B(n47616), .Z(n47618) );
  NOR U67929 ( .A(n58206), .B(n47618), .Z(n47622) );
  XOR U67930 ( .A(n50240), .B(n47622), .Z(n47619) );
  NOR U67931 ( .A(n47620), .B(n47619), .Z(n47634) );
  IV U67932 ( .A(n47621), .Z(n47625) );
  IV U67933 ( .A(n47622), .Z(n50241) );
  NOR U67934 ( .A(n47628), .B(n50241), .Z(n47623) );
  IV U67935 ( .A(n47623), .Z(n47624) );
  NOR U67936 ( .A(n47625), .B(n47624), .Z(n58214) );
  IV U67937 ( .A(n47626), .Z(n47631) );
  NOR U67938 ( .A(n47628), .B(n47627), .Z(n47629) );
  IV U67939 ( .A(n47629), .Z(n47630) );
  NOR U67940 ( .A(n47631), .B(n47630), .Z(n58211) );
  NOR U67941 ( .A(n58214), .B(n58211), .Z(n47632) );
  IV U67942 ( .A(n47632), .Z(n47633) );
  NOR U67943 ( .A(n47634), .B(n47633), .Z(n47635) );
  IV U67944 ( .A(n47635), .Z(n55457) );
  XOR U67945 ( .A(n58219), .B(n55457), .Z(n50237) );
  IV U67946 ( .A(n50237), .Z(n47643) );
  IV U67947 ( .A(n47636), .Z(n47638) );
  NOR U67948 ( .A(n47638), .B(n47637), .Z(n55456) );
  IV U67949 ( .A(n47639), .Z(n47641) );
  NOR U67950 ( .A(n47641), .B(n47640), .Z(n50236) );
  NOR U67951 ( .A(n55456), .B(n50236), .Z(n47642) );
  XOR U67952 ( .A(n47643), .B(n47642), .Z(n50232) );
  XOR U67953 ( .A(n50230), .B(n50232), .Z(n50234) );
  XOR U67954 ( .A(n47644), .B(n50234), .Z(n50227) );
  XOR U67955 ( .A(n50229), .B(n50227), .Z(n53013) );
  IV U67956 ( .A(n47645), .Z(n47648) );
  IV U67957 ( .A(n47646), .Z(n47647) );
  NOR U67958 ( .A(n47648), .B(n47647), .Z(n53011) );
  XOR U67959 ( .A(n53013), .B(n53011), .Z(n50223) );
  XOR U67960 ( .A(n50222), .B(n50223), .Z(n50217) );
  IV U67961 ( .A(n47649), .Z(n47650) );
  NOR U67962 ( .A(n47650), .B(n47652), .Z(n50214) );
  NOR U67963 ( .A(n50221), .B(n50219), .Z(n47654) );
  IV U67964 ( .A(n47651), .Z(n47653) );
  NOR U67965 ( .A(n47653), .B(n47652), .Z(n50216) );
  NOR U67966 ( .A(n47654), .B(n50216), .Z(n47655) );
  IV U67967 ( .A(n47655), .Z(n47656) );
  NOR U67968 ( .A(n50214), .B(n47656), .Z(n47657) );
  XOR U67969 ( .A(n50217), .B(n47657), .Z(n47666) );
  IV U67970 ( .A(n47666), .Z(n55430) );
  IV U67971 ( .A(n47658), .Z(n47660) );
  NOR U67972 ( .A(n47660), .B(n47659), .Z(n50209) );
  XOR U67973 ( .A(n55430), .B(n50209), .Z(n47661) );
  NOR U67974 ( .A(n47662), .B(n47661), .Z(n63517) );
  IV U67975 ( .A(n47663), .Z(n55433) );
  NOR U67976 ( .A(n55433), .B(n47664), .Z(n50211) );
  NOR U67977 ( .A(n50211), .B(n50209), .Z(n47665) );
  XOR U67978 ( .A(n47666), .B(n47665), .Z(n50205) );
  IV U67979 ( .A(n50205), .Z(n47667) );
  NOR U67980 ( .A(n47668), .B(n47667), .Z(n47669) );
  NOR U67981 ( .A(n63517), .B(n47669), .Z(n47670) );
  IV U67982 ( .A(n47670), .Z(n50207) );
  IV U67983 ( .A(n47671), .Z(n47672) );
  NOR U67984 ( .A(n47672), .B(n47674), .Z(n50206) );
  IV U67985 ( .A(n47673), .Z(n47677) );
  XOR U67986 ( .A(n47675), .B(n47674), .Z(n47676) );
  NOR U67987 ( .A(n47677), .B(n47676), .Z(n50203) );
  NOR U67988 ( .A(n50206), .B(n50203), .Z(n47678) );
  XOR U67989 ( .A(n50207), .B(n47678), .Z(n50197) );
  IV U67990 ( .A(n47679), .Z(n47680) );
  NOR U67991 ( .A(n47688), .B(n47680), .Z(n50198) );
  IV U67992 ( .A(n47681), .Z(n47684) );
  IV U67993 ( .A(n47682), .Z(n47683) );
  NOR U67994 ( .A(n47684), .B(n47683), .Z(n50200) );
  NOR U67995 ( .A(n50198), .B(n50200), .Z(n47685) );
  XOR U67996 ( .A(n50197), .B(n47685), .Z(n50192) );
  IV U67997 ( .A(n47686), .Z(n47687) );
  NOR U67998 ( .A(n47688), .B(n47687), .Z(n50190) );
  XOR U67999 ( .A(n50192), .B(n50190), .Z(n55414) );
  IV U68000 ( .A(n47689), .Z(n50187) );
  NOR U68001 ( .A(n47690), .B(n50187), .Z(n47703) );
  IV U68002 ( .A(n47691), .Z(n47692) );
  NOR U68003 ( .A(n55417), .B(n47692), .Z(n50184) );
  NOR U68004 ( .A(n47703), .B(n50184), .Z(n47693) );
  XOR U68005 ( .A(n55414), .B(n47693), .Z(n47701) );
  IV U68006 ( .A(n47701), .Z(n47694) );
  NOR U68007 ( .A(n47695), .B(n47694), .Z(n50183) );
  IV U68008 ( .A(n47696), .Z(n47697) );
  NOR U68009 ( .A(n47697), .B(n47699), .Z(n53024) );
  IV U68010 ( .A(n47698), .Z(n47700) );
  NOR U68011 ( .A(n47700), .B(n47699), .Z(n47702) );
  NOR U68012 ( .A(n47702), .B(n47701), .Z(n47706) );
  IV U68013 ( .A(n47702), .Z(n47705) );
  XOR U68014 ( .A(n47703), .B(n55414), .Z(n47704) );
  NOR U68015 ( .A(n47705), .B(n47704), .Z(n55407) );
  NOR U68016 ( .A(n47706), .B(n55407), .Z(n53025) );
  XOR U68017 ( .A(n53024), .B(n53025), .Z(n47707) );
  NOR U68018 ( .A(n47708), .B(n47707), .Z(n47709) );
  NOR U68019 ( .A(n50183), .B(n47709), .Z(n50177) );
  IV U68020 ( .A(n47710), .Z(n47712) );
  NOR U68021 ( .A(n47712), .B(n47711), .Z(n47713) );
  IV U68022 ( .A(n47713), .Z(n50179) );
  XOR U68023 ( .A(n50177), .B(n50179), .Z(n50182) );
  XOR U68024 ( .A(n50180), .B(n50182), .Z(n50172) );
  XOR U68025 ( .A(n50171), .B(n50172), .Z(n50160) );
  XOR U68026 ( .A(n47714), .B(n50160), .Z(n55389) );
  NOR U68027 ( .A(n47723), .B(n55389), .Z(n58282) );
  NOR U68028 ( .A(n47715), .B(n50161), .Z(n47719) );
  IV U68029 ( .A(n47716), .Z(n47718) );
  NOR U68030 ( .A(n47718), .B(n47717), .Z(n55388) );
  NOR U68031 ( .A(n47719), .B(n55388), .Z(n47720) );
  XOR U68032 ( .A(n47720), .B(n55389), .Z(n53036) );
  IV U68033 ( .A(n47721), .Z(n47722) );
  NOR U68034 ( .A(n47722), .B(n47731), .Z(n53037) );
  XOR U68035 ( .A(n53036), .B(n53037), .Z(n47725) );
  NOR U68036 ( .A(n53037), .B(n47723), .Z(n47724) );
  NOR U68037 ( .A(n47725), .B(n47724), .Z(n47726) );
  NOR U68038 ( .A(n58282), .B(n47726), .Z(n47744) );
  IV U68039 ( .A(n47744), .Z(n53046) );
  IV U68040 ( .A(n47727), .Z(n47729) );
  IV U68041 ( .A(n47728), .Z(n47734) );
  NOR U68042 ( .A(n47729), .B(n47734), .Z(n53043) );
  IV U68043 ( .A(n47730), .Z(n47732) );
  NOR U68044 ( .A(n47732), .B(n47731), .Z(n53040) );
  IV U68045 ( .A(n47733), .Z(n47735) );
  NOR U68046 ( .A(n47735), .B(n47734), .Z(n53045) );
  NOR U68047 ( .A(n53040), .B(n53045), .Z(n47743) );
  IV U68048 ( .A(n47743), .Z(n47736) );
  NOR U68049 ( .A(n53043), .B(n47736), .Z(n47737) );
  XOR U68050 ( .A(n53046), .B(n47737), .Z(n47742) );
  IV U68051 ( .A(n47742), .Z(n47738) );
  NOR U68052 ( .A(n47749), .B(n47738), .Z(n58292) );
  IV U68053 ( .A(n47739), .Z(n47741) );
  NOR U68054 ( .A(n47741), .B(n47740), .Z(n47745) );
  NOR U68055 ( .A(n47745), .B(n47742), .Z(n47748) );
  XOR U68056 ( .A(n47744), .B(n47743), .Z(n47747) );
  IV U68057 ( .A(n47745), .Z(n47746) );
  NOR U68058 ( .A(n47747), .B(n47746), .Z(n60666) );
  NOR U68059 ( .A(n47748), .B(n60666), .Z(n53050) );
  XOR U68060 ( .A(n53049), .B(n53050), .Z(n47751) );
  NOR U68061 ( .A(n53050), .B(n47749), .Z(n47750) );
  NOR U68062 ( .A(n47751), .B(n47750), .Z(n47752) );
  NOR U68063 ( .A(n58292), .B(n47752), .Z(n50155) );
  IV U68064 ( .A(n47753), .Z(n50156) );
  NOR U68065 ( .A(n50158), .B(n50156), .Z(n47756) );
  IV U68066 ( .A(n47754), .Z(n47755) );
  NOR U68067 ( .A(n47755), .B(n47759), .Z(n53058) );
  NOR U68068 ( .A(n47756), .B(n53058), .Z(n47757) );
  XOR U68069 ( .A(n50155), .B(n47757), .Z(n50153) );
  IV U68070 ( .A(n47758), .Z(n47760) );
  NOR U68071 ( .A(n47760), .B(n47759), .Z(n50151) );
  XOR U68072 ( .A(n50153), .B(n50151), .Z(n53057) );
  XOR U68073 ( .A(n53055), .B(n53057), .Z(n50150) );
  XOR U68074 ( .A(n47761), .B(n50150), .Z(n53070) );
  IV U68075 ( .A(n47762), .Z(n47763) );
  NOR U68076 ( .A(n47764), .B(n47763), .Z(n47767) );
  IV U68077 ( .A(n53075), .Z(n47766) );
  NOR U68078 ( .A(n47766), .B(n47765), .Z(n50143) );
  NOR U68079 ( .A(n47767), .B(n50143), .Z(n53072) );
  XOR U68080 ( .A(n53070), .B(n53072), .Z(n53068) );
  XOR U68081 ( .A(n53067), .B(n53068), .Z(n50142) );
  XOR U68082 ( .A(n50140), .B(n50142), .Z(n53082) );
  XOR U68083 ( .A(n53080), .B(n53082), .Z(n50138) );
  XOR U68084 ( .A(n47768), .B(n50138), .Z(n53087) );
  XOR U68085 ( .A(n53088), .B(n53087), .Z(n50132) );
  XOR U68086 ( .A(n47780), .B(n50132), .Z(n47773) );
  IV U68087 ( .A(n47769), .Z(n47771) );
  NOR U68088 ( .A(n47771), .B(n47770), .Z(n47784) );
  IV U68089 ( .A(n47784), .Z(n47772) );
  NOR U68090 ( .A(n47773), .B(n47772), .Z(n55345) );
  IV U68091 ( .A(n47774), .Z(n47777) );
  NOR U68092 ( .A(n47775), .B(n47777), .Z(n50131) );
  IV U68093 ( .A(n47776), .Z(n47778) );
  NOR U68094 ( .A(n47778), .B(n47777), .Z(n50129) );
  NOR U68095 ( .A(n50131), .B(n50129), .Z(n47779) );
  IV U68096 ( .A(n47779), .Z(n47781) );
  NOR U68097 ( .A(n47781), .B(n47780), .Z(n47782) );
  XOR U68098 ( .A(n50132), .B(n47782), .Z(n47783) );
  NOR U68099 ( .A(n47784), .B(n47783), .Z(n53099) );
  NOR U68100 ( .A(n55345), .B(n53099), .Z(n50128) );
  XOR U68101 ( .A(n47785), .B(n50128), .Z(n50126) );
  XOR U68102 ( .A(n50124), .B(n50126), .Z(n50119) );
  XOR U68103 ( .A(n50118), .B(n50119), .Z(n50122) );
  XOR U68104 ( .A(n50121), .B(n50122), .Z(n47786) );
  XOR U68105 ( .A(n47787), .B(n47786), .Z(n53117) );
  IV U68106 ( .A(n47788), .Z(n47790) );
  NOR U68107 ( .A(n47790), .B(n47789), .Z(n53115) );
  IV U68108 ( .A(n47791), .Z(n53112) );
  NOR U68109 ( .A(n47792), .B(n53112), .Z(n47793) );
  NOR U68110 ( .A(n53115), .B(n47793), .Z(n47794) );
  XOR U68111 ( .A(n53117), .B(n47794), .Z(n50111) );
  IV U68112 ( .A(n47795), .Z(n47796) );
  NOR U68113 ( .A(n47796), .B(n47798), .Z(n53124) );
  IV U68114 ( .A(n47797), .Z(n47799) );
  NOR U68115 ( .A(n47799), .B(n47798), .Z(n53130) );
  NOR U68116 ( .A(n53124), .B(n53130), .Z(n50112) );
  XOR U68117 ( .A(n50111), .B(n50112), .Z(n53139) );
  XOR U68118 ( .A(n53138), .B(n53139), .Z(n47807) );
  IV U68119 ( .A(n47807), .Z(n53144) );
  XOR U68120 ( .A(n53140), .B(n53144), .Z(n47800) );
  NOR U68121 ( .A(n47801), .B(n47800), .Z(n58341) );
  IV U68122 ( .A(n47802), .Z(n47803) );
  NOR U68123 ( .A(n47806), .B(n47803), .Z(n47804) );
  IV U68124 ( .A(n47804), .Z(n53147) );
  NOR U68125 ( .A(n47806), .B(n47805), .Z(n53143) );
  NOR U68126 ( .A(n53143), .B(n53140), .Z(n47808) );
  XOR U68127 ( .A(n47808), .B(n47807), .Z(n53146) );
  XOR U68128 ( .A(n53147), .B(n53146), .Z(n47809) );
  NOR U68129 ( .A(n47810), .B(n47809), .Z(n47811) );
  NOR U68130 ( .A(n58341), .B(n47811), .Z(n47827) );
  IV U68131 ( .A(n47827), .Z(n55312) );
  XOR U68132 ( .A(n53149), .B(n55312), .Z(n47812) );
  NOR U68133 ( .A(n47826), .B(n47812), .Z(n47813) );
  IV U68134 ( .A(n47813), .Z(n47814) );
  NOR U68135 ( .A(n47815), .B(n47814), .Z(n47816) );
  IV U68136 ( .A(n47816), .Z(n55298) );
  NOR U68137 ( .A(n47825), .B(n55298), .Z(n53153) );
  IV U68138 ( .A(n47817), .Z(n47818) );
  NOR U68139 ( .A(n47818), .B(n47820), .Z(n50101) );
  IV U68140 ( .A(n47819), .Z(n47821) );
  NOR U68141 ( .A(n47821), .B(n47820), .Z(n50099) );
  NOR U68142 ( .A(n50101), .B(n50099), .Z(n47833) );
  IV U68143 ( .A(n47833), .Z(n47822) );
  NOR U68144 ( .A(n53153), .B(n47822), .Z(n47823) );
  IV U68145 ( .A(n47823), .Z(n47831) );
  NOR U68146 ( .A(n47825), .B(n47824), .Z(n47829) );
  NOR U68147 ( .A(n53149), .B(n47826), .Z(n47828) );
  XOR U68148 ( .A(n47828), .B(n47827), .Z(n50103) );
  IV U68149 ( .A(n50103), .Z(n47832) );
  NOR U68150 ( .A(n47829), .B(n47832), .Z(n47830) );
  NOR U68151 ( .A(n47831), .B(n47830), .Z(n47835) );
  NOR U68152 ( .A(n47833), .B(n47832), .Z(n47834) );
  NOR U68153 ( .A(n47835), .B(n47834), .Z(n53159) );
  IV U68154 ( .A(n47836), .Z(n47846) );
  IV U68155 ( .A(n47837), .Z(n47838) );
  NOR U68156 ( .A(n47846), .B(n47838), .Z(n53155) );
  IV U68157 ( .A(n47839), .Z(n47841) );
  NOR U68158 ( .A(n47841), .B(n47840), .Z(n53157) );
  NOR U68159 ( .A(n53155), .B(n53157), .Z(n47842) );
  XOR U68160 ( .A(n53159), .B(n47842), .Z(n47843) );
  IV U68161 ( .A(n47843), .Z(n50098) );
  IV U68162 ( .A(n47844), .Z(n47845) );
  NOR U68163 ( .A(n47846), .B(n47845), .Z(n50096) );
  XOR U68164 ( .A(n50098), .B(n50096), .Z(n53172) );
  NOR U68165 ( .A(n47848), .B(n47847), .Z(n53165) );
  NOR U68166 ( .A(n53165), .B(n47849), .Z(n47850) );
  XOR U68167 ( .A(n53172), .B(n47850), .Z(n47851) );
  IV U68168 ( .A(n47851), .Z(n53170) );
  IV U68169 ( .A(n47852), .Z(n47853) );
  NOR U68170 ( .A(n47853), .B(n47856), .Z(n47860) );
  IV U68171 ( .A(n47860), .Z(n47854) );
  NOR U68172 ( .A(n53170), .B(n47854), .Z(n58366) );
  IV U68173 ( .A(n47855), .Z(n47857) );
  NOR U68174 ( .A(n47857), .B(n47856), .Z(n47858) );
  IV U68175 ( .A(n47858), .Z(n53169) );
  XOR U68176 ( .A(n53170), .B(n53169), .Z(n47859) );
  NOR U68177 ( .A(n47860), .B(n47859), .Z(n53180) );
  IV U68178 ( .A(n47861), .Z(n47863) );
  NOR U68179 ( .A(n47863), .B(n47862), .Z(n53178) );
  XOR U68180 ( .A(n53180), .B(n53178), .Z(n47864) );
  NOR U68181 ( .A(n58366), .B(n47864), .Z(n53176) );
  IV U68182 ( .A(n47865), .Z(n47866) );
  NOR U68183 ( .A(n47869), .B(n47866), .Z(n53175) );
  IV U68184 ( .A(n47867), .Z(n47868) );
  NOR U68185 ( .A(n47869), .B(n47868), .Z(n53184) );
  NOR U68186 ( .A(n53175), .B(n53184), .Z(n47870) );
  XOR U68187 ( .A(n53176), .B(n47870), .Z(n53192) );
  IV U68188 ( .A(n47871), .Z(n47880) );
  IV U68189 ( .A(n47872), .Z(n47873) );
  NOR U68190 ( .A(n47880), .B(n47873), .Z(n53190) );
  IV U68191 ( .A(n47874), .Z(n47876) );
  NOR U68192 ( .A(n47876), .B(n47875), .Z(n53187) );
  NOR U68193 ( .A(n53190), .B(n53187), .Z(n47877) );
  XOR U68194 ( .A(n53192), .B(n47877), .Z(n53193) );
  IV U68195 ( .A(n47878), .Z(n47879) );
  NOR U68196 ( .A(n47880), .B(n47879), .Z(n47881) );
  IV U68197 ( .A(n47881), .Z(n53194) );
  XOR U68198 ( .A(n53193), .B(n53194), .Z(n53197) );
  XOR U68199 ( .A(n53196), .B(n53197), .Z(n50091) );
  XOR U68200 ( .A(n50093), .B(n50091), .Z(n55265) );
  IV U68201 ( .A(n47882), .Z(n53217) );
  NOR U68202 ( .A(n47883), .B(n53217), .Z(n47887) );
  IV U68203 ( .A(n47884), .Z(n47886) );
  NOR U68204 ( .A(n47886), .B(n47885), .Z(n55268) );
  NOR U68205 ( .A(n47887), .B(n55268), .Z(n47888) );
  XOR U68206 ( .A(n55265), .B(n47888), .Z(n47889) );
  IV U68207 ( .A(n47889), .Z(n53215) );
  XOR U68208 ( .A(n53213), .B(n53215), .Z(n50082) );
  XOR U68209 ( .A(n50081), .B(n50082), .Z(n58396) );
  XOR U68210 ( .A(n47890), .B(n58396), .Z(n47891) );
  IV U68211 ( .A(n47891), .Z(n50074) );
  XOR U68212 ( .A(n50073), .B(n50074), .Z(n47892) );
  XOR U68213 ( .A(n47893), .B(n47892), .Z(n50068) );
  IV U68214 ( .A(n47894), .Z(n47897) );
  IV U68215 ( .A(n47895), .Z(n47896) );
  NOR U68216 ( .A(n47897), .B(n47896), .Z(n47898) );
  IV U68217 ( .A(n47898), .Z(n50069) );
  XOR U68218 ( .A(n50068), .B(n50069), .Z(n50067) );
  IV U68219 ( .A(n47899), .Z(n47902) );
  IV U68220 ( .A(n47900), .Z(n47901) );
  NOR U68221 ( .A(n47902), .B(n47901), .Z(n50065) );
  IV U68222 ( .A(n47903), .Z(n47904) );
  NOR U68223 ( .A(n47905), .B(n47904), .Z(n50063) );
  NOR U68224 ( .A(n50065), .B(n50063), .Z(n47906) );
  XOR U68225 ( .A(n50067), .B(n47906), .Z(n47907) );
  IV U68226 ( .A(n47907), .Z(n50062) );
  XOR U68227 ( .A(n50060), .B(n50062), .Z(n55252) );
  IV U68228 ( .A(n47908), .Z(n47911) );
  NOR U68229 ( .A(n47909), .B(n47911), .Z(n58421) );
  IV U68230 ( .A(n47910), .Z(n47912) );
  NOR U68231 ( .A(n47912), .B(n47911), .Z(n55251) );
  NOR U68232 ( .A(n58421), .B(n55251), .Z(n50059) );
  XOR U68233 ( .A(n55252), .B(n50059), .Z(n47913) );
  IV U68234 ( .A(n47913), .Z(n53228) );
  XOR U68235 ( .A(n53227), .B(n53228), .Z(n53231) );
  XOR U68236 ( .A(n53230), .B(n53231), .Z(n55241) );
  XOR U68237 ( .A(n50055), .B(n55241), .Z(n47914) );
  NOR U68238 ( .A(n47915), .B(n47914), .Z(n55244) );
  IV U68239 ( .A(n47916), .Z(n47917) );
  NOR U68240 ( .A(n47917), .B(n47919), .Z(n55248) );
  IV U68241 ( .A(n47918), .Z(n47920) );
  NOR U68242 ( .A(n47920), .B(n47919), .Z(n55239) );
  NOR U68243 ( .A(n55248), .B(n55239), .Z(n50054) );
  IV U68244 ( .A(n50054), .Z(n47921) );
  NOR U68245 ( .A(n50055), .B(n47921), .Z(n47922) );
  XOR U68246 ( .A(n55241), .B(n47922), .Z(n50046) );
  NOR U68247 ( .A(n47923), .B(n50046), .Z(n47924) );
  NOR U68248 ( .A(n55244), .B(n47924), .Z(n50051) );
  IV U68249 ( .A(n47925), .Z(n47928) );
  IV U68250 ( .A(n47926), .Z(n47927) );
  NOR U68251 ( .A(n47928), .B(n47927), .Z(n50047) );
  NOR U68252 ( .A(n50050), .B(n50047), .Z(n47929) );
  XOR U68253 ( .A(n50051), .B(n47929), .Z(n50045) );
  IV U68254 ( .A(n47930), .Z(n47931) );
  NOR U68255 ( .A(n47932), .B(n47931), .Z(n50041) );
  IV U68256 ( .A(n47933), .Z(n47936) );
  IV U68257 ( .A(n47934), .Z(n47935) );
  NOR U68258 ( .A(n47936), .B(n47935), .Z(n50043) );
  NOR U68259 ( .A(n50041), .B(n50043), .Z(n47937) );
  XOR U68260 ( .A(n50045), .B(n47937), .Z(n47938) );
  NOR U68261 ( .A(n47939), .B(n47938), .Z(n47942) );
  IV U68262 ( .A(n47939), .Z(n47941) );
  XOR U68263 ( .A(n50045), .B(n50043), .Z(n47940) );
  NOR U68264 ( .A(n47941), .B(n47940), .Z(n58453) );
  NOR U68265 ( .A(n47942), .B(n58453), .Z(n53244) );
  IV U68266 ( .A(n47943), .Z(n47944) );
  NOR U68267 ( .A(n47944), .B(n47946), .Z(n53248) );
  IV U68268 ( .A(n47945), .Z(n47947) );
  NOR U68269 ( .A(n47947), .B(n47946), .Z(n53243) );
  NOR U68270 ( .A(n53248), .B(n53243), .Z(n47948) );
  XOR U68271 ( .A(n53244), .B(n47948), .Z(n53252) );
  XOR U68272 ( .A(n53251), .B(n53252), .Z(n47952) );
  IV U68273 ( .A(n47952), .Z(n53258) );
  XOR U68274 ( .A(n53256), .B(n53258), .Z(n58479) );
  NOR U68275 ( .A(n47949), .B(n58479), .Z(n58474) );
  IV U68276 ( .A(n47950), .Z(n47951) );
  NOR U68277 ( .A(n47956), .B(n47951), .Z(n53254) );
  NOR U68278 ( .A(n53254), .B(n53256), .Z(n47953) );
  XOR U68279 ( .A(n47953), .B(n47952), .Z(n50040) );
  IV U68280 ( .A(n47954), .Z(n47955) );
  NOR U68281 ( .A(n47956), .B(n47955), .Z(n47957) );
  IV U68282 ( .A(n47957), .Z(n50039) );
  XOR U68283 ( .A(n50040), .B(n50039), .Z(n47958) );
  NOR U68284 ( .A(n47959), .B(n47958), .Z(n47960) );
  NOR U68285 ( .A(n58474), .B(n47960), .Z(n50034) );
  XOR U68286 ( .A(n58482), .B(n50034), .Z(n55221) );
  NOR U68287 ( .A(n47961), .B(n55221), .Z(n55214) );
  IV U68288 ( .A(n47962), .Z(n47963) );
  NOR U68289 ( .A(n47967), .B(n47963), .Z(n47964) );
  IV U68290 ( .A(n47964), .Z(n55217) );
  IV U68291 ( .A(n47965), .Z(n47966) );
  NOR U68292 ( .A(n47967), .B(n47966), .Z(n55220) );
  XOR U68293 ( .A(n55220), .B(n55221), .Z(n55216) );
  XOR U68294 ( .A(n55217), .B(n55216), .Z(n50036) );
  NOR U68295 ( .A(n47968), .B(n50036), .Z(n47969) );
  NOR U68296 ( .A(n55214), .B(n47969), .Z(n53261) );
  XOR U68297 ( .A(n53262), .B(n53261), .Z(n53266) );
  XOR U68298 ( .A(n53265), .B(n53266), .Z(n55205) );
  IV U68299 ( .A(n47970), .Z(n55208) );
  NOR U68300 ( .A(n47971), .B(n55208), .Z(n50032) );
  IV U68301 ( .A(n47972), .Z(n47974) );
  NOR U68302 ( .A(n47974), .B(n47973), .Z(n53268) );
  NOR U68303 ( .A(n50032), .B(n53268), .Z(n47975) );
  XOR U68304 ( .A(n55205), .B(n47975), .Z(n47985) );
  IV U68305 ( .A(n47985), .Z(n47976) );
  NOR U68306 ( .A(n47988), .B(n47976), .Z(n55200) );
  IV U68307 ( .A(n47977), .Z(n47980) );
  XOR U68308 ( .A(n47978), .B(n47981), .Z(n47979) );
  NOR U68309 ( .A(n47980), .B(n47979), .Z(n50029) );
  NOR U68310 ( .A(n47982), .B(n47981), .Z(n47986) );
  IV U68311 ( .A(n47986), .Z(n47984) );
  XOR U68312 ( .A(n53268), .B(n55205), .Z(n47983) );
  NOR U68313 ( .A(n47984), .B(n47983), .Z(n58496) );
  NOR U68314 ( .A(n47986), .B(n47985), .Z(n47987) );
  NOR U68315 ( .A(n58496), .B(n47987), .Z(n47996) );
  XOR U68316 ( .A(n50029), .B(n47996), .Z(n47990) );
  NOR U68317 ( .A(n47996), .B(n47988), .Z(n47989) );
  NOR U68318 ( .A(n47990), .B(n47989), .Z(n47991) );
  NOR U68319 ( .A(n55200), .B(n47991), .Z(n48002) );
  IV U68320 ( .A(n48002), .Z(n48012) );
  IV U68321 ( .A(n47992), .Z(n47999) );
  IV U68322 ( .A(n47993), .Z(n47994) );
  NOR U68323 ( .A(n47999), .B(n47994), .Z(n48005) );
  IV U68324 ( .A(n48005), .Z(n47995) );
  NOR U68325 ( .A(n48012), .B(n47995), .Z(n58517) );
  IV U68326 ( .A(n47996), .Z(n50030) );
  IV U68327 ( .A(n47997), .Z(n47998) );
  NOR U68328 ( .A(n47999), .B(n47998), .Z(n48001) );
  IV U68329 ( .A(n48001), .Z(n48000) );
  NOR U68330 ( .A(n50030), .B(n48000), .Z(n55199) );
  NOR U68331 ( .A(n48002), .B(n48001), .Z(n48003) );
  NOR U68332 ( .A(n55199), .B(n48003), .Z(n48004) );
  NOR U68333 ( .A(n48005), .B(n48004), .Z(n48006) );
  NOR U68334 ( .A(n58517), .B(n48006), .Z(n48014) );
  IV U68335 ( .A(n48014), .Z(n48007) );
  NOR U68336 ( .A(n48008), .B(n48007), .Z(n55193) );
  IV U68337 ( .A(n48009), .Z(n48011) );
  NOR U68338 ( .A(n48011), .B(n48010), .Z(n48015) );
  IV U68339 ( .A(n48015), .Z(n48013) );
  NOR U68340 ( .A(n48013), .B(n48012), .Z(n58518) );
  NOR U68341 ( .A(n48015), .B(n48014), .Z(n48016) );
  NOR U68342 ( .A(n58518), .B(n48016), .Z(n48024) );
  NOR U68343 ( .A(n48017), .B(n48024), .Z(n48018) );
  NOR U68344 ( .A(n55193), .B(n48018), .Z(n50026) );
  IV U68345 ( .A(n48019), .Z(n48020) );
  NOR U68346 ( .A(n48020), .B(n48022), .Z(n48031) );
  IV U68347 ( .A(n48031), .Z(n50028) );
  NOR U68348 ( .A(n50026), .B(n50028), .Z(n48033) );
  IV U68349 ( .A(n48021), .Z(n48023) );
  NOR U68350 ( .A(n48023), .B(n48022), .Z(n48027) );
  IV U68351 ( .A(n48027), .Z(n48026) );
  IV U68352 ( .A(n48024), .Z(n48025) );
  NOR U68353 ( .A(n48026), .B(n48025), .Z(n55196) );
  NOR U68354 ( .A(n50026), .B(n48027), .Z(n48028) );
  NOR U68355 ( .A(n55196), .B(n48028), .Z(n48029) );
  IV U68356 ( .A(n48029), .Z(n48030) );
  NOR U68357 ( .A(n48031), .B(n48030), .Z(n48032) );
  NOR U68358 ( .A(n48033), .B(n48032), .Z(n53280) );
  XOR U68359 ( .A(n53279), .B(n53280), .Z(n50025) );
  IV U68360 ( .A(n48034), .Z(n48039) );
  IV U68361 ( .A(n48035), .Z(n48036) );
  NOR U68362 ( .A(n48039), .B(n48036), .Z(n50023) );
  XOR U68363 ( .A(n50025), .B(n50023), .Z(n50021) );
  IV U68364 ( .A(n48037), .Z(n48038) );
  NOR U68365 ( .A(n48039), .B(n48038), .Z(n50019) );
  XOR U68366 ( .A(n50021), .B(n50019), .Z(n48044) );
  NOR U68367 ( .A(n48040), .B(n48044), .Z(n50013) );
  IV U68368 ( .A(n48041), .Z(n48042) );
  NOR U68369 ( .A(n48042), .B(n55188), .Z(n48046) );
  IV U68370 ( .A(n48046), .Z(n48043) );
  NOR U68371 ( .A(n48043), .B(n50025), .Z(n50022) );
  IV U68372 ( .A(n48044), .Z(n48045) );
  NOR U68373 ( .A(n48046), .B(n48045), .Z(n48047) );
  NOR U68374 ( .A(n50022), .B(n48047), .Z(n48053) );
  NOR U68375 ( .A(n48048), .B(n48053), .Z(n48049) );
  NOR U68376 ( .A(n50013), .B(n48049), .Z(n48065) );
  IV U68377 ( .A(n48050), .Z(n48052) );
  IV U68378 ( .A(n48051), .Z(n55176) );
  NOR U68379 ( .A(n48052), .B(n55176), .Z(n48054) );
  NOR U68380 ( .A(n48065), .B(n48054), .Z(n48062) );
  IV U68381 ( .A(n48053), .Z(n55177) );
  IV U68382 ( .A(n48054), .Z(n48055) );
  NOR U68383 ( .A(n55177), .B(n48055), .Z(n58529) );
  IV U68384 ( .A(n48056), .Z(n48058) );
  NOR U68385 ( .A(n48058), .B(n48057), .Z(n48068) );
  IV U68386 ( .A(n48068), .Z(n48059) );
  NOR U68387 ( .A(n58529), .B(n48059), .Z(n48060) );
  IV U68388 ( .A(n48060), .Z(n48061) );
  NOR U68389 ( .A(n48062), .B(n48061), .Z(n55167) );
  NOR U68390 ( .A(n48063), .B(n55176), .Z(n48066) );
  IV U68391 ( .A(n48066), .Z(n48064) );
  NOR U68392 ( .A(n48064), .B(n55177), .Z(n53290) );
  NOR U68393 ( .A(n48066), .B(n48065), .Z(n48067) );
  NOR U68394 ( .A(n53290), .B(n48067), .Z(n48071) );
  NOR U68395 ( .A(n48068), .B(n48071), .Z(n48069) );
  NOR U68396 ( .A(n55167), .B(n48069), .Z(n48070) );
  NOR U68397 ( .A(n48072), .B(n48070), .Z(n48075) );
  IV U68398 ( .A(n48071), .Z(n48074) );
  IV U68399 ( .A(n48072), .Z(n48073) );
  NOR U68400 ( .A(n48074), .B(n48073), .Z(n55170) );
  NOR U68401 ( .A(n48075), .B(n55170), .Z(n50011) );
  IV U68402 ( .A(n48076), .Z(n48078) );
  NOR U68403 ( .A(n48078), .B(n48077), .Z(n48088) );
  IV U68404 ( .A(n48088), .Z(n50012) );
  XOR U68405 ( .A(n50011), .B(n50012), .Z(n53298) );
  IV U68406 ( .A(n53298), .Z(n48084) );
  IV U68407 ( .A(n48079), .Z(n48080) );
  NOR U68408 ( .A(n48080), .B(n48082), .Z(n50008) );
  IV U68409 ( .A(n48081), .Z(n48083) );
  NOR U68410 ( .A(n48083), .B(n48082), .Z(n53296) );
  NOR U68411 ( .A(n50008), .B(n53296), .Z(n48085) );
  NOR U68412 ( .A(n48084), .B(n48085), .Z(n48093) );
  IV U68413 ( .A(n48085), .Z(n48091) );
  IV U68414 ( .A(n48086), .Z(n55159) );
  NOR U68415 ( .A(n55159), .B(n48087), .Z(n53293) );
  NOR U68416 ( .A(n53293), .B(n48088), .Z(n48089) );
  XOR U68417 ( .A(n50011), .B(n48089), .Z(n48090) );
  NOR U68418 ( .A(n48091), .B(n48090), .Z(n48092) );
  NOR U68419 ( .A(n48093), .B(n48092), .Z(n53300) );
  XOR U68420 ( .A(n48094), .B(n53300), .Z(n49999) );
  XOR U68421 ( .A(n50000), .B(n49999), .Z(n49998) );
  IV U68422 ( .A(n48095), .Z(n48107) );
  IV U68423 ( .A(n48096), .Z(n48097) );
  NOR U68424 ( .A(n48107), .B(n48097), .Z(n49996) );
  IV U68425 ( .A(n48098), .Z(n48100) );
  NOR U68426 ( .A(n48100), .B(n48099), .Z(n50001) );
  NOR U68427 ( .A(n49996), .B(n50001), .Z(n48101) );
  XOR U68428 ( .A(n49998), .B(n48101), .Z(n53308) );
  IV U68429 ( .A(n48102), .Z(n48104) );
  NOR U68430 ( .A(n48104), .B(n48103), .Z(n55125) );
  IV U68431 ( .A(n48105), .Z(n48106) );
  NOR U68432 ( .A(n48107), .B(n48106), .Z(n53311) );
  NOR U68433 ( .A(n55125), .B(n53311), .Z(n48108) );
  XOR U68434 ( .A(n53308), .B(n48108), .Z(n58539) );
  XOR U68435 ( .A(n53310), .B(n58539), .Z(n49995) );
  XOR U68436 ( .A(n49993), .B(n49995), .Z(n49989) );
  XOR U68437 ( .A(n48109), .B(n49989), .Z(n48110) );
  IV U68438 ( .A(n48110), .Z(n49974) );
  XOR U68439 ( .A(n49972), .B(n49974), .Z(n49977) );
  IV U68440 ( .A(n48111), .Z(n48113) );
  NOR U68441 ( .A(n48113), .B(n48112), .Z(n49975) );
  XOR U68442 ( .A(n49977), .B(n49975), .Z(n49963) );
  XOR U68443 ( .A(n49964), .B(n49963), .Z(n48119) );
  IV U68444 ( .A(n48119), .Z(n58578) );
  NOR U68445 ( .A(n48114), .B(n58578), .Z(n53322) );
  IV U68446 ( .A(n48115), .Z(n48117) );
  NOR U68447 ( .A(n48117), .B(n48116), .Z(n48120) );
  IV U68448 ( .A(n48120), .Z(n48118) );
  NOR U68449 ( .A(n48118), .B(n49963), .Z(n58573) );
  NOR U68450 ( .A(n48120), .B(n48119), .Z(n48121) );
  NOR U68451 ( .A(n58573), .B(n48121), .Z(n48126) );
  NOR U68452 ( .A(n48122), .B(n48126), .Z(n48123) );
  NOR U68453 ( .A(n53322), .B(n48123), .Z(n48124) );
  NOR U68454 ( .A(n48125), .B(n48124), .Z(n48129) );
  IV U68455 ( .A(n48125), .Z(n48128) );
  IV U68456 ( .A(n48126), .Z(n48127) );
  NOR U68457 ( .A(n48128), .B(n48127), .Z(n60447) );
  NOR U68458 ( .A(n48129), .B(n60447), .Z(n48130) );
  IV U68459 ( .A(n48130), .Z(n49961) );
  XOR U68460 ( .A(n49960), .B(n49961), .Z(n53324) );
  IV U68461 ( .A(n53324), .Z(n48146) );
  NOR U68462 ( .A(n48131), .B(n48146), .Z(n48141) );
  IV U68463 ( .A(n48132), .Z(n48135) );
  NOR U68464 ( .A(n48133), .B(n49961), .Z(n48134) );
  IV U68465 ( .A(n48134), .Z(n48137) );
  NOR U68466 ( .A(n48135), .B(n48137), .Z(n49959) );
  IV U68467 ( .A(n48136), .Z(n48138) );
  NOR U68468 ( .A(n48138), .B(n48137), .Z(n58592) );
  NOR U68469 ( .A(n49959), .B(n58592), .Z(n48139) );
  IV U68470 ( .A(n48139), .Z(n48140) );
  NOR U68471 ( .A(n48141), .B(n48140), .Z(n48142) );
  IV U68472 ( .A(n48142), .Z(n49952) );
  IV U68473 ( .A(n48143), .Z(n49953) );
  XOR U68474 ( .A(n49949), .B(n53339), .Z(n53335) );
  XOR U68475 ( .A(n53334), .B(n53335), .Z(n49942) );
  IV U68476 ( .A(n48147), .Z(n53338) );
  NOR U68477 ( .A(n48148), .B(n53338), .Z(n48151) );
  NOR U68478 ( .A(n48149), .B(n49943), .Z(n48150) );
  NOR U68479 ( .A(n48151), .B(n48150), .Z(n48152) );
  XOR U68480 ( .A(n49942), .B(n48152), .Z(n48166) );
  IV U68481 ( .A(n48166), .Z(n55083) );
  XOR U68482 ( .A(n49939), .B(n55083), .Z(n48157) );
  IV U68483 ( .A(n48153), .Z(n48155) );
  XOR U68484 ( .A(n48160), .B(n48161), .Z(n48154) );
  NOR U68485 ( .A(n48155), .B(n48154), .Z(n48167) );
  IV U68486 ( .A(n48167), .Z(n48156) );
  NOR U68487 ( .A(n48157), .B(n48156), .Z(n58617) );
  IV U68488 ( .A(n48158), .Z(n48159) );
  NOR U68489 ( .A(n48159), .B(n48161), .Z(n49935) );
  IV U68490 ( .A(n48160), .Z(n48162) );
  NOR U68491 ( .A(n48162), .B(n48161), .Z(n49937) );
  NOR U68492 ( .A(n49935), .B(n49937), .Z(n48163) );
  IV U68493 ( .A(n48163), .Z(n48164) );
  NOR U68494 ( .A(n49939), .B(n48164), .Z(n48165) );
  XOR U68495 ( .A(n48166), .B(n48165), .Z(n48173) );
  IV U68496 ( .A(n48173), .Z(n48168) );
  NOR U68497 ( .A(n48168), .B(n48167), .Z(n48169) );
  NOR U68498 ( .A(n58617), .B(n48169), .Z(n48170) );
  NOR U68499 ( .A(n48171), .B(n48170), .Z(n48174) );
  IV U68500 ( .A(n48171), .Z(n48172) );
  NOR U68501 ( .A(n48173), .B(n48172), .Z(n55072) );
  NOR U68502 ( .A(n48174), .B(n55072), .Z(n53350) );
  IV U68503 ( .A(n48178), .Z(n48175) );
  NOR U68504 ( .A(n48176), .B(n48175), .Z(n55073) );
  NOR U68505 ( .A(n48178), .B(n48177), .Z(n48181) );
  IV U68506 ( .A(n48179), .Z(n48180) );
  NOR U68507 ( .A(n48181), .B(n48180), .Z(n55068) );
  NOR U68508 ( .A(n55073), .B(n55068), .Z(n53351) );
  XOR U68509 ( .A(n53350), .B(n53351), .Z(n49934) );
  XOR U68510 ( .A(n49932), .B(n49934), .Z(n53363) );
  XOR U68511 ( .A(n48188), .B(n53363), .Z(n48182) );
  NOR U68512 ( .A(n48190), .B(n48182), .Z(n58635) );
  IV U68513 ( .A(n48183), .Z(n48184) );
  NOR U68514 ( .A(n48184), .B(n48186), .Z(n49924) );
  IV U68515 ( .A(n48185), .Z(n48187) );
  NOR U68516 ( .A(n48187), .B(n48186), .Z(n53362) );
  NOR U68517 ( .A(n48188), .B(n53362), .Z(n48189) );
  XOR U68518 ( .A(n48189), .B(n53363), .Z(n49925) );
  XOR U68519 ( .A(n49924), .B(n49925), .Z(n48192) );
  NOR U68520 ( .A(n49925), .B(n48190), .Z(n48191) );
  NOR U68521 ( .A(n48192), .B(n48191), .Z(n48193) );
  NOR U68522 ( .A(n58635), .B(n48193), .Z(n49920) );
  IV U68523 ( .A(n48194), .Z(n48196) );
  NOR U68524 ( .A(n48196), .B(n48195), .Z(n48197) );
  IV U68525 ( .A(n48197), .Z(n49922) );
  XOR U68526 ( .A(n49920), .B(n49922), .Z(n53377) );
  XOR U68527 ( .A(n48198), .B(n53377), .Z(n49913) );
  IV U68528 ( .A(n48199), .Z(n48201) );
  NOR U68529 ( .A(n48201), .B(n48200), .Z(n49917) );
  IV U68530 ( .A(n48202), .Z(n48204) );
  NOR U68531 ( .A(n48204), .B(n48203), .Z(n49915) );
  NOR U68532 ( .A(n49917), .B(n49915), .Z(n48205) );
  XOR U68533 ( .A(n49913), .B(n48205), .Z(n49905) );
  XOR U68534 ( .A(n48206), .B(n49905), .Z(n49901) );
  XOR U68535 ( .A(n48207), .B(n49901), .Z(n49899) );
  XOR U68536 ( .A(n49897), .B(n49899), .Z(n49896) );
  IV U68537 ( .A(n48208), .Z(n48216) );
  IV U68538 ( .A(n48209), .Z(n48210) );
  NOR U68539 ( .A(n48216), .B(n48210), .Z(n48211) );
  IV U68540 ( .A(n48211), .Z(n48217) );
  NOR U68541 ( .A(n49896), .B(n48217), .Z(n58659) );
  IV U68542 ( .A(n48212), .Z(n48213) );
  NOR U68543 ( .A(n48213), .B(n48223), .Z(n49891) );
  IV U68544 ( .A(n48214), .Z(n48215) );
  NOR U68545 ( .A(n48216), .B(n48215), .Z(n49894) );
  XOR U68546 ( .A(n49896), .B(n49894), .Z(n49892) );
  IV U68547 ( .A(n49892), .Z(n48218) );
  XOR U68548 ( .A(n49891), .B(n48218), .Z(n48220) );
  NOR U68549 ( .A(n48218), .B(n48217), .Z(n48219) );
  NOR U68550 ( .A(n48220), .B(n48219), .Z(n48221) );
  NOR U68551 ( .A(n58659), .B(n48221), .Z(n49886) );
  IV U68552 ( .A(n48222), .Z(n48224) );
  NOR U68553 ( .A(n48224), .B(n48223), .Z(n49889) );
  IV U68554 ( .A(n48225), .Z(n48229) );
  NOR U68555 ( .A(n48226), .B(n48229), .Z(n49885) );
  NOR U68556 ( .A(n49889), .B(n49885), .Z(n48227) );
  XOR U68557 ( .A(n49886), .B(n48227), .Z(n49884) );
  IV U68558 ( .A(n48228), .Z(n48230) );
  NOR U68559 ( .A(n48230), .B(n48229), .Z(n49882) );
  XOR U68560 ( .A(n49884), .B(n49882), .Z(n55039) );
  XOR U68561 ( .A(n49880), .B(n55039), .Z(n49876) );
  XOR U68562 ( .A(n48231), .B(n49876), .Z(n53394) );
  XOR U68563 ( .A(n53393), .B(n53394), .Z(n53401) );
  XOR U68564 ( .A(n53400), .B(n53401), .Z(n53405) );
  XOR U68565 ( .A(n53403), .B(n53405), .Z(n49866) );
  XOR U68566 ( .A(n49863), .B(n49866), .Z(n49861) );
  XOR U68567 ( .A(n49859), .B(n49861), .Z(n48232) );
  XOR U68568 ( .A(n48233), .B(n48232), .Z(n49858) );
  XOR U68569 ( .A(n48234), .B(n49858), .Z(n48235) );
  IV U68570 ( .A(n48235), .Z(n49852) );
  XOR U68571 ( .A(n48236), .B(n49852), .Z(n49843) );
  IV U68572 ( .A(n48237), .Z(n48238) );
  NOR U68573 ( .A(n48239), .B(n48238), .Z(n49844) );
  IV U68574 ( .A(n48240), .Z(n48243) );
  IV U68575 ( .A(n48241), .Z(n48242) );
  NOR U68576 ( .A(n48243), .B(n48242), .Z(n49848) );
  NOR U68577 ( .A(n49844), .B(n49848), .Z(n48244) );
  XOR U68578 ( .A(n49843), .B(n48244), .Z(n49842) );
  XOR U68579 ( .A(n49840), .B(n49842), .Z(n53412) );
  XOR U68580 ( .A(n48245), .B(n53412), .Z(n48246) );
  IV U68581 ( .A(n48246), .Z(n53415) );
  XOR U68582 ( .A(n53414), .B(n53415), .Z(n48252) );
  IV U68583 ( .A(n48252), .Z(n48247) );
  NOR U68584 ( .A(n48248), .B(n48247), .Z(n48255) );
  IV U68585 ( .A(n48249), .Z(n48250) );
  NOR U68586 ( .A(n48250), .B(n53415), .Z(n58726) );
  IV U68587 ( .A(n48251), .Z(n48253) );
  NOR U68588 ( .A(n48253), .B(n48252), .Z(n55002) );
  NOR U68589 ( .A(n58726), .B(n55002), .Z(n48254) );
  IV U68590 ( .A(n48254), .Z(n53418) );
  NOR U68591 ( .A(n48255), .B(n53418), .Z(n53419) );
  XOR U68592 ( .A(n53420), .B(n53419), .Z(n53422) );
  XOR U68593 ( .A(n48256), .B(n53422), .Z(n53442) );
  XOR U68594 ( .A(n48257), .B(n53442), .Z(n53454) );
  XOR U68595 ( .A(n53455), .B(n53454), .Z(n53458) );
  IV U68596 ( .A(n48258), .Z(n48259) );
  NOR U68597 ( .A(n48260), .B(n48259), .Z(n49828) );
  IV U68598 ( .A(n48261), .Z(n48263) );
  NOR U68599 ( .A(n48263), .B(n48262), .Z(n53456) );
  NOR U68600 ( .A(n49828), .B(n53456), .Z(n48264) );
  XOR U68601 ( .A(n53458), .B(n48264), .Z(n49825) );
  XOR U68602 ( .A(n48265), .B(n49825), .Z(n53470) );
  IV U68603 ( .A(n48266), .Z(n48267) );
  NOR U68604 ( .A(n48277), .B(n48267), .Z(n48274) );
  IV U68605 ( .A(n48274), .Z(n53474) );
  NOR U68606 ( .A(n53470), .B(n53474), .Z(n49821) );
  IV U68607 ( .A(n48268), .Z(n48271) );
  IV U68608 ( .A(n48269), .Z(n48270) );
  NOR U68609 ( .A(n48271), .B(n48270), .Z(n48272) );
  IV U68610 ( .A(n48272), .Z(n54988) );
  XOR U68611 ( .A(n53470), .B(n54988), .Z(n48273) );
  NOR U68612 ( .A(n48274), .B(n48273), .Z(n49820) );
  IV U68613 ( .A(n48275), .Z(n48276) );
  NOR U68614 ( .A(n48277), .B(n48276), .Z(n49819) );
  XOR U68615 ( .A(n49820), .B(n49819), .Z(n48278) );
  NOR U68616 ( .A(n49821), .B(n48278), .Z(n48279) );
  IV U68617 ( .A(n48279), .Z(n53480) );
  IV U68618 ( .A(n48280), .Z(n48282) );
  NOR U68619 ( .A(n48282), .B(n48281), .Z(n53478) );
  XOR U68620 ( .A(n53480), .B(n53478), .Z(n49803) );
  IV U68621 ( .A(n48283), .Z(n48284) );
  NOR U68622 ( .A(n48284), .B(n49812), .Z(n48287) );
  NOR U68623 ( .A(n48285), .B(n49804), .Z(n48286) );
  NOR U68624 ( .A(n48287), .B(n48286), .Z(n48288) );
  XOR U68625 ( .A(n49803), .B(n48288), .Z(n53486) );
  XOR U68626 ( .A(n49800), .B(n53486), .Z(n49798) );
  IV U68627 ( .A(n48289), .Z(n48290) );
  NOR U68628 ( .A(n48292), .B(n48290), .Z(n49797) );
  IV U68629 ( .A(n48291), .Z(n48295) );
  XOR U68630 ( .A(n48293), .B(n48292), .Z(n48294) );
  NOR U68631 ( .A(n48295), .B(n48294), .Z(n53484) );
  NOR U68632 ( .A(n49797), .B(n53484), .Z(n48296) );
  XOR U68633 ( .A(n49798), .B(n48296), .Z(n48297) );
  IV U68634 ( .A(n48297), .Z(n49793) );
  IV U68635 ( .A(n48298), .Z(n48301) );
  IV U68636 ( .A(n48299), .Z(n48300) );
  NOR U68637 ( .A(n48301), .B(n48300), .Z(n49791) );
  XOR U68638 ( .A(n49793), .B(n49791), .Z(n49795) );
  XOR U68639 ( .A(n48302), .B(n49795), .Z(n69264) );
  IV U68640 ( .A(n48303), .Z(n48312) );
  IV U68641 ( .A(n48304), .Z(n48305) );
  NOR U68642 ( .A(n48312), .B(n48305), .Z(n49782) );
  IV U68643 ( .A(n48306), .Z(n48308) );
  NOR U68644 ( .A(n48308), .B(n48307), .Z(n49786) );
  NOR U68645 ( .A(n49782), .B(n49786), .Z(n48309) );
  XOR U68646 ( .A(n69264), .B(n48309), .Z(n49779) );
  IV U68647 ( .A(n48310), .Z(n48311) );
  NOR U68648 ( .A(n48312), .B(n48311), .Z(n49784) );
  IV U68649 ( .A(n48313), .Z(n48315) );
  NOR U68650 ( .A(n48315), .B(n48314), .Z(n49780) );
  NOR U68651 ( .A(n49784), .B(n49780), .Z(n48316) );
  XOR U68652 ( .A(n49779), .B(n48316), .Z(n49777) );
  XOR U68653 ( .A(n49776), .B(n49777), .Z(n49774) );
  XOR U68654 ( .A(n49769), .B(n49774), .Z(n48317) );
  XOR U68655 ( .A(n48318), .B(n48317), .Z(n49762) );
  IV U68656 ( .A(n48319), .Z(n48321) );
  IV U68657 ( .A(n48320), .Z(n48323) );
  NOR U68658 ( .A(n48321), .B(n48323), .Z(n53495) );
  NOR U68659 ( .A(n48322), .B(n49763), .Z(n48325) );
  NOR U68660 ( .A(n48324), .B(n48323), .Z(n53490) );
  NOR U68661 ( .A(n48325), .B(n53490), .Z(n48326) );
  IV U68662 ( .A(n48326), .Z(n48327) );
  NOR U68663 ( .A(n53495), .B(n48327), .Z(n48328) );
  XOR U68664 ( .A(n49762), .B(n48328), .Z(n53507) );
  XOR U68665 ( .A(n53493), .B(n53507), .Z(n53501) );
  IV U68666 ( .A(n48329), .Z(n53508) );
  NOR U68667 ( .A(n48330), .B(n53508), .Z(n48333) );
  NOR U68668 ( .A(n48331), .B(n49755), .Z(n48332) );
  NOR U68669 ( .A(n48333), .B(n48332), .Z(n48334) );
  XOR U68670 ( .A(n53501), .B(n48334), .Z(n49747) );
  IV U68671 ( .A(n48335), .Z(n48336) );
  NOR U68672 ( .A(n48336), .B(n48340), .Z(n53522) );
  IV U68673 ( .A(n48337), .Z(n49751) );
  NOR U68674 ( .A(n48338), .B(n49751), .Z(n48342) );
  IV U68675 ( .A(n48339), .Z(n48341) );
  NOR U68676 ( .A(n48341), .B(n48340), .Z(n49748) );
  NOR U68677 ( .A(n48342), .B(n49748), .Z(n48343) );
  IV U68678 ( .A(n48343), .Z(n48344) );
  NOR U68679 ( .A(n53522), .B(n48344), .Z(n48345) );
  XOR U68680 ( .A(n49747), .B(n48345), .Z(n53520) );
  XOR U68681 ( .A(n53519), .B(n53520), .Z(n49746) );
  IV U68682 ( .A(n48346), .Z(n48349) );
  IV U68683 ( .A(n48347), .Z(n48348) );
  NOR U68684 ( .A(n48349), .B(n48348), .Z(n49744) );
  XOR U68685 ( .A(n49746), .B(n49744), .Z(n53532) );
  XOR U68686 ( .A(n53531), .B(n53532), .Z(n53543) );
  NOR U68687 ( .A(n48356), .B(n48350), .Z(n53527) );
  XOR U68688 ( .A(n48351), .B(n48356), .Z(n48352) );
  NOR U68689 ( .A(n48353), .B(n48352), .Z(n53542) );
  IV U68690 ( .A(n48354), .Z(n48355) );
  NOR U68691 ( .A(n48356), .B(n48355), .Z(n49742) );
  NOR U68692 ( .A(n53542), .B(n49742), .Z(n48357) );
  IV U68693 ( .A(n48357), .Z(n48358) );
  NOR U68694 ( .A(n53527), .B(n48358), .Z(n48359) );
  XOR U68695 ( .A(n53543), .B(n48359), .Z(n48360) );
  IV U68696 ( .A(n48360), .Z(n53541) );
  IV U68697 ( .A(n48361), .Z(n54941) );
  NOR U68698 ( .A(n48362), .B(n54941), .Z(n48370) );
  IV U68699 ( .A(n48370), .Z(n48363) );
  NOR U68700 ( .A(n53541), .B(n48363), .Z(n49738) );
  IV U68701 ( .A(n48364), .Z(n48365) );
  NOR U68702 ( .A(n48368), .B(n48365), .Z(n53539) );
  XOR U68703 ( .A(n53539), .B(n53541), .Z(n49741) );
  IV U68704 ( .A(n48366), .Z(n48367) );
  NOR U68705 ( .A(n48368), .B(n48367), .Z(n49739) );
  XOR U68706 ( .A(n49741), .B(n49739), .Z(n54939) );
  IV U68707 ( .A(n54939), .Z(n48369) );
  NOR U68708 ( .A(n48370), .B(n48369), .Z(n48371) );
  NOR U68709 ( .A(n49738), .B(n48371), .Z(n49731) );
  NOR U68710 ( .A(n48372), .B(n60256), .Z(n49736) );
  IV U68711 ( .A(n48373), .Z(n48375) );
  IV U68712 ( .A(n48374), .Z(n48381) );
  NOR U68713 ( .A(n48375), .B(n48381), .Z(n49732) );
  NOR U68714 ( .A(n49736), .B(n49732), .Z(n48376) );
  XOR U68715 ( .A(n49731), .B(n48376), .Z(n54935) );
  IV U68716 ( .A(n48377), .Z(n48378) );
  NOR U68717 ( .A(n48379), .B(n48378), .Z(n54933) );
  IV U68718 ( .A(n48380), .Z(n48382) );
  NOR U68719 ( .A(n48382), .B(n48381), .Z(n58854) );
  NOR U68720 ( .A(n54933), .B(n58854), .Z(n49730) );
  XOR U68721 ( .A(n54935), .B(n49730), .Z(n48383) );
  IV U68722 ( .A(n48383), .Z(n49727) );
  XOR U68723 ( .A(n49726), .B(n49727), .Z(n53552) );
  XOR U68724 ( .A(n53551), .B(n53552), .Z(n53567) );
  IV U68725 ( .A(n48384), .Z(n48385) );
  NOR U68726 ( .A(n48385), .B(n48389), .Z(n53565) );
  IV U68727 ( .A(n48386), .Z(n54925) );
  NOR U68728 ( .A(n54925), .B(n48387), .Z(n53558) );
  IV U68729 ( .A(n48388), .Z(n48390) );
  NOR U68730 ( .A(n48390), .B(n48389), .Z(n49725) );
  NOR U68731 ( .A(n53558), .B(n49725), .Z(n48391) );
  IV U68732 ( .A(n48391), .Z(n48392) );
  NOR U68733 ( .A(n53565), .B(n48392), .Z(n48393) );
  XOR U68734 ( .A(n53567), .B(n48393), .Z(n49721) );
  IV U68735 ( .A(n48394), .Z(n49722) );
  NOR U68736 ( .A(n49722), .B(n48395), .Z(n48399) );
  IV U68737 ( .A(n48396), .Z(n48398) );
  NOR U68738 ( .A(n48398), .B(n48397), .Z(n53568) );
  NOR U68739 ( .A(n48399), .B(n53568), .Z(n48400) );
  XOR U68740 ( .A(n49721), .B(n48400), .Z(n54916) );
  XOR U68741 ( .A(n48401), .B(n54916), .Z(n53588) );
  XOR U68742 ( .A(n53586), .B(n53588), .Z(n49713) );
  XOR U68743 ( .A(n49712), .B(n49713), .Z(n49717) );
  XOR U68744 ( .A(n49715), .B(n49717), .Z(n53603) );
  XOR U68745 ( .A(n48402), .B(n53603), .Z(n53598) );
  XOR U68746 ( .A(n48403), .B(n53598), .Z(n53609) );
  XOR U68747 ( .A(n53608), .B(n53609), .Z(n53613) );
  XOR U68748 ( .A(n53612), .B(n53613), .Z(n58891) );
  XOR U68749 ( .A(n53615), .B(n58891), .Z(n49709) );
  XOR U68750 ( .A(n48404), .B(n49709), .Z(n53626) );
  XOR U68751 ( .A(n48405), .B(n53626), .Z(n53623) );
  XOR U68752 ( .A(n48406), .B(n53623), .Z(n49703) );
  XOR U68753 ( .A(n48407), .B(n49703), .Z(n53642) );
  NOR U68754 ( .A(n53641), .B(n53644), .Z(n48408) );
  XOR U68755 ( .A(n53642), .B(n48408), .Z(n53650) );
  XOR U68756 ( .A(n53648), .B(n53650), .Z(n53651) );
  XOR U68757 ( .A(n53652), .B(n53651), .Z(n48409) );
  NOR U68758 ( .A(n48410), .B(n48409), .Z(n53656) );
  IV U68759 ( .A(n48410), .Z(n48411) );
  NOR U68760 ( .A(n53650), .B(n48411), .Z(n54867) );
  NOR U68761 ( .A(n53656), .B(n54867), .Z(n49697) );
  IV U68762 ( .A(n48412), .Z(n48413) );
  NOR U68763 ( .A(n48413), .B(n48422), .Z(n49696) );
  IV U68764 ( .A(n48414), .Z(n48415) );
  NOR U68765 ( .A(n48418), .B(n48415), .Z(n54862) );
  IV U68766 ( .A(n48416), .Z(n48417) );
  NOR U68767 ( .A(n48418), .B(n48417), .Z(n54870) );
  NOR U68768 ( .A(n54862), .B(n54870), .Z(n48419) );
  IV U68769 ( .A(n48419), .Z(n53654) );
  NOR U68770 ( .A(n49696), .B(n53654), .Z(n48420) );
  XOR U68771 ( .A(n49697), .B(n48420), .Z(n49692) );
  IV U68772 ( .A(n48421), .Z(n48423) );
  NOR U68773 ( .A(n48423), .B(n48422), .Z(n49690) );
  XOR U68774 ( .A(n49692), .B(n49690), .Z(n49695) );
  XOR U68775 ( .A(n49693), .B(n49695), .Z(n54855) );
  IV U68776 ( .A(n48424), .Z(n48425) );
  NOR U68777 ( .A(n48428), .B(n48425), .Z(n54858) );
  IV U68778 ( .A(n48426), .Z(n48427) );
  NOR U68779 ( .A(n48428), .B(n48427), .Z(n54854) );
  NOR U68780 ( .A(n54858), .B(n54854), .Z(n49689) );
  IV U68781 ( .A(n49689), .Z(n48431) );
  NOR U68782 ( .A(n49687), .B(n48431), .Z(n48429) );
  XOR U68783 ( .A(n54855), .B(n48429), .Z(n48430) );
  NOR U68784 ( .A(n48432), .B(n48430), .Z(n48435) );
  XOR U68785 ( .A(n54855), .B(n48431), .Z(n48434) );
  IV U68786 ( .A(n48432), .Z(n48433) );
  NOR U68787 ( .A(n48434), .B(n48433), .Z(n58915) );
  NOR U68788 ( .A(n48435), .B(n58915), .Z(n53660) );
  XOR U68789 ( .A(n53662), .B(n53660), .Z(n53666) );
  XOR U68790 ( .A(n49683), .B(n53666), .Z(n48436) );
  IV U68791 ( .A(n48436), .Z(n49681) );
  XOR U68792 ( .A(n49680), .B(n49681), .Z(n53670) );
  XOR U68793 ( .A(n53669), .B(n53670), .Z(n53673) );
  XOR U68794 ( .A(n53672), .B(n53673), .Z(n49678) );
  IV U68795 ( .A(n48437), .Z(n48440) );
  IV U68796 ( .A(n48438), .Z(n48439) );
  NOR U68797 ( .A(n48440), .B(n48439), .Z(n49676) );
  XOR U68798 ( .A(n49678), .B(n49676), .Z(n54832) );
  NOR U68799 ( .A(n54834), .B(n48441), .Z(n48445) );
  IV U68800 ( .A(n48442), .Z(n48444) );
  IV U68801 ( .A(n48443), .Z(n48448) );
  NOR U68802 ( .A(n48444), .B(n48448), .Z(n60169) );
  NOR U68803 ( .A(n48445), .B(n60169), .Z(n48446) );
  XOR U68804 ( .A(n54832), .B(n48446), .Z(n49671) );
  IV U68805 ( .A(n48447), .Z(n48449) );
  NOR U68806 ( .A(n48449), .B(n48448), .Z(n60164) );
  NOR U68807 ( .A(n48450), .B(n54825), .Z(n49672) );
  NOR U68808 ( .A(n60164), .B(n49672), .Z(n48451) );
  XOR U68809 ( .A(n49671), .B(n48451), .Z(n53691) );
  IV U68810 ( .A(n48452), .Z(n53680) );
  NOR U68811 ( .A(n48453), .B(n53680), .Z(n48456) );
  IV U68812 ( .A(n48454), .Z(n48455) );
  NOR U68813 ( .A(n48455), .B(n48459), .Z(n53690) );
  NOR U68814 ( .A(n48456), .B(n53690), .Z(n48457) );
  XOR U68815 ( .A(n53691), .B(n48457), .Z(n53687) );
  IV U68816 ( .A(n48458), .Z(n48460) );
  NOR U68817 ( .A(n48460), .B(n48459), .Z(n53688) );
  IV U68818 ( .A(n48461), .Z(n48462) );
  NOR U68819 ( .A(n48462), .B(n48465), .Z(n53702) );
  NOR U68820 ( .A(n53688), .B(n53702), .Z(n48463) );
  XOR U68821 ( .A(n53687), .B(n48463), .Z(n53701) );
  IV U68822 ( .A(n48464), .Z(n48466) );
  NOR U68823 ( .A(n48466), .B(n48465), .Z(n53699) );
  XOR U68824 ( .A(n53701), .B(n53699), .Z(n49661) );
  XOR U68825 ( .A(n48467), .B(n49661), .Z(n53714) );
  XOR U68826 ( .A(n48468), .B(n53714), .Z(n53718) );
  XOR U68827 ( .A(n48469), .B(n53718), .Z(n53731) );
  XOR U68828 ( .A(n53727), .B(n53731), .Z(n53736) );
  XOR U68829 ( .A(n48470), .B(n53736), .Z(n53742) );
  XOR U68830 ( .A(n48471), .B(n53742), .Z(n49645) );
  XOR U68831 ( .A(n49648), .B(n49645), .Z(n49643) );
  IV U68832 ( .A(n48472), .Z(n48473) );
  NOR U68833 ( .A(n48474), .B(n48473), .Z(n48475) );
  IV U68834 ( .A(n48475), .Z(n49641) );
  XOR U68835 ( .A(n49643), .B(n49641), .Z(n48476) );
  XOR U68836 ( .A(n48477), .B(n48476), .Z(n54791) );
  IV U68837 ( .A(n54791), .Z(n48483) );
  NOR U68838 ( .A(n48478), .B(n54794), .Z(n49639) );
  IV U68839 ( .A(n48479), .Z(n49633) );
  NOR U68840 ( .A(n48480), .B(n49633), .Z(n48481) );
  NOR U68841 ( .A(n49639), .B(n48481), .Z(n48482) );
  XOR U68842 ( .A(n48483), .B(n48482), .Z(n59009) );
  XOR U68843 ( .A(n49631), .B(n59009), .Z(n48484) );
  XOR U68844 ( .A(n48491), .B(n48484), .Z(n48488) );
  IV U68845 ( .A(n48485), .Z(n48486) );
  NOR U68846 ( .A(n48486), .B(n48497), .Z(n48494) );
  IV U68847 ( .A(n48494), .Z(n48487) );
  NOR U68848 ( .A(n48488), .B(n48487), .Z(n54784) );
  IV U68849 ( .A(n48489), .Z(n48490) );
  NOR U68850 ( .A(n49626), .B(n48490), .Z(n59007) );
  XOR U68851 ( .A(n49631), .B(n48491), .Z(n48492) );
  NOR U68852 ( .A(n59007), .B(n48492), .Z(n48493) );
  XOR U68853 ( .A(n48493), .B(n59009), .Z(n48504) );
  NOR U68854 ( .A(n48494), .B(n48504), .Z(n48495) );
  NOR U68855 ( .A(n54784), .B(n48495), .Z(n53748) );
  IV U68856 ( .A(n48496), .Z(n48498) );
  NOR U68857 ( .A(n48498), .B(n48497), .Z(n48499) );
  IV U68858 ( .A(n48499), .Z(n53749) );
  XOR U68859 ( .A(n53748), .B(n53749), .Z(n54778) );
  IV U68860 ( .A(n54778), .Z(n48503) );
  IV U68861 ( .A(n48500), .Z(n48502) );
  NOR U68862 ( .A(n48502), .B(n48501), .Z(n48505) );
  NOR U68863 ( .A(n48503), .B(n48505), .Z(n48508) );
  IV U68864 ( .A(n48504), .Z(n48507) );
  IV U68865 ( .A(n48505), .Z(n48506) );
  NOR U68866 ( .A(n48507), .B(n48506), .Z(n53752) );
  NOR U68867 ( .A(n48508), .B(n53752), .Z(n48515) );
  IV U68868 ( .A(n48515), .Z(n49621) );
  NOR U68869 ( .A(n48509), .B(n49621), .Z(n59023) );
  IV U68870 ( .A(n48510), .Z(n54781) );
  NOR U68871 ( .A(n54781), .B(n48511), .Z(n49623) );
  IV U68872 ( .A(n48512), .Z(n48514) );
  NOR U68873 ( .A(n48514), .B(n48513), .Z(n49620) );
  NOR U68874 ( .A(n49623), .B(n49620), .Z(n48516) );
  XOR U68875 ( .A(n48516), .B(n48515), .Z(n48529) );
  IV U68876 ( .A(n48529), .Z(n48517) );
  NOR U68877 ( .A(n48518), .B(n48517), .Z(n48519) );
  NOR U68878 ( .A(n59023), .B(n48519), .Z(n48531) );
  IV U68879 ( .A(n48531), .Z(n48524) );
  IV U68880 ( .A(n48520), .Z(n48522) );
  IV U68881 ( .A(n48521), .Z(n48526) );
  NOR U68882 ( .A(n48522), .B(n48526), .Z(n48534) );
  IV U68883 ( .A(n48534), .Z(n48523) );
  NOR U68884 ( .A(n48524), .B(n48523), .Z(n65369) );
  IV U68885 ( .A(n48525), .Z(n48527) );
  NOR U68886 ( .A(n48527), .B(n48526), .Z(n48530) );
  IV U68887 ( .A(n48530), .Z(n48528) );
  NOR U68888 ( .A(n48529), .B(n48528), .Z(n49619) );
  NOR U68889 ( .A(n48531), .B(n48530), .Z(n48532) );
  NOR U68890 ( .A(n49619), .B(n48532), .Z(n48533) );
  NOR U68891 ( .A(n48534), .B(n48533), .Z(n48535) );
  NOR U68892 ( .A(n65369), .B(n48535), .Z(n49617) );
  XOR U68893 ( .A(n48536), .B(n49617), .Z(n53768) );
  XOR U68894 ( .A(n53766), .B(n53768), .Z(n53770) );
  XOR U68895 ( .A(n53769), .B(n53770), .Z(n53778) );
  XOR U68896 ( .A(n53777), .B(n53778), .Z(n49613) );
  XOR U68897 ( .A(n49612), .B(n49613), .Z(n53775) );
  XOR U68898 ( .A(n53774), .B(n53775), .Z(n49610) );
  IV U68899 ( .A(n48537), .Z(n48538) );
  NOR U68900 ( .A(n48541), .B(n48538), .Z(n49608) );
  XOR U68901 ( .A(n49610), .B(n49608), .Z(n53787) );
  IV U68902 ( .A(n48539), .Z(n48540) );
  NOR U68903 ( .A(n48541), .B(n48540), .Z(n53785) );
  XOR U68904 ( .A(n53787), .B(n53785), .Z(n53793) );
  IV U68905 ( .A(n48542), .Z(n49605) );
  NOR U68906 ( .A(n48543), .B(n49605), .Z(n48551) );
  IV U68907 ( .A(n48544), .Z(n48545) );
  NOR U68908 ( .A(n48545), .B(n48547), .Z(n53792) );
  IV U68909 ( .A(n48546), .Z(n48548) );
  NOR U68910 ( .A(n48548), .B(n48547), .Z(n53788) );
  NOR U68911 ( .A(n53792), .B(n53788), .Z(n48549) );
  IV U68912 ( .A(n48549), .Z(n48550) );
  NOR U68913 ( .A(n48551), .B(n48550), .Z(n48552) );
  XOR U68914 ( .A(n53793), .B(n48552), .Z(n48553) );
  IV U68915 ( .A(n48553), .Z(n53797) );
  IV U68916 ( .A(n48554), .Z(n48556) );
  NOR U68917 ( .A(n48556), .B(n48555), .Z(n48565) );
  IV U68918 ( .A(n48565), .Z(n48557) );
  NOR U68919 ( .A(n53797), .B(n48557), .Z(n59058) );
  IV U68920 ( .A(n48558), .Z(n48559) );
  NOR U68921 ( .A(n48559), .B(n48562), .Z(n48560) );
  IV U68922 ( .A(n48560), .Z(n49603) );
  IV U68923 ( .A(n48561), .Z(n48563) );
  NOR U68924 ( .A(n48563), .B(n48562), .Z(n53795) );
  XOR U68925 ( .A(n53795), .B(n53797), .Z(n49602) );
  XOR U68926 ( .A(n49603), .B(n49602), .Z(n48564) );
  NOR U68927 ( .A(n48565), .B(n48564), .Z(n53809) );
  NOR U68928 ( .A(n59058), .B(n53809), .Z(n49600) );
  XOR U68929 ( .A(n48566), .B(n49600), .Z(n53813) );
  XOR U68930 ( .A(n53811), .B(n53813), .Z(n53816) );
  IV U68931 ( .A(n48567), .Z(n48569) );
  NOR U68932 ( .A(n48569), .B(n48568), .Z(n53814) );
  XOR U68933 ( .A(n53816), .B(n53814), .Z(n53820) );
  NOR U68934 ( .A(n53821), .B(n48570), .Z(n49595) );
  IV U68935 ( .A(n48571), .Z(n49589) );
  NOR U68936 ( .A(n48572), .B(n49589), .Z(n48573) );
  NOR U68937 ( .A(n49595), .B(n48573), .Z(n48574) );
  XOR U68938 ( .A(n53820), .B(n48574), .Z(n48583) );
  IV U68939 ( .A(n48583), .Z(n59074) );
  XOR U68940 ( .A(n48581), .B(n59074), .Z(n48578) );
  IV U68941 ( .A(n48575), .Z(n48576) );
  NOR U68942 ( .A(n48576), .B(n48588), .Z(n48585) );
  IV U68943 ( .A(n48585), .Z(n48577) );
  NOR U68944 ( .A(n48578), .B(n48577), .Z(n49576) );
  IV U68945 ( .A(n48579), .Z(n59077) );
  NOR U68946 ( .A(n48580), .B(n59077), .Z(n49577) );
  NOR U68947 ( .A(n48581), .B(n49577), .Z(n48582) );
  XOR U68948 ( .A(n48583), .B(n48582), .Z(n53827) );
  IV U68949 ( .A(n53827), .Z(n48584) );
  NOR U68950 ( .A(n48585), .B(n48584), .Z(n48586) );
  NOR U68951 ( .A(n49576), .B(n48586), .Z(n53831) );
  IV U68952 ( .A(n48587), .Z(n48589) );
  NOR U68953 ( .A(n48589), .B(n48588), .Z(n53826) );
  NOR U68954 ( .A(n48591), .B(n48590), .Z(n48592) );
  IV U68955 ( .A(n48592), .Z(n48594) );
  NOR U68956 ( .A(n48594), .B(n48593), .Z(n53832) );
  NOR U68957 ( .A(n53826), .B(n53832), .Z(n48595) );
  XOR U68958 ( .A(n53831), .B(n48595), .Z(n53842) );
  XOR U68959 ( .A(n53840), .B(n53842), .Z(n53844) );
  XOR U68960 ( .A(n53843), .B(n53844), .Z(n49574) );
  IV U68961 ( .A(n48596), .Z(n48597) );
  NOR U68962 ( .A(n48597), .B(n48602), .Z(n49573) );
  IV U68963 ( .A(n48598), .Z(n48599) );
  NOR U68964 ( .A(n48600), .B(n48599), .Z(n48601) );
  IV U68965 ( .A(n48601), .Z(n48603) );
  NOR U68966 ( .A(n48603), .B(n48602), .Z(n49567) );
  NOR U68967 ( .A(n49573), .B(n49567), .Z(n48604) );
  XOR U68968 ( .A(n49574), .B(n48604), .Z(n48605) );
  IV U68969 ( .A(n48605), .Z(n49571) );
  XOR U68970 ( .A(n49569), .B(n49571), .Z(n53849) );
  XOR U68971 ( .A(n53848), .B(n53849), .Z(n53853) );
  XOR U68972 ( .A(n53851), .B(n53853), .Z(n53855) );
  XOR U68973 ( .A(n53856), .B(n53855), .Z(n48617) );
  IV U68974 ( .A(n48617), .Z(n48606) );
  NOR U68975 ( .A(n48607), .B(n48606), .Z(n59094) );
  IV U68976 ( .A(n48608), .Z(n48611) );
  IV U68977 ( .A(n48609), .Z(n48616) );
  NOR U68978 ( .A(n48616), .B(n53855), .Z(n48610) );
  IV U68979 ( .A(n48610), .Z(n48613) );
  NOR U68980 ( .A(n48611), .B(n48613), .Z(n54692) );
  IV U68981 ( .A(n48612), .Z(n48614) );
  NOR U68982 ( .A(n48614), .B(n48613), .Z(n59091) );
  NOR U68983 ( .A(n48616), .B(n48615), .Z(n48618) );
  NOR U68984 ( .A(n48618), .B(n48617), .Z(n48619) );
  NOR U68985 ( .A(n59091), .B(n48619), .Z(n48620) );
  IV U68986 ( .A(n48620), .Z(n48621) );
  NOR U68987 ( .A(n54692), .B(n48621), .Z(n53862) );
  NOR U68988 ( .A(n48622), .B(n53862), .Z(n48623) );
  NOR U68989 ( .A(n59094), .B(n48623), .Z(n48624) );
  IV U68990 ( .A(n48624), .Z(n53859) );
  XOR U68991 ( .A(n53858), .B(n53859), .Z(n49565) );
  IV U68992 ( .A(n48625), .Z(n53864) );
  NOR U68993 ( .A(n48626), .B(n53864), .Z(n48630) );
  IV U68994 ( .A(n48627), .Z(n48629) );
  NOR U68995 ( .A(n48629), .B(n48628), .Z(n49564) );
  NOR U68996 ( .A(n48630), .B(n49564), .Z(n48631) );
  XOR U68997 ( .A(n49565), .B(n48631), .Z(n49556) );
  XOR U68998 ( .A(n49562), .B(n49556), .Z(n48632) );
  NOR U68999 ( .A(n48633), .B(n48632), .Z(n64338) );
  IV U69000 ( .A(n48634), .Z(n48636) );
  IV U69001 ( .A(n48635), .Z(n48643) );
  NOR U69002 ( .A(n48636), .B(n48643), .Z(n49557) );
  NOR U69003 ( .A(n48637), .B(n49557), .Z(n48638) );
  XOR U69004 ( .A(n48638), .B(n49556), .Z(n49561) );
  IV U69005 ( .A(n48639), .Z(n48640) );
  NOR U69006 ( .A(n48641), .B(n48640), .Z(n49554) );
  IV U69007 ( .A(n48642), .Z(n48644) );
  NOR U69008 ( .A(n48644), .B(n48643), .Z(n49559) );
  NOR U69009 ( .A(n49554), .B(n49559), .Z(n48645) );
  XOR U69010 ( .A(n49561), .B(n48645), .Z(n48646) );
  NOR U69011 ( .A(n48647), .B(n48646), .Z(n48648) );
  NOR U69012 ( .A(n64338), .B(n48648), .Z(n49549) );
  IV U69013 ( .A(n48649), .Z(n48650) );
  NOR U69014 ( .A(n48657), .B(n48650), .Z(n49548) );
  IV U69015 ( .A(n48651), .Z(n48653) );
  NOR U69016 ( .A(n48653), .B(n48652), .Z(n49551) );
  NOR U69017 ( .A(n49548), .B(n49551), .Z(n48654) );
  XOR U69018 ( .A(n49549), .B(n48654), .Z(n54653) );
  IV U69019 ( .A(n48655), .Z(n48656) );
  NOR U69020 ( .A(n48657), .B(n48656), .Z(n54654) );
  IV U69021 ( .A(n48658), .Z(n48661) );
  IV U69022 ( .A(n48659), .Z(n48660) );
  NOR U69023 ( .A(n48661), .B(n48660), .Z(n54647) );
  NOR U69024 ( .A(n54655), .B(n54647), .Z(n53875) );
  IV U69025 ( .A(n53875), .Z(n48662) );
  NOR U69026 ( .A(n54654), .B(n48662), .Z(n48663) );
  XOR U69027 ( .A(n54653), .B(n48663), .Z(n53876) );
  IV U69028 ( .A(n48664), .Z(n48665) );
  NOR U69029 ( .A(n48673), .B(n48665), .Z(n53881) );
  IV U69030 ( .A(n48666), .Z(n48669) );
  IV U69031 ( .A(n48667), .Z(n48668) );
  NOR U69032 ( .A(n48669), .B(n48668), .Z(n53877) );
  NOR U69033 ( .A(n53881), .B(n53877), .Z(n48670) );
  XOR U69034 ( .A(n53876), .B(n48670), .Z(n49540) );
  IV U69035 ( .A(n48671), .Z(n48672) );
  NOR U69036 ( .A(n48673), .B(n48672), .Z(n49539) );
  XOR U69037 ( .A(n49540), .B(n49539), .Z(n49542) );
  XOR U69038 ( .A(n48674), .B(n49542), .Z(n53886) );
  IV U69039 ( .A(n48675), .Z(n48677) );
  IV U69040 ( .A(n48676), .Z(n48679) );
  NOR U69041 ( .A(n48677), .B(n48679), .Z(n54635) );
  IV U69042 ( .A(n48678), .Z(n48680) );
  NOR U69043 ( .A(n48680), .B(n48679), .Z(n59116) );
  NOR U69044 ( .A(n54635), .B(n59116), .Z(n48682) );
  IV U69045 ( .A(n48682), .Z(n48681) );
  NOR U69046 ( .A(n53886), .B(n48681), .Z(n48683) );
  XOR U69047 ( .A(n49541), .B(n49542), .Z(n54637) );
  NOR U69048 ( .A(n48682), .B(n54637), .Z(n53884) );
  NOR U69049 ( .A(n48683), .B(n53884), .Z(n49524) );
  XOR U69050 ( .A(n49523), .B(n49524), .Z(n49521) );
  XOR U69051 ( .A(n48684), .B(n49521), .Z(n48695) );
  IV U69052 ( .A(n48695), .Z(n53898) );
  NOR U69053 ( .A(n48685), .B(n53898), .Z(n49512) );
  IV U69054 ( .A(n48686), .Z(n48691) );
  IV U69055 ( .A(n48687), .Z(n48688) );
  NOR U69056 ( .A(n48691), .B(n48688), .Z(n49513) );
  IV U69057 ( .A(n48689), .Z(n48690) );
  NOR U69058 ( .A(n48691), .B(n48690), .Z(n48696) );
  IV U69059 ( .A(n48696), .Z(n48694) );
  XOR U69060 ( .A(n48692), .B(n49521), .Z(n48693) );
  NOR U69061 ( .A(n48694), .B(n48693), .Z(n59953) );
  NOR U69062 ( .A(n48696), .B(n48695), .Z(n48697) );
  NOR U69063 ( .A(n59953), .B(n48697), .Z(n49514) );
  XOR U69064 ( .A(n49513), .B(n49514), .Z(n48698) );
  NOR U69065 ( .A(n48699), .B(n48698), .Z(n48700) );
  NOR U69066 ( .A(n49512), .B(n48700), .Z(n48701) );
  IV U69067 ( .A(n48701), .Z(n53900) );
  IV U69068 ( .A(n48702), .Z(n48704) );
  NOR U69069 ( .A(n48704), .B(n48703), .Z(n49511) );
  XOR U69070 ( .A(n53900), .B(n49511), .Z(n53906) );
  XOR U69071 ( .A(n48705), .B(n53906), .Z(n48713) );
  NOR U69072 ( .A(n48706), .B(n48713), .Z(n48709) );
  IV U69073 ( .A(n48706), .Z(n48708) );
  XOR U69074 ( .A(n49509), .B(n53906), .Z(n48707) );
  NOR U69075 ( .A(n48708), .B(n48707), .Z(n49506) );
  NOR U69076 ( .A(n48709), .B(n49506), .Z(n48717) );
  IV U69077 ( .A(n48717), .Z(n48710) );
  NOR U69078 ( .A(n48711), .B(n48710), .Z(n54621) );
  IV U69079 ( .A(n48712), .Z(n48715) );
  IV U69080 ( .A(n48713), .Z(n53911) );
  NOR U69081 ( .A(n48715), .B(n53911), .Z(n48714) );
  IV U69082 ( .A(n48714), .Z(n54626) );
  NOR U69083 ( .A(n48716), .B(n54626), .Z(n53917) );
  NOR U69084 ( .A(n48716), .B(n48715), .Z(n48718) );
  NOR U69085 ( .A(n48718), .B(n48717), .Z(n48719) );
  NOR U69086 ( .A(n53917), .B(n48719), .Z(n48728) );
  NOR U69087 ( .A(n48720), .B(n48728), .Z(n48721) );
  NOR U69088 ( .A(n54621), .B(n48721), .Z(n49503) );
  IV U69089 ( .A(n48722), .Z(n48724) );
  NOR U69090 ( .A(n48724), .B(n48723), .Z(n49502) );
  XOR U69091 ( .A(n49503), .B(n49502), .Z(n48735) );
  IV U69092 ( .A(n48735), .Z(n49498) );
  IV U69093 ( .A(n48725), .Z(n48726) );
  NOR U69094 ( .A(n48743), .B(n48726), .Z(n48746) );
  IV U69095 ( .A(n48746), .Z(n48727) );
  NOR U69096 ( .A(n49498), .B(n48727), .Z(n54610) );
  IV U69097 ( .A(n48728), .Z(n48733) );
  IV U69098 ( .A(n48729), .Z(n48731) );
  IV U69099 ( .A(n48730), .Z(n48739) );
  NOR U69100 ( .A(n48731), .B(n48739), .Z(n48734) );
  IV U69101 ( .A(n48734), .Z(n48732) );
  NOR U69102 ( .A(n48733), .B(n48732), .Z(n54616) );
  NOR U69103 ( .A(n48735), .B(n48734), .Z(n48736) );
  NOR U69104 ( .A(n54616), .B(n48736), .Z(n48737) );
  IV U69105 ( .A(n48737), .Z(n49501) );
  IV U69106 ( .A(n48738), .Z(n48740) );
  NOR U69107 ( .A(n48740), .B(n48739), .Z(n49499) );
  IV U69108 ( .A(n48741), .Z(n48742) );
  NOR U69109 ( .A(n48743), .B(n48742), .Z(n49496) );
  NOR U69110 ( .A(n49499), .B(n49496), .Z(n48744) );
  XOR U69111 ( .A(n49501), .B(n48744), .Z(n48745) );
  NOR U69112 ( .A(n48746), .B(n48745), .Z(n48747) );
  NOR U69113 ( .A(n54610), .B(n48747), .Z(n49483) );
  NOR U69114 ( .A(n48749), .B(n48748), .Z(n49493) );
  NOR U69115 ( .A(n49493), .B(n48750), .Z(n48751) );
  XOR U69116 ( .A(n49483), .B(n48751), .Z(n49480) );
  XOR U69117 ( .A(n48752), .B(n49480), .Z(n53926) );
  XOR U69118 ( .A(n53924), .B(n53926), .Z(n53929) );
  IV U69119 ( .A(n48753), .Z(n48754) );
  NOR U69120 ( .A(n48762), .B(n48754), .Z(n49477) );
  IV U69121 ( .A(n48755), .Z(n48757) );
  NOR U69122 ( .A(n48757), .B(n48756), .Z(n53927) );
  NOR U69123 ( .A(n49477), .B(n53927), .Z(n48758) );
  XOR U69124 ( .A(n53929), .B(n48758), .Z(n48759) );
  IV U69125 ( .A(n48759), .Z(n49474) );
  IV U69126 ( .A(n48760), .Z(n48761) );
  NOR U69127 ( .A(n48762), .B(n48761), .Z(n49472) );
  XOR U69128 ( .A(n49474), .B(n49472), .Z(n49470) );
  XOR U69129 ( .A(n48763), .B(n49470), .Z(n48764) );
  IV U69130 ( .A(n48764), .Z(n49465) );
  NOR U69131 ( .A(n48766), .B(n48765), .Z(n48767) );
  IV U69132 ( .A(n48767), .Z(n48769) );
  NOR U69133 ( .A(n48769), .B(n48768), .Z(n49463) );
  XOR U69134 ( .A(n49465), .B(n49463), .Z(n49457) );
  XOR U69135 ( .A(n48770), .B(n49457), .Z(n49448) );
  IV U69136 ( .A(n48771), .Z(n48773) );
  IV U69137 ( .A(n48772), .Z(n48777) );
  NOR U69138 ( .A(n48773), .B(n48777), .Z(n48774) );
  IV U69139 ( .A(n48774), .Z(n48784) );
  NOR U69140 ( .A(n49448), .B(n48784), .Z(n49446) );
  NOR U69141 ( .A(n48775), .B(n49451), .Z(n48779) );
  IV U69142 ( .A(n48776), .Z(n48778) );
  NOR U69143 ( .A(n48778), .B(n48777), .Z(n49447) );
  NOR U69144 ( .A(n48779), .B(n49447), .Z(n48780) );
  XOR U69145 ( .A(n48780), .B(n49448), .Z(n48781) );
  IV U69146 ( .A(n48781), .Z(n53936) );
  IV U69147 ( .A(n48782), .Z(n48783) );
  NOR U69148 ( .A(n48794), .B(n48783), .Z(n48785) );
  IV U69149 ( .A(n48785), .Z(n53935) );
  XOR U69150 ( .A(n53936), .B(n53935), .Z(n48787) );
  NOR U69151 ( .A(n48785), .B(n48784), .Z(n48786) );
  NOR U69152 ( .A(n48787), .B(n48786), .Z(n48788) );
  NOR U69153 ( .A(n49446), .B(n48788), .Z(n49439) );
  IV U69154 ( .A(n48789), .Z(n48791) );
  NOR U69155 ( .A(n48791), .B(n48790), .Z(n48792) );
  IV U69156 ( .A(n48792), .Z(n48793) );
  NOR U69157 ( .A(n48794), .B(n48793), .Z(n48795) );
  IV U69158 ( .A(n48795), .Z(n53937) );
  XOR U69159 ( .A(n49439), .B(n53937), .Z(n49436) );
  NOR U69160 ( .A(n49440), .B(n48796), .Z(n48799) );
  IV U69161 ( .A(n48797), .Z(n48802) );
  NOR U69162 ( .A(n48798), .B(n48802), .Z(n49435) );
  NOR U69163 ( .A(n48799), .B(n49435), .Z(n48800) );
  XOR U69164 ( .A(n49436), .B(n48800), .Z(n49423) );
  IV U69165 ( .A(n48801), .Z(n48803) );
  NOR U69166 ( .A(n48803), .B(n48802), .Z(n48804) );
  IV U69167 ( .A(n48804), .Z(n49430) );
  XOR U69168 ( .A(n49423), .B(n49430), .Z(n49433) );
  XOR U69169 ( .A(n49432), .B(n49433), .Z(n49420) );
  IV U69170 ( .A(n48805), .Z(n48807) );
  NOR U69171 ( .A(n48807), .B(n48806), .Z(n48808) );
  IV U69172 ( .A(n48808), .Z(n49418) );
  XOR U69173 ( .A(n49420), .B(n49418), .Z(n48809) );
  XOR U69174 ( .A(n48810), .B(n48809), .Z(n53947) );
  XOR U69175 ( .A(n48811), .B(n53947), .Z(n65162) );
  XOR U69176 ( .A(n48812), .B(n65162), .Z(n53950) );
  XOR U69177 ( .A(n53949), .B(n53950), .Z(n53973) );
  XOR U69178 ( .A(n48813), .B(n53973), .Z(n49400) );
  NOR U69179 ( .A(n48815), .B(n48814), .Z(n48816) );
  IV U69180 ( .A(n48816), .Z(n48817) );
  NOR U69181 ( .A(n48817), .B(n48821), .Z(n53995) );
  IV U69182 ( .A(n48818), .Z(n49403) );
  NOR U69183 ( .A(n48819), .B(n49403), .Z(n48823) );
  IV U69184 ( .A(n48820), .Z(n48822) );
  NOR U69185 ( .A(n48822), .B(n48821), .Z(n49399) );
  NOR U69186 ( .A(n48823), .B(n49399), .Z(n48824) );
  IV U69187 ( .A(n48824), .Z(n48825) );
  NOR U69188 ( .A(n53995), .B(n48825), .Z(n48826) );
  XOR U69189 ( .A(n49400), .B(n48826), .Z(n49398) );
  IV U69190 ( .A(n48827), .Z(n48829) );
  NOR U69191 ( .A(n48829), .B(n48828), .Z(n48830) );
  IV U69192 ( .A(n48830), .Z(n48831) );
  NOR U69193 ( .A(n48832), .B(n48831), .Z(n49396) );
  XOR U69194 ( .A(n49398), .B(n49396), .Z(n54012) );
  XOR U69195 ( .A(n54013), .B(n54012), .Z(n54022) );
  XOR U69196 ( .A(n48833), .B(n54022), .Z(n48846) );
  IV U69197 ( .A(n48846), .Z(n48837) );
  IV U69198 ( .A(n48834), .Z(n48835) );
  NOR U69199 ( .A(n48835), .B(n48852), .Z(n48849) );
  IV U69200 ( .A(n48849), .Z(n48836) );
  NOR U69201 ( .A(n48837), .B(n48836), .Z(n54543) );
  IV U69202 ( .A(n48838), .Z(n48840) );
  NOR U69203 ( .A(n48840), .B(n48839), .Z(n48841) );
  IV U69204 ( .A(n48841), .Z(n48843) );
  NOR U69205 ( .A(n48843), .B(n48842), .Z(n48845) );
  IV U69206 ( .A(n48845), .Z(n48844) );
  NOR U69207 ( .A(n54022), .B(n48844), .Z(n54554) );
  NOR U69208 ( .A(n48846), .B(n48845), .Z(n48847) );
  NOR U69209 ( .A(n54554), .B(n48847), .Z(n48848) );
  NOR U69210 ( .A(n48849), .B(n48848), .Z(n48850) );
  NOR U69211 ( .A(n54543), .B(n48850), .Z(n49392) );
  IV U69212 ( .A(n48851), .Z(n48853) );
  NOR U69213 ( .A(n48853), .B(n48852), .Z(n54023) );
  IV U69214 ( .A(n48854), .Z(n48855) );
  NOR U69215 ( .A(n48858), .B(n48855), .Z(n49394) );
  IV U69216 ( .A(n48856), .Z(n48857) );
  NOR U69217 ( .A(n48858), .B(n48857), .Z(n49391) );
  NOR U69218 ( .A(n49394), .B(n49391), .Z(n48859) );
  IV U69219 ( .A(n48859), .Z(n48860) );
  NOR U69220 ( .A(n54023), .B(n48860), .Z(n48861) );
  XOR U69221 ( .A(n49392), .B(n48861), .Z(n54030) );
  XOR U69222 ( .A(n54030), .B(n54028), .Z(n54032) );
  XOR U69223 ( .A(n54031), .B(n54032), .Z(n54524) );
  XOR U69224 ( .A(n49388), .B(n54524), .Z(n49385) );
  NOR U69225 ( .A(n54527), .B(n54529), .Z(n48865) );
  IV U69226 ( .A(n48862), .Z(n48864) );
  IV U69227 ( .A(n48863), .Z(n48868) );
  NOR U69228 ( .A(n48864), .B(n48868), .Z(n49383) );
  NOR U69229 ( .A(n48865), .B(n49383), .Z(n48866) );
  XOR U69230 ( .A(n49385), .B(n48866), .Z(n49377) );
  IV U69231 ( .A(n48867), .Z(n48869) );
  NOR U69232 ( .A(n48869), .B(n48868), .Z(n49380) );
  IV U69233 ( .A(n48870), .Z(n48871) );
  NOR U69234 ( .A(n48875), .B(n48871), .Z(n49378) );
  NOR U69235 ( .A(n49380), .B(n49378), .Z(n48872) );
  XOR U69236 ( .A(n49377), .B(n48872), .Z(n49376) );
  IV U69237 ( .A(n48873), .Z(n48874) );
  NOR U69238 ( .A(n48875), .B(n48874), .Z(n49374) );
  XOR U69239 ( .A(n49376), .B(n49374), .Z(n49370) );
  XOR U69240 ( .A(n49369), .B(n49370), .Z(n49372) );
  XOR U69241 ( .A(n49373), .B(n49372), .Z(n48876) );
  NOR U69242 ( .A(n48877), .B(n48876), .Z(n54038) );
  IV U69243 ( .A(n48877), .Z(n48878) );
  NOR U69244 ( .A(n48878), .B(n49370), .Z(n54517) );
  NOR U69245 ( .A(n54038), .B(n54517), .Z(n54041) );
  IV U69246 ( .A(n48879), .Z(n59828) );
  NOR U69247 ( .A(n48880), .B(n59828), .Z(n59318) );
  IV U69248 ( .A(n48881), .Z(n48882) );
  NOR U69249 ( .A(n48882), .B(n48885), .Z(n54040) );
  NOR U69250 ( .A(n59318), .B(n54040), .Z(n48883) );
  XOR U69251 ( .A(n54041), .B(n48883), .Z(n49368) );
  IV U69252 ( .A(n48884), .Z(n48886) );
  NOR U69253 ( .A(n48886), .B(n48885), .Z(n49366) );
  XOR U69254 ( .A(n49368), .B(n49366), .Z(n54046) );
  XOR U69255 ( .A(n54043), .B(n54046), .Z(n49364) );
  XOR U69256 ( .A(n48887), .B(n49364), .Z(n49357) );
  XOR U69257 ( .A(n48888), .B(n49357), .Z(n49347) );
  XOR U69258 ( .A(n49345), .B(n49347), .Z(n49342) );
  IV U69259 ( .A(n48889), .Z(n48890) );
  NOR U69260 ( .A(n48891), .B(n48890), .Z(n49340) );
  XOR U69261 ( .A(n49342), .B(n49340), .Z(n54060) );
  IV U69262 ( .A(n48892), .Z(n48894) );
  NOR U69263 ( .A(n48894), .B(n48893), .Z(n49343) );
  NOR U69264 ( .A(n49343), .B(n49330), .Z(n48895) );
  XOR U69265 ( .A(n54060), .B(n48895), .Z(n49322) );
  IV U69266 ( .A(n48896), .Z(n48897) );
  NOR U69267 ( .A(n48898), .B(n48897), .Z(n48901) );
  IV U69268 ( .A(n48899), .Z(n48900) );
  NOR U69269 ( .A(n48900), .B(n48904), .Z(n49325) );
  NOR U69270 ( .A(n48901), .B(n49325), .Z(n48902) );
  XOR U69271 ( .A(n49322), .B(n48902), .Z(n49320) );
  IV U69272 ( .A(n48903), .Z(n48905) );
  NOR U69273 ( .A(n48905), .B(n48904), .Z(n49323) );
  IV U69274 ( .A(n48906), .Z(n48908) );
  NOR U69275 ( .A(n48908), .B(n48907), .Z(n49319) );
  NOR U69276 ( .A(n49323), .B(n49319), .Z(n48909) );
  XOR U69277 ( .A(n49320), .B(n48909), .Z(n54066) );
  XOR U69278 ( .A(n54067), .B(n54066), .Z(n54070) );
  XOR U69279 ( .A(n48910), .B(n54070), .Z(n48911) );
  NOR U69280 ( .A(n48912), .B(n48911), .Z(n48922) );
  IV U69281 ( .A(n48913), .Z(n48916) );
  XOR U69282 ( .A(n54069), .B(n54070), .Z(n49314) );
  NOR U69283 ( .A(n48914), .B(n49314), .Z(n48915) );
  IV U69284 ( .A(n48915), .Z(n48918) );
  NOR U69285 ( .A(n48916), .B(n48918), .Z(n54468) );
  IV U69286 ( .A(n48917), .Z(n48919) );
  NOR U69287 ( .A(n48919), .B(n48918), .Z(n54465) );
  NOR U69288 ( .A(n54468), .B(n54465), .Z(n48920) );
  IV U69289 ( .A(n48920), .Z(n48921) );
  NOR U69290 ( .A(n48922), .B(n48921), .Z(n49302) );
  NOR U69291 ( .A(n48923), .B(n49303), .Z(n48927) );
  IV U69292 ( .A(n48924), .Z(n48926) );
  NOR U69293 ( .A(n48926), .B(n48925), .Z(n54076) );
  NOR U69294 ( .A(n48927), .B(n54076), .Z(n48928) );
  XOR U69295 ( .A(n49302), .B(n48928), .Z(n54083) );
  XOR U69296 ( .A(n54079), .B(n54083), .Z(n48929) );
  NOR U69297 ( .A(n48930), .B(n48929), .Z(n54448) );
  IV U69298 ( .A(n48931), .Z(n48932) );
  NOR U69299 ( .A(n48932), .B(n48934), .Z(n54081) );
  IV U69300 ( .A(n48933), .Z(n48935) );
  NOR U69301 ( .A(n48935), .B(n48934), .Z(n49299) );
  NOR U69302 ( .A(n54081), .B(n49299), .Z(n48936) );
  IV U69303 ( .A(n48936), .Z(n48937) );
  NOR U69304 ( .A(n48937), .B(n54079), .Z(n48938) );
  XOR U69305 ( .A(n54083), .B(n48938), .Z(n48939) );
  NOR U69306 ( .A(n48940), .B(n48939), .Z(n48941) );
  NOR U69307 ( .A(n54448), .B(n48941), .Z(n49294) );
  IV U69308 ( .A(n48942), .Z(n54442) );
  NOR U69309 ( .A(n54442), .B(n48943), .Z(n49296) );
  IV U69310 ( .A(n48944), .Z(n48946) );
  NOR U69311 ( .A(n48946), .B(n48945), .Z(n49293) );
  NOR U69312 ( .A(n49296), .B(n49293), .Z(n48947) );
  XOR U69313 ( .A(n49294), .B(n48947), .Z(n54089) );
  XOR U69314 ( .A(n54088), .B(n54089), .Z(n54092) );
  XOR U69315 ( .A(n48948), .B(n54092), .Z(n49285) );
  XOR U69316 ( .A(n49289), .B(n49285), .Z(n54099) );
  NOR U69317 ( .A(n49286), .B(n49288), .Z(n48952) );
  IV U69318 ( .A(n48949), .Z(n48951) );
  NOR U69319 ( .A(n48951), .B(n48950), .Z(n54098) );
  NOR U69320 ( .A(n48952), .B(n54098), .Z(n48953) );
  XOR U69321 ( .A(n54099), .B(n48953), .Z(n54095) );
  IV U69322 ( .A(n48954), .Z(n48955) );
  NOR U69323 ( .A(n48955), .B(n48959), .Z(n54102) );
  NOR U69324 ( .A(n54102), .B(n48956), .Z(n48957) );
  XOR U69325 ( .A(n54095), .B(n48957), .Z(n54110) );
  IV U69326 ( .A(n48958), .Z(n48960) );
  NOR U69327 ( .A(n48960), .B(n48959), .Z(n54108) );
  XOR U69328 ( .A(n54110), .B(n54108), .Z(n54112) );
  XOR U69329 ( .A(n54111), .B(n54112), .Z(n54131) );
  XOR U69330 ( .A(n54121), .B(n54131), .Z(n54116) );
  IV U69331 ( .A(n48961), .Z(n48962) );
  NOR U69332 ( .A(n48962), .B(n48967), .Z(n49283) );
  IV U69333 ( .A(n48963), .Z(n48964) );
  NOR U69334 ( .A(n48965), .B(n48964), .Z(n54115) );
  IV U69335 ( .A(n48966), .Z(n48968) );
  NOR U69336 ( .A(n48968), .B(n48967), .Z(n54130) );
  NOR U69337 ( .A(n54115), .B(n54130), .Z(n48969) );
  IV U69338 ( .A(n48969), .Z(n48970) );
  NOR U69339 ( .A(n49283), .B(n48970), .Z(n48971) );
  XOR U69340 ( .A(n54116), .B(n48971), .Z(n54135) );
  IV U69341 ( .A(n48972), .Z(n48974) );
  NOR U69342 ( .A(n48974), .B(n48973), .Z(n48975) );
  IV U69343 ( .A(n48975), .Z(n54134) );
  XOR U69344 ( .A(n54135), .B(n54134), .Z(n49276) );
  XOR U69345 ( .A(n48976), .B(n49276), .Z(n49279) );
  IV U69346 ( .A(n48977), .Z(n48979) );
  NOR U69347 ( .A(n48979), .B(n48978), .Z(n48980) );
  IV U69348 ( .A(n48980), .Z(n49278) );
  XOR U69349 ( .A(n49279), .B(n49278), .Z(n48981) );
  NOR U69350 ( .A(n48982), .B(n48981), .Z(n48986) );
  IV U69351 ( .A(n48982), .Z(n48985) );
  IV U69352 ( .A(n48983), .Z(n54137) );
  XOR U69353 ( .A(n54137), .B(n49276), .Z(n49281) );
  XOR U69354 ( .A(n49280), .B(n49281), .Z(n48984) );
  NOR U69355 ( .A(n48985), .B(n48984), .Z(n59377) );
  NOR U69356 ( .A(n48986), .B(n59377), .Z(n48987) );
  IV U69357 ( .A(n48987), .Z(n49268) );
  XOR U69358 ( .A(n48988), .B(n49268), .Z(n54389) );
  NOR U69359 ( .A(n48989), .B(n49269), .Z(n48992) );
  IV U69360 ( .A(n48990), .Z(n54392) );
  NOR U69361 ( .A(n48991), .B(n54392), .Z(n54146) );
  NOR U69362 ( .A(n48992), .B(n54146), .Z(n48993) );
  XOR U69363 ( .A(n54389), .B(n48993), .Z(n54149) );
  IV U69364 ( .A(n48994), .Z(n48996) );
  IV U69365 ( .A(n48995), .Z(n49009) );
  NOR U69366 ( .A(n48996), .B(n49009), .Z(n54153) );
  IV U69367 ( .A(n48997), .Z(n48998) );
  NOR U69368 ( .A(n48998), .B(n49000), .Z(n54150) );
  IV U69369 ( .A(n48999), .Z(n49001) );
  NOR U69370 ( .A(n49001), .B(n49000), .Z(n54155) );
  NOR U69371 ( .A(n54150), .B(n54155), .Z(n49002) );
  IV U69372 ( .A(n49002), .Z(n49003) );
  NOR U69373 ( .A(n54153), .B(n49003), .Z(n49004) );
  XOR U69374 ( .A(n54149), .B(n49004), .Z(n49262) );
  IV U69375 ( .A(n49005), .Z(n49006) );
  NOR U69376 ( .A(n49007), .B(n49006), .Z(n49255) );
  IV U69377 ( .A(n49008), .Z(n49010) );
  NOR U69378 ( .A(n49010), .B(n49009), .Z(n49260) );
  NOR U69379 ( .A(n49255), .B(n49260), .Z(n49011) );
  XOR U69380 ( .A(n49262), .B(n49011), .Z(n49257) );
  XOR U69381 ( .A(n49259), .B(n49257), .Z(n49254) );
  XOR U69382 ( .A(n49012), .B(n49254), .Z(n49240) );
  NOR U69383 ( .A(n49013), .B(n49244), .Z(n49016) );
  IV U69384 ( .A(n49014), .Z(n49019) );
  NOR U69385 ( .A(n49015), .B(n49019), .Z(n49239) );
  NOR U69386 ( .A(n49016), .B(n49239), .Z(n49017) );
  XOR U69387 ( .A(n49240), .B(n49017), .Z(n49238) );
  IV U69388 ( .A(n49018), .Z(n49020) );
  NOR U69389 ( .A(n49020), .B(n49019), .Z(n49236) );
  XOR U69390 ( .A(n49238), .B(n49236), .Z(n54165) );
  XOR U69391 ( .A(n54164), .B(n54165), .Z(n49022) );
  IV U69392 ( .A(n49022), .Z(n54167) );
  XOR U69393 ( .A(n54166), .B(n54167), .Z(n65004) );
  NOR U69394 ( .A(n49021), .B(n65004), .Z(n54353) );
  IV U69395 ( .A(n49021), .Z(n49029) );
  NOR U69396 ( .A(n54166), .B(n54162), .Z(n49023) );
  XOR U69397 ( .A(n49023), .B(n49022), .Z(n49234) );
  IV U69398 ( .A(n49024), .Z(n49026) );
  NOR U69399 ( .A(n49026), .B(n49025), .Z(n49027) );
  IV U69400 ( .A(n49027), .Z(n49235) );
  XOR U69401 ( .A(n49234), .B(n49235), .Z(n49028) );
  NOR U69402 ( .A(n49029), .B(n49028), .Z(n49030) );
  NOR U69403 ( .A(n54353), .B(n49030), .Z(n49031) );
  IV U69404 ( .A(n49031), .Z(n49232) );
  XOR U69405 ( .A(n49231), .B(n49232), .Z(n54175) );
  IV U69406 ( .A(n49032), .Z(n49034) );
  NOR U69407 ( .A(n49034), .B(n49033), .Z(n54173) );
  XOR U69408 ( .A(n54175), .B(n54173), .Z(n54177) );
  IV U69409 ( .A(n49035), .Z(n49038) );
  IV U69410 ( .A(n49036), .Z(n49037) );
  NOR U69411 ( .A(n49038), .B(n49037), .Z(n49039) );
  IV U69412 ( .A(n49039), .Z(n54176) );
  XOR U69413 ( .A(n54177), .B(n54176), .Z(n49224) );
  NOR U69414 ( .A(n49228), .B(n49040), .Z(n49043) );
  IV U69415 ( .A(n49049), .Z(n49042) );
  IV U69416 ( .A(n49041), .Z(n49048) );
  NOR U69417 ( .A(n49042), .B(n49048), .Z(n49223) );
  NOR U69418 ( .A(n49043), .B(n49223), .Z(n49044) );
  XOR U69419 ( .A(n49224), .B(n49044), .Z(n54185) );
  IV U69420 ( .A(n49045), .Z(n49046) );
  NOR U69421 ( .A(n49046), .B(n49048), .Z(n49221) );
  IV U69422 ( .A(n49047), .Z(n49051) );
  XOR U69423 ( .A(n49049), .B(n49048), .Z(n49050) );
  NOR U69424 ( .A(n49051), .B(n49050), .Z(n54183) );
  NOR U69425 ( .A(n49221), .B(n54183), .Z(n49052) );
  XOR U69426 ( .A(n54185), .B(n49052), .Z(n49211) );
  IV U69427 ( .A(n49053), .Z(n54327) );
  NOR U69428 ( .A(n49054), .B(n54327), .Z(n49219) );
  IV U69429 ( .A(n49055), .Z(n49057) );
  NOR U69430 ( .A(n49057), .B(n49056), .Z(n54186) );
  NOR U69431 ( .A(n49219), .B(n54186), .Z(n49058) );
  XOR U69432 ( .A(n49211), .B(n49058), .Z(n49203) );
  XOR U69433 ( .A(n49059), .B(n49203), .Z(n49201) );
  IV U69434 ( .A(n49060), .Z(n49062) );
  NOR U69435 ( .A(n49062), .B(n49061), .Z(n49197) );
  XOR U69436 ( .A(n49201), .B(n49197), .Z(n49063) );
  XOR U69437 ( .A(n49064), .B(n49063), .Z(n49194) );
  XOR U69438 ( .A(n49065), .B(n49194), .Z(n49190) );
  XOR U69439 ( .A(n49188), .B(n49190), .Z(n49184) );
  IV U69440 ( .A(n49070), .Z(n49066) );
  NOR U69441 ( .A(n49066), .B(n59457), .Z(n49189) );
  XOR U69442 ( .A(n49068), .B(n49067), .Z(n49069) );
  NOR U69443 ( .A(n49070), .B(n49069), .Z(n49073) );
  IV U69444 ( .A(n49071), .Z(n49072) );
  NOR U69445 ( .A(n49073), .B(n49072), .Z(n49185) );
  NOR U69446 ( .A(n49189), .B(n49185), .Z(n49074) );
  XOR U69447 ( .A(n49184), .B(n49074), .Z(n54199) );
  XOR U69448 ( .A(n54192), .B(n54199), .Z(n49075) );
  XOR U69449 ( .A(n49076), .B(n49075), .Z(n49077) );
  IV U69450 ( .A(n49077), .Z(n59481) );
  IV U69451 ( .A(n49078), .Z(n49088) );
  IV U69452 ( .A(n49079), .Z(n49080) );
  NOR U69453 ( .A(n49088), .B(n49080), .Z(n59484) );
  IV U69454 ( .A(n49081), .Z(n49083) );
  NOR U69455 ( .A(n49083), .B(n49082), .Z(n59479) );
  NOR U69456 ( .A(n59484), .B(n59479), .Z(n49183) );
  XOR U69457 ( .A(n59481), .B(n49183), .Z(n49178) );
  IV U69458 ( .A(n49084), .Z(n49085) );
  NOR U69459 ( .A(n49085), .B(n49091), .Z(n49177) );
  IV U69460 ( .A(n49086), .Z(n49087) );
  NOR U69461 ( .A(n49088), .B(n49087), .Z(n49181) );
  NOR U69462 ( .A(n49177), .B(n49181), .Z(n49089) );
  XOR U69463 ( .A(n49178), .B(n49089), .Z(n49176) );
  IV U69464 ( .A(n49090), .Z(n49092) );
  NOR U69465 ( .A(n49092), .B(n49091), .Z(n49174) );
  XOR U69466 ( .A(n49176), .B(n49174), .Z(n54295) );
  XOR U69467 ( .A(n49093), .B(n54295), .Z(n49159) );
  XOR U69468 ( .A(n49094), .B(n49159), .Z(n49157) );
  XOR U69469 ( .A(n49095), .B(n49157), .Z(n49149) );
  XOR U69470 ( .A(n49147), .B(n49149), .Z(n49154) );
  NOR U69471 ( .A(n49096), .B(n49150), .Z(n49099) );
  NOR U69472 ( .A(n49143), .B(n49097), .Z(n49098) );
  NOR U69473 ( .A(n49099), .B(n49098), .Z(n49100) );
  XOR U69474 ( .A(n49154), .B(n49100), .Z(n54219) );
  NOR U69475 ( .A(n49101), .B(n54208), .Z(n49105) );
  IV U69476 ( .A(n49102), .Z(n49104) );
  IV U69477 ( .A(n49103), .Z(n49111) );
  NOR U69478 ( .A(n49104), .B(n49111), .Z(n54218) );
  NOR U69479 ( .A(n49105), .B(n54218), .Z(n49106) );
  XOR U69480 ( .A(n54219), .B(n49106), .Z(n54214) );
  IV U69481 ( .A(n49107), .Z(n49108) );
  NOR U69482 ( .A(n49109), .B(n49108), .Z(n54215) );
  IV U69483 ( .A(n49110), .Z(n49112) );
  NOR U69484 ( .A(n49112), .B(n49111), .Z(n49140) );
  NOR U69485 ( .A(n54215), .B(n49140), .Z(n49113) );
  XOR U69486 ( .A(n54214), .B(n49113), .Z(n54226) );
  XOR U69487 ( .A(n54225), .B(n54226), .Z(n49137) );
  XOR U69488 ( .A(n49136), .B(n49137), .Z(n54235) );
  IV U69489 ( .A(n49114), .Z(n49115) );
  NOR U69490 ( .A(n49118), .B(n49115), .Z(n54233) );
  IV U69491 ( .A(n49116), .Z(n49117) );
  NOR U69492 ( .A(n49118), .B(n49117), .Z(n54223) );
  NOR U69493 ( .A(n54233), .B(n54223), .Z(n49119) );
  XOR U69494 ( .A(n54235), .B(n49119), .Z(n49120) );
  IV U69495 ( .A(n49120), .Z(n54238) );
  XOR U69496 ( .A(n54236), .B(n54238), .Z(n54242) );
  XOR U69497 ( .A(n54240), .B(n54242), .Z(n49132) );
  XOR U69498 ( .A(n49130), .B(n49132), .Z(n49135) );
  XOR U69499 ( .A(n49133), .B(n49135), .Z(n59544) );
  NOR U69500 ( .A(n49122), .B(n49121), .Z(n49123) );
  XOR U69501 ( .A(n49124), .B(n49123), .Z(n54251) );
  NOR U69502 ( .A(n49126), .B(n49125), .Z(n54252) );
  IV U69503 ( .A(n54252), .Z(n49127) );
  NOR U69504 ( .A(n54251), .B(n49127), .Z(n54248) );
  IV U69505 ( .A(n54248), .Z(n49128) );
  NOR U69506 ( .A(n59544), .B(n49128), .Z(n49129) );
  IV U69507 ( .A(n49129), .Z(n54259) );
  IV U69508 ( .A(n49130), .Z(n49131) );
  NOR U69509 ( .A(n49132), .B(n49131), .Z(n54261) );
  IV U69510 ( .A(n49133), .Z(n49134) );
  NOR U69511 ( .A(n49135), .B(n49134), .Z(n59547) );
  NOR U69512 ( .A(n54261), .B(n59547), .Z(n54243) );
  IV U69513 ( .A(n49136), .Z(n49138) );
  NOR U69514 ( .A(n49138), .B(n49137), .Z(n49139) );
  IV U69515 ( .A(n49139), .Z(n54228) );
  IV U69516 ( .A(n49140), .Z(n49141) );
  NOR U69517 ( .A(n49141), .B(n54219), .Z(n59531) );
  IV U69518 ( .A(n49142), .Z(n49145) );
  NOR U69519 ( .A(n49143), .B(n49154), .Z(n49144) );
  IV U69520 ( .A(n49144), .Z(n54205) );
  NOR U69521 ( .A(n49145), .B(n54205), .Z(n49146) );
  IV U69522 ( .A(n49146), .Z(n54278) );
  IV U69523 ( .A(n49147), .Z(n49148) );
  NOR U69524 ( .A(n49149), .B(n49148), .Z(n59519) );
  IV U69525 ( .A(n49150), .Z(n49152) );
  NOR U69526 ( .A(n49152), .B(n49151), .Z(n49153) );
  IV U69527 ( .A(n49153), .Z(n49155) );
  NOR U69528 ( .A(n49155), .B(n49154), .Z(n54283) );
  NOR U69529 ( .A(n59519), .B(n54283), .Z(n54203) );
  IV U69530 ( .A(n49156), .Z(n49158) );
  NOR U69531 ( .A(n49158), .B(n49157), .Z(n59516) );
  NOR U69532 ( .A(n54285), .B(n59503), .Z(n49160) );
  IV U69533 ( .A(n49159), .Z(n54287) );
  NOR U69534 ( .A(n49160), .B(n54287), .Z(n54202) );
  IV U69535 ( .A(n49161), .Z(n49162) );
  NOR U69536 ( .A(n54287), .B(n49162), .Z(n59508) );
  IV U69537 ( .A(n49163), .Z(n49164) );
  NOR U69538 ( .A(n54287), .B(n49164), .Z(n54290) );
  IV U69539 ( .A(n49165), .Z(n49166) );
  NOR U69540 ( .A(n49166), .B(n54295), .Z(n54201) );
  IV U69541 ( .A(n49167), .Z(n49170) );
  NOR U69542 ( .A(n49168), .B(n49176), .Z(n49169) );
  IV U69543 ( .A(n49169), .Z(n49172) );
  NOR U69544 ( .A(n49170), .B(n49172), .Z(n59495) );
  IV U69545 ( .A(n49171), .Z(n49173) );
  NOR U69546 ( .A(n49173), .B(n49172), .Z(n59492) );
  IV U69547 ( .A(n49174), .Z(n49175) );
  NOR U69548 ( .A(n49176), .B(n49175), .Z(n54301) );
  IV U69549 ( .A(n49177), .Z(n49180) );
  IV U69550 ( .A(n49178), .Z(n49179) );
  NOR U69551 ( .A(n49180), .B(n49179), .Z(n59476) );
  IV U69552 ( .A(n49181), .Z(n49182) );
  NOR U69553 ( .A(n59481), .B(n49182), .Z(n59472) );
  NOR U69554 ( .A(n59481), .B(n49183), .Z(n54200) );
  IV U69555 ( .A(n49184), .Z(n49187) );
  IV U69556 ( .A(n49185), .Z(n49186) );
  NOR U69557 ( .A(n49187), .B(n49186), .Z(n54305) );
  NOR U69558 ( .A(n49188), .B(n49190), .Z(n59453) );
  IV U69559 ( .A(n49189), .Z(n49191) );
  NOR U69560 ( .A(n49191), .B(n49190), .Z(n59460) );
  XOR U69561 ( .A(n59453), .B(n59460), .Z(n49192) );
  NOR U69562 ( .A(n54305), .B(n49192), .Z(n54191) );
  IV U69563 ( .A(n49193), .Z(n54314) );
  IV U69564 ( .A(n49194), .Z(n69928) );
  NOR U69565 ( .A(n54314), .B(n69928), .Z(n54190) );
  IV U69566 ( .A(n49195), .Z(n49196) );
  NOR U69567 ( .A(n69928), .B(n49196), .Z(n59447) );
  IV U69568 ( .A(n49197), .Z(n49198) );
  NOR U69569 ( .A(n49201), .B(n49198), .Z(n54315) );
  IV U69570 ( .A(n49199), .Z(n49200) );
  NOR U69571 ( .A(n49201), .B(n49200), .Z(n59441) );
  IV U69572 ( .A(n49202), .Z(n49206) );
  NOR U69573 ( .A(n49204), .B(n49203), .Z(n49205) );
  IV U69574 ( .A(n49205), .Z(n49208) );
  NOR U69575 ( .A(n49206), .B(n49208), .Z(n59438) );
  IV U69576 ( .A(n49207), .Z(n49209) );
  NOR U69577 ( .A(n49209), .B(n49208), .Z(n59427) );
  IV U69578 ( .A(n49210), .Z(n49215) );
  IV U69579 ( .A(n49211), .Z(n54323) );
  XOR U69580 ( .A(n54186), .B(n54323), .Z(n49212) );
  NOR U69581 ( .A(n49213), .B(n49212), .Z(n49214) );
  IV U69582 ( .A(n49214), .Z(n49217) );
  NOR U69583 ( .A(n49215), .B(n49217), .Z(n54318) );
  IV U69584 ( .A(n49216), .Z(n49218) );
  NOR U69585 ( .A(n49218), .B(n49217), .Z(n59430) );
  IV U69586 ( .A(n49219), .Z(n49220) );
  NOR U69587 ( .A(n49220), .B(n54323), .Z(n54189) );
  IV U69588 ( .A(n49221), .Z(n49222) );
  NOR U69589 ( .A(n54185), .B(n49222), .Z(n54339) );
  IV U69590 ( .A(n49223), .Z(n49225) );
  IV U69591 ( .A(n49224), .Z(n49227) );
  NOR U69592 ( .A(n49225), .B(n49227), .Z(n54341) );
  NOR U69593 ( .A(n54339), .B(n54341), .Z(n54182) );
  IV U69594 ( .A(n49226), .Z(n49230) );
  NOR U69595 ( .A(n49228), .B(n49227), .Z(n49229) );
  IV U69596 ( .A(n49229), .Z(n54180) );
  NOR U69597 ( .A(n49230), .B(n54180), .Z(n59422) );
  IV U69598 ( .A(n49231), .Z(n49233) );
  NOR U69599 ( .A(n49233), .B(n49232), .Z(n54351) );
  NOR U69600 ( .A(n54353), .B(n54351), .Z(n54172) );
  NOR U69601 ( .A(n49235), .B(n49234), .Z(n54355) );
  IV U69602 ( .A(n49236), .Z(n49237) );
  NOR U69603 ( .A(n49238), .B(n49237), .Z(n54368) );
  IV U69604 ( .A(n49239), .Z(n49241) );
  IV U69605 ( .A(n49240), .Z(n49243) );
  NOR U69606 ( .A(n49241), .B(n49243), .Z(n54366) );
  NOR U69607 ( .A(n54368), .B(n54366), .Z(n54161) );
  IV U69608 ( .A(n49242), .Z(n49246) );
  NOR U69609 ( .A(n49244), .B(n49243), .Z(n49245) );
  IV U69610 ( .A(n49245), .Z(n49248) );
  NOR U69611 ( .A(n49246), .B(n49248), .Z(n59406) );
  IV U69612 ( .A(n49247), .Z(n49249) );
  NOR U69613 ( .A(n49249), .B(n49248), .Z(n54372) );
  IV U69614 ( .A(n49250), .Z(n49251) );
  NOR U69615 ( .A(n49254), .B(n49251), .Z(n59409) );
  IV U69616 ( .A(n49252), .Z(n49253) );
  NOR U69617 ( .A(n49254), .B(n49253), .Z(n54377) );
  NOR U69618 ( .A(n59409), .B(n54377), .Z(n54160) );
  IV U69619 ( .A(n49255), .Z(n49256) );
  NOR U69620 ( .A(n49256), .B(n49262), .Z(n59403) );
  IV U69621 ( .A(n49257), .Z(n49258) );
  NOR U69622 ( .A(n49259), .B(n49258), .Z(n54379) );
  NOR U69623 ( .A(n59403), .B(n54379), .Z(n54159) );
  IV U69624 ( .A(n49260), .Z(n49261) );
  NOR U69625 ( .A(n49262), .B(n49261), .Z(n59399) );
  IV U69626 ( .A(n49263), .Z(n49266) );
  NOR U69627 ( .A(n49264), .B(n49268), .Z(n49265) );
  IV U69628 ( .A(n49265), .Z(n49273) );
  NOR U69629 ( .A(n49266), .B(n49273), .Z(n59729) );
  IV U69630 ( .A(n49267), .Z(n49271) );
  NOR U69631 ( .A(n49269), .B(n49268), .Z(n49270) );
  IV U69632 ( .A(n49270), .Z(n54143) );
  NOR U69633 ( .A(n49271), .B(n54143), .Z(n59725) );
  NOR U69634 ( .A(n59729), .B(n59725), .Z(n59384) );
  IV U69635 ( .A(n49272), .Z(n49274) );
  NOR U69636 ( .A(n49274), .B(n49273), .Z(n54399) );
  NOR U69637 ( .A(n59377), .B(n54399), .Z(n54141) );
  IV U69638 ( .A(n49275), .Z(n49277) );
  IV U69639 ( .A(n49276), .Z(n54136) );
  NOR U69640 ( .A(n49277), .B(n54136), .Z(n54404) );
  NOR U69641 ( .A(n49279), .B(n49278), .Z(n59380) );
  NOR U69642 ( .A(n54404), .B(n59380), .Z(n54140) );
  IV U69643 ( .A(n49280), .Z(n49282) );
  NOR U69644 ( .A(n49282), .B(n49281), .Z(n54401) );
  IV U69645 ( .A(n49283), .Z(n49284) );
  NOR U69646 ( .A(n54131), .B(n49284), .Z(n59374) );
  IV U69647 ( .A(n49285), .Z(n49290) );
  NOR U69648 ( .A(n49286), .B(n49290), .Z(n49287) );
  IV U69649 ( .A(n49287), .Z(n59753) );
  NOR U69650 ( .A(n49288), .B(n59753), .Z(n54420) );
  NOR U69651 ( .A(n49290), .B(n49289), .Z(n59756) );
  IV U69652 ( .A(n49291), .Z(n49292) );
  NOR U69653 ( .A(n54089), .B(n49292), .Z(n64586) );
  NOR U69654 ( .A(n59756), .B(n64586), .Z(n54427) );
  IV U69655 ( .A(n49293), .Z(n49295) );
  IV U69656 ( .A(n49294), .Z(n54439) );
  NOR U69657 ( .A(n49295), .B(n54439), .Z(n54435) );
  IV U69658 ( .A(n49296), .Z(n49297) );
  NOR U69659 ( .A(n49297), .B(n54439), .Z(n49298) );
  IV U69660 ( .A(n49298), .Z(n54087) );
  IV U69661 ( .A(n49299), .Z(n49300) );
  NOR U69662 ( .A(n54083), .B(n49300), .Z(n54452) );
  NOR U69663 ( .A(n54448), .B(n54452), .Z(n54085) );
  IV U69664 ( .A(n49301), .Z(n49305) );
  IV U69665 ( .A(n49302), .Z(n54077) );
  NOR U69666 ( .A(n49303), .B(n54077), .Z(n49304) );
  IV U69667 ( .A(n49304), .Z(n49307) );
  NOR U69668 ( .A(n49305), .B(n49307), .Z(n54460) );
  IV U69669 ( .A(n49306), .Z(n49308) );
  NOR U69670 ( .A(n49308), .B(n49307), .Z(n54463) );
  NOR U69671 ( .A(n54468), .B(n54463), .Z(n54074) );
  IV U69672 ( .A(n49309), .Z(n49310) );
  NOR U69673 ( .A(n49310), .B(n54070), .Z(n49311) );
  IV U69674 ( .A(n49311), .Z(n49312) );
  NOR U69675 ( .A(n49313), .B(n49312), .Z(n54471) );
  IV U69676 ( .A(n49313), .Z(n49318) );
  NOR U69677 ( .A(n49315), .B(n49314), .Z(n49316) );
  IV U69678 ( .A(n49316), .Z(n49317) );
  NOR U69679 ( .A(n49318), .B(n49317), .Z(n54476) );
  IV U69680 ( .A(n49319), .Z(n49321) );
  NOR U69681 ( .A(n49321), .B(n49320), .Z(n54479) );
  IV U69682 ( .A(n49322), .Z(n49327) );
  IV U69683 ( .A(n49323), .Z(n49324) );
  NOR U69684 ( .A(n49327), .B(n49324), .Z(n54485) );
  IV U69685 ( .A(n49325), .Z(n49326) );
  NOR U69686 ( .A(n49327), .B(n49326), .Z(n49328) );
  IV U69687 ( .A(n49328), .Z(n54488) );
  IV U69688 ( .A(n49329), .Z(n49335) );
  XOR U69689 ( .A(n49343), .B(n54060), .Z(n49338) );
  NOR U69690 ( .A(n49330), .B(n49338), .Z(n49331) );
  IV U69691 ( .A(n49331), .Z(n49332) );
  NOR U69692 ( .A(n49333), .B(n49332), .Z(n49334) );
  IV U69693 ( .A(n49334), .Z(n54063) );
  NOR U69694 ( .A(n49335), .B(n54063), .Z(n49336) );
  IV U69695 ( .A(n49336), .Z(n59352) );
  IV U69696 ( .A(n49337), .Z(n49339) );
  NOR U69697 ( .A(n49339), .B(n49338), .Z(n54490) );
  IV U69698 ( .A(n49340), .Z(n49341) );
  NOR U69699 ( .A(n49342), .B(n49341), .Z(n54493) );
  IV U69700 ( .A(n49343), .Z(n49344) );
  NOR U69701 ( .A(n49344), .B(n54060), .Z(n59340) );
  NOR U69702 ( .A(n54493), .B(n59340), .Z(n54057) );
  IV U69703 ( .A(n49345), .Z(n49346) );
  NOR U69704 ( .A(n49347), .B(n49346), .Z(n54496) );
  IV U69705 ( .A(n49348), .Z(n49351) );
  NOR U69706 ( .A(n49357), .B(n49349), .Z(n49350) );
  IV U69707 ( .A(n49350), .Z(n49359) );
  NOR U69708 ( .A(n49351), .B(n49359), .Z(n54498) );
  NOR U69709 ( .A(n54496), .B(n54498), .Z(n54056) );
  IV U69710 ( .A(n49352), .Z(n49354) );
  NOR U69711 ( .A(n49354), .B(n49353), .Z(n49355) );
  IV U69712 ( .A(n49355), .Z(n49356) );
  NOR U69713 ( .A(n49357), .B(n49356), .Z(n54506) );
  IV U69714 ( .A(n49358), .Z(n49360) );
  NOR U69715 ( .A(n49360), .B(n49359), .Z(n54501) );
  NOR U69716 ( .A(n54506), .B(n54501), .Z(n54055) );
  IV U69717 ( .A(n49361), .Z(n49362) );
  NOR U69718 ( .A(n49362), .B(n49364), .Z(n54503) );
  IV U69719 ( .A(n49363), .Z(n49365) );
  NOR U69720 ( .A(n49365), .B(n49364), .Z(n54509) );
  IV U69721 ( .A(n49366), .Z(n49367) );
  NOR U69722 ( .A(n49368), .B(n49367), .Z(n59313) );
  IV U69723 ( .A(n49369), .Z(n49371) );
  NOR U69724 ( .A(n49371), .B(n49370), .Z(n59836) );
  NOR U69725 ( .A(n49373), .B(n49372), .Z(n59831) );
  NOR U69726 ( .A(n59836), .B(n59831), .Z(n54516) );
  IV U69727 ( .A(n54516), .Z(n54036) );
  IV U69728 ( .A(n49374), .Z(n49375) );
  NOR U69729 ( .A(n49376), .B(n49375), .Z(n59307) );
  IV U69730 ( .A(n49377), .Z(n49382) );
  IV U69731 ( .A(n49378), .Z(n49379) );
  NOR U69732 ( .A(n49382), .B(n49379), .Z(n59304) );
  IV U69733 ( .A(n49380), .Z(n49381) );
  NOR U69734 ( .A(n49382), .B(n49381), .Z(n54520) );
  IV U69735 ( .A(n49383), .Z(n49384) );
  NOR U69736 ( .A(n49385), .B(n49384), .Z(n59291) );
  NOR U69737 ( .A(n54524), .B(n54527), .Z(n49386) );
  IV U69738 ( .A(n49386), .Z(n49387) );
  NOR U69739 ( .A(n54529), .B(n49387), .Z(n54035) );
  IV U69740 ( .A(n49388), .Z(n49389) );
  NOR U69741 ( .A(n49389), .B(n54524), .Z(n49390) );
  IV U69742 ( .A(n49390), .Z(n54534) );
  IV U69743 ( .A(n49391), .Z(n49393) );
  IV U69744 ( .A(n49392), .Z(n54025) );
  NOR U69745 ( .A(n49393), .B(n54025), .Z(n54538) );
  IV U69746 ( .A(n49394), .Z(n49395) );
  NOR U69747 ( .A(n49395), .B(n54025), .Z(n54547) );
  NOR U69748 ( .A(n54538), .B(n54547), .Z(n54027) );
  IV U69749 ( .A(n49396), .Z(n49397) );
  NOR U69750 ( .A(n49398), .B(n49397), .Z(n54000) );
  IV U69751 ( .A(n54000), .Z(n53994) );
  IV U69752 ( .A(n49399), .Z(n49401) );
  IV U69753 ( .A(n49400), .Z(n53996) );
  NOR U69754 ( .A(n49401), .B(n53996), .Z(n54574) );
  IV U69755 ( .A(n49402), .Z(n49406) );
  XOR U69756 ( .A(n53974), .B(n53973), .Z(n49404) );
  NOR U69757 ( .A(n49404), .B(n49403), .Z(n49405) );
  IV U69758 ( .A(n49405), .Z(n53991) );
  NOR U69759 ( .A(n49406), .B(n53991), .Z(n53985) );
  IV U69760 ( .A(n49407), .Z(n49410) );
  NOR U69761 ( .A(n49408), .B(n53950), .Z(n49409) );
  IV U69762 ( .A(n49409), .Z(n53966) );
  NOR U69763 ( .A(n49410), .B(n53966), .Z(n59273) );
  IV U69764 ( .A(n49411), .Z(n49412) );
  NOR U69765 ( .A(n65162), .B(n49412), .Z(n59260) );
  IV U69766 ( .A(n53956), .Z(n49413) );
  NOR U69767 ( .A(n65162), .B(n49413), .Z(n59256) );
  IV U69768 ( .A(n49414), .Z(n49415) );
  NOR U69769 ( .A(n53947), .B(n49415), .Z(n59253) );
  IV U69770 ( .A(n49416), .Z(n49417) );
  NOR U69771 ( .A(n53947), .B(n49417), .Z(n59249) );
  NOR U69772 ( .A(n49420), .B(n49418), .Z(n59239) );
  IV U69773 ( .A(n49419), .Z(n49421) );
  NOR U69774 ( .A(n49421), .B(n49420), .Z(n59235) );
  IV U69775 ( .A(n49422), .Z(n49426) );
  IV U69776 ( .A(n49423), .Z(n49431) );
  NOR U69777 ( .A(n49424), .B(n49431), .Z(n49425) );
  IV U69778 ( .A(n49425), .Z(n49428) );
  NOR U69779 ( .A(n49426), .B(n49428), .Z(n59232) );
  IV U69780 ( .A(n49427), .Z(n49429) );
  NOR U69781 ( .A(n49429), .B(n49428), .Z(n59227) );
  NOR U69782 ( .A(n49431), .B(n49430), .Z(n59219) );
  IV U69783 ( .A(n49432), .Z(n49434) );
  NOR U69784 ( .A(n49434), .B(n49433), .Z(n54579) );
  NOR U69785 ( .A(n59219), .B(n54579), .Z(n53941) );
  IV U69786 ( .A(n49435), .Z(n49437) );
  NOR U69787 ( .A(n49437), .B(n49436), .Z(n59216) );
  IV U69788 ( .A(n49438), .Z(n49442) );
  IV U69789 ( .A(n49439), .Z(n53938) );
  NOR U69790 ( .A(n49440), .B(n53938), .Z(n49441) );
  IV U69791 ( .A(n49441), .Z(n49444) );
  NOR U69792 ( .A(n49442), .B(n49444), .Z(n59213) );
  IV U69793 ( .A(n49443), .Z(n49445) );
  NOR U69794 ( .A(n49445), .B(n49444), .Z(n54582) );
  IV U69795 ( .A(n49446), .Z(n54590) );
  IV U69796 ( .A(n49447), .Z(n49449) );
  NOR U69797 ( .A(n49449), .B(n49448), .Z(n54594) );
  IV U69798 ( .A(n49450), .Z(n49453) );
  NOR U69799 ( .A(n49451), .B(n49457), .Z(n49452) );
  IV U69800 ( .A(n49452), .Z(n49455) );
  NOR U69801 ( .A(n49453), .B(n49455), .Z(n54596) );
  NOR U69802 ( .A(n54594), .B(n54596), .Z(n53934) );
  IV U69803 ( .A(n49454), .Z(n49456) );
  NOR U69804 ( .A(n49456), .B(n49455), .Z(n59202) );
  NOR U69805 ( .A(n49458), .B(n49457), .Z(n49459) );
  IV U69806 ( .A(n49459), .Z(n59199) );
  NOR U69807 ( .A(n49460), .B(n59199), .Z(n53933) );
  IV U69808 ( .A(n49461), .Z(n49462) );
  NOR U69809 ( .A(n49462), .B(n49470), .Z(n59191) );
  IV U69810 ( .A(n49463), .Z(n49464) );
  NOR U69811 ( .A(n49465), .B(n49464), .Z(n59194) );
  NOR U69812 ( .A(n59191), .B(n59194), .Z(n53932) );
  IV U69813 ( .A(n49466), .Z(n49468) );
  XOR U69814 ( .A(n49469), .B(n49470), .Z(n49467) );
  NOR U69815 ( .A(n49468), .B(n49467), .Z(n59187) );
  IV U69816 ( .A(n49469), .Z(n49471) );
  NOR U69817 ( .A(n49471), .B(n49470), .Z(n59178) );
  IV U69818 ( .A(n49472), .Z(n49473) );
  NOR U69819 ( .A(n49474), .B(n49473), .Z(n59183) );
  NOR U69820 ( .A(n59178), .B(n59183), .Z(n49475) );
  IV U69821 ( .A(n49475), .Z(n49476) );
  NOR U69822 ( .A(n59187), .B(n49476), .Z(n53931) );
  IV U69823 ( .A(n49477), .Z(n49478) );
  NOR U69824 ( .A(n53929), .B(n49478), .Z(n59180) );
  IV U69825 ( .A(n49479), .Z(n49481) );
  NOR U69826 ( .A(n49481), .B(n49480), .Z(n59171) );
  IV U69827 ( .A(n49482), .Z(n49486) );
  IV U69828 ( .A(n49483), .Z(n49494) );
  XOR U69829 ( .A(n49493), .B(n49494), .Z(n49490) );
  NOR U69830 ( .A(n49484), .B(n49490), .Z(n49485) );
  IV U69831 ( .A(n49485), .Z(n53922) );
  NOR U69832 ( .A(n49486), .B(n53922), .Z(n54599) );
  IV U69833 ( .A(n49487), .Z(n49488) );
  NOR U69834 ( .A(n49488), .B(n49494), .Z(n59166) );
  IV U69835 ( .A(n49489), .Z(n49491) );
  NOR U69836 ( .A(n49491), .B(n49490), .Z(n49492) );
  IV U69837 ( .A(n49492), .Z(n59164) );
  IV U69838 ( .A(n49493), .Z(n49495) );
  NOR U69839 ( .A(n49495), .B(n49494), .Z(n54605) );
  NOR U69840 ( .A(n54610), .B(n54605), .Z(n53920) );
  IV U69841 ( .A(n49496), .Z(n49497) );
  NOR U69842 ( .A(n49498), .B(n49497), .Z(n54607) );
  IV U69843 ( .A(n49499), .Z(n49500) );
  NOR U69844 ( .A(n49501), .B(n49500), .Z(n54614) );
  NOR U69845 ( .A(n54616), .B(n54614), .Z(n53919) );
  IV U69846 ( .A(n49502), .Z(n49505) );
  IV U69847 ( .A(n49503), .Z(n49504) );
  NOR U69848 ( .A(n49505), .B(n49504), .Z(n54619) );
  NOR U69849 ( .A(n54621), .B(n54619), .Z(n53918) );
  IV U69850 ( .A(n49506), .Z(n49507) );
  NOR U69851 ( .A(n53908), .B(n49507), .Z(n49508) );
  IV U69852 ( .A(n49508), .Z(n59156) );
  IV U69853 ( .A(n49509), .Z(n49510) );
  NOR U69854 ( .A(n49510), .B(n53906), .Z(n59140) );
  IV U69855 ( .A(n49511), .Z(n53899) );
  IV U69856 ( .A(n49512), .Z(n59136) );
  IV U69857 ( .A(n49513), .Z(n49516) );
  IV U69858 ( .A(n49514), .Z(n49515) );
  NOR U69859 ( .A(n49516), .B(n49515), .Z(n59946) );
  NOR U69860 ( .A(n59953), .B(n59946), .Z(n59134) );
  IV U69861 ( .A(n59134), .Z(n53894) );
  IV U69862 ( .A(n49517), .Z(n49518) );
  NOR U69863 ( .A(n49521), .B(n49518), .Z(n54629) );
  IV U69864 ( .A(n49519), .Z(n49520) );
  NOR U69865 ( .A(n49521), .B(n49520), .Z(n54632) );
  IV U69866 ( .A(n49522), .Z(n49528) );
  IV U69867 ( .A(n49523), .Z(n49525) );
  IV U69868 ( .A(n49524), .Z(n49530) );
  NOR U69869 ( .A(n49525), .B(n49530), .Z(n49526) );
  IV U69870 ( .A(n49526), .Z(n49527) );
  NOR U69871 ( .A(n49528), .B(n49527), .Z(n59130) );
  IV U69872 ( .A(n49529), .Z(n49531) );
  NOR U69873 ( .A(n49531), .B(n49530), .Z(n59127) );
  IV U69874 ( .A(n49532), .Z(n49535) );
  NOR U69875 ( .A(n49533), .B(n49542), .Z(n49534) );
  IV U69876 ( .A(n49534), .Z(n49537) );
  NOR U69877 ( .A(n49535), .B(n49537), .Z(n59113) );
  IV U69878 ( .A(n49536), .Z(n49538) );
  NOR U69879 ( .A(n49538), .B(n49537), .Z(n59106) );
  IV U69880 ( .A(n49539), .Z(n54640) );
  NOR U69881 ( .A(n49540), .B(n54640), .Z(n49544) );
  IV U69882 ( .A(n49541), .Z(n49543) );
  NOR U69883 ( .A(n49543), .B(n49542), .Z(n59109) );
  NOR U69884 ( .A(n49544), .B(n59109), .Z(n49545) );
  IV U69885 ( .A(n49545), .Z(n53883) );
  IV U69886 ( .A(n54654), .Z(n49546) );
  NOR U69887 ( .A(n54653), .B(n49546), .Z(n49547) );
  IV U69888 ( .A(n49547), .Z(n54665) );
  IV U69889 ( .A(n49548), .Z(n49550) );
  IV U69890 ( .A(n49549), .Z(n49553) );
  NOR U69891 ( .A(n49550), .B(n49553), .Z(n54661) );
  IV U69892 ( .A(n49551), .Z(n49552) );
  NOR U69893 ( .A(n49553), .B(n49552), .Z(n64343) );
  NOR U69894 ( .A(n64338), .B(n64343), .Z(n54669) );
  IV U69895 ( .A(n49554), .Z(n49555) );
  NOR U69896 ( .A(n49555), .B(n49561), .Z(n54666) );
  IV U69897 ( .A(n49556), .Z(n49563) );
  IV U69898 ( .A(n49557), .Z(n49558) );
  NOR U69899 ( .A(n49563), .B(n49558), .Z(n54674) );
  IV U69900 ( .A(n49559), .Z(n49560) );
  NOR U69901 ( .A(n49561), .B(n49560), .Z(n54672) );
  NOR U69902 ( .A(n54674), .B(n54672), .Z(n53873) );
  NOR U69903 ( .A(n49563), .B(n49562), .Z(n54677) );
  IV U69904 ( .A(n49564), .Z(n49566) );
  NOR U69905 ( .A(n49566), .B(n49565), .Z(n54682) );
  NOR U69906 ( .A(n54677), .B(n54682), .Z(n53872) );
  IV U69907 ( .A(n49567), .Z(n49568) );
  NOR U69908 ( .A(n49568), .B(n49574), .Z(n59087) );
  IV U69909 ( .A(n49569), .Z(n49570) );
  NOR U69910 ( .A(n49571), .B(n49570), .Z(n49572) );
  NOR U69911 ( .A(n59087), .B(n49572), .Z(n54704) );
  IV U69912 ( .A(n49573), .Z(n49575) );
  NOR U69913 ( .A(n49575), .B(n49574), .Z(n59085) );
  IV U69914 ( .A(n49576), .Z(n53835) );
  IV U69915 ( .A(n49577), .Z(n49578) );
  NOR U69916 ( .A(n59074), .B(n49578), .Z(n54722) );
  IV U69917 ( .A(n49579), .Z(n49583) );
  XOR U69918 ( .A(n49595), .B(n53820), .Z(n49581) );
  NOR U69919 ( .A(n49581), .B(n49580), .Z(n49582) );
  IV U69920 ( .A(n49582), .Z(n49586) );
  NOR U69921 ( .A(n49583), .B(n49586), .Z(n49584) );
  IV U69922 ( .A(n49584), .Z(n59071) );
  IV U69923 ( .A(n49585), .Z(n49587) );
  NOR U69924 ( .A(n49587), .B(n49586), .Z(n54730) );
  IV U69925 ( .A(n49588), .Z(n49591) );
  NOR U69926 ( .A(n49589), .B(n53820), .Z(n49590) );
  IV U69927 ( .A(n49590), .Z(n49593) );
  NOR U69928 ( .A(n49591), .B(n49593), .Z(n54727) );
  IV U69929 ( .A(n49592), .Z(n49594) );
  NOR U69930 ( .A(n49594), .B(n49593), .Z(n54736) );
  IV U69931 ( .A(n49595), .Z(n49596) );
  NOR U69932 ( .A(n49596), .B(n53820), .Z(n49597) );
  IV U69933 ( .A(n49597), .Z(n49598) );
  NOR U69934 ( .A(n53819), .B(n49598), .Z(n54733) );
  IV U69935 ( .A(n49599), .Z(n49601) );
  IV U69936 ( .A(n49600), .Z(n59063) );
  NOR U69937 ( .A(n49601), .B(n59063), .Z(n54747) );
  NOR U69938 ( .A(n49603), .B(n49602), .Z(n53803) );
  IV U69939 ( .A(n49604), .Z(n49607) );
  NOR U69940 ( .A(n49605), .B(n53793), .Z(n49606) );
  IV U69941 ( .A(n49606), .Z(n53799) );
  NOR U69942 ( .A(n49607), .B(n53799), .Z(n54753) );
  IV U69943 ( .A(n49608), .Z(n49609) );
  NOR U69944 ( .A(n49610), .B(n49609), .Z(n49611) );
  IV U69945 ( .A(n49611), .Z(n54761) );
  IV U69946 ( .A(n49612), .Z(n49614) );
  NOR U69947 ( .A(n49614), .B(n49613), .Z(n49615) );
  IV U69948 ( .A(n49615), .Z(n53780) );
  IV U69949 ( .A(n49616), .Z(n49618) );
  IV U69950 ( .A(n49617), .Z(n53757) );
  NOR U69951 ( .A(n49618), .B(n53757), .Z(n54765) );
  IV U69952 ( .A(n49619), .Z(n59027) );
  IV U69953 ( .A(n49620), .Z(n49622) );
  NOR U69954 ( .A(n49622), .B(n49621), .Z(n54773) );
  IV U69955 ( .A(n49623), .Z(n49624) );
  NOR U69956 ( .A(n49624), .B(n54778), .Z(n53755) );
  IV U69957 ( .A(n53752), .Z(n65380) );
  NOR U69958 ( .A(n49626), .B(n49625), .Z(n49627) );
  IV U69959 ( .A(n49627), .Z(n49628) );
  NOR U69960 ( .A(n49628), .B(n59009), .Z(n53746) );
  IV U69961 ( .A(n49629), .Z(n49630) );
  NOR U69962 ( .A(n59009), .B(n49630), .Z(n59003) );
  NOR U69963 ( .A(n59009), .B(n49631), .Z(n59000) );
  IV U69964 ( .A(n49632), .Z(n49635) );
  NOR U69965 ( .A(n54791), .B(n49633), .Z(n49634) );
  IV U69966 ( .A(n49634), .Z(n49637) );
  NOR U69967 ( .A(n49635), .B(n49637), .Z(n58996) );
  IV U69968 ( .A(n49636), .Z(n49638) );
  NOR U69969 ( .A(n49638), .B(n49637), .Z(n58993) );
  IV U69970 ( .A(n49639), .Z(n49640) );
  NOR U69971 ( .A(n49640), .B(n54791), .Z(n53745) );
  NOR U69972 ( .A(n49643), .B(n49641), .Z(n58981) );
  IV U69973 ( .A(n49642), .Z(n49644) );
  NOR U69974 ( .A(n49644), .B(n49643), .Z(n58977) );
  IV U69975 ( .A(n49645), .Z(n49649) );
  IV U69976 ( .A(n49646), .Z(n49647) );
  NOR U69977 ( .A(n49649), .B(n49647), .Z(n58984) );
  NOR U69978 ( .A(n49649), .B(n49648), .Z(n60120) );
  IV U69979 ( .A(n49650), .Z(n49651) );
  NOR U69980 ( .A(n49651), .B(n53742), .Z(n64228) );
  NOR U69981 ( .A(n60120), .B(n64228), .Z(n58974) );
  IV U69982 ( .A(n58974), .Z(n53744) );
  NOR U69983 ( .A(n49653), .B(n49652), .Z(n49654) );
  IV U69984 ( .A(n49654), .Z(n49658) );
  NOR U69985 ( .A(n49655), .B(n53731), .Z(n49656) );
  IV U69986 ( .A(n49656), .Z(n49657) );
  NOR U69987 ( .A(n49658), .B(n49657), .Z(n58965) );
  IV U69988 ( .A(n49659), .Z(n49663) );
  NOR U69989 ( .A(n49661), .B(n49660), .Z(n49662) );
  IV U69990 ( .A(n49662), .Z(n49669) );
  NOR U69991 ( .A(n49663), .B(n49669), .Z(n58947) );
  IV U69992 ( .A(n49664), .Z(n49667) );
  NOR U69993 ( .A(n49665), .B(n53701), .Z(n49666) );
  IV U69994 ( .A(n49666), .Z(n53695) );
  NOR U69995 ( .A(n49667), .B(n53695), .Z(n58944) );
  IV U69996 ( .A(n49668), .Z(n49670) );
  NOR U69997 ( .A(n49670), .B(n49669), .Z(n58950) );
  NOR U69998 ( .A(n58944), .B(n58950), .Z(n53712) );
  IV U69999 ( .A(n49671), .Z(n54822) );
  IV U70000 ( .A(n49672), .Z(n49673) );
  NOR U70001 ( .A(n54822), .B(n49673), .Z(n53678) );
  XOR U70002 ( .A(n60164), .B(n54822), .Z(n53681) );
  IV U70003 ( .A(n53681), .Z(n49674) );
  NOR U70004 ( .A(n49674), .B(n54832), .Z(n49675) );
  IV U70005 ( .A(n49675), .Z(n53677) );
  IV U70006 ( .A(n49676), .Z(n49677) );
  NOR U70007 ( .A(n49678), .B(n49677), .Z(n49679) );
  IV U70008 ( .A(n49679), .Z(n54837) );
  IV U70009 ( .A(n49680), .Z(n49682) );
  NOR U70010 ( .A(n49682), .B(n49681), .Z(n54848) );
  NOR U70011 ( .A(n49683), .B(n53666), .Z(n49684) );
  IV U70012 ( .A(n49684), .Z(n49685) );
  NOR U70013 ( .A(n49686), .B(n49685), .Z(n58924) );
  NOR U70014 ( .A(n54848), .B(n58924), .Z(n53668) );
  IV U70015 ( .A(n49687), .Z(n49688) );
  NOR U70016 ( .A(n49688), .B(n54855), .Z(n54851) );
  NOR U70017 ( .A(n49689), .B(n54855), .Z(n53659) );
  IV U70018 ( .A(n49690), .Z(n49691) );
  NOR U70019 ( .A(n49692), .B(n49691), .Z(n70528) );
  IV U70020 ( .A(n49693), .Z(n49694) );
  NOR U70021 ( .A(n49695), .B(n49694), .Z(n70515) );
  NOR U70022 ( .A(n70528), .B(n70515), .Z(n65487) );
  IV U70023 ( .A(n49696), .Z(n49698) );
  IV U70024 ( .A(n49697), .Z(n54863) );
  NOR U70025 ( .A(n49698), .B(n54863), .Z(n58910) );
  IV U70026 ( .A(n49699), .Z(n49700) );
  NOR U70027 ( .A(n49703), .B(n49700), .Z(n54873) );
  IV U70028 ( .A(n49701), .Z(n49702) );
  NOR U70029 ( .A(n49703), .B(n49702), .Z(n54879) );
  IV U70030 ( .A(n49704), .Z(n49707) );
  NOR U70031 ( .A(n49705), .B(n53623), .Z(n49706) );
  IV U70032 ( .A(n49706), .Z(n53638) );
  NOR U70033 ( .A(n49707), .B(n53638), .Z(n58896) );
  IV U70034 ( .A(n49708), .Z(n58888) );
  NOR U70035 ( .A(n49709), .B(n58888), .Z(n53621) );
  IV U70036 ( .A(n49710), .Z(n49711) );
  NOR U70037 ( .A(n49713), .B(n49711), .Z(n54903) );
  IV U70038 ( .A(n49712), .Z(n49714) );
  NOR U70039 ( .A(n49714), .B(n49713), .Z(n54912) );
  IV U70040 ( .A(n49715), .Z(n49716) );
  NOR U70041 ( .A(n49717), .B(n49716), .Z(n54906) );
  NOR U70042 ( .A(n54912), .B(n54906), .Z(n53597) );
  IV U70043 ( .A(n49718), .Z(n49719) );
  NOR U70044 ( .A(n49719), .B(n54916), .Z(n53576) );
  IV U70045 ( .A(n49720), .Z(n49724) );
  IV U70046 ( .A(n49721), .Z(n53570) );
  NOR U70047 ( .A(n49722), .B(n53570), .Z(n49723) );
  IV U70048 ( .A(n49723), .Z(n53574) );
  NOR U70049 ( .A(n49724), .B(n53574), .Z(n58869) );
  IV U70050 ( .A(n49725), .Z(n53562) );
  IV U70051 ( .A(n49726), .Z(n49728) );
  NOR U70052 ( .A(n49728), .B(n49727), .Z(n49729) );
  IV U70053 ( .A(n49729), .Z(n54932) );
  NOR U70054 ( .A(n54935), .B(n49730), .Z(n49735) );
  IV U70055 ( .A(n49731), .Z(n49734) );
  IV U70056 ( .A(n49732), .Z(n49733) );
  NOR U70057 ( .A(n49734), .B(n49733), .Z(n58848) );
  NOR U70058 ( .A(n49735), .B(n58848), .Z(n53549) );
  IV U70059 ( .A(n49736), .Z(n58852) );
  NOR U70060 ( .A(n58852), .B(n54939), .Z(n49737) );
  NOR U70061 ( .A(n49738), .B(n49737), .Z(n53548) );
  IV U70062 ( .A(n49739), .Z(n49740) );
  NOR U70063 ( .A(n49741), .B(n49740), .Z(n58842) );
  IV U70064 ( .A(n49742), .Z(n49743) );
  NOR U70065 ( .A(n49743), .B(n53543), .Z(n54951) );
  IV U70066 ( .A(n49744), .Z(n49745) );
  NOR U70067 ( .A(n49746), .B(n49745), .Z(n54956) );
  IV U70068 ( .A(n49747), .Z(n53524) );
  IV U70069 ( .A(n49748), .Z(n49749) );
  NOR U70070 ( .A(n53524), .B(n49749), .Z(n58834) );
  IV U70071 ( .A(n49750), .Z(n49753) );
  NOR U70072 ( .A(n53524), .B(n49751), .Z(n49752) );
  IV U70073 ( .A(n49752), .Z(n53517) );
  NOR U70074 ( .A(n49753), .B(n53517), .Z(n58827) );
  IV U70075 ( .A(n49754), .Z(n49757) );
  NOR U70076 ( .A(n49755), .B(n53501), .Z(n49756) );
  IV U70077 ( .A(n49756), .Z(n49759) );
  NOR U70078 ( .A(n49757), .B(n49759), .Z(n58824) );
  NOR U70079 ( .A(n58827), .B(n58824), .Z(n53515) );
  IV U70080 ( .A(n49758), .Z(n49760) );
  NOR U70081 ( .A(n49760), .B(n49759), .Z(n53513) );
  IV U70082 ( .A(n53513), .Z(n65602) );
  IV U70083 ( .A(n49761), .Z(n49765) );
  IV U70084 ( .A(n49762), .Z(n53497) );
  NOR U70085 ( .A(n53497), .B(n49763), .Z(n49764) );
  IV U70086 ( .A(n49764), .Z(n49767) );
  NOR U70087 ( .A(n49765), .B(n49767), .Z(n58807) );
  IV U70088 ( .A(n49766), .Z(n49768) );
  NOR U70089 ( .A(n49768), .B(n49767), .Z(n65623) );
  NOR U70090 ( .A(n58807), .B(n65623), .Z(n53489) );
  IV U70091 ( .A(n49769), .Z(n49770) );
  NOR U70092 ( .A(n49770), .B(n49774), .Z(n58796) );
  IV U70093 ( .A(n49771), .Z(n49772) );
  NOR U70094 ( .A(n49772), .B(n49774), .Z(n54973) );
  IV U70095 ( .A(n49773), .Z(n49775) );
  NOR U70096 ( .A(n49775), .B(n49774), .Z(n58799) );
  IV U70097 ( .A(n49776), .Z(n49778) );
  NOR U70098 ( .A(n49778), .B(n49777), .Z(n54978) );
  IV U70099 ( .A(n49779), .Z(n49785) );
  IV U70100 ( .A(n49780), .Z(n49781) );
  NOR U70101 ( .A(n49785), .B(n49781), .Z(n58790) );
  NOR U70102 ( .A(n54978), .B(n58790), .Z(n53488) );
  IV U70103 ( .A(n49782), .Z(n49783) );
  NOR U70104 ( .A(n49783), .B(n69264), .Z(n58783) );
  IV U70105 ( .A(n49784), .Z(n69261) );
  NOR U70106 ( .A(n49785), .B(n69261), .Z(n58793) );
  NOR U70107 ( .A(n58783), .B(n58793), .Z(n53487) );
  IV U70108 ( .A(n49786), .Z(n49787) );
  NOR U70109 ( .A(n49787), .B(n69264), .Z(n58776) );
  IV U70110 ( .A(n49788), .Z(n49789) );
  NOR U70111 ( .A(n49789), .B(n49795), .Z(n49790) );
  IV U70112 ( .A(n49790), .Z(n58782) );
  IV U70113 ( .A(n49791), .Z(n49792) );
  NOR U70114 ( .A(n49793), .B(n49792), .Z(n64000) );
  IV U70115 ( .A(n49794), .Z(n49796) );
  NOR U70116 ( .A(n49796), .B(n49795), .Z(n64005) );
  NOR U70117 ( .A(n64000), .B(n64005), .Z(n58773) );
  IV U70118 ( .A(n49797), .Z(n49799) );
  NOR U70119 ( .A(n49799), .B(n49798), .Z(n58757) );
  IV U70120 ( .A(n49800), .Z(n49801) );
  NOR U70121 ( .A(n49801), .B(n53486), .Z(n58760) );
  IV U70122 ( .A(n49802), .Z(n49806) );
  NOR U70123 ( .A(n49804), .B(n49803), .Z(n49805) );
  IV U70124 ( .A(n49805), .Z(n49809) );
  NOR U70125 ( .A(n49806), .B(n49809), .Z(n58762) );
  XOR U70126 ( .A(n58760), .B(n58762), .Z(n49807) );
  NOR U70127 ( .A(n58757), .B(n49807), .Z(n53482) );
  IV U70128 ( .A(n49808), .Z(n49810) );
  NOR U70129 ( .A(n49810), .B(n49809), .Z(n58765) );
  IV U70130 ( .A(n49811), .Z(n49815) );
  IV U70131 ( .A(n49812), .Z(n49813) );
  NOR U70132 ( .A(n49813), .B(n53480), .Z(n49814) );
  IV U70133 ( .A(n49814), .Z(n49817) );
  NOR U70134 ( .A(n49815), .B(n49817), .Z(n58753) );
  IV U70135 ( .A(n49816), .Z(n49818) );
  NOR U70136 ( .A(n49818), .B(n49817), .Z(n58750) );
  IV U70137 ( .A(n49819), .Z(n53472) );
  NOR U70138 ( .A(n53472), .B(n49820), .Z(n49822) );
  NOR U70139 ( .A(n49822), .B(n49821), .Z(n49823) );
  IV U70140 ( .A(n49823), .Z(n53467) );
  IV U70141 ( .A(n49824), .Z(n49826) );
  IV U70142 ( .A(n49825), .Z(n53463) );
  NOR U70143 ( .A(n49826), .B(n53463), .Z(n54993) );
  IV U70144 ( .A(n54984), .Z(n49827) );
  XOR U70145 ( .A(n49826), .B(n49825), .Z(n54983) );
  NOR U70146 ( .A(n49827), .B(n54983), .Z(n54991) );
  NOR U70147 ( .A(n54993), .B(n54991), .Z(n53460) );
  IV U70148 ( .A(n49828), .Z(n49829) );
  NOR U70149 ( .A(n49829), .B(n53458), .Z(n54996) );
  IV U70150 ( .A(n49830), .Z(n49831) );
  NOR U70151 ( .A(n53442), .B(n49831), .Z(n53440) );
  NOR U70152 ( .A(n49832), .B(n53422), .Z(n49833) );
  IV U70153 ( .A(n49833), .Z(n58734) );
  NOR U70154 ( .A(n58734), .B(n49834), .Z(n53438) );
  IV U70155 ( .A(n49837), .Z(n49835) );
  NOR U70156 ( .A(n53412), .B(n49835), .Z(n55013) );
  IV U70157 ( .A(n49836), .Z(n49839) );
  XOR U70158 ( .A(n49837), .B(n53412), .Z(n49838) );
  NOR U70159 ( .A(n49839), .B(n49838), .Z(n55008) );
  NOR U70160 ( .A(n55013), .B(n55008), .Z(n53410) );
  IV U70161 ( .A(n49840), .Z(n49841) );
  NOR U70162 ( .A(n49842), .B(n49841), .Z(n55017) );
  IV U70163 ( .A(n49843), .Z(n49850) );
  IV U70164 ( .A(n49844), .Z(n49845) );
  NOR U70165 ( .A(n49850), .B(n49845), .Z(n58717) );
  NOR U70166 ( .A(n55017), .B(n58717), .Z(n53409) );
  IV U70167 ( .A(n49846), .Z(n49847) );
  NOR U70168 ( .A(n49847), .B(n49852), .Z(n58714) );
  IV U70169 ( .A(n49848), .Z(n49849) );
  NOR U70170 ( .A(n49850), .B(n49849), .Z(n58720) );
  NOR U70171 ( .A(n58714), .B(n58720), .Z(n53408) );
  IV U70172 ( .A(n49851), .Z(n49853) );
  NOR U70173 ( .A(n49853), .B(n49852), .Z(n55019) );
  IV U70174 ( .A(n49854), .Z(n49855) );
  NOR U70175 ( .A(n49858), .B(n49855), .Z(n58697) );
  IV U70176 ( .A(n49856), .Z(n49857) );
  NOR U70177 ( .A(n49858), .B(n49857), .Z(n55021) );
  NOR U70178 ( .A(n49859), .B(n49861), .Z(n58700) );
  IV U70179 ( .A(n49860), .Z(n49862) );
  NOR U70180 ( .A(n49862), .B(n49861), .Z(n55025) );
  IV U70181 ( .A(n49863), .Z(n49864) );
  NOR U70182 ( .A(n49864), .B(n49866), .Z(n60375) );
  IV U70183 ( .A(n49865), .Z(n49869) );
  NOR U70184 ( .A(n49867), .B(n49866), .Z(n49868) );
  IV U70185 ( .A(n49868), .Z(n49871) );
  NOR U70186 ( .A(n49869), .B(n49871), .Z(n60369) );
  IV U70187 ( .A(n49870), .Z(n49872) );
  NOR U70188 ( .A(n49872), .B(n49871), .Z(n60373) );
  NOR U70189 ( .A(n60369), .B(n60373), .Z(n49873) );
  IV U70190 ( .A(n49873), .Z(n49874) );
  NOR U70191 ( .A(n60375), .B(n49874), .Z(n58691) );
  IV U70192 ( .A(n58691), .Z(n53407) );
  IV U70193 ( .A(n49875), .Z(n49879) );
  NOR U70194 ( .A(n49877), .B(n49876), .Z(n49878) );
  IV U70195 ( .A(n49878), .Z(n53397) );
  NOR U70196 ( .A(n49879), .B(n53397), .Z(n58682) );
  IV U70197 ( .A(n49880), .Z(n49881) );
  NOR U70198 ( .A(n55039), .B(n49881), .Z(n55045) );
  IV U70199 ( .A(n49882), .Z(n49883) );
  NOR U70200 ( .A(n49884), .B(n49883), .Z(n55048) );
  IV U70201 ( .A(n49885), .Z(n49888) );
  IV U70202 ( .A(n49886), .Z(n49887) );
  NOR U70203 ( .A(n49888), .B(n49887), .Z(n58671) );
  NOR U70204 ( .A(n55048), .B(n58671), .Z(n53387) );
  IV U70205 ( .A(n49889), .Z(n49890) );
  NOR U70206 ( .A(n49890), .B(n49892), .Z(n58664) );
  IV U70207 ( .A(n49891), .Z(n49893) );
  NOR U70208 ( .A(n49893), .B(n49892), .Z(n58668) );
  IV U70209 ( .A(n49894), .Z(n49895) );
  NOR U70210 ( .A(n49896), .B(n49895), .Z(n58656) );
  IV U70211 ( .A(n49897), .Z(n49898) );
  NOR U70212 ( .A(n49899), .B(n49898), .Z(n49900) );
  IV U70213 ( .A(n49900), .Z(n55051) );
  IV U70214 ( .A(n49901), .Z(n53383) );
  IV U70215 ( .A(n49902), .Z(n49903) );
  NOR U70216 ( .A(n53383), .B(n49903), .Z(n58653) );
  IV U70217 ( .A(n49904), .Z(n49908) );
  NOR U70218 ( .A(n49906), .B(n49905), .Z(n49907) );
  IV U70219 ( .A(n49907), .Z(n49910) );
  NOR U70220 ( .A(n49908), .B(n49910), .Z(n58650) );
  NOR U70221 ( .A(n58653), .B(n58650), .Z(n53386) );
  IV U70222 ( .A(n49909), .Z(n49911) );
  NOR U70223 ( .A(n49911), .B(n49910), .Z(n58647) );
  IV U70224 ( .A(n49912), .Z(n49914) );
  IV U70225 ( .A(n49913), .Z(n49918) );
  NOR U70226 ( .A(n49914), .B(n49918), .Z(n58643) );
  NOR U70227 ( .A(n58647), .B(n58643), .Z(n53380) );
  IV U70228 ( .A(n49915), .Z(n49916) );
  NOR U70229 ( .A(n49916), .B(n49918), .Z(n58641) );
  IV U70230 ( .A(n49917), .Z(n49919) );
  NOR U70231 ( .A(n49919), .B(n49918), .Z(n55058) );
  IV U70232 ( .A(n49920), .Z(n49921) );
  NOR U70233 ( .A(n49922), .B(n49921), .Z(n49923) );
  IV U70234 ( .A(n49923), .Z(n53371) );
  IV U70235 ( .A(n49924), .Z(n49927) );
  IV U70236 ( .A(n49925), .Z(n49926) );
  NOR U70237 ( .A(n49927), .B(n49926), .Z(n58632) );
  IV U70238 ( .A(n49928), .Z(n49931) );
  NOR U70239 ( .A(n49929), .B(n49934), .Z(n49930) );
  IV U70240 ( .A(n49930), .Z(n53366) );
  NOR U70241 ( .A(n49931), .B(n53366), .Z(n53358) );
  IV U70242 ( .A(n49932), .Z(n49933) );
  NOR U70243 ( .A(n49934), .B(n49933), .Z(n53355) );
  IV U70244 ( .A(n53355), .Z(n53349) );
  NOR U70245 ( .A(n58617), .B(n55072), .Z(n53347) );
  IV U70246 ( .A(n49935), .Z(n49936) );
  NOR U70247 ( .A(n55083), .B(n49936), .Z(n55077) );
  IV U70248 ( .A(n49937), .Z(n49938) );
  NOR U70249 ( .A(n55083), .B(n49938), .Z(n58620) );
  IV U70250 ( .A(n49939), .Z(n49940) );
  NOR U70251 ( .A(n55083), .B(n49940), .Z(n53346) );
  IV U70252 ( .A(n49941), .Z(n49945) );
  NOR U70253 ( .A(n49943), .B(n49942), .Z(n49944) );
  IV U70254 ( .A(n49944), .Z(n49947) );
  NOR U70255 ( .A(n49945), .B(n49947), .Z(n58602) );
  IV U70256 ( .A(n49946), .Z(n49948) );
  NOR U70257 ( .A(n49948), .B(n49947), .Z(n55089) );
  IV U70258 ( .A(n49949), .Z(n49950) );
  NOR U70259 ( .A(n53339), .B(n49950), .Z(n55099) );
  IV U70260 ( .A(n49951), .Z(n49955) );
  NOR U70261 ( .A(n49953), .B(n49952), .Z(n49954) );
  IV U70262 ( .A(n49954), .Z(n49957) );
  NOR U70263 ( .A(n49955), .B(n49957), .Z(n55104) );
  NOR U70264 ( .A(n55099), .B(n55104), .Z(n53333) );
  IV U70265 ( .A(n49956), .Z(n49958) );
  NOR U70266 ( .A(n49958), .B(n49957), .Z(n55101) );
  IV U70267 ( .A(n49959), .Z(n55115) );
  IV U70268 ( .A(n49960), .Z(n49962) );
  NOR U70269 ( .A(n49962), .B(n49961), .Z(n60443) );
  NOR U70270 ( .A(n60447), .B(n60443), .Z(n58589) );
  NOR U70271 ( .A(n49964), .B(n49963), .Z(n49965) );
  IV U70272 ( .A(n49965), .Z(n49966) );
  NOR U70273 ( .A(n49967), .B(n49966), .Z(n55117) );
  IV U70274 ( .A(n49968), .Z(n49971) );
  NOR U70275 ( .A(n49969), .B(n49974), .Z(n49970) );
  IV U70276 ( .A(n49970), .Z(n53320) );
  NOR U70277 ( .A(n49971), .B(n53320), .Z(n58569) );
  IV U70278 ( .A(n49972), .Z(n49973) );
  NOR U70279 ( .A(n49974), .B(n49973), .Z(n58560) );
  IV U70280 ( .A(n49975), .Z(n49976) );
  NOR U70281 ( .A(n49977), .B(n49976), .Z(n58557) );
  NOR U70282 ( .A(n58560), .B(n58557), .Z(n53318) );
  IV U70283 ( .A(n49978), .Z(n49981) );
  NOR U70284 ( .A(n49979), .B(n49989), .Z(n49980) );
  IV U70285 ( .A(n49980), .Z(n49984) );
  NOR U70286 ( .A(n49981), .B(n49984), .Z(n49982) );
  IV U70287 ( .A(n49982), .Z(n58556) );
  IV U70288 ( .A(n49983), .Z(n49985) );
  NOR U70289 ( .A(n49985), .B(n49984), .Z(n49986) );
  IV U70290 ( .A(n49986), .Z(n55121) );
  IV U70291 ( .A(n49990), .Z(n49987) );
  NOR U70292 ( .A(n49987), .B(n49989), .Z(n58552) );
  IV U70293 ( .A(n49988), .Z(n49992) );
  XOR U70294 ( .A(n49990), .B(n49989), .Z(n49991) );
  NOR U70295 ( .A(n49992), .B(n49991), .Z(n55122) );
  NOR U70296 ( .A(n58552), .B(n55122), .Z(n53316) );
  IV U70297 ( .A(n49993), .Z(n49994) );
  NOR U70298 ( .A(n49995), .B(n49994), .Z(n58550) );
  IV U70299 ( .A(n49996), .Z(n49997) );
  NOR U70300 ( .A(n49998), .B(n49997), .Z(n55130) );
  IV U70301 ( .A(n49999), .Z(n50003) );
  NOR U70302 ( .A(n50003), .B(n50000), .Z(n55139) );
  IV U70303 ( .A(n50001), .Z(n50002) );
  NOR U70304 ( .A(n50003), .B(n50002), .Z(n55134) );
  NOR U70305 ( .A(n55139), .B(n55134), .Z(n53306) );
  IV U70306 ( .A(n50004), .Z(n50007) );
  NOR U70307 ( .A(n50005), .B(n53300), .Z(n50006) );
  IV U70308 ( .A(n50006), .Z(n53304) );
  NOR U70309 ( .A(n50007), .B(n53304), .Z(n55136) );
  IV U70310 ( .A(n50008), .Z(n50009) );
  NOR U70311 ( .A(n50009), .B(n53298), .Z(n50010) );
  IV U70312 ( .A(n50010), .Z(n55151) );
  IV U70313 ( .A(n50011), .Z(n55156) );
  NOR U70314 ( .A(n55156), .B(n50012), .Z(n55165) );
  NOR U70315 ( .A(n55170), .B(n55165), .Z(n53291) );
  IV U70316 ( .A(n50013), .Z(n50014) );
  NOR U70317 ( .A(n50015), .B(n50014), .Z(n58526) );
  IV U70318 ( .A(n50015), .Z(n50018) );
  NOR U70319 ( .A(n55188), .B(n55177), .Z(n50016) );
  IV U70320 ( .A(n50016), .Z(n50017) );
  NOR U70321 ( .A(n50018), .B(n50017), .Z(n55181) );
  IV U70322 ( .A(n50019), .Z(n50020) );
  NOR U70323 ( .A(n50021), .B(n50020), .Z(n55189) );
  NOR U70324 ( .A(n55189), .B(n50022), .Z(n55185) );
  IV U70325 ( .A(n50023), .Z(n50024) );
  NOR U70326 ( .A(n50025), .B(n50024), .Z(n53288) );
  IV U70327 ( .A(n53288), .Z(n53278) );
  IV U70328 ( .A(n50026), .Z(n50027) );
  NOR U70329 ( .A(n50028), .B(n50027), .Z(n53275) );
  IV U70330 ( .A(n53275), .Z(n53273) );
  IV U70331 ( .A(n50029), .Z(n50031) );
  NOR U70332 ( .A(n50031), .B(n50030), .Z(n58505) );
  IV U70333 ( .A(n50032), .Z(n50033) );
  NOR U70334 ( .A(n50033), .B(n55205), .Z(n53271) );
  IV U70335 ( .A(n50034), .Z(n50035) );
  NOR U70336 ( .A(n50036), .B(n50035), .Z(n50037) );
  NOR U70337 ( .A(n58474), .B(n50037), .Z(n50038) );
  IV U70338 ( .A(n50038), .Z(n53260) );
  NOR U70339 ( .A(n50040), .B(n50039), .Z(n58471) );
  IV U70340 ( .A(n50041), .Z(n50042) );
  NOR U70341 ( .A(n50045), .B(n50042), .Z(n55231) );
  IV U70342 ( .A(n50043), .Z(n50044) );
  NOR U70343 ( .A(n50045), .B(n50044), .Z(n58441) );
  IV U70344 ( .A(n50046), .Z(n50049) );
  IV U70345 ( .A(n50047), .Z(n50048) );
  NOR U70346 ( .A(n50049), .B(n50048), .Z(n55234) );
  IV U70347 ( .A(n50050), .Z(n50053) );
  IV U70348 ( .A(n50051), .Z(n50052) );
  NOR U70349 ( .A(n50053), .B(n50052), .Z(n55237) );
  NOR U70350 ( .A(n55244), .B(n55237), .Z(n53241) );
  NOR U70351 ( .A(n50054), .B(n55241), .Z(n53240) );
  IV U70352 ( .A(n50055), .Z(n50056) );
  NOR U70353 ( .A(n50056), .B(n55241), .Z(n50057) );
  IV U70354 ( .A(n50057), .Z(n50058) );
  NOR U70355 ( .A(n53234), .B(n50058), .Z(n58432) );
  NOR U70356 ( .A(n50059), .B(n55252), .Z(n53226) );
  IV U70357 ( .A(n50060), .Z(n50061) );
  NOR U70358 ( .A(n50062), .B(n50061), .Z(n60562) );
  IV U70359 ( .A(n50063), .Z(n50064) );
  NOR U70360 ( .A(n50067), .B(n50064), .Z(n63727) );
  NOR U70361 ( .A(n60562), .B(n63727), .Z(n58418) );
  IV U70362 ( .A(n58418), .Z(n53225) );
  IV U70363 ( .A(n50065), .Z(n50066) );
  NOR U70364 ( .A(n50067), .B(n50066), .Z(n58415) );
  IV U70365 ( .A(n50068), .Z(n50070) );
  NOR U70366 ( .A(n50070), .B(n50069), .Z(n58412) );
  IV U70367 ( .A(n50071), .Z(n50072) );
  NOR U70368 ( .A(n50072), .B(n50074), .Z(n58410) );
  NOR U70369 ( .A(n58412), .B(n58410), .Z(n53224) );
  IV U70370 ( .A(n50073), .Z(n50075) );
  NOR U70371 ( .A(n50075), .B(n50074), .Z(n55258) );
  IV U70372 ( .A(n50076), .Z(n50078) );
  XOR U70373 ( .A(n50084), .B(n58396), .Z(n50077) );
  NOR U70374 ( .A(n50078), .B(n50077), .Z(n58406) );
  NOR U70375 ( .A(n55258), .B(n58406), .Z(n53223) );
  IV U70376 ( .A(n50079), .Z(n50080) );
  NOR U70377 ( .A(n50080), .B(n58396), .Z(n55260) );
  IV U70378 ( .A(n50081), .Z(n50083) );
  NOR U70379 ( .A(n50083), .B(n50082), .Z(n58384) );
  IV U70380 ( .A(n50084), .Z(n50085) );
  NOR U70381 ( .A(n50085), .B(n58396), .Z(n58379) );
  NOR U70382 ( .A(n58384), .B(n58379), .Z(n53222) );
  IV U70383 ( .A(n50093), .Z(n50086) );
  NOR U70384 ( .A(n50086), .B(n50091), .Z(n55271) );
  IV U70385 ( .A(n50087), .Z(n50088) );
  NOR U70386 ( .A(n53217), .B(n50088), .Z(n55264) );
  NOR U70387 ( .A(n55268), .B(n55264), .Z(n50089) );
  IV U70388 ( .A(n50089), .Z(n50090) );
  NOR U70389 ( .A(n55271), .B(n50090), .Z(n50095) );
  IV U70390 ( .A(n50091), .Z(n50092) );
  NOR U70391 ( .A(n50093), .B(n50092), .Z(n50094) );
  NOR U70392 ( .A(n50095), .B(n50094), .Z(n53212) );
  IV U70393 ( .A(n50096), .Z(n50097) );
  NOR U70394 ( .A(n50098), .B(n50097), .Z(n53161) );
  IV U70395 ( .A(n53161), .Z(n53154) );
  IV U70396 ( .A(n50099), .Z(n50100) );
  NOR U70397 ( .A(n50103), .B(n50100), .Z(n55292) );
  IV U70398 ( .A(n50101), .Z(n50102) );
  NOR U70399 ( .A(n50103), .B(n50102), .Z(n58350) );
  IV U70400 ( .A(n50104), .Z(n50107) );
  NOR U70401 ( .A(n50105), .B(n55312), .Z(n50106) );
  IV U70402 ( .A(n50106), .Z(n50109) );
  NOR U70403 ( .A(n50107), .B(n50109), .Z(n55301) );
  IV U70404 ( .A(n50108), .Z(n50110) );
  NOR U70405 ( .A(n50110), .B(n50109), .Z(n55307) );
  IV U70406 ( .A(n50111), .Z(n53131) );
  NOR U70407 ( .A(n50112), .B(n53131), .Z(n53123) );
  IV U70408 ( .A(n50113), .Z(n50114) );
  NOR U70409 ( .A(n50114), .B(n50122), .Z(n50115) );
  IV U70410 ( .A(n50115), .Z(n55325) );
  IV U70411 ( .A(n50116), .Z(n50117) );
  NOR U70412 ( .A(n50117), .B(n50122), .Z(n55330) );
  IV U70413 ( .A(n50118), .Z(n50120) );
  NOR U70414 ( .A(n50120), .B(n50119), .Z(n58321) );
  IV U70415 ( .A(n50121), .Z(n50123) );
  NOR U70416 ( .A(n50123), .B(n50122), .Z(n55333) );
  NOR U70417 ( .A(n58321), .B(n55333), .Z(n53110) );
  IV U70418 ( .A(n50124), .Z(n50125) );
  NOR U70419 ( .A(n50126), .B(n50125), .Z(n53106) );
  IV U70420 ( .A(n50127), .Z(n53102) );
  IV U70421 ( .A(n50128), .Z(n53101) );
  IV U70422 ( .A(n50129), .Z(n50130) );
  NOR U70423 ( .A(n50132), .B(n50130), .Z(n55342) );
  IV U70424 ( .A(n50131), .Z(n50133) );
  NOR U70425 ( .A(n50133), .B(n50132), .Z(n55351) );
  IV U70426 ( .A(n50134), .Z(n50135) );
  NOR U70427 ( .A(n50135), .B(n50138), .Z(n50136) );
  IV U70428 ( .A(n50136), .Z(n55356) );
  IV U70429 ( .A(n50137), .Z(n50139) );
  NOR U70430 ( .A(n50139), .B(n50138), .Z(n53085) );
  IV U70431 ( .A(n53085), .Z(n53079) );
  IV U70432 ( .A(n50140), .Z(n50141) );
  NOR U70433 ( .A(n50142), .B(n50141), .Z(n55357) );
  XOR U70434 ( .A(n50148), .B(n50150), .Z(n50145) );
  IV U70435 ( .A(n50143), .Z(n50144) );
  NOR U70436 ( .A(n50145), .B(n50144), .Z(n55364) );
  IV U70437 ( .A(n50146), .Z(n50147) );
  NOR U70438 ( .A(n50150), .B(n50147), .Z(n55371) );
  IV U70439 ( .A(n50148), .Z(n50149) );
  NOR U70440 ( .A(n50150), .B(n50149), .Z(n55374) );
  NOR U70441 ( .A(n55371), .B(n55374), .Z(n53066) );
  IV U70442 ( .A(n50151), .Z(n50152) );
  NOR U70443 ( .A(n50153), .B(n50152), .Z(n50154) );
  IV U70444 ( .A(n50154), .Z(n53061) );
  IV U70445 ( .A(n50155), .Z(n53059) );
  NOR U70446 ( .A(n50156), .B(n53059), .Z(n50157) );
  IV U70447 ( .A(n50157), .Z(n58298) );
  NOR U70448 ( .A(n58298), .B(n50158), .Z(n53054) );
  IV U70449 ( .A(n50159), .Z(n50163) );
  NOR U70450 ( .A(n50161), .B(n50160), .Z(n50162) );
  IV U70451 ( .A(n50162), .Z(n50169) );
  NOR U70452 ( .A(n50163), .B(n50169), .Z(n55385) );
  IV U70453 ( .A(n50164), .Z(n50167) );
  NOR U70454 ( .A(n50165), .B(n50172), .Z(n50166) );
  IV U70455 ( .A(n50166), .Z(n50175) );
  NOR U70456 ( .A(n50167), .B(n50175), .Z(n55398) );
  IV U70457 ( .A(n50168), .Z(n50170) );
  NOR U70458 ( .A(n50170), .B(n50169), .Z(n55393) );
  NOR U70459 ( .A(n55398), .B(n55393), .Z(n53031) );
  IV U70460 ( .A(n50171), .Z(n50173) );
  NOR U70461 ( .A(n50173), .B(n50172), .Z(n55401) );
  IV U70462 ( .A(n50174), .Z(n50176) );
  NOR U70463 ( .A(n50176), .B(n50175), .Z(n55396) );
  NOR U70464 ( .A(n55401), .B(n55396), .Z(n53030) );
  IV U70465 ( .A(n50177), .Z(n50178) );
  NOR U70466 ( .A(n50179), .B(n50178), .Z(n58276) );
  IV U70467 ( .A(n50180), .Z(n50181) );
  NOR U70468 ( .A(n50182), .B(n50181), .Z(n55404) );
  NOR U70469 ( .A(n58276), .B(n55404), .Z(n53029) );
  IV U70470 ( .A(n50183), .Z(n58271) );
  IV U70471 ( .A(n50184), .Z(n50185) );
  NOR U70472 ( .A(n50185), .B(n55414), .Z(n53023) );
  IV U70473 ( .A(n50186), .Z(n50189) );
  NOR U70474 ( .A(n50187), .B(n50192), .Z(n50188) );
  IV U70475 ( .A(n50188), .Z(n50194) );
  NOR U70476 ( .A(n50189), .B(n50194), .Z(n55420) );
  IV U70477 ( .A(n50190), .Z(n50191) );
  NOR U70478 ( .A(n50192), .B(n50191), .Z(n58256) );
  IV U70479 ( .A(n50193), .Z(n50195) );
  NOR U70480 ( .A(n50195), .B(n50194), .Z(n58258) );
  NOR U70481 ( .A(n58256), .B(n58258), .Z(n50196) );
  IV U70482 ( .A(n50196), .Z(n53022) );
  IV U70483 ( .A(n50197), .Z(n50202) );
  IV U70484 ( .A(n50198), .Z(n50199) );
  NOR U70485 ( .A(n50202), .B(n50199), .Z(n58253) );
  IV U70486 ( .A(n50200), .Z(n50201) );
  NOR U70487 ( .A(n50202), .B(n50201), .Z(n58243) );
  IV U70488 ( .A(n50203), .Z(n50204) );
  NOR U70489 ( .A(n50205), .B(n50204), .Z(n55424) );
  IV U70490 ( .A(n50206), .Z(n50208) );
  NOR U70491 ( .A(n50208), .B(n50207), .Z(n60702) );
  NOR U70492 ( .A(n63517), .B(n60702), .Z(n58247) );
  IV U70493 ( .A(n50209), .Z(n50210) );
  NOR U70494 ( .A(n55430), .B(n50210), .Z(n58236) );
  IV U70495 ( .A(n50211), .Z(n50212) );
  NOR U70496 ( .A(n55430), .B(n50212), .Z(n50213) );
  NOR U70497 ( .A(n58236), .B(n50213), .Z(n53021) );
  IV U70498 ( .A(n50214), .Z(n50215) );
  NOR U70499 ( .A(n50217), .B(n50215), .Z(n55439) );
  IV U70500 ( .A(n50216), .Z(n50218) );
  NOR U70501 ( .A(n50218), .B(n50217), .Z(n55436) );
  NOR U70502 ( .A(n50219), .B(n50223), .Z(n50220) );
  IV U70503 ( .A(n50220), .Z(n55443) );
  NOR U70504 ( .A(n55443), .B(n50221), .Z(n53020) );
  IV U70505 ( .A(n50222), .Z(n50224) );
  NOR U70506 ( .A(n50224), .B(n50223), .Z(n53017) );
  IV U70507 ( .A(n53017), .Z(n53008) );
  IV U70508 ( .A(n50225), .Z(n50226) );
  NOR U70509 ( .A(n50226), .B(n50234), .Z(n58226) );
  IV U70510 ( .A(n50227), .Z(n50228) );
  NOR U70511 ( .A(n50229), .B(n50228), .Z(n58228) );
  NOR U70512 ( .A(n58226), .B(n58228), .Z(n53010) );
  IV U70513 ( .A(n50230), .Z(n50231) );
  NOR U70514 ( .A(n50232), .B(n50231), .Z(n55452) );
  IV U70515 ( .A(n50233), .Z(n50235) );
  NOR U70516 ( .A(n50235), .B(n50234), .Z(n58223) );
  NOR U70517 ( .A(n55452), .B(n58223), .Z(n53007) );
  IV U70518 ( .A(n50236), .Z(n50238) );
  NOR U70519 ( .A(n50238), .B(n50237), .Z(n55450) );
  NOR U70520 ( .A(n58219), .B(n55456), .Z(n50239) );
  NOR U70521 ( .A(n55457), .B(n50239), .Z(n53006) );
  IV U70522 ( .A(n50240), .Z(n50242) );
  NOR U70523 ( .A(n50242), .B(n50241), .Z(n58208) );
  NOR U70524 ( .A(n58206), .B(n58208), .Z(n50243) );
  IV U70525 ( .A(n50243), .Z(n53004) );
  IV U70526 ( .A(n50244), .Z(n50245) );
  NOR U70527 ( .A(n50246), .B(n50245), .Z(n58188) );
  IV U70528 ( .A(n50247), .Z(n50248) );
  NOR U70529 ( .A(n50249), .B(n50248), .Z(n58203) );
  NOR U70530 ( .A(n58188), .B(n58203), .Z(n53003) );
  IV U70531 ( .A(n50250), .Z(n50251) );
  NOR U70532 ( .A(n50252), .B(n50251), .Z(n58194) );
  NOR U70533 ( .A(n58192), .B(n58194), .Z(n53002) );
  NOR U70534 ( .A(n50254), .B(n50253), .Z(n53001) );
  IV U70535 ( .A(n50255), .Z(n50258) );
  IV U70536 ( .A(n50256), .Z(n50257) );
  NOR U70537 ( .A(n50258), .B(n50257), .Z(n58176) );
  NOR U70538 ( .A(n58169), .B(n58176), .Z(n52999) );
  IV U70539 ( .A(n50259), .Z(n50263) );
  NOR U70540 ( .A(n50261), .B(n50260), .Z(n50262) );
  IV U70541 ( .A(n50262), .Z(n50265) );
  NOR U70542 ( .A(n50263), .B(n50265), .Z(n55464) );
  IV U70543 ( .A(n50264), .Z(n50266) );
  NOR U70544 ( .A(n50266), .B(n50265), .Z(n50267) );
  IV U70545 ( .A(n50267), .Z(n58168) );
  IV U70546 ( .A(n50268), .Z(n50269) );
  NOR U70547 ( .A(n50269), .B(n52987), .Z(n52983) );
  IV U70548 ( .A(n50270), .Z(n50271) );
  NOR U70549 ( .A(n52987), .B(n50271), .Z(n50272) );
  IV U70550 ( .A(n50272), .Z(n58164) );
  IV U70551 ( .A(n50273), .Z(n50278) );
  IV U70552 ( .A(n50274), .Z(n50275) );
  NOR U70553 ( .A(n50278), .B(n50275), .Z(n58159) );
  IV U70554 ( .A(n50276), .Z(n50277) );
  NOR U70555 ( .A(n50278), .B(n50277), .Z(n55468) );
  IV U70556 ( .A(n50279), .Z(n50282) );
  NOR U70557 ( .A(n50280), .B(n50288), .Z(n50281) );
  IV U70558 ( .A(n50281), .Z(n50284) );
  NOR U70559 ( .A(n50282), .B(n50284), .Z(n58153) );
  IV U70560 ( .A(n50283), .Z(n50285) );
  NOR U70561 ( .A(n50285), .B(n50284), .Z(n55471) );
  IV U70562 ( .A(n50286), .Z(n50287) );
  NOR U70563 ( .A(n50288), .B(n50287), .Z(n58148) );
  IV U70564 ( .A(n50289), .Z(n50290) );
  NOR U70565 ( .A(n50290), .B(n50292), .Z(n63443) );
  IV U70566 ( .A(n50291), .Z(n50293) );
  NOR U70567 ( .A(n50293), .B(n50292), .Z(n63447) );
  NOR U70568 ( .A(n63443), .B(n63447), .Z(n55475) );
  IV U70569 ( .A(n50294), .Z(n50297) );
  NOR U70570 ( .A(n50295), .B(n52969), .Z(n50296) );
  IV U70571 ( .A(n50296), .Z(n52975) );
  NOR U70572 ( .A(n50297), .B(n52975), .Z(n55479) );
  IV U70573 ( .A(n50298), .Z(n50299) );
  NOR U70574 ( .A(n50311), .B(n50299), .Z(n55490) );
  IV U70575 ( .A(n50300), .Z(n50302) );
  NOR U70576 ( .A(n50302), .B(n50301), .Z(n55485) );
  NOR U70577 ( .A(n55490), .B(n55485), .Z(n52966) );
  XOR U70578 ( .A(n50309), .B(n50311), .Z(n50305) );
  IV U70579 ( .A(n50303), .Z(n50304) );
  NOR U70580 ( .A(n50305), .B(n50304), .Z(n55496) );
  IV U70581 ( .A(n50306), .Z(n50307) );
  NOR U70582 ( .A(n50308), .B(n50307), .Z(n55499) );
  IV U70583 ( .A(n50309), .Z(n50310) );
  NOR U70584 ( .A(n50311), .B(n50310), .Z(n55494) );
  NOR U70585 ( .A(n55499), .B(n55494), .Z(n52965) );
  IV U70586 ( .A(n50312), .Z(n50314) );
  NOR U70587 ( .A(n50314), .B(n50313), .Z(n55507) );
  IV U70588 ( .A(n50315), .Z(n50317) );
  NOR U70589 ( .A(n50317), .B(n50316), .Z(n55504) );
  IV U70590 ( .A(n50318), .Z(n50320) );
  NOR U70591 ( .A(n50320), .B(n50319), .Z(n55502) );
  NOR U70592 ( .A(n55504), .B(n55502), .Z(n50321) );
  IV U70593 ( .A(n50321), .Z(n50322) );
  NOR U70594 ( .A(n55507), .B(n50322), .Z(n52964) );
  IV U70595 ( .A(n50323), .Z(n50325) );
  IV U70596 ( .A(n50324), .Z(n50327) );
  NOR U70597 ( .A(n50325), .B(n50327), .Z(n55510) );
  IV U70598 ( .A(n50326), .Z(n50328) );
  NOR U70599 ( .A(n50328), .B(n50327), .Z(n58129) );
  NOR U70600 ( .A(n58131), .B(n58129), .Z(n52963) );
  IV U70601 ( .A(n50329), .Z(n50330) );
  NOR U70602 ( .A(n50330), .B(n50338), .Z(n58121) );
  NOR U70603 ( .A(n50332), .B(n50331), .Z(n58124) );
  NOR U70604 ( .A(n58121), .B(n58124), .Z(n52962) );
  IV U70605 ( .A(n50333), .Z(n50334) );
  NOR U70606 ( .A(n50334), .B(n50338), .Z(n50335) );
  IV U70607 ( .A(n50335), .Z(n50336) );
  NOR U70608 ( .A(n50337), .B(n50336), .Z(n58118) );
  IV U70609 ( .A(n50337), .Z(n50342) );
  NOR U70610 ( .A(n50339), .B(n50338), .Z(n50340) );
  IV U70611 ( .A(n50340), .Z(n50341) );
  NOR U70612 ( .A(n50342), .B(n50341), .Z(n58114) );
  NOR U70613 ( .A(n50344), .B(n50343), .Z(n50345) );
  IV U70614 ( .A(n50345), .Z(n58112) );
  IV U70615 ( .A(n50346), .Z(n52953) );
  NOR U70616 ( .A(n52953), .B(n50347), .Z(n58108) );
  IV U70617 ( .A(n50348), .Z(n50350) );
  NOR U70618 ( .A(n50350), .B(n50349), .Z(n55522) );
  NOR U70619 ( .A(n58108), .B(n55522), .Z(n52950) );
  IV U70620 ( .A(n50351), .Z(n50355) );
  NOR U70621 ( .A(n50353), .B(n50352), .Z(n50354) );
  IV U70622 ( .A(n50354), .Z(n50357) );
  NOR U70623 ( .A(n50355), .B(n50357), .Z(n58105) );
  IV U70624 ( .A(n50356), .Z(n50358) );
  NOR U70625 ( .A(n50358), .B(n50357), .Z(n55527) );
  IV U70626 ( .A(n50359), .Z(n50363) );
  IV U70627 ( .A(n50360), .Z(n50372) );
  NOR U70628 ( .A(n50372), .B(n50361), .Z(n50362) );
  IV U70629 ( .A(n50362), .Z(n50365) );
  NOR U70630 ( .A(n50363), .B(n50365), .Z(n55524) );
  IV U70631 ( .A(n50364), .Z(n50366) );
  NOR U70632 ( .A(n50366), .B(n50365), .Z(n55531) );
  NOR U70633 ( .A(n50372), .B(n50367), .Z(n50368) );
  IV U70634 ( .A(n50368), .Z(n50369) );
  NOR U70635 ( .A(n50370), .B(n50369), .Z(n55533) );
  NOR U70636 ( .A(n55531), .B(n55533), .Z(n52949) );
  IV U70637 ( .A(n50370), .Z(n50375) );
  NOR U70638 ( .A(n50372), .B(n50371), .Z(n50373) );
  IV U70639 ( .A(n50373), .Z(n50374) );
  NOR U70640 ( .A(n50375), .B(n50374), .Z(n55536) );
  IV U70641 ( .A(n50376), .Z(n50380) );
  NOR U70642 ( .A(n50378), .B(n50377), .Z(n50379) );
  IV U70643 ( .A(n50379), .Z(n50382) );
  NOR U70644 ( .A(n50380), .B(n50382), .Z(n58101) );
  NOR U70645 ( .A(n55536), .B(n58101), .Z(n52948) );
  IV U70646 ( .A(n50381), .Z(n50383) );
  NOR U70647 ( .A(n50383), .B(n50382), .Z(n58098) );
  IV U70648 ( .A(n50384), .Z(n50388) );
  NOR U70649 ( .A(n50386), .B(n50385), .Z(n50387) );
  IV U70650 ( .A(n50387), .Z(n50390) );
  NOR U70651 ( .A(n50388), .B(n50390), .Z(n55541) );
  IV U70652 ( .A(n50389), .Z(n50391) );
  NOR U70653 ( .A(n50391), .B(n50390), .Z(n55538) );
  IV U70654 ( .A(n50392), .Z(n50396) );
  IV U70655 ( .A(n50393), .Z(n52941) );
  NOR U70656 ( .A(n50394), .B(n52941), .Z(n50395) );
  IV U70657 ( .A(n50395), .Z(n52946) );
  NOR U70658 ( .A(n50396), .B(n52946), .Z(n58094) );
  IV U70659 ( .A(n50397), .Z(n50404) );
  NOR U70660 ( .A(n50404), .B(n50398), .Z(n55558) );
  IV U70661 ( .A(n50399), .Z(n50401) );
  NOR U70662 ( .A(n50401), .B(n50400), .Z(n55555) );
  NOR U70663 ( .A(n55558), .B(n55555), .Z(n52937) );
  IV U70664 ( .A(n50402), .Z(n50403) );
  NOR U70665 ( .A(n50404), .B(n50403), .Z(n55553) );
  IV U70666 ( .A(n50405), .Z(n50409) );
  NOR U70667 ( .A(n52935), .B(n50406), .Z(n50407) );
  IV U70668 ( .A(n50407), .Z(n50408) );
  NOR U70669 ( .A(n50409), .B(n50408), .Z(n58085) );
  NOR U70670 ( .A(n52909), .B(n50410), .Z(n50411) );
  IV U70671 ( .A(n50411), .Z(n55581) );
  NOR U70672 ( .A(n55581), .B(n50412), .Z(n52899) );
  IV U70673 ( .A(n50413), .Z(n50416) );
  NOR U70674 ( .A(n50414), .B(n55593), .Z(n50415) );
  IV U70675 ( .A(n50415), .Z(n50418) );
  NOR U70676 ( .A(n50416), .B(n50418), .Z(n55588) );
  IV U70677 ( .A(n50417), .Z(n50419) );
  NOR U70678 ( .A(n50419), .B(n50418), .Z(n55585) );
  NOR U70679 ( .A(n55593), .B(n50420), .Z(n52898) );
  IV U70680 ( .A(n50421), .Z(n50422) );
  NOR U70681 ( .A(n50423), .B(n50422), .Z(n50424) );
  IV U70682 ( .A(n50424), .Z(n55601) );
  NOR U70683 ( .A(n55601), .B(n50425), .Z(n52897) );
  NOR U70684 ( .A(n50427), .B(n50426), .Z(n50428) );
  IV U70685 ( .A(n50428), .Z(n55607) );
  NOR U70686 ( .A(n55607), .B(n50429), .Z(n52896) );
  IV U70687 ( .A(n50430), .Z(n50435) );
  XOR U70688 ( .A(n50431), .B(n52889), .Z(n50432) );
  NOR U70689 ( .A(n50433), .B(n50432), .Z(n50434) );
  IV U70690 ( .A(n50434), .Z(n50437) );
  NOR U70691 ( .A(n50435), .B(n50437), .Z(n55612) );
  IV U70692 ( .A(n50436), .Z(n50438) );
  NOR U70693 ( .A(n50438), .B(n50437), .Z(n55617) );
  IV U70694 ( .A(n50439), .Z(n50441) );
  NOR U70695 ( .A(n50441), .B(n50440), .Z(n55619) );
  XOR U70696 ( .A(n55617), .B(n55619), .Z(n50442) );
  NOR U70697 ( .A(n55612), .B(n50442), .Z(n52895) );
  IV U70698 ( .A(n50443), .Z(n50446) );
  NOR U70699 ( .A(n50444), .B(n50449), .Z(n50445) );
  IV U70700 ( .A(n50445), .Z(n52892) );
  NOR U70701 ( .A(n50446), .B(n52892), .Z(n58060) );
  IV U70702 ( .A(n50447), .Z(n50448) );
  NOR U70703 ( .A(n50449), .B(n50448), .Z(n52885) );
  IV U70704 ( .A(n52885), .Z(n52876) );
  IV U70705 ( .A(n50450), .Z(n50452) );
  NOR U70706 ( .A(n50452), .B(n50451), .Z(n60864) );
  IV U70707 ( .A(n50453), .Z(n50454) );
  NOR U70708 ( .A(n50454), .B(n52870), .Z(n63304) );
  NOR U70709 ( .A(n60864), .B(n63304), .Z(n58054) );
  IV U70710 ( .A(n50455), .Z(n50456) );
  NOR U70711 ( .A(n50457), .B(n50456), .Z(n58050) );
  IV U70712 ( .A(n50458), .Z(n50459) );
  NOR U70713 ( .A(n50459), .B(n52861), .Z(n58047) );
  IV U70714 ( .A(n50460), .Z(n50465) );
  IV U70715 ( .A(n50461), .Z(n50462) );
  NOR U70716 ( .A(n50465), .B(n50462), .Z(n55636) );
  IV U70717 ( .A(n50463), .Z(n50467) );
  NOR U70718 ( .A(n50465), .B(n50464), .Z(n50466) );
  IV U70719 ( .A(n50466), .Z(n50469) );
  NOR U70720 ( .A(n50467), .B(n50469), .Z(n58042) );
  NOR U70721 ( .A(n55636), .B(n58042), .Z(n52859) );
  IV U70722 ( .A(n50468), .Z(n50470) );
  NOR U70723 ( .A(n50470), .B(n50469), .Z(n58039) );
  NOR U70724 ( .A(n50471), .B(n50478), .Z(n50472) );
  IV U70725 ( .A(n50472), .Z(n55639) );
  NOR U70726 ( .A(n55639), .B(n50473), .Z(n52858) );
  IV U70727 ( .A(n50474), .Z(n50475) );
  NOR U70728 ( .A(n50478), .B(n50475), .Z(n58029) );
  IV U70729 ( .A(n50476), .Z(n50477) );
  NOR U70730 ( .A(n50478), .B(n50477), .Z(n52852) );
  IV U70731 ( .A(n50479), .Z(n50481) );
  NOR U70732 ( .A(n50481), .B(n50480), .Z(n52849) );
  IV U70733 ( .A(n52849), .Z(n52840) );
  IV U70734 ( .A(n50482), .Z(n50484) );
  NOR U70735 ( .A(n50484), .B(n50483), .Z(n58020) );
  NOR U70736 ( .A(n55649), .B(n58020), .Z(n52838) );
  NOR U70737 ( .A(n50486), .B(n50485), .Z(n55646) );
  IV U70738 ( .A(n50487), .Z(n50488) );
  NOR U70739 ( .A(n50488), .B(n50490), .Z(n55652) );
  IV U70740 ( .A(n50489), .Z(n50491) );
  NOR U70741 ( .A(n50491), .B(n50490), .Z(n55654) );
  NOR U70742 ( .A(n55652), .B(n55654), .Z(n52837) );
  IV U70743 ( .A(n50492), .Z(n50493) );
  NOR U70744 ( .A(n50494), .B(n50493), .Z(n55657) );
  IV U70745 ( .A(n50495), .Z(n50498) );
  NOR U70746 ( .A(n50504), .B(n50496), .Z(n50497) );
  IV U70747 ( .A(n50497), .Z(n50500) );
  NOR U70748 ( .A(n50498), .B(n50500), .Z(n55662) );
  NOR U70749 ( .A(n55657), .B(n55662), .Z(n52836) );
  IV U70750 ( .A(n50499), .Z(n50501) );
  NOR U70751 ( .A(n50501), .B(n50500), .Z(n55659) );
  IV U70752 ( .A(n50502), .Z(n50506) );
  NOR U70753 ( .A(n50504), .B(n50503), .Z(n50505) );
  IV U70754 ( .A(n50505), .Z(n52830) );
  NOR U70755 ( .A(n50506), .B(n52830), .Z(n50507) );
  IV U70756 ( .A(n50507), .Z(n58015) );
  IV U70757 ( .A(n50508), .Z(n50513) );
  IV U70758 ( .A(n50509), .Z(n50510) );
  NOR U70759 ( .A(n50511), .B(n50510), .Z(n50512) );
  IV U70760 ( .A(n50512), .Z(n52833) );
  NOR U70761 ( .A(n50513), .B(n52833), .Z(n50514) );
  IV U70762 ( .A(n50514), .Z(n58005) );
  IV U70763 ( .A(n50515), .Z(n50516) );
  NOR U70764 ( .A(n50517), .B(n50516), .Z(n58000) );
  NOR U70765 ( .A(n57999), .B(n58000), .Z(n52828) );
  IV U70766 ( .A(n50518), .Z(n50519) );
  NOR U70767 ( .A(n50519), .B(n55670), .Z(n55665) );
  NOR U70768 ( .A(n50520), .B(n55667), .Z(n50521) );
  NOR U70769 ( .A(n55665), .B(n50521), .Z(n52827) );
  IV U70770 ( .A(n50522), .Z(n50523) );
  NOR U70771 ( .A(n50524), .B(n50523), .Z(n57990) );
  IV U70772 ( .A(n50525), .Z(n50528) );
  IV U70773 ( .A(n50526), .Z(n50527) );
  NOR U70774 ( .A(n50528), .B(n50527), .Z(n55677) );
  XOR U70775 ( .A(n50529), .B(n52810), .Z(n50531) );
  NOR U70776 ( .A(n50531), .B(n50530), .Z(n50532) );
  IV U70777 ( .A(n50532), .Z(n55681) );
  NOR U70778 ( .A(n55681), .B(n50533), .Z(n52821) );
  IV U70779 ( .A(n50534), .Z(n50537) );
  NOR U70780 ( .A(n50535), .B(n50540), .Z(n50536) );
  IV U70781 ( .A(n50536), .Z(n52814) );
  NOR U70782 ( .A(n50537), .B(n52814), .Z(n55685) );
  IV U70783 ( .A(n50538), .Z(n50539) );
  NOR U70784 ( .A(n50540), .B(n50539), .Z(n57969) );
  IV U70785 ( .A(n50541), .Z(n50546) );
  IV U70786 ( .A(n50542), .Z(n50543) );
  NOR U70787 ( .A(n50546), .B(n50543), .Z(n55687) );
  IV U70788 ( .A(n50544), .Z(n50545) );
  NOR U70789 ( .A(n50546), .B(n50545), .Z(n55693) );
  IV U70790 ( .A(n50547), .Z(n52806) );
  NOR U70791 ( .A(n52806), .B(n50548), .Z(n55690) );
  IV U70792 ( .A(n50549), .Z(n50552) );
  NOR U70793 ( .A(n50550), .B(n52806), .Z(n50551) );
  IV U70794 ( .A(n50551), .Z(n52803) );
  NOR U70795 ( .A(n50552), .B(n52803), .Z(n55696) );
  IV U70796 ( .A(n50553), .Z(n50554) );
  NOR U70797 ( .A(n50554), .B(n50557), .Z(n57958) );
  IV U70798 ( .A(n50555), .Z(n50556) );
  NOR U70799 ( .A(n50557), .B(n50556), .Z(n55702) );
  IV U70800 ( .A(n50558), .Z(n50559) );
  NOR U70801 ( .A(n50560), .B(n50559), .Z(n55705) );
  IV U70802 ( .A(n50561), .Z(n50562) );
  NOR U70803 ( .A(n50562), .B(n52797), .Z(n55707) );
  NOR U70804 ( .A(n55705), .B(n55707), .Z(n52800) );
  IV U70805 ( .A(n50563), .Z(n50564) );
  NOR U70806 ( .A(n50565), .B(n50564), .Z(n55717) );
  IV U70807 ( .A(n50566), .Z(n50570) );
  NOR U70808 ( .A(n50568), .B(n50567), .Z(n50569) );
  IV U70809 ( .A(n50569), .Z(n50572) );
  NOR U70810 ( .A(n50570), .B(n50572), .Z(n55719) );
  NOR U70811 ( .A(n55717), .B(n55719), .Z(n52794) );
  IV U70812 ( .A(n50571), .Z(n50573) );
  NOR U70813 ( .A(n50573), .B(n50572), .Z(n57952) );
  IV U70814 ( .A(n50574), .Z(n52788) );
  NOR U70815 ( .A(n52788), .B(n50575), .Z(n52785) );
  IV U70816 ( .A(n52785), .Z(n52776) );
  IV U70817 ( .A(n50576), .Z(n50578) );
  NOR U70818 ( .A(n50578), .B(n50577), .Z(n55727) );
  IV U70819 ( .A(n50579), .Z(n50580) );
  NOR U70820 ( .A(n52733), .B(n50580), .Z(n50581) );
  IV U70821 ( .A(n50581), .Z(n57915) );
  IV U70822 ( .A(n50582), .Z(n50583) );
  NOR U70823 ( .A(n50584), .B(n50583), .Z(n57911) );
  IV U70824 ( .A(n50585), .Z(n50586) );
  NOR U70825 ( .A(n50587), .B(n50586), .Z(n57917) );
  NOR U70826 ( .A(n57911), .B(n57917), .Z(n52732) );
  IV U70827 ( .A(n50588), .Z(n50590) );
  NOR U70828 ( .A(n50590), .B(n50589), .Z(n55759) );
  IV U70829 ( .A(n50591), .Z(n50592) );
  NOR U70830 ( .A(n50592), .B(n50596), .Z(n50593) );
  IV U70831 ( .A(n50593), .Z(n57907) );
  IV U70832 ( .A(n50594), .Z(n50595) );
  NOR U70833 ( .A(n50596), .B(n50595), .Z(n57903) );
  IV U70834 ( .A(n50597), .Z(n50598) );
  NOR U70835 ( .A(n50599), .B(n50598), .Z(n55776) );
  IV U70836 ( .A(n50600), .Z(n50603) );
  IV U70837 ( .A(n50601), .Z(n50602) );
  NOR U70838 ( .A(n50603), .B(n50602), .Z(n55778) );
  NOR U70839 ( .A(n55776), .B(n55778), .Z(n52719) );
  IV U70840 ( .A(n50604), .Z(n50605) );
  NOR U70841 ( .A(n50605), .B(n52714), .Z(n57897) );
  NOR U70842 ( .A(n50607), .B(n50606), .Z(n55786) );
  NOR U70843 ( .A(n57897), .B(n55786), .Z(n50608) );
  IV U70844 ( .A(n50608), .Z(n52713) );
  IV U70845 ( .A(n50609), .Z(n50610) );
  NOR U70846 ( .A(n50611), .B(n50610), .Z(n57900) );
  IV U70847 ( .A(n50612), .Z(n50613) );
  NOR U70848 ( .A(n52703), .B(n50613), .Z(n55791) );
  NOR U70849 ( .A(n57900), .B(n55791), .Z(n52712) );
  IV U70850 ( .A(n50614), .Z(n50616) );
  NOR U70851 ( .A(n50616), .B(n50615), .Z(n52709) );
  IV U70852 ( .A(n50617), .Z(n50622) );
  IV U70853 ( .A(n50618), .Z(n50619) );
  NOR U70854 ( .A(n50620), .B(n50619), .Z(n50621) );
  IV U70855 ( .A(n50621), .Z(n52705) );
  NOR U70856 ( .A(n50622), .B(n52705), .Z(n57885) );
  IV U70857 ( .A(n50623), .Z(n50624) );
  NOR U70858 ( .A(n50624), .B(n50630), .Z(n57865) );
  IV U70859 ( .A(n50625), .Z(n50628) );
  NOR U70860 ( .A(n50631), .B(n50638), .Z(n50626) );
  IV U70861 ( .A(n50626), .Z(n50627) );
  NOR U70862 ( .A(n50628), .B(n50627), .Z(n57869) );
  IV U70863 ( .A(n50629), .Z(n50634) );
  NOR U70864 ( .A(n50631), .B(n50630), .Z(n50632) );
  IV U70865 ( .A(n50632), .Z(n50633) );
  NOR U70866 ( .A(n50634), .B(n50633), .Z(n57857) );
  IV U70867 ( .A(n50635), .Z(n55798) );
  NOR U70868 ( .A(n50636), .B(n55798), .Z(n50640) );
  IV U70869 ( .A(n50637), .Z(n50639) );
  NOR U70870 ( .A(n50639), .B(n50638), .Z(n57860) );
  NOR U70871 ( .A(n50640), .B(n57860), .Z(n52690) );
  IV U70872 ( .A(n50641), .Z(n55795) );
  IV U70873 ( .A(n50642), .Z(n50643) );
  NOR U70874 ( .A(n50646), .B(n50643), .Z(n55803) );
  NOR U70875 ( .A(n55801), .B(n55803), .Z(n52689) );
  IV U70876 ( .A(n50644), .Z(n50645) );
  NOR U70877 ( .A(n50646), .B(n50645), .Z(n55811) );
  IV U70878 ( .A(n50647), .Z(n50649) );
  NOR U70879 ( .A(n50649), .B(n50648), .Z(n55806) );
  NOR U70880 ( .A(n55811), .B(n55806), .Z(n52688) );
  IV U70881 ( .A(n50650), .Z(n50652) );
  NOR U70882 ( .A(n50652), .B(n50651), .Z(n60989) );
  IV U70883 ( .A(n50653), .Z(n50654) );
  NOR U70884 ( .A(n50654), .B(n63050), .Z(n63043) );
  NOR U70885 ( .A(n60989), .B(n63043), .Z(n55819) );
  IV U70886 ( .A(n50655), .Z(n50657) );
  IV U70887 ( .A(n50656), .Z(n50661) );
  NOR U70888 ( .A(n50657), .B(n50661), .Z(n60998) );
  IV U70889 ( .A(n50658), .Z(n50659) );
  NOR U70890 ( .A(n50659), .B(n50661), .Z(n60993) );
  NOR U70891 ( .A(n60998), .B(n60993), .Z(n55824) );
  IV U70892 ( .A(n50660), .Z(n55828) );
  NOR U70893 ( .A(n50661), .B(n55828), .Z(n52679) );
  IV U70894 ( .A(n50662), .Z(n50664) );
  NOR U70895 ( .A(n50664), .B(n50663), .Z(n55837) );
  IV U70896 ( .A(n50665), .Z(n50666) );
  NOR U70897 ( .A(n55825), .B(n50666), .Z(n55831) );
  NOR U70898 ( .A(n55837), .B(n55831), .Z(n52674) );
  IV U70899 ( .A(n50667), .Z(n50669) );
  NOR U70900 ( .A(n50669), .B(n50668), .Z(n55839) );
  IV U70901 ( .A(n50670), .Z(n50671) );
  NOR U70902 ( .A(n50672), .B(n50671), .Z(n50673) );
  IV U70903 ( .A(n50673), .Z(n52662) );
  IV U70904 ( .A(n50674), .Z(n50676) );
  NOR U70905 ( .A(n50676), .B(n50675), .Z(n55853) );
  IV U70906 ( .A(n50677), .Z(n50678) );
  NOR U70907 ( .A(n50679), .B(n50678), .Z(n57837) );
  NOR U70908 ( .A(n55853), .B(n57837), .Z(n52655) );
  IV U70909 ( .A(n50680), .Z(n50681) );
  NOR U70910 ( .A(n50682), .B(n50681), .Z(n55850) );
  IV U70911 ( .A(n50683), .Z(n50685) );
  XOR U70912 ( .A(n50691), .B(n50689), .Z(n50684) );
  NOR U70913 ( .A(n50685), .B(n50684), .Z(n55855) );
  NOR U70914 ( .A(n55850), .B(n55855), .Z(n52654) );
  IV U70915 ( .A(n50686), .Z(n50687) );
  NOR U70916 ( .A(n50689), .B(n50687), .Z(n57833) );
  IV U70917 ( .A(n50688), .Z(n50690) );
  NOR U70918 ( .A(n50690), .B(n50689), .Z(n57830) );
  IV U70919 ( .A(n50691), .Z(n50692) );
  NOR U70920 ( .A(n50692), .B(n55860), .Z(n52653) );
  NOR U70921 ( .A(n50693), .B(n55860), .Z(n55869) );
  IV U70922 ( .A(n50694), .Z(n50695) );
  NOR U70923 ( .A(n50695), .B(n52638), .Z(n52642) );
  IV U70924 ( .A(n50696), .Z(n50698) );
  NOR U70925 ( .A(n50698), .B(n50697), .Z(n55878) );
  NOR U70926 ( .A(n50700), .B(n50699), .Z(n55876) );
  NOR U70927 ( .A(n55878), .B(n55876), .Z(n52636) );
  IV U70928 ( .A(n50701), .Z(n61059) );
  NOR U70929 ( .A(n50702), .B(n61059), .Z(n55881) );
  NOR U70930 ( .A(n50703), .B(n50712), .Z(n50704) );
  IV U70931 ( .A(n50704), .Z(n50705) );
  NOR U70932 ( .A(n50706), .B(n50705), .Z(n55889) );
  IV U70933 ( .A(n50707), .Z(n50709) );
  NOR U70934 ( .A(n50709), .B(n50708), .Z(n55892) );
  IV U70935 ( .A(n50710), .Z(n50711) );
  NOR U70936 ( .A(n50712), .B(n50711), .Z(n55887) );
  NOR U70937 ( .A(n55892), .B(n55887), .Z(n50713) );
  IV U70938 ( .A(n50713), .Z(n52635) );
  IV U70939 ( .A(n50714), .Z(n50716) );
  NOR U70940 ( .A(n50716), .B(n50715), .Z(n57819) );
  IV U70941 ( .A(n50717), .Z(n50719) );
  NOR U70942 ( .A(n50719), .B(n50718), .Z(n55895) );
  NOR U70943 ( .A(n57819), .B(n55895), .Z(n52634) );
  IV U70944 ( .A(n50720), .Z(n50721) );
  NOR U70945 ( .A(n50721), .B(n50727), .Z(n57817) );
  IV U70946 ( .A(n50722), .Z(n50723) );
  NOR U70947 ( .A(n50724), .B(n50723), .Z(n57822) );
  NOR U70948 ( .A(n57817), .B(n57822), .Z(n52633) );
  IV U70949 ( .A(n50728), .Z(n50725) );
  NOR U70950 ( .A(n50725), .B(n50727), .Z(n55903) );
  IV U70951 ( .A(n50726), .Z(n50730) );
  XOR U70952 ( .A(n50728), .B(n50727), .Z(n50729) );
  NOR U70953 ( .A(n50730), .B(n50729), .Z(n55898) );
  NOR U70954 ( .A(n55903), .B(n55898), .Z(n52632) );
  IV U70955 ( .A(n50731), .Z(n50732) );
  NOR U70956 ( .A(n50732), .B(n50734), .Z(n55919) );
  IV U70957 ( .A(n50733), .Z(n50735) );
  NOR U70958 ( .A(n50735), .B(n50734), .Z(n55921) );
  NOR U70959 ( .A(n55919), .B(n55921), .Z(n52607) );
  IV U70960 ( .A(n50736), .Z(n50737) );
  NOR U70961 ( .A(n50737), .B(n57803), .Z(n55932) );
  IV U70962 ( .A(n50738), .Z(n50739) );
  NOR U70963 ( .A(n57803), .B(n50739), .Z(n55929) );
  IV U70964 ( .A(n50740), .Z(n50741) );
  NOR U70965 ( .A(n50742), .B(n50741), .Z(n55935) );
  IV U70966 ( .A(n50743), .Z(n50746) );
  IV U70967 ( .A(n50744), .Z(n50745) );
  NOR U70968 ( .A(n50746), .B(n50745), .Z(n55937) );
  NOR U70969 ( .A(n55935), .B(n55937), .Z(n52593) );
  IV U70970 ( .A(n50747), .Z(n50748) );
  NOR U70971 ( .A(n50748), .B(n50750), .Z(n57798) );
  IV U70972 ( .A(n50749), .Z(n50751) );
  NOR U70973 ( .A(n50751), .B(n50750), .Z(n57795) );
  IV U70974 ( .A(n50752), .Z(n50755) );
  NOR U70975 ( .A(n50764), .B(n50753), .Z(n50754) );
  IV U70976 ( .A(n50754), .Z(n50757) );
  NOR U70977 ( .A(n50755), .B(n50757), .Z(n57784) );
  IV U70978 ( .A(n50756), .Z(n50758) );
  NOR U70979 ( .A(n50758), .B(n50757), .Z(n55940) );
  IV U70980 ( .A(n50759), .Z(n50760) );
  NOR U70981 ( .A(n50764), .B(n50760), .Z(n50761) );
  IV U70982 ( .A(n50761), .Z(n50762) );
  NOR U70983 ( .A(n50763), .B(n50762), .Z(n57787) );
  IV U70984 ( .A(n50763), .Z(n50768) );
  NOR U70985 ( .A(n50765), .B(n50764), .Z(n50766) );
  IV U70986 ( .A(n50766), .Z(n50767) );
  NOR U70987 ( .A(n50768), .B(n50767), .Z(n57780) );
  IV U70988 ( .A(n50769), .Z(n50771) );
  NOR U70989 ( .A(n50771), .B(n50770), .Z(n57777) );
  IV U70990 ( .A(n50772), .Z(n50773) );
  NOR U70991 ( .A(n50776), .B(n50773), .Z(n55947) );
  IV U70992 ( .A(n50774), .Z(n50775) );
  NOR U70993 ( .A(n50776), .B(n50775), .Z(n50777) );
  IV U70994 ( .A(n50777), .Z(n50778) );
  NOR U70995 ( .A(n50779), .B(n50778), .Z(n55944) );
  IV U70996 ( .A(n50780), .Z(n50794) );
  XOR U70997 ( .A(n50794), .B(n50786), .Z(n50798) );
  XOR U70998 ( .A(n50796), .B(n50798), .Z(n50781) );
  NOR U70999 ( .A(n50782), .B(n50781), .Z(n50783) );
  IV U71000 ( .A(n50783), .Z(n57767) );
  NOR U71001 ( .A(n57767), .B(n50784), .Z(n52592) );
  IV U71002 ( .A(n50785), .Z(n50789) );
  IV U71003 ( .A(n50786), .Z(n50795) );
  NOR U71004 ( .A(n50787), .B(n50795), .Z(n50788) );
  IV U71005 ( .A(n50788), .Z(n50791) );
  NOR U71006 ( .A(n50789), .B(n50791), .Z(n57763) );
  IV U71007 ( .A(n50790), .Z(n50792) );
  NOR U71008 ( .A(n50792), .B(n50791), .Z(n50793) );
  IV U71009 ( .A(n50793), .Z(n55951) );
  NOR U71010 ( .A(n50795), .B(n50794), .Z(n55953) );
  IV U71011 ( .A(n50796), .Z(n50797) );
  NOR U71012 ( .A(n50798), .B(n50797), .Z(n57760) );
  NOR U71013 ( .A(n55953), .B(n57760), .Z(n52591) );
  NOR U71014 ( .A(n50800), .B(n50799), .Z(n55959) );
  NOR U71015 ( .A(n55955), .B(n55959), .Z(n52590) );
  IV U71016 ( .A(n50801), .Z(n50802) );
  NOR U71017 ( .A(n50802), .B(n50804), .Z(n55979) );
  IV U71018 ( .A(n50803), .Z(n50805) );
  NOR U71019 ( .A(n50805), .B(n50804), .Z(n55974) );
  NOR U71020 ( .A(n55979), .B(n55974), .Z(n52563) );
  IV U71021 ( .A(n50806), .Z(n50811) );
  IV U71022 ( .A(n50807), .Z(n50808) );
  NOR U71023 ( .A(n50811), .B(n50808), .Z(n57743) );
  IV U71024 ( .A(n50809), .Z(n50810) );
  NOR U71025 ( .A(n50811), .B(n50810), .Z(n57740) );
  IV U71026 ( .A(n50812), .Z(n50813) );
  NOR U71027 ( .A(n52560), .B(n50813), .Z(n55985) );
  IV U71028 ( .A(n50814), .Z(n50815) );
  NOR U71029 ( .A(n50815), .B(n52560), .Z(n55982) );
  IV U71030 ( .A(n50816), .Z(n50820) );
  NOR U71031 ( .A(n50817), .B(n52549), .Z(n50818) );
  IV U71032 ( .A(n50818), .Z(n50819) );
  NOR U71033 ( .A(n50820), .B(n50819), .Z(n50821) );
  IV U71034 ( .A(n50821), .Z(n57733) );
  IV U71035 ( .A(n50822), .Z(n50823) );
  NOR U71036 ( .A(n50824), .B(n50823), .Z(n50825) );
  IV U71037 ( .A(n50825), .Z(n56006) );
  IV U71038 ( .A(n50826), .Z(n50828) );
  NOR U71039 ( .A(n50828), .B(n50827), .Z(n56009) );
  IV U71040 ( .A(n50829), .Z(n50830) );
  NOR U71041 ( .A(n50830), .B(n50832), .Z(n57726) );
  NOR U71042 ( .A(n56009), .B(n57726), .Z(n52534) );
  IV U71043 ( .A(n50831), .Z(n50833) );
  NOR U71044 ( .A(n50833), .B(n50832), .Z(n57723) );
  IV U71045 ( .A(n50834), .Z(n50835) );
  NOR U71046 ( .A(n50836), .B(n50835), .Z(n56014) );
  IV U71047 ( .A(n50837), .Z(n50840) );
  IV U71048 ( .A(n50838), .Z(n50839) );
  NOR U71049 ( .A(n50840), .B(n50839), .Z(n56011) );
  IV U71050 ( .A(n50841), .Z(n50846) );
  IV U71051 ( .A(n50842), .Z(n50843) );
  NOR U71052 ( .A(n50844), .B(n50843), .Z(n50845) );
  IV U71053 ( .A(n50845), .Z(n50848) );
  NOR U71054 ( .A(n50846), .B(n50848), .Z(n57718) );
  IV U71055 ( .A(n50847), .Z(n50849) );
  NOR U71056 ( .A(n50849), .B(n50848), .Z(n57715) );
  IV U71057 ( .A(n50850), .Z(n50851) );
  NOR U71058 ( .A(n50852), .B(n50851), .Z(n56017) );
  IV U71059 ( .A(n50852), .Z(n50854) );
  NOR U71060 ( .A(n50854), .B(n50853), .Z(n56019) );
  NOR U71061 ( .A(n56017), .B(n56019), .Z(n52532) );
  IV U71062 ( .A(n50855), .Z(n50856) );
  NOR U71063 ( .A(n50857), .B(n50856), .Z(n52525) );
  IV U71064 ( .A(n50858), .Z(n50860) );
  NOR U71065 ( .A(n50860), .B(n50859), .Z(n50861) );
  IV U71066 ( .A(n50861), .Z(n56033) );
  IV U71067 ( .A(n50862), .Z(n61203) );
  NOR U71068 ( .A(n50863), .B(n61203), .Z(n50864) );
  NOR U71069 ( .A(n62893), .B(n50864), .Z(n56031) );
  NOR U71070 ( .A(n50866), .B(n50865), .Z(n57707) );
  IV U71071 ( .A(n50867), .Z(n50868) );
  NOR U71072 ( .A(n50869), .B(n50868), .Z(n56035) );
  NOR U71073 ( .A(n57707), .B(n56035), .Z(n52516) );
  IV U71074 ( .A(n50870), .Z(n50871) );
  NOR U71075 ( .A(n52510), .B(n50871), .Z(n56038) );
  IV U71076 ( .A(n50872), .Z(n50873) );
  NOR U71077 ( .A(n52510), .B(n50873), .Z(n56042) );
  NOR U71078 ( .A(n56038), .B(n56042), .Z(n52512) );
  IV U71079 ( .A(n50874), .Z(n50878) );
  NOR U71080 ( .A(n50876), .B(n50875), .Z(n50877) );
  IV U71081 ( .A(n50877), .Z(n52506) );
  NOR U71082 ( .A(n50878), .B(n52506), .Z(n56054) );
  IV U71083 ( .A(n50879), .Z(n50882) );
  IV U71084 ( .A(n50880), .Z(n50885) );
  XOR U71085 ( .A(n50883), .B(n50885), .Z(n50881) );
  NOR U71086 ( .A(n50882), .B(n50881), .Z(n56051) );
  IV U71087 ( .A(n50883), .Z(n62858) );
  NOR U71088 ( .A(n62858), .B(n50884), .Z(n56060) );
  NOR U71089 ( .A(n62858), .B(n50885), .Z(n56057) );
  IV U71090 ( .A(n50886), .Z(n50887) );
  NOR U71091 ( .A(n50888), .B(n50887), .Z(n57697) );
  IV U71092 ( .A(n50889), .Z(n50890) );
  NOR U71093 ( .A(n50890), .B(n50892), .Z(n68276) );
  IV U71094 ( .A(n50891), .Z(n50893) );
  NOR U71095 ( .A(n50893), .B(n50892), .Z(n57696) );
  NOR U71096 ( .A(n68276), .B(n57696), .Z(n52503) );
  IV U71097 ( .A(n50894), .Z(n50895) );
  NOR U71098 ( .A(n50895), .B(n52500), .Z(n56064) );
  IV U71099 ( .A(n50896), .Z(n50897) );
  NOR U71100 ( .A(n50901), .B(n50897), .Z(n50898) );
  IV U71101 ( .A(n50898), .Z(n57684) );
  NOR U71102 ( .A(n50899), .B(n50901), .Z(n61216) );
  IV U71103 ( .A(n50900), .Z(n50902) );
  NOR U71104 ( .A(n50902), .B(n50901), .Z(n61207) );
  NOR U71105 ( .A(n61216), .B(n61207), .Z(n56068) );
  IV U71106 ( .A(n50903), .Z(n50904) );
  NOR U71107 ( .A(n50905), .B(n50904), .Z(n56069) );
  IV U71108 ( .A(n50906), .Z(n50908) );
  IV U71109 ( .A(n50907), .Z(n52492) );
  NOR U71110 ( .A(n50908), .B(n52492), .Z(n56071) );
  NOR U71111 ( .A(n56069), .B(n56071), .Z(n52495) );
  IV U71112 ( .A(n50909), .Z(n50910) );
  NOR U71113 ( .A(n50910), .B(n50915), .Z(n57672) );
  IV U71114 ( .A(n50911), .Z(n50912) );
  NOR U71115 ( .A(n50913), .B(n50912), .Z(n56079) );
  IV U71116 ( .A(n50914), .Z(n50916) );
  NOR U71117 ( .A(n50916), .B(n50915), .Z(n56074) );
  NOR U71118 ( .A(n56079), .B(n56074), .Z(n50917) );
  IV U71119 ( .A(n50917), .Z(n52490) );
  IV U71120 ( .A(n50918), .Z(n50919) );
  NOR U71121 ( .A(n50920), .B(n50919), .Z(n56077) );
  IV U71122 ( .A(n50921), .Z(n50923) );
  IV U71123 ( .A(n50922), .Z(n50924) );
  NOR U71124 ( .A(n50923), .B(n50924), .Z(n57665) );
  NOR U71125 ( .A(n56077), .B(n57665), .Z(n52489) );
  NOR U71126 ( .A(n50925), .B(n50924), .Z(n50926) );
  IV U71127 ( .A(n50926), .Z(n56083) );
  NOR U71128 ( .A(n50927), .B(n56083), .Z(n50930) );
  IV U71129 ( .A(n50928), .Z(n50929) );
  NOR U71130 ( .A(n50929), .B(n52484), .Z(n56086) );
  NOR U71131 ( .A(n50930), .B(n56086), .Z(n52488) );
  IV U71132 ( .A(n50931), .Z(n50933) );
  XOR U71133 ( .A(n52483), .B(n52484), .Z(n50932) );
  NOR U71134 ( .A(n50933), .B(n50932), .Z(n56090) );
  IV U71135 ( .A(n50934), .Z(n57647) );
  IV U71136 ( .A(n50935), .Z(n50936) );
  NOR U71137 ( .A(n57647), .B(n50936), .Z(n56110) );
  IV U71138 ( .A(n50937), .Z(n50938) );
  NOR U71139 ( .A(n57647), .B(n50938), .Z(n56115) );
  IV U71140 ( .A(n50939), .Z(n50940) );
  NOR U71141 ( .A(n50940), .B(n56120), .Z(n57641) );
  IV U71142 ( .A(n50941), .Z(n50942) );
  NOR U71143 ( .A(n50942), .B(n56120), .Z(n57638) );
  IV U71144 ( .A(n50943), .Z(n50944) );
  NOR U71145 ( .A(n50945), .B(n50944), .Z(n56129) );
  IV U71146 ( .A(n50946), .Z(n50947) );
  NOR U71147 ( .A(n50947), .B(n56120), .Z(n50948) );
  NOR U71148 ( .A(n56129), .B(n50948), .Z(n52461) );
  IV U71149 ( .A(n50949), .Z(n50950) );
  NOR U71150 ( .A(n50950), .B(n50959), .Z(n57629) );
  IV U71151 ( .A(n50951), .Z(n50953) );
  NOR U71152 ( .A(n50953), .B(n50952), .Z(n57623) );
  NOR U71153 ( .A(n57629), .B(n57623), .Z(n52446) );
  IV U71154 ( .A(n50954), .Z(n50956) );
  NOR U71155 ( .A(n50956), .B(n50955), .Z(n62785) );
  IV U71156 ( .A(n50957), .Z(n50958) );
  NOR U71157 ( .A(n50959), .B(n50958), .Z(n62798) );
  NOR U71158 ( .A(n62785), .B(n62798), .Z(n57619) );
  IV U71159 ( .A(n50960), .Z(n50961) );
  NOR U71160 ( .A(n57615), .B(n50961), .Z(n50965) );
  IV U71161 ( .A(n50962), .Z(n50964) );
  NOR U71162 ( .A(n50964), .B(n50963), .Z(n56136) );
  NOR U71163 ( .A(n50965), .B(n56136), .Z(n52445) );
  IV U71164 ( .A(n50966), .Z(n50967) );
  NOR U71165 ( .A(n50967), .B(n57612), .Z(n57608) );
  IV U71166 ( .A(n50968), .Z(n50969) );
  NOR U71167 ( .A(n50970), .B(n50969), .Z(n57597) );
  IV U71168 ( .A(n50971), .Z(n50973) );
  NOR U71169 ( .A(n50973), .B(n50972), .Z(n61297) );
  IV U71170 ( .A(n50974), .Z(n50975) );
  NOR U71171 ( .A(n50975), .B(n52437), .Z(n62770) );
  NOR U71172 ( .A(n61297), .B(n62770), .Z(n57596) );
  IV U71173 ( .A(n57596), .Z(n52435) );
  IV U71174 ( .A(n50976), .Z(n50981) );
  IV U71175 ( .A(n50977), .Z(n50978) );
  NOR U71176 ( .A(n50981), .B(n50978), .Z(n56141) );
  IV U71177 ( .A(n50979), .Z(n50983) );
  NOR U71178 ( .A(n50981), .B(n50980), .Z(n50982) );
  IV U71179 ( .A(n50982), .Z(n50985) );
  NOR U71180 ( .A(n50983), .B(n50985), .Z(n56138) );
  IV U71181 ( .A(n50984), .Z(n50986) );
  NOR U71182 ( .A(n50986), .B(n50985), .Z(n57585) );
  NOR U71183 ( .A(n50988), .B(n50987), .Z(n50989) );
  IV U71184 ( .A(n50989), .Z(n57580) );
  NOR U71185 ( .A(n57580), .B(n50990), .Z(n52434) );
  IV U71186 ( .A(n50991), .Z(n50995) );
  NOR U71187 ( .A(n50993), .B(n50992), .Z(n50994) );
  IV U71188 ( .A(n50994), .Z(n50997) );
  NOR U71189 ( .A(n50995), .B(n50997), .Z(n57576) );
  IV U71190 ( .A(n50996), .Z(n50998) );
  NOR U71191 ( .A(n50998), .B(n50997), .Z(n57571) );
  IV U71192 ( .A(n50999), .Z(n51000) );
  NOR U71193 ( .A(n51000), .B(n56146), .Z(n52429) );
  IV U71194 ( .A(n51001), .Z(n51002) );
  NOR U71195 ( .A(n56146), .B(n51002), .Z(n56153) );
  IV U71196 ( .A(n51003), .Z(n51004) );
  NOR U71197 ( .A(n51006), .B(n51004), .Z(n57562) );
  IV U71198 ( .A(n51005), .Z(n51007) );
  NOR U71199 ( .A(n51007), .B(n51006), .Z(n57564) );
  XOR U71200 ( .A(n57562), .B(n57564), .Z(n51008) );
  NOR U71201 ( .A(n56153), .B(n51008), .Z(n52428) );
  IV U71202 ( .A(n51009), .Z(n56172) );
  NOR U71203 ( .A(n56172), .B(n51010), .Z(n52420) );
  IV U71204 ( .A(n51011), .Z(n51015) );
  NOR U71205 ( .A(n51013), .B(n51012), .Z(n51014) );
  IV U71206 ( .A(n51014), .Z(n52391) );
  NOR U71207 ( .A(n51015), .B(n52391), .Z(n56204) );
  IV U71208 ( .A(n51016), .Z(n51019) );
  NOR U71209 ( .A(n51017), .B(n51027), .Z(n51018) );
  IV U71210 ( .A(n51018), .Z(n51021) );
  NOR U71211 ( .A(n51019), .B(n51021), .Z(n56214) );
  IV U71212 ( .A(n51020), .Z(n51022) );
  NOR U71213 ( .A(n51022), .B(n51021), .Z(n56211) );
  IV U71214 ( .A(n51023), .Z(n51025) );
  IV U71215 ( .A(n51024), .Z(n56222) );
  NOR U71216 ( .A(n51025), .B(n56222), .Z(n56217) );
  IV U71217 ( .A(n51026), .Z(n56225) );
  NOR U71218 ( .A(n56225), .B(n51027), .Z(n51028) );
  NOR U71219 ( .A(n56217), .B(n51028), .Z(n52389) );
  IV U71220 ( .A(n51029), .Z(n51030) );
  NOR U71221 ( .A(n51031), .B(n51030), .Z(n56226) );
  NOR U71222 ( .A(n56226), .B(n56228), .Z(n51032) );
  IV U71223 ( .A(n51032), .Z(n51035) );
  IV U71224 ( .A(n51033), .Z(n51034) );
  NOR U71225 ( .A(n56222), .B(n51034), .Z(n57555) );
  NOR U71226 ( .A(n51035), .B(n57555), .Z(n52388) );
  IV U71227 ( .A(n51036), .Z(n51037) );
  NOR U71228 ( .A(n51038), .B(n51037), .Z(n56234) );
  NOR U71229 ( .A(n51040), .B(n51039), .Z(n56230) );
  NOR U71230 ( .A(n56234), .B(n56230), .Z(n52387) );
  IV U71231 ( .A(n51041), .Z(n51042) );
  NOR U71232 ( .A(n52377), .B(n51042), .Z(n56245) );
  IV U71233 ( .A(n51043), .Z(n52375) );
  NOR U71234 ( .A(n51044), .B(n52375), .Z(n57543) );
  NOR U71235 ( .A(n57532), .B(n57543), .Z(n52372) );
  IV U71236 ( .A(n51045), .Z(n51046) );
  NOR U71237 ( .A(n57540), .B(n51046), .Z(n57528) );
  NOR U71238 ( .A(n57523), .B(n57528), .Z(n51047) );
  IV U71239 ( .A(n51047), .Z(n51052) );
  IV U71240 ( .A(n51048), .Z(n51051) );
  IV U71241 ( .A(n51049), .Z(n51050) );
  NOR U71242 ( .A(n51051), .B(n51050), .Z(n57526) );
  NOR U71243 ( .A(n51052), .B(n57526), .Z(n52371) );
  IV U71244 ( .A(n51053), .Z(n51057) );
  NOR U71245 ( .A(n51054), .B(n52361), .Z(n51055) );
  IV U71246 ( .A(n51055), .Z(n51056) );
  NOR U71247 ( .A(n51057), .B(n51056), .Z(n57520) );
  NOR U71248 ( .A(n51059), .B(n51058), .Z(n51060) );
  IV U71249 ( .A(n51060), .Z(n51061) );
  NOR U71250 ( .A(n51062), .B(n51061), .Z(n57511) );
  IV U71251 ( .A(n51063), .Z(n51064) );
  NOR U71252 ( .A(n51067), .B(n51064), .Z(n68093) );
  IV U71253 ( .A(n51065), .Z(n51066) );
  NOR U71254 ( .A(n51067), .B(n51066), .Z(n57510) );
  NOR U71255 ( .A(n68093), .B(n57510), .Z(n52356) );
  IV U71256 ( .A(n51068), .Z(n51072) );
  NOR U71257 ( .A(n51070), .B(n51069), .Z(n51071) );
  IV U71258 ( .A(n51071), .Z(n52354) );
  NOR U71259 ( .A(n51072), .B(n52354), .Z(n52350) );
  IV U71260 ( .A(n52350), .Z(n52344) );
  IV U71261 ( .A(n51073), .Z(n51077) );
  IV U71262 ( .A(n51074), .Z(n51079) );
  NOR U71263 ( .A(n51075), .B(n51079), .Z(n51076) );
  IV U71264 ( .A(n51076), .Z(n52346) );
  NOR U71265 ( .A(n51077), .B(n52346), .Z(n56270) );
  NOR U71266 ( .A(n51079), .B(n51078), .Z(n56267) );
  IV U71267 ( .A(n51080), .Z(n51083) );
  IV U71268 ( .A(n51081), .Z(n51082) );
  NOR U71269 ( .A(n51083), .B(n51082), .Z(n56274) );
  XOR U71270 ( .A(n61363), .B(n57505), .Z(n51084) );
  NOR U71271 ( .A(n56273), .B(n51084), .Z(n51085) );
  IV U71272 ( .A(n51085), .Z(n52342) );
  IV U71273 ( .A(n51086), .Z(n51087) );
  NOR U71274 ( .A(n51088), .B(n51087), .Z(n61375) );
  IV U71275 ( .A(n51089), .Z(n51092) );
  NOR U71276 ( .A(n52331), .B(n51090), .Z(n51091) );
  IV U71277 ( .A(n51091), .Z(n52335) );
  NOR U71278 ( .A(n51092), .B(n52335), .Z(n62611) );
  NOR U71279 ( .A(n61375), .B(n62611), .Z(n56286) );
  IV U71280 ( .A(n56286), .Z(n51096) );
  IV U71281 ( .A(n51093), .Z(n51095) );
  NOR U71282 ( .A(n51095), .B(n51094), .Z(n56278) );
  NOR U71283 ( .A(n51096), .B(n56278), .Z(n52341) );
  NOR U71284 ( .A(n51097), .B(n51104), .Z(n57493) );
  IV U71285 ( .A(n51098), .Z(n51099) );
  NOR U71286 ( .A(n51099), .B(n51104), .Z(n57490) );
  IV U71287 ( .A(n51100), .Z(n51101) );
  NOR U71288 ( .A(n51102), .B(n51101), .Z(n56299) );
  IV U71289 ( .A(n51103), .Z(n51105) );
  NOR U71290 ( .A(n51105), .B(n51104), .Z(n56296) );
  NOR U71291 ( .A(n56299), .B(n56296), .Z(n52326) );
  IV U71292 ( .A(n51106), .Z(n51107) );
  NOR U71293 ( .A(n51107), .B(n52323), .Z(n57487) );
  IV U71294 ( .A(n51108), .Z(n52315) );
  IV U71295 ( .A(n51109), .Z(n51110) );
  NOR U71296 ( .A(n52315), .B(n51110), .Z(n51111) );
  IV U71297 ( .A(n51111), .Z(n57476) );
  IV U71298 ( .A(n51112), .Z(n51113) );
  NOR U71299 ( .A(n51114), .B(n51113), .Z(n57471) );
  IV U71300 ( .A(n51115), .Z(n51116) );
  NOR U71301 ( .A(n52304), .B(n51116), .Z(n57460) );
  IV U71302 ( .A(n51117), .Z(n51118) );
  NOR U71303 ( .A(n66966), .B(n51118), .Z(n62552) );
  IV U71304 ( .A(n51119), .Z(n51120) );
  NOR U71305 ( .A(n66966), .B(n51120), .Z(n61391) );
  NOR U71306 ( .A(n62552), .B(n61391), .Z(n57453) );
  IV U71307 ( .A(n51121), .Z(n51123) );
  NOR U71308 ( .A(n51123), .B(n51122), .Z(n57450) );
  IV U71309 ( .A(n51124), .Z(n51125) );
  NOR U71310 ( .A(n57432), .B(n51125), .Z(n52283) );
  IV U71311 ( .A(n51126), .Z(n51136) );
  NOR U71312 ( .A(n51128), .B(n51127), .Z(n51134) );
  IV U71313 ( .A(n51129), .Z(n57412) );
  XOR U71314 ( .A(n51144), .B(n57412), .Z(n51130) );
  NOR U71315 ( .A(n51131), .B(n51130), .Z(n51132) );
  IV U71316 ( .A(n51132), .Z(n51133) );
  NOR U71317 ( .A(n51134), .B(n51133), .Z(n51135) );
  IV U71318 ( .A(n51135), .Z(n52281) );
  NOR U71319 ( .A(n51136), .B(n52281), .Z(n57425) );
  IV U71320 ( .A(n51137), .Z(n51140) );
  NOR U71321 ( .A(n51138), .B(n57412), .Z(n51139) );
  IV U71322 ( .A(n51139), .Z(n51142) );
  NOR U71323 ( .A(n51140), .B(n51142), .Z(n56315) );
  IV U71324 ( .A(n51141), .Z(n51143) );
  NOR U71325 ( .A(n51143), .B(n51142), .Z(n56321) );
  IV U71326 ( .A(n51144), .Z(n51145) );
  NOR U71327 ( .A(n51145), .B(n57412), .Z(n57402) );
  IV U71328 ( .A(n51146), .Z(n51147) );
  NOR U71329 ( .A(n52269), .B(n51147), .Z(n56327) );
  IV U71330 ( .A(n51148), .Z(n51149) );
  NOR U71331 ( .A(n51150), .B(n51149), .Z(n51151) );
  IV U71332 ( .A(n51151), .Z(n52264) );
  NOR U71333 ( .A(n51152), .B(n52258), .Z(n51153) );
  IV U71334 ( .A(n51153), .Z(n51154) );
  NOR U71335 ( .A(n51155), .B(n51154), .Z(n56337) );
  IV U71336 ( .A(n51156), .Z(n51165) );
  IV U71337 ( .A(n51170), .Z(n51158) );
  NOR U71338 ( .A(n51158), .B(n51157), .Z(n51163) );
  NOR U71339 ( .A(n51160), .B(n51159), .Z(n51161) );
  IV U71340 ( .A(n51161), .Z(n51162) );
  NOR U71341 ( .A(n51163), .B(n51162), .Z(n51164) );
  IV U71342 ( .A(n51164), .Z(n51167) );
  NOR U71343 ( .A(n51165), .B(n51167), .Z(n56370) );
  IV U71344 ( .A(n51166), .Z(n51168) );
  NOR U71345 ( .A(n51168), .B(n51167), .Z(n56376) );
  IV U71346 ( .A(n51169), .Z(n51172) );
  NOR U71347 ( .A(n51170), .B(n51175), .Z(n51171) );
  IV U71348 ( .A(n51171), .Z(n52234) );
  NOR U71349 ( .A(n51172), .B(n52234), .Z(n57384) );
  IV U71350 ( .A(n51173), .Z(n51174) );
  NOR U71351 ( .A(n51175), .B(n51174), .Z(n56382) );
  IV U71352 ( .A(n51176), .Z(n51178) );
  IV U71353 ( .A(n51177), .Z(n51180) );
  NOR U71354 ( .A(n51178), .B(n51180), .Z(n56379) );
  IV U71355 ( .A(n51179), .Z(n57379) );
  NOR U71356 ( .A(n51180), .B(n57379), .Z(n51181) );
  NOR U71357 ( .A(n57377), .B(n51181), .Z(n52231) );
  NOR U71358 ( .A(n51183), .B(n51182), .Z(n56385) );
  IV U71359 ( .A(n51184), .Z(n51186) );
  NOR U71360 ( .A(n51186), .B(n51185), .Z(n57367) );
  IV U71361 ( .A(n51187), .Z(n51188) );
  NOR U71362 ( .A(n51188), .B(n51191), .Z(n57365) );
  NOR U71363 ( .A(n57367), .B(n57365), .Z(n52230) );
  IV U71364 ( .A(n51189), .Z(n57358) );
  NOR U71365 ( .A(n57358), .B(n57356), .Z(n51193) );
  IV U71366 ( .A(n51190), .Z(n57363) );
  NOR U71367 ( .A(n57363), .B(n51191), .Z(n51192) );
  NOR U71368 ( .A(n51193), .B(n51192), .Z(n52229) );
  IV U71369 ( .A(n51194), .Z(n51198) );
  IV U71370 ( .A(n51195), .Z(n51201) );
  NOR U71371 ( .A(n51201), .B(n51196), .Z(n51197) );
  IV U71372 ( .A(n51197), .Z(n52210) );
  NOR U71373 ( .A(n51198), .B(n52210), .Z(n56400) );
  IV U71374 ( .A(n51199), .Z(n51200) );
  NOR U71375 ( .A(n51201), .B(n51200), .Z(n56402) );
  NOR U71376 ( .A(n56400), .B(n56402), .Z(n52208) );
  IV U71377 ( .A(n51202), .Z(n51207) );
  NOR U71378 ( .A(n51217), .B(n51214), .Z(n51203) );
  XOR U71379 ( .A(n51212), .B(n51203), .Z(n51205) );
  NOR U71380 ( .A(n51205), .B(n51204), .Z(n51206) );
  IV U71381 ( .A(n51206), .Z(n51209) );
  NOR U71382 ( .A(n51207), .B(n51209), .Z(n56410) );
  IV U71383 ( .A(n51208), .Z(n51210) );
  NOR U71384 ( .A(n51210), .B(n51209), .Z(n56419) );
  IV U71385 ( .A(n51211), .Z(n51213) );
  IV U71386 ( .A(n51212), .Z(n51215) );
  NOR U71387 ( .A(n51213), .B(n51215), .Z(n56416) );
  IV U71388 ( .A(n51214), .Z(n51216) );
  NOR U71389 ( .A(n51216), .B(n51215), .Z(n56422) );
  IV U71390 ( .A(n51217), .Z(n51219) );
  XOR U71391 ( .A(n51218), .B(n51221), .Z(n56427) );
  NOR U71392 ( .A(n51219), .B(n56427), .Z(n52202) );
  IV U71393 ( .A(n51220), .Z(n51224) );
  NOR U71394 ( .A(n51222), .B(n51221), .Z(n51223) );
  IV U71395 ( .A(n51223), .Z(n51226) );
  NOR U71396 ( .A(n51224), .B(n51226), .Z(n57341) );
  IV U71397 ( .A(n51225), .Z(n51227) );
  NOR U71398 ( .A(n51227), .B(n51226), .Z(n57338) );
  IV U71399 ( .A(n51228), .Z(n51231) );
  NOR U71400 ( .A(n51229), .B(n52193), .Z(n51230) );
  IV U71401 ( .A(n51230), .Z(n52200) );
  NOR U71402 ( .A(n51231), .B(n52200), .Z(n56436) );
  IV U71403 ( .A(n51232), .Z(n51237) );
  IV U71404 ( .A(n51233), .Z(n52184) );
  NOR U71405 ( .A(n51234), .B(n52184), .Z(n51235) );
  IV U71406 ( .A(n51235), .Z(n51236) );
  NOR U71407 ( .A(n51237), .B(n51236), .Z(n56442) );
  IV U71408 ( .A(n51238), .Z(n51239) );
  NOR U71409 ( .A(n51239), .B(n51244), .Z(n57329) );
  IV U71410 ( .A(n51240), .Z(n51241) );
  NOR U71411 ( .A(n51241), .B(n51244), .Z(n57334) );
  NOR U71412 ( .A(n57329), .B(n57334), .Z(n52180) );
  IV U71413 ( .A(n51242), .Z(n51243) );
  NOR U71414 ( .A(n51244), .B(n51243), .Z(n57326) );
  IV U71415 ( .A(n51245), .Z(n51247) );
  NOR U71416 ( .A(n51247), .B(n51246), .Z(n56451) );
  IV U71417 ( .A(n51248), .Z(n51250) );
  NOR U71418 ( .A(n51250), .B(n51249), .Z(n57323) );
  NOR U71419 ( .A(n56451), .B(n57323), .Z(n52179) );
  NOR U71420 ( .A(n56462), .B(n51251), .Z(n51252) );
  IV U71421 ( .A(n51252), .Z(n51254) );
  IV U71422 ( .A(n51253), .Z(n52149) );
  XOR U71423 ( .A(n52147), .B(n52149), .Z(n56459) );
  NOR U71424 ( .A(n51254), .B(n56459), .Z(n52157) );
  IV U71425 ( .A(n51255), .Z(n51256) );
  NOR U71426 ( .A(n51256), .B(n52149), .Z(n56470) );
  IV U71427 ( .A(n51257), .Z(n51258) );
  NOR U71428 ( .A(n52150), .B(n51258), .Z(n56473) );
  IV U71429 ( .A(n51259), .Z(n51264) );
  IV U71430 ( .A(n51260), .Z(n51261) );
  NOR U71431 ( .A(n51262), .B(n51261), .Z(n51263) );
  IV U71432 ( .A(n51263), .Z(n51266) );
  NOR U71433 ( .A(n51264), .B(n51266), .Z(n57315) );
  IV U71434 ( .A(n51265), .Z(n51267) );
  NOR U71435 ( .A(n51267), .B(n51266), .Z(n57312) );
  IV U71436 ( .A(n51268), .Z(n51272) );
  NOR U71437 ( .A(n51270), .B(n51269), .Z(n51271) );
  IV U71438 ( .A(n51271), .Z(n51274) );
  NOR U71439 ( .A(n51272), .B(n51274), .Z(n56498) );
  IV U71440 ( .A(n51273), .Z(n51275) );
  NOR U71441 ( .A(n51275), .B(n51274), .Z(n56496) );
  IV U71442 ( .A(n51276), .Z(n51277) );
  NOR U71443 ( .A(n51277), .B(n51284), .Z(n51278) );
  IV U71444 ( .A(n51278), .Z(n51279) );
  NOR U71445 ( .A(n51283), .B(n51279), .Z(n56501) );
  NOR U71446 ( .A(n56496), .B(n56501), .Z(n51280) );
  IV U71447 ( .A(n51280), .Z(n52137) );
  IV U71448 ( .A(n51281), .Z(n51282) );
  NOR U71449 ( .A(n51284), .B(n51282), .Z(n56508) );
  IV U71450 ( .A(n51283), .Z(n51288) );
  NOR U71451 ( .A(n51285), .B(n51284), .Z(n51286) );
  IV U71452 ( .A(n51286), .Z(n51287) );
  NOR U71453 ( .A(n51288), .B(n51287), .Z(n56505) );
  NOR U71454 ( .A(n56508), .B(n56505), .Z(n52136) );
  IV U71455 ( .A(n51289), .Z(n51290) );
  NOR U71456 ( .A(n51291), .B(n51290), .Z(n57304) );
  IV U71457 ( .A(n51292), .Z(n51293) );
  NOR U71458 ( .A(n51294), .B(n51293), .Z(n56512) );
  NOR U71459 ( .A(n57304), .B(n56512), .Z(n52129) );
  IV U71460 ( .A(n51295), .Z(n51297) );
  NOR U71461 ( .A(n51297), .B(n51296), .Z(n56517) );
  IV U71462 ( .A(n51298), .Z(n51301) );
  NOR U71463 ( .A(n51299), .B(n56537), .Z(n51300) );
  IV U71464 ( .A(n51300), .Z(n51303) );
  NOR U71465 ( .A(n51301), .B(n51303), .Z(n56524) );
  IV U71466 ( .A(n51302), .Z(n51304) );
  NOR U71467 ( .A(n51304), .B(n51303), .Z(n56521) );
  IV U71468 ( .A(n51305), .Z(n51306) );
  NOR U71469 ( .A(n51306), .B(n56537), .Z(n56531) );
  IV U71470 ( .A(n51307), .Z(n51311) );
  NOR U71471 ( .A(n51309), .B(n51308), .Z(n51310) );
  IV U71472 ( .A(n51310), .Z(n51313) );
  NOR U71473 ( .A(n51311), .B(n51313), .Z(n56545) );
  IV U71474 ( .A(n51312), .Z(n51314) );
  NOR U71475 ( .A(n51314), .B(n51313), .Z(n56548) );
  IV U71476 ( .A(n51315), .Z(n51316) );
  NOR U71477 ( .A(n51317), .B(n51316), .Z(n51318) );
  IV U71478 ( .A(n51318), .Z(n51327) );
  NOR U71479 ( .A(n51320), .B(n51319), .Z(n51325) );
  NOR U71480 ( .A(n51322), .B(n51321), .Z(n51323) );
  IV U71481 ( .A(n51323), .Z(n51324) );
  NOR U71482 ( .A(n51325), .B(n51324), .Z(n51326) );
  IV U71483 ( .A(n51326), .Z(n51329) );
  NOR U71484 ( .A(n51327), .B(n51329), .Z(n56550) );
  NOR U71485 ( .A(n56548), .B(n56550), .Z(n52126) );
  IV U71486 ( .A(n51328), .Z(n51330) );
  NOR U71487 ( .A(n51330), .B(n51329), .Z(n56556) );
  IV U71488 ( .A(n51331), .Z(n51334) );
  NOR U71489 ( .A(n51332), .B(n51337), .Z(n51333) );
  IV U71490 ( .A(n51333), .Z(n52124) );
  NOR U71491 ( .A(n51334), .B(n52124), .Z(n56553) );
  IV U71492 ( .A(n51335), .Z(n51336) );
  NOR U71493 ( .A(n51337), .B(n51336), .Z(n56562) );
  IV U71494 ( .A(n51338), .Z(n51339) );
  NOR U71495 ( .A(n52119), .B(n51339), .Z(n56566) );
  NOR U71496 ( .A(n56562), .B(n56566), .Z(n52122) );
  IV U71497 ( .A(n51340), .Z(n51341) );
  NOR U71498 ( .A(n52110), .B(n51341), .Z(n57282) );
  IV U71499 ( .A(n51342), .Z(n51343) );
  NOR U71500 ( .A(n51344), .B(n51343), .Z(n56576) );
  IV U71501 ( .A(n51345), .Z(n51347) );
  NOR U71502 ( .A(n51347), .B(n51346), .Z(n56581) );
  NOR U71503 ( .A(n56576), .B(n56581), .Z(n51348) );
  IV U71504 ( .A(n51348), .Z(n52108) );
  IV U71505 ( .A(n51349), .Z(n57275) );
  IV U71506 ( .A(n51350), .Z(n51351) );
  NOR U71507 ( .A(n51351), .B(n52071), .Z(n56615) );
  IV U71508 ( .A(n51352), .Z(n51354) );
  NOR U71509 ( .A(n51354), .B(n51353), .Z(n51355) );
  IV U71510 ( .A(n51355), .Z(n56626) );
  IV U71511 ( .A(n51356), .Z(n51357) );
  NOR U71512 ( .A(n51358), .B(n51357), .Z(n51359) );
  IV U71513 ( .A(n51359), .Z(n52075) );
  IV U71514 ( .A(n51360), .Z(n52056) );
  IV U71515 ( .A(n51361), .Z(n51363) );
  NOR U71516 ( .A(n51363), .B(n51362), .Z(n51364) );
  IV U71517 ( .A(n51364), .Z(n57261) );
  NOR U71518 ( .A(n51365), .B(n51370), .Z(n51366) );
  IV U71519 ( .A(n51366), .Z(n56641) );
  NOR U71520 ( .A(n51367), .B(n56641), .Z(n52055) );
  IV U71521 ( .A(n51368), .Z(n51369) );
  NOR U71522 ( .A(n51370), .B(n51369), .Z(n56644) );
  IV U71523 ( .A(n51371), .Z(n51374) );
  IV U71524 ( .A(n51372), .Z(n51373) );
  NOR U71525 ( .A(n51374), .B(n51373), .Z(n56650) );
  IV U71526 ( .A(n51375), .Z(n51376) );
  NOR U71527 ( .A(n51376), .B(n51378), .Z(n57250) );
  IV U71528 ( .A(n51377), .Z(n51379) );
  NOR U71529 ( .A(n51379), .B(n51378), .Z(n57247) );
  IV U71530 ( .A(n51380), .Z(n51383) );
  NOR U71531 ( .A(n51381), .B(n52049), .Z(n51382) );
  IV U71532 ( .A(n51382), .Z(n52053) );
  NOR U71533 ( .A(n51383), .B(n52053), .Z(n57243) );
  IV U71534 ( .A(n51384), .Z(n51385) );
  NOR U71535 ( .A(n51386), .B(n51385), .Z(n57234) );
  NOR U71536 ( .A(n51387), .B(n52042), .Z(n57231) );
  IV U71537 ( .A(n51388), .Z(n51389) );
  NOR U71538 ( .A(n52042), .B(n51389), .Z(n57224) );
  IV U71539 ( .A(n51390), .Z(n51391) );
  NOR U71540 ( .A(n51391), .B(n51399), .Z(n51392) );
  IV U71541 ( .A(n51392), .Z(n51393) );
  NOR U71542 ( .A(n51394), .B(n51393), .Z(n56657) );
  IV U71543 ( .A(n51395), .Z(n51397) );
  NOR U71544 ( .A(n51397), .B(n51396), .Z(n51398) );
  IV U71545 ( .A(n51398), .Z(n51400) );
  NOR U71546 ( .A(n51400), .B(n51399), .Z(n56659) );
  NOR U71547 ( .A(n56657), .B(n56659), .Z(n52039) );
  IV U71548 ( .A(n51401), .Z(n51402) );
  NOR U71549 ( .A(n51402), .B(n56664), .Z(n52038) );
  IV U71550 ( .A(n51403), .Z(n51404) );
  NOR U71551 ( .A(n51404), .B(n56664), .Z(n57214) );
  IV U71552 ( .A(n51405), .Z(n51409) );
  NOR U71553 ( .A(n51407), .B(n51406), .Z(n51408) );
  IV U71554 ( .A(n51408), .Z(n52008) );
  NOR U71555 ( .A(n51409), .B(n52008), .Z(n57206) );
  NOR U71556 ( .A(n51411), .B(n51410), .Z(n56687) );
  NOR U71557 ( .A(n51413), .B(n51412), .Z(n56695) );
  IV U71558 ( .A(n51414), .Z(n51415) );
  NOR U71559 ( .A(n51415), .B(n51420), .Z(n51416) );
  IV U71560 ( .A(n51416), .Z(n51417) );
  NOR U71561 ( .A(n51419), .B(n51417), .Z(n57192) );
  NOR U71562 ( .A(n56695), .B(n57192), .Z(n51996) );
  IV U71563 ( .A(n51421), .Z(n51418) );
  NOR U71564 ( .A(n51418), .B(n51420), .Z(n57185) );
  IV U71565 ( .A(n51419), .Z(n51426) );
  XOR U71566 ( .A(n51421), .B(n51420), .Z(n51422) );
  NOR U71567 ( .A(n51423), .B(n51422), .Z(n51424) );
  IV U71568 ( .A(n51424), .Z(n51425) );
  NOR U71569 ( .A(n51426), .B(n51425), .Z(n57196) );
  NOR U71570 ( .A(n57185), .B(n57196), .Z(n51995) );
  IV U71571 ( .A(n51427), .Z(n51428) );
  NOR U71572 ( .A(n57182), .B(n51428), .Z(n51432) );
  IV U71573 ( .A(n51429), .Z(n51430) );
  NOR U71574 ( .A(n51431), .B(n51430), .Z(n57187) );
  NOR U71575 ( .A(n51432), .B(n57187), .Z(n51994) );
  IV U71576 ( .A(n51433), .Z(n51435) );
  NOR U71577 ( .A(n51435), .B(n51434), .Z(n62204) );
  NOR U71578 ( .A(n51437), .B(n51436), .Z(n61691) );
  NOR U71579 ( .A(n62204), .B(n61691), .Z(n56701) );
  IV U71580 ( .A(n51438), .Z(n51439) );
  NOR U71581 ( .A(n56711), .B(n51439), .Z(n51443) );
  IV U71582 ( .A(n51440), .Z(n51442) );
  NOR U71583 ( .A(n51442), .B(n51441), .Z(n56702) );
  NOR U71584 ( .A(n51443), .B(n56702), .Z(n51993) );
  IV U71585 ( .A(n51444), .Z(n51445) );
  NOR U71586 ( .A(n51446), .B(n51445), .Z(n51447) );
  IV U71587 ( .A(n51447), .Z(n56714) );
  IV U71588 ( .A(n51448), .Z(n51452) );
  NOR U71589 ( .A(n51450), .B(n51449), .Z(n51451) );
  IV U71590 ( .A(n51451), .Z(n51454) );
  NOR U71591 ( .A(n51452), .B(n51454), .Z(n56723) );
  IV U71592 ( .A(n51453), .Z(n51455) );
  NOR U71593 ( .A(n51455), .B(n51454), .Z(n51456) );
  IV U71594 ( .A(n51456), .Z(n56731) );
  IV U71595 ( .A(n51457), .Z(n51458) );
  NOR U71596 ( .A(n51458), .B(n51972), .Z(n51979) );
  IV U71597 ( .A(n51979), .Z(n51971) );
  IV U71598 ( .A(n51976), .Z(n51462) );
  NOR U71599 ( .A(n51459), .B(n51972), .Z(n51460) );
  IV U71600 ( .A(n51460), .Z(n51461) );
  NOR U71601 ( .A(n51462), .B(n51461), .Z(n57160) );
  IV U71602 ( .A(n51463), .Z(n51467) );
  IV U71603 ( .A(n51464), .Z(n56739) );
  NOR U71604 ( .A(n56739), .B(n51465), .Z(n51466) );
  IV U71605 ( .A(n51466), .Z(n51469) );
  NOR U71606 ( .A(n51467), .B(n51469), .Z(n57157) );
  IV U71607 ( .A(n51468), .Z(n51470) );
  NOR U71608 ( .A(n51470), .B(n51469), .Z(n56734) );
  IV U71609 ( .A(n51471), .Z(n51472) );
  NOR U71610 ( .A(n51472), .B(n56739), .Z(n51969) );
  NOR U71611 ( .A(n57146), .B(n57151), .Z(n51473) );
  NOR U71612 ( .A(n57148), .B(n51473), .Z(n51968) );
  IV U71613 ( .A(n51474), .Z(n56751) );
  XOR U71614 ( .A(n51961), .B(n56751), .Z(n51964) );
  NOR U71615 ( .A(n56745), .B(n56750), .Z(n51475) );
  NOR U71616 ( .A(n51964), .B(n51475), .Z(n51967) );
  IV U71617 ( .A(n51476), .Z(n51477) );
  NOR U71618 ( .A(n51477), .B(n51479), .Z(n56761) );
  IV U71619 ( .A(n51478), .Z(n51480) );
  NOR U71620 ( .A(n51480), .B(n51479), .Z(n57130) );
  NOR U71621 ( .A(n56761), .B(n57130), .Z(n51958) );
  IV U71622 ( .A(n51481), .Z(n51483) );
  NOR U71623 ( .A(n51483), .B(n51482), .Z(n57128) );
  IV U71624 ( .A(n51484), .Z(n51943) );
  IV U71625 ( .A(n51485), .Z(n51486) );
  NOR U71626 ( .A(n51943), .B(n51486), .Z(n57121) );
  IV U71627 ( .A(n51487), .Z(n51488) );
  NOR U71628 ( .A(n51488), .B(n51490), .Z(n57110) );
  NOR U71629 ( .A(n57121), .B(n57110), .Z(n51937) );
  IV U71630 ( .A(n51489), .Z(n51491) );
  NOR U71631 ( .A(n51491), .B(n51490), .Z(n56772) );
  IV U71632 ( .A(n51492), .Z(n51495) );
  NOR U71633 ( .A(n51493), .B(n51500), .Z(n51494) );
  IV U71634 ( .A(n51494), .Z(n51497) );
  NOR U71635 ( .A(n51495), .B(n51497), .Z(n57112) );
  IV U71636 ( .A(n51496), .Z(n51498) );
  NOR U71637 ( .A(n51498), .B(n51497), .Z(n56776) );
  IV U71638 ( .A(n51499), .Z(n51503) );
  NOR U71639 ( .A(n51501), .B(n51500), .Z(n51502) );
  IV U71640 ( .A(n51502), .Z(n51509) );
  NOR U71641 ( .A(n51503), .B(n51509), .Z(n57103) );
  NOR U71642 ( .A(n56776), .B(n57103), .Z(n51504) );
  IV U71643 ( .A(n51504), .Z(n51936) );
  IV U71644 ( .A(n51505), .Z(n51507) );
  NOR U71645 ( .A(n51507), .B(n51506), .Z(n56778) );
  IV U71646 ( .A(n51508), .Z(n51510) );
  NOR U71647 ( .A(n51510), .B(n51509), .Z(n57106) );
  NOR U71648 ( .A(n56778), .B(n57106), .Z(n51935) );
  IV U71649 ( .A(n51511), .Z(n51512) );
  NOR U71650 ( .A(n51919), .B(n51512), .Z(n51926) );
  IV U71651 ( .A(n51926), .Z(n51916) );
  IV U71652 ( .A(n51513), .Z(n51514) );
  NOR U71653 ( .A(n51514), .B(n51922), .Z(n57098) );
  NOR U71654 ( .A(n51922), .B(n51515), .Z(n57095) );
  IV U71655 ( .A(n51516), .Z(n51518) );
  IV U71656 ( .A(n51517), .Z(n51905) );
  NOR U71657 ( .A(n51518), .B(n51905), .Z(n56787) );
  IV U71658 ( .A(n51519), .Z(n51520) );
  NOR U71659 ( .A(n51520), .B(n51896), .Z(n56797) );
  IV U71660 ( .A(n51521), .Z(n51523) );
  NOR U71661 ( .A(n51523), .B(n51522), .Z(n51524) );
  IV U71662 ( .A(n51524), .Z(n56809) );
  IV U71663 ( .A(n51525), .Z(n51885) );
  NOR U71664 ( .A(n51885), .B(n51526), .Z(n56806) );
  IV U71665 ( .A(n51527), .Z(n51531) );
  NOR U71666 ( .A(n51529), .B(n51528), .Z(n51530) );
  IV U71667 ( .A(n51530), .Z(n51533) );
  NOR U71668 ( .A(n51531), .B(n51533), .Z(n67310) );
  NOR U71669 ( .A(n56806), .B(n67310), .Z(n51883) );
  IV U71670 ( .A(n51532), .Z(n51534) );
  NOR U71671 ( .A(n51534), .B(n51533), .Z(n56810) );
  IV U71672 ( .A(n51535), .Z(n51536) );
  NOR U71673 ( .A(n51537), .B(n51536), .Z(n56814) );
  IV U71674 ( .A(n51538), .Z(n51541) );
  IV U71675 ( .A(n51539), .Z(n51540) );
  NOR U71676 ( .A(n51541), .B(n51540), .Z(n56815) );
  NOR U71677 ( .A(n56814), .B(n56815), .Z(n51882) );
  NOR U71678 ( .A(n51542), .B(n51541), .Z(n56822) );
  NOR U71679 ( .A(n57079), .B(n56822), .Z(n51881) );
  IV U71680 ( .A(n51543), .Z(n51546) );
  IV U71681 ( .A(n51544), .Z(n51545) );
  NOR U71682 ( .A(n51546), .B(n51545), .Z(n62068) );
  NOR U71683 ( .A(n61786), .B(n62068), .Z(n57076) );
  IV U71684 ( .A(n51547), .Z(n51549) );
  NOR U71685 ( .A(n51549), .B(n51548), .Z(n51879) );
  IV U71686 ( .A(n51879), .Z(n51869) );
  IV U71687 ( .A(n51550), .Z(n51552) );
  NOR U71688 ( .A(n51552), .B(n51551), .Z(n51866) );
  IV U71689 ( .A(n51866), .Z(n51856) );
  IV U71690 ( .A(n51553), .Z(n51854) );
  IV U71691 ( .A(n51554), .Z(n51555) );
  NOR U71692 ( .A(n51854), .B(n51555), .Z(n56824) );
  NOR U71693 ( .A(n51557), .B(n51556), .Z(n51558) );
  IV U71694 ( .A(n51558), .Z(n51559) );
  NOR U71695 ( .A(n51560), .B(n51559), .Z(n51847) );
  IV U71696 ( .A(n51561), .Z(n51562) );
  NOR U71697 ( .A(n51565), .B(n51562), .Z(n56836) );
  IV U71698 ( .A(n51566), .Z(n51563) );
  NOR U71699 ( .A(n51563), .B(n51565), .Z(n57049) );
  IV U71700 ( .A(n51564), .Z(n51568) );
  XOR U71701 ( .A(n51566), .B(n51565), .Z(n51567) );
  NOR U71702 ( .A(n51568), .B(n51567), .Z(n56841) );
  NOR U71703 ( .A(n57049), .B(n56841), .Z(n51822) );
  IV U71704 ( .A(n51569), .Z(n51570) );
  NOR U71705 ( .A(n51571), .B(n51570), .Z(n51820) );
  IV U71706 ( .A(n51820), .Z(n51814) );
  IV U71707 ( .A(n51572), .Z(n51573) );
  NOR U71708 ( .A(n51574), .B(n51573), .Z(n57043) );
  IV U71709 ( .A(n51575), .Z(n51585) );
  NOR U71710 ( .A(n51577), .B(n51576), .Z(n51583) );
  IV U71711 ( .A(n51578), .Z(n51810) );
  XOR U71712 ( .A(n51810), .B(n51809), .Z(n51579) );
  NOR U71713 ( .A(n51580), .B(n51579), .Z(n51581) );
  IV U71714 ( .A(n51581), .Z(n51582) );
  NOR U71715 ( .A(n51583), .B(n51582), .Z(n51584) );
  IV U71716 ( .A(n51584), .Z(n51587) );
  NOR U71717 ( .A(n51585), .B(n51587), .Z(n57039) );
  IV U71718 ( .A(n51586), .Z(n51588) );
  NOR U71719 ( .A(n51588), .B(n51587), .Z(n57036) );
  IV U71720 ( .A(n51589), .Z(n51592) );
  NOR U71721 ( .A(n51590), .B(n51810), .Z(n51591) );
  IV U71722 ( .A(n51591), .Z(n51594) );
  NOR U71723 ( .A(n51592), .B(n51594), .Z(n57032) );
  IV U71724 ( .A(n51593), .Z(n51595) );
  NOR U71725 ( .A(n51595), .B(n51594), .Z(n51596) );
  IV U71726 ( .A(n51596), .Z(n57030) );
  NOR U71727 ( .A(n51598), .B(n51597), .Z(n57015) );
  IV U71728 ( .A(n51599), .Z(n51600) );
  NOR U71729 ( .A(n51600), .B(n51603), .Z(n61978) );
  IV U71730 ( .A(n51601), .Z(n51602) );
  NOR U71731 ( .A(n51603), .B(n51602), .Z(n61825) );
  NOR U71732 ( .A(n61978), .B(n61825), .Z(n57014) );
  IV U71733 ( .A(n51604), .Z(n51611) );
  IV U71734 ( .A(n51605), .Z(n51606) );
  NOR U71735 ( .A(n51611), .B(n51606), .Z(n61842) );
  IV U71736 ( .A(n51607), .Z(n51608) );
  NOR U71737 ( .A(n51608), .B(n51806), .Z(n61837) );
  NOR U71738 ( .A(n61842), .B(n61837), .Z(n56844) );
  IV U71739 ( .A(n51609), .Z(n51610) );
  NOR U71740 ( .A(n51611), .B(n51610), .Z(n56851) );
  IV U71741 ( .A(n51612), .Z(n51613) );
  NOR U71742 ( .A(n51785), .B(n51613), .Z(n56865) );
  IV U71743 ( .A(n51614), .Z(n51617) );
  NOR U71744 ( .A(n51615), .B(n51772), .Z(n51616) );
  IV U71745 ( .A(n51616), .Z(n51765) );
  NOR U71746 ( .A(n51617), .B(n51765), .Z(n57008) );
  NOR U71747 ( .A(n56865), .B(n57008), .Z(n51783) );
  IV U71748 ( .A(n51618), .Z(n51622) );
  NOR U71749 ( .A(n51620), .B(n51619), .Z(n51621) );
  IV U71750 ( .A(n51621), .Z(n51761) );
  NOR U71751 ( .A(n51622), .B(n51761), .Z(n57000) );
  IV U71752 ( .A(n51623), .Z(n51626) );
  NOR U71753 ( .A(n51624), .B(n51632), .Z(n51625) );
  IV U71754 ( .A(n51625), .Z(n51629) );
  NOR U71755 ( .A(n51626), .B(n51629), .Z(n56885) );
  IV U71756 ( .A(n51751), .Z(n51627) );
  XOR U71757 ( .A(n51631), .B(n51632), .Z(n51750) );
  NOR U71758 ( .A(n51627), .B(n51750), .Z(n56894) );
  IV U71759 ( .A(n51628), .Z(n51630) );
  NOR U71760 ( .A(n51630), .B(n51629), .Z(n56891) );
  NOR U71761 ( .A(n56894), .B(n56891), .Z(n51747) );
  IV U71762 ( .A(n51631), .Z(n51633) );
  NOR U71763 ( .A(n51633), .B(n51632), .Z(n56993) );
  IV U71764 ( .A(n51634), .Z(n51637) );
  IV U71765 ( .A(n51635), .Z(n51636) );
  NOR U71766 ( .A(n51637), .B(n51636), .Z(n61889) );
  NOR U71767 ( .A(n61947), .B(n61889), .Z(n56903) );
  IV U71768 ( .A(n51638), .Z(n51639) );
  NOR U71769 ( .A(n51639), .B(n51732), .Z(n51640) );
  IV U71770 ( .A(n51640), .Z(n51641) );
  NOR U71771 ( .A(n51735), .B(n51641), .Z(n56989) );
  IV U71772 ( .A(n51642), .Z(n51644) );
  NOR U71773 ( .A(n51644), .B(n51643), .Z(n56910) );
  IV U71774 ( .A(n51645), .Z(n51647) );
  NOR U71775 ( .A(n51647), .B(n51646), .Z(n56913) );
  IV U71776 ( .A(n51648), .Z(n51650) );
  IV U71777 ( .A(n51649), .Z(n51652) );
  NOR U71778 ( .A(n51650), .B(n51652), .Z(n56925) );
  IV U71779 ( .A(n56925), .Z(n56923) );
  IV U71780 ( .A(n51651), .Z(n51653) );
  NOR U71781 ( .A(n51653), .B(n51652), .Z(n51654) );
  IV U71782 ( .A(n51654), .Z(n56933) );
  IV U71783 ( .A(n51655), .Z(n51656) );
  NOR U71784 ( .A(n51656), .B(n51658), .Z(n56978) );
  IV U71785 ( .A(n56978), .Z(n56975) );
  IV U71786 ( .A(n51657), .Z(n51659) );
  NOR U71787 ( .A(n51659), .B(n51658), .Z(n56947) );
  IV U71788 ( .A(n51660), .Z(n51662) );
  NOR U71789 ( .A(n51662), .B(n51661), .Z(n56941) );
  NOR U71790 ( .A(n56947), .B(n56941), .Z(n51702) );
  IV U71791 ( .A(n51663), .Z(n51664) );
  NOR U71792 ( .A(n51665), .B(n51664), .Z(n56949) );
  IV U71793 ( .A(n51666), .Z(n51668) );
  NOR U71794 ( .A(n51668), .B(n51667), .Z(n56946) );
  NOR U71795 ( .A(n56949), .B(n56946), .Z(n51669) );
  IV U71796 ( .A(n51669), .Z(n51701) );
  IV U71797 ( .A(n51670), .Z(n51672) );
  IV U71798 ( .A(n51671), .Z(n51674) );
  NOR U71799 ( .A(n51672), .B(n51674), .Z(n56962) );
  IV U71800 ( .A(n51673), .Z(n51677) );
  NOR U71801 ( .A(n51675), .B(n51674), .Z(n51676) );
  IV U71802 ( .A(n51676), .Z(n51681) );
  NOR U71803 ( .A(n51677), .B(n51681), .Z(n51678) );
  NOR U71804 ( .A(n56962), .B(n51678), .Z(n51679) );
  IV U71805 ( .A(n51679), .Z(n56945) );
  IV U71806 ( .A(n51680), .Z(n51682) );
  NOR U71807 ( .A(n51682), .B(n51681), .Z(n51683) );
  NOR U71808 ( .A(n56963), .B(n51683), .Z(n51684) );
  IV U71809 ( .A(n51684), .Z(n51700) );
  IV U71810 ( .A(n51685), .Z(n51686) );
  NOR U71811 ( .A(n51687), .B(n51686), .Z(n51689) );
  NOR U71812 ( .A(n51689), .B(n51688), .Z(n51690) );
  IV U71813 ( .A(n51690), .Z(n51699) );
  NOR U71814 ( .A(n51692), .B(n51691), .Z(n51694) );
  NOR U71815 ( .A(n51694), .B(n51693), .Z(n51695) );
  NOR U71816 ( .A(n51696), .B(n51695), .Z(n51697) );
  IV U71817 ( .A(n51697), .Z(n51698) );
  NOR U71818 ( .A(n51699), .B(n51698), .Z(n56971) );
  XOR U71819 ( .A(n51700), .B(n56971), .Z(n56944) );
  XOR U71820 ( .A(n56945), .B(n56944), .Z(n56957) );
  XOR U71821 ( .A(n51701), .B(n56957), .Z(n56943) );
  XOR U71822 ( .A(n51702), .B(n56943), .Z(n56977) );
  XOR U71823 ( .A(n56975), .B(n56977), .Z(n56938) );
  IV U71824 ( .A(n51703), .Z(n51704) );
  NOR U71825 ( .A(n51715), .B(n51704), .Z(n56935) );
  IV U71826 ( .A(n51705), .Z(n51707) );
  NOR U71827 ( .A(n51707), .B(n51706), .Z(n56979) );
  IV U71828 ( .A(n51708), .Z(n51709) );
  NOR U71829 ( .A(n51710), .B(n51709), .Z(n56937) );
  NOR U71830 ( .A(n56979), .B(n56937), .Z(n51711) );
  IV U71831 ( .A(n51711), .Z(n51712) );
  NOR U71832 ( .A(n56935), .B(n51712), .Z(n51713) );
  XOR U71833 ( .A(n56938), .B(n51713), .Z(n51714) );
  IV U71834 ( .A(n51714), .Z(n56932) );
  NOR U71835 ( .A(n51716), .B(n51715), .Z(n51717) );
  IV U71836 ( .A(n51717), .Z(n51718) );
  NOR U71837 ( .A(n51719), .B(n51718), .Z(n56930) );
  XOR U71838 ( .A(n56932), .B(n56930), .Z(n56934) );
  XOR U71839 ( .A(n56933), .B(n56934), .Z(n56924) );
  XOR U71840 ( .A(n56923), .B(n56924), .Z(n56920) );
  IV U71841 ( .A(n51720), .Z(n51721) );
  NOR U71842 ( .A(n51722), .B(n51721), .Z(n56926) );
  IV U71843 ( .A(n51723), .Z(n51725) );
  NOR U71844 ( .A(n51725), .B(n51724), .Z(n56919) );
  NOR U71845 ( .A(n56926), .B(n56919), .Z(n51726) );
  XOR U71846 ( .A(n56920), .B(n51726), .Z(n51727) );
  IV U71847 ( .A(n51727), .Z(n56915) );
  XOR U71848 ( .A(n56913), .B(n56915), .Z(n56911) );
  XOR U71849 ( .A(n56910), .B(n56911), .Z(n56906) );
  IV U71850 ( .A(n51728), .Z(n51730) );
  NOR U71851 ( .A(n51730), .B(n51729), .Z(n56908) );
  IV U71852 ( .A(n51731), .Z(n51733) );
  NOR U71853 ( .A(n51733), .B(n51732), .Z(n56905) );
  NOR U71854 ( .A(n56908), .B(n56905), .Z(n51734) );
  XOR U71855 ( .A(n56906), .B(n51734), .Z(n56986) );
  IV U71856 ( .A(n51735), .Z(n51741) );
  IV U71857 ( .A(n51736), .Z(n51738) );
  NOR U71858 ( .A(n51738), .B(n51737), .Z(n51739) );
  IV U71859 ( .A(n51739), .Z(n51740) );
  NOR U71860 ( .A(n51741), .B(n51740), .Z(n51742) );
  IV U71861 ( .A(n51742), .Z(n56987) );
  XOR U71862 ( .A(n56986), .B(n56987), .Z(n56990) );
  XOR U71863 ( .A(n56989), .B(n56990), .Z(n56901) );
  XOR U71864 ( .A(n56900), .B(n56901), .Z(n61891) );
  XOR U71865 ( .A(n56903), .B(n61891), .Z(n56898) );
  IV U71866 ( .A(n51743), .Z(n51744) );
  NOR U71867 ( .A(n51745), .B(n51744), .Z(n56996) );
  NOR U71868 ( .A(n56897), .B(n56996), .Z(n51746) );
  XOR U71869 ( .A(n56898), .B(n51746), .Z(n56995) );
  XOR U71870 ( .A(n56993), .B(n56995), .Z(n56893) );
  XOR U71871 ( .A(n51747), .B(n56893), .Z(n51748) );
  IV U71872 ( .A(n51748), .Z(n56887) );
  XOR U71873 ( .A(n56885), .B(n56887), .Z(n56881) );
  IV U71874 ( .A(n51749), .Z(n51753) );
  XOR U71875 ( .A(n51751), .B(n51750), .Z(n51752) );
  NOR U71876 ( .A(n51753), .B(n51752), .Z(n51754) );
  IV U71877 ( .A(n51754), .Z(n56880) );
  NOR U71878 ( .A(n51755), .B(n56880), .Z(n51756) );
  XOR U71879 ( .A(n56881), .B(n51756), .Z(n57001) );
  XOR U71880 ( .A(n57000), .B(n57001), .Z(n57005) );
  IV U71881 ( .A(n51757), .Z(n51758) );
  NOR U71882 ( .A(n51759), .B(n51758), .Z(n56876) );
  IV U71883 ( .A(n51760), .Z(n51762) );
  NOR U71884 ( .A(n51762), .B(n51761), .Z(n57003) );
  NOR U71885 ( .A(n56876), .B(n57003), .Z(n51763) );
  XOR U71886 ( .A(n57005), .B(n51763), .Z(n51775) );
  IV U71887 ( .A(n51775), .Z(n56874) );
  IV U71888 ( .A(n51764), .Z(n51766) );
  NOR U71889 ( .A(n51766), .B(n51765), .Z(n51781) );
  IV U71890 ( .A(n51781), .Z(n51767) );
  NOR U71891 ( .A(n56874), .B(n51767), .Z(n61864) );
  IV U71892 ( .A(n51768), .Z(n51770) );
  NOR U71893 ( .A(n51770), .B(n51769), .Z(n56870) );
  IV U71894 ( .A(n51771), .Z(n51773) );
  NOR U71895 ( .A(n51773), .B(n51772), .Z(n56872) );
  NOR U71896 ( .A(n56870), .B(n56872), .Z(n51774) );
  XOR U71897 ( .A(n51775), .B(n51774), .Z(n56868) );
  IV U71898 ( .A(n51776), .Z(n51778) );
  NOR U71899 ( .A(n51778), .B(n51777), .Z(n51779) );
  IV U71900 ( .A(n51779), .Z(n56869) );
  XOR U71901 ( .A(n56868), .B(n56869), .Z(n51780) );
  NOR U71902 ( .A(n51781), .B(n51780), .Z(n51782) );
  NOR U71903 ( .A(n61864), .B(n51782), .Z(n56866) );
  XOR U71904 ( .A(n51783), .B(n56866), .Z(n56864) );
  IV U71905 ( .A(n51784), .Z(n51786) );
  NOR U71906 ( .A(n51786), .B(n51785), .Z(n56862) );
  XOR U71907 ( .A(n56864), .B(n56862), .Z(n56861) );
  IV U71908 ( .A(n51787), .Z(n51792) );
  IV U71909 ( .A(n51788), .Z(n51789) );
  NOR U71910 ( .A(n51790), .B(n51789), .Z(n51791) );
  IV U71911 ( .A(n51791), .Z(n51796) );
  NOR U71912 ( .A(n51792), .B(n51796), .Z(n56859) );
  XOR U71913 ( .A(n56861), .B(n56859), .Z(n56856) );
  IV U71914 ( .A(n51793), .Z(n51794) );
  NOR U71915 ( .A(n51794), .B(n51801), .Z(n56854) );
  IV U71916 ( .A(n51795), .Z(n51797) );
  NOR U71917 ( .A(n51797), .B(n51796), .Z(n56857) );
  NOR U71918 ( .A(n56854), .B(n56857), .Z(n51798) );
  XOR U71919 ( .A(n56856), .B(n51798), .Z(n51799) );
  IV U71920 ( .A(n51799), .Z(n56850) );
  IV U71921 ( .A(n51800), .Z(n51802) );
  NOR U71922 ( .A(n51802), .B(n51801), .Z(n56848) );
  XOR U71923 ( .A(n56850), .B(n56848), .Z(n56853) );
  XOR U71924 ( .A(n56851), .B(n56853), .Z(n61838) );
  XOR U71925 ( .A(n56844), .B(n61838), .Z(n56845) );
  NOR U71926 ( .A(n51804), .B(n51803), .Z(n61975) );
  IV U71927 ( .A(n51805), .Z(n51807) );
  NOR U71928 ( .A(n51807), .B(n51806), .Z(n61832) );
  NOR U71929 ( .A(n61975), .B(n61832), .Z(n56846) );
  XOR U71930 ( .A(n56845), .B(n56846), .Z(n61828) );
  XOR U71931 ( .A(n57014), .B(n61828), .Z(n51808) );
  IV U71932 ( .A(n51808), .Z(n57016) );
  XOR U71933 ( .A(n57015), .B(n57016), .Z(n57021) );
  IV U71934 ( .A(n51809), .Z(n57024) );
  NOR U71935 ( .A(n51810), .B(n57024), .Z(n51811) );
  NOR U71936 ( .A(n57022), .B(n51811), .Z(n51812) );
  XOR U71937 ( .A(n57021), .B(n51812), .Z(n57029) );
  XOR U71938 ( .A(n57030), .B(n57029), .Z(n57033) );
  XOR U71939 ( .A(n57032), .B(n57033), .Z(n57037) );
  XOR U71940 ( .A(n57036), .B(n57037), .Z(n57040) );
  XOR U71941 ( .A(n57039), .B(n57040), .Z(n57046) );
  XOR U71942 ( .A(n57043), .B(n57046), .Z(n51813) );
  NOR U71943 ( .A(n51814), .B(n51813), .Z(n67357) );
  IV U71944 ( .A(n51815), .Z(n51816) );
  NOR U71945 ( .A(n51817), .B(n51816), .Z(n57045) );
  NOR U71946 ( .A(n57045), .B(n57043), .Z(n51818) );
  XOR U71947 ( .A(n57046), .B(n51818), .Z(n51819) );
  NOR U71948 ( .A(n51820), .B(n51819), .Z(n51821) );
  NOR U71949 ( .A(n67357), .B(n51821), .Z(n56842) );
  XOR U71950 ( .A(n51822), .B(n56842), .Z(n56839) );
  XOR U71951 ( .A(n56836), .B(n56839), .Z(n56834) );
  IV U71952 ( .A(n51823), .Z(n51824) );
  NOR U71953 ( .A(n51825), .B(n51824), .Z(n56838) );
  IV U71954 ( .A(n51835), .Z(n51829) );
  NOR U71955 ( .A(n51826), .B(n51838), .Z(n51827) );
  IV U71956 ( .A(n51827), .Z(n51828) );
  NOR U71957 ( .A(n51829), .B(n51828), .Z(n56832) );
  NOR U71958 ( .A(n56838), .B(n56832), .Z(n51830) );
  XOR U71959 ( .A(n56834), .B(n51830), .Z(n57053) );
  IV U71960 ( .A(n51831), .Z(n51832) );
  NOR U71961 ( .A(n51832), .B(n51838), .Z(n51833) );
  IV U71962 ( .A(n51833), .Z(n51834) );
  NOR U71963 ( .A(n51835), .B(n51834), .Z(n51836) );
  IV U71964 ( .A(n51836), .Z(n57054) );
  XOR U71965 ( .A(n57053), .B(n57054), .Z(n57058) );
  IV U71966 ( .A(n51837), .Z(n51841) );
  NOR U71967 ( .A(n51839), .B(n51838), .Z(n51840) );
  IV U71968 ( .A(n51840), .Z(n51843) );
  NOR U71969 ( .A(n51841), .B(n51843), .Z(n56830) );
  IV U71970 ( .A(n51842), .Z(n51844) );
  NOR U71971 ( .A(n51844), .B(n51843), .Z(n57056) );
  NOR U71972 ( .A(n56830), .B(n57056), .Z(n51845) );
  XOR U71973 ( .A(n57058), .B(n51845), .Z(n51846) );
  NOR U71974 ( .A(n51847), .B(n51846), .Z(n51850) );
  IV U71975 ( .A(n51847), .Z(n51849) );
  XOR U71976 ( .A(n57056), .B(n57058), .Z(n51848) );
  NOR U71977 ( .A(n51849), .B(n51848), .Z(n62031) );
  NOR U71978 ( .A(n51850), .B(n62031), .Z(n56827) );
  IV U71979 ( .A(n51853), .Z(n51851) );
  NOR U71980 ( .A(n51854), .B(n51851), .Z(n62025) );
  IV U71981 ( .A(n51852), .Z(n51855) );
  XOR U71982 ( .A(n51854), .B(n51853), .Z(n51860) );
  NOR U71983 ( .A(n51855), .B(n51860), .Z(n61800) );
  NOR U71984 ( .A(n62025), .B(n61800), .Z(n56828) );
  XOR U71985 ( .A(n56827), .B(n56828), .Z(n56825) );
  XOR U71986 ( .A(n56824), .B(n56825), .Z(n57064) );
  NOR U71987 ( .A(n51856), .B(n57064), .Z(n61796) );
  IV U71988 ( .A(n51857), .Z(n51858) );
  NOR U71989 ( .A(n51859), .B(n51858), .Z(n57067) );
  NOR U71990 ( .A(n51861), .B(n51860), .Z(n51862) );
  IV U71991 ( .A(n51862), .Z(n57063) );
  NOR U71992 ( .A(n51863), .B(n57063), .Z(n51864) );
  XOR U71993 ( .A(n57064), .B(n51864), .Z(n57068) );
  XOR U71994 ( .A(n57067), .B(n57068), .Z(n51873) );
  IV U71995 ( .A(n51873), .Z(n51865) );
  NOR U71996 ( .A(n51866), .B(n51865), .Z(n51867) );
  NOR U71997 ( .A(n61796), .B(n51867), .Z(n51875) );
  IV U71998 ( .A(n51875), .Z(n51868) );
  NOR U71999 ( .A(n51869), .B(n51868), .Z(n61793) );
  IV U72000 ( .A(n51870), .Z(n51872) );
  NOR U72001 ( .A(n51872), .B(n51871), .Z(n51876) );
  IV U72002 ( .A(n51876), .Z(n51874) );
  NOR U72003 ( .A(n51874), .B(n51873), .Z(n61790) );
  NOR U72004 ( .A(n51876), .B(n51875), .Z(n51877) );
  NOR U72005 ( .A(n61790), .B(n51877), .Z(n51878) );
  NOR U72006 ( .A(n51879), .B(n51878), .Z(n51880) );
  NOR U72007 ( .A(n61793), .B(n51880), .Z(n57075) );
  XOR U72008 ( .A(n57076), .B(n57075), .Z(n57080) );
  XOR U72009 ( .A(n51881), .B(n57080), .Z(n56819) );
  XOR U72010 ( .A(n51882), .B(n56819), .Z(n56812) );
  XOR U72011 ( .A(n56810), .B(n56812), .Z(n67309) );
  XOR U72012 ( .A(n51883), .B(n67309), .Z(n56807) );
  XOR U72013 ( .A(n56809), .B(n56807), .Z(n56802) );
  IV U72014 ( .A(n51893), .Z(n51888) );
  NOR U72015 ( .A(n51885), .B(n51884), .Z(n51886) );
  IV U72016 ( .A(n51886), .Z(n51887) );
  NOR U72017 ( .A(n51888), .B(n51887), .Z(n56800) );
  XOR U72018 ( .A(n56802), .B(n56800), .Z(n56805) );
  IV U72019 ( .A(n51889), .Z(n51890) );
  NOR U72020 ( .A(n51890), .B(n51896), .Z(n51891) );
  IV U72021 ( .A(n51891), .Z(n51892) );
  NOR U72022 ( .A(n51893), .B(n51892), .Z(n56803) );
  XOR U72023 ( .A(n56805), .B(n56803), .Z(n56798) );
  XOR U72024 ( .A(n56797), .B(n56798), .Z(n56795) );
  IV U72025 ( .A(n51894), .Z(n51895) );
  NOR U72026 ( .A(n51896), .B(n51895), .Z(n56793) );
  XOR U72027 ( .A(n56795), .B(n56793), .Z(n61766) );
  IV U72028 ( .A(n51897), .Z(n51898) );
  NOR U72029 ( .A(n51899), .B(n51898), .Z(n61767) );
  NOR U72030 ( .A(n61767), .B(n57086), .Z(n51900) );
  XOR U72031 ( .A(n61766), .B(n51900), .Z(n57088) );
  IV U72032 ( .A(n51901), .Z(n51903) );
  NOR U72033 ( .A(n51903), .B(n51902), .Z(n57087) );
  IV U72034 ( .A(n51904), .Z(n51906) );
  NOR U72035 ( .A(n51906), .B(n51905), .Z(n57091) );
  NOR U72036 ( .A(n57087), .B(n57091), .Z(n51907) );
  XOR U72037 ( .A(n57088), .B(n51907), .Z(n56789) );
  XOR U72038 ( .A(n56787), .B(n56789), .Z(n56791) );
  IV U72039 ( .A(n51908), .Z(n51910) );
  NOR U72040 ( .A(n51910), .B(n51909), .Z(n56790) );
  IV U72041 ( .A(n51911), .Z(n51912) );
  NOR U72042 ( .A(n51913), .B(n51912), .Z(n56784) );
  NOR U72043 ( .A(n56790), .B(n56784), .Z(n51914) );
  XOR U72044 ( .A(n56791), .B(n51914), .Z(n51915) );
  IV U72045 ( .A(n51915), .Z(n57096) );
  XOR U72046 ( .A(n57095), .B(n57096), .Z(n57100) );
  XOR U72047 ( .A(n57098), .B(n57100), .Z(n56781) );
  NOR U72048 ( .A(n51916), .B(n56781), .Z(n57102) );
  IV U72049 ( .A(n57102), .Z(n61754) );
  NOR U72050 ( .A(n61754), .B(n51917), .Z(n51934) );
  IV U72051 ( .A(n51917), .Z(n51918) );
  NOR U72052 ( .A(n51919), .B(n51918), .Z(n51927) );
  IV U72053 ( .A(n51927), .Z(n51925) );
  IV U72054 ( .A(n51920), .Z(n51921) );
  NOR U72055 ( .A(n51922), .B(n51921), .Z(n51923) );
  IV U72056 ( .A(n51923), .Z(n56782) );
  XOR U72057 ( .A(n56782), .B(n56781), .Z(n51930) );
  IV U72058 ( .A(n51930), .Z(n51924) );
  NOR U72059 ( .A(n51925), .B(n51924), .Z(n67270) );
  NOR U72060 ( .A(n51927), .B(n51926), .Z(n51928) );
  IV U72061 ( .A(n51928), .Z(n51929) );
  NOR U72062 ( .A(n51930), .B(n51929), .Z(n51931) );
  NOR U72063 ( .A(n67270), .B(n51931), .Z(n51932) );
  IV U72064 ( .A(n51932), .Z(n51933) );
  NOR U72065 ( .A(n51934), .B(n51933), .Z(n56779) );
  XOR U72066 ( .A(n51935), .B(n56779), .Z(n57105) );
  XOR U72067 ( .A(n51936), .B(n57105), .Z(n57113) );
  XOR U72068 ( .A(n57112), .B(n57113), .Z(n56774) );
  XOR U72069 ( .A(n56772), .B(n56774), .Z(n57122) );
  XOR U72070 ( .A(n51937), .B(n57122), .Z(n51938) );
  IV U72071 ( .A(n51938), .Z(n56768) );
  IV U72072 ( .A(n51939), .Z(n51940) );
  NOR U72073 ( .A(n51943), .B(n51940), .Z(n56766) );
  XOR U72074 ( .A(n56768), .B(n56766), .Z(n56771) );
  IV U72075 ( .A(n51941), .Z(n51948) );
  NOR U72076 ( .A(n51943), .B(n51942), .Z(n51944) );
  IV U72077 ( .A(n51944), .Z(n51945) );
  NOR U72078 ( .A(n51946), .B(n51945), .Z(n51947) );
  IV U72079 ( .A(n51947), .Z(n51950) );
  NOR U72080 ( .A(n51948), .B(n51950), .Z(n56769) );
  XOR U72081 ( .A(n56771), .B(n56769), .Z(n57126) );
  IV U72082 ( .A(n51949), .Z(n51951) );
  NOR U72083 ( .A(n51951), .B(n51950), .Z(n56763) );
  IV U72084 ( .A(n51952), .Z(n51953) );
  NOR U72085 ( .A(n51954), .B(n51953), .Z(n57125) );
  NOR U72086 ( .A(n56763), .B(n57125), .Z(n51955) );
  XOR U72087 ( .A(n57126), .B(n51955), .Z(n51956) );
  IV U72088 ( .A(n51956), .Z(n57132) );
  XOR U72089 ( .A(n57128), .B(n57132), .Z(n51957) );
  XOR U72090 ( .A(n51958), .B(n51957), .Z(n56757) );
  XOR U72091 ( .A(n57137), .B(n57139), .Z(n51959) );
  NOR U72092 ( .A(n56758), .B(n51959), .Z(n51960) );
  XOR U72093 ( .A(n56757), .B(n51960), .Z(n62153) );
  IV U72094 ( .A(n62153), .Z(n51966) );
  IV U72095 ( .A(n51961), .Z(n51962) );
  NOR U72096 ( .A(n56751), .B(n51962), .Z(n62150) );
  IV U72097 ( .A(n51963), .Z(n51965) );
  NOR U72098 ( .A(n51965), .B(n51964), .Z(n62157) );
  NOR U72099 ( .A(n62150), .B(n62157), .Z(n56749) );
  XOR U72100 ( .A(n51966), .B(n56749), .Z(n56754) );
  XOR U72101 ( .A(n51967), .B(n56754), .Z(n57147) );
  XOR U72102 ( .A(n51968), .B(n57147), .Z(n56738) );
  XOR U72103 ( .A(n51969), .B(n56738), .Z(n56735) );
  XOR U72104 ( .A(n56734), .B(n56735), .Z(n57159) );
  XOR U72105 ( .A(n57157), .B(n57159), .Z(n57161) );
  XOR U72106 ( .A(n57160), .B(n57161), .Z(n51970) );
  NOR U72107 ( .A(n51971), .B(n51970), .Z(n62176) );
  NOR U72108 ( .A(n51973), .B(n51972), .Z(n51974) );
  IV U72109 ( .A(n51974), .Z(n51975) );
  NOR U72110 ( .A(n51976), .B(n51975), .Z(n56732) );
  NOR U72111 ( .A(n57160), .B(n56732), .Z(n51977) );
  XOR U72112 ( .A(n57161), .B(n51977), .Z(n51978) );
  NOR U72113 ( .A(n51979), .B(n51978), .Z(n51980) );
  NOR U72114 ( .A(n62176), .B(n51980), .Z(n56729) );
  XOR U72115 ( .A(n56731), .B(n56729), .Z(n56724) );
  XOR U72116 ( .A(n56723), .B(n56724), .Z(n56728) );
  IV U72117 ( .A(n51981), .Z(n51985) );
  NOR U72118 ( .A(n51983), .B(n51982), .Z(n51984) );
  IV U72119 ( .A(n51984), .Z(n51990) );
  NOR U72120 ( .A(n51985), .B(n51990), .Z(n56726) );
  XOR U72121 ( .A(n56728), .B(n56726), .Z(n56722) );
  IV U72122 ( .A(n51986), .Z(n51987) );
  NOR U72123 ( .A(n51988), .B(n51987), .Z(n56718) );
  IV U72124 ( .A(n51989), .Z(n51991) );
  NOR U72125 ( .A(n51991), .B(n51990), .Z(n56720) );
  NOR U72126 ( .A(n56718), .B(n56720), .Z(n51992) );
  XOR U72127 ( .A(n56722), .B(n51992), .Z(n56712) );
  XOR U72128 ( .A(n56714), .B(n56712), .Z(n56716) );
  XOR U72129 ( .A(n56715), .B(n56716), .Z(n56705) );
  XOR U72130 ( .A(n56704), .B(n56705), .Z(n56707) );
  XOR U72131 ( .A(n51993), .B(n56707), .Z(n56700) );
  XOR U72132 ( .A(n56701), .B(n56700), .Z(n57172) );
  XOR U72133 ( .A(n57171), .B(n57172), .Z(n56698) );
  XOR U72134 ( .A(n56697), .B(n56698), .Z(n57188) );
  XOR U72135 ( .A(n51994), .B(n57188), .Z(n57184) );
  XOR U72136 ( .A(n51995), .B(n57184), .Z(n57193) );
  XOR U72137 ( .A(n51996), .B(n57193), .Z(n51997) );
  IV U72138 ( .A(n51997), .Z(n56694) );
  XOR U72139 ( .A(n51998), .B(n56694), .Z(n56688) );
  XOR U72140 ( .A(n56687), .B(n56688), .Z(n56691) );
  NOR U72141 ( .A(n51999), .B(n56681), .Z(n52000) );
  NOR U72142 ( .A(n56690), .B(n52000), .Z(n52001) );
  XOR U72143 ( .A(n56691), .B(n52001), .Z(n52002) );
  IV U72144 ( .A(n52002), .Z(n56679) );
  IV U72145 ( .A(n52003), .Z(n52005) );
  NOR U72146 ( .A(n52005), .B(n52004), .Z(n52006) );
  IV U72147 ( .A(n52006), .Z(n52010) );
  NOR U72148 ( .A(n56679), .B(n52010), .Z(n61663) );
  IV U72149 ( .A(n52007), .Z(n52009) );
  NOR U72150 ( .A(n52009), .B(n52008), .Z(n56674) );
  XOR U72151 ( .A(n56677), .B(n56679), .Z(n56675) );
  IV U72152 ( .A(n56675), .Z(n52011) );
  XOR U72153 ( .A(n56674), .B(n52011), .Z(n52013) );
  NOR U72154 ( .A(n52011), .B(n52010), .Z(n52012) );
  NOR U72155 ( .A(n52013), .B(n52012), .Z(n52014) );
  NOR U72156 ( .A(n61663), .B(n52014), .Z(n57207) );
  XOR U72157 ( .A(n57206), .B(n57207), .Z(n52019) );
  IV U72158 ( .A(n52015), .Z(n52016) );
  NOR U72159 ( .A(n52016), .B(n52021), .Z(n52017) );
  NOR U72160 ( .A(n52019), .B(n52017), .Z(n52032) );
  IV U72161 ( .A(n52018), .Z(n52026) );
  IV U72162 ( .A(n52019), .Z(n52020) );
  NOR U72163 ( .A(n52021), .B(n52020), .Z(n52022) );
  IV U72164 ( .A(n52022), .Z(n52023) );
  NOR U72165 ( .A(n52024), .B(n52023), .Z(n52025) );
  IV U72166 ( .A(n52025), .Z(n52028) );
  NOR U72167 ( .A(n52026), .B(n52028), .Z(n56673) );
  IV U72168 ( .A(n52027), .Z(n52029) );
  NOR U72169 ( .A(n52029), .B(n52028), .Z(n62231) );
  NOR U72170 ( .A(n56673), .B(n62231), .Z(n52030) );
  IV U72171 ( .A(n52030), .Z(n52031) );
  NOR U72172 ( .A(n52032), .B(n52031), .Z(n52033) );
  IV U72173 ( .A(n52033), .Z(n57213) );
  IV U72174 ( .A(n52034), .Z(n52037) );
  IV U72175 ( .A(n52035), .Z(n52036) );
  NOR U72176 ( .A(n52037), .B(n52036), .Z(n57211) );
  XOR U72177 ( .A(n57213), .B(n57211), .Z(n57215) );
  XOR U72178 ( .A(n57214), .B(n57215), .Z(n56663) );
  XOR U72179 ( .A(n52038), .B(n56663), .Z(n56661) );
  XOR U72180 ( .A(n52039), .B(n56661), .Z(n52040) );
  IV U72181 ( .A(n52040), .Z(n57225) );
  XOR U72182 ( .A(n57224), .B(n57225), .Z(n57229) );
  IV U72183 ( .A(n52041), .Z(n52043) );
  NOR U72184 ( .A(n52043), .B(n52042), .Z(n57227) );
  XOR U72185 ( .A(n57229), .B(n57227), .Z(n57232) );
  XOR U72186 ( .A(n57231), .B(n57232), .Z(n57238) );
  XOR U72187 ( .A(n57234), .B(n57238), .Z(n56654) );
  IV U72188 ( .A(n52044), .Z(n52046) );
  NOR U72189 ( .A(n52046), .B(n52045), .Z(n57237) );
  IV U72190 ( .A(n52047), .Z(n52048) );
  NOR U72191 ( .A(n52049), .B(n52048), .Z(n56653) );
  NOR U72192 ( .A(n57237), .B(n56653), .Z(n52050) );
  XOR U72193 ( .A(n56654), .B(n52050), .Z(n52051) );
  IV U72194 ( .A(n52051), .Z(n57242) );
  IV U72195 ( .A(n52052), .Z(n52054) );
  NOR U72196 ( .A(n52054), .B(n52053), .Z(n57240) );
  XOR U72197 ( .A(n57242), .B(n57240), .Z(n57244) );
  XOR U72198 ( .A(n57243), .B(n57244), .Z(n57249) );
  XOR U72199 ( .A(n57247), .B(n57249), .Z(n57251) );
  XOR U72200 ( .A(n57250), .B(n57251), .Z(n56651) );
  XOR U72201 ( .A(n56650), .B(n56651), .Z(n56645) );
  XOR U72202 ( .A(n56644), .B(n56645), .Z(n56640) );
  XOR U72203 ( .A(n52055), .B(n56640), .Z(n57260) );
  XOR U72204 ( .A(n57261), .B(n57260), .Z(n52065) );
  IV U72205 ( .A(n52065), .Z(n57263) );
  NOR U72206 ( .A(n52056), .B(n57263), .Z(n52057) );
  IV U72207 ( .A(n52057), .Z(n56637) );
  IV U72208 ( .A(n52058), .Z(n52059) );
  NOR U72209 ( .A(n52060), .B(n52059), .Z(n52067) );
  IV U72210 ( .A(n52067), .Z(n52061) );
  NOR U72211 ( .A(n56637), .B(n52061), .Z(n61623) );
  NOR U72212 ( .A(n56636), .B(n57262), .Z(n52062) );
  NOR U72213 ( .A(n52063), .B(n52062), .Z(n52064) );
  XOR U72214 ( .A(n52065), .B(n52064), .Z(n52066) );
  NOR U72215 ( .A(n52067), .B(n52066), .Z(n52068) );
  NOR U72216 ( .A(n61623), .B(n52068), .Z(n52069) );
  IV U72217 ( .A(n52069), .Z(n56629) );
  NOR U72218 ( .A(n52075), .B(n56629), .Z(n56627) );
  IV U72219 ( .A(n52070), .Z(n52072) );
  NOR U72220 ( .A(n52072), .B(n52071), .Z(n56621) );
  NOR U72221 ( .A(n52073), .B(n56630), .Z(n52074) );
  XOR U72222 ( .A(n52074), .B(n56629), .Z(n56622) );
  IV U72223 ( .A(n56622), .Z(n52076) );
  XOR U72224 ( .A(n56621), .B(n52076), .Z(n52078) );
  NOR U72225 ( .A(n52076), .B(n52075), .Z(n52077) );
  NOR U72226 ( .A(n52078), .B(n52077), .Z(n52079) );
  NOR U72227 ( .A(n56627), .B(n52079), .Z(n56624) );
  XOR U72228 ( .A(n56626), .B(n56624), .Z(n56617) );
  XOR U72229 ( .A(n56615), .B(n56617), .Z(n56610) );
  IV U72230 ( .A(n52080), .Z(n56611) );
  NOR U72231 ( .A(n52081), .B(n56611), .Z(n52082) );
  XOR U72232 ( .A(n56610), .B(n52082), .Z(n61610) );
  IV U72233 ( .A(n61610), .Z(n52095) );
  IV U72234 ( .A(n52083), .Z(n52087) );
  NOR U72235 ( .A(n52085), .B(n52084), .Z(n52086) );
  IV U72236 ( .A(n52086), .Z(n52097) );
  NOR U72237 ( .A(n52087), .B(n52097), .Z(n56606) );
  IV U72238 ( .A(n52088), .Z(n52090) );
  NOR U72239 ( .A(n52090), .B(n52089), .Z(n61608) );
  IV U72240 ( .A(n52091), .Z(n52092) );
  NOR U72241 ( .A(n56611), .B(n52092), .Z(n62296) );
  NOR U72242 ( .A(n61608), .B(n62296), .Z(n56605) );
  IV U72243 ( .A(n56605), .Z(n52093) );
  NOR U72244 ( .A(n56606), .B(n52093), .Z(n52094) );
  XOR U72245 ( .A(n52095), .B(n52094), .Z(n56600) );
  IV U72246 ( .A(n52096), .Z(n52098) );
  NOR U72247 ( .A(n52098), .B(n52097), .Z(n56599) );
  NOR U72248 ( .A(n52099), .B(n56593), .Z(n52100) );
  XOR U72249 ( .A(n56599), .B(n52100), .Z(n52101) );
  XOR U72250 ( .A(n56600), .B(n52101), .Z(n56590) );
  XOR U72251 ( .A(n56589), .B(n56590), .Z(n57274) );
  XOR U72252 ( .A(n57275), .B(n57274), .Z(n56584) );
  IV U72253 ( .A(n52102), .Z(n62323) );
  NOR U72254 ( .A(n62323), .B(n56588), .Z(n52103) );
  NOR U72255 ( .A(n52104), .B(n52103), .Z(n52105) );
  XOR U72256 ( .A(n56584), .B(n52105), .Z(n62312) );
  IV U72257 ( .A(n52106), .Z(n52107) );
  NOR U72258 ( .A(n52107), .B(n62323), .Z(n56579) );
  XOR U72259 ( .A(n62312), .B(n56579), .Z(n56583) );
  XOR U72260 ( .A(n52108), .B(n56583), .Z(n57284) );
  XOR U72261 ( .A(n57282), .B(n57284), .Z(n57287) );
  IV U72262 ( .A(n52109), .Z(n52113) );
  NOR U72263 ( .A(n52111), .B(n52110), .Z(n52112) );
  IV U72264 ( .A(n52112), .Z(n52115) );
  NOR U72265 ( .A(n52113), .B(n52115), .Z(n57285) );
  XOR U72266 ( .A(n57287), .B(n57285), .Z(n57281) );
  IV U72267 ( .A(n52114), .Z(n52116) );
  NOR U72268 ( .A(n52116), .B(n52115), .Z(n57279) );
  XOR U72269 ( .A(n57281), .B(n57279), .Z(n56572) );
  XOR U72270 ( .A(n56564), .B(n56572), .Z(n56570) );
  IV U72271 ( .A(n52117), .Z(n52118) );
  NOR U72272 ( .A(n52119), .B(n52118), .Z(n52120) );
  IV U72273 ( .A(n52120), .Z(n56569) );
  XOR U72274 ( .A(n56570), .B(n56569), .Z(n52121) );
  XOR U72275 ( .A(n52122), .B(n52121), .Z(n56561) );
  IV U72276 ( .A(n52123), .Z(n52125) );
  NOR U72277 ( .A(n52125), .B(n52124), .Z(n56559) );
  XOR U72278 ( .A(n56561), .B(n56559), .Z(n56554) );
  XOR U72279 ( .A(n56553), .B(n56554), .Z(n56558) );
  XOR U72280 ( .A(n56556), .B(n56558), .Z(n56552) );
  XOR U72281 ( .A(n52126), .B(n56552), .Z(n52127) );
  IV U72282 ( .A(n52127), .Z(n56547) );
  XOR U72283 ( .A(n56545), .B(n56547), .Z(n56532) );
  XOR U72284 ( .A(n56531), .B(n56532), .Z(n56522) );
  XOR U72285 ( .A(n56521), .B(n56522), .Z(n56525) );
  XOR U72286 ( .A(n56524), .B(n56525), .Z(n56518) );
  XOR U72287 ( .A(n56517), .B(n56518), .Z(n57302) );
  XOR U72288 ( .A(n57302), .B(n52128), .Z(n56513) );
  XOR U72289 ( .A(n52129), .B(n56513), .Z(n61556) );
  IV U72290 ( .A(n52130), .Z(n52132) );
  NOR U72291 ( .A(n52132), .B(n52131), .Z(n61559) );
  IV U72292 ( .A(n52133), .Z(n52135) );
  NOR U72293 ( .A(n52135), .B(n52134), .Z(n61555) );
  NOR U72294 ( .A(n61559), .B(n61555), .Z(n56507) );
  XOR U72295 ( .A(n61556), .B(n56507), .Z(n56504) );
  XOR U72296 ( .A(n52136), .B(n56504), .Z(n56503) );
  XOR U72297 ( .A(n52137), .B(n56503), .Z(n56499) );
  XOR U72298 ( .A(n56498), .B(n56499), .Z(n56486) );
  XOR U72299 ( .A(n52138), .B(n56486), .Z(n57314) );
  XOR U72300 ( .A(n57312), .B(n57314), .Z(n57316) );
  XOR U72301 ( .A(n57315), .B(n57316), .Z(n56482) );
  IV U72302 ( .A(n52139), .Z(n52140) );
  NOR U72303 ( .A(n52141), .B(n52140), .Z(n56481) );
  IV U72304 ( .A(n52142), .Z(n52143) );
  NOR U72305 ( .A(n52144), .B(n52143), .Z(n56479) );
  NOR U72306 ( .A(n56481), .B(n56479), .Z(n52145) );
  XOR U72307 ( .A(n56482), .B(n52145), .Z(n52146) );
  IV U72308 ( .A(n52146), .Z(n56475) );
  XOR U72309 ( .A(n56473), .B(n56475), .Z(n56478) );
  IV U72310 ( .A(n56478), .Z(n52156) );
  IV U72311 ( .A(n52147), .Z(n52148) );
  NOR U72312 ( .A(n52149), .B(n52148), .Z(n56468) );
  NOR U72313 ( .A(n52151), .B(n52150), .Z(n52152) );
  IV U72314 ( .A(n52152), .Z(n52153) );
  NOR U72315 ( .A(n52154), .B(n52153), .Z(n56476) );
  NOR U72316 ( .A(n56468), .B(n56476), .Z(n52155) );
  XOR U72317 ( .A(n52156), .B(n52155), .Z(n56471) );
  XOR U72318 ( .A(n56470), .B(n56471), .Z(n56458) );
  XOR U72319 ( .A(n52157), .B(n56458), .Z(n56455) );
  XOR U72320 ( .A(n52159), .B(n52158), .Z(n52160) );
  NOR U72321 ( .A(n52161), .B(n52160), .Z(n52162) );
  IV U72322 ( .A(n52162), .Z(n52166) );
  NOR U72323 ( .A(n52164), .B(n52163), .Z(n52165) );
  IV U72324 ( .A(n52165), .Z(n52172) );
  NOR U72325 ( .A(n52166), .B(n52172), .Z(n52167) );
  IV U72326 ( .A(n52167), .Z(n52174) );
  NOR U72327 ( .A(n56455), .B(n52174), .Z(n67856) );
  IV U72328 ( .A(n52168), .Z(n52170) );
  NOR U72329 ( .A(n52170), .B(n52169), .Z(n56448) );
  IV U72330 ( .A(n52171), .Z(n52173) );
  NOR U72331 ( .A(n52173), .B(n52172), .Z(n56454) );
  XOR U72332 ( .A(n56454), .B(n56455), .Z(n56449) );
  IV U72333 ( .A(n56449), .Z(n52175) );
  XOR U72334 ( .A(n56448), .B(n52175), .Z(n52177) );
  NOR U72335 ( .A(n52175), .B(n52174), .Z(n52176) );
  NOR U72336 ( .A(n52177), .B(n52176), .Z(n52178) );
  NOR U72337 ( .A(n67856), .B(n52178), .Z(n56452) );
  XOR U72338 ( .A(n52179), .B(n56452), .Z(n57328) );
  XOR U72339 ( .A(n57326), .B(n57328), .Z(n57335) );
  XOR U72340 ( .A(n52180), .B(n57335), .Z(n57332) );
  IV U72341 ( .A(n52185), .Z(n52181) );
  NOR U72342 ( .A(n52181), .B(n52184), .Z(n61513) );
  IV U72343 ( .A(n52182), .Z(n52189) );
  IV U72344 ( .A(n52183), .Z(n52187) );
  XOR U72345 ( .A(n52185), .B(n52184), .Z(n52186) );
  NOR U72346 ( .A(n52187), .B(n52186), .Z(n52188) );
  IV U72347 ( .A(n52188), .Z(n62427) );
  NOR U72348 ( .A(n52189), .B(n62427), .Z(n52190) );
  NOR U72349 ( .A(n61513), .B(n52190), .Z(n57333) );
  XOR U72350 ( .A(n57332), .B(n57333), .Z(n56443) );
  XOR U72351 ( .A(n56442), .B(n56443), .Z(n56446) );
  IV U72352 ( .A(n52191), .Z(n52192) );
  NOR U72353 ( .A(n52193), .B(n52192), .Z(n56445) );
  IV U72354 ( .A(n52194), .Z(n52196) );
  NOR U72355 ( .A(n52196), .B(n52195), .Z(n56439) );
  NOR U72356 ( .A(n56445), .B(n56439), .Z(n52197) );
  XOR U72357 ( .A(n56446), .B(n52197), .Z(n52198) );
  IV U72358 ( .A(n52198), .Z(n56435) );
  IV U72359 ( .A(n52199), .Z(n52201) );
  NOR U72360 ( .A(n52201), .B(n52200), .Z(n56433) );
  XOR U72361 ( .A(n56435), .B(n56433), .Z(n56438) );
  XOR U72362 ( .A(n56436), .B(n56438), .Z(n57339) );
  XOR U72363 ( .A(n57338), .B(n57339), .Z(n57342) );
  XOR U72364 ( .A(n57341), .B(n57342), .Z(n56426) );
  XOR U72365 ( .A(n52202), .B(n56426), .Z(n56424) );
  XOR U72366 ( .A(n56422), .B(n56424), .Z(n56417) );
  XOR U72367 ( .A(n56416), .B(n56417), .Z(n56420) );
  XOR U72368 ( .A(n56419), .B(n56420), .Z(n56412) );
  XOR U72369 ( .A(n56410), .B(n56412), .Z(n56407) );
  NOR U72370 ( .A(n52204), .B(n52203), .Z(n52205) );
  IV U72371 ( .A(n52205), .Z(n56406) );
  NOR U72372 ( .A(n52206), .B(n56406), .Z(n52207) );
  XOR U72373 ( .A(n56407), .B(n52207), .Z(n56404) );
  XOR U72374 ( .A(n52208), .B(n56404), .Z(n56395) );
  IV U72375 ( .A(n52209), .Z(n52211) );
  NOR U72376 ( .A(n52211), .B(n52210), .Z(n56397) );
  IV U72377 ( .A(n52212), .Z(n52215) );
  NOR U72378 ( .A(n52213), .B(n52218), .Z(n52214) );
  IV U72379 ( .A(n52214), .Z(n52221) );
  NOR U72380 ( .A(n52215), .B(n52221), .Z(n56394) );
  NOR U72381 ( .A(n56397), .B(n56394), .Z(n52216) );
  XOR U72382 ( .A(n56395), .B(n52216), .Z(n56393) );
  IV U72383 ( .A(n52217), .Z(n52219) );
  NOR U72384 ( .A(n52219), .B(n52218), .Z(n56388) );
  IV U72385 ( .A(n52220), .Z(n52222) );
  NOR U72386 ( .A(n52222), .B(n52221), .Z(n56391) );
  NOR U72387 ( .A(n56388), .B(n56391), .Z(n52223) );
  XOR U72388 ( .A(n56393), .B(n52223), .Z(n57353) );
  IV U72389 ( .A(n52224), .Z(n52226) );
  NOR U72390 ( .A(n52226), .B(n52225), .Z(n61465) );
  IV U72391 ( .A(n52227), .Z(n52228) );
  NOR U72392 ( .A(n57356), .B(n52228), .Z(n61460) );
  NOR U72393 ( .A(n61465), .B(n61460), .Z(n57354) );
  XOR U72394 ( .A(n57353), .B(n57354), .Z(n57355) );
  XOR U72395 ( .A(n52229), .B(n57355), .Z(n57364) );
  XOR U72396 ( .A(n52230), .B(n57364), .Z(n56386) );
  XOR U72397 ( .A(n56385), .B(n56386), .Z(n57376) );
  XOR U72398 ( .A(n52231), .B(n57376), .Z(n52232) );
  IV U72399 ( .A(n52232), .Z(n56381) );
  XOR U72400 ( .A(n56379), .B(n56381), .Z(n56383) );
  XOR U72401 ( .A(n56382), .B(n56383), .Z(n57385) );
  XOR U72402 ( .A(n57384), .B(n57385), .Z(n57389) );
  IV U72403 ( .A(n52233), .Z(n52235) );
  NOR U72404 ( .A(n52235), .B(n52234), .Z(n57387) );
  XOR U72405 ( .A(n57389), .B(n57387), .Z(n56377) );
  XOR U72406 ( .A(n56376), .B(n56377), .Z(n56371) );
  XOR U72407 ( .A(n56370), .B(n56371), .Z(n56375) );
  IV U72408 ( .A(n52236), .Z(n52237) );
  NOR U72409 ( .A(n52238), .B(n52237), .Z(n56373) );
  XOR U72410 ( .A(n56375), .B(n56373), .Z(n56365) );
  NOR U72411 ( .A(n52239), .B(n56358), .Z(n56364) );
  NOR U72412 ( .A(n56364), .B(n52240), .Z(n52241) );
  XOR U72413 ( .A(n56365), .B(n52241), .Z(n52242) );
  IV U72414 ( .A(n52242), .Z(n56355) );
  IV U72415 ( .A(n52243), .Z(n52245) );
  NOR U72416 ( .A(n52245), .B(n52244), .Z(n56353) );
  IV U72417 ( .A(n52246), .Z(n52248) );
  IV U72418 ( .A(n52247), .Z(n56345) );
  NOR U72419 ( .A(n52248), .B(n56345), .Z(n56351) );
  NOR U72420 ( .A(n56353), .B(n56351), .Z(n52249) );
  XOR U72421 ( .A(n56355), .B(n52249), .Z(n56341) );
  NOR U72422 ( .A(n52250), .B(n56345), .Z(n52254) );
  IV U72423 ( .A(n52251), .Z(n52253) );
  NOR U72424 ( .A(n52253), .B(n52252), .Z(n56340) );
  NOR U72425 ( .A(n52254), .B(n56340), .Z(n52255) );
  XOR U72426 ( .A(n56341), .B(n52255), .Z(n56336) );
  IV U72427 ( .A(n52256), .Z(n52257) );
  NOR U72428 ( .A(n52258), .B(n52257), .Z(n56334) );
  XOR U72429 ( .A(n56336), .B(n56334), .Z(n56339) );
  XOR U72430 ( .A(n56337), .B(n56339), .Z(n57393) );
  NOR U72431 ( .A(n52264), .B(n57393), .Z(n62513) );
  NOR U72432 ( .A(n52260), .B(n52259), .Z(n56331) );
  IV U72433 ( .A(n52261), .Z(n52262) );
  NOR U72434 ( .A(n52263), .B(n52262), .Z(n57392) );
  XOR U72435 ( .A(n57392), .B(n57393), .Z(n56332) );
  IV U72436 ( .A(n56332), .Z(n52265) );
  XOR U72437 ( .A(n56331), .B(n52265), .Z(n52267) );
  NOR U72438 ( .A(n52265), .B(n52264), .Z(n52266) );
  NOR U72439 ( .A(n52267), .B(n52266), .Z(n52268) );
  NOR U72440 ( .A(n62513), .B(n52268), .Z(n56324) );
  IV U72441 ( .A(n52269), .Z(n52277) );
  XOR U72442 ( .A(n52271), .B(n52270), .Z(n52274) );
  IV U72443 ( .A(n52272), .Z(n52273) );
  NOR U72444 ( .A(n52274), .B(n52273), .Z(n52275) );
  IV U72445 ( .A(n52275), .Z(n52276) );
  NOR U72446 ( .A(n52277), .B(n52276), .Z(n56325) );
  NOR U72447 ( .A(n56325), .B(n52278), .Z(n52279) );
  XOR U72448 ( .A(n56324), .B(n52279), .Z(n56328) );
  XOR U72449 ( .A(n56327), .B(n56328), .Z(n57409) );
  XOR U72450 ( .A(n57402), .B(n57409), .Z(n56322) );
  XOR U72451 ( .A(n56321), .B(n56322), .Z(n56316) );
  XOR U72452 ( .A(n56315), .B(n56316), .Z(n56320) );
  IV U72453 ( .A(n52280), .Z(n52282) );
  NOR U72454 ( .A(n52282), .B(n52281), .Z(n56318) );
  XOR U72455 ( .A(n56320), .B(n56318), .Z(n57426) );
  XOR U72456 ( .A(n57425), .B(n57426), .Z(n57435) );
  XOR U72457 ( .A(n52283), .B(n57435), .Z(n56313) );
  XOR U72458 ( .A(n56310), .B(n56313), .Z(n56308) );
  IV U72459 ( .A(n52284), .Z(n52287) );
  NOR U72460 ( .A(n52285), .B(n52287), .Z(n56312) );
  IV U72461 ( .A(n52286), .Z(n52290) );
  NOR U72462 ( .A(n52288), .B(n52287), .Z(n52289) );
  IV U72463 ( .A(n52289), .Z(n52293) );
  NOR U72464 ( .A(n52290), .B(n52293), .Z(n56306) );
  NOR U72465 ( .A(n56312), .B(n56306), .Z(n52291) );
  XOR U72466 ( .A(n56308), .B(n52291), .Z(n57447) );
  IV U72467 ( .A(n52292), .Z(n52294) );
  NOR U72468 ( .A(n52294), .B(n52293), .Z(n52295) );
  IV U72469 ( .A(n52295), .Z(n57448) );
  XOR U72470 ( .A(n57447), .B(n57448), .Z(n57451) );
  XOR U72471 ( .A(n57450), .B(n57451), .Z(n61393) );
  XOR U72472 ( .A(n57453), .B(n61393), .Z(n56303) );
  IV U72473 ( .A(n52296), .Z(n52297) );
  NOR U72474 ( .A(n52299), .B(n52297), .Z(n56302) );
  IV U72475 ( .A(n52298), .Z(n52300) );
  NOR U72476 ( .A(n52300), .B(n52299), .Z(n57454) );
  NOR U72477 ( .A(n56302), .B(n57454), .Z(n52301) );
  XOR U72478 ( .A(n56303), .B(n52301), .Z(n57468) );
  XOR U72479 ( .A(n57460), .B(n57468), .Z(n57475) );
  IV U72480 ( .A(n52302), .Z(n52303) );
  NOR U72481 ( .A(n52304), .B(n52303), .Z(n52311) );
  IV U72482 ( .A(n52311), .Z(n52305) );
  NOR U72483 ( .A(n57475), .B(n52305), .Z(n62565) );
  IV U72484 ( .A(n52306), .Z(n52308) );
  NOR U72485 ( .A(n52308), .B(n52307), .Z(n57467) );
  NOR U72486 ( .A(n57460), .B(n57467), .Z(n52309) );
  XOR U72487 ( .A(n57468), .B(n52309), .Z(n52310) );
  NOR U72488 ( .A(n52311), .B(n52310), .Z(n52312) );
  NOR U72489 ( .A(n62565), .B(n52312), .Z(n57472) );
  XOR U72490 ( .A(n57471), .B(n57472), .Z(n52313) );
  XOR U72491 ( .A(n57476), .B(n52313), .Z(n57482) );
  NOR U72492 ( .A(n52315), .B(n52314), .Z(n52316) );
  IV U72493 ( .A(n52316), .Z(n52317) );
  NOR U72494 ( .A(n52318), .B(n52317), .Z(n57479) );
  IV U72495 ( .A(n52319), .Z(n52320) );
  NOR U72496 ( .A(n52323), .B(n52320), .Z(n57481) );
  NOR U72497 ( .A(n57479), .B(n57481), .Z(n52321) );
  XOR U72498 ( .A(n57482), .B(n52321), .Z(n57484) );
  IV U72499 ( .A(n52322), .Z(n52324) );
  NOR U72500 ( .A(n52324), .B(n52323), .Z(n52325) );
  IV U72501 ( .A(n52325), .Z(n57485) );
  XOR U72502 ( .A(n57484), .B(n57485), .Z(n57489) );
  XOR U72503 ( .A(n57487), .B(n57489), .Z(n56298) );
  XOR U72504 ( .A(n52326), .B(n56298), .Z(n52327) );
  IV U72505 ( .A(n52327), .Z(n57492) );
  XOR U72506 ( .A(n57490), .B(n57492), .Z(n57494) );
  XOR U72507 ( .A(n57493), .B(n57494), .Z(n56295) );
  IV U72508 ( .A(n52328), .Z(n52333) );
  IV U72509 ( .A(n52329), .Z(n52330) );
  NOR U72510 ( .A(n52331), .B(n52330), .Z(n52332) );
  IV U72511 ( .A(n52332), .Z(n52338) );
  NOR U72512 ( .A(n52333), .B(n52338), .Z(n56293) );
  XOR U72513 ( .A(n56295), .B(n56293), .Z(n56291) );
  IV U72514 ( .A(n52334), .Z(n52336) );
  NOR U72515 ( .A(n52336), .B(n52335), .Z(n56282) );
  IV U72516 ( .A(n52337), .Z(n52339) );
  NOR U72517 ( .A(n52339), .B(n52338), .Z(n56283) );
  NOR U72518 ( .A(n56282), .B(n56283), .Z(n52340) );
  XOR U72519 ( .A(n56291), .B(n52340), .Z(n56279) );
  XOR U72520 ( .A(n52341), .B(n56279), .Z(n57504) );
  XOR U72521 ( .A(n52342), .B(n57504), .Z(n56275) );
  XOR U72522 ( .A(n56274), .B(n56275), .Z(n56268) );
  XOR U72523 ( .A(n56267), .B(n56268), .Z(n56271) );
  XOR U72524 ( .A(n56270), .B(n56271), .Z(n52343) );
  NOR U72525 ( .A(n52344), .B(n52343), .Z(n66921) );
  IV U72526 ( .A(n52345), .Z(n52347) );
  NOR U72527 ( .A(n52347), .B(n52346), .Z(n56264) );
  NOR U72528 ( .A(n56270), .B(n56264), .Z(n52348) );
  XOR U72529 ( .A(n56271), .B(n52348), .Z(n52349) );
  NOR U72530 ( .A(n52350), .B(n52349), .Z(n52351) );
  NOR U72531 ( .A(n66921), .B(n52351), .Z(n52352) );
  IV U72532 ( .A(n52352), .Z(n56263) );
  IV U72533 ( .A(n52353), .Z(n52355) );
  NOR U72534 ( .A(n52355), .B(n52354), .Z(n56261) );
  XOR U72535 ( .A(n56263), .B(n56261), .Z(n68092) );
  XOR U72536 ( .A(n52356), .B(n68092), .Z(n52357) );
  IV U72537 ( .A(n52357), .Z(n57512) );
  XOR U72538 ( .A(n57511), .B(n57512), .Z(n57517) );
  IV U72539 ( .A(n52358), .Z(n52365) );
  NOR U72540 ( .A(n52365), .B(n52359), .Z(n57516) );
  IV U72541 ( .A(n52360), .Z(n52362) );
  NOR U72542 ( .A(n52362), .B(n52361), .Z(n56258) );
  NOR U72543 ( .A(n57516), .B(n56258), .Z(n52363) );
  XOR U72544 ( .A(n57517), .B(n52363), .Z(n56255) );
  IV U72545 ( .A(n52364), .Z(n52369) );
  NOR U72546 ( .A(n52366), .B(n52365), .Z(n52367) );
  IV U72547 ( .A(n52367), .Z(n52368) );
  NOR U72548 ( .A(n52369), .B(n52368), .Z(n52370) );
  IV U72549 ( .A(n52370), .Z(n56256) );
  XOR U72550 ( .A(n56255), .B(n56256), .Z(n57522) );
  XOR U72551 ( .A(n57520), .B(n57522), .Z(n57529) );
  XOR U72552 ( .A(n52371), .B(n57529), .Z(n57534) );
  XOR U72553 ( .A(n52372), .B(n57534), .Z(n62659) );
  IV U72554 ( .A(n52373), .Z(n52374) );
  NOR U72555 ( .A(n52375), .B(n52374), .Z(n62658) );
  IV U72556 ( .A(n52376), .Z(n52380) );
  NOR U72557 ( .A(n52378), .B(n52377), .Z(n52379) );
  IV U72558 ( .A(n52379), .Z(n52382) );
  NOR U72559 ( .A(n52380), .B(n52382), .Z(n62676) );
  NOR U72560 ( .A(n62658), .B(n62676), .Z(n56253) );
  IV U72561 ( .A(n52381), .Z(n52383) );
  NOR U72562 ( .A(n52383), .B(n52382), .Z(n56251) );
  XOR U72563 ( .A(n56253), .B(n56251), .Z(n52384) );
  XOR U72564 ( .A(n62659), .B(n52384), .Z(n52385) );
  IV U72565 ( .A(n52385), .Z(n56247) );
  XOR U72566 ( .A(n56245), .B(n56247), .Z(n56249) );
  XOR U72567 ( .A(n56248), .B(n56249), .Z(n56240) );
  XOR U72568 ( .A(n56239), .B(n56240), .Z(n56243) );
  NOR U72569 ( .A(n56242), .B(n56237), .Z(n52386) );
  XOR U72570 ( .A(n56243), .B(n52386), .Z(n56231) );
  XOR U72571 ( .A(n52387), .B(n56231), .Z(n57557) );
  XOR U72572 ( .A(n52388), .B(n57557), .Z(n56219) );
  XOR U72573 ( .A(n52389), .B(n56219), .Z(n56213) );
  XOR U72574 ( .A(n56211), .B(n56213), .Z(n56215) );
  XOR U72575 ( .A(n56214), .B(n56215), .Z(n56205) );
  XOR U72576 ( .A(n56204), .B(n56205), .Z(n56209) );
  IV U72577 ( .A(n52390), .Z(n52392) );
  NOR U72578 ( .A(n52392), .B(n52391), .Z(n56207) );
  XOR U72579 ( .A(n56209), .B(n56207), .Z(n56202) );
  IV U72580 ( .A(n52393), .Z(n56199) );
  XOR U72581 ( .A(n52394), .B(n56199), .Z(n52395) );
  NOR U72582 ( .A(n56200), .B(n52395), .Z(n52396) );
  XOR U72583 ( .A(n56202), .B(n52396), .Z(n56188) );
  IV U72584 ( .A(n52397), .Z(n52399) );
  NOR U72585 ( .A(n52399), .B(n52398), .Z(n56181) );
  IV U72586 ( .A(n52400), .Z(n52402) );
  NOR U72587 ( .A(n52402), .B(n52401), .Z(n56187) );
  NOR U72588 ( .A(n56181), .B(n56187), .Z(n52403) );
  XOR U72589 ( .A(n56188), .B(n52403), .Z(n56176) );
  IV U72590 ( .A(n52404), .Z(n52406) );
  NOR U72591 ( .A(n52406), .B(n52405), .Z(n56183) );
  IV U72592 ( .A(n52407), .Z(n52410) );
  NOR U72593 ( .A(n52408), .B(n52418), .Z(n52409) );
  IV U72594 ( .A(n52409), .Z(n52412) );
  NOR U72595 ( .A(n52410), .B(n52412), .Z(n56177) );
  IV U72596 ( .A(n52411), .Z(n52413) );
  NOR U72597 ( .A(n52413), .B(n52412), .Z(n56179) );
  NOR U72598 ( .A(n56177), .B(n56179), .Z(n52414) );
  IV U72599 ( .A(n52414), .Z(n52415) );
  NOR U72600 ( .A(n56183), .B(n52415), .Z(n52416) );
  XOR U72601 ( .A(n56176), .B(n52416), .Z(n56171) );
  IV U72602 ( .A(n52417), .Z(n52419) );
  NOR U72603 ( .A(n52419), .B(n52418), .Z(n56168) );
  XOR U72604 ( .A(n56171), .B(n56168), .Z(n56164) );
  XOR U72605 ( .A(n52420), .B(n56164), .Z(n56161) );
  IV U72606 ( .A(n52421), .Z(n52423) );
  NOR U72607 ( .A(n52423), .B(n52422), .Z(n56160) );
  IV U72608 ( .A(n52424), .Z(n52425) );
  NOR U72609 ( .A(n52426), .B(n52425), .Z(n56158) );
  NOR U72610 ( .A(n56160), .B(n56158), .Z(n52427) );
  XOR U72611 ( .A(n56161), .B(n52427), .Z(n57565) );
  XOR U72612 ( .A(n52428), .B(n57565), .Z(n56145) );
  XOR U72613 ( .A(n52429), .B(n56145), .Z(n61311) );
  IV U72614 ( .A(n52430), .Z(n52432) );
  NOR U72615 ( .A(n52432), .B(n52431), .Z(n61309) );
  NOR U72616 ( .A(n61314), .B(n61309), .Z(n57570) );
  XOR U72617 ( .A(n61311), .B(n57570), .Z(n52433) );
  IV U72618 ( .A(n52433), .Z(n57572) );
  XOR U72619 ( .A(n57571), .B(n57572), .Z(n57577) );
  XOR U72620 ( .A(n57576), .B(n57577), .Z(n57581) );
  XOR U72621 ( .A(n52434), .B(n57581), .Z(n57587) );
  XOR U72622 ( .A(n57585), .B(n57587), .Z(n56139) );
  XOR U72623 ( .A(n56138), .B(n56139), .Z(n56143) );
  XOR U72624 ( .A(n56141), .B(n56143), .Z(n61299) );
  XOR U72625 ( .A(n52435), .B(n61299), .Z(n57598) );
  XOR U72626 ( .A(n57597), .B(n57598), .Z(n57604) );
  IV U72627 ( .A(n52436), .Z(n52438) );
  NOR U72628 ( .A(n52438), .B(n52437), .Z(n57602) );
  XOR U72629 ( .A(n57604), .B(n57602), .Z(n61290) );
  IV U72630 ( .A(n52439), .Z(n52440) );
  NOR U72631 ( .A(n52441), .B(n52440), .Z(n62781) );
  IV U72632 ( .A(n52442), .Z(n52443) );
  NOR U72633 ( .A(n57612), .B(n52443), .Z(n61289) );
  NOR U72634 ( .A(n62781), .B(n61289), .Z(n57605) );
  XOR U72635 ( .A(n61290), .B(n57605), .Z(n52444) );
  IV U72636 ( .A(n52444), .Z(n57609) );
  XOR U72637 ( .A(n57608), .B(n57609), .Z(n57611) );
  XOR U72638 ( .A(n52445), .B(n57611), .Z(n57618) );
  XOR U72639 ( .A(n57619), .B(n57618), .Z(n57628) );
  XOR U72640 ( .A(n52446), .B(n57628), .Z(n57624) );
  IV U72641 ( .A(n52447), .Z(n52448) );
  NOR U72642 ( .A(n52448), .B(n52451), .Z(n52449) );
  IV U72643 ( .A(n52449), .Z(n57625) );
  XOR U72644 ( .A(n57624), .B(n57625), .Z(n56134) );
  IV U72645 ( .A(n52450), .Z(n52452) );
  NOR U72646 ( .A(n52452), .B(n52451), .Z(n57630) );
  IV U72647 ( .A(n52453), .Z(n52460) );
  IV U72648 ( .A(n52454), .Z(n52455) );
  NOR U72649 ( .A(n52460), .B(n52455), .Z(n56132) );
  NOR U72650 ( .A(n57630), .B(n56132), .Z(n52456) );
  XOR U72651 ( .A(n56134), .B(n52456), .Z(n52457) );
  IV U72652 ( .A(n52457), .Z(n56128) );
  IV U72653 ( .A(n52458), .Z(n52459) );
  NOR U72654 ( .A(n52460), .B(n52459), .Z(n56126) );
  XOR U72655 ( .A(n56128), .B(n56126), .Z(n56130) );
  XOR U72656 ( .A(n52461), .B(n56130), .Z(n52462) );
  IV U72657 ( .A(n52462), .Z(n57640) );
  XOR U72658 ( .A(n57638), .B(n57640), .Z(n57642) );
  XOR U72659 ( .A(n57641), .B(n57642), .Z(n57646) );
  XOR U72660 ( .A(n56115), .B(n57646), .Z(n56111) );
  XOR U72661 ( .A(n56110), .B(n56111), .Z(n57661) );
  IV U72662 ( .A(n52463), .Z(n52464) );
  NOR U72663 ( .A(n57647), .B(n52464), .Z(n56113) );
  NOR U72664 ( .A(n52466), .B(n52465), .Z(n57660) );
  NOR U72665 ( .A(n56113), .B(n57660), .Z(n52467) );
  XOR U72666 ( .A(n57661), .B(n52467), .Z(n52468) );
  IV U72667 ( .A(n52468), .Z(n57659) );
  IV U72668 ( .A(n52473), .Z(n52470) );
  IV U72669 ( .A(n52469), .Z(n56098) );
  NOR U72670 ( .A(n52470), .B(n56098), .Z(n52471) );
  IV U72671 ( .A(n52471), .Z(n52476) );
  NOR U72672 ( .A(n57659), .B(n52476), .Z(n61248) );
  IV U72673 ( .A(n52472), .Z(n52475) );
  XOR U72674 ( .A(n52473), .B(n56098), .Z(n52474) );
  NOR U72675 ( .A(n52475), .B(n52474), .Z(n56107) );
  XOR U72676 ( .A(n57657), .B(n57659), .Z(n56108) );
  IV U72677 ( .A(n56108), .Z(n52477) );
  XOR U72678 ( .A(n56107), .B(n52477), .Z(n52479) );
  NOR U72679 ( .A(n52477), .B(n52476), .Z(n52478) );
  NOR U72680 ( .A(n52479), .B(n52478), .Z(n52480) );
  NOR U72681 ( .A(n61248), .B(n52480), .Z(n56094) );
  IV U72682 ( .A(n52481), .Z(n52482) );
  NOR U72683 ( .A(n52482), .B(n56098), .Z(n52486) );
  IV U72684 ( .A(n52483), .Z(n52485) );
  NOR U72685 ( .A(n52485), .B(n52484), .Z(n56093) );
  NOR U72686 ( .A(n52486), .B(n56093), .Z(n52487) );
  XOR U72687 ( .A(n56094), .B(n52487), .Z(n56092) );
  XOR U72688 ( .A(n56090), .B(n56092), .Z(n56087) );
  XOR U72689 ( .A(n52488), .B(n56087), .Z(n56076) );
  XOR U72690 ( .A(n52489), .B(n56076), .Z(n56080) );
  XOR U72691 ( .A(n52490), .B(n56080), .Z(n57674) );
  XOR U72692 ( .A(n57672), .B(n57674), .Z(n57677) );
  IV U72693 ( .A(n52491), .Z(n52493) );
  NOR U72694 ( .A(n52493), .B(n52492), .Z(n57675) );
  XOR U72695 ( .A(n57677), .B(n57675), .Z(n52494) );
  XOR U72696 ( .A(n52495), .B(n52494), .Z(n56067) );
  XOR U72697 ( .A(n56068), .B(n56067), .Z(n57683) );
  XOR U72698 ( .A(n57684), .B(n57683), .Z(n57681) );
  IV U72699 ( .A(n52496), .Z(n52497) );
  NOR U72700 ( .A(n52498), .B(n52497), .Z(n57685) );
  IV U72701 ( .A(n52499), .Z(n52501) );
  NOR U72702 ( .A(n52501), .B(n52500), .Z(n57680) );
  NOR U72703 ( .A(n57685), .B(n57680), .Z(n52502) );
  XOR U72704 ( .A(n57681), .B(n52502), .Z(n56066) );
  XOR U72705 ( .A(n56064), .B(n56066), .Z(n68275) );
  XOR U72706 ( .A(n52503), .B(n68275), .Z(n52504) );
  IV U72707 ( .A(n52504), .Z(n57698) );
  XOR U72708 ( .A(n57697), .B(n57698), .Z(n56058) );
  XOR U72709 ( .A(n56057), .B(n56058), .Z(n62855) );
  XOR U72710 ( .A(n56060), .B(n62855), .Z(n56052) );
  XOR U72711 ( .A(n56051), .B(n56052), .Z(n56055) );
  XOR U72712 ( .A(n56054), .B(n56055), .Z(n56046) );
  IV U72713 ( .A(n52505), .Z(n52507) );
  NOR U72714 ( .A(n52507), .B(n52506), .Z(n56047) );
  IV U72715 ( .A(n52508), .Z(n52509) );
  NOR U72716 ( .A(n52510), .B(n52509), .Z(n56048) );
  NOR U72717 ( .A(n56047), .B(n56048), .Z(n52511) );
  XOR U72718 ( .A(n56046), .B(n52511), .Z(n56039) );
  XOR U72719 ( .A(n52512), .B(n56039), .Z(n66706) );
  NOR U72720 ( .A(n52514), .B(n52513), .Z(n66707) );
  NOR U72721 ( .A(n66707), .B(n57703), .Z(n52515) );
  XOR U72722 ( .A(n66706), .B(n52515), .Z(n56036) );
  XOR U72723 ( .A(n52516), .B(n56036), .Z(n62895) );
  XOR U72724 ( .A(n56031), .B(n62895), .Z(n56032) );
  XOR U72725 ( .A(n56033), .B(n56032), .Z(n56029) );
  IV U72726 ( .A(n52517), .Z(n52518) );
  NOR U72727 ( .A(n52519), .B(n52518), .Z(n57711) );
  IV U72728 ( .A(n52520), .Z(n52521) );
  NOR U72729 ( .A(n52522), .B(n52521), .Z(n56028) );
  NOR U72730 ( .A(n57711), .B(n56028), .Z(n52523) );
  XOR U72731 ( .A(n56029), .B(n52523), .Z(n52524) );
  NOR U72732 ( .A(n52525), .B(n52524), .Z(n52528) );
  IV U72733 ( .A(n52525), .Z(n52527) );
  XOR U72734 ( .A(n57711), .B(n56029), .Z(n52526) );
  NOR U72735 ( .A(n52527), .B(n52526), .Z(n68306) );
  NOR U72736 ( .A(n52528), .B(n68306), .Z(n56023) );
  NOR U72737 ( .A(n52530), .B(n52529), .Z(n56025) );
  NOR U72738 ( .A(n56022), .B(n56025), .Z(n52531) );
  XOR U72739 ( .A(n56023), .B(n52531), .Z(n56021) );
  XOR U72740 ( .A(n52532), .B(n56021), .Z(n52533) );
  IV U72741 ( .A(n52533), .Z(n57717) );
  XOR U72742 ( .A(n57715), .B(n57717), .Z(n57719) );
  XOR U72743 ( .A(n57718), .B(n57719), .Z(n56013) );
  XOR U72744 ( .A(n56011), .B(n56013), .Z(n56015) );
  XOR U72745 ( .A(n56014), .B(n56015), .Z(n57725) );
  XOR U72746 ( .A(n57723), .B(n57725), .Z(n57728) );
  XOR U72747 ( .A(n52534), .B(n57728), .Z(n56003) );
  XOR U72748 ( .A(n56006), .B(n56003), .Z(n55998) );
  IV U72749 ( .A(n52535), .Z(n52537) );
  NOR U72750 ( .A(n52537), .B(n52536), .Z(n56004) );
  IV U72751 ( .A(n52538), .Z(n52540) );
  NOR U72752 ( .A(n52540), .B(n52539), .Z(n55997) );
  NOR U72753 ( .A(n56004), .B(n55997), .Z(n52541) );
  XOR U72754 ( .A(n55998), .B(n52541), .Z(n55994) );
  IV U72755 ( .A(n52542), .Z(n52544) );
  NOR U72756 ( .A(n52544), .B(n52543), .Z(n56000) );
  IV U72757 ( .A(n52550), .Z(n52545) );
  NOR U72758 ( .A(n52545), .B(n52549), .Z(n55995) );
  NOR U72759 ( .A(n56000), .B(n55995), .Z(n52546) );
  XOR U72760 ( .A(n55994), .B(n52546), .Z(n55993) );
  IV U72761 ( .A(n52547), .Z(n52555) );
  IV U72762 ( .A(n52548), .Z(n52552) );
  XOR U72763 ( .A(n52550), .B(n52549), .Z(n52551) );
  NOR U72764 ( .A(n52552), .B(n52551), .Z(n52553) );
  IV U72765 ( .A(n52553), .Z(n52554) );
  NOR U72766 ( .A(n52555), .B(n52554), .Z(n55991) );
  XOR U72767 ( .A(n55993), .B(n55991), .Z(n57732) );
  XOR U72768 ( .A(n57733), .B(n57732), .Z(n55988) );
  IV U72769 ( .A(n52556), .Z(n52558) );
  NOR U72770 ( .A(n52558), .B(n52557), .Z(n57734) );
  IV U72771 ( .A(n52559), .Z(n52561) );
  NOR U72772 ( .A(n52561), .B(n52560), .Z(n55989) );
  NOR U72773 ( .A(n57734), .B(n55989), .Z(n52562) );
  XOR U72774 ( .A(n55988), .B(n52562), .Z(n55983) );
  XOR U72775 ( .A(n55982), .B(n55983), .Z(n55986) );
  XOR U72776 ( .A(n55985), .B(n55986), .Z(n57741) );
  XOR U72777 ( .A(n57740), .B(n57741), .Z(n57744) );
  XOR U72778 ( .A(n57743), .B(n57744), .Z(n55980) );
  XOR U72779 ( .A(n52563), .B(n55980), .Z(n52564) );
  IV U72780 ( .A(n52564), .Z(n55978) );
  IV U72781 ( .A(n52565), .Z(n52567) );
  NOR U72782 ( .A(n52567), .B(n52566), .Z(n55976) );
  XOR U72783 ( .A(n55978), .B(n55976), .Z(n57750) );
  IV U72784 ( .A(n52568), .Z(n52569) );
  NOR U72785 ( .A(n52570), .B(n52569), .Z(n55972) );
  NOR U72786 ( .A(n52572), .B(n52571), .Z(n57749) );
  NOR U72787 ( .A(n55972), .B(n57749), .Z(n52573) );
  XOR U72788 ( .A(n57750), .B(n52573), .Z(n55964) );
  NOR U72789 ( .A(n52575), .B(n52574), .Z(n55965) );
  IV U72790 ( .A(n52576), .Z(n52578) );
  IV U72791 ( .A(n52577), .Z(n52581) );
  NOR U72792 ( .A(n52578), .B(n52581), .Z(n57753) );
  IV U72793 ( .A(n52579), .Z(n52580) );
  NOR U72794 ( .A(n52581), .B(n52580), .Z(n57755) );
  XOR U72795 ( .A(n57753), .B(n57755), .Z(n52582) );
  NOR U72796 ( .A(n55965), .B(n52582), .Z(n52583) );
  XOR U72797 ( .A(n55964), .B(n52583), .Z(n55968) );
  IV U72798 ( .A(n52584), .Z(n52585) );
  NOR U72799 ( .A(n52585), .B(n52587), .Z(n55962) );
  IV U72800 ( .A(n52586), .Z(n52588) );
  NOR U72801 ( .A(n52588), .B(n52587), .Z(n55967) );
  NOR U72802 ( .A(n55962), .B(n55967), .Z(n52589) );
  XOR U72803 ( .A(n55968), .B(n52589), .Z(n55956) );
  XOR U72804 ( .A(n52590), .B(n55956), .Z(n57762) );
  XOR U72805 ( .A(n52591), .B(n57762), .Z(n55950) );
  XOR U72806 ( .A(n55951), .B(n55950), .Z(n57764) );
  XOR U72807 ( .A(n57763), .B(n57764), .Z(n57768) );
  XOR U72808 ( .A(n52592), .B(n57768), .Z(n55946) );
  XOR U72809 ( .A(n55944), .B(n55946), .Z(n55948) );
  XOR U72810 ( .A(n55947), .B(n55948), .Z(n57779) );
  XOR U72811 ( .A(n57777), .B(n57779), .Z(n57781) );
  XOR U72812 ( .A(n57780), .B(n57781), .Z(n57788) );
  XOR U72813 ( .A(n57787), .B(n57788), .Z(n55942) );
  XOR U72814 ( .A(n55940), .B(n55942), .Z(n57786) );
  XOR U72815 ( .A(n57784), .B(n57786), .Z(n57796) );
  XOR U72816 ( .A(n57795), .B(n57796), .Z(n57799) );
  XOR U72817 ( .A(n57798), .B(n57799), .Z(n55938) );
  XOR U72818 ( .A(n52593), .B(n55938), .Z(n52594) );
  IV U72819 ( .A(n52594), .Z(n55930) );
  XOR U72820 ( .A(n55929), .B(n55930), .Z(n55933) );
  XOR U72821 ( .A(n55932), .B(n55933), .Z(n57812) );
  IV U72822 ( .A(n52595), .Z(n57806) );
  NOR U72823 ( .A(n57806), .B(n52597), .Z(n52601) );
  IV U72824 ( .A(n52596), .Z(n52600) );
  NOR U72825 ( .A(n52598), .B(n52597), .Z(n52599) );
  IV U72826 ( .A(n52599), .Z(n52604) );
  NOR U72827 ( .A(n52600), .B(n52604), .Z(n57810) );
  NOR U72828 ( .A(n52601), .B(n57810), .Z(n52602) );
  XOR U72829 ( .A(n57812), .B(n52602), .Z(n57807) );
  IV U72830 ( .A(n52603), .Z(n52605) );
  NOR U72831 ( .A(n52605), .B(n52604), .Z(n52606) );
  IV U72832 ( .A(n52606), .Z(n57808) );
  XOR U72833 ( .A(n57807), .B(n57808), .Z(n55922) );
  XOR U72834 ( .A(n52607), .B(n55922), .Z(n55917) );
  IV U72835 ( .A(n52608), .Z(n52610) );
  NOR U72836 ( .A(n52610), .B(n52609), .Z(n55916) );
  IV U72837 ( .A(n52611), .Z(n52613) );
  NOR U72838 ( .A(n52613), .B(n52612), .Z(n52614) );
  IV U72839 ( .A(n52614), .Z(n52615) );
  NOR U72840 ( .A(n52616), .B(n52615), .Z(n55925) );
  NOR U72841 ( .A(n55916), .B(n55925), .Z(n52617) );
  XOR U72842 ( .A(n55917), .B(n52617), .Z(n55909) );
  IV U72843 ( .A(n52618), .Z(n52620) );
  NOR U72844 ( .A(n52620), .B(n52619), .Z(n52621) );
  IV U72845 ( .A(n52621), .Z(n52627) );
  NOR U72846 ( .A(n55909), .B(n52627), .Z(n62978) );
  NOR U72847 ( .A(n52622), .B(n55908), .Z(n52623) );
  XOR U72848 ( .A(n52623), .B(n55909), .Z(n55902) );
  IV U72849 ( .A(n52624), .Z(n52626) );
  NOR U72850 ( .A(n52626), .B(n52625), .Z(n52628) );
  IV U72851 ( .A(n52628), .Z(n55901) );
  XOR U72852 ( .A(n55902), .B(n55901), .Z(n52630) );
  NOR U72853 ( .A(n52628), .B(n52627), .Z(n52629) );
  NOR U72854 ( .A(n52630), .B(n52629), .Z(n52631) );
  NOR U72855 ( .A(n62978), .B(n52631), .Z(n55899) );
  XOR U72856 ( .A(n52632), .B(n55899), .Z(n57824) );
  XOR U72857 ( .A(n52633), .B(n57824), .Z(n55896) );
  XOR U72858 ( .A(n52634), .B(n55896), .Z(n55894) );
  XOR U72859 ( .A(n52635), .B(n55894), .Z(n61068) );
  XOR U72860 ( .A(n55889), .B(n61068), .Z(n55882) );
  XOR U72861 ( .A(n55881), .B(n55882), .Z(n55879) );
  XOR U72862 ( .A(n52636), .B(n55879), .Z(n52650) );
  NOR U72863 ( .A(n52642), .B(n52650), .Z(n52646) );
  IV U72864 ( .A(n52637), .Z(n52639) );
  NOR U72865 ( .A(n52639), .B(n52638), .Z(n52640) );
  IV U72866 ( .A(n52640), .Z(n52647) );
  IV U72867 ( .A(n52650), .Z(n52641) );
  NOR U72868 ( .A(n52647), .B(n52641), .Z(n61047) );
  IV U72869 ( .A(n52642), .Z(n52644) );
  XOR U72870 ( .A(n55878), .B(n55879), .Z(n52643) );
  NOR U72871 ( .A(n52644), .B(n52643), .Z(n61050) );
  NOR U72872 ( .A(n61047), .B(n61050), .Z(n57828) );
  IV U72873 ( .A(n57828), .Z(n52645) );
  NOR U72874 ( .A(n52646), .B(n52645), .Z(n55870) );
  XOR U72875 ( .A(n55869), .B(n55870), .Z(n52652) );
  NOR U72876 ( .A(n55869), .B(n52647), .Z(n52648) );
  IV U72877 ( .A(n52648), .Z(n52649) );
  NOR U72878 ( .A(n52650), .B(n52649), .Z(n52651) );
  NOR U72879 ( .A(n52652), .B(n52651), .Z(n55874) );
  XOR U72880 ( .A(n55873), .B(n55874), .Z(n55859) );
  XOR U72881 ( .A(n52653), .B(n55859), .Z(n57831) );
  XOR U72882 ( .A(n57830), .B(n57831), .Z(n57834) );
  XOR U72883 ( .A(n57833), .B(n57834), .Z(n55857) );
  XOR U72884 ( .A(n52654), .B(n55857), .Z(n55852) );
  XOR U72885 ( .A(n52655), .B(n55852), .Z(n57841) );
  NOR U72886 ( .A(n52662), .B(n57841), .Z(n63034) );
  IV U72887 ( .A(n52656), .Z(n52657) );
  NOR U72888 ( .A(n52658), .B(n52657), .Z(n55844) );
  IV U72889 ( .A(n52659), .Z(n52661) );
  NOR U72890 ( .A(n52661), .B(n52660), .Z(n57843) );
  XOR U72891 ( .A(n57840), .B(n57841), .Z(n57844) );
  XOR U72892 ( .A(n57843), .B(n57844), .Z(n55845) );
  IV U72893 ( .A(n55845), .Z(n52663) );
  XOR U72894 ( .A(n55844), .B(n52663), .Z(n52665) );
  NOR U72895 ( .A(n52663), .B(n52662), .Z(n52664) );
  NOR U72896 ( .A(n52665), .B(n52664), .Z(n52666) );
  NOR U72897 ( .A(n63034), .B(n52666), .Z(n55835) );
  IV U72898 ( .A(n52667), .Z(n52669) );
  NOR U72899 ( .A(n52669), .B(n52668), .Z(n55847) );
  IV U72900 ( .A(n52670), .Z(n52672) );
  NOR U72901 ( .A(n52672), .B(n52671), .Z(n55834) );
  NOR U72902 ( .A(n55847), .B(n55834), .Z(n52673) );
  XOR U72903 ( .A(n55835), .B(n52673), .Z(n55841) );
  XOR U72904 ( .A(n55839), .B(n55841), .Z(n55832) );
  XOR U72905 ( .A(n52674), .B(n55832), .Z(n52675) );
  IV U72906 ( .A(n52675), .Z(n55826) );
  IV U72907 ( .A(n52676), .Z(n55830) );
  NOR U72908 ( .A(n55830), .B(n55825), .Z(n52677) );
  XOR U72909 ( .A(n55826), .B(n52677), .Z(n52678) );
  XOR U72910 ( .A(n52679), .B(n52678), .Z(n60995) );
  XOR U72911 ( .A(n55824), .B(n60995), .Z(n55818) );
  XOR U72912 ( .A(n55819), .B(n55818), .Z(n63051) );
  IV U72913 ( .A(n52680), .Z(n52681) );
  NOR U72914 ( .A(n52681), .B(n63050), .Z(n55820) );
  XOR U72915 ( .A(n63051), .B(n55820), .Z(n55816) );
  IV U72916 ( .A(n52682), .Z(n52683) );
  NOR U72917 ( .A(n52683), .B(n52685), .Z(n55809) );
  IV U72918 ( .A(n52684), .Z(n52686) );
  NOR U72919 ( .A(n52686), .B(n52685), .Z(n55814) );
  NOR U72920 ( .A(n55809), .B(n55814), .Z(n52687) );
  XOR U72921 ( .A(n55816), .B(n52687), .Z(n55807) );
  XOR U72922 ( .A(n52688), .B(n55807), .Z(n55805) );
  XOR U72923 ( .A(n52689), .B(n55805), .Z(n55794) );
  XOR U72924 ( .A(n55795), .B(n55794), .Z(n57861) );
  XOR U72925 ( .A(n52690), .B(n57861), .Z(n52691) );
  IV U72926 ( .A(n52691), .Z(n57859) );
  XOR U72927 ( .A(n57857), .B(n57859), .Z(n57870) );
  XOR U72928 ( .A(n57869), .B(n57870), .Z(n57866) );
  XOR U72929 ( .A(n57865), .B(n57866), .Z(n57883) );
  IV U72930 ( .A(n52692), .Z(n52694) );
  NOR U72931 ( .A(n52694), .B(n52693), .Z(n57872) );
  NOR U72932 ( .A(n52698), .B(n52695), .Z(n57882) );
  NOR U72933 ( .A(n57872), .B(n57882), .Z(n52696) );
  XOR U72934 ( .A(n57883), .B(n52696), .Z(n57879) );
  IV U72935 ( .A(n52697), .Z(n52699) );
  NOR U72936 ( .A(n52699), .B(n52698), .Z(n52700) );
  IV U72937 ( .A(n52700), .Z(n57880) );
  XOR U72938 ( .A(n57879), .B(n57880), .Z(n57886) );
  XOR U72939 ( .A(n57885), .B(n57886), .Z(n57892) );
  IV U72940 ( .A(n52701), .Z(n52702) );
  NOR U72941 ( .A(n52703), .B(n52702), .Z(n57888) );
  IV U72942 ( .A(n52704), .Z(n52706) );
  NOR U72943 ( .A(n52706), .B(n52705), .Z(n57890) );
  NOR U72944 ( .A(n57888), .B(n57890), .Z(n52707) );
  XOR U72945 ( .A(n57892), .B(n52707), .Z(n52708) );
  NOR U72946 ( .A(n52709), .B(n52708), .Z(n55793) );
  IV U72947 ( .A(n52709), .Z(n52711) );
  XOR U72948 ( .A(n57890), .B(n57892), .Z(n52710) );
  NOR U72949 ( .A(n52711), .B(n52710), .Z(n66466) );
  NOR U72950 ( .A(n55793), .B(n66466), .Z(n57901) );
  XOR U72951 ( .A(n52712), .B(n57901), .Z(n57899) );
  XOR U72952 ( .A(n52713), .B(n57899), .Z(n55782) );
  NOR U72953 ( .A(n52715), .B(n52714), .Z(n52716) );
  IV U72954 ( .A(n52716), .Z(n55783) );
  NOR U72955 ( .A(n52717), .B(n55783), .Z(n52718) );
  XOR U72956 ( .A(n55782), .B(n52718), .Z(n55780) );
  XOR U72957 ( .A(n52719), .B(n55780), .Z(n52720) );
  IV U72958 ( .A(n52720), .Z(n57904) );
  XOR U72959 ( .A(n57903), .B(n57904), .Z(n57906) );
  XOR U72960 ( .A(n57907), .B(n57906), .Z(n55770) );
  IV U72961 ( .A(n52721), .Z(n52722) );
  NOR U72962 ( .A(n52723), .B(n52722), .Z(n55774) );
  IV U72963 ( .A(n52724), .Z(n52725) );
  NOR U72964 ( .A(n52727), .B(n52725), .Z(n55769) );
  NOR U72965 ( .A(n55774), .B(n55769), .Z(n52726) );
  XOR U72966 ( .A(n55770), .B(n52726), .Z(n55763) );
  NOR U72967 ( .A(n52728), .B(n52727), .Z(n52729) );
  IV U72968 ( .A(n52729), .Z(n55762) );
  NOR U72969 ( .A(n52730), .B(n55762), .Z(n52731) );
  XOR U72970 ( .A(n55763), .B(n52731), .Z(n57913) );
  XOR U72971 ( .A(n55759), .B(n57913), .Z(n57918) );
  XOR U72972 ( .A(n52732), .B(n57918), .Z(n57914) );
  XOR U72973 ( .A(n57915), .B(n57914), .Z(n55758) );
  NOR U72974 ( .A(n52734), .B(n52733), .Z(n52735) );
  IV U72975 ( .A(n52735), .Z(n52736) );
  NOR U72976 ( .A(n52737), .B(n52736), .Z(n55756) );
  XOR U72977 ( .A(n55758), .B(n55756), .Z(n55752) );
  IV U72978 ( .A(n52738), .Z(n52740) );
  NOR U72979 ( .A(n52740), .B(n52739), .Z(n55754) );
  IV U72980 ( .A(n52741), .Z(n52742) );
  NOR U72981 ( .A(n52742), .B(n52747), .Z(n55751) );
  NOR U72982 ( .A(n55754), .B(n55751), .Z(n52743) );
  XOR U72983 ( .A(n55752), .B(n52743), .Z(n55745) );
  IV U72984 ( .A(n52744), .Z(n52745) );
  NOR U72985 ( .A(n52745), .B(n52747), .Z(n55748) );
  IV U72986 ( .A(n52746), .Z(n52748) );
  NOR U72987 ( .A(n52748), .B(n52747), .Z(n55744) );
  NOR U72988 ( .A(n55748), .B(n55744), .Z(n52749) );
  XOR U72989 ( .A(n55745), .B(n52749), .Z(n55742) );
  IV U72990 ( .A(n52750), .Z(n52757) );
  NOR U72991 ( .A(n52751), .B(n52757), .Z(n55736) );
  NOR U72992 ( .A(n55741), .B(n55736), .Z(n52752) );
  XOR U72993 ( .A(n55742), .B(n52752), .Z(n55732) );
  IV U72994 ( .A(n52753), .Z(n52754) );
  NOR U72995 ( .A(n52755), .B(n52754), .Z(n55738) );
  IV U72996 ( .A(n52756), .Z(n52760) );
  NOR U72997 ( .A(n52758), .B(n52757), .Z(n52759) );
  IV U72998 ( .A(n52759), .Z(n52763) );
  NOR U72999 ( .A(n52760), .B(n52763), .Z(n55733) );
  NOR U73000 ( .A(n55738), .B(n55733), .Z(n52761) );
  XOR U73001 ( .A(n55732), .B(n52761), .Z(n55731) );
  IV U73002 ( .A(n52762), .Z(n52764) );
  NOR U73003 ( .A(n52764), .B(n52763), .Z(n55729) );
  XOR U73004 ( .A(n55731), .B(n55729), .Z(n57926) );
  XOR U73005 ( .A(n55727), .B(n57926), .Z(n57929) );
  IV U73006 ( .A(n57929), .Z(n52771) );
  IV U73007 ( .A(n52765), .Z(n52767) );
  NOR U73008 ( .A(n52767), .B(n52766), .Z(n57925) );
  NOR U73009 ( .A(n52769), .B(n52768), .Z(n57928) );
  NOR U73010 ( .A(n57925), .B(n57928), .Z(n52770) );
  XOR U73011 ( .A(n52771), .B(n52770), .Z(n57938) );
  NOR U73012 ( .A(n52773), .B(n52772), .Z(n52774) );
  XOR U73013 ( .A(n57938), .B(n52774), .Z(n57941) );
  XOR U73014 ( .A(n55722), .B(n57941), .Z(n52775) );
  NOR U73015 ( .A(n52776), .B(n52775), .Z(n66406) );
  IV U73016 ( .A(n52777), .Z(n57943) );
  IV U73017 ( .A(n52778), .Z(n52781) );
  IV U73018 ( .A(n52779), .Z(n52780) );
  NOR U73019 ( .A(n52781), .B(n52780), .Z(n57939) );
  NOR U73020 ( .A(n55722), .B(n57939), .Z(n52782) );
  XOR U73021 ( .A(n57941), .B(n52782), .Z(n52783) );
  IV U73022 ( .A(n52783), .Z(n57942) );
  XOR U73023 ( .A(n57943), .B(n57942), .Z(n52784) );
  NOR U73024 ( .A(n52785), .B(n52784), .Z(n52786) );
  NOR U73025 ( .A(n66406), .B(n52786), .Z(n57947) );
  IV U73026 ( .A(n52787), .Z(n52789) );
  NOR U73027 ( .A(n52789), .B(n52788), .Z(n57946) );
  IV U73028 ( .A(n52790), .Z(n52792) );
  NOR U73029 ( .A(n52792), .B(n52791), .Z(n57949) );
  NOR U73030 ( .A(n57946), .B(n57949), .Z(n52793) );
  XOR U73031 ( .A(n57947), .B(n52793), .Z(n57954) );
  XOR U73032 ( .A(n57952), .B(n57954), .Z(n55721) );
  XOR U73033 ( .A(n52794), .B(n55721), .Z(n55711) );
  NOR U73034 ( .A(n52797), .B(n52795), .Z(n55710) );
  IV U73035 ( .A(n52796), .Z(n52798) );
  NOR U73036 ( .A(n52798), .B(n52797), .Z(n55713) );
  NOR U73037 ( .A(n55710), .B(n55713), .Z(n52799) );
  XOR U73038 ( .A(n55711), .B(n52799), .Z(n55709) );
  XOR U73039 ( .A(n52800), .B(n55709), .Z(n52801) );
  IV U73040 ( .A(n52801), .Z(n55703) );
  XOR U73041 ( .A(n55702), .B(n55703), .Z(n57959) );
  XOR U73042 ( .A(n57958), .B(n57959), .Z(n57963) );
  IV U73043 ( .A(n52802), .Z(n52804) );
  NOR U73044 ( .A(n52804), .B(n52803), .Z(n57961) );
  XOR U73045 ( .A(n57963), .B(n57961), .Z(n55697) );
  XOR U73046 ( .A(n55696), .B(n55697), .Z(n55701) );
  IV U73047 ( .A(n52805), .Z(n52807) );
  NOR U73048 ( .A(n52807), .B(n52806), .Z(n55699) );
  XOR U73049 ( .A(n55701), .B(n55699), .Z(n55691) );
  XOR U73050 ( .A(n55690), .B(n55691), .Z(n55694) );
  XOR U73051 ( .A(n55693), .B(n55694), .Z(n55688) );
  XOR U73052 ( .A(n55687), .B(n55688), .Z(n57970) );
  XOR U73053 ( .A(n57969), .B(n57970), .Z(n57979) );
  XOR U73054 ( .A(n55685), .B(n57979), .Z(n57982) );
  IV U73055 ( .A(n52808), .Z(n52812) );
  NOR U73056 ( .A(n52810), .B(n52809), .Z(n52811) );
  IV U73057 ( .A(n52811), .Z(n52819) );
  NOR U73058 ( .A(n52812), .B(n52819), .Z(n57980) );
  IV U73059 ( .A(n52813), .Z(n52815) );
  NOR U73060 ( .A(n52815), .B(n52814), .Z(n57977) );
  NOR U73061 ( .A(n57980), .B(n57977), .Z(n52816) );
  XOR U73062 ( .A(n57982), .B(n52816), .Z(n52817) );
  IV U73063 ( .A(n52817), .Z(n57985) );
  IV U73064 ( .A(n52818), .Z(n52820) );
  NOR U73065 ( .A(n52820), .B(n52819), .Z(n57983) );
  XOR U73066 ( .A(n57985), .B(n57983), .Z(n55682) );
  XOR U73067 ( .A(n52821), .B(n55682), .Z(n55678) );
  XOR U73068 ( .A(n55677), .B(n55678), .Z(n57993) );
  XOR U73069 ( .A(n57990), .B(n57993), .Z(n55675) );
  NOR U73070 ( .A(n52823), .B(n52822), .Z(n57992) );
  IV U73071 ( .A(n52824), .Z(n52825) );
  NOR U73072 ( .A(n55670), .B(n52825), .Z(n55674) );
  NOR U73073 ( .A(n57992), .B(n55674), .Z(n52826) );
  XOR U73074 ( .A(n55675), .B(n52826), .Z(n55671) );
  XOR U73075 ( .A(n52827), .B(n55671), .Z(n57998) );
  XOR U73076 ( .A(n52828), .B(n57998), .Z(n58004) );
  XOR U73077 ( .A(n58005), .B(n58004), .Z(n58011) );
  IV U73078 ( .A(n52829), .Z(n52831) );
  NOR U73079 ( .A(n52831), .B(n52830), .Z(n58010) );
  IV U73080 ( .A(n52832), .Z(n52834) );
  NOR U73081 ( .A(n52834), .B(n52833), .Z(n58007) );
  NOR U73082 ( .A(n58010), .B(n58007), .Z(n52835) );
  XOR U73083 ( .A(n58011), .B(n52835), .Z(n58013) );
  XOR U73084 ( .A(n58015), .B(n58013), .Z(n55660) );
  XOR U73085 ( .A(n55659), .B(n55660), .Z(n55664) );
  XOR U73086 ( .A(n52836), .B(n55664), .Z(n55651) );
  XOR U73087 ( .A(n52837), .B(n55651), .Z(n55647) );
  XOR U73088 ( .A(n55646), .B(n55647), .Z(n58021) );
  XOR U73089 ( .A(n52838), .B(n58021), .Z(n52844) );
  IV U73090 ( .A(n52844), .Z(n52839) );
  NOR U73091 ( .A(n52840), .B(n52839), .Z(n63268) );
  IV U73092 ( .A(n52841), .Z(n52842) );
  NOR U73093 ( .A(n52843), .B(n52842), .Z(n52845) );
  NOR U73094 ( .A(n52845), .B(n52844), .Z(n52848) );
  IV U73095 ( .A(n52845), .Z(n52847) );
  XOR U73096 ( .A(n55649), .B(n58021), .Z(n52846) );
  NOR U73097 ( .A(n52847), .B(n52846), .Z(n58026) );
  NOR U73098 ( .A(n52848), .B(n58026), .Z(n52853) );
  NOR U73099 ( .A(n52849), .B(n52853), .Z(n52850) );
  NOR U73100 ( .A(n63268), .B(n52850), .Z(n52851) );
  NOR U73101 ( .A(n52852), .B(n52851), .Z(n52856) );
  IV U73102 ( .A(n52852), .Z(n52855) );
  IV U73103 ( .A(n52853), .Z(n52854) );
  NOR U73104 ( .A(n52855), .B(n52854), .Z(n63271) );
  NOR U73105 ( .A(n52856), .B(n63271), .Z(n52857) );
  IV U73106 ( .A(n52857), .Z(n58030) );
  XOR U73107 ( .A(n58029), .B(n58030), .Z(n55640) );
  XOR U73108 ( .A(n52858), .B(n55640), .Z(n58041) );
  XOR U73109 ( .A(n58039), .B(n58041), .Z(n58044) );
  XOR U73110 ( .A(n52859), .B(n58044), .Z(n55630) );
  IV U73111 ( .A(n52860), .Z(n52862) );
  NOR U73112 ( .A(n52862), .B(n52861), .Z(n55633) );
  IV U73113 ( .A(n52863), .Z(n52865) );
  NOR U73114 ( .A(n52865), .B(n52864), .Z(n55631) );
  NOR U73115 ( .A(n55633), .B(n55631), .Z(n52866) );
  XOR U73116 ( .A(n55630), .B(n52866), .Z(n58049) );
  XOR U73117 ( .A(n58047), .B(n58049), .Z(n58051) );
  XOR U73118 ( .A(n58050), .B(n58051), .Z(n60866) );
  XOR U73119 ( .A(n58054), .B(n60866), .Z(n52867) );
  IV U73120 ( .A(n52867), .Z(n58056) );
  IV U73121 ( .A(n52868), .Z(n52869) );
  NOR U73122 ( .A(n52870), .B(n52869), .Z(n58055) );
  IV U73123 ( .A(n52871), .Z(n52873) );
  IV U73124 ( .A(n52872), .Z(n52879) );
  NOR U73125 ( .A(n52873), .B(n52879), .Z(n55628) );
  NOR U73126 ( .A(n58055), .B(n55628), .Z(n52874) );
  XOR U73127 ( .A(n58056), .B(n52874), .Z(n52881) );
  IV U73128 ( .A(n52881), .Z(n52875) );
  NOR U73129 ( .A(n52876), .B(n52875), .Z(n73646) );
  IV U73130 ( .A(n52877), .Z(n52878) );
  NOR U73131 ( .A(n52879), .B(n52878), .Z(n52882) );
  IV U73132 ( .A(n52882), .Z(n52880) );
  NOR U73133 ( .A(n58056), .B(n52880), .Z(n63311) );
  NOR U73134 ( .A(n52882), .B(n52881), .Z(n52883) );
  NOR U73135 ( .A(n63311), .B(n52883), .Z(n52884) );
  NOR U73136 ( .A(n52885), .B(n52884), .Z(n52886) );
  NOR U73137 ( .A(n73646), .B(n52886), .Z(n52887) );
  IV U73138 ( .A(n52887), .Z(n58061) );
  XOR U73139 ( .A(n58060), .B(n58061), .Z(n55626) );
  IV U73140 ( .A(n52888), .Z(n52890) );
  NOR U73141 ( .A(n52890), .B(n52889), .Z(n55622) );
  IV U73142 ( .A(n52891), .Z(n52893) );
  NOR U73143 ( .A(n52893), .B(n52892), .Z(n55624) );
  NOR U73144 ( .A(n55622), .B(n55624), .Z(n52894) );
  XOR U73145 ( .A(n55626), .B(n52894), .Z(n55611) );
  XOR U73146 ( .A(n52895), .B(n55611), .Z(n55608) );
  XOR U73147 ( .A(n52896), .B(n55608), .Z(n55600) );
  XOR U73148 ( .A(n52897), .B(n55600), .Z(n55592) );
  XOR U73149 ( .A(n52898), .B(n55592), .Z(n55587) );
  XOR U73150 ( .A(n55585), .B(n55587), .Z(n55590) );
  XOR U73151 ( .A(n55588), .B(n55590), .Z(n55582) );
  XOR U73152 ( .A(n52899), .B(n55582), .Z(n55577) );
  IV U73153 ( .A(n52900), .Z(n52904) );
  XOR U73154 ( .A(n52902), .B(n52901), .Z(n52903) );
  NOR U73155 ( .A(n52904), .B(n52903), .Z(n52911) );
  IV U73156 ( .A(n52911), .Z(n66260) );
  NOR U73157 ( .A(n55577), .B(n66260), .Z(n63330) );
  IV U73158 ( .A(n52905), .Z(n52906) );
  NOR U73159 ( .A(n52909), .B(n52906), .Z(n55572) );
  IV U73160 ( .A(n52907), .Z(n52908) );
  NOR U73161 ( .A(n52909), .B(n52908), .Z(n55575) );
  XOR U73162 ( .A(n55577), .B(n55575), .Z(n55573) );
  XOR U73163 ( .A(n55572), .B(n55573), .Z(n66265) );
  IV U73164 ( .A(n66265), .Z(n52910) );
  NOR U73165 ( .A(n52911), .B(n52910), .Z(n52912) );
  NOR U73166 ( .A(n63330), .B(n52912), .Z(n55569) );
  IV U73167 ( .A(n52913), .Z(n52918) );
  IV U73168 ( .A(n52914), .Z(n52915) );
  NOR U73169 ( .A(n52916), .B(n52915), .Z(n52917) );
  IV U73170 ( .A(n52917), .Z(n52921) );
  NOR U73171 ( .A(n52918), .B(n52921), .Z(n52919) );
  IV U73172 ( .A(n52919), .Z(n55570) );
  XOR U73173 ( .A(n55569), .B(n55570), .Z(n58077) );
  IV U73174 ( .A(n52920), .Z(n52922) );
  NOR U73175 ( .A(n52922), .B(n52921), .Z(n58075) );
  XOR U73176 ( .A(n58077), .B(n58075), .Z(n58079) );
  IV U73177 ( .A(n52923), .Z(n52924) );
  NOR U73178 ( .A(n52931), .B(n52924), .Z(n58078) );
  IV U73179 ( .A(n52925), .Z(n52927) );
  NOR U73180 ( .A(n52927), .B(n52926), .Z(n55567) );
  NOR U73181 ( .A(n58078), .B(n55567), .Z(n52928) );
  XOR U73182 ( .A(n58079), .B(n52928), .Z(n55561) );
  IV U73183 ( .A(n52929), .Z(n52930) );
  NOR U73184 ( .A(n52931), .B(n52930), .Z(n55562) );
  NOR U73185 ( .A(n55564), .B(n55562), .Z(n52932) );
  XOR U73186 ( .A(n55561), .B(n52932), .Z(n58084) );
  IV U73187 ( .A(n52933), .Z(n52934) );
  NOR U73188 ( .A(n52935), .B(n52934), .Z(n58082) );
  XOR U73189 ( .A(n58084), .B(n58082), .Z(n58086) );
  XOR U73190 ( .A(n58085), .B(n58086), .Z(n55559) );
  XOR U73191 ( .A(n55553), .B(n55559), .Z(n52936) );
  XOR U73192 ( .A(n52937), .B(n52936), .Z(n55547) );
  NOR U73193 ( .A(n52939), .B(n52938), .Z(n52940) );
  IV U73194 ( .A(n52940), .Z(n55548) );
  XOR U73195 ( .A(n55547), .B(n55548), .Z(n55551) );
  NOR U73196 ( .A(n52942), .B(n52941), .Z(n55544) );
  NOR U73197 ( .A(n55550), .B(n55544), .Z(n52943) );
  XOR U73198 ( .A(n55551), .B(n52943), .Z(n52944) );
  IV U73199 ( .A(n52944), .Z(n58093) );
  IV U73200 ( .A(n52945), .Z(n52947) );
  NOR U73201 ( .A(n52947), .B(n52946), .Z(n58091) );
  XOR U73202 ( .A(n58093), .B(n58091), .Z(n58096) );
  XOR U73203 ( .A(n58094), .B(n58096), .Z(n55540) );
  XOR U73204 ( .A(n55538), .B(n55540), .Z(n55543) );
  XOR U73205 ( .A(n55541), .B(n55543), .Z(n58100) );
  XOR U73206 ( .A(n58098), .B(n58100), .Z(n58103) );
  XOR U73207 ( .A(n52948), .B(n58103), .Z(n55530) );
  XOR U73208 ( .A(n52949), .B(n55530), .Z(n55526) );
  XOR U73209 ( .A(n55524), .B(n55526), .Z(n55529) );
  XOR U73210 ( .A(n55527), .B(n55529), .Z(n58106) );
  XOR U73211 ( .A(n58105), .B(n58106), .Z(n58109) );
  XOR U73212 ( .A(n52950), .B(n58109), .Z(n55516) );
  IV U73213 ( .A(n52951), .Z(n52952) );
  NOR U73214 ( .A(n52953), .B(n52952), .Z(n52954) );
  IV U73215 ( .A(n52954), .Z(n55517) );
  XOR U73216 ( .A(n55516), .B(n55517), .Z(n55520) );
  IV U73217 ( .A(n52955), .Z(n52956) );
  NOR U73218 ( .A(n52957), .B(n52956), .Z(n55519) );
  IV U73219 ( .A(n52958), .Z(n52960) );
  NOR U73220 ( .A(n52960), .B(n52959), .Z(n55513) );
  NOR U73221 ( .A(n55519), .B(n55513), .Z(n52961) );
  XOR U73222 ( .A(n55520), .B(n52961), .Z(n58111) );
  XOR U73223 ( .A(n58112), .B(n58111), .Z(n58115) );
  XOR U73224 ( .A(n58114), .B(n58115), .Z(n58119) );
  XOR U73225 ( .A(n58118), .B(n58119), .Z(n58125) );
  XOR U73226 ( .A(n52962), .B(n58125), .Z(n58128) );
  XOR U73227 ( .A(n52963), .B(n58128), .Z(n55511) );
  XOR U73228 ( .A(n55510), .B(n55511), .Z(n55508) );
  XOR U73229 ( .A(n52964), .B(n55508), .Z(n55493) );
  XOR U73230 ( .A(n52965), .B(n55493), .Z(n55497) );
  XOR U73231 ( .A(n55496), .B(n55497), .Z(n55491) );
  XOR U73232 ( .A(n52966), .B(n55491), .Z(n55483) );
  IV U73233 ( .A(n52967), .Z(n52968) );
  NOR U73234 ( .A(n52969), .B(n52968), .Z(n55487) );
  IV U73235 ( .A(n52970), .Z(n52971) );
  NOR U73236 ( .A(n52972), .B(n52971), .Z(n55482) );
  NOR U73237 ( .A(n55487), .B(n55482), .Z(n52973) );
  XOR U73238 ( .A(n55483), .B(n52973), .Z(n55478) );
  IV U73239 ( .A(n52974), .Z(n52976) );
  NOR U73240 ( .A(n52976), .B(n52975), .Z(n55476) );
  XOR U73241 ( .A(n55478), .B(n55476), .Z(n55480) );
  XOR U73242 ( .A(n55479), .B(n55480), .Z(n63444) );
  XOR U73243 ( .A(n55475), .B(n63444), .Z(n58146) );
  IV U73244 ( .A(n52977), .Z(n52978) );
  NOR U73245 ( .A(n52979), .B(n52978), .Z(n68814) );
  IV U73246 ( .A(n52980), .Z(n52981) );
  NOR U73247 ( .A(n52982), .B(n52981), .Z(n66186) );
  NOR U73248 ( .A(n68814), .B(n66186), .Z(n58147) );
  XOR U73249 ( .A(n58146), .B(n58147), .Z(n58150) );
  XOR U73250 ( .A(n58148), .B(n58150), .Z(n55472) );
  XOR U73251 ( .A(n55471), .B(n55472), .Z(n58155) );
  XOR U73252 ( .A(n58153), .B(n58155), .Z(n55470) );
  XOR U73253 ( .A(n55468), .B(n55470), .Z(n58161) );
  XOR U73254 ( .A(n58159), .B(n58161), .Z(n58163) );
  XOR U73255 ( .A(n58164), .B(n58163), .Z(n52985) );
  NOR U73256 ( .A(n52983), .B(n52985), .Z(n52998) );
  IV U73257 ( .A(n52984), .Z(n52992) );
  IV U73258 ( .A(n52985), .Z(n52986) );
  NOR U73259 ( .A(n52987), .B(n52986), .Z(n52988) );
  IV U73260 ( .A(n52988), .Z(n52989) );
  NOR U73261 ( .A(n52990), .B(n52989), .Z(n52991) );
  IV U73262 ( .A(n52991), .Z(n52994) );
  NOR U73263 ( .A(n52992), .B(n52994), .Z(n60762) );
  IV U73264 ( .A(n52993), .Z(n52995) );
  NOR U73265 ( .A(n52995), .B(n52994), .Z(n60760) );
  NOR U73266 ( .A(n60762), .B(n60760), .Z(n52996) );
  IV U73267 ( .A(n52996), .Z(n52997) );
  NOR U73268 ( .A(n52998), .B(n52997), .Z(n58166) );
  XOR U73269 ( .A(n58168), .B(n58166), .Z(n55466) );
  XOR U73270 ( .A(n55464), .B(n55466), .Z(n58177) );
  XOR U73271 ( .A(n52999), .B(n58177), .Z(n53000) );
  IV U73272 ( .A(n53000), .Z(n58187) );
  XOR U73273 ( .A(n53001), .B(n58187), .Z(n58196) );
  XOR U73274 ( .A(n53002), .B(n58196), .Z(n58189) );
  XOR U73275 ( .A(n53003), .B(n58189), .Z(n58210) );
  XOR U73276 ( .A(n53004), .B(n58210), .Z(n58212) );
  XOR U73277 ( .A(n58211), .B(n58212), .Z(n58215) );
  XOR U73278 ( .A(n58214), .B(n58215), .Z(n53005) );
  XOR U73279 ( .A(n53006), .B(n53005), .Z(n55453) );
  XOR U73280 ( .A(n55450), .B(n55453), .Z(n58224) );
  XOR U73281 ( .A(n53007), .B(n58224), .Z(n53009) );
  XOR U73282 ( .A(n53010), .B(n53009), .Z(n55448) );
  NOR U73283 ( .A(n53008), .B(n55448), .Z(n66153) );
  IV U73284 ( .A(n53009), .Z(n58230) );
  IV U73285 ( .A(n53010), .Z(n53014) );
  IV U73286 ( .A(n53011), .Z(n53012) );
  NOR U73287 ( .A(n53013), .B(n53012), .Z(n55447) );
  NOR U73288 ( .A(n53014), .B(n55447), .Z(n53015) );
  XOR U73289 ( .A(n58230), .B(n53015), .Z(n53016) );
  NOR U73290 ( .A(n53017), .B(n53016), .Z(n53018) );
  NOR U73291 ( .A(n66153), .B(n53018), .Z(n53019) );
  IV U73292 ( .A(n53019), .Z(n55444) );
  XOR U73293 ( .A(n53020), .B(n55444), .Z(n55437) );
  XOR U73294 ( .A(n55436), .B(n55437), .Z(n55440) );
  XOR U73295 ( .A(n55439), .B(n55440), .Z(n58237) );
  XOR U73296 ( .A(n53021), .B(n58237), .Z(n58246) );
  XOR U73297 ( .A(n58247), .B(n58246), .Z(n55426) );
  XOR U73298 ( .A(n55424), .B(n55426), .Z(n58245) );
  XOR U73299 ( .A(n58243), .B(n58245), .Z(n58254) );
  XOR U73300 ( .A(n58253), .B(n58254), .Z(n58260) );
  XOR U73301 ( .A(n53022), .B(n58260), .Z(n55422) );
  XOR U73302 ( .A(n55420), .B(n55422), .Z(n55413) );
  XOR U73303 ( .A(n53023), .B(n55413), .Z(n58273) );
  IV U73304 ( .A(n53024), .Z(n53027) );
  IV U73305 ( .A(n53025), .Z(n53026) );
  NOR U73306 ( .A(n53027), .B(n53026), .Z(n58272) );
  NOR U73307 ( .A(n55407), .B(n58272), .Z(n53028) );
  XOR U73308 ( .A(n58273), .B(n53028), .Z(n58270) );
  XOR U73309 ( .A(n58271), .B(n58270), .Z(n55405) );
  XOR U73310 ( .A(n53029), .B(n55405), .Z(n55395) );
  XOR U73311 ( .A(n53030), .B(n55395), .Z(n55399) );
  XOR U73312 ( .A(n53031), .B(n55399), .Z(n53032) );
  IV U73313 ( .A(n53032), .Z(n55387) );
  XOR U73314 ( .A(n55385), .B(n55387), .Z(n58283) );
  NOR U73315 ( .A(n53033), .B(n55388), .Z(n53034) );
  NOR U73316 ( .A(n53034), .B(n55389), .Z(n53035) );
  XOR U73317 ( .A(n58283), .B(n53035), .Z(n58286) );
  IV U73318 ( .A(n53036), .Z(n53039) );
  IV U73319 ( .A(n53037), .Z(n53038) );
  NOR U73320 ( .A(n53039), .B(n53038), .Z(n55383) );
  IV U73321 ( .A(n53040), .Z(n53041) );
  NOR U73322 ( .A(n53041), .B(n53046), .Z(n58285) );
  NOR U73323 ( .A(n55383), .B(n58285), .Z(n53042) );
  XOR U73324 ( .A(n58286), .B(n53042), .Z(n55380) );
  IV U73325 ( .A(n53043), .Z(n53044) );
  NOR U73326 ( .A(n53044), .B(n53046), .Z(n55381) );
  IV U73327 ( .A(n53045), .Z(n53047) );
  NOR U73328 ( .A(n53047), .B(n53046), .Z(n58288) );
  NOR U73329 ( .A(n55381), .B(n58288), .Z(n53048) );
  XOR U73330 ( .A(n55380), .B(n53048), .Z(n60660) );
  IV U73331 ( .A(n60660), .Z(n53053) );
  IV U73332 ( .A(n53049), .Z(n53052) );
  IV U73333 ( .A(n53050), .Z(n53051) );
  NOR U73334 ( .A(n53052), .B(n53051), .Z(n60659) );
  NOR U73335 ( .A(n60666), .B(n60659), .Z(n58291) );
  XOR U73336 ( .A(n53053), .B(n58291), .Z(n58293) );
  XOR U73337 ( .A(n58292), .B(n58293), .Z(n58299) );
  XOR U73338 ( .A(n53054), .B(n58299), .Z(n58308) );
  NOR U73339 ( .A(n53061), .B(n58308), .Z(n63576) );
  IV U73340 ( .A(n53055), .Z(n53056) );
  NOR U73341 ( .A(n53057), .B(n53056), .Z(n55377) );
  IV U73342 ( .A(n53058), .Z(n53060) );
  NOR U73343 ( .A(n53060), .B(n53059), .Z(n58306) );
  XOR U73344 ( .A(n58308), .B(n58306), .Z(n55378) );
  IV U73345 ( .A(n55378), .Z(n53062) );
  XOR U73346 ( .A(n55377), .B(n53062), .Z(n53064) );
  NOR U73347 ( .A(n53062), .B(n53061), .Z(n53063) );
  NOR U73348 ( .A(n53064), .B(n53063), .Z(n53065) );
  NOR U73349 ( .A(n63576), .B(n53065), .Z(n55372) );
  XOR U73350 ( .A(n53066), .B(n55372), .Z(n55366) );
  XOR U73351 ( .A(n55364), .B(n55366), .Z(n55369) );
  IV U73352 ( .A(n53067), .Z(n53069) );
  NOR U73353 ( .A(n53069), .B(n53068), .Z(n55362) );
  IV U73354 ( .A(n53070), .Z(n53071) );
  NOR U73355 ( .A(n53072), .B(n53071), .Z(n53073) );
  IV U73356 ( .A(n53073), .Z(n53074) );
  NOR U73357 ( .A(n53075), .B(n53074), .Z(n55367) );
  NOR U73358 ( .A(n55362), .B(n55367), .Z(n53076) );
  XOR U73359 ( .A(n55369), .B(n53076), .Z(n53077) );
  IV U73360 ( .A(n53077), .Z(n55361) );
  XOR U73361 ( .A(n55357), .B(n55361), .Z(n53078) );
  NOR U73362 ( .A(n53079), .B(n53078), .Z(n66073) );
  IV U73363 ( .A(n53080), .Z(n53081) );
  NOR U73364 ( .A(n53082), .B(n53081), .Z(n55359) );
  NOR U73365 ( .A(n55357), .B(n55359), .Z(n53083) );
  XOR U73366 ( .A(n55361), .B(n53083), .Z(n53084) );
  NOR U73367 ( .A(n53085), .B(n53084), .Z(n53086) );
  NOR U73368 ( .A(n66073), .B(n53086), .Z(n55354) );
  XOR U73369 ( .A(n55356), .B(n55354), .Z(n58316) );
  IV U73370 ( .A(n53087), .Z(n53094) );
  NOR U73371 ( .A(n53088), .B(n53094), .Z(n58312) );
  IV U73372 ( .A(n53089), .Z(n53090) );
  NOR U73373 ( .A(n53090), .B(n53094), .Z(n58314) );
  NOR U73374 ( .A(n58312), .B(n58314), .Z(n53091) );
  XOR U73375 ( .A(n58316), .B(n53091), .Z(n53092) );
  IV U73376 ( .A(n53092), .Z(n55350) );
  IV U73377 ( .A(n53093), .Z(n53095) );
  NOR U73378 ( .A(n53095), .B(n53094), .Z(n55348) );
  XOR U73379 ( .A(n55350), .B(n55348), .Z(n55353) );
  XOR U73380 ( .A(n55351), .B(n55353), .Z(n55343) );
  XOR U73381 ( .A(n55342), .B(n55343), .Z(n55346) );
  NOR U73382 ( .A(n53101), .B(n55346), .Z(n53096) );
  IV U73383 ( .A(n53096), .Z(n55338) );
  NOR U73384 ( .A(n53102), .B(n55338), .Z(n60634) );
  NOR U73385 ( .A(n53097), .B(n55345), .Z(n53098) );
  NOR U73386 ( .A(n53099), .B(n53098), .Z(n53100) );
  XOR U73387 ( .A(n55346), .B(n53100), .Z(n53107) );
  IV U73388 ( .A(n53107), .Z(n53104) );
  NOR U73389 ( .A(n53102), .B(n53101), .Z(n53103) );
  NOR U73390 ( .A(n53104), .B(n53103), .Z(n53105) );
  NOR U73391 ( .A(n60634), .B(n53105), .Z(n58322) );
  NOR U73392 ( .A(n53106), .B(n58322), .Z(n53109) );
  IV U73393 ( .A(n53106), .Z(n53108) );
  NOR U73394 ( .A(n53108), .B(n53107), .Z(n63624) );
  NOR U73395 ( .A(n53109), .B(n63624), .Z(n55334) );
  XOR U73396 ( .A(n53110), .B(n55334), .Z(n55332) );
  XOR U73397 ( .A(n55330), .B(n55332), .Z(n55324) );
  XOR U73398 ( .A(n55325), .B(n55324), .Z(n55326) );
  IV U73399 ( .A(n53111), .Z(n53114) );
  NOR U73400 ( .A(n53117), .B(n53112), .Z(n53113) );
  IV U73401 ( .A(n53113), .Z(n53120) );
  NOR U73402 ( .A(n53114), .B(n53120), .Z(n58327) );
  IV U73403 ( .A(n53115), .Z(n53116) );
  NOR U73404 ( .A(n53117), .B(n53116), .Z(n55327) );
  NOR U73405 ( .A(n58327), .B(n55327), .Z(n53118) );
  XOR U73406 ( .A(n55326), .B(n53118), .Z(n58331) );
  IV U73407 ( .A(n53119), .Z(n53121) );
  NOR U73408 ( .A(n53121), .B(n53120), .Z(n53122) );
  IV U73409 ( .A(n53122), .Z(n58330) );
  XOR U73410 ( .A(n58331), .B(n58330), .Z(n53125) );
  NOR U73411 ( .A(n53123), .B(n53125), .Z(n53137) );
  IV U73412 ( .A(n53124), .Z(n53129) );
  IV U73413 ( .A(n53125), .Z(n53126) );
  NOR U73414 ( .A(n53131), .B(n53126), .Z(n53127) );
  IV U73415 ( .A(n53127), .Z(n53128) );
  NOR U73416 ( .A(n53129), .B(n53128), .Z(n68946) );
  IV U73417 ( .A(n53130), .Z(n53134) );
  NOR U73418 ( .A(n58331), .B(n53131), .Z(n53132) );
  IV U73419 ( .A(n53132), .Z(n53133) );
  NOR U73420 ( .A(n53134), .B(n53133), .Z(n63646) );
  NOR U73421 ( .A(n68946), .B(n63646), .Z(n53135) );
  IV U73422 ( .A(n53135), .Z(n53136) );
  NOR U73423 ( .A(n53137), .B(n53136), .Z(n55322) );
  NOR U73424 ( .A(n53139), .B(n53138), .Z(n55321) );
  IV U73425 ( .A(n53140), .Z(n53141) );
  NOR U73426 ( .A(n53144), .B(n53141), .Z(n58333) );
  NOR U73427 ( .A(n55321), .B(n58333), .Z(n53142) );
  XOR U73428 ( .A(n55322), .B(n53142), .Z(n58340) );
  IV U73429 ( .A(n53143), .Z(n53145) );
  NOR U73430 ( .A(n53145), .B(n53144), .Z(n58336) );
  NOR U73431 ( .A(n53147), .B(n53146), .Z(n58338) );
  NOR U73432 ( .A(n58336), .B(n58338), .Z(n53148) );
  XOR U73433 ( .A(n58340), .B(n53148), .Z(n55311) );
  IV U73434 ( .A(n53149), .Z(n53150) );
  NOR U73435 ( .A(n53150), .B(n55312), .Z(n53151) );
  NOR U73436 ( .A(n58341), .B(n53151), .Z(n53152) );
  XOR U73437 ( .A(n55311), .B(n53152), .Z(n55309) );
  XOR U73438 ( .A(n55307), .B(n55309), .Z(n55302) );
  XOR U73439 ( .A(n55301), .B(n55302), .Z(n55297) );
  XOR U73440 ( .A(n53153), .B(n55297), .Z(n58351) );
  XOR U73441 ( .A(n58350), .B(n58351), .Z(n55294) );
  XOR U73442 ( .A(n55292), .B(n55294), .Z(n58349) );
  NOR U73443 ( .A(n53154), .B(n58349), .Z(n63679) );
  IV U73444 ( .A(n53155), .Z(n53156) );
  NOR U73445 ( .A(n53159), .B(n53156), .Z(n58359) );
  IV U73446 ( .A(n53157), .Z(n53158) );
  NOR U73447 ( .A(n53159), .B(n53158), .Z(n58347) );
  XOR U73448 ( .A(n58349), .B(n58347), .Z(n58360) );
  XOR U73449 ( .A(n58359), .B(n58360), .Z(n55286) );
  IV U73450 ( .A(n55286), .Z(n53160) );
  NOR U73451 ( .A(n53161), .B(n53160), .Z(n53162) );
  NOR U73452 ( .A(n63679), .B(n53162), .Z(n55288) );
  IV U73453 ( .A(n53165), .Z(n53163) );
  NOR U73454 ( .A(n53163), .B(n53172), .Z(n55287) );
  IV U73455 ( .A(n53164), .Z(n53167) );
  XOR U73456 ( .A(n53165), .B(n53172), .Z(n53166) );
  NOR U73457 ( .A(n53167), .B(n53166), .Z(n55284) );
  NOR U73458 ( .A(n55287), .B(n55284), .Z(n53168) );
  XOR U73459 ( .A(n55288), .B(n53168), .Z(n58365) );
  NOR U73460 ( .A(n53170), .B(n53169), .Z(n58363) );
  IV U73461 ( .A(n53171), .Z(n53173) );
  NOR U73462 ( .A(n53173), .B(n53172), .Z(n55282) );
  NOR U73463 ( .A(n58363), .B(n55282), .Z(n53174) );
  XOR U73464 ( .A(n58365), .B(n53174), .Z(n55280) );
  IV U73465 ( .A(n53175), .Z(n53177) );
  IV U73466 ( .A(n53176), .Z(n53186) );
  NOR U73467 ( .A(n53177), .B(n53186), .Z(n58371) );
  IV U73468 ( .A(n53178), .Z(n53179) );
  NOR U73469 ( .A(n53180), .B(n53179), .Z(n55279) );
  NOR U73470 ( .A(n55279), .B(n58366), .Z(n53181) );
  IV U73471 ( .A(n53181), .Z(n53182) );
  NOR U73472 ( .A(n58371), .B(n53182), .Z(n53183) );
  XOR U73473 ( .A(n55280), .B(n53183), .Z(n58370) );
  IV U73474 ( .A(n53184), .Z(n53185) );
  NOR U73475 ( .A(n53186), .B(n53185), .Z(n58368) );
  IV U73476 ( .A(n53187), .Z(n53188) );
  NOR U73477 ( .A(n53192), .B(n53188), .Z(n55277) );
  NOR U73478 ( .A(n58368), .B(n55277), .Z(n53189) );
  XOR U73479 ( .A(n58370), .B(n53189), .Z(n55274) );
  IV U73480 ( .A(n53190), .Z(n53191) );
  NOR U73481 ( .A(n53192), .B(n53191), .Z(n53205) );
  IV U73482 ( .A(n53205), .Z(n55275) );
  XOR U73483 ( .A(n55274), .B(n55275), .Z(n53203) );
  IV U73484 ( .A(n53203), .Z(n53201) );
  IV U73485 ( .A(n53193), .Z(n53195) );
  NOR U73486 ( .A(n53195), .B(n53194), .Z(n53206) );
  IV U73487 ( .A(n53196), .Z(n53198) );
  NOR U73488 ( .A(n53198), .B(n53197), .Z(n53202) );
  NOR U73489 ( .A(n53206), .B(n53202), .Z(n53199) );
  IV U73490 ( .A(n53199), .Z(n53200) );
  NOR U73491 ( .A(n53201), .B(n53200), .Z(n53210) );
  IV U73492 ( .A(n53202), .Z(n53204) );
  NOR U73493 ( .A(n53204), .B(n53203), .Z(n65985) );
  NOR U73494 ( .A(n55274), .B(n53205), .Z(n53208) );
  IV U73495 ( .A(n53206), .Z(n53207) );
  NOR U73496 ( .A(n53208), .B(n53207), .Z(n65990) );
  NOR U73497 ( .A(n65985), .B(n65990), .Z(n63698) );
  IV U73498 ( .A(n63698), .Z(n53209) );
  NOR U73499 ( .A(n53210), .B(n53209), .Z(n53211) );
  IV U73500 ( .A(n53211), .Z(n55272) );
  XOR U73501 ( .A(n53212), .B(n55272), .Z(n58388) );
  IV U73502 ( .A(n53213), .Z(n53214) );
  NOR U73503 ( .A(n53215), .B(n53214), .Z(n58382) );
  IV U73504 ( .A(n53216), .Z(n53220) );
  NOR U73505 ( .A(n53217), .B(n55265), .Z(n53218) );
  IV U73506 ( .A(n53218), .Z(n53219) );
  NOR U73507 ( .A(n53220), .B(n53219), .Z(n58387) );
  NOR U73508 ( .A(n58382), .B(n58387), .Z(n53221) );
  XOR U73509 ( .A(n58388), .B(n53221), .Z(n58378) );
  XOR U73510 ( .A(n53222), .B(n58378), .Z(n58395) );
  XOR U73511 ( .A(n55260), .B(n58395), .Z(n58408) );
  XOR U73512 ( .A(n53223), .B(n58408), .Z(n58409) );
  XOR U73513 ( .A(n53224), .B(n58409), .Z(n58417) );
  XOR U73514 ( .A(n58415), .B(n58417), .Z(n60563) );
  XOR U73515 ( .A(n53225), .B(n60563), .Z(n55256) );
  XOR U73516 ( .A(n53226), .B(n55256), .Z(n58427) );
  IV U73517 ( .A(n53227), .Z(n53229) );
  NOR U73518 ( .A(n53229), .B(n53228), .Z(n55255) );
  IV U73519 ( .A(n53230), .Z(n53232) );
  NOR U73520 ( .A(n53232), .B(n53231), .Z(n58426) );
  NOR U73521 ( .A(n55255), .B(n58426), .Z(n53233) );
  XOR U73522 ( .A(n58427), .B(n53233), .Z(n58429) );
  IV U73523 ( .A(n53234), .Z(n53238) );
  NOR U73524 ( .A(n53235), .B(n55241), .Z(n53236) );
  IV U73525 ( .A(n53236), .Z(n53237) );
  NOR U73526 ( .A(n53238), .B(n53237), .Z(n53239) );
  IV U73527 ( .A(n53239), .Z(n58430) );
  XOR U73528 ( .A(n58429), .B(n58430), .Z(n58434) );
  XOR U73529 ( .A(n58432), .B(n58434), .Z(n55240) );
  XOR U73530 ( .A(n53240), .B(n55240), .Z(n55245) );
  XOR U73531 ( .A(n53241), .B(n55245), .Z(n53242) );
  IV U73532 ( .A(n53242), .Z(n55236) );
  XOR U73533 ( .A(n55234), .B(n55236), .Z(n58442) );
  XOR U73534 ( .A(n58441), .B(n58442), .Z(n55232) );
  XOR U73535 ( .A(n55231), .B(n55232), .Z(n58454) );
  IV U73536 ( .A(n53243), .Z(n53245) );
  IV U73537 ( .A(n53244), .Z(n53249) );
  NOR U73538 ( .A(n53245), .B(n53249), .Z(n55229) );
  NOR U73539 ( .A(n58453), .B(n55229), .Z(n53246) );
  XOR U73540 ( .A(n58454), .B(n53246), .Z(n53247) );
  IV U73541 ( .A(n53247), .Z(n58464) );
  IV U73542 ( .A(n53248), .Z(n53250) );
  NOR U73543 ( .A(n53250), .B(n53249), .Z(n58462) );
  NOR U73544 ( .A(n53252), .B(n53251), .Z(n58460) );
  NOR U73545 ( .A(n58462), .B(n58460), .Z(n53253) );
  XOR U73546 ( .A(n58464), .B(n53253), .Z(n55227) );
  IV U73547 ( .A(n53254), .Z(n53255) );
  NOR U73548 ( .A(n53258), .B(n53255), .Z(n55226) );
  IV U73549 ( .A(n53256), .Z(n53257) );
  NOR U73550 ( .A(n53258), .B(n53257), .Z(n58456) );
  NOR U73551 ( .A(n55226), .B(n58456), .Z(n53259) );
  XOR U73552 ( .A(n55227), .B(n53259), .Z(n58473) );
  XOR U73553 ( .A(n58471), .B(n58473), .Z(n58478) );
  XOR U73554 ( .A(n53260), .B(n58478), .Z(n58485) );
  IV U73555 ( .A(n53261), .Z(n58486) );
  NOR U73556 ( .A(n53262), .B(n58486), .Z(n53263) );
  NOR U73557 ( .A(n55214), .B(n53263), .Z(n53264) );
  XOR U73558 ( .A(n58485), .B(n53264), .Z(n55211) );
  IV U73559 ( .A(n53265), .Z(n53267) );
  NOR U73560 ( .A(n53267), .B(n53266), .Z(n58493) );
  IV U73561 ( .A(n53268), .Z(n53269) );
  NOR U73562 ( .A(n53269), .B(n55205), .Z(n55212) );
  NOR U73563 ( .A(n58493), .B(n55212), .Z(n53270) );
  XOR U73564 ( .A(n55211), .B(n53270), .Z(n55204) );
  XOR U73565 ( .A(n53271), .B(n55204), .Z(n58497) );
  XOR U73566 ( .A(n58496), .B(n58497), .Z(n55201) );
  XOR U73567 ( .A(n55200), .B(n55201), .Z(n58506) );
  XOR U73568 ( .A(n58505), .B(n58506), .Z(n65875) );
  IV U73569 ( .A(n65875), .Z(n79544) );
  NOR U73570 ( .A(n58517), .B(n55199), .Z(n53272) );
  XOR U73571 ( .A(n79544), .B(n53272), .Z(n58519) );
  XOR U73572 ( .A(n58518), .B(n58519), .Z(n55194) );
  NOR U73573 ( .A(n53273), .B(n55194), .Z(n60515) );
  XOR U73574 ( .A(n55193), .B(n55194), .Z(n55197) );
  XOR U73575 ( .A(n55196), .B(n55197), .Z(n53282) );
  IV U73576 ( .A(n53282), .Z(n53274) );
  NOR U73577 ( .A(n53275), .B(n53274), .Z(n53276) );
  NOR U73578 ( .A(n60515), .B(n53276), .Z(n53284) );
  IV U73579 ( .A(n53284), .Z(n53277) );
  NOR U73580 ( .A(n53278), .B(n53277), .Z(n60507) );
  IV U73581 ( .A(n53279), .Z(n53281) );
  NOR U73582 ( .A(n53281), .B(n53280), .Z(n53285) );
  IV U73583 ( .A(n53285), .Z(n53283) );
  NOR U73584 ( .A(n53283), .B(n53282), .Z(n60510) );
  NOR U73585 ( .A(n53285), .B(n53284), .Z(n53286) );
  NOR U73586 ( .A(n60510), .B(n53286), .Z(n53287) );
  NOR U73587 ( .A(n53288), .B(n53287), .Z(n53289) );
  NOR U73588 ( .A(n60507), .B(n53289), .Z(n55184) );
  XOR U73589 ( .A(n55185), .B(n55184), .Z(n55182) );
  XOR U73590 ( .A(n55181), .B(n55182), .Z(n58527) );
  XOR U73591 ( .A(n58526), .B(n58527), .Z(n58530) );
  XOR U73592 ( .A(n53290), .B(n58530), .Z(n55168) );
  XOR U73593 ( .A(n55167), .B(n55168), .Z(n55171) );
  XOR U73594 ( .A(n53291), .B(n55171), .Z(n53292) );
  IV U73595 ( .A(n53292), .Z(n55155) );
  IV U73596 ( .A(n53293), .Z(n53294) );
  NOR U73597 ( .A(n55156), .B(n53294), .Z(n53295) );
  XOR U73598 ( .A(n55155), .B(n53295), .Z(n55150) );
  XOR U73599 ( .A(n55151), .B(n55150), .Z(n55146) );
  IV U73600 ( .A(n53296), .Z(n53297) );
  NOR U73601 ( .A(n53298), .B(n53297), .Z(n55152) );
  IV U73602 ( .A(n53299), .Z(n53301) );
  NOR U73603 ( .A(n53301), .B(n53300), .Z(n55147) );
  NOR U73604 ( .A(n55152), .B(n55147), .Z(n53302) );
  XOR U73605 ( .A(n55146), .B(n53302), .Z(n55145) );
  IV U73606 ( .A(n53303), .Z(n53305) );
  NOR U73607 ( .A(n53305), .B(n53304), .Z(n55143) );
  XOR U73608 ( .A(n55145), .B(n55143), .Z(n55137) );
  XOR U73609 ( .A(n55136), .B(n55137), .Z(n55140) );
  XOR U73610 ( .A(n53306), .B(n55140), .Z(n53307) );
  IV U73611 ( .A(n53307), .Z(n55131) );
  XOR U73612 ( .A(n55130), .B(n55131), .Z(n58544) );
  IV U73613 ( .A(n53308), .Z(n55127) );
  IV U73614 ( .A(n53311), .Z(n53309) );
  NOR U73615 ( .A(n55127), .B(n53309), .Z(n58537) );
  NOR U73616 ( .A(n53310), .B(n58539), .Z(n53312) );
  XOR U73617 ( .A(n55127), .B(n53311), .Z(n58545) );
  NOR U73618 ( .A(n53312), .B(n58545), .Z(n53313) );
  NOR U73619 ( .A(n58537), .B(n53313), .Z(n53314) );
  XOR U73620 ( .A(n58544), .B(n53314), .Z(n53315) );
  IV U73621 ( .A(n53315), .Z(n58554) );
  XOR U73622 ( .A(n58550), .B(n58554), .Z(n55123) );
  XOR U73623 ( .A(n53316), .B(n55123), .Z(n55120) );
  XOR U73624 ( .A(n55121), .B(n55120), .Z(n58561) );
  XOR U73625 ( .A(n58556), .B(n58561), .Z(n53317) );
  XOR U73626 ( .A(n53318), .B(n53317), .Z(n58568) );
  IV U73627 ( .A(n53319), .Z(n53321) );
  NOR U73628 ( .A(n53321), .B(n53320), .Z(n58566) );
  XOR U73629 ( .A(n58568), .B(n58566), .Z(n58570) );
  XOR U73630 ( .A(n58569), .B(n58570), .Z(n55119) );
  XOR U73631 ( .A(n55117), .B(n55119), .Z(n58574) );
  XOR U73632 ( .A(n58573), .B(n58574), .Z(n58577) );
  XOR U73633 ( .A(n53322), .B(n58577), .Z(n60444) );
  XOR U73634 ( .A(n58589), .B(n60444), .Z(n55113) );
  XOR U73635 ( .A(n55115), .B(n55113), .Z(n58593) );
  IV U73636 ( .A(n58593), .Z(n53329) );
  IV U73637 ( .A(n53323), .Z(n53327) );
  NOR U73638 ( .A(n53325), .B(n53324), .Z(n53326) );
  IV U73639 ( .A(n53326), .Z(n53331) );
  NOR U73640 ( .A(n53327), .B(n53331), .Z(n55111) );
  NOR U73641 ( .A(n58592), .B(n55111), .Z(n53328) );
  XOR U73642 ( .A(n53329), .B(n53328), .Z(n55110) );
  IV U73643 ( .A(n53330), .Z(n53332) );
  NOR U73644 ( .A(n53332), .B(n53331), .Z(n55108) );
  XOR U73645 ( .A(n55110), .B(n55108), .Z(n55102) );
  XOR U73646 ( .A(n55101), .B(n55102), .Z(n55106) );
  XOR U73647 ( .A(n53333), .B(n55106), .Z(n55094) );
  IV U73648 ( .A(n53334), .Z(n53336) );
  NOR U73649 ( .A(n53336), .B(n53335), .Z(n55096) );
  IV U73650 ( .A(n53337), .Z(n53341) );
  NOR U73651 ( .A(n53339), .B(n53338), .Z(n53340) );
  IV U73652 ( .A(n53340), .Z(n53344) );
  NOR U73653 ( .A(n53341), .B(n53344), .Z(n55093) );
  NOR U73654 ( .A(n55096), .B(n55093), .Z(n53342) );
  XOR U73655 ( .A(n55094), .B(n53342), .Z(n58607) );
  IV U73656 ( .A(n53343), .Z(n53345) );
  NOR U73657 ( .A(n53345), .B(n53344), .Z(n58605) );
  XOR U73658 ( .A(n58607), .B(n58605), .Z(n55091) );
  XOR U73659 ( .A(n55089), .B(n55091), .Z(n58603) );
  XOR U73660 ( .A(n58602), .B(n58603), .Z(n55082) );
  XOR U73661 ( .A(n53346), .B(n55082), .Z(n58622) );
  XOR U73662 ( .A(n58620), .B(n58622), .Z(n55078) );
  XOR U73663 ( .A(n55077), .B(n55078), .Z(n58618) );
  XOR U73664 ( .A(n53347), .B(n58618), .Z(n53348) );
  IV U73665 ( .A(n53348), .Z(n53352) );
  NOR U73666 ( .A(n53349), .B(n53352), .Z(n60420) );
  IV U73667 ( .A(n53350), .Z(n55069) );
  NOR U73668 ( .A(n53351), .B(n55069), .Z(n53353) );
  XOR U73669 ( .A(n53353), .B(n53352), .Z(n53360) );
  IV U73670 ( .A(n53360), .Z(n53354) );
  NOR U73671 ( .A(n53355), .B(n53354), .Z(n53356) );
  NOR U73672 ( .A(n60420), .B(n53356), .Z(n53357) );
  NOR U73673 ( .A(n53358), .B(n53357), .Z(n53361) );
  IV U73674 ( .A(n53358), .Z(n53359) );
  NOR U73675 ( .A(n53360), .B(n53359), .Z(n74225) );
  NOR U73676 ( .A(n53361), .B(n74225), .Z(n55065) );
  IV U73677 ( .A(n53362), .Z(n53364) );
  NOR U73678 ( .A(n53364), .B(n53363), .Z(n58628) );
  IV U73679 ( .A(n53365), .Z(n53367) );
  NOR U73680 ( .A(n53367), .B(n53366), .Z(n55066) );
  NOR U73681 ( .A(n58628), .B(n55066), .Z(n53368) );
  XOR U73682 ( .A(n55065), .B(n53368), .Z(n58634) );
  XOR U73683 ( .A(n58632), .B(n58634), .Z(n58636) );
  NOR U73684 ( .A(n53371), .B(n58636), .Z(n55064) );
  IV U73685 ( .A(n53369), .Z(n53370) );
  NOR U73686 ( .A(n53370), .B(n53377), .Z(n55061) );
  XOR U73687 ( .A(n58635), .B(n58636), .Z(n55062) );
  IV U73688 ( .A(n55062), .Z(n53372) );
  XOR U73689 ( .A(n55061), .B(n53372), .Z(n53374) );
  NOR U73690 ( .A(n53372), .B(n53371), .Z(n53373) );
  NOR U73691 ( .A(n53374), .B(n53373), .Z(n53375) );
  NOR U73692 ( .A(n55064), .B(n53375), .Z(n55055) );
  IV U73693 ( .A(n53376), .Z(n53378) );
  NOR U73694 ( .A(n53378), .B(n53377), .Z(n53379) );
  IV U73695 ( .A(n53379), .Z(n55057) );
  XOR U73696 ( .A(n55055), .B(n55057), .Z(n55059) );
  XOR U73697 ( .A(n55058), .B(n55059), .Z(n58645) );
  XOR U73698 ( .A(n58641), .B(n58645), .Z(n58649) );
  XOR U73699 ( .A(n53380), .B(n58649), .Z(n55053) );
  IV U73700 ( .A(n53381), .Z(n53382) );
  NOR U73701 ( .A(n53383), .B(n53382), .Z(n53384) );
  IV U73702 ( .A(n53384), .Z(n55054) );
  XOR U73703 ( .A(n55053), .B(n55054), .Z(n53385) );
  XOR U73704 ( .A(n53386), .B(n53385), .Z(n55050) );
  XOR U73705 ( .A(n55051), .B(n55050), .Z(n58657) );
  XOR U73706 ( .A(n58656), .B(n58657), .Z(n58660) );
  XOR U73707 ( .A(n58659), .B(n58660), .Z(n58669) );
  XOR U73708 ( .A(n58668), .B(n58669), .Z(n58666) );
  XOR U73709 ( .A(n58664), .B(n58666), .Z(n58673) );
  XOR U73710 ( .A(n53387), .B(n58673), .Z(n53388) );
  IV U73711 ( .A(n53388), .Z(n55047) );
  XOR U73712 ( .A(n55045), .B(n55047), .Z(n55038) );
  NOR U73713 ( .A(n55042), .B(n53389), .Z(n53390) );
  IV U73714 ( .A(n53390), .Z(n53391) );
  NOR U73715 ( .A(n55039), .B(n53391), .Z(n53392) );
  XOR U73716 ( .A(n55038), .B(n53392), .Z(n58683) );
  XOR U73717 ( .A(n58682), .B(n58683), .Z(n58687) );
  IV U73718 ( .A(n53393), .Z(n53395) );
  NOR U73719 ( .A(n53395), .B(n53394), .Z(n55034) );
  IV U73720 ( .A(n53396), .Z(n53398) );
  NOR U73721 ( .A(n53398), .B(n53397), .Z(n58685) );
  NOR U73722 ( .A(n55034), .B(n58685), .Z(n53399) );
  XOR U73723 ( .A(n58687), .B(n53399), .Z(n55029) );
  IV U73724 ( .A(n53400), .Z(n53402) );
  NOR U73725 ( .A(n53402), .B(n53401), .Z(n55031) );
  IV U73726 ( .A(n53403), .Z(n53404) );
  NOR U73727 ( .A(n53405), .B(n53404), .Z(n55028) );
  NOR U73728 ( .A(n55031), .B(n55028), .Z(n53406) );
  XOR U73729 ( .A(n55029), .B(n53406), .Z(n60370) );
  XOR U73730 ( .A(n53407), .B(n60370), .Z(n55026) );
  XOR U73731 ( .A(n55025), .B(n55026), .Z(n58701) );
  XOR U73732 ( .A(n58700), .B(n58701), .Z(n55022) );
  XOR U73733 ( .A(n55021), .B(n55022), .Z(n58698) );
  XOR U73734 ( .A(n58697), .B(n58698), .Z(n58716) );
  XOR U73735 ( .A(n55019), .B(n58716), .Z(n58722) );
  XOR U73736 ( .A(n53408), .B(n58722), .Z(n55016) );
  XOR U73737 ( .A(n53409), .B(n55016), .Z(n55014) );
  XOR U73738 ( .A(n53410), .B(n55014), .Z(n55006) );
  IV U73739 ( .A(n53411), .Z(n53413) );
  NOR U73740 ( .A(n53413), .B(n53412), .Z(n55010) );
  IV U73741 ( .A(n53414), .Z(n53416) );
  NOR U73742 ( .A(n53416), .B(n53415), .Z(n55005) );
  NOR U73743 ( .A(n55010), .B(n55005), .Z(n53417) );
  XOR U73744 ( .A(n55006), .B(n53417), .Z(n55004) );
  XOR U73745 ( .A(n53418), .B(n55004), .Z(n53428) );
  IV U73746 ( .A(n53428), .Z(n53426) );
  IV U73747 ( .A(n53419), .Z(n53436) );
  NOR U73748 ( .A(n53420), .B(n53436), .Z(n53430) );
  IV U73749 ( .A(n53421), .Z(n53423) );
  NOR U73750 ( .A(n53423), .B(n53422), .Z(n53427) );
  NOR U73751 ( .A(n53430), .B(n53427), .Z(n53424) );
  IV U73752 ( .A(n53424), .Z(n53425) );
  NOR U73753 ( .A(n53426), .B(n53425), .Z(n53433) );
  IV U73754 ( .A(n53427), .Z(n53429) );
  NOR U73755 ( .A(n53429), .B(n53428), .Z(n63962) );
  IV U73756 ( .A(n53430), .Z(n53431) );
  NOR U73757 ( .A(n55004), .B(n53431), .Z(n60348) );
  NOR U73758 ( .A(n63962), .B(n60348), .Z(n53432) );
  IV U73759 ( .A(n53432), .Z(n58729) );
  NOR U73760 ( .A(n53433), .B(n58729), .Z(n53434) );
  IV U73761 ( .A(n53434), .Z(n58732) );
  IV U73762 ( .A(n53435), .Z(n53437) );
  NOR U73763 ( .A(n53437), .B(n53436), .Z(n58730) );
  XOR U73764 ( .A(n58732), .B(n58730), .Z(n58735) );
  XOR U73765 ( .A(n53438), .B(n58735), .Z(n60333) );
  IV U73766 ( .A(n60333), .Z(n53439) );
  NOR U73767 ( .A(n53440), .B(n53439), .Z(n53453) );
  IV U73768 ( .A(n53441), .Z(n53447) );
  NOR U73769 ( .A(n53442), .B(n60333), .Z(n53443) );
  IV U73770 ( .A(n53443), .Z(n53444) );
  NOR U73771 ( .A(n53445), .B(n53444), .Z(n53446) );
  IV U73772 ( .A(n53446), .Z(n53449) );
  NOR U73773 ( .A(n53447), .B(n53449), .Z(n60339) );
  IV U73774 ( .A(n53448), .Z(n53450) );
  NOR U73775 ( .A(n53450), .B(n53449), .Z(n63970) );
  NOR U73776 ( .A(n60339), .B(n63970), .Z(n53451) );
  IV U73777 ( .A(n53451), .Z(n53452) );
  NOR U73778 ( .A(n53453), .B(n53452), .Z(n55000) );
  IV U73779 ( .A(n53454), .Z(n60336) );
  NOR U73780 ( .A(n53455), .B(n60336), .Z(n58743) );
  IV U73781 ( .A(n53456), .Z(n53457) );
  NOR U73782 ( .A(n53458), .B(n53457), .Z(n54999) );
  NOR U73783 ( .A(n58743), .B(n54999), .Z(n53459) );
  XOR U73784 ( .A(n55000), .B(n53459), .Z(n54998) );
  XOR U73785 ( .A(n54996), .B(n54998), .Z(n54994) );
  XOR U73786 ( .A(n53460), .B(n54994), .Z(n53461) );
  IV U73787 ( .A(n53461), .Z(n54986) );
  IV U73788 ( .A(n53462), .Z(n54990) );
  NOR U73789 ( .A(n53463), .B(n54990), .Z(n53465) );
  NOR U73790 ( .A(n53470), .B(n54988), .Z(n53464) );
  NOR U73791 ( .A(n53465), .B(n53464), .Z(n53466) );
  XOR U73792 ( .A(n54986), .B(n53466), .Z(n53468) );
  NOR U73793 ( .A(n53467), .B(n53468), .Z(n53477) );
  IV U73794 ( .A(n53468), .Z(n53469) );
  NOR U73795 ( .A(n53470), .B(n53469), .Z(n53471) );
  IV U73796 ( .A(n53471), .Z(n53473) );
  NOR U73797 ( .A(n53472), .B(n53473), .Z(n60317) );
  NOR U73798 ( .A(n53474), .B(n53473), .Z(n60325) );
  NOR U73799 ( .A(n60317), .B(n60325), .Z(n53475) );
  IV U73800 ( .A(n53475), .Z(n53476) );
  NOR U73801 ( .A(n53477), .B(n53476), .Z(n54980) );
  IV U73802 ( .A(n53478), .Z(n53479) );
  NOR U73803 ( .A(n53480), .B(n53479), .Z(n53481) );
  IV U73804 ( .A(n53481), .Z(n54982) );
  XOR U73805 ( .A(n54980), .B(n54982), .Z(n58752) );
  XOR U73806 ( .A(n58750), .B(n58752), .Z(n58755) );
  XOR U73807 ( .A(n58753), .B(n58755), .Z(n58766) );
  XOR U73808 ( .A(n58765), .B(n58766), .Z(n58761) );
  XOR U73809 ( .A(n53482), .B(n58761), .Z(n53483) );
  IV U73810 ( .A(n53483), .Z(n58772) );
  IV U73811 ( .A(n53484), .Z(n53485) );
  NOR U73812 ( .A(n53486), .B(n53485), .Z(n58770) );
  XOR U73813 ( .A(n58772), .B(n58770), .Z(n64002) );
  XOR U73814 ( .A(n58773), .B(n64002), .Z(n58780) );
  XOR U73815 ( .A(n58782), .B(n58780), .Z(n58777) );
  XOR U73816 ( .A(n58776), .B(n58777), .Z(n69271) );
  XOR U73817 ( .A(n53487), .B(n69271), .Z(n54977) );
  XOR U73818 ( .A(n53488), .B(n54977), .Z(n58801) );
  XOR U73819 ( .A(n58799), .B(n58801), .Z(n54974) );
  XOR U73820 ( .A(n54973), .B(n54974), .Z(n58797) );
  XOR U73821 ( .A(n58796), .B(n58797), .Z(n65622) );
  XOR U73822 ( .A(n53489), .B(n65622), .Z(n54967) );
  IV U73823 ( .A(n53490), .Z(n53491) );
  NOR U73824 ( .A(n53497), .B(n53491), .Z(n53492) );
  IV U73825 ( .A(n53492), .Z(n54968) );
  XOR U73826 ( .A(n54967), .B(n54968), .Z(n58810) );
  IV U73827 ( .A(n53493), .Z(n53494) );
  NOR U73828 ( .A(n53494), .B(n53507), .Z(n54964) );
  IV U73829 ( .A(n53495), .Z(n53496) );
  NOR U73830 ( .A(n53497), .B(n53496), .Z(n58808) );
  NOR U73831 ( .A(n54964), .B(n58808), .Z(n53498) );
  XOR U73832 ( .A(n58810), .B(n53498), .Z(n53499) );
  IV U73833 ( .A(n53499), .Z(n58819) );
  IV U73834 ( .A(n53500), .Z(n53505) );
  NOR U73835 ( .A(n53502), .B(n53501), .Z(n53503) );
  IV U73836 ( .A(n53503), .Z(n53504) );
  NOR U73837 ( .A(n53505), .B(n53504), .Z(n58817) );
  XOR U73838 ( .A(n58819), .B(n58817), .Z(n54963) );
  NOR U73839 ( .A(n65602), .B(n54963), .Z(n64040) );
  IV U73840 ( .A(n53506), .Z(n53511) );
  NOR U73841 ( .A(n53508), .B(n53507), .Z(n53509) );
  IV U73842 ( .A(n53509), .Z(n53510) );
  NOR U73843 ( .A(n53511), .B(n53510), .Z(n54961) );
  XOR U73844 ( .A(n54963), .B(n54961), .Z(n65604) );
  IV U73845 ( .A(n65604), .Z(n53512) );
  NOR U73846 ( .A(n53513), .B(n53512), .Z(n53514) );
  NOR U73847 ( .A(n64040), .B(n53514), .Z(n58823) );
  XOR U73848 ( .A(n53515), .B(n58823), .Z(n58832) );
  IV U73849 ( .A(n53516), .Z(n53518) );
  NOR U73850 ( .A(n53518), .B(n53517), .Z(n58830) );
  XOR U73851 ( .A(n58832), .B(n58830), .Z(n58835) );
  XOR U73852 ( .A(n58834), .B(n58835), .Z(n58839) );
  IV U73853 ( .A(n53519), .Z(n53521) );
  NOR U73854 ( .A(n53521), .B(n53520), .Z(n54959) );
  IV U73855 ( .A(n53522), .Z(n53523) );
  NOR U73856 ( .A(n53524), .B(n53523), .Z(n58837) );
  NOR U73857 ( .A(n54959), .B(n58837), .Z(n53525) );
  XOR U73858 ( .A(n58839), .B(n53525), .Z(n53526) );
  IV U73859 ( .A(n53526), .Z(n54958) );
  XOR U73860 ( .A(n54956), .B(n54958), .Z(n53530) );
  IV U73861 ( .A(n53527), .Z(n53528) );
  NOR U73862 ( .A(n53528), .B(n53543), .Z(n53536) );
  IV U73863 ( .A(n53536), .Z(n53529) );
  NOR U73864 ( .A(n53530), .B(n53529), .Z(n60270) );
  IV U73865 ( .A(n53531), .Z(n53533) );
  NOR U73866 ( .A(n53533), .B(n53532), .Z(n54954) );
  NOR U73867 ( .A(n54956), .B(n54954), .Z(n53534) );
  XOR U73868 ( .A(n54958), .B(n53534), .Z(n53535) );
  NOR U73869 ( .A(n53536), .B(n53535), .Z(n53537) );
  NOR U73870 ( .A(n60270), .B(n53537), .Z(n53538) );
  IV U73871 ( .A(n53538), .Z(n54952) );
  XOR U73872 ( .A(n54951), .B(n54952), .Z(n58846) );
  IV U73873 ( .A(n58846), .Z(n53546) );
  IV U73874 ( .A(n53539), .Z(n53540) );
  NOR U73875 ( .A(n53541), .B(n53540), .Z(n58845) );
  IV U73876 ( .A(n53542), .Z(n53544) );
  NOR U73877 ( .A(n53544), .B(n53543), .Z(n54948) );
  NOR U73878 ( .A(n58845), .B(n54948), .Z(n53545) );
  XOR U73879 ( .A(n53546), .B(n53545), .Z(n58844) );
  XOR U73880 ( .A(n58842), .B(n58844), .Z(n53547) );
  XOR U73881 ( .A(n53548), .B(n53547), .Z(n54934) );
  XOR U73882 ( .A(n53549), .B(n54934), .Z(n54931) );
  XOR U73883 ( .A(n54932), .B(n54931), .Z(n53555) );
  IV U73884 ( .A(n53555), .Z(n58865) );
  NOR U73885 ( .A(n53567), .B(n58865), .Z(n53550) );
  IV U73886 ( .A(n53550), .Z(n54924) );
  NOR U73887 ( .A(n53562), .B(n54924), .Z(n64070) );
  IV U73888 ( .A(n53551), .Z(n53553) );
  NOR U73889 ( .A(n53553), .B(n53552), .Z(n53556) );
  IV U73890 ( .A(n53556), .Z(n53554) );
  NOR U73891 ( .A(n53554), .B(n54931), .Z(n64060) );
  NOR U73892 ( .A(n53556), .B(n53555), .Z(n53557) );
  NOR U73893 ( .A(n64060), .B(n53557), .Z(n53561) );
  IV U73894 ( .A(n53558), .Z(n53559) );
  NOR U73895 ( .A(n53567), .B(n53559), .Z(n53560) );
  XOR U73896 ( .A(n53561), .B(n53560), .Z(n54919) );
  NOR U73897 ( .A(n53562), .B(n53567), .Z(n53563) );
  NOR U73898 ( .A(n54919), .B(n53563), .Z(n53564) );
  NOR U73899 ( .A(n64070), .B(n53564), .Z(n53572) );
  IV U73900 ( .A(n53565), .Z(n53566) );
  NOR U73901 ( .A(n53567), .B(n53566), .Z(n58863) );
  IV U73902 ( .A(n53568), .Z(n53569) );
  NOR U73903 ( .A(n53570), .B(n53569), .Z(n54920) );
  NOR U73904 ( .A(n58863), .B(n54920), .Z(n53571) );
  XOR U73905 ( .A(n53572), .B(n53571), .Z(n58868) );
  IV U73906 ( .A(n53573), .Z(n53575) );
  NOR U73907 ( .A(n53575), .B(n53574), .Z(n58866) );
  XOR U73908 ( .A(n58868), .B(n58866), .Z(n58870) );
  XOR U73909 ( .A(n58869), .B(n58870), .Z(n54915) );
  XOR U73910 ( .A(n53576), .B(n54915), .Z(n64095) );
  XOR U73911 ( .A(n53578), .B(n53577), .Z(n53579) );
  NOR U73912 ( .A(n53580), .B(n53579), .Z(n53581) );
  IV U73913 ( .A(n53581), .Z(n53584) );
  NOR U73914 ( .A(n53582), .B(n54916), .Z(n53583) );
  IV U73915 ( .A(n53583), .Z(n53590) );
  NOR U73916 ( .A(n53584), .B(n53590), .Z(n53585) );
  IV U73917 ( .A(n53585), .Z(n53592) );
  NOR U73918 ( .A(n64095), .B(n53592), .Z(n64115) );
  IV U73919 ( .A(n53586), .Z(n53587) );
  NOR U73920 ( .A(n53588), .B(n53587), .Z(n54909) );
  IV U73921 ( .A(n53589), .Z(n53591) );
  NOR U73922 ( .A(n53591), .B(n53590), .Z(n64094) );
  XOR U73923 ( .A(n64094), .B(n64095), .Z(n54910) );
  IV U73924 ( .A(n54910), .Z(n53593) );
  XOR U73925 ( .A(n54909), .B(n53593), .Z(n53595) );
  NOR U73926 ( .A(n53593), .B(n53592), .Z(n53594) );
  NOR U73927 ( .A(n53595), .B(n53594), .Z(n53596) );
  NOR U73928 ( .A(n64115), .B(n53596), .Z(n54907) );
  XOR U73929 ( .A(n53597), .B(n54907), .Z(n54905) );
  XOR U73930 ( .A(n54903), .B(n54905), .Z(n54902) );
  IV U73931 ( .A(n53598), .Z(n53607) );
  IV U73932 ( .A(n53599), .Z(n53600) );
  NOR U73933 ( .A(n53607), .B(n53600), .Z(n54898) );
  IV U73934 ( .A(n53601), .Z(n53602) );
  NOR U73935 ( .A(n53603), .B(n53602), .Z(n54900) );
  NOR U73936 ( .A(n54898), .B(n54900), .Z(n53604) );
  XOR U73937 ( .A(n54902), .B(n53604), .Z(n54893) );
  IV U73938 ( .A(n53605), .Z(n53606) );
  NOR U73939 ( .A(n53607), .B(n53606), .Z(n54890) );
  IV U73940 ( .A(n53608), .Z(n53610) );
  NOR U73941 ( .A(n53610), .B(n53609), .Z(n54894) );
  NOR U73942 ( .A(n54890), .B(n54894), .Z(n53611) );
  XOR U73943 ( .A(n54893), .B(n53611), .Z(n58883) );
  IV U73944 ( .A(n53612), .Z(n53614) );
  NOR U73945 ( .A(n53614), .B(n53613), .Z(n54889) );
  IV U73946 ( .A(n53615), .Z(n53616) );
  NOR U73947 ( .A(n53616), .B(n58891), .Z(n58882) );
  NOR U73948 ( .A(n54889), .B(n58882), .Z(n53617) );
  XOR U73949 ( .A(n58883), .B(n53617), .Z(n58879) );
  IV U73950 ( .A(n53618), .Z(n53619) );
  NOR U73951 ( .A(n53619), .B(n58891), .Z(n53620) );
  IV U73952 ( .A(n53620), .Z(n58880) );
  XOR U73953 ( .A(n58879), .B(n58880), .Z(n58887) );
  XOR U73954 ( .A(n53621), .B(n58887), .Z(n54884) );
  IV U73955 ( .A(n53622), .Z(n53624) );
  NOR U73956 ( .A(n53624), .B(n53623), .Z(n53625) );
  IV U73957 ( .A(n53625), .Z(n53632) );
  NOR U73958 ( .A(n54884), .B(n53632), .Z(n54882) );
  IV U73959 ( .A(n53626), .Z(n53631) );
  IV U73960 ( .A(n53627), .Z(n53628) );
  NOR U73961 ( .A(n53631), .B(n53628), .Z(n54886) );
  IV U73962 ( .A(n53629), .Z(n53630) );
  NOR U73963 ( .A(n53631), .B(n53630), .Z(n54883) );
  XOR U73964 ( .A(n54883), .B(n54884), .Z(n54887) );
  IV U73965 ( .A(n54887), .Z(n53633) );
  XOR U73966 ( .A(n54886), .B(n53633), .Z(n53635) );
  NOR U73967 ( .A(n53633), .B(n53632), .Z(n53634) );
  NOR U73968 ( .A(n53635), .B(n53634), .Z(n53636) );
  NOR U73969 ( .A(n54882), .B(n53636), .Z(n58893) );
  IV U73970 ( .A(n53637), .Z(n53639) );
  NOR U73971 ( .A(n53639), .B(n53638), .Z(n53640) );
  IV U73972 ( .A(n53640), .Z(n58894) );
  XOR U73973 ( .A(n58893), .B(n58894), .Z(n58897) );
  XOR U73974 ( .A(n58896), .B(n58897), .Z(n54880) );
  XOR U73975 ( .A(n54879), .B(n54880), .Z(n54874) );
  XOR U73976 ( .A(n54873), .B(n54874), .Z(n54878) );
  IV U73977 ( .A(n53641), .Z(n53643) );
  IV U73978 ( .A(n53642), .Z(n53645) );
  NOR U73979 ( .A(n53643), .B(n53645), .Z(n54876) );
  XOR U73980 ( .A(n54878), .B(n54876), .Z(n58902) );
  IV U73981 ( .A(n53644), .Z(n53646) );
  NOR U73982 ( .A(n53646), .B(n53645), .Z(n53647) );
  IV U73983 ( .A(n53647), .Z(n58901) );
  XOR U73984 ( .A(n58902), .B(n58901), .Z(n58904) );
  IV U73985 ( .A(n53648), .Z(n53649) );
  NOR U73986 ( .A(n53650), .B(n53649), .Z(n58903) );
  NOR U73987 ( .A(n53652), .B(n53651), .Z(n58907) );
  NOR U73988 ( .A(n58903), .B(n58907), .Z(n53653) );
  XOR U73989 ( .A(n58904), .B(n53653), .Z(n54869) );
  NOR U73990 ( .A(n53654), .B(n54867), .Z(n53655) );
  NOR U73991 ( .A(n53656), .B(n53655), .Z(n53657) );
  XOR U73992 ( .A(n54869), .B(n53657), .Z(n75892) );
  XOR U73993 ( .A(n58910), .B(n75892), .Z(n65485) );
  XOR U73994 ( .A(n65487), .B(n65485), .Z(n53658) );
  IV U73995 ( .A(n53658), .Z(n58916) );
  XOR U73996 ( .A(n53659), .B(n58916), .Z(n54852) );
  XOR U73997 ( .A(n54851), .B(n54852), .Z(n58919) );
  IV U73998 ( .A(n58919), .Z(n53664) );
  IV U73999 ( .A(n53660), .Z(n53661) );
  NOR U74000 ( .A(n53662), .B(n53661), .Z(n58918) );
  NOR U74001 ( .A(n58915), .B(n58918), .Z(n53663) );
  XOR U74002 ( .A(n53664), .B(n53663), .Z(n58923) );
  IV U74003 ( .A(n53665), .Z(n53667) );
  NOR U74004 ( .A(n53667), .B(n53666), .Z(n58921) );
  XOR U74005 ( .A(n58923), .B(n58921), .Z(n58926) );
  XOR U74006 ( .A(n53668), .B(n58926), .Z(n54843) );
  IV U74007 ( .A(n53669), .Z(n53671) );
  NOR U74008 ( .A(n53671), .B(n53670), .Z(n54845) );
  IV U74009 ( .A(n53672), .Z(n53674) );
  NOR U74010 ( .A(n53674), .B(n53673), .Z(n54842) );
  NOR U74011 ( .A(n54845), .B(n54842), .Z(n53675) );
  XOR U74012 ( .A(n54843), .B(n53675), .Z(n54838) );
  XOR U74013 ( .A(n54837), .B(n54838), .Z(n53676) );
  XOR U74014 ( .A(n53677), .B(n53676), .Z(n54821) );
  XOR U74015 ( .A(n53678), .B(n54821), .Z(n54819) );
  IV U74016 ( .A(n53679), .Z(n53683) );
  NOR U74017 ( .A(n53681), .B(n53680), .Z(n53682) );
  IV U74018 ( .A(n53682), .Z(n53685) );
  NOR U74019 ( .A(n53683), .B(n53685), .Z(n54817) );
  XOR U74020 ( .A(n54819), .B(n54817), .Z(n58934) );
  IV U74021 ( .A(n53684), .Z(n53686) );
  NOR U74022 ( .A(n53686), .B(n53685), .Z(n58932) );
  XOR U74023 ( .A(n58934), .B(n58932), .Z(n58940) );
  IV U74024 ( .A(n53687), .Z(n53704) );
  IV U74025 ( .A(n53688), .Z(n53689) );
  NOR U74026 ( .A(n53704), .B(n53689), .Z(n58939) );
  IV U74027 ( .A(n53690), .Z(n53692) );
  NOR U74028 ( .A(n53692), .B(n53691), .Z(n58935) );
  NOR U74029 ( .A(n58939), .B(n58935), .Z(n53693) );
  XOR U74030 ( .A(n58940), .B(n53693), .Z(n53706) );
  IV U74031 ( .A(n53706), .Z(n53698) );
  IV U74032 ( .A(n53694), .Z(n53696) );
  NOR U74033 ( .A(n53696), .B(n53695), .Z(n53710) );
  IV U74034 ( .A(n53710), .Z(n53697) );
  NOR U74035 ( .A(n53698), .B(n53697), .Z(n64203) );
  IV U74036 ( .A(n53699), .Z(n53700) );
  NOR U74037 ( .A(n53701), .B(n53700), .Z(n54813) );
  IV U74038 ( .A(n53702), .Z(n53703) );
  NOR U74039 ( .A(n53704), .B(n53703), .Z(n53707) );
  IV U74040 ( .A(n53707), .Z(n53705) );
  NOR U74041 ( .A(n53705), .B(n58940), .Z(n60158) );
  NOR U74042 ( .A(n53707), .B(n53706), .Z(n53708) );
  NOR U74043 ( .A(n60158), .B(n53708), .Z(n54814) );
  XOR U74044 ( .A(n54813), .B(n54814), .Z(n53709) );
  NOR U74045 ( .A(n53710), .B(n53709), .Z(n53711) );
  NOR U74046 ( .A(n64203), .B(n53711), .Z(n58943) );
  XOR U74047 ( .A(n53712), .B(n58943), .Z(n58949) );
  XOR U74048 ( .A(n58947), .B(n58949), .Z(n60152) );
  NOR U74049 ( .A(n53714), .B(n53713), .Z(n53715) );
  IV U74050 ( .A(n53715), .Z(n60146) );
  NOR U74051 ( .A(n53716), .B(n60146), .Z(n58954) );
  XOR U74052 ( .A(n60152), .B(n58954), .Z(n58961) );
  IV U74053 ( .A(n53717), .Z(n53719) );
  IV U74054 ( .A(n53718), .Z(n53726) );
  NOR U74055 ( .A(n53719), .B(n53726), .Z(n58956) );
  XOR U74056 ( .A(n53719), .B(n53718), .Z(n53722) );
  IV U74057 ( .A(n53720), .Z(n53721) );
  NOR U74058 ( .A(n53722), .B(n53721), .Z(n58960) );
  NOR U74059 ( .A(n58956), .B(n58960), .Z(n53723) );
  XOR U74060 ( .A(n58961), .B(n53723), .Z(n54807) );
  IV U74061 ( .A(n53724), .Z(n53725) );
  NOR U74062 ( .A(n53726), .B(n53725), .Z(n54810) );
  IV U74063 ( .A(n53727), .Z(n53728) );
  NOR U74064 ( .A(n53728), .B(n53731), .Z(n54808) );
  NOR U74065 ( .A(n54810), .B(n54808), .Z(n53729) );
  XOR U74066 ( .A(n54807), .B(n53729), .Z(n54806) );
  IV U74067 ( .A(n53730), .Z(n53735) );
  NOR U74068 ( .A(n53732), .B(n53731), .Z(n53733) );
  IV U74069 ( .A(n53733), .Z(n53734) );
  NOR U74070 ( .A(n53735), .B(n53734), .Z(n54804) );
  XOR U74071 ( .A(n54806), .B(n54804), .Z(n58966) );
  XOR U74072 ( .A(n58965), .B(n58966), .Z(n54800) );
  NOR U74073 ( .A(n53737), .B(n53736), .Z(n53738) );
  IV U74074 ( .A(n53738), .Z(n54801) );
  IV U74075 ( .A(n53739), .Z(n54803) );
  NOR U74076 ( .A(n54801), .B(n54803), .Z(n53740) );
  XOR U74077 ( .A(n54800), .B(n53740), .Z(n58973) );
  IV U74078 ( .A(n53741), .Z(n53743) );
  NOR U74079 ( .A(n53743), .B(n53742), .Z(n58971) );
  XOR U74080 ( .A(n58973), .B(n58971), .Z(n60122) );
  XOR U74081 ( .A(n53744), .B(n60122), .Z(n58985) );
  XOR U74082 ( .A(n58984), .B(n58985), .Z(n58979) );
  XOR U74083 ( .A(n58977), .B(n58979), .Z(n58982) );
  XOR U74084 ( .A(n58981), .B(n58982), .Z(n54790) );
  XOR U74085 ( .A(n53745), .B(n54790), .Z(n58995) );
  XOR U74086 ( .A(n58993), .B(n58995), .Z(n58998) );
  XOR U74087 ( .A(n58996), .B(n58998), .Z(n59001) );
  XOR U74088 ( .A(n59000), .B(n59001), .Z(n59004) );
  XOR U74089 ( .A(n59003), .B(n59004), .Z(n59008) );
  XOR U74090 ( .A(n53746), .B(n59008), .Z(n54787) );
  XOR U74091 ( .A(n54784), .B(n54787), .Z(n53747) );
  NOR U74092 ( .A(n65380), .B(n53747), .Z(n64238) );
  IV U74093 ( .A(n53748), .Z(n53750) );
  NOR U74094 ( .A(n53750), .B(n53749), .Z(n54786) );
  NOR U74095 ( .A(n54784), .B(n54786), .Z(n53751) );
  XOR U74096 ( .A(n53751), .B(n54787), .Z(n65383) );
  NOR U74097 ( .A(n53752), .B(n65383), .Z(n53753) );
  NOR U74098 ( .A(n64238), .B(n53753), .Z(n53754) );
  IV U74099 ( .A(n53754), .Z(n54777) );
  XOR U74100 ( .A(n53755), .B(n54777), .Z(n54775) );
  XOR U74101 ( .A(n54773), .B(n54775), .Z(n59024) );
  XOR U74102 ( .A(n59023), .B(n59024), .Z(n59026) );
  XOR U74103 ( .A(n59027), .B(n59026), .Z(n54770) );
  IV U74104 ( .A(n53756), .Z(n53760) );
  NOR U74105 ( .A(n53758), .B(n53757), .Z(n53759) );
  IV U74106 ( .A(n53759), .Z(n53762) );
  NOR U74107 ( .A(n53760), .B(n53762), .Z(n54771) );
  IV U74108 ( .A(n53761), .Z(n53763) );
  NOR U74109 ( .A(n53763), .B(n53762), .Z(n65363) );
  NOR U74110 ( .A(n65369), .B(n65363), .Z(n60081) );
  IV U74111 ( .A(n60081), .Z(n53764) );
  NOR U74112 ( .A(n54771), .B(n53764), .Z(n53765) );
  XOR U74113 ( .A(n54770), .B(n53765), .Z(n54766) );
  XOR U74114 ( .A(n54765), .B(n54766), .Z(n59032) );
  IV U74115 ( .A(n53766), .Z(n53767) );
  NOR U74116 ( .A(n53768), .B(n53767), .Z(n54768) );
  IV U74117 ( .A(n53769), .Z(n53771) );
  NOR U74118 ( .A(n53771), .B(n53770), .Z(n59031) );
  NOR U74119 ( .A(n54768), .B(n59031), .Z(n53772) );
  XOR U74120 ( .A(n59032), .B(n53772), .Z(n53773) );
  IV U74121 ( .A(n53773), .Z(n59034) );
  NOR U74122 ( .A(n53780), .B(n59034), .Z(n59041) );
  IV U74123 ( .A(n53774), .Z(n53776) );
  NOR U74124 ( .A(n53776), .B(n53775), .Z(n59038) );
  IV U74125 ( .A(n53777), .Z(n53779) );
  NOR U74126 ( .A(n53779), .B(n53778), .Z(n59033) );
  XOR U74127 ( .A(n59033), .B(n59034), .Z(n59039) );
  IV U74128 ( .A(n59039), .Z(n53781) );
  XOR U74129 ( .A(n59038), .B(n53781), .Z(n53783) );
  NOR U74130 ( .A(n53781), .B(n53780), .Z(n53782) );
  NOR U74131 ( .A(n53783), .B(n53782), .Z(n53784) );
  NOR U74132 ( .A(n59041), .B(n53784), .Z(n54760) );
  XOR U74133 ( .A(n54761), .B(n54760), .Z(n54759) );
  IV U74134 ( .A(n53785), .Z(n53786) );
  NOR U74135 ( .A(n53787), .B(n53786), .Z(n54762) );
  IV U74136 ( .A(n53788), .Z(n53789) );
  NOR U74137 ( .A(n53789), .B(n53793), .Z(n54757) );
  NOR U74138 ( .A(n54762), .B(n54757), .Z(n53790) );
  XOR U74139 ( .A(n54759), .B(n53790), .Z(n53791) );
  IV U74140 ( .A(n53791), .Z(n59051) );
  IV U74141 ( .A(n53792), .Z(n53794) );
  NOR U74142 ( .A(n53794), .B(n53793), .Z(n59049) );
  XOR U74143 ( .A(n59051), .B(n59049), .Z(n54755) );
  XOR U74144 ( .A(n54753), .B(n54755), .Z(n59048) );
  IV U74145 ( .A(n53795), .Z(n53796) );
  NOR U74146 ( .A(n53797), .B(n53796), .Z(n54751) );
  IV U74147 ( .A(n53798), .Z(n53800) );
  NOR U74148 ( .A(n53800), .B(n53799), .Z(n59046) );
  NOR U74149 ( .A(n54751), .B(n59046), .Z(n53801) );
  XOR U74150 ( .A(n59048), .B(n53801), .Z(n53802) );
  NOR U74151 ( .A(n53803), .B(n53802), .Z(n53806) );
  IV U74152 ( .A(n53803), .Z(n53805) );
  XOR U74153 ( .A(n59046), .B(n59048), .Z(n53804) );
  NOR U74154 ( .A(n53805), .B(n53804), .Z(n60053) );
  NOR U74155 ( .A(n53806), .B(n60053), .Z(n53807) );
  IV U74156 ( .A(n53807), .Z(n59062) );
  NOR U74157 ( .A(n59065), .B(n59058), .Z(n53808) );
  NOR U74158 ( .A(n53809), .B(n53808), .Z(n53810) );
  XOR U74159 ( .A(n59062), .B(n53810), .Z(n54748) );
  XOR U74160 ( .A(n54747), .B(n54748), .Z(n54743) );
  IV U74161 ( .A(n53811), .Z(n53812) );
  NOR U74162 ( .A(n53813), .B(n53812), .Z(n54745) );
  IV U74163 ( .A(n53814), .Z(n53815) );
  NOR U74164 ( .A(n53816), .B(n53815), .Z(n54742) );
  NOR U74165 ( .A(n54745), .B(n54742), .Z(n53817) );
  XOR U74166 ( .A(n54743), .B(n53817), .Z(n53818) );
  IV U74167 ( .A(n53818), .Z(n54741) );
  IV U74168 ( .A(n53819), .Z(n53824) );
  NOR U74169 ( .A(n53821), .B(n53820), .Z(n53822) );
  IV U74170 ( .A(n53822), .Z(n53823) );
  NOR U74171 ( .A(n53824), .B(n53823), .Z(n54739) );
  XOR U74172 ( .A(n54741), .B(n54739), .Z(n54735) );
  XOR U74173 ( .A(n54733), .B(n54735), .Z(n54737) );
  XOR U74174 ( .A(n54736), .B(n54737), .Z(n54729) );
  XOR U74175 ( .A(n54727), .B(n54729), .Z(n54732) );
  XOR U74176 ( .A(n54730), .B(n54732), .Z(n59072) );
  XOR U74177 ( .A(n59071), .B(n59072), .Z(n53829) );
  IV U74178 ( .A(n53829), .Z(n59073) );
  XOR U74179 ( .A(n54722), .B(n59073), .Z(n53825) );
  NOR U74180 ( .A(n53835), .B(n53825), .Z(n64280) );
  IV U74181 ( .A(n53826), .Z(n53828) );
  NOR U74182 ( .A(n53828), .B(n53827), .Z(n54719) );
  NOR U74183 ( .A(n54722), .B(n54719), .Z(n53830) );
  XOR U74184 ( .A(n53830), .B(n53829), .Z(n54718) );
  IV U74185 ( .A(n53831), .Z(n53834) );
  IV U74186 ( .A(n53832), .Z(n53833) );
  NOR U74187 ( .A(n53834), .B(n53833), .Z(n53836) );
  IV U74188 ( .A(n53836), .Z(n54717) );
  XOR U74189 ( .A(n54718), .B(n54717), .Z(n53838) );
  NOR U74190 ( .A(n53836), .B(n53835), .Z(n53837) );
  NOR U74191 ( .A(n53838), .B(n53837), .Z(n53839) );
  NOR U74192 ( .A(n64280), .B(n53839), .Z(n54709) );
  IV U74193 ( .A(n53840), .Z(n53841) );
  NOR U74194 ( .A(n53842), .B(n53841), .Z(n54714) );
  IV U74195 ( .A(n53843), .Z(n53845) );
  NOR U74196 ( .A(n53845), .B(n53844), .Z(n53846) );
  NOR U74197 ( .A(n54714), .B(n53846), .Z(n54710) );
  XOR U74198 ( .A(n54709), .B(n54710), .Z(n59088) );
  XOR U74199 ( .A(n59085), .B(n59088), .Z(n54703) );
  XOR U74200 ( .A(n54704), .B(n54703), .Z(n53847) );
  IV U74201 ( .A(n53847), .Z(n54701) );
  IV U74202 ( .A(n53848), .Z(n53850) );
  NOR U74203 ( .A(n53850), .B(n53849), .Z(n54700) );
  IV U74204 ( .A(n53851), .Z(n53852) );
  NOR U74205 ( .A(n53853), .B(n53852), .Z(n54698) );
  NOR U74206 ( .A(n54700), .B(n54698), .Z(n53854) );
  XOR U74207 ( .A(n54701), .B(n53854), .Z(n54691) );
  NOR U74208 ( .A(n53856), .B(n53855), .Z(n54695) );
  NOR U74209 ( .A(n54695), .B(n54692), .Z(n53857) );
  XOR U74210 ( .A(n54691), .B(n53857), .Z(n59092) );
  XOR U74211 ( .A(n59091), .B(n59092), .Z(n59095) );
  XOR U74212 ( .A(n59094), .B(n59095), .Z(n54687) );
  IV U74213 ( .A(n53858), .Z(n53860) );
  NOR U74214 ( .A(n53860), .B(n53859), .Z(n54688) );
  IV U74215 ( .A(n53861), .Z(n53866) );
  IV U74216 ( .A(n53862), .Z(n53863) );
  NOR U74217 ( .A(n53864), .B(n53863), .Z(n53865) );
  IV U74218 ( .A(n53865), .Z(n53869) );
  NOR U74219 ( .A(n53866), .B(n53869), .Z(n54685) );
  NOR U74220 ( .A(n54688), .B(n54685), .Z(n53867) );
  XOR U74221 ( .A(n54687), .B(n53867), .Z(n54679) );
  IV U74222 ( .A(n53868), .Z(n53870) );
  NOR U74223 ( .A(n53870), .B(n53869), .Z(n53871) );
  IV U74224 ( .A(n53871), .Z(n54680) );
  XOR U74225 ( .A(n54679), .B(n54680), .Z(n54684) );
  XOR U74226 ( .A(n53872), .B(n54684), .Z(n54671) );
  XOR U74227 ( .A(n53873), .B(n54671), .Z(n54668) );
  XOR U74228 ( .A(n54666), .B(n54668), .Z(n64340) );
  XOR U74229 ( .A(n54669), .B(n64340), .Z(n53874) );
  IV U74230 ( .A(n53874), .Z(n54662) );
  XOR U74231 ( .A(n54661), .B(n54662), .Z(n54664) );
  XOR U74232 ( .A(n54665), .B(n54664), .Z(n54648) );
  NOR U74233 ( .A(n54653), .B(n53875), .Z(n53879) );
  IV U74234 ( .A(n53876), .Z(n54643) );
  IV U74235 ( .A(n53877), .Z(n53878) );
  NOR U74236 ( .A(n54643), .B(n53878), .Z(n59103) );
  NOR U74237 ( .A(n53879), .B(n59103), .Z(n53880) );
  XOR U74238 ( .A(n54648), .B(n53880), .Z(n54646) );
  IV U74239 ( .A(n53881), .Z(n53882) );
  NOR U74240 ( .A(n54643), .B(n53882), .Z(n54644) );
  XOR U74241 ( .A(n54646), .B(n54644), .Z(n59110) );
  XOR U74242 ( .A(n53883), .B(n59110), .Z(n59108) );
  XOR U74243 ( .A(n59106), .B(n59108), .Z(n59114) );
  XOR U74244 ( .A(n59113), .B(n59114), .Z(n54636) );
  XOR U74245 ( .A(n53884), .B(n54636), .Z(n59122) );
  IV U74246 ( .A(n53885), .Z(n53890) );
  IV U74247 ( .A(n53886), .Z(n53887) );
  NOR U74248 ( .A(n53888), .B(n53887), .Z(n53889) );
  IV U74249 ( .A(n53889), .Z(n53892) );
  NOR U74250 ( .A(n53890), .B(n53892), .Z(n59120) );
  XOR U74251 ( .A(n59122), .B(n59120), .Z(n59125) );
  IV U74252 ( .A(n53891), .Z(n53893) );
  NOR U74253 ( .A(n53893), .B(n53892), .Z(n59123) );
  XOR U74254 ( .A(n59125), .B(n59123), .Z(n59128) );
  XOR U74255 ( .A(n59127), .B(n59128), .Z(n59131) );
  XOR U74256 ( .A(n59130), .B(n59131), .Z(n54633) );
  XOR U74257 ( .A(n54632), .B(n54633), .Z(n54630) );
  XOR U74258 ( .A(n54629), .B(n54630), .Z(n59947) );
  XOR U74259 ( .A(n53894), .B(n59947), .Z(n59135) );
  XOR U74260 ( .A(n59136), .B(n59135), .Z(n53901) );
  IV U74261 ( .A(n53901), .Z(n53895) );
  NOR U74262 ( .A(n53899), .B(n53895), .Z(n53896) );
  IV U74263 ( .A(n53896), .Z(n53897) );
  NOR U74264 ( .A(n53898), .B(n53897), .Z(n59940) );
  NOR U74265 ( .A(n53900), .B(n53899), .Z(n53902) );
  NOR U74266 ( .A(n53902), .B(n53901), .Z(n53903) );
  NOR U74267 ( .A(n59940), .B(n53903), .Z(n53904) );
  IV U74268 ( .A(n53904), .Z(n59141) );
  XOR U74269 ( .A(n59140), .B(n59141), .Z(n59153) );
  IV U74270 ( .A(n53905), .Z(n53907) );
  NOR U74271 ( .A(n53907), .B(n53906), .Z(n59144) );
  IV U74272 ( .A(n53908), .Z(n53915) );
  XOR U74273 ( .A(n53910), .B(n53909), .Z(n53912) );
  NOR U74274 ( .A(n53912), .B(n53911), .Z(n53913) );
  IV U74275 ( .A(n53913), .Z(n53914) );
  NOR U74276 ( .A(n53915), .B(n53914), .Z(n59151) );
  NOR U74277 ( .A(n59144), .B(n59151), .Z(n53916) );
  XOR U74278 ( .A(n59153), .B(n53916), .Z(n59154) );
  XOR U74279 ( .A(n59156), .B(n59154), .Z(n54625) );
  XOR U74280 ( .A(n53917), .B(n54625), .Z(n54622) );
  XOR U74281 ( .A(n53918), .B(n54622), .Z(n54613) );
  XOR U74282 ( .A(n53919), .B(n54613), .Z(n54608) );
  XOR U74283 ( .A(n54607), .B(n54608), .Z(n54611) );
  XOR U74284 ( .A(n53920), .B(n54611), .Z(n59163) );
  XOR U74285 ( .A(n59164), .B(n59163), .Z(n59167) );
  XOR U74286 ( .A(n59166), .B(n59167), .Z(n54600) );
  XOR U74287 ( .A(n54599), .B(n54600), .Z(n54604) );
  IV U74288 ( .A(n53921), .Z(n53923) );
  NOR U74289 ( .A(n53923), .B(n53922), .Z(n54602) );
  XOR U74290 ( .A(n54604), .B(n54602), .Z(n59172) );
  XOR U74291 ( .A(n59171), .B(n59172), .Z(n59904) );
  IV U74292 ( .A(n59904), .Z(n53930) );
  IV U74293 ( .A(n53924), .Z(n53925) );
  NOR U74294 ( .A(n53926), .B(n53925), .Z(n59907) );
  IV U74295 ( .A(n53927), .Z(n53928) );
  NOR U74296 ( .A(n53929), .B(n53928), .Z(n59903) );
  NOR U74297 ( .A(n59907), .B(n59903), .Z(n59174) );
  XOR U74298 ( .A(n53930), .B(n59174), .Z(n59181) );
  XOR U74299 ( .A(n59180), .B(n59181), .Z(n59188) );
  XOR U74300 ( .A(n53931), .B(n59188), .Z(n59190) );
  XOR U74301 ( .A(n53932), .B(n59190), .Z(n59198) );
  XOR U74302 ( .A(n53933), .B(n59198), .Z(n59203) );
  XOR U74303 ( .A(n59202), .B(n59203), .Z(n54598) );
  XOR U74304 ( .A(n53934), .B(n54598), .Z(n54588) );
  XOR U74305 ( .A(n54590), .B(n54588), .Z(n54592) );
  NOR U74306 ( .A(n53936), .B(n53935), .Z(n54591) );
  NOR U74307 ( .A(n53938), .B(n53937), .Z(n54586) );
  NOR U74308 ( .A(n54591), .B(n54586), .Z(n53939) );
  XOR U74309 ( .A(n54592), .B(n53939), .Z(n53940) );
  IV U74310 ( .A(n53940), .Z(n54584) );
  XOR U74311 ( .A(n54582), .B(n54584), .Z(n59215) );
  XOR U74312 ( .A(n59213), .B(n59215), .Z(n59220) );
  XOR U74313 ( .A(n59216), .B(n59220), .Z(n54580) );
  XOR U74314 ( .A(n53941), .B(n54580), .Z(n53942) );
  IV U74315 ( .A(n53942), .Z(n59229) );
  XOR U74316 ( .A(n59227), .B(n59229), .Z(n59233) );
  XOR U74317 ( .A(n59232), .B(n59233), .Z(n59236) );
  XOR U74318 ( .A(n59235), .B(n59236), .Z(n59240) );
  XOR U74319 ( .A(n59239), .B(n59240), .Z(n59244) );
  IV U74320 ( .A(n53943), .Z(n53944) );
  NOR U74321 ( .A(n53947), .B(n53944), .Z(n59242) );
  XOR U74322 ( .A(n59244), .B(n59242), .Z(n59248) );
  IV U74323 ( .A(n53945), .Z(n53946) );
  NOR U74324 ( .A(n53947), .B(n53946), .Z(n59246) );
  XOR U74325 ( .A(n59248), .B(n59246), .Z(n59250) );
  XOR U74326 ( .A(n59249), .B(n59250), .Z(n59254) );
  XOR U74327 ( .A(n59253), .B(n59254), .Z(n59257) );
  XOR U74328 ( .A(n59256), .B(n59257), .Z(n59261) );
  XOR U74329 ( .A(n59260), .B(n59261), .Z(n53961) );
  IV U74330 ( .A(n53961), .Z(n53955) );
  IV U74331 ( .A(n53948), .Z(n53957) );
  NOR U74332 ( .A(n65162), .B(n53957), .Z(n53952) );
  IV U74333 ( .A(n53949), .Z(n53951) );
  NOR U74334 ( .A(n53951), .B(n53950), .Z(n53960) );
  NOR U74335 ( .A(n53952), .B(n53960), .Z(n53953) );
  IV U74336 ( .A(n53953), .Z(n53954) );
  NOR U74337 ( .A(n53955), .B(n53954), .Z(n53964) );
  XOR U74338 ( .A(n53956), .B(n65162), .Z(n53959) );
  NOR U74339 ( .A(n53957), .B(n53961), .Z(n53958) );
  IV U74340 ( .A(n53958), .Z(n65168) );
  NOR U74341 ( .A(n53959), .B(n65168), .Z(n59263) );
  IV U74342 ( .A(n53960), .Z(n53962) );
  NOR U74343 ( .A(n53962), .B(n53961), .Z(n69650) );
  NOR U74344 ( .A(n59263), .B(n69650), .Z(n64479) );
  IV U74345 ( .A(n64479), .Z(n53963) );
  NOR U74346 ( .A(n53964), .B(n53963), .Z(n59265) );
  IV U74347 ( .A(n53965), .Z(n53967) );
  NOR U74348 ( .A(n53967), .B(n53966), .Z(n53968) );
  IV U74349 ( .A(n53968), .Z(n59266) );
  XOR U74350 ( .A(n59265), .B(n59266), .Z(n59275) );
  XOR U74351 ( .A(n59273), .B(n59275), .Z(n59277) );
  IV U74352 ( .A(n53969), .Z(n53979) );
  IV U74353 ( .A(n53970), .Z(n53971) );
  NOR U74354 ( .A(n53972), .B(n53971), .Z(n53977) );
  NOR U74355 ( .A(n53974), .B(n53973), .Z(n53975) );
  IV U74356 ( .A(n53975), .Z(n53976) );
  NOR U74357 ( .A(n53977), .B(n53976), .Z(n53978) );
  IV U74358 ( .A(n53978), .Z(n53981) );
  NOR U74359 ( .A(n53979), .B(n53981), .Z(n59270) );
  IV U74360 ( .A(n53980), .Z(n53982) );
  NOR U74361 ( .A(n53982), .B(n53981), .Z(n59276) );
  NOR U74362 ( .A(n59270), .B(n59276), .Z(n53983) );
  XOR U74363 ( .A(n59277), .B(n53983), .Z(n53984) );
  NOR U74364 ( .A(n53985), .B(n53984), .Z(n53988) );
  XOR U74365 ( .A(n59276), .B(n59277), .Z(n53987) );
  IV U74366 ( .A(n53985), .Z(n53986) );
  NOR U74367 ( .A(n53987), .B(n53986), .Z(n59870) );
  NOR U74368 ( .A(n53988), .B(n59870), .Z(n53989) );
  IV U74369 ( .A(n53989), .Z(n59282) );
  IV U74370 ( .A(n53990), .Z(n53992) );
  NOR U74371 ( .A(n53992), .B(n53991), .Z(n59280) );
  XOR U74372 ( .A(n59282), .B(n59280), .Z(n54578) );
  XOR U74373 ( .A(n54574), .B(n54578), .Z(n53993) );
  NOR U74374 ( .A(n53994), .B(n53993), .Z(n59864) );
  IV U74375 ( .A(n53995), .Z(n53997) );
  NOR U74376 ( .A(n53997), .B(n53996), .Z(n54576) );
  NOR U74377 ( .A(n54574), .B(n54576), .Z(n53998) );
  XOR U74378 ( .A(n54578), .B(n53998), .Z(n53999) );
  NOR U74379 ( .A(n54000), .B(n53999), .Z(n54001) );
  NOR U74380 ( .A(n59864), .B(n54001), .Z(n54571) );
  IV U74381 ( .A(n54002), .Z(n54003) );
  NOR U74382 ( .A(n54003), .B(n54012), .Z(n54004) );
  IV U74383 ( .A(n54004), .Z(n54572) );
  XOR U74384 ( .A(n54571), .B(n54572), .Z(n54564) );
  IV U74385 ( .A(n54005), .Z(n54006) );
  NOR U74386 ( .A(n54006), .B(n54012), .Z(n54562) );
  XOR U74387 ( .A(n54564), .B(n54562), .Z(n54567) );
  NOR U74388 ( .A(n54008), .B(n54007), .Z(n54009) );
  IV U74389 ( .A(n54009), .Z(n54010) );
  NOR U74390 ( .A(n54011), .B(n54010), .Z(n54016) );
  NOR U74391 ( .A(n54013), .B(n54012), .Z(n54014) );
  IV U74392 ( .A(n54014), .Z(n54015) );
  NOR U74393 ( .A(n54016), .B(n54015), .Z(n54017) );
  IV U74394 ( .A(n54017), .Z(n54566) );
  NOR U74395 ( .A(n54018), .B(n54566), .Z(n54019) );
  XOR U74396 ( .A(n54567), .B(n54019), .Z(n54553) );
  IV U74397 ( .A(n54020), .Z(n54021) );
  NOR U74398 ( .A(n54022), .B(n54021), .Z(n54551) );
  XOR U74399 ( .A(n54553), .B(n54551), .Z(n54555) );
  XOR U74400 ( .A(n54554), .B(n54555), .Z(n54544) );
  IV U74401 ( .A(n54023), .Z(n54024) );
  NOR U74402 ( .A(n54025), .B(n54024), .Z(n54541) );
  NOR U74403 ( .A(n54543), .B(n54541), .Z(n54026) );
  XOR U74404 ( .A(n54544), .B(n54026), .Z(n54539) );
  XOR U74405 ( .A(n54027), .B(n54539), .Z(n54536) );
  IV U74406 ( .A(n54028), .Z(n54029) );
  NOR U74407 ( .A(n54030), .B(n54029), .Z(n54535) );
  IV U74408 ( .A(n54031), .Z(n54033) );
  NOR U74409 ( .A(n54033), .B(n54032), .Z(n54530) );
  NOR U74410 ( .A(n54535), .B(n54530), .Z(n54034) );
  XOR U74411 ( .A(n54536), .B(n54034), .Z(n54532) );
  XOR U74412 ( .A(n54534), .B(n54532), .Z(n54523) );
  XOR U74413 ( .A(n54035), .B(n54523), .Z(n59293) );
  XOR U74414 ( .A(n59291), .B(n59293), .Z(n54521) );
  XOR U74415 ( .A(n54520), .B(n54521), .Z(n59306) );
  XOR U74416 ( .A(n59304), .B(n59306), .Z(n59308) );
  XOR U74417 ( .A(n59307), .B(n59308), .Z(n59832) );
  XOR U74418 ( .A(n54036), .B(n59832), .Z(n59315) );
  NOR U74419 ( .A(n59318), .B(n54517), .Z(n54037) );
  NOR U74420 ( .A(n54038), .B(n54037), .Z(n54039) );
  XOR U74421 ( .A(n59315), .B(n54039), .Z(n54514) );
  IV U74422 ( .A(n54040), .Z(n54042) );
  IV U74423 ( .A(n54041), .Z(n59316) );
  NOR U74424 ( .A(n54042), .B(n59316), .Z(n54512) );
  XOR U74425 ( .A(n54514), .B(n54512), .Z(n59327) );
  XOR U74426 ( .A(n59313), .B(n59327), .Z(n59335) );
  IV U74427 ( .A(n59335), .Z(n54051) );
  IV U74428 ( .A(n54043), .Z(n54044) );
  NOR U74429 ( .A(n54044), .B(n54046), .Z(n59326) );
  IV U74430 ( .A(n54045), .Z(n54049) );
  NOR U74431 ( .A(n54047), .B(n54046), .Z(n54048) );
  IV U74432 ( .A(n54048), .Z(n54053) );
  NOR U74433 ( .A(n54049), .B(n54053), .Z(n59333) );
  NOR U74434 ( .A(n59326), .B(n59333), .Z(n54050) );
  XOR U74435 ( .A(n54051), .B(n54050), .Z(n59332) );
  IV U74436 ( .A(n54052), .Z(n54054) );
  NOR U74437 ( .A(n54054), .B(n54053), .Z(n59330) );
  XOR U74438 ( .A(n59332), .B(n59330), .Z(n54510) );
  XOR U74439 ( .A(n54509), .B(n54510), .Z(n54505) );
  XOR U74440 ( .A(n54503), .B(n54505), .Z(n54508) );
  XOR U74441 ( .A(n54055), .B(n54508), .Z(n54495) );
  XOR U74442 ( .A(n54056), .B(n54495), .Z(n59341) );
  XOR U74443 ( .A(n54057), .B(n59341), .Z(n54058) );
  IV U74444 ( .A(n54058), .Z(n54492) );
  XOR U74445 ( .A(n54490), .B(n54492), .Z(n59346) );
  IV U74446 ( .A(n54059), .Z(n54061) );
  NOR U74447 ( .A(n54061), .B(n54060), .Z(n59344) );
  XOR U74448 ( .A(n59346), .B(n59344), .Z(n59351) );
  IV U74449 ( .A(n54062), .Z(n54064) );
  NOR U74450 ( .A(n54064), .B(n54063), .Z(n59347) );
  XOR U74451 ( .A(n59351), .B(n59347), .Z(n54489) );
  XOR U74452 ( .A(n59352), .B(n54489), .Z(n54065) );
  XOR U74453 ( .A(n54488), .B(n54065), .Z(n54486) );
  XOR U74454 ( .A(n54485), .B(n54486), .Z(n54480) );
  XOR U74455 ( .A(n54479), .B(n54480), .Z(n54483) );
  IV U74456 ( .A(n54066), .Z(n54068) );
  NOR U74457 ( .A(n54068), .B(n54067), .Z(n54482) );
  IV U74458 ( .A(n54069), .Z(n54071) );
  NOR U74459 ( .A(n54071), .B(n54070), .Z(n54474) );
  NOR U74460 ( .A(n54482), .B(n54474), .Z(n54072) );
  XOR U74461 ( .A(n54483), .B(n54072), .Z(n54073) );
  IV U74462 ( .A(n54073), .Z(n54477) );
  XOR U74463 ( .A(n54476), .B(n54477), .Z(n54472) );
  XOR U74464 ( .A(n54471), .B(n54472), .Z(n54466) );
  XOR U74465 ( .A(n54465), .B(n54466), .Z(n54469) );
  XOR U74466 ( .A(n54074), .B(n54469), .Z(n54075) );
  IV U74467 ( .A(n54075), .Z(n54462) );
  XOR U74468 ( .A(n54460), .B(n54462), .Z(n54457) );
  IV U74469 ( .A(n54076), .Z(n54078) );
  NOR U74470 ( .A(n54078), .B(n54077), .Z(n54455) );
  XOR U74471 ( .A(n54457), .B(n54455), .Z(n54459) );
  IV U74472 ( .A(n54459), .Z(n70169) );
  IV U74473 ( .A(n54079), .Z(n54080) );
  NOR U74474 ( .A(n54083), .B(n54080), .Z(n54458) );
  IV U74475 ( .A(n54081), .Z(n54082) );
  NOR U74476 ( .A(n54083), .B(n54082), .Z(n54451) );
  NOR U74477 ( .A(n54458), .B(n54451), .Z(n54084) );
  XOR U74478 ( .A(n70169), .B(n54084), .Z(n54453) );
  XOR U74479 ( .A(n54085), .B(n54453), .Z(n54086) );
  XOR U74480 ( .A(n54087), .B(n54086), .Z(n54437) );
  XOR U74481 ( .A(n54435), .B(n54437), .Z(n54432) );
  IV U74482 ( .A(n54088), .Z(n54090) );
  NOR U74483 ( .A(n54090), .B(n54089), .Z(n54428) );
  IV U74484 ( .A(n54091), .Z(n54093) );
  NOR U74485 ( .A(n54093), .B(n54092), .Z(n54430) );
  NOR U74486 ( .A(n54428), .B(n54430), .Z(n54094) );
  XOR U74487 ( .A(n54432), .B(n54094), .Z(n54426) );
  XOR U74488 ( .A(n54427), .B(n54426), .Z(n59749) );
  XOR U74489 ( .A(n54420), .B(n59749), .Z(n54424) );
  IV U74490 ( .A(n54095), .Z(n54106) );
  IV U74491 ( .A(n54096), .Z(n54097) );
  NOR U74492 ( .A(n54106), .B(n54097), .Z(n54418) );
  IV U74493 ( .A(n54098), .Z(n54100) );
  NOR U74494 ( .A(n54100), .B(n54099), .Z(n54422) );
  NOR U74495 ( .A(n54418), .B(n54422), .Z(n54101) );
  XOR U74496 ( .A(n54424), .B(n54101), .Z(n54412) );
  IV U74497 ( .A(n54102), .Z(n54103) );
  NOR U74498 ( .A(n54106), .B(n54103), .Z(n54413) );
  IV U74499 ( .A(n54104), .Z(n54105) );
  NOR U74500 ( .A(n54106), .B(n54105), .Z(n54415) );
  NOR U74501 ( .A(n54413), .B(n54415), .Z(n54107) );
  XOR U74502 ( .A(n54412), .B(n54107), .Z(n59365) );
  IV U74503 ( .A(n54108), .Z(n54109) );
  NOR U74504 ( .A(n54110), .B(n54109), .Z(n59364) );
  IV U74505 ( .A(n54111), .Z(n54113) );
  NOR U74506 ( .A(n54113), .B(n54112), .Z(n59363) );
  NOR U74507 ( .A(n59364), .B(n59363), .Z(n54114) );
  XOR U74508 ( .A(n59365), .B(n54114), .Z(n54124) );
  IV U74509 ( .A(n54124), .Z(n54120) );
  IV U74510 ( .A(n54115), .Z(n54118) );
  IV U74511 ( .A(n54116), .Z(n54117) );
  NOR U74512 ( .A(n54118), .B(n54117), .Z(n54128) );
  IV U74513 ( .A(n54128), .Z(n54119) );
  NOR U74514 ( .A(n54120), .B(n54119), .Z(n59735) );
  NOR U74515 ( .A(n54121), .B(n54131), .Z(n54125) );
  IV U74516 ( .A(n54125), .Z(n54123) );
  XOR U74517 ( .A(n59364), .B(n59365), .Z(n54122) );
  NOR U74518 ( .A(n54123), .B(n54122), .Z(n64593) );
  NOR U74519 ( .A(n54125), .B(n54124), .Z(n54126) );
  NOR U74520 ( .A(n64593), .B(n54126), .Z(n54127) );
  NOR U74521 ( .A(n54128), .B(n54127), .Z(n54129) );
  NOR U74522 ( .A(n59735), .B(n54129), .Z(n59371) );
  IV U74523 ( .A(n54130), .Z(n54132) );
  NOR U74524 ( .A(n54132), .B(n54131), .Z(n54133) );
  IV U74525 ( .A(n54133), .Z(n59372) );
  XOR U74526 ( .A(n59371), .B(n59372), .Z(n59375) );
  XOR U74527 ( .A(n59374), .B(n59375), .Z(n54409) );
  IV U74528 ( .A(n54409), .Z(n54139) );
  NOR U74529 ( .A(n54135), .B(n54134), .Z(n54408) );
  NOR U74530 ( .A(n54137), .B(n54136), .Z(n54406) );
  NOR U74531 ( .A(n54408), .B(n54406), .Z(n54138) );
  XOR U74532 ( .A(n54139), .B(n54138), .Z(n54402) );
  XOR U74533 ( .A(n54401), .B(n54402), .Z(n59381) );
  XOR U74534 ( .A(n54140), .B(n59381), .Z(n54398) );
  XOR U74535 ( .A(n54141), .B(n54398), .Z(n59726) );
  XOR U74536 ( .A(n59384), .B(n59726), .Z(n59385) );
  IV U74537 ( .A(n54142), .Z(n54144) );
  NOR U74538 ( .A(n54144), .B(n54143), .Z(n54145) );
  IV U74539 ( .A(n54145), .Z(n59386) );
  XOR U74540 ( .A(n59385), .B(n59386), .Z(n54388) );
  IV U74541 ( .A(n54146), .Z(n54147) );
  NOR U74542 ( .A(n54389), .B(n54147), .Z(n54148) );
  XOR U74543 ( .A(n54388), .B(n54148), .Z(n54386) );
  IV U74544 ( .A(n54149), .Z(n54157) );
  IV U74545 ( .A(n54150), .Z(n54151) );
  NOR U74546 ( .A(n54157), .B(n54151), .Z(n54152) );
  IV U74547 ( .A(n54152), .Z(n54385) );
  XOR U74548 ( .A(n54386), .B(n54385), .Z(n54382) );
  IV U74549 ( .A(n54153), .Z(n54154) );
  NOR U74550 ( .A(n54157), .B(n54154), .Z(n59396) );
  IV U74551 ( .A(n54155), .Z(n54156) );
  NOR U74552 ( .A(n54157), .B(n54156), .Z(n54383) );
  NOR U74553 ( .A(n59396), .B(n54383), .Z(n54158) );
  XOR U74554 ( .A(n54382), .B(n54158), .Z(n59404) );
  XOR U74555 ( .A(n59399), .B(n59404), .Z(n54380) );
  XOR U74556 ( .A(n54159), .B(n54380), .Z(n54376) );
  XOR U74557 ( .A(n54160), .B(n54376), .Z(n54374) );
  XOR U74558 ( .A(n54372), .B(n54374), .Z(n59408) );
  XOR U74559 ( .A(n59406), .B(n59408), .Z(n54369) );
  XOR U74560 ( .A(n54161), .B(n54369), .Z(n54359) );
  IV U74561 ( .A(n54162), .Z(n54163) );
  NOR U74562 ( .A(n54163), .B(n54167), .Z(n54358) );
  NOR U74563 ( .A(n54165), .B(n54164), .Z(n54363) );
  IV U74564 ( .A(n54166), .Z(n54168) );
  NOR U74565 ( .A(n54168), .B(n54167), .Z(n54361) );
  NOR U74566 ( .A(n54363), .B(n54361), .Z(n54169) );
  IV U74567 ( .A(n54169), .Z(n54170) );
  NOR U74568 ( .A(n54358), .B(n54170), .Z(n54171) );
  XOR U74569 ( .A(n54359), .B(n54171), .Z(n54357) );
  XOR U74570 ( .A(n54355), .B(n54357), .Z(n65003) );
  XOR U74571 ( .A(n54172), .B(n65003), .Z(n54345) );
  IV U74572 ( .A(n54173), .Z(n54174) );
  NOR U74573 ( .A(n54175), .B(n54174), .Z(n54348) );
  NOR U74574 ( .A(n54177), .B(n54176), .Z(n54344) );
  NOR U74575 ( .A(n54348), .B(n54344), .Z(n54178) );
  XOR U74576 ( .A(n54345), .B(n54178), .Z(n59421) );
  IV U74577 ( .A(n54179), .Z(n54181) );
  NOR U74578 ( .A(n54181), .B(n54180), .Z(n59419) );
  XOR U74579 ( .A(n59421), .B(n59419), .Z(n59424) );
  XOR U74580 ( .A(n59422), .B(n59424), .Z(n54343) );
  XOR U74581 ( .A(n54182), .B(n54343), .Z(n54334) );
  IV U74582 ( .A(n54183), .Z(n54184) );
  NOR U74583 ( .A(n54185), .B(n54184), .Z(n54336) );
  IV U74584 ( .A(n54186), .Z(n54187) );
  NOR U74585 ( .A(n54187), .B(n54323), .Z(n54333) );
  NOR U74586 ( .A(n54336), .B(n54333), .Z(n54188) );
  XOR U74587 ( .A(n54334), .B(n54188), .Z(n54324) );
  XOR U74588 ( .A(n54189), .B(n54324), .Z(n59432) );
  XOR U74589 ( .A(n59430), .B(n59432), .Z(n54320) );
  XOR U74590 ( .A(n54318), .B(n54320), .Z(n59428) );
  XOR U74591 ( .A(n59427), .B(n59428), .Z(n59439) );
  XOR U74592 ( .A(n59438), .B(n59439), .Z(n59442) );
  XOR U74593 ( .A(n59441), .B(n59442), .Z(n54316) );
  XOR U74594 ( .A(n54315), .B(n54316), .Z(n59448) );
  XOR U74595 ( .A(n59447), .B(n59448), .Z(n54309) );
  XOR U74596 ( .A(n54190), .B(n54309), .Z(n69941) );
  XOR U74597 ( .A(n54191), .B(n69941), .Z(n59467) );
  IV U74598 ( .A(n54192), .Z(n54193) );
  NOR U74599 ( .A(n54199), .B(n54193), .Z(n59466) );
  IV U74600 ( .A(n54194), .Z(n54195) );
  NOR U74601 ( .A(n54199), .B(n54195), .Z(n59458) );
  NOR U74602 ( .A(n59466), .B(n59458), .Z(n54196) );
  XOR U74603 ( .A(n59467), .B(n54196), .Z(n59465) );
  IV U74604 ( .A(n54197), .Z(n54198) );
  NOR U74605 ( .A(n54199), .B(n54198), .Z(n59463) );
  XOR U74606 ( .A(n59465), .B(n59463), .Z(n59480) );
  XOR U74607 ( .A(n54200), .B(n59480), .Z(n59474) );
  XOR U74608 ( .A(n59472), .B(n59474), .Z(n59477) );
  XOR U74609 ( .A(n59476), .B(n59477), .Z(n54302) );
  XOR U74610 ( .A(n54301), .B(n54302), .Z(n59493) );
  XOR U74611 ( .A(n59492), .B(n59493), .Z(n59497) );
  XOR U74612 ( .A(n59495), .B(n59497), .Z(n54294) );
  XOR U74613 ( .A(n54201), .B(n54294), .Z(n54292) );
  XOR U74614 ( .A(n54290), .B(n54292), .Z(n59510) );
  XOR U74615 ( .A(n59508), .B(n59510), .Z(n54286) );
  XOR U74616 ( .A(n54202), .B(n54286), .Z(n59517) );
  XOR U74617 ( .A(n59516), .B(n59517), .Z(n59520) );
  XOR U74618 ( .A(n54203), .B(n59520), .Z(n54277) );
  XOR U74619 ( .A(n54278), .B(n54277), .Z(n54282) );
  IV U74620 ( .A(n54204), .Z(n54206) );
  NOR U74621 ( .A(n54206), .B(n54205), .Z(n54280) );
  XOR U74622 ( .A(n54282), .B(n54280), .Z(n59526) );
  IV U74623 ( .A(n54207), .Z(n54210) );
  NOR U74624 ( .A(n54208), .B(n54219), .Z(n54209) );
  IV U74625 ( .A(n54209), .Z(n54212) );
  NOR U74626 ( .A(n54210), .B(n54212), .Z(n59524) );
  XOR U74627 ( .A(n59526), .B(n59524), .Z(n59529) );
  IV U74628 ( .A(n54211), .Z(n54213) );
  NOR U74629 ( .A(n54213), .B(n54212), .Z(n59527) );
  XOR U74630 ( .A(n59529), .B(n59527), .Z(n59532) );
  XOR U74631 ( .A(n59531), .B(n59532), .Z(n59536) );
  IV U74632 ( .A(n54214), .Z(n54217) );
  IV U74633 ( .A(n54215), .Z(n54216) );
  NOR U74634 ( .A(n54217), .B(n54216), .Z(n54275) );
  IV U74635 ( .A(n54218), .Z(n54220) );
  NOR U74636 ( .A(n54220), .B(n54219), .Z(n59534) );
  NOR U74637 ( .A(n54275), .B(n59534), .Z(n54221) );
  XOR U74638 ( .A(n59536), .B(n54221), .Z(n54222) );
  IV U74639 ( .A(n54222), .Z(n59539) );
  NOR U74640 ( .A(n54228), .B(n59539), .Z(n59668) );
  IV U74641 ( .A(n54223), .Z(n54224) );
  NOR U74642 ( .A(n54235), .B(n54224), .Z(n54272) );
  IV U74643 ( .A(n54225), .Z(n54227) );
  NOR U74644 ( .A(n54227), .B(n54226), .Z(n59538) );
  XOR U74645 ( .A(n59538), .B(n59539), .Z(n54273) );
  IV U74646 ( .A(n54273), .Z(n54229) );
  XOR U74647 ( .A(n54272), .B(n54229), .Z(n54231) );
  NOR U74648 ( .A(n54229), .B(n54228), .Z(n54230) );
  NOR U74649 ( .A(n54231), .B(n54230), .Z(n54232) );
  NOR U74650 ( .A(n59668), .B(n54232), .Z(n54267) );
  IV U74651 ( .A(n54233), .Z(n54234) );
  NOR U74652 ( .A(n54235), .B(n54234), .Z(n54270) );
  IV U74653 ( .A(n54236), .Z(n54237) );
  NOR U74654 ( .A(n54238), .B(n54237), .Z(n54266) );
  NOR U74655 ( .A(n54270), .B(n54266), .Z(n54239) );
  XOR U74656 ( .A(n54267), .B(n54239), .Z(n54265) );
  IV U74657 ( .A(n54240), .Z(n54241) );
  NOR U74658 ( .A(n54242), .B(n54241), .Z(n54263) );
  XOR U74659 ( .A(n54265), .B(n54263), .Z(n59549) );
  XOR U74660 ( .A(n54243), .B(n59549), .Z(n54258) );
  XOR U74661 ( .A(n54259), .B(n54258), .Z(n59556) );
  IV U74662 ( .A(n54244), .Z(n54245) );
  NOR U74663 ( .A(n54246), .B(n54245), .Z(n54247) );
  IV U74664 ( .A(n54247), .Z(n59569) );
  NOR U74665 ( .A(n54251), .B(n59569), .Z(n59574) );
  NOR U74666 ( .A(n54248), .B(n59574), .Z(n54249) );
  XOR U74667 ( .A(n59544), .B(n54249), .Z(n54250) );
  IV U74668 ( .A(n54250), .Z(n69988) );
  XOR U74669 ( .A(n54252), .B(n54251), .Z(n59568) );
  IV U74670 ( .A(n54253), .Z(n54255) );
  NOR U74671 ( .A(n54255), .B(n54254), .Z(n59570) );
  IV U74672 ( .A(n59570), .Z(n59567) );
  NOR U74673 ( .A(n59568), .B(n59567), .Z(n59599) );
  IV U74674 ( .A(n59599), .Z(n54256) );
  NOR U74675 ( .A(n69988), .B(n54256), .Z(n59557) );
  IV U74676 ( .A(n59557), .Z(n54257) );
  NOR U74677 ( .A(n59556), .B(n54257), .Z(n64832) );
  IV U74678 ( .A(n54258), .Z(n59546) );
  NOR U74679 ( .A(n59546), .B(n54259), .Z(n54260) );
  IV U74680 ( .A(n54260), .Z(n59550) );
  IV U74681 ( .A(n54261), .Z(n54262) );
  NOR U74682 ( .A(n54265), .B(n54262), .Z(n64817) );
  IV U74683 ( .A(n54263), .Z(n54264) );
  NOR U74684 ( .A(n54265), .B(n54264), .Z(n64813) );
  IV U74685 ( .A(n54266), .Z(n54269) );
  IV U74686 ( .A(n54267), .Z(n54268) );
  NOR U74687 ( .A(n54269), .B(n54268), .Z(n64820) );
  IV U74688 ( .A(n54270), .Z(n54271) );
  NOR U74689 ( .A(n54271), .B(n54273), .Z(n64808) );
  IV U74690 ( .A(n54272), .Z(n54274) );
  NOR U74691 ( .A(n54274), .B(n54273), .Z(n64805) );
  IV U74692 ( .A(n54275), .Z(n54276) );
  NOR U74693 ( .A(n59536), .B(n54276), .Z(n59670) );
  IV U74694 ( .A(n54277), .Z(n54279) );
  NOR U74695 ( .A(n54279), .B(n54278), .Z(n64917) );
  IV U74696 ( .A(n54280), .Z(n54281) );
  NOR U74697 ( .A(n54282), .B(n54281), .Z(n64910) );
  NOR U74698 ( .A(n64917), .B(n64910), .Z(n64784) );
  IV U74699 ( .A(n64784), .Z(n59523) );
  IV U74700 ( .A(n54283), .Z(n54284) );
  NOR U74701 ( .A(n59520), .B(n54284), .Z(n64780) );
  IV U74702 ( .A(n54285), .Z(n54289) );
  NOR U74703 ( .A(n54287), .B(n54286), .Z(n54288) );
  IV U74704 ( .A(n54288), .Z(n59504) );
  NOR U74705 ( .A(n54289), .B(n59504), .Z(n64775) );
  IV U74706 ( .A(n54290), .Z(n54291) );
  NOR U74707 ( .A(n54292), .B(n54291), .Z(n64769) );
  IV U74708 ( .A(n54293), .Z(n54300) );
  NOR U74709 ( .A(n54295), .B(n54294), .Z(n54296) );
  IV U74710 ( .A(n54296), .Z(n54297) );
  NOR U74711 ( .A(n54298), .B(n54297), .Z(n54299) );
  IV U74712 ( .A(n54299), .Z(n59501) );
  NOR U74713 ( .A(n54300), .B(n59501), .Z(n64765) );
  IV U74714 ( .A(n54301), .Z(n54303) );
  NOR U74715 ( .A(n54303), .B(n54302), .Z(n54304) );
  IV U74716 ( .A(n54304), .Z(n64754) );
  IV U74717 ( .A(n54305), .Z(n54306) );
  NOR U74718 ( .A(n69941), .B(n54306), .Z(n64728) );
  IV U74719 ( .A(n59460), .Z(n54307) );
  XOR U74720 ( .A(n59453), .B(n69941), .Z(n59459) );
  NOR U74721 ( .A(n54307), .B(n59459), .Z(n59686) );
  IV U74722 ( .A(n54308), .Z(n54311) );
  NOR U74723 ( .A(n69928), .B(n54309), .Z(n54310) );
  IV U74724 ( .A(n54310), .Z(n54313) );
  NOR U74725 ( .A(n54311), .B(n54313), .Z(n54312) );
  IV U74726 ( .A(n54312), .Z(n64725) );
  NOR U74727 ( .A(n54314), .B(n54313), .Z(n59451) );
  IV U74728 ( .A(n59451), .Z(n59446) );
  IV U74729 ( .A(n54315), .Z(n54317) );
  NOR U74730 ( .A(n54317), .B(n54316), .Z(n64711) );
  IV U74731 ( .A(n54318), .Z(n54319) );
  NOR U74732 ( .A(n54320), .B(n54319), .Z(n54321) );
  IV U74733 ( .A(n54321), .Z(n59433) );
  IV U74734 ( .A(n54322), .Z(n54329) );
  NOR U74735 ( .A(n54324), .B(n54323), .Z(n54325) );
  IV U74736 ( .A(n54325), .Z(n54326) );
  NOR U74737 ( .A(n54327), .B(n54326), .Z(n54328) );
  IV U74738 ( .A(n54328), .Z(n54331) );
  NOR U74739 ( .A(n54329), .B(n54331), .Z(n64702) );
  IV U74740 ( .A(n54330), .Z(n54332) );
  NOR U74741 ( .A(n54332), .B(n54331), .Z(n59696) );
  IV U74742 ( .A(n54333), .Z(n54335) );
  IV U74743 ( .A(n54334), .Z(n54337) );
  NOR U74744 ( .A(n54335), .B(n54337), .Z(n64690) );
  IV U74745 ( .A(n54336), .Z(n54338) );
  NOR U74746 ( .A(n54338), .B(n54337), .Z(n59699) );
  IV U74747 ( .A(n54339), .Z(n54340) );
  NOR U74748 ( .A(n54340), .B(n54343), .Z(n64693) );
  IV U74749 ( .A(n54341), .Z(n54342) );
  NOR U74750 ( .A(n54343), .B(n54342), .Z(n64686) );
  IV U74751 ( .A(n54344), .Z(n54347) );
  IV U74752 ( .A(n54345), .Z(n54346) );
  NOR U74753 ( .A(n54347), .B(n54346), .Z(n64678) );
  IV U74754 ( .A(n54348), .Z(n54350) );
  XOR U74755 ( .A(n54353), .B(n65003), .Z(n54349) );
  NOR U74756 ( .A(n54350), .B(n54349), .Z(n64674) );
  IV U74757 ( .A(n54351), .Z(n54352) );
  NOR U74758 ( .A(n54352), .B(n65003), .Z(n64671) );
  IV U74759 ( .A(n54353), .Z(n54354) );
  NOR U74760 ( .A(n54354), .B(n65003), .Z(n64666) );
  IV U74761 ( .A(n54355), .Z(n54356) );
  NOR U74762 ( .A(n54357), .B(n54356), .Z(n69894) );
  IV U74763 ( .A(n54358), .Z(n54360) );
  IV U74764 ( .A(n54359), .Z(n54364) );
  NOR U74765 ( .A(n54360), .B(n54364), .Z(n69889) );
  NOR U74766 ( .A(n69894), .B(n69889), .Z(n64665) );
  IV U74767 ( .A(n54361), .Z(n54362) );
  NOR U74768 ( .A(n54362), .B(n54364), .Z(n64662) );
  IV U74769 ( .A(n54363), .Z(n54365) );
  NOR U74770 ( .A(n54365), .B(n54364), .Z(n64659) );
  IV U74771 ( .A(n54366), .Z(n54367) );
  NOR U74772 ( .A(n54369), .B(n54367), .Z(n59706) );
  IV U74773 ( .A(n54368), .Z(n54370) );
  NOR U74774 ( .A(n54370), .B(n54369), .Z(n59705) );
  XOR U74775 ( .A(n59706), .B(n59705), .Z(n54371) );
  NOR U74776 ( .A(n64659), .B(n54371), .Z(n59417) );
  IV U74777 ( .A(n54372), .Z(n54373) );
  NOR U74778 ( .A(n54374), .B(n54373), .Z(n54375) );
  IV U74779 ( .A(n54375), .Z(n59412) );
  IV U74780 ( .A(n54376), .Z(n59411) );
  IV U74781 ( .A(n54377), .Z(n54378) );
  NOR U74782 ( .A(n59411), .B(n54378), .Z(n64638) );
  IV U74783 ( .A(n54379), .Z(n54381) );
  NOR U74784 ( .A(n54381), .B(n54380), .Z(n59715) );
  IV U74785 ( .A(n54382), .Z(n59397) );
  IV U74786 ( .A(n54383), .Z(n54384) );
  NOR U74787 ( .A(n59397), .B(n54384), .Z(n64625) );
  NOR U74788 ( .A(n54386), .B(n54385), .Z(n59718) );
  IV U74789 ( .A(n54387), .Z(n54394) );
  NOR U74790 ( .A(n54389), .B(n54388), .Z(n54390) );
  IV U74791 ( .A(n54390), .Z(n54391) );
  NOR U74792 ( .A(n54392), .B(n54391), .Z(n54393) );
  IV U74793 ( .A(n54393), .Z(n54396) );
  NOR U74794 ( .A(n54394), .B(n54396), .Z(n64621) );
  NOR U74795 ( .A(n59718), .B(n64621), .Z(n59395) );
  IV U74796 ( .A(n54395), .Z(n54397) );
  NOR U74797 ( .A(n54397), .B(n54396), .Z(n59390) );
  IV U74798 ( .A(n54398), .Z(n59379) );
  IV U74799 ( .A(n54399), .Z(n54400) );
  NOR U74800 ( .A(n59379), .B(n54400), .Z(n64616) );
  IV U74801 ( .A(n54401), .Z(n54403) );
  NOR U74802 ( .A(n54403), .B(n54402), .Z(n69832) );
  IV U74803 ( .A(n54404), .Z(n54405) );
  NOR U74804 ( .A(n54405), .B(n59381), .Z(n65036) );
  NOR U74805 ( .A(n69832), .B(n65036), .Z(n64609) );
  IV U74806 ( .A(n54406), .Z(n54407) );
  NOR U74807 ( .A(n54407), .B(n54409), .Z(n64606) );
  IV U74808 ( .A(n54408), .Z(n54410) );
  NOR U74809 ( .A(n54410), .B(n54409), .Z(n54411) );
  IV U74810 ( .A(n54411), .Z(n64603) );
  IV U74811 ( .A(n54412), .Z(n54417) );
  IV U74812 ( .A(n54413), .Z(n54414) );
  NOR U74813 ( .A(n54417), .B(n54414), .Z(n59741) );
  IV U74814 ( .A(n54415), .Z(n54416) );
  NOR U74815 ( .A(n54417), .B(n54416), .Z(n59738) );
  IV U74816 ( .A(n54418), .Z(n54419) );
  NOR U74817 ( .A(n54424), .B(n54419), .Z(n59743) );
  IV U74818 ( .A(n54420), .Z(n54421) );
  NOR U74819 ( .A(n54421), .B(n59749), .Z(n54425) );
  IV U74820 ( .A(n54422), .Z(n54423) );
  NOR U74821 ( .A(n54424), .B(n54423), .Z(n59746) );
  NOR U74822 ( .A(n54425), .B(n59746), .Z(n59361) );
  IV U74823 ( .A(n54426), .Z(n59758) );
  NOR U74824 ( .A(n54427), .B(n59758), .Z(n54434) );
  IV U74825 ( .A(n54428), .Z(n54429) );
  NOR U74826 ( .A(n54429), .B(n54432), .Z(n64583) );
  IV U74827 ( .A(n54430), .Z(n54431) );
  NOR U74828 ( .A(n54432), .B(n54431), .Z(n64581) );
  XOR U74829 ( .A(n64583), .B(n64581), .Z(n54433) );
  NOR U74830 ( .A(n54434), .B(n54433), .Z(n59360) );
  IV U74831 ( .A(n54435), .Z(n54436) );
  NOR U74832 ( .A(n54437), .B(n54436), .Z(n64577) );
  IV U74833 ( .A(n54438), .Z(n54444) );
  XOR U74834 ( .A(n54452), .B(n54453), .Z(n54449) );
  NOR U74835 ( .A(n54439), .B(n54449), .Z(n54440) );
  IV U74836 ( .A(n54440), .Z(n54441) );
  NOR U74837 ( .A(n54442), .B(n54441), .Z(n54443) );
  IV U74838 ( .A(n54443), .Z(n54446) );
  NOR U74839 ( .A(n54444), .B(n54446), .Z(n64569) );
  NOR U74840 ( .A(n64577), .B(n64569), .Z(n59359) );
  IV U74841 ( .A(n54445), .Z(n54447) );
  NOR U74842 ( .A(n54447), .B(n54446), .Z(n59764) );
  IV U74843 ( .A(n54448), .Z(n54450) );
  NOR U74844 ( .A(n54450), .B(n54449), .Z(n64564) );
  IV U74845 ( .A(n54451), .Z(n70166) );
  NOR U74846 ( .A(n70166), .B(n54459), .Z(n64557) );
  IV U74847 ( .A(n54452), .Z(n54454) );
  NOR U74848 ( .A(n54454), .B(n54453), .Z(n59769) );
  NOR U74849 ( .A(n64557), .B(n59769), .Z(n59358) );
  IV U74850 ( .A(n54455), .Z(n54456) );
  NOR U74851 ( .A(n54457), .B(n54456), .Z(n59774) );
  IV U74852 ( .A(n54458), .Z(n70170) );
  NOR U74853 ( .A(n70170), .B(n54459), .Z(n64559) );
  NOR U74854 ( .A(n59774), .B(n64559), .Z(n59357) );
  IV U74855 ( .A(n54460), .Z(n54461) );
  NOR U74856 ( .A(n54462), .B(n54461), .Z(n59772) );
  IV U74857 ( .A(n54463), .Z(n54464) );
  NOR U74858 ( .A(n54469), .B(n54464), .Z(n59776) );
  NOR U74859 ( .A(n59772), .B(n59776), .Z(n59356) );
  IV U74860 ( .A(n54465), .Z(n54467) );
  NOR U74861 ( .A(n54467), .B(n54466), .Z(n64553) );
  IV U74862 ( .A(n54468), .Z(n54470) );
  NOR U74863 ( .A(n54470), .B(n54469), .Z(n59779) );
  NOR U74864 ( .A(n64553), .B(n59779), .Z(n59355) );
  IV U74865 ( .A(n54471), .Z(n54473) );
  NOR U74866 ( .A(n54473), .B(n54472), .Z(n64551) );
  IV U74867 ( .A(n54474), .Z(n54475) );
  NOR U74868 ( .A(n54475), .B(n54483), .Z(n59787) );
  IV U74869 ( .A(n54476), .Z(n54478) );
  NOR U74870 ( .A(n54478), .B(n54477), .Z(n59784) );
  NOR U74871 ( .A(n59787), .B(n59784), .Z(n59354) );
  IV U74872 ( .A(n54479), .Z(n54481) );
  NOR U74873 ( .A(n54481), .B(n54480), .Z(n59793) );
  IV U74874 ( .A(n54482), .Z(n54484) );
  NOR U74875 ( .A(n54484), .B(n54483), .Z(n59790) );
  NOR U74876 ( .A(n59793), .B(n59790), .Z(n59353) );
  IV U74877 ( .A(n54485), .Z(n54487) );
  NOR U74878 ( .A(n54487), .B(n54486), .Z(n64546) );
  NOR U74879 ( .A(n54489), .B(n54488), .Z(n64543) );
  IV U74880 ( .A(n54490), .Z(n54491) );
  NOR U74881 ( .A(n54492), .B(n54491), .Z(n64531) );
  IV U74882 ( .A(n54493), .Z(n54494) );
  NOR U74883 ( .A(n54494), .B(n59341), .Z(n59795) );
  IV U74884 ( .A(n54495), .Z(n54500) );
  IV U74885 ( .A(n54496), .Z(n54497) );
  NOR U74886 ( .A(n54500), .B(n54497), .Z(n64523) );
  NOR U74887 ( .A(n59795), .B(n64523), .Z(n59339) );
  IV U74888 ( .A(n54498), .Z(n54499) );
  NOR U74889 ( .A(n54500), .B(n54499), .Z(n64526) );
  IV U74890 ( .A(n54501), .Z(n54502) );
  NOR U74891 ( .A(n54508), .B(n54502), .Z(n59801) );
  NOR U74892 ( .A(n64526), .B(n59801), .Z(n59338) );
  IV U74893 ( .A(n54503), .Z(n54504) );
  NOR U74894 ( .A(n54505), .B(n54504), .Z(n59806) );
  IV U74895 ( .A(n54506), .Z(n54507) );
  NOR U74896 ( .A(n54508), .B(n54507), .Z(n59803) );
  NOR U74897 ( .A(n59806), .B(n59803), .Z(n59337) );
  IV U74898 ( .A(n54509), .Z(n54511) );
  NOR U74899 ( .A(n54511), .B(n54510), .Z(n59808) );
  IV U74900 ( .A(n54512), .Z(n54513) );
  NOR U74901 ( .A(n54514), .B(n54513), .Z(n54515) );
  IV U74902 ( .A(n54515), .Z(n59321) );
  NOR U74903 ( .A(n54516), .B(n59832), .Z(n54519) );
  IV U74904 ( .A(n54517), .Z(n54518) );
  NOR U74905 ( .A(n54518), .B(n59315), .Z(n59821) );
  NOR U74906 ( .A(n54519), .B(n59821), .Z(n59311) );
  IV U74907 ( .A(n54520), .Z(n54522) );
  NOR U74908 ( .A(n54522), .B(n54521), .Z(n59299) );
  NOR U74909 ( .A(n54524), .B(n54523), .Z(n54525) );
  IV U74910 ( .A(n54525), .Z(n54526) );
  NOR U74911 ( .A(n54527), .B(n54526), .Z(n54528) );
  IV U74912 ( .A(n54528), .Z(n59840) );
  NOR U74913 ( .A(n54529), .B(n59840), .Z(n59290) );
  IV U74914 ( .A(n54530), .Z(n54531) );
  NOR U74915 ( .A(n54531), .B(n54536), .Z(n65116) );
  IV U74916 ( .A(n54532), .Z(n54533) );
  NOR U74917 ( .A(n54534), .B(n54533), .Z(n59844) );
  NOR U74918 ( .A(n65116), .B(n59844), .Z(n59288) );
  IV U74919 ( .A(n54535), .Z(n54537) );
  NOR U74920 ( .A(n54537), .B(n54536), .Z(n65120) );
  IV U74921 ( .A(n54538), .Z(n54540) );
  IV U74922 ( .A(n54539), .Z(n54549) );
  NOR U74923 ( .A(n54540), .B(n54549), .Z(n59848) );
  IV U74924 ( .A(n54541), .Z(n54542) );
  NOR U74925 ( .A(n54542), .B(n54544), .Z(n59854) );
  IV U74926 ( .A(n54543), .Z(n54545) );
  NOR U74927 ( .A(n54545), .B(n54544), .Z(n59856) );
  NOR U74928 ( .A(n59854), .B(n59856), .Z(n54546) );
  IV U74929 ( .A(n54546), .Z(n54550) );
  IV U74930 ( .A(n54547), .Z(n54548) );
  NOR U74931 ( .A(n54549), .B(n54548), .Z(n59852) );
  NOR U74932 ( .A(n54550), .B(n59852), .Z(n59287) );
  IV U74933 ( .A(n54551), .Z(n54552) );
  NOR U74934 ( .A(n54553), .B(n54552), .Z(n64492) );
  IV U74935 ( .A(n54554), .Z(n54556) );
  NOR U74936 ( .A(n54556), .B(n54555), .Z(n64495) );
  NOR U74937 ( .A(n64492), .B(n64495), .Z(n59286) );
  IV U74938 ( .A(n54557), .Z(n54559) );
  XOR U74939 ( .A(n54565), .B(n54567), .Z(n54558) );
  NOR U74940 ( .A(n54559), .B(n54558), .Z(n54560) );
  IV U74941 ( .A(n54560), .Z(n54561) );
  NOR U74942 ( .A(n54566), .B(n54561), .Z(n64489) );
  IV U74943 ( .A(n54562), .Z(n54563) );
  NOR U74944 ( .A(n54564), .B(n54563), .Z(n64484) );
  IV U74945 ( .A(n54565), .Z(n54570) );
  NOR U74946 ( .A(n54567), .B(n54566), .Z(n54568) );
  IV U74947 ( .A(n54568), .Z(n54569) );
  NOR U74948 ( .A(n54570), .B(n54569), .Z(n64486) );
  NOR U74949 ( .A(n64484), .B(n64486), .Z(n59285) );
  IV U74950 ( .A(n54571), .Z(n54573) );
  NOR U74951 ( .A(n54573), .B(n54572), .Z(n59859) );
  NOR U74952 ( .A(n59864), .B(n59859), .Z(n59284) );
  IV U74953 ( .A(n54574), .Z(n54575) );
  NOR U74954 ( .A(n54578), .B(n54575), .Z(n69664) );
  IV U74955 ( .A(n54576), .Z(n54577) );
  NOR U74956 ( .A(n54578), .B(n54577), .Z(n65147) );
  NOR U74957 ( .A(n69664), .B(n65147), .Z(n59863) );
  IV U74958 ( .A(n54579), .Z(n54581) );
  NOR U74959 ( .A(n54581), .B(n54580), .Z(n59226) );
  IV U74960 ( .A(n59226), .Z(n59224) );
  IV U74961 ( .A(n54582), .Z(n54583) );
  NOR U74962 ( .A(n54584), .B(n54583), .Z(n54585) );
  IV U74963 ( .A(n54585), .Z(n64441) );
  IV U74964 ( .A(n54586), .Z(n54587) );
  NOR U74965 ( .A(n54587), .B(n54592), .Z(n64437) );
  IV U74966 ( .A(n54588), .Z(n54589) );
  NOR U74967 ( .A(n54590), .B(n54589), .Z(n59898) );
  IV U74968 ( .A(n54591), .Z(n54593) );
  NOR U74969 ( .A(n54593), .B(n54592), .Z(n59896) );
  NOR U74970 ( .A(n59898), .B(n59896), .Z(n59211) );
  IV U74971 ( .A(n54594), .Z(n54595) );
  NOR U74972 ( .A(n54595), .B(n54598), .Z(n64433) );
  IV U74973 ( .A(n54596), .Z(n54597) );
  NOR U74974 ( .A(n54598), .B(n54597), .Z(n64430) );
  IV U74975 ( .A(n54599), .Z(n54601) );
  NOR U74976 ( .A(n54601), .B(n54600), .Z(n59916) );
  IV U74977 ( .A(n54602), .Z(n54603) );
  NOR U74978 ( .A(n54604), .B(n54603), .Z(n59913) );
  NOR U74979 ( .A(n59916), .B(n59913), .Z(n59170) );
  IV U74980 ( .A(n54605), .Z(n54606) );
  NOR U74981 ( .A(n54606), .B(n54611), .Z(n59921) );
  IV U74982 ( .A(n54607), .Z(n54609) );
  NOR U74983 ( .A(n54609), .B(n54608), .Z(n64384) );
  IV U74984 ( .A(n54610), .Z(n54612) );
  NOR U74985 ( .A(n54612), .B(n54611), .Z(n64388) );
  NOR U74986 ( .A(n64384), .B(n64388), .Z(n59161) );
  IV U74987 ( .A(n54613), .Z(n54618) );
  IV U74988 ( .A(n54614), .Z(n54615) );
  NOR U74989 ( .A(n54618), .B(n54615), .Z(n59928) );
  IV U74990 ( .A(n54616), .Z(n54617) );
  NOR U74991 ( .A(n54618), .B(n54617), .Z(n59925) );
  IV U74992 ( .A(n54619), .Z(n54620) );
  NOR U74993 ( .A(n54620), .B(n54622), .Z(n59934) );
  IV U74994 ( .A(n54621), .Z(n54623) );
  NOR U74995 ( .A(n54623), .B(n54622), .Z(n59931) );
  IV U74996 ( .A(n54624), .Z(n54628) );
  NOR U74997 ( .A(n54626), .B(n54625), .Z(n54627) );
  IV U74998 ( .A(n54627), .Z(n59159) );
  NOR U74999 ( .A(n54628), .B(n59159), .Z(n64379) );
  IV U75000 ( .A(n54629), .Z(n54631) );
  NOR U75001 ( .A(n54631), .B(n54630), .Z(n59950) );
  IV U75002 ( .A(n54632), .Z(n54634) );
  NOR U75003 ( .A(n54634), .B(n54633), .Z(n59957) );
  IV U75004 ( .A(n54635), .Z(n54639) );
  NOR U75005 ( .A(n54637), .B(n54636), .Z(n54638) );
  IV U75006 ( .A(n54638), .Z(n59117) );
  NOR U75007 ( .A(n54639), .B(n59117), .Z(n64355) );
  NOR U75008 ( .A(n54640), .B(n59110), .Z(n54641) );
  IV U75009 ( .A(n54641), .Z(n54642) );
  NOR U75010 ( .A(n54643), .B(n54642), .Z(n59981) );
  IV U75011 ( .A(n54644), .Z(n54645) );
  NOR U75012 ( .A(n54646), .B(n54645), .Z(n59978) );
  IV U75013 ( .A(n54647), .Z(n54650) );
  IV U75014 ( .A(n54648), .Z(n59105) );
  XOR U75015 ( .A(n54655), .B(n59105), .Z(n54649) );
  NOR U75016 ( .A(n54650), .B(n54649), .Z(n54651) );
  IV U75017 ( .A(n54651), .Z(n54652) );
  NOR U75018 ( .A(n54653), .B(n54652), .Z(n59984) );
  XOR U75019 ( .A(n54654), .B(n54653), .Z(n54659) );
  IV U75020 ( .A(n54655), .Z(n54656) );
  NOR U75021 ( .A(n54656), .B(n59105), .Z(n54657) );
  IV U75022 ( .A(n54657), .Z(n54658) );
  NOR U75023 ( .A(n54659), .B(n54658), .Z(n64349) );
  NOR U75024 ( .A(n59984), .B(n64349), .Z(n54660) );
  IV U75025 ( .A(n54660), .Z(n59102) );
  IV U75026 ( .A(n54661), .Z(n54663) );
  NOR U75027 ( .A(n54663), .B(n54662), .Z(n59990) );
  NOR U75028 ( .A(n54665), .B(n54664), .Z(n64346) );
  NOR U75029 ( .A(n59990), .B(n64346), .Z(n59101) );
  IV U75030 ( .A(n54666), .Z(n54667) );
  NOR U75031 ( .A(n54668), .B(n54667), .Z(n64335) );
  NOR U75032 ( .A(n54669), .B(n64340), .Z(n54670) );
  NOR U75033 ( .A(n64335), .B(n54670), .Z(n59100) );
  IV U75034 ( .A(n54671), .Z(n54676) );
  IV U75035 ( .A(n54672), .Z(n54673) );
  NOR U75036 ( .A(n54676), .B(n54673), .Z(n59992) );
  IV U75037 ( .A(n54674), .Z(n54675) );
  NOR U75038 ( .A(n54676), .B(n54675), .Z(n64328) );
  IV U75039 ( .A(n54677), .Z(n54678) );
  NOR U75040 ( .A(n54678), .B(n54684), .Z(n59996) );
  NOR U75041 ( .A(n64328), .B(n59996), .Z(n59099) );
  IV U75042 ( .A(n54679), .Z(n54681) );
  NOR U75043 ( .A(n54681), .B(n54680), .Z(n64311) );
  IV U75044 ( .A(n54682), .Z(n54683) );
  NOR U75045 ( .A(n54684), .B(n54683), .Z(n64323) );
  NOR U75046 ( .A(n64311), .B(n64323), .Z(n59098) );
  IV U75047 ( .A(n54685), .Z(n54686) );
  NOR U75048 ( .A(n54687), .B(n54686), .Z(n64315) );
  IV U75049 ( .A(n54688), .Z(n54689) );
  NOR U75050 ( .A(n54689), .B(n59095), .Z(n54690) );
  IV U75051 ( .A(n54690), .Z(n60000) );
  IV U75052 ( .A(n54691), .Z(n54697) );
  IV U75053 ( .A(n54692), .Z(n54693) );
  NOR U75054 ( .A(n54697), .B(n54693), .Z(n54694) );
  IV U75055 ( .A(n54694), .Z(n64306) );
  IV U75056 ( .A(n54695), .Z(n54696) );
  NOR U75057 ( .A(n54697), .B(n54696), .Z(n60004) );
  IV U75058 ( .A(n54698), .Z(n54699) );
  NOR U75059 ( .A(n54699), .B(n54701), .Z(n60006) );
  NOR U75060 ( .A(n60004), .B(n60006), .Z(n59090) );
  IV U75061 ( .A(n54700), .Z(n54702) );
  NOR U75062 ( .A(n54702), .B(n54701), .Z(n64293) );
  NOR U75063 ( .A(n54704), .B(n54703), .Z(n54705) );
  IV U75064 ( .A(n54705), .Z(n54706) );
  NOR U75065 ( .A(n54707), .B(n54706), .Z(n54708) );
  IV U75066 ( .A(n54708), .Z(n64299) );
  IV U75067 ( .A(n54709), .Z(n54715) );
  NOR U75068 ( .A(n54710), .B(n54715), .Z(n54711) );
  IV U75069 ( .A(n54711), .Z(n54712) );
  NOR U75070 ( .A(n54713), .B(n54712), .Z(n64289) );
  IV U75071 ( .A(n54714), .Z(n54716) );
  NOR U75072 ( .A(n54716), .B(n54715), .Z(n64286) );
  NOR U75073 ( .A(n54718), .B(n54717), .Z(n64281) );
  IV U75074 ( .A(n54719), .Z(n54720) );
  NOR U75075 ( .A(n54720), .B(n59073), .Z(n69483) );
  NOR U75076 ( .A(n69483), .B(n64280), .Z(n59083) );
  IV U75077 ( .A(n54721), .Z(n54726) );
  IV U75078 ( .A(n54722), .Z(n54723) );
  NOR U75079 ( .A(n54723), .B(n59073), .Z(n54724) );
  IV U75080 ( .A(n54724), .Z(n54725) );
  NOR U75081 ( .A(n54726), .B(n54725), .Z(n64275) );
  IV U75082 ( .A(n54727), .Z(n54728) );
  NOR U75083 ( .A(n54729), .B(n54728), .Z(n60017) );
  IV U75084 ( .A(n54730), .Z(n54731) );
  NOR U75085 ( .A(n54732), .B(n54731), .Z(n60015) );
  NOR U75086 ( .A(n60017), .B(n60015), .Z(n59070) );
  IV U75087 ( .A(n54733), .Z(n54734) );
  NOR U75088 ( .A(n54735), .B(n54734), .Z(n60023) );
  IV U75089 ( .A(n54736), .Z(n54738) );
  NOR U75090 ( .A(n54738), .B(n54737), .Z(n60021) );
  NOR U75091 ( .A(n60023), .B(n60021), .Z(n59069) );
  IV U75092 ( .A(n54739), .Z(n54740) );
  NOR U75093 ( .A(n54741), .B(n54740), .Z(n64272) );
  IV U75094 ( .A(n54742), .Z(n54744) );
  NOR U75095 ( .A(n54744), .B(n54743), .Z(n60030) );
  NOR U75096 ( .A(n64272), .B(n60030), .Z(n59068) );
  IV U75097 ( .A(n54745), .Z(n54746) );
  NOR U75098 ( .A(n54746), .B(n54748), .Z(n60028) );
  IV U75099 ( .A(n54747), .Z(n54749) );
  NOR U75100 ( .A(n54749), .B(n54748), .Z(n54750) );
  IV U75101 ( .A(n54750), .Z(n60034) );
  IV U75102 ( .A(n54751), .Z(n54752) );
  NOR U75103 ( .A(n54752), .B(n59048), .Z(n60050) );
  IV U75104 ( .A(n54753), .Z(n54754) );
  NOR U75105 ( .A(n54755), .B(n54754), .Z(n54756) );
  IV U75106 ( .A(n54756), .Z(n59052) );
  IV U75107 ( .A(n54757), .Z(n54758) );
  NOR U75108 ( .A(n54759), .B(n54758), .Z(n64256) );
  IV U75109 ( .A(n54760), .Z(n54763) );
  NOR U75110 ( .A(n54761), .B(n54763), .Z(n60062) );
  IV U75111 ( .A(n54762), .Z(n54764) );
  NOR U75112 ( .A(n54764), .B(n54763), .Z(n60060) );
  NOR U75113 ( .A(n60062), .B(n60060), .Z(n59037) );
  IV U75114 ( .A(n54765), .Z(n54767) );
  NOR U75115 ( .A(n54767), .B(n54766), .Z(n60074) );
  IV U75116 ( .A(n54768), .Z(n54769) );
  NOR U75117 ( .A(n54769), .B(n59032), .Z(n64251) );
  NOR U75118 ( .A(n60074), .B(n64251), .Z(n69435) );
  IV U75119 ( .A(n54770), .Z(n60078) );
  IV U75120 ( .A(n54771), .Z(n54772) );
  NOR U75121 ( .A(n60078), .B(n54772), .Z(n60072) );
  IV U75122 ( .A(n54773), .Z(n54774) );
  NOR U75123 ( .A(n54775), .B(n54774), .Z(n64246) );
  IV U75124 ( .A(n54776), .Z(n54783) );
  NOR U75125 ( .A(n54778), .B(n54777), .Z(n54779) );
  IV U75126 ( .A(n54779), .Z(n54780) );
  NOR U75127 ( .A(n54781), .B(n54780), .Z(n54782) );
  IV U75128 ( .A(n54782), .Z(n59019) );
  NOR U75129 ( .A(n54783), .B(n59019), .Z(n64241) );
  NOR U75130 ( .A(n64246), .B(n64241), .Z(n59022) );
  IV U75131 ( .A(n54784), .Z(n54785) );
  NOR U75132 ( .A(n54785), .B(n54787), .Z(n60092) );
  IV U75133 ( .A(n54786), .Z(n54788) );
  NOR U75134 ( .A(n54788), .B(n54787), .Z(n60089) );
  NOR U75135 ( .A(n60092), .B(n60089), .Z(n59017) );
  IV U75136 ( .A(n54789), .Z(n54796) );
  NOR U75137 ( .A(n54791), .B(n54790), .Z(n54792) );
  IV U75138 ( .A(n54792), .Z(n54793) );
  NOR U75139 ( .A(n54794), .B(n54793), .Z(n54795) );
  IV U75140 ( .A(n54795), .Z(n54798) );
  NOR U75141 ( .A(n54796), .B(n54798), .Z(n60105) );
  IV U75142 ( .A(n54797), .Z(n54799) );
  NOR U75143 ( .A(n54799), .B(n54798), .Z(n60114) );
  NOR U75144 ( .A(n54801), .B(n54800), .Z(n54802) );
  IV U75145 ( .A(n54802), .Z(n75821) );
  NOR U75146 ( .A(n54803), .B(n75821), .Z(n58970) );
  IV U75147 ( .A(n58970), .Z(n58964) );
  IV U75148 ( .A(n54804), .Z(n54805) );
  NOR U75149 ( .A(n54806), .B(n54805), .Z(n60131) );
  IV U75150 ( .A(n54807), .Z(n54812) );
  IV U75151 ( .A(n54808), .Z(n54809) );
  NOR U75152 ( .A(n54812), .B(n54809), .Z(n60128) );
  IV U75153 ( .A(n54810), .Z(n54811) );
  NOR U75154 ( .A(n54812), .B(n54811), .Z(n60134) );
  IV U75155 ( .A(n54813), .Z(n54816) );
  IV U75156 ( .A(n54814), .Z(n54815) );
  NOR U75157 ( .A(n54816), .B(n54815), .Z(n60155) );
  NOR U75158 ( .A(n60158), .B(n60155), .Z(n58942) );
  IV U75159 ( .A(n54817), .Z(n54818) );
  NOR U75160 ( .A(n54819), .B(n54818), .Z(n60159) );
  IV U75161 ( .A(n54820), .Z(n54827) );
  NOR U75162 ( .A(n54822), .B(n54821), .Z(n54823) );
  IV U75163 ( .A(n54823), .Z(n54824) );
  NOR U75164 ( .A(n54825), .B(n54824), .Z(n54826) );
  IV U75165 ( .A(n54826), .Z(n54829) );
  NOR U75166 ( .A(n54827), .B(n54829), .Z(n64183) );
  IV U75167 ( .A(n54828), .Z(n54830) );
  NOR U75168 ( .A(n54830), .B(n54829), .Z(n64180) );
  IV U75169 ( .A(n54831), .Z(n54836) );
  NOR U75170 ( .A(n54838), .B(n54832), .Z(n54833) );
  IV U75171 ( .A(n54833), .Z(n60166) );
  NOR U75172 ( .A(n54834), .B(n60166), .Z(n54835) );
  IV U75173 ( .A(n54835), .Z(n54840) );
  NOR U75174 ( .A(n54836), .B(n54840), .Z(n60172) );
  NOR U75175 ( .A(n54838), .B(n54837), .Z(n60181) );
  IV U75176 ( .A(n54839), .Z(n54841) );
  NOR U75177 ( .A(n54841), .B(n54840), .Z(n60175) );
  NOR U75178 ( .A(n60181), .B(n60175), .Z(n58928) );
  IV U75179 ( .A(n54842), .Z(n54844) );
  IV U75180 ( .A(n54843), .Z(n54846) );
  NOR U75181 ( .A(n54844), .B(n54846), .Z(n60178) );
  IV U75182 ( .A(n54845), .Z(n54847) );
  NOR U75183 ( .A(n54847), .B(n54846), .Z(n60187) );
  IV U75184 ( .A(n54848), .Z(n54849) );
  NOR U75185 ( .A(n54849), .B(n58926), .Z(n54850) );
  IV U75186 ( .A(n54850), .Z(n60185) );
  IV U75187 ( .A(n54851), .Z(n54853) );
  NOR U75188 ( .A(n54853), .B(n54852), .Z(n64161) );
  IV U75189 ( .A(n54854), .Z(n54857) );
  NOR U75190 ( .A(n54855), .B(n58916), .Z(n54856) );
  IV U75191 ( .A(n54856), .Z(n54859) );
  NOR U75192 ( .A(n54857), .B(n54859), .Z(n64156) );
  IV U75193 ( .A(n54858), .Z(n54860) );
  NOR U75194 ( .A(n54860), .B(n54859), .Z(n64157) );
  XOR U75195 ( .A(n64156), .B(n64157), .Z(n54861) );
  NOR U75196 ( .A(n64161), .B(n54861), .Z(n58914) );
  IV U75197 ( .A(n54862), .Z(n54865) );
  NOR U75198 ( .A(n54869), .B(n54863), .Z(n54864) );
  IV U75199 ( .A(n54864), .Z(n54871) );
  NOR U75200 ( .A(n54865), .B(n54871), .Z(n54866) );
  IV U75201 ( .A(n54866), .Z(n64144) );
  IV U75202 ( .A(n54867), .Z(n54868) );
  NOR U75203 ( .A(n54869), .B(n54868), .Z(n65499) );
  IV U75204 ( .A(n54870), .Z(n54872) );
  NOR U75205 ( .A(n54872), .B(n54871), .Z(n65490) );
  NOR U75206 ( .A(n65499), .B(n65490), .Z(n60191) );
  IV U75207 ( .A(n54873), .Z(n54875) );
  NOR U75208 ( .A(n54875), .B(n54874), .Z(n65512) );
  IV U75209 ( .A(n54876), .Z(n54877) );
  NOR U75210 ( .A(n54878), .B(n54877), .Z(n65508) );
  NOR U75211 ( .A(n65512), .B(n65508), .Z(n64133) );
  IV U75212 ( .A(n54879), .Z(n54881) );
  NOR U75213 ( .A(n54881), .B(n54880), .Z(n60198) );
  IV U75214 ( .A(n54882), .Z(n64129) );
  IV U75215 ( .A(n54883), .Z(n54885) );
  NOR U75216 ( .A(n54885), .B(n54884), .Z(n60211) );
  IV U75217 ( .A(n54886), .Z(n54888) );
  NOR U75218 ( .A(n54888), .B(n54887), .Z(n60205) );
  NOR U75219 ( .A(n60211), .B(n60205), .Z(n58892) );
  IV U75220 ( .A(n54889), .Z(n54892) );
  IV U75221 ( .A(n54890), .Z(n54896) );
  XOR U75222 ( .A(n54896), .B(n54893), .Z(n54891) );
  NOR U75223 ( .A(n54892), .B(n54891), .Z(n64124) );
  IV U75224 ( .A(n54893), .Z(n54897) );
  IV U75225 ( .A(n54894), .Z(n54895) );
  NOR U75226 ( .A(n54897), .B(n54895), .Z(n64121) );
  NOR U75227 ( .A(n54897), .B(n54896), .Z(n60220) );
  IV U75228 ( .A(n54898), .Z(n54899) );
  NOR U75229 ( .A(n54899), .B(n54902), .Z(n60222) );
  NOR U75230 ( .A(n60220), .B(n60222), .Z(n58877) );
  IV U75231 ( .A(n54900), .Z(n54901) );
  NOR U75232 ( .A(n54902), .B(n54901), .Z(n60225) );
  IV U75233 ( .A(n54903), .Z(n54904) );
  NOR U75234 ( .A(n54905), .B(n54904), .Z(n60229) );
  IV U75235 ( .A(n54906), .Z(n54908) );
  IV U75236 ( .A(n54907), .Z(n54913) );
  NOR U75237 ( .A(n54908), .B(n54913), .Z(n60231) );
  NOR U75238 ( .A(n60229), .B(n60231), .Z(n58876) );
  IV U75239 ( .A(n54909), .Z(n54911) );
  NOR U75240 ( .A(n54911), .B(n54910), .Z(n64112) );
  IV U75241 ( .A(n54912), .Z(n54914) );
  NOR U75242 ( .A(n54914), .B(n54913), .Z(n60234) );
  NOR U75243 ( .A(n64112), .B(n60234), .Z(n58875) );
  NOR U75244 ( .A(n54916), .B(n54915), .Z(n54917) );
  IV U75245 ( .A(n54917), .Z(n64086) );
  NOR U75246 ( .A(n64086), .B(n54918), .Z(n58874) );
  IV U75247 ( .A(n54919), .Z(n54922) );
  IV U75248 ( .A(n54920), .Z(n54921) );
  NOR U75249 ( .A(n54922), .B(n54921), .Z(n64074) );
  IV U75250 ( .A(n54923), .Z(n54927) );
  NOR U75251 ( .A(n54925), .B(n54924), .Z(n54926) );
  IV U75252 ( .A(n54926), .Z(n54929) );
  NOR U75253 ( .A(n54927), .B(n54929), .Z(n64067) );
  IV U75254 ( .A(n54928), .Z(n54930) );
  NOR U75255 ( .A(n54930), .B(n54929), .Z(n64063) );
  NOR U75256 ( .A(n54932), .B(n54931), .Z(n60242) );
  IV U75257 ( .A(n54933), .Z(n54937) );
  IV U75258 ( .A(n54934), .Z(n58850) );
  NOR U75259 ( .A(n54935), .B(n58850), .Z(n54936) );
  IV U75260 ( .A(n54936), .Z(n58855) );
  NOR U75261 ( .A(n54937), .B(n58855), .Z(n60248) );
  NOR U75262 ( .A(n60242), .B(n60248), .Z(n58862) );
  IV U75263 ( .A(n54938), .Z(n54943) );
  NOR U75264 ( .A(n58844), .B(n54939), .Z(n54940) );
  IV U75265 ( .A(n54940), .Z(n60253) );
  NOR U75266 ( .A(n54941), .B(n60253), .Z(n54942) );
  IV U75267 ( .A(n54942), .Z(n54945) );
  NOR U75268 ( .A(n54943), .B(n54945), .Z(n60262) );
  IV U75269 ( .A(n54944), .Z(n54946) );
  NOR U75270 ( .A(n54946), .B(n54945), .Z(n54947) );
  IV U75271 ( .A(n54947), .Z(n64056) );
  IV U75272 ( .A(n54948), .Z(n54949) );
  NOR U75273 ( .A(n58846), .B(n54949), .Z(n54950) );
  IV U75274 ( .A(n54950), .Z(n60266) );
  IV U75275 ( .A(n54951), .Z(n54953) );
  NOR U75276 ( .A(n54953), .B(n54952), .Z(n60268) );
  NOR U75277 ( .A(n60270), .B(n60268), .Z(n58841) );
  IV U75278 ( .A(n54954), .Z(n54955) );
  NOR U75279 ( .A(n54958), .B(n54955), .Z(n60276) );
  IV U75280 ( .A(n54956), .Z(n54957) );
  NOR U75281 ( .A(n54958), .B(n54957), .Z(n60273) );
  IV U75282 ( .A(n54959), .Z(n54960) );
  NOR U75283 ( .A(n54960), .B(n58839), .Z(n64048) );
  IV U75284 ( .A(n54961), .Z(n54962) );
  NOR U75285 ( .A(n54963), .B(n54962), .Z(n58822) );
  IV U75286 ( .A(n58822), .Z(n58816) );
  IV U75287 ( .A(n54964), .Z(n54965) );
  NOR U75288 ( .A(n54965), .B(n58810), .Z(n54966) );
  IV U75289 ( .A(n54966), .Z(n60292) );
  IV U75290 ( .A(n54967), .Z(n54969) );
  NOR U75291 ( .A(n54969), .B(n54968), .Z(n54970) );
  IV U75292 ( .A(n54970), .Z(n58811) );
  IV U75293 ( .A(n65623), .Z(n54971) );
  NOR U75294 ( .A(n65622), .B(n54971), .Z(n54972) );
  IV U75295 ( .A(n54972), .Z(n64032) );
  IV U75296 ( .A(n54973), .Z(n54975) );
  NOR U75297 ( .A(n54975), .B(n54974), .Z(n54976) );
  IV U75298 ( .A(n54976), .Z(n58802) );
  IV U75299 ( .A(n54977), .Z(n58792) );
  IV U75300 ( .A(n54978), .Z(n54979) );
  NOR U75301 ( .A(n58792), .B(n54979), .Z(n64021) );
  IV U75302 ( .A(n54980), .Z(n54981) );
  NOR U75303 ( .A(n54982), .B(n54981), .Z(n60319) );
  NOR U75304 ( .A(n60317), .B(n60319), .Z(n58749) );
  XOR U75305 ( .A(n54984), .B(n54983), .Z(n54985) );
  NOR U75306 ( .A(n54986), .B(n54985), .Z(n54987) );
  IV U75307 ( .A(n54987), .Z(n54989) );
  NOR U75308 ( .A(n54988), .B(n54989), .Z(n60322) );
  NOR U75309 ( .A(n54990), .B(n54989), .Z(n63985) );
  IV U75310 ( .A(n54991), .Z(n54992) );
  NOR U75311 ( .A(n54992), .B(n54994), .Z(n60328) );
  IV U75312 ( .A(n54993), .Z(n54995) );
  NOR U75313 ( .A(n54995), .B(n54994), .Z(n63988) );
  IV U75314 ( .A(n54996), .Z(n54997) );
  NOR U75315 ( .A(n54998), .B(n54997), .Z(n63982) );
  IV U75316 ( .A(n54999), .Z(n55001) );
  IV U75317 ( .A(n55000), .Z(n58744) );
  NOR U75318 ( .A(n55001), .B(n58744), .Z(n63975) );
  NOR U75319 ( .A(n63982), .B(n63975), .Z(n58748) );
  IV U75320 ( .A(n55002), .Z(n55003) );
  NOR U75321 ( .A(n55004), .B(n55003), .Z(n63943) );
  IV U75322 ( .A(n55005), .Z(n55007) );
  IV U75323 ( .A(n55006), .Z(n58727) );
  NOR U75324 ( .A(n55007), .B(n58727), .Z(n63946) );
  NOR U75325 ( .A(n63943), .B(n63946), .Z(n60351) );
  IV U75326 ( .A(n55008), .Z(n55009) );
  NOR U75327 ( .A(n55009), .B(n55014), .Z(n63948) );
  IV U75328 ( .A(n55010), .Z(n55012) );
  XOR U75329 ( .A(n55013), .B(n55014), .Z(n55011) );
  NOR U75330 ( .A(n55012), .B(n55011), .Z(n63930) );
  NOR U75331 ( .A(n63948), .B(n63930), .Z(n58725) );
  IV U75332 ( .A(n55013), .Z(n55015) );
  NOR U75333 ( .A(n55015), .B(n55014), .Z(n60352) );
  IV U75334 ( .A(n55016), .Z(n58719) );
  IV U75335 ( .A(n55017), .Z(n55018) );
  NOR U75336 ( .A(n58719), .B(n55018), .Z(n60357) );
  NOR U75337 ( .A(n60352), .B(n60357), .Z(n58724) );
  IV U75338 ( .A(n55019), .Z(n55020) );
  NOR U75339 ( .A(n55020), .B(n58716), .Z(n60366) );
  IV U75340 ( .A(n55021), .Z(n55023) );
  NOR U75341 ( .A(n55023), .B(n55022), .Z(n55024) );
  IV U75342 ( .A(n55024), .Z(n58709) );
  IV U75343 ( .A(n55025), .Z(n55027) );
  NOR U75344 ( .A(n55027), .B(n55026), .Z(n58694) );
  IV U75345 ( .A(n58694), .Z(n58690) );
  IV U75346 ( .A(n55028), .Z(n55030) );
  IV U75347 ( .A(n55029), .Z(n55032) );
  NOR U75348 ( .A(n55030), .B(n55032), .Z(n60378) );
  IV U75349 ( .A(n55031), .Z(n55033) );
  NOR U75350 ( .A(n55033), .B(n55032), .Z(n63915) );
  IV U75351 ( .A(n55034), .Z(n55035) );
  NOR U75352 ( .A(n55035), .B(n58687), .Z(n55036) );
  IV U75353 ( .A(n55036), .Z(n63914) );
  IV U75354 ( .A(n55037), .Z(n55044) );
  NOR U75355 ( .A(n55039), .B(n55038), .Z(n55040) );
  IV U75356 ( .A(n55040), .Z(n55041) );
  NOR U75357 ( .A(n55042), .B(n55041), .Z(n55043) );
  IV U75358 ( .A(n55043), .Z(n58680) );
  NOR U75359 ( .A(n55044), .B(n58680), .Z(n63899) );
  IV U75360 ( .A(n55045), .Z(n55046) );
  NOR U75361 ( .A(n55047), .B(n55046), .Z(n60386) );
  IV U75362 ( .A(n55048), .Z(n55049) );
  NOR U75363 ( .A(n55049), .B(n58673), .Z(n63895) );
  NOR U75364 ( .A(n60386), .B(n63895), .Z(n58678) );
  IV U75365 ( .A(n55050), .Z(n55052) );
  NOR U75366 ( .A(n55052), .B(n55051), .Z(n63880) );
  IV U75367 ( .A(n55053), .Z(n58655) );
  NOR U75368 ( .A(n58655), .B(n55054), .Z(n63877) );
  IV U75369 ( .A(n55055), .Z(n55056) );
  NOR U75370 ( .A(n55057), .B(n55056), .Z(n60406) );
  IV U75371 ( .A(n55058), .Z(n55060) );
  NOR U75372 ( .A(n55060), .B(n55059), .Z(n60404) );
  NOR U75373 ( .A(n60406), .B(n60404), .Z(n58639) );
  IV U75374 ( .A(n55061), .Z(n55063) );
  NOR U75375 ( .A(n55063), .B(n55062), .Z(n60413) );
  IV U75376 ( .A(n55064), .Z(n60411) );
  IV U75377 ( .A(n55065), .Z(n58629) );
  IV U75378 ( .A(n55066), .Z(n55067) );
  NOR U75379 ( .A(n58629), .B(n55067), .Z(n74234) );
  NOR U75380 ( .A(n74225), .B(n74234), .Z(n60416) );
  IV U75381 ( .A(n55068), .Z(n55071) );
  XOR U75382 ( .A(n58617), .B(n58618), .Z(n69145) );
  NOR U75383 ( .A(n55069), .B(n69145), .Z(n55070) );
  IV U75384 ( .A(n55070), .Z(n55074) );
  NOR U75385 ( .A(n55071), .B(n55074), .Z(n60417) );
  IV U75386 ( .A(n55072), .Z(n69148) );
  NOR U75387 ( .A(n69148), .B(n58618), .Z(n55076) );
  IV U75388 ( .A(n55073), .Z(n55075) );
  NOR U75389 ( .A(n55075), .B(n55074), .Z(n65776) );
  NOR U75390 ( .A(n55076), .B(n65776), .Z(n63860) );
  IV U75391 ( .A(n55077), .Z(n55079) );
  NOR U75392 ( .A(n55079), .B(n55078), .Z(n55080) );
  IV U75393 ( .A(n55080), .Z(n58623) );
  IV U75394 ( .A(n55081), .Z(n55088) );
  NOR U75395 ( .A(n55083), .B(n55082), .Z(n55084) );
  IV U75396 ( .A(n55084), .Z(n55085) );
  NOR U75397 ( .A(n55086), .B(n55085), .Z(n55087) );
  IV U75398 ( .A(n55087), .Z(n58615) );
  NOR U75399 ( .A(n55088), .B(n58615), .Z(n63849) );
  IV U75400 ( .A(n55089), .Z(n55090) );
  NOR U75401 ( .A(n55091), .B(n55090), .Z(n55092) );
  IV U75402 ( .A(n55092), .Z(n58608) );
  IV U75403 ( .A(n55093), .Z(n55095) );
  IV U75404 ( .A(n55094), .Z(n55097) );
  NOR U75405 ( .A(n55095), .B(n55097), .Z(n60432) );
  IV U75406 ( .A(n55096), .Z(n55098) );
  NOR U75407 ( .A(n55098), .B(n55097), .Z(n60429) );
  IV U75408 ( .A(n55099), .Z(n55100) );
  NOR U75409 ( .A(n55100), .B(n55106), .Z(n60435) );
  IV U75410 ( .A(n55101), .Z(n55103) );
  NOR U75411 ( .A(n55103), .B(n55102), .Z(n63838) );
  IV U75412 ( .A(n55104), .Z(n55105) );
  NOR U75413 ( .A(n55106), .B(n55105), .Z(n63841) );
  NOR U75414 ( .A(n63838), .B(n63841), .Z(n55107) );
  IV U75415 ( .A(n55107), .Z(n58601) );
  IV U75416 ( .A(n55108), .Z(n55109) );
  NOR U75417 ( .A(n55110), .B(n55109), .Z(n63835) );
  IV U75418 ( .A(n55111), .Z(n55112) );
  NOR U75419 ( .A(n58593), .B(n55112), .Z(n60440) );
  NOR U75420 ( .A(n63835), .B(n60440), .Z(n58600) );
  IV U75421 ( .A(n55113), .Z(n55114) );
  NOR U75422 ( .A(n55115), .B(n55114), .Z(n55116) );
  IV U75423 ( .A(n55116), .Z(n58595) );
  IV U75424 ( .A(n55117), .Z(n55118) );
  NOR U75425 ( .A(n55119), .B(n55118), .Z(n60455) );
  IV U75426 ( .A(n55120), .Z(n58559) );
  NOR U75427 ( .A(n58559), .B(n55121), .Z(n60464) );
  IV U75428 ( .A(n55122), .Z(n55124) );
  NOR U75429 ( .A(n55124), .B(n55123), .Z(n63821) );
  IV U75430 ( .A(n55125), .Z(n55126) );
  NOR U75431 ( .A(n55127), .B(n55126), .Z(n55128) );
  IV U75432 ( .A(n55128), .Z(n55129) );
  NOR U75433 ( .A(n55129), .B(n58544), .Z(n63810) );
  IV U75434 ( .A(n55130), .Z(n55132) );
  NOR U75435 ( .A(n55132), .B(n55131), .Z(n60473) );
  IV U75436 ( .A(n58537), .Z(n55133) );
  NOR U75437 ( .A(n55133), .B(n58544), .Z(n63807) );
  NOR U75438 ( .A(n60473), .B(n63807), .Z(n58535) );
  IV U75439 ( .A(n55134), .Z(n55135) );
  NOR U75440 ( .A(n55140), .B(n55135), .Z(n69084) );
  IV U75441 ( .A(n55136), .Z(n55138) );
  NOR U75442 ( .A(n55138), .B(n55137), .Z(n74118) );
  IV U75443 ( .A(n55139), .Z(n55141) );
  NOR U75444 ( .A(n55141), .B(n55140), .Z(n70792) );
  NOR U75445 ( .A(n74118), .B(n70792), .Z(n65828) );
  IV U75446 ( .A(n65828), .Z(n55142) );
  NOR U75447 ( .A(n69084), .B(n55142), .Z(n60476) );
  IV U75448 ( .A(n55143), .Z(n55144) );
  NOR U75449 ( .A(n55145), .B(n55144), .Z(n60477) );
  IV U75450 ( .A(n55146), .Z(n55149) );
  IV U75451 ( .A(n55147), .Z(n55148) );
  NOR U75452 ( .A(n55149), .B(n55148), .Z(n63795) );
  NOR U75453 ( .A(n60477), .B(n63795), .Z(n58534) );
  NOR U75454 ( .A(n55151), .B(n55150), .Z(n69074) );
  IV U75455 ( .A(n55152), .Z(n55153) );
  NOR U75456 ( .A(n55153), .B(n55155), .Z(n65832) );
  NOR U75457 ( .A(n69074), .B(n65832), .Z(n63800) );
  IV U75458 ( .A(n55154), .Z(n55161) );
  NOR U75459 ( .A(n55156), .B(n55155), .Z(n55157) );
  IV U75460 ( .A(n55157), .Z(n55158) );
  NOR U75461 ( .A(n55159), .B(n55158), .Z(n55160) );
  IV U75462 ( .A(n55160), .Z(n55163) );
  NOR U75463 ( .A(n55161), .B(n55163), .Z(n60481) );
  IV U75464 ( .A(n55162), .Z(n55164) );
  NOR U75465 ( .A(n55164), .B(n55163), .Z(n60486) );
  IV U75466 ( .A(n55165), .Z(n55166) );
  NOR U75467 ( .A(n55166), .B(n55171), .Z(n65836) );
  IV U75468 ( .A(n55167), .Z(n55169) );
  NOR U75469 ( .A(n55169), .B(n55168), .Z(n65844) );
  IV U75470 ( .A(n55170), .Z(n55172) );
  NOR U75471 ( .A(n55172), .B(n55171), .Z(n70815) );
  NOR U75472 ( .A(n65844), .B(n70815), .Z(n60489) );
  IV U75473 ( .A(n55173), .Z(n55174) );
  NOR U75474 ( .A(n58530), .B(n55174), .Z(n55175) );
  IV U75475 ( .A(n55175), .Z(n55180) );
  NOR U75476 ( .A(n55177), .B(n55176), .Z(n55178) );
  IV U75477 ( .A(n55178), .Z(n55179) );
  NOR U75478 ( .A(n55180), .B(n55179), .Z(n60490) );
  IV U75479 ( .A(n55181), .Z(n55183) );
  NOR U75480 ( .A(n55183), .B(n55182), .Z(n60500) );
  IV U75481 ( .A(n55184), .Z(n55190) );
  NOR U75482 ( .A(n55185), .B(n55190), .Z(n55186) );
  IV U75483 ( .A(n55186), .Z(n55187) );
  NOR U75484 ( .A(n55188), .B(n55187), .Z(n60502) );
  NOR U75485 ( .A(n60500), .B(n60502), .Z(n58525) );
  IV U75486 ( .A(n55189), .Z(n55191) );
  NOR U75487 ( .A(n55191), .B(n55190), .Z(n60505) );
  NOR U75488 ( .A(n60507), .B(n60505), .Z(n55192) );
  IV U75489 ( .A(n55192), .Z(n58524) );
  NOR U75490 ( .A(n60515), .B(n60510), .Z(n58523) );
  IV U75491 ( .A(n55193), .Z(n55195) );
  NOR U75492 ( .A(n55195), .B(n55194), .Z(n65861) );
  IV U75493 ( .A(n55196), .Z(n55198) );
  NOR U75494 ( .A(n55198), .B(n55197), .Z(n60513) );
  NOR U75495 ( .A(n65861), .B(n60513), .Z(n58522) );
  IV U75496 ( .A(n55199), .Z(n79545) );
  NOR U75497 ( .A(n79545), .B(n65875), .Z(n58510) );
  IV U75498 ( .A(n58510), .Z(n58504) );
  IV U75499 ( .A(n55200), .Z(n55202) );
  NOR U75500 ( .A(n55202), .B(n55201), .Z(n60525) );
  IV U75501 ( .A(n55203), .Z(n55210) );
  NOR U75502 ( .A(n55205), .B(n55204), .Z(n55206) );
  IV U75503 ( .A(n55206), .Z(n55207) );
  NOR U75504 ( .A(n55208), .B(n55207), .Z(n55209) );
  IV U75505 ( .A(n55209), .Z(n58500) );
  NOR U75506 ( .A(n55210), .B(n58500), .Z(n60534) );
  IV U75507 ( .A(n55211), .Z(n58495) );
  IV U75508 ( .A(n55212), .Z(n55213) );
  NOR U75509 ( .A(n58495), .B(n55213), .Z(n60531) );
  IV U75510 ( .A(n55214), .Z(n55215) );
  NOR U75511 ( .A(n55215), .B(n58485), .Z(n60537) );
  NOR U75512 ( .A(n55217), .B(n55216), .Z(n55218) );
  IV U75513 ( .A(n55218), .Z(n55219) );
  XOR U75514 ( .A(n58474), .B(n58478), .Z(n55224) );
  NOR U75515 ( .A(n55219), .B(n55224), .Z(n60545) );
  NOR U75516 ( .A(n60537), .B(n60545), .Z(n58483) );
  IV U75517 ( .A(n55220), .Z(n55222) );
  NOR U75518 ( .A(n55222), .B(n55221), .Z(n55223) );
  IV U75519 ( .A(n55223), .Z(n55225) );
  NOR U75520 ( .A(n55225), .B(n55224), .Z(n60542) );
  IV U75521 ( .A(n55226), .Z(n55228) );
  IV U75522 ( .A(n55227), .Z(n58457) );
  NOR U75523 ( .A(n55228), .B(n58457), .Z(n63766) );
  IV U75524 ( .A(n55229), .Z(n55230) );
  NOR U75525 ( .A(n55230), .B(n58454), .Z(n63755) );
  IV U75526 ( .A(n55231), .Z(n55233) );
  NOR U75527 ( .A(n55233), .B(n55232), .Z(n58450) );
  IV U75528 ( .A(n58450), .Z(n58440) );
  IV U75529 ( .A(n55234), .Z(n55235) );
  NOR U75530 ( .A(n55236), .B(n55235), .Z(n63748) );
  IV U75531 ( .A(n55237), .Z(n55238) );
  NOR U75532 ( .A(n55238), .B(n55245), .Z(n63746) );
  NOR U75533 ( .A(n63748), .B(n63746), .Z(n58438) );
  IV U75534 ( .A(n55239), .Z(n55243) );
  NOR U75535 ( .A(n55241), .B(n55240), .Z(n55242) );
  IV U75536 ( .A(n55242), .Z(n55249) );
  NOR U75537 ( .A(n55243), .B(n55249), .Z(n63737) );
  IV U75538 ( .A(n55244), .Z(n55246) );
  NOR U75539 ( .A(n55246), .B(n55245), .Z(n63741) );
  NOR U75540 ( .A(n63737), .B(n63741), .Z(n55247) );
  IV U75541 ( .A(n55247), .Z(n58437) );
  IV U75542 ( .A(n55248), .Z(n55250) );
  NOR U75543 ( .A(n55250), .B(n55249), .Z(n63739) );
  IV U75544 ( .A(n55251), .Z(n55254) );
  NOR U75545 ( .A(n55252), .B(n55256), .Z(n55253) );
  IV U75546 ( .A(n55253), .Z(n58422) );
  NOR U75547 ( .A(n55254), .B(n58422), .Z(n65940) );
  IV U75548 ( .A(n55255), .Z(n55257) );
  NOR U75549 ( .A(n55257), .B(n55256), .Z(n69019) );
  NOR U75550 ( .A(n65940), .B(n69019), .Z(n63731) );
  IV U75551 ( .A(n55258), .Z(n55259) );
  NOR U75552 ( .A(n55259), .B(n58395), .Z(n63710) );
  IV U75553 ( .A(n55260), .Z(n55261) );
  NOR U75554 ( .A(n55261), .B(n58395), .Z(n55262) );
  IV U75555 ( .A(n55262), .Z(n55263) );
  NOR U75556 ( .A(n58391), .B(n55263), .Z(n79421) );
  NOR U75557 ( .A(n63710), .B(n79421), .Z(n58405) );
  IV U75558 ( .A(n55264), .Z(n55267) );
  NOR U75559 ( .A(n55265), .B(n55272), .Z(n55266) );
  IV U75560 ( .A(n55266), .Z(n55269) );
  NOR U75561 ( .A(n55267), .B(n55269), .Z(n63701) );
  IV U75562 ( .A(n55268), .Z(n55270) );
  NOR U75563 ( .A(n55270), .B(n55269), .Z(n60575) );
  IV U75564 ( .A(n55271), .Z(n55273) );
  NOR U75565 ( .A(n55273), .B(n55272), .Z(n60579) );
  NOR U75566 ( .A(n65985), .B(n60579), .Z(n58377) );
  IV U75567 ( .A(n55274), .Z(n55276) );
  NOR U75568 ( .A(n55276), .B(n55275), .Z(n63694) );
  NOR U75569 ( .A(n63694), .B(n65990), .Z(n58376) );
  IV U75570 ( .A(n55277), .Z(n55278) );
  NOR U75571 ( .A(n58370), .B(n55278), .Z(n63692) );
  IV U75572 ( .A(n55279), .Z(n55281) );
  IV U75573 ( .A(n55280), .Z(n58372) );
  NOR U75574 ( .A(n55281), .B(n58372), .Z(n60584) );
  IV U75575 ( .A(n55282), .Z(n55283) );
  NOR U75576 ( .A(n58365), .B(n55283), .Z(n60593) );
  IV U75577 ( .A(n55284), .Z(n55285) );
  NOR U75578 ( .A(n55286), .B(n55285), .Z(n60590) );
  IV U75579 ( .A(n55287), .Z(n55290) );
  IV U75580 ( .A(n55288), .Z(n55289) );
  NOR U75581 ( .A(n55290), .B(n55289), .Z(n60596) );
  NOR U75582 ( .A(n63679), .B(n60596), .Z(n55291) );
  IV U75583 ( .A(n55291), .Z(n58362) );
  IV U75584 ( .A(n55292), .Z(n55293) );
  NOR U75585 ( .A(n55294), .B(n55293), .Z(n55295) );
  IV U75586 ( .A(n55295), .Z(n58353) );
  IV U75587 ( .A(n55296), .Z(n55300) );
  NOR U75588 ( .A(n55298), .B(n55297), .Z(n55299) );
  IV U75589 ( .A(n55299), .Z(n55305) );
  NOR U75590 ( .A(n55300), .B(n55305), .Z(n60602) );
  IV U75591 ( .A(n55301), .Z(n55303) );
  NOR U75592 ( .A(n55303), .B(n55302), .Z(n60609) );
  IV U75593 ( .A(n55304), .Z(n55306) );
  NOR U75594 ( .A(n55306), .B(n55305), .Z(n63672) );
  NOR U75595 ( .A(n60609), .B(n63672), .Z(n58346) );
  IV U75596 ( .A(n55307), .Z(n55308) );
  NOR U75597 ( .A(n55309), .B(n55308), .Z(n60611) );
  IV U75598 ( .A(n55310), .Z(n55317) );
  IV U75599 ( .A(n55311), .Z(n58342) );
  NOR U75600 ( .A(n55312), .B(n58342), .Z(n55313) );
  IV U75601 ( .A(n55313), .Z(n55314) );
  NOR U75602 ( .A(n55315), .B(n55314), .Z(n55316) );
  IV U75603 ( .A(n55316), .Z(n55319) );
  NOR U75604 ( .A(n55317), .B(n55319), .Z(n63655) );
  NOR U75605 ( .A(n60611), .B(n63655), .Z(n58345) );
  IV U75606 ( .A(n55318), .Z(n55320) );
  NOR U75607 ( .A(n55320), .B(n55319), .Z(n60614) );
  IV U75608 ( .A(n55321), .Z(n55323) );
  IV U75609 ( .A(n55322), .Z(n58334) );
  NOR U75610 ( .A(n55323), .B(n58334), .Z(n68953) );
  NOR U75611 ( .A(n68946), .B(n68953), .Z(n60624) );
  NOR U75612 ( .A(n55325), .B(n55324), .Z(n60625) );
  IV U75613 ( .A(n55326), .Z(n58329) );
  IV U75614 ( .A(n55327), .Z(n55328) );
  NOR U75615 ( .A(n58329), .B(n55328), .Z(n63629) );
  NOR U75616 ( .A(n60625), .B(n63629), .Z(n55329) );
  IV U75617 ( .A(n55329), .Z(n58326) );
  IV U75618 ( .A(n55330), .Z(n55331) );
  NOR U75619 ( .A(n55332), .B(n55331), .Z(n60631) );
  IV U75620 ( .A(n55333), .Z(n55336) );
  IV U75621 ( .A(n55334), .Z(n55335) );
  NOR U75622 ( .A(n55336), .B(n55335), .Z(n60628) );
  IV U75623 ( .A(n55337), .Z(n55341) );
  NOR U75624 ( .A(n55339), .B(n55338), .Z(n55340) );
  IV U75625 ( .A(n55340), .Z(n58318) );
  NOR U75626 ( .A(n55341), .B(n58318), .Z(n60638) );
  IV U75627 ( .A(n55342), .Z(n55344) );
  NOR U75628 ( .A(n55344), .B(n55343), .Z(n66050) );
  IV U75629 ( .A(n55345), .Z(n55347) );
  NOR U75630 ( .A(n55347), .B(n55346), .Z(n66046) );
  NOR U75631 ( .A(n66050), .B(n66046), .Z(n60637) );
  IV U75632 ( .A(n55348), .Z(n55349) );
  NOR U75633 ( .A(n55350), .B(n55349), .Z(n66058) );
  IV U75634 ( .A(n55351), .Z(n55352) );
  NOR U75635 ( .A(n55353), .B(n55352), .Z(n66053) );
  NOR U75636 ( .A(n66058), .B(n66053), .Z(n60641) );
  IV U75637 ( .A(n55354), .Z(n55355) );
  NOR U75638 ( .A(n55356), .B(n55355), .Z(n66069) );
  NOR U75639 ( .A(n66073), .B(n66069), .Z(n63595) );
  IV U75640 ( .A(n55357), .Z(n55358) );
  NOR U75641 ( .A(n55361), .B(n55358), .Z(n66081) );
  IV U75642 ( .A(n55359), .Z(n55360) );
  NOR U75643 ( .A(n55361), .B(n55360), .Z(n66076) );
  NOR U75644 ( .A(n66081), .B(n66076), .Z(n63593) );
  IV U75645 ( .A(n55362), .Z(n55363) );
  NOR U75646 ( .A(n55363), .B(n55369), .Z(n60644) );
  IV U75647 ( .A(n55364), .Z(n55365) );
  NOR U75648 ( .A(n55366), .B(n55365), .Z(n60647) );
  IV U75649 ( .A(n55367), .Z(n55368) );
  NOR U75650 ( .A(n55369), .B(n55368), .Z(n60642) );
  NOR U75651 ( .A(n60647), .B(n60642), .Z(n55370) );
  IV U75652 ( .A(n55370), .Z(n58311) );
  IV U75653 ( .A(n55371), .Z(n55373) );
  IV U75654 ( .A(n55372), .Z(n55375) );
  NOR U75655 ( .A(n55373), .B(n55375), .Z(n63579) );
  IV U75656 ( .A(n55374), .Z(n55376) );
  NOR U75657 ( .A(n55376), .B(n55375), .Z(n60651) );
  IV U75658 ( .A(n55377), .Z(n55379) );
  NOR U75659 ( .A(n55379), .B(n55378), .Z(n63582) );
  IV U75660 ( .A(n55380), .Z(n58290) );
  IV U75661 ( .A(n55381), .Z(n55382) );
  NOR U75662 ( .A(n58290), .B(n55382), .Z(n60663) );
  IV U75663 ( .A(n55383), .Z(n55384) );
  NOR U75664 ( .A(n55384), .B(n58286), .Z(n60669) );
  IV U75665 ( .A(n55385), .Z(n55386) );
  NOR U75666 ( .A(n55387), .B(n55386), .Z(n60674) );
  IV U75667 ( .A(n55388), .Z(n55392) );
  NOR U75668 ( .A(n55389), .B(n58283), .Z(n55390) );
  IV U75669 ( .A(n55390), .Z(n55391) );
  NOR U75670 ( .A(n55392), .B(n55391), .Z(n63557) );
  NOR U75671 ( .A(n60674), .B(n63557), .Z(n68917) );
  IV U75672 ( .A(n68917), .Z(n58281) );
  IV U75673 ( .A(n55393), .Z(n55394) );
  NOR U75674 ( .A(n55394), .B(n55399), .Z(n60672) );
  IV U75675 ( .A(n55395), .Z(n55403) );
  IV U75676 ( .A(n55396), .Z(n55397) );
  NOR U75677 ( .A(n55403), .B(n55397), .Z(n63548) );
  IV U75678 ( .A(n55398), .Z(n55400) );
  NOR U75679 ( .A(n55400), .B(n55399), .Z(n63543) );
  NOR U75680 ( .A(n63548), .B(n63543), .Z(n60679) );
  IV U75681 ( .A(n55401), .Z(n55402) );
  NOR U75682 ( .A(n55403), .B(n55402), .Z(n60680) );
  IV U75683 ( .A(n55404), .Z(n55406) );
  NOR U75684 ( .A(n55406), .B(n55405), .Z(n60683) );
  NOR U75685 ( .A(n60680), .B(n60683), .Z(n58280) );
  IV U75686 ( .A(n55407), .Z(n55408) );
  NOR U75687 ( .A(n55408), .B(n58273), .Z(n60694) );
  IV U75688 ( .A(n55409), .Z(n55411) );
  NOR U75689 ( .A(n55411), .B(n55410), .Z(n55412) );
  IV U75690 ( .A(n55412), .Z(n55419) );
  NOR U75691 ( .A(n55414), .B(n55413), .Z(n55415) );
  IV U75692 ( .A(n55415), .Z(n55416) );
  NOR U75693 ( .A(n55417), .B(n55416), .Z(n55418) );
  IV U75694 ( .A(n55418), .Z(n58262) );
  NOR U75695 ( .A(n55419), .B(n58262), .Z(n63531) );
  NOR U75696 ( .A(n60694), .B(n63531), .Z(n58269) );
  IV U75697 ( .A(n55420), .Z(n55421) );
  NOR U75698 ( .A(n55422), .B(n55421), .Z(n55423) );
  IV U75699 ( .A(n55423), .Z(n58264) );
  IV U75700 ( .A(n55424), .Z(n55425) );
  NOR U75701 ( .A(n55426), .B(n55425), .Z(n55427) );
  IV U75702 ( .A(n55427), .Z(n58248) );
  IV U75703 ( .A(n55428), .Z(n55435) );
  XOR U75704 ( .A(n58236), .B(n58237), .Z(n55429) );
  NOR U75705 ( .A(n55430), .B(n55429), .Z(n55431) );
  IV U75706 ( .A(n55431), .Z(n55432) );
  NOR U75707 ( .A(n55433), .B(n55432), .Z(n55434) );
  IV U75708 ( .A(n55434), .Z(n58240) );
  NOR U75709 ( .A(n55435), .B(n58240), .Z(n60708) );
  IV U75710 ( .A(n55436), .Z(n55438) );
  NOR U75711 ( .A(n55438), .B(n55437), .Z(n60722) );
  IV U75712 ( .A(n55439), .Z(n55441) );
  NOR U75713 ( .A(n55441), .B(n55440), .Z(n60714) );
  NOR U75714 ( .A(n60722), .B(n60714), .Z(n58235) );
  IV U75715 ( .A(n55442), .Z(n55446) );
  NOR U75716 ( .A(n55444), .B(n55443), .Z(n55445) );
  IV U75717 ( .A(n55445), .Z(n58232) );
  NOR U75718 ( .A(n55446), .B(n58232), .Z(n60719) );
  IV U75719 ( .A(n55447), .Z(n55449) );
  NOR U75720 ( .A(n55449), .B(n55448), .Z(n60725) );
  IV U75721 ( .A(n55450), .Z(n55451) );
  NOR U75722 ( .A(n55451), .B(n55453), .Z(n60743) );
  IV U75723 ( .A(n55452), .Z(n55454) );
  NOR U75724 ( .A(n55454), .B(n55453), .Z(n60740) );
  NOR U75725 ( .A(n60743), .B(n60740), .Z(n55455) );
  IV U75726 ( .A(n55455), .Z(n58222) );
  IV U75727 ( .A(n55456), .Z(n55459) );
  NOR U75728 ( .A(n55457), .B(n58212), .Z(n55458) );
  IV U75729 ( .A(n55458), .Z(n58220) );
  NOR U75730 ( .A(n55459), .B(n58220), .Z(n60739) );
  IV U75731 ( .A(n55460), .Z(n55461) );
  NOR U75732 ( .A(n55461), .B(n58183), .Z(n55462) );
  IV U75733 ( .A(n55462), .Z(n55463) );
  NOR U75734 ( .A(n58187), .B(n55463), .Z(n63485) );
  IV U75735 ( .A(n55464), .Z(n55465) );
  NOR U75736 ( .A(n55466), .B(n55465), .Z(n55467) );
  IV U75737 ( .A(n55467), .Z(n58171) );
  IV U75738 ( .A(n55468), .Z(n55469) );
  NOR U75739 ( .A(n55470), .B(n55469), .Z(n58158) );
  IV U75740 ( .A(n58158), .Z(n58152) );
  IV U75741 ( .A(n55471), .Z(n55473) );
  NOR U75742 ( .A(n55473), .B(n55472), .Z(n55474) );
  IV U75743 ( .A(n55474), .Z(n60773) );
  NOR U75744 ( .A(n55475), .B(n63444), .Z(n58145) );
  IV U75745 ( .A(n55476), .Z(n55477) );
  NOR U75746 ( .A(n55478), .B(n55477), .Z(n66199) );
  IV U75747 ( .A(n55479), .Z(n55481) );
  NOR U75748 ( .A(n55481), .B(n55480), .Z(n66193) );
  NOR U75749 ( .A(n66199), .B(n66193), .Z(n63440) );
  IV U75750 ( .A(n63440), .Z(n58144) );
  IV U75751 ( .A(n55482), .Z(n55484) );
  IV U75752 ( .A(n55483), .Z(n55488) );
  NOR U75753 ( .A(n55484), .B(n55488), .Z(n63437) );
  IV U75754 ( .A(n55485), .Z(n55486) );
  NOR U75755 ( .A(n55486), .B(n55491), .Z(n66211) );
  IV U75756 ( .A(n55487), .Z(n55489) );
  NOR U75757 ( .A(n55489), .B(n55488), .Z(n66202) );
  NOR U75758 ( .A(n66211), .B(n66202), .Z(n60777) );
  IV U75759 ( .A(n55490), .Z(n55492) );
  NOR U75760 ( .A(n55492), .B(n55491), .Z(n60778) );
  IV U75761 ( .A(n55493), .Z(n55501) );
  IV U75762 ( .A(n55494), .Z(n55495) );
  NOR U75763 ( .A(n55501), .B(n55495), .Z(n63430) );
  IV U75764 ( .A(n55496), .Z(n55498) );
  NOR U75765 ( .A(n55498), .B(n55497), .Z(n60781) );
  NOR U75766 ( .A(n63430), .B(n60781), .Z(n58142) );
  IV U75767 ( .A(n55499), .Z(n55500) );
  NOR U75768 ( .A(n55501), .B(n55500), .Z(n68796) );
  IV U75769 ( .A(n55502), .Z(n55503) );
  NOR U75770 ( .A(n55503), .B(n55508), .Z(n66216) );
  NOR U75771 ( .A(n68796), .B(n66216), .Z(n63429) );
  IV U75772 ( .A(n55504), .Z(n55505) );
  NOR U75773 ( .A(n55505), .B(n55508), .Z(n55506) );
  IV U75774 ( .A(n55506), .Z(n63427) );
  IV U75775 ( .A(n55507), .Z(n55509) );
  NOR U75776 ( .A(n55509), .B(n55508), .Z(n58138) );
  IV U75777 ( .A(n55510), .Z(n55512) );
  NOR U75778 ( .A(n55512), .B(n55511), .Z(n58135) );
  IV U75779 ( .A(n58135), .Z(n58127) );
  IV U75780 ( .A(n55513), .Z(n55514) );
  NOR U75781 ( .A(n55514), .B(n55520), .Z(n55515) );
  IV U75782 ( .A(n55515), .Z(n63397) );
  IV U75783 ( .A(n55516), .Z(n55518) );
  NOR U75784 ( .A(n55518), .B(n55517), .Z(n68766) );
  IV U75785 ( .A(n55519), .Z(n55521) );
  NOR U75786 ( .A(n55521), .B(n55520), .Z(n68775) );
  NOR U75787 ( .A(n68766), .B(n68775), .Z(n63394) );
  IV U75788 ( .A(n55522), .Z(n55523) );
  NOR U75789 ( .A(n55523), .B(n58109), .Z(n63389) );
  IV U75790 ( .A(n55524), .Z(n55525) );
  NOR U75791 ( .A(n55526), .B(n55525), .Z(n68751) );
  IV U75792 ( .A(n55527), .Z(n55528) );
  NOR U75793 ( .A(n55529), .B(n55528), .Z(n68756) );
  NOR U75794 ( .A(n68751), .B(n68756), .Z(n63384) );
  IV U75795 ( .A(n55530), .Z(n55535) );
  IV U75796 ( .A(n55531), .Z(n55532) );
  NOR U75797 ( .A(n55535), .B(n55532), .Z(n63381) );
  IV U75798 ( .A(n55533), .Z(n55534) );
  NOR U75799 ( .A(n55535), .B(n55534), .Z(n60787) );
  IV U75800 ( .A(n55536), .Z(n55537) );
  NOR U75801 ( .A(n58103), .B(n55537), .Z(n60784) );
  IV U75802 ( .A(n55538), .Z(n55539) );
  NOR U75803 ( .A(n55540), .B(n55539), .Z(n60791) );
  IV U75804 ( .A(n55541), .Z(n55542) );
  NOR U75805 ( .A(n55543), .B(n55542), .Z(n60794) );
  NOR U75806 ( .A(n60791), .B(n60794), .Z(n58097) );
  IV U75807 ( .A(n55544), .Z(n55545) );
  NOR U75808 ( .A(n55545), .B(n55551), .Z(n55546) );
  IV U75809 ( .A(n55546), .Z(n60799) );
  IV U75810 ( .A(n55547), .Z(n55549) );
  NOR U75811 ( .A(n55549), .B(n55548), .Z(n63374) );
  IV U75812 ( .A(n55550), .Z(n55552) );
  NOR U75813 ( .A(n55552), .B(n55551), .Z(n60803) );
  NOR U75814 ( .A(n63374), .B(n60803), .Z(n58090) );
  IV U75815 ( .A(n55553), .Z(n55554) );
  NOR U75816 ( .A(n55554), .B(n55559), .Z(n63373) );
  IV U75817 ( .A(n63373), .Z(n63371) );
  IV U75818 ( .A(n55555), .Z(n55556) );
  NOR U75819 ( .A(n55556), .B(n55559), .Z(n55557) );
  IV U75820 ( .A(n55557), .Z(n63360) );
  IV U75821 ( .A(n55558), .Z(n55560) );
  NOR U75822 ( .A(n55560), .B(n55559), .Z(n60807) );
  IV U75823 ( .A(n55561), .Z(n55566) );
  IV U75824 ( .A(n55562), .Z(n55563) );
  NOR U75825 ( .A(n55566), .B(n55563), .Z(n63349) );
  IV U75826 ( .A(n55564), .Z(n55565) );
  NOR U75827 ( .A(n55566), .B(n55565), .Z(n60813) );
  IV U75828 ( .A(n55567), .Z(n55568) );
  NOR U75829 ( .A(n55568), .B(n58079), .Z(n60816) );
  IV U75830 ( .A(n55569), .Z(n55571) );
  NOR U75831 ( .A(n55571), .B(n55570), .Z(n60823) );
  IV U75832 ( .A(n55572), .Z(n55574) );
  NOR U75833 ( .A(n55574), .B(n55573), .Z(n63332) );
  IV U75834 ( .A(n55575), .Z(n55576) );
  NOR U75835 ( .A(n55577), .B(n55576), .Z(n66264) );
  NOR U75836 ( .A(n63330), .B(n66264), .Z(n55578) );
  IV U75837 ( .A(n55578), .Z(n55579) );
  NOR U75838 ( .A(n63332), .B(n55579), .Z(n58074) );
  IV U75839 ( .A(n55580), .Z(n55584) );
  NOR U75840 ( .A(n55582), .B(n55581), .Z(n55583) );
  IV U75841 ( .A(n55583), .Z(n58071) );
  NOR U75842 ( .A(n55584), .B(n58071), .Z(n58066) );
  IV U75843 ( .A(n55585), .Z(n55586) );
  NOR U75844 ( .A(n55587), .B(n55586), .Z(n60830) );
  IV U75845 ( .A(n55588), .Z(n55589) );
  NOR U75846 ( .A(n55590), .B(n55589), .Z(n60832) );
  NOR U75847 ( .A(n60830), .B(n60832), .Z(n58065) );
  IV U75848 ( .A(n55591), .Z(n55595) );
  NOR U75849 ( .A(n55593), .B(n55592), .Z(n55594) );
  IV U75850 ( .A(n55594), .Z(n55597) );
  NOR U75851 ( .A(n55595), .B(n55597), .Z(n60840) );
  IV U75852 ( .A(n55596), .Z(n55598) );
  NOR U75853 ( .A(n55598), .B(n55597), .Z(n60837) );
  IV U75854 ( .A(n55599), .Z(n55603) );
  NOR U75855 ( .A(n55601), .B(n55600), .Z(n55602) );
  IV U75856 ( .A(n55602), .Z(n55605) );
  NOR U75857 ( .A(n55603), .B(n55605), .Z(n60846) );
  IV U75858 ( .A(n55604), .Z(n55606) );
  NOR U75859 ( .A(n55606), .B(n55605), .Z(n60843) );
  NOR U75860 ( .A(n55608), .B(n55607), .Z(n55609) );
  IV U75861 ( .A(n55609), .Z(n55614) );
  NOR U75862 ( .A(n55610), .B(n55614), .Z(n60849) );
  IV U75863 ( .A(n55611), .Z(n55618) );
  IV U75864 ( .A(n55612), .Z(n55613) );
  NOR U75865 ( .A(n55618), .B(n55613), .Z(n63320) );
  NOR U75866 ( .A(n55615), .B(n55614), .Z(n60853) );
  NOR U75867 ( .A(n63320), .B(n60853), .Z(n58064) );
  IV U75868 ( .A(n55619), .Z(n55616) );
  NOR U75869 ( .A(n55616), .B(n55618), .Z(n60858) );
  IV U75870 ( .A(n55617), .Z(n55621) );
  XOR U75871 ( .A(n55619), .B(n55618), .Z(n55620) );
  NOR U75872 ( .A(n55621), .B(n55620), .Z(n63317) );
  NOR U75873 ( .A(n60858), .B(n63317), .Z(n58063) );
  IV U75874 ( .A(n55622), .Z(n55623) );
  NOR U75875 ( .A(n55623), .B(n55626), .Z(n60855) );
  IV U75876 ( .A(n55624), .Z(n55625) );
  NOR U75877 ( .A(n55626), .B(n55625), .Z(n55627) );
  IV U75878 ( .A(n55627), .Z(n60863) );
  IV U75879 ( .A(n55628), .Z(n55629) );
  NOR U75880 ( .A(n58056), .B(n55629), .Z(n63308) );
  IV U75881 ( .A(n55630), .Z(n55635) );
  IV U75882 ( .A(n55631), .Z(n55632) );
  NOR U75883 ( .A(n55635), .B(n55632), .Z(n60869) );
  IV U75884 ( .A(n55633), .Z(n55634) );
  NOR U75885 ( .A(n55635), .B(n55634), .Z(n60873) );
  IV U75886 ( .A(n55636), .Z(n55637) );
  NOR U75887 ( .A(n58044), .B(n55637), .Z(n63284) );
  NOR U75888 ( .A(n60873), .B(n63284), .Z(n58046) );
  IV U75889 ( .A(n55638), .Z(n55642) );
  NOR U75890 ( .A(n55640), .B(n55639), .Z(n55641) );
  IV U75891 ( .A(n55641), .Z(n55644) );
  NOR U75892 ( .A(n55642), .B(n55644), .Z(n63277) );
  IV U75893 ( .A(n55643), .Z(n55645) );
  NOR U75894 ( .A(n55645), .B(n55644), .Z(n58034) );
  IV U75895 ( .A(n58026), .Z(n58019) );
  IV U75896 ( .A(n55646), .Z(n55648) );
  NOR U75897 ( .A(n55648), .B(n55647), .Z(n66327) );
  IV U75898 ( .A(n55649), .Z(n55650) );
  NOR U75899 ( .A(n55650), .B(n58021), .Z(n66321) );
  NOR U75900 ( .A(n66327), .B(n66321), .Z(n63258) );
  IV U75901 ( .A(n63258), .Z(n58023) );
  IV U75902 ( .A(n55651), .Z(n55656) );
  IV U75903 ( .A(n55652), .Z(n55653) );
  NOR U75904 ( .A(n55656), .B(n55653), .Z(n60878) );
  IV U75905 ( .A(n55654), .Z(n55655) );
  NOR U75906 ( .A(n55656), .B(n55655), .Z(n63251) );
  IV U75907 ( .A(n55657), .Z(n55658) );
  NOR U75908 ( .A(n55664), .B(n55658), .Z(n63248) );
  IV U75909 ( .A(n55659), .Z(n55661) );
  NOR U75910 ( .A(n55661), .B(n55660), .Z(n60887) );
  IV U75911 ( .A(n55662), .Z(n55663) );
  NOR U75912 ( .A(n55664), .B(n55663), .Z(n60882) );
  NOR U75913 ( .A(n60887), .B(n60882), .Z(n58017) );
  IV U75914 ( .A(n55665), .Z(n55672) );
  XOR U75915 ( .A(n55672), .B(n55671), .Z(n55666) );
  NOR U75916 ( .A(n55667), .B(n55666), .Z(n55668) );
  IV U75917 ( .A(n55668), .Z(n55669) );
  NOR U75918 ( .A(n55670), .B(n55669), .Z(n63240) );
  IV U75919 ( .A(n55671), .Z(n55673) );
  NOR U75920 ( .A(n55673), .B(n55672), .Z(n63237) );
  IV U75921 ( .A(n55674), .Z(n55676) );
  NOR U75922 ( .A(n55676), .B(n55675), .Z(n60902) );
  NOR U75923 ( .A(n63237), .B(n60902), .Z(n57996) );
  IV U75924 ( .A(n55677), .Z(n55679) );
  NOR U75925 ( .A(n55679), .B(n55678), .Z(n60907) );
  IV U75926 ( .A(n55680), .Z(n55684) );
  NOR U75927 ( .A(n55682), .B(n55681), .Z(n55683) );
  IV U75928 ( .A(n55683), .Z(n57987) );
  NOR U75929 ( .A(n55684), .B(n57987), .Z(n60914) );
  NOR U75930 ( .A(n60907), .B(n60914), .Z(n57989) );
  IV U75931 ( .A(n55685), .Z(n55686) );
  NOR U75932 ( .A(n55686), .B(n57979), .Z(n57974) );
  IV U75933 ( .A(n57974), .Z(n57968) );
  IV U75934 ( .A(n55687), .Z(n55689) );
  NOR U75935 ( .A(n55689), .B(n55688), .Z(n63223) );
  IV U75936 ( .A(n55690), .Z(n55692) );
  NOR U75937 ( .A(n55692), .B(n55691), .Z(n66378) );
  IV U75938 ( .A(n55693), .Z(n55695) );
  NOR U75939 ( .A(n55695), .B(n55694), .Z(n66374) );
  NOR U75940 ( .A(n66378), .B(n66374), .Z(n63222) );
  IV U75941 ( .A(n63222), .Z(n57966) );
  IV U75942 ( .A(n55696), .Z(n55698) );
  NOR U75943 ( .A(n55698), .B(n55697), .Z(n63215) );
  IV U75944 ( .A(n55699), .Z(n55700) );
  NOR U75945 ( .A(n55701), .B(n55700), .Z(n63219) );
  NOR U75946 ( .A(n63215), .B(n63219), .Z(n57965) );
  IV U75947 ( .A(n55702), .Z(n55704) );
  NOR U75948 ( .A(n55704), .B(n55703), .Z(n63206) );
  IV U75949 ( .A(n55705), .Z(n55706) );
  NOR U75950 ( .A(n55706), .B(n55709), .Z(n60924) );
  IV U75951 ( .A(n55707), .Z(n55708) );
  NOR U75952 ( .A(n55709), .B(n55708), .Z(n60922) );
  IV U75953 ( .A(n55710), .Z(n55712) );
  IV U75954 ( .A(n55711), .Z(n55714) );
  NOR U75955 ( .A(n55712), .B(n55714), .Z(n60930) );
  IV U75956 ( .A(n55713), .Z(n55715) );
  NOR U75957 ( .A(n55715), .B(n55714), .Z(n60928) );
  XOR U75958 ( .A(n60930), .B(n60928), .Z(n55716) );
  NOR U75959 ( .A(n60922), .B(n55716), .Z(n57956) );
  IV U75960 ( .A(n55717), .Z(n55718) );
  NOR U75961 ( .A(n55718), .B(n55721), .Z(n60936) );
  IV U75962 ( .A(n55719), .Z(n55720) );
  NOR U75963 ( .A(n55721), .B(n55720), .Z(n60933) );
  IV U75964 ( .A(n55722), .Z(n55723) );
  NOR U75965 ( .A(n57941), .B(n55723), .Z(n63191) );
  NOR U75966 ( .A(n57938), .B(n55724), .Z(n55725) );
  IV U75967 ( .A(n55725), .Z(n57931) );
  NOR U75968 ( .A(n55726), .B(n57931), .Z(n60945) );
  IV U75969 ( .A(n55727), .Z(n55728) );
  NOR U75970 ( .A(n55728), .B(n57926), .Z(n60957) );
  IV U75971 ( .A(n55729), .Z(n55730) );
  NOR U75972 ( .A(n55731), .B(n55730), .Z(n63182) );
  IV U75973 ( .A(n55732), .Z(n55740) );
  IV U75974 ( .A(n55733), .Z(n55734) );
  NOR U75975 ( .A(n55740), .B(n55734), .Z(n63180) );
  XOR U75976 ( .A(n63182), .B(n63180), .Z(n55735) );
  NOR U75977 ( .A(n60957), .B(n55735), .Z(n57924) );
  IV U75978 ( .A(n55736), .Z(n55737) );
  NOR U75979 ( .A(n55737), .B(n55742), .Z(n71358) );
  IV U75980 ( .A(n55738), .Z(n55739) );
  NOR U75981 ( .A(n55740), .B(n55739), .Z(n71348) );
  NOR U75982 ( .A(n71358), .B(n71348), .Z(n60962) );
  IV U75983 ( .A(n55741), .Z(n55743) );
  NOR U75984 ( .A(n55743), .B(n55742), .Z(n60963) );
  IV U75985 ( .A(n55744), .Z(n55747) );
  IV U75986 ( .A(n55745), .Z(n55750) );
  XOR U75987 ( .A(n55748), .B(n55750), .Z(n55746) );
  NOR U75988 ( .A(n55747), .B(n55746), .Z(n63157) );
  IV U75989 ( .A(n55748), .Z(n55749) );
  NOR U75990 ( .A(n55750), .B(n55749), .Z(n63154) );
  IV U75991 ( .A(n55751), .Z(n55753) );
  NOR U75992 ( .A(n55753), .B(n55752), .Z(n63160) );
  NOR U75993 ( .A(n63154), .B(n63160), .Z(n57922) );
  IV U75994 ( .A(n55754), .Z(n55755) );
  NOR U75995 ( .A(n55755), .B(n55758), .Z(n63163) );
  IV U75996 ( .A(n55756), .Z(n55757) );
  NOR U75997 ( .A(n55758), .B(n55757), .Z(n63147) );
  IV U75998 ( .A(n55759), .Z(n55760) );
  NOR U75999 ( .A(n57913), .B(n55760), .Z(n63138) );
  IV U76000 ( .A(n55761), .Z(n55765) );
  NOR U76001 ( .A(n55763), .B(n55762), .Z(n55764) );
  IV U76002 ( .A(n55764), .Z(n55767) );
  NOR U76003 ( .A(n55765), .B(n55767), .Z(n63135) );
  IV U76004 ( .A(n55766), .Z(n55768) );
  NOR U76005 ( .A(n55768), .B(n55767), .Z(n63132) );
  IV U76006 ( .A(n55769), .Z(n55772) );
  IV U76007 ( .A(n55770), .Z(n55771) );
  NOR U76008 ( .A(n55772), .B(n55771), .Z(n63130) );
  NOR U76009 ( .A(n63132), .B(n63130), .Z(n55773) );
  IV U76010 ( .A(n55773), .Z(n57910) );
  IV U76011 ( .A(n55774), .Z(n55775) );
  NOR U76012 ( .A(n55775), .B(n57906), .Z(n60968) );
  IV U76013 ( .A(n55776), .Z(n55777) );
  NOR U76014 ( .A(n55777), .B(n55780), .Z(n63123) );
  IV U76015 ( .A(n55778), .Z(n55779) );
  NOR U76016 ( .A(n55780), .B(n55779), .Z(n63107) );
  IV U76017 ( .A(n55781), .Z(n55785) );
  NOR U76018 ( .A(n55783), .B(n55782), .Z(n55784) );
  IV U76019 ( .A(n55784), .Z(n55789) );
  NOR U76020 ( .A(n55785), .B(n55789), .Z(n63110) );
  IV U76021 ( .A(n55786), .Z(n55787) );
  NOR U76022 ( .A(n57899), .B(n55787), .Z(n66454) );
  IV U76023 ( .A(n55788), .Z(n55790) );
  NOR U76024 ( .A(n55790), .B(n55789), .Z(n68522) );
  NOR U76025 ( .A(n66454), .B(n68522), .Z(n63102) );
  NOR U76026 ( .A(n66466), .B(n55791), .Z(n55792) );
  NOR U76027 ( .A(n55793), .B(n55792), .Z(n63098) );
  IV U76028 ( .A(n55794), .Z(n55797) );
  NOR U76029 ( .A(n55795), .B(n55797), .Z(n68490) );
  IV U76030 ( .A(n55796), .Z(n55800) );
  NOR U76031 ( .A(n55798), .B(n55797), .Z(n55799) );
  IV U76032 ( .A(n55799), .Z(n57855) );
  NOR U76033 ( .A(n55800), .B(n57855), .Z(n68496) );
  NOR U76034 ( .A(n68490), .B(n68496), .Z(n60981) );
  IV U76035 ( .A(n60981), .Z(n57853) );
  IV U76036 ( .A(n55801), .Z(n55802) );
  NOR U76037 ( .A(n55805), .B(n55802), .Z(n60986) );
  IV U76038 ( .A(n55803), .Z(n55804) );
  NOR U76039 ( .A(n55805), .B(n55804), .Z(n63073) );
  IV U76040 ( .A(n55806), .Z(n55808) );
  IV U76041 ( .A(n55807), .Z(n55812) );
  NOR U76042 ( .A(n55808), .B(n55812), .Z(n63067) );
  IV U76043 ( .A(n55809), .Z(n55810) );
  NOR U76044 ( .A(n55810), .B(n55816), .Z(n66490) );
  IV U76045 ( .A(n55811), .Z(n55813) );
  NOR U76046 ( .A(n55813), .B(n55812), .Z(n68483) );
  NOR U76047 ( .A(n66490), .B(n68483), .Z(n63066) );
  IV U76048 ( .A(n55814), .Z(n55815) );
  NOR U76049 ( .A(n55816), .B(n55815), .Z(n55817) );
  IV U76050 ( .A(n55817), .Z(n63059) );
  IV U76051 ( .A(n55818), .Z(n60990) );
  NOR U76052 ( .A(n55819), .B(n60990), .Z(n55823) );
  IV U76053 ( .A(n55820), .Z(n55821) );
  NOR U76054 ( .A(n63051), .B(n55821), .Z(n55822) );
  NOR U76055 ( .A(n55823), .B(n55822), .Z(n57851) );
  NOR U76056 ( .A(n55824), .B(n60995), .Z(n57850) );
  NOR U76057 ( .A(n55826), .B(n55825), .Z(n55827) );
  IV U76058 ( .A(n55827), .Z(n55829) );
  NOR U76059 ( .A(n55828), .B(n55829), .Z(n61004) );
  NOR U76060 ( .A(n55830), .B(n55829), .Z(n61001) );
  IV U76061 ( .A(n55831), .Z(n55833) );
  NOR U76062 ( .A(n55833), .B(n55832), .Z(n61007) );
  IV U76063 ( .A(n55834), .Z(n55836) );
  IV U76064 ( .A(n55835), .Z(n55848) );
  NOR U76065 ( .A(n55836), .B(n55848), .Z(n61015) );
  IV U76066 ( .A(n55837), .Z(n55838) );
  NOR U76067 ( .A(n55841), .B(n55838), .Z(n61011) );
  IV U76068 ( .A(n55839), .Z(n55840) );
  NOR U76069 ( .A(n55841), .B(n55840), .Z(n61013) );
  NOR U76070 ( .A(n61011), .B(n61013), .Z(n55842) );
  IV U76071 ( .A(n55842), .Z(n55843) );
  NOR U76072 ( .A(n61015), .B(n55843), .Z(n57849) );
  IV U76073 ( .A(n55844), .Z(n55846) );
  NOR U76074 ( .A(n55846), .B(n55845), .Z(n63037) );
  IV U76075 ( .A(n55847), .Z(n55849) );
  NOR U76076 ( .A(n55849), .B(n55848), .Z(n61018) );
  NOR U76077 ( .A(n63037), .B(n61018), .Z(n57848) );
  IV U76078 ( .A(n55850), .Z(n55851) );
  NOR U76079 ( .A(n55851), .B(n55857), .Z(n66525) );
  IV U76080 ( .A(n55852), .Z(n57839) );
  IV U76081 ( .A(n55853), .Z(n55854) );
  NOR U76082 ( .A(n57839), .B(n55854), .Z(n66521) );
  NOR U76083 ( .A(n66525), .B(n66521), .Z(n61034) );
  IV U76084 ( .A(n55855), .Z(n55856) );
  NOR U76085 ( .A(n55857), .B(n55856), .Z(n61031) );
  IV U76086 ( .A(n55858), .Z(n55865) );
  NOR U76087 ( .A(n55860), .B(n55859), .Z(n55861) );
  IV U76088 ( .A(n55861), .Z(n55862) );
  NOR U76089 ( .A(n55863), .B(n55862), .Z(n55864) );
  IV U76090 ( .A(n55864), .Z(n55867) );
  NOR U76091 ( .A(n55865), .B(n55867), .Z(n61037) );
  IV U76092 ( .A(n55866), .Z(n55868) );
  NOR U76093 ( .A(n55868), .B(n55867), .Z(n63021) );
  IV U76094 ( .A(n55869), .Z(n55872) );
  IV U76095 ( .A(n55870), .Z(n55871) );
  NOR U76096 ( .A(n55872), .B(n55871), .Z(n61044) );
  IV U76097 ( .A(n55873), .Z(n55875) );
  NOR U76098 ( .A(n55875), .B(n55874), .Z(n61040) );
  NOR U76099 ( .A(n61044), .B(n61040), .Z(n57829) );
  IV U76100 ( .A(n55876), .Z(n55877) );
  NOR U76101 ( .A(n55877), .B(n55879), .Z(n61053) );
  IV U76102 ( .A(n55878), .Z(n55880) );
  NOR U76103 ( .A(n55880), .B(n55879), .Z(n63015) );
  IV U76104 ( .A(n55881), .Z(n55883) );
  NOR U76105 ( .A(n55883), .B(n55882), .Z(n55884) );
  NOR U76106 ( .A(n63015), .B(n55884), .Z(n55885) );
  IV U76107 ( .A(n55885), .Z(n55886) );
  NOR U76108 ( .A(n61053), .B(n55886), .Z(n57827) );
  IV U76109 ( .A(n55887), .Z(n55888) );
  NOR U76110 ( .A(n55894), .B(n55888), .Z(n63006) );
  IV U76111 ( .A(n55889), .Z(n55890) );
  NOR U76112 ( .A(n55890), .B(n61068), .Z(n55891) );
  NOR U76113 ( .A(n63006), .B(n55891), .Z(n61065) );
  IV U76114 ( .A(n55892), .Z(n55893) );
  NOR U76115 ( .A(n55894), .B(n55893), .Z(n62999) );
  IV U76116 ( .A(n55895), .Z(n55897) );
  IV U76117 ( .A(n55896), .Z(n57820) );
  NOR U76118 ( .A(n55897), .B(n57820), .Z(n63003) );
  NOR U76119 ( .A(n62999), .B(n63003), .Z(n57826) );
  IV U76120 ( .A(n55898), .Z(n55900) );
  IV U76121 ( .A(n55899), .Z(n55904) );
  NOR U76122 ( .A(n55900), .B(n55904), .Z(n62985) );
  NOR U76123 ( .A(n55902), .B(n55901), .Z(n62981) );
  IV U76124 ( .A(n55903), .Z(n55905) );
  NOR U76125 ( .A(n55905), .B(n55904), .Z(n62988) );
  NOR U76126 ( .A(n62981), .B(n62988), .Z(n55906) );
  IV U76127 ( .A(n55906), .Z(n57816) );
  IV U76128 ( .A(n55907), .Z(n55911) );
  NOR U76129 ( .A(n55909), .B(n55908), .Z(n55910) );
  IV U76130 ( .A(n55910), .Z(n55914) );
  NOR U76131 ( .A(n55911), .B(n55914), .Z(n55912) );
  IV U76132 ( .A(n55912), .Z(n61073) );
  IV U76133 ( .A(n55913), .Z(n55915) );
  NOR U76134 ( .A(n55915), .B(n55914), .Z(n61074) );
  IV U76135 ( .A(n55916), .Z(n55918) );
  IV U76136 ( .A(n55917), .Z(n55926) );
  NOR U76137 ( .A(n55918), .B(n55926), .Z(n61076) );
  NOR U76138 ( .A(n61074), .B(n61076), .Z(n57815) );
  IV U76139 ( .A(n55919), .Z(n55920) );
  NOR U76140 ( .A(n55920), .B(n55922), .Z(n62973) );
  IV U76141 ( .A(n55921), .Z(n55923) );
  NOR U76142 ( .A(n55923), .B(n55922), .Z(n62970) );
  NOR U76143 ( .A(n62973), .B(n62970), .Z(n55924) );
  IV U76144 ( .A(n55924), .Z(n55928) );
  IV U76145 ( .A(n55925), .Z(n55927) );
  NOR U76146 ( .A(n55927), .B(n55926), .Z(n61079) );
  NOR U76147 ( .A(n55928), .B(n61079), .Z(n57814) );
  IV U76148 ( .A(n55929), .Z(n55931) );
  NOR U76149 ( .A(n55931), .B(n55930), .Z(n66582) );
  IV U76150 ( .A(n55932), .Z(n55934) );
  NOR U76151 ( .A(n55934), .B(n55933), .Z(n66578) );
  NOR U76152 ( .A(n66582), .B(n66578), .Z(n61090) );
  IV U76153 ( .A(n55935), .Z(n55936) );
  NOR U76154 ( .A(n55936), .B(n55938), .Z(n61087) );
  IV U76155 ( .A(n55937), .Z(n55939) );
  NOR U76156 ( .A(n55939), .B(n55938), .Z(n61093) );
  IV U76157 ( .A(n55940), .Z(n55941) );
  NOR U76158 ( .A(n55942), .B(n55941), .Z(n55943) );
  IV U76159 ( .A(n55943), .Z(n57790) );
  IV U76160 ( .A(n55944), .Z(n55945) );
  NOR U76161 ( .A(n55946), .B(n55945), .Z(n61110) );
  IV U76162 ( .A(n55947), .Z(n55949) );
  NOR U76163 ( .A(n55949), .B(n55948), .Z(n61105) );
  NOR U76164 ( .A(n61110), .B(n61105), .Z(n57776) );
  IV U76165 ( .A(n55950), .Z(n55952) );
  NOR U76166 ( .A(n55952), .B(n55951), .Z(n62943) );
  IV U76167 ( .A(n55953), .Z(n55954) );
  NOR U76168 ( .A(n57762), .B(n55954), .Z(n66618) );
  IV U76169 ( .A(n55955), .Z(n55958) );
  IV U76170 ( .A(n55956), .Z(n55957) );
  NOR U76171 ( .A(n55958), .B(n55957), .Z(n66623) );
  NOR U76172 ( .A(n66618), .B(n66623), .Z(n61119) );
  IV U76173 ( .A(n61119), .Z(n57759) );
  IV U76174 ( .A(n55959), .Z(n55961) );
  XOR U76175 ( .A(n55962), .B(n55968), .Z(n55960) );
  NOR U76176 ( .A(n55961), .B(n55960), .Z(n61125) );
  IV U76177 ( .A(n55962), .Z(n55963) );
  NOR U76178 ( .A(n55963), .B(n55968), .Z(n66629) );
  IV U76179 ( .A(n55964), .Z(n57754) );
  IV U76180 ( .A(n55965), .Z(n55966) );
  NOR U76181 ( .A(n57754), .B(n55966), .Z(n66630) );
  IV U76182 ( .A(n55967), .Z(n55969) );
  NOR U76183 ( .A(n55969), .B(n55968), .Z(n61124) );
  NOR U76184 ( .A(n66630), .B(n61124), .Z(n55970) );
  IV U76185 ( .A(n55970), .Z(n55971) );
  NOR U76186 ( .A(n66629), .B(n55971), .Z(n57758) );
  IV U76187 ( .A(n55972), .Z(n55973) );
  NOR U76188 ( .A(n55973), .B(n55978), .Z(n61134) );
  IV U76189 ( .A(n55974), .Z(n55975) );
  NOR U76190 ( .A(n55975), .B(n55980), .Z(n62934) );
  IV U76191 ( .A(n55976), .Z(n55977) );
  NOR U76192 ( .A(n55978), .B(n55977), .Z(n61140) );
  NOR U76193 ( .A(n62934), .B(n61140), .Z(n57747) );
  IV U76194 ( .A(n55979), .Z(n55981) );
  NOR U76195 ( .A(n55981), .B(n55980), .Z(n62931) );
  IV U76196 ( .A(n55982), .Z(n55984) );
  NOR U76197 ( .A(n55984), .B(n55983), .Z(n61148) );
  IV U76198 ( .A(n55985), .Z(n55987) );
  NOR U76199 ( .A(n55987), .B(n55986), .Z(n61150) );
  NOR U76200 ( .A(n61148), .B(n61150), .Z(n57739) );
  IV U76201 ( .A(n55988), .Z(n57735) );
  IV U76202 ( .A(n55989), .Z(n55990) );
  NOR U76203 ( .A(n57735), .B(n55990), .Z(n61154) );
  IV U76204 ( .A(n55991), .Z(n55992) );
  NOR U76205 ( .A(n55993), .B(n55992), .Z(n61160) );
  IV U76206 ( .A(n55994), .Z(n56002) );
  IV U76207 ( .A(n55995), .Z(n55996) );
  NOR U76208 ( .A(n56002), .B(n55996), .Z(n61165) );
  IV U76209 ( .A(n55997), .Z(n55999) );
  NOR U76210 ( .A(n55999), .B(n55998), .Z(n61173) );
  IV U76211 ( .A(n56000), .Z(n56001) );
  NOR U76212 ( .A(n56002), .B(n56001), .Z(n61168) );
  NOR U76213 ( .A(n61173), .B(n61168), .Z(n57730) );
  IV U76214 ( .A(n56003), .Z(n56007) );
  IV U76215 ( .A(n56004), .Z(n56005) );
  NOR U76216 ( .A(n56007), .B(n56005), .Z(n61170) );
  NOR U76217 ( .A(n56007), .B(n56006), .Z(n56008) );
  IV U76218 ( .A(n56008), .Z(n62920) );
  IV U76219 ( .A(n56009), .Z(n56010) );
  NOR U76220 ( .A(n56010), .B(n56015), .Z(n62910) );
  IV U76221 ( .A(n56011), .Z(n56012) );
  NOR U76222 ( .A(n56013), .B(n56012), .Z(n62906) );
  IV U76223 ( .A(n56014), .Z(n56016) );
  NOR U76224 ( .A(n56016), .B(n56015), .Z(n62913) );
  NOR U76225 ( .A(n62906), .B(n62913), .Z(n57722) );
  IV U76226 ( .A(n56017), .Z(n56018) );
  NOR U76227 ( .A(n56021), .B(n56018), .Z(n61179) );
  IV U76228 ( .A(n56019), .Z(n56020) );
  NOR U76229 ( .A(n56021), .B(n56020), .Z(n61183) );
  IV U76230 ( .A(n56022), .Z(n56024) );
  IV U76231 ( .A(n56023), .Z(n56026) );
  NOR U76232 ( .A(n56024), .B(n56026), .Z(n61185) );
  NOR U76233 ( .A(n61183), .B(n61185), .Z(n57714) );
  IV U76234 ( .A(n56025), .Z(n56027) );
  NOR U76235 ( .A(n56027), .B(n56026), .Z(n68313) );
  NOR U76236 ( .A(n68306), .B(n68313), .Z(n61191) );
  IV U76237 ( .A(n56028), .Z(n56030) );
  NOR U76238 ( .A(n56030), .B(n56029), .Z(n61188) );
  NOR U76239 ( .A(n62895), .B(n56031), .Z(n61198) );
  IV U76240 ( .A(n56032), .Z(n57712) );
  NOR U76241 ( .A(n57712), .B(n56033), .Z(n61193) );
  NOR U76242 ( .A(n61198), .B(n61193), .Z(n56034) );
  IV U76243 ( .A(n56034), .Z(n57710) );
  IV U76244 ( .A(n56035), .Z(n56037) );
  IV U76245 ( .A(n56036), .Z(n57708) );
  NOR U76246 ( .A(n56037), .B(n57708), .Z(n62891) );
  IV U76247 ( .A(n56038), .Z(n56040) );
  IV U76248 ( .A(n56039), .Z(n56044) );
  NOR U76249 ( .A(n56040), .B(n56044), .Z(n56041) );
  IV U76250 ( .A(n56041), .Z(n62878) );
  IV U76251 ( .A(n56042), .Z(n56043) );
  NOR U76252 ( .A(n56044), .B(n56043), .Z(n62873) );
  IV U76253 ( .A(n56047), .Z(n56045) );
  NOR U76254 ( .A(n56046), .B(n56045), .Z(n62865) );
  XOR U76255 ( .A(n56047), .B(n56046), .Z(n56050) );
  IV U76256 ( .A(n56048), .Z(n56049) );
  NOR U76257 ( .A(n56050), .B(n56049), .Z(n62870) );
  NOR U76258 ( .A(n62865), .B(n62870), .Z(n57702) );
  IV U76259 ( .A(n56051), .Z(n56053) );
  NOR U76260 ( .A(n56053), .B(n56052), .Z(n68293) );
  IV U76261 ( .A(n56054), .Z(n56056) );
  NOR U76262 ( .A(n56056), .B(n56055), .Z(n68299) );
  NOR U76263 ( .A(n68293), .B(n68299), .Z(n62864) );
  IV U76264 ( .A(n56057), .Z(n56059) );
  NOR U76265 ( .A(n56059), .B(n56058), .Z(n62848) );
  IV U76266 ( .A(n56060), .Z(n56061) );
  NOR U76267 ( .A(n56061), .B(n62855), .Z(n56062) );
  NOR U76268 ( .A(n62848), .B(n56062), .Z(n57701) );
  IV U76269 ( .A(n68276), .Z(n56063) );
  NOR U76270 ( .A(n56063), .B(n68275), .Z(n62843) );
  IV U76271 ( .A(n56064), .Z(n56065) );
  NOR U76272 ( .A(n56066), .B(n56065), .Z(n57690) );
  IV U76273 ( .A(n56067), .Z(n61209) );
  NOR U76274 ( .A(n56068), .B(n61209), .Z(n57679) );
  IV U76275 ( .A(n56069), .Z(n56070) );
  NOR U76276 ( .A(n56070), .B(n57677), .Z(n61213) );
  IV U76277 ( .A(n56071), .Z(n56072) );
  NOR U76278 ( .A(n57677), .B(n56072), .Z(n56073) );
  IV U76279 ( .A(n56073), .Z(n61222) );
  IV U76280 ( .A(n56074), .Z(n56075) );
  NOR U76281 ( .A(n56075), .B(n56080), .Z(n61224) );
  IV U76282 ( .A(n56076), .Z(n57667) );
  IV U76283 ( .A(n56077), .Z(n56078) );
  NOR U76284 ( .A(n57667), .B(n56078), .Z(n61229) );
  IV U76285 ( .A(n56079), .Z(n56081) );
  NOR U76286 ( .A(n56081), .B(n56080), .Z(n62832) );
  NOR U76287 ( .A(n61229), .B(n62832), .Z(n57671) );
  IV U76288 ( .A(n56082), .Z(n56085) );
  NOR U76289 ( .A(n56087), .B(n56083), .Z(n56084) );
  IV U76290 ( .A(n56084), .Z(n57669) );
  NOR U76291 ( .A(n56085), .B(n57669), .Z(n61236) );
  IV U76292 ( .A(n56086), .Z(n56088) );
  NOR U76293 ( .A(n56088), .B(n56087), .Z(n56089) );
  IV U76294 ( .A(n56089), .Z(n61234) );
  IV U76295 ( .A(n56090), .Z(n56091) );
  NOR U76296 ( .A(n56092), .B(n56091), .Z(n61239) );
  IV U76297 ( .A(n56093), .Z(n56095) );
  IV U76298 ( .A(n56094), .Z(n56097) );
  NOR U76299 ( .A(n56095), .B(n56097), .Z(n62823) );
  NOR U76300 ( .A(n61239), .B(n62823), .Z(n57664) );
  IV U76301 ( .A(n56096), .Z(n56103) );
  NOR U76302 ( .A(n56098), .B(n56097), .Z(n56099) );
  IV U76303 ( .A(n56099), .Z(n56100) );
  NOR U76304 ( .A(n56101), .B(n56100), .Z(n56102) );
  IV U76305 ( .A(n56102), .Z(n56105) );
  NOR U76306 ( .A(n56103), .B(n56105), .Z(n62819) );
  IV U76307 ( .A(n56104), .Z(n56106) );
  NOR U76308 ( .A(n56106), .B(n56105), .Z(n62816) );
  IV U76309 ( .A(n56107), .Z(n56109) );
  NOR U76310 ( .A(n56109), .B(n56108), .Z(n61241) );
  IV U76311 ( .A(n56110), .Z(n56112) );
  NOR U76312 ( .A(n56112), .B(n56111), .Z(n66778) );
  IV U76313 ( .A(n56113), .Z(n56114) );
  NOR U76314 ( .A(n56114), .B(n57661), .Z(n66772) );
  NOR U76315 ( .A(n66778), .B(n66772), .Z(n62812) );
  IV U76316 ( .A(n56115), .Z(n56116) );
  NOR U76317 ( .A(n56116), .B(n57646), .Z(n56117) );
  IV U76318 ( .A(n56117), .Z(n56118) );
  NOR U76319 ( .A(n57649), .B(n56118), .Z(n62809) );
  IV U76320 ( .A(n56119), .Z(n56125) );
  NOR U76321 ( .A(n56120), .B(n56130), .Z(n56121) );
  IV U76322 ( .A(n56121), .Z(n56122) );
  NOR U76323 ( .A(n56123), .B(n56122), .Z(n56124) );
  IV U76324 ( .A(n56124), .Z(n57636) );
  NOR U76325 ( .A(n56125), .B(n57636), .Z(n61266) );
  IV U76326 ( .A(n56126), .Z(n56127) );
  NOR U76327 ( .A(n56128), .B(n56127), .Z(n61274) );
  IV U76328 ( .A(n56129), .Z(n56131) );
  NOR U76329 ( .A(n56131), .B(n56130), .Z(n61269) );
  NOR U76330 ( .A(n61274), .B(n61269), .Z(n57633) );
  IV U76331 ( .A(n56132), .Z(n56133) );
  NOR U76332 ( .A(n56134), .B(n56133), .Z(n61271) );
  IV U76333 ( .A(n57629), .Z(n56135) );
  NOR U76334 ( .A(n56135), .B(n57628), .Z(n57622) );
  IV U76335 ( .A(n57622), .Z(n57617) );
  IV U76336 ( .A(n56136), .Z(n56137) );
  NOR U76337 ( .A(n56137), .B(n57611), .Z(n62792) );
  IV U76338 ( .A(n56138), .Z(n56140) );
  NOR U76339 ( .A(n56140), .B(n56139), .Z(n66827) );
  IV U76340 ( .A(n56141), .Z(n56142) );
  NOR U76341 ( .A(n56143), .B(n56142), .Z(n66823) );
  NOR U76342 ( .A(n66827), .B(n66823), .Z(n61296) );
  IV U76343 ( .A(n56144), .Z(n56151) );
  NOR U76344 ( .A(n56146), .B(n56145), .Z(n56147) );
  IV U76345 ( .A(n56147), .Z(n56148) );
  NOR U76346 ( .A(n56149), .B(n56148), .Z(n56150) );
  IV U76347 ( .A(n56150), .Z(n56156) );
  NOR U76348 ( .A(n56151), .B(n56156), .Z(n56152) );
  IV U76349 ( .A(n56152), .Z(n62749) );
  IV U76350 ( .A(n56153), .Z(n56154) );
  IV U76351 ( .A(n57565), .Z(n57563) );
  NOR U76352 ( .A(n56154), .B(n57563), .Z(n66847) );
  IV U76353 ( .A(n56155), .Z(n56157) );
  NOR U76354 ( .A(n56157), .B(n56156), .Z(n68190) );
  NOR U76355 ( .A(n66847), .B(n68190), .Z(n62747) );
  IV U76356 ( .A(n56158), .Z(n56159) );
  NOR U76357 ( .A(n56159), .B(n56161), .Z(n61319) );
  IV U76358 ( .A(n56160), .Z(n56162) );
  NOR U76359 ( .A(n56162), .B(n56161), .Z(n62741) );
  IV U76360 ( .A(n56163), .Z(n56167) );
  NOR U76361 ( .A(n56172), .B(n56164), .Z(n56165) );
  IV U76362 ( .A(n56165), .Z(n56166) );
  NOR U76363 ( .A(n56167), .B(n56166), .Z(n62738) );
  IV U76364 ( .A(n56168), .Z(n56169) );
  NOR U76365 ( .A(n56171), .B(n56169), .Z(n61328) );
  IV U76366 ( .A(n56170), .Z(n56175) );
  NOR U76367 ( .A(n56172), .B(n56171), .Z(n56173) );
  IV U76368 ( .A(n56173), .Z(n56174) );
  NOR U76369 ( .A(n56175), .B(n56174), .Z(n61325) );
  NOR U76370 ( .A(n61328), .B(n61325), .Z(n57561) );
  IV U76371 ( .A(n56176), .Z(n56185) );
  IV U76372 ( .A(n56177), .Z(n56178) );
  NOR U76373 ( .A(n56185), .B(n56178), .Z(n62735) );
  IV U76374 ( .A(n56179), .Z(n56180) );
  NOR U76375 ( .A(n56185), .B(n56180), .Z(n66865) );
  NOR U76376 ( .A(n62735), .B(n66865), .Z(n57560) );
  IV U76377 ( .A(n56181), .Z(n56182) );
  NOR U76378 ( .A(n56182), .B(n56188), .Z(n66872) );
  IV U76379 ( .A(n56183), .Z(n56184) );
  NOR U76380 ( .A(n56185), .B(n56184), .Z(n66870) );
  NOR U76381 ( .A(n66872), .B(n66870), .Z(n56186) );
  IV U76382 ( .A(n56186), .Z(n62732) );
  IV U76383 ( .A(n56187), .Z(n56189) );
  NOR U76384 ( .A(n56189), .B(n56188), .Z(n62728) );
  IV U76385 ( .A(n56190), .Z(n56195) );
  NOR U76386 ( .A(n56200), .B(n56202), .Z(n56191) );
  IV U76387 ( .A(n56191), .Z(n56192) );
  NOR U76388 ( .A(n56193), .B(n56192), .Z(n56194) );
  IV U76389 ( .A(n56194), .Z(n56197) );
  NOR U76390 ( .A(n56195), .B(n56197), .Z(n62725) );
  IV U76391 ( .A(n56196), .Z(n56198) );
  NOR U76392 ( .A(n56198), .B(n56197), .Z(n62721) );
  NOR U76393 ( .A(n56200), .B(n56199), .Z(n56201) );
  IV U76394 ( .A(n56201), .Z(n56203) );
  NOR U76395 ( .A(n56203), .B(n56202), .Z(n62718) );
  IV U76396 ( .A(n56204), .Z(n56206) );
  NOR U76397 ( .A(n56206), .B(n56205), .Z(n62709) );
  IV U76398 ( .A(n56207), .Z(n56208) );
  NOR U76399 ( .A(n56209), .B(n56208), .Z(n62715) );
  NOR U76400 ( .A(n62709), .B(n62715), .Z(n56210) );
  IV U76401 ( .A(n56210), .Z(n57559) );
  IV U76402 ( .A(n56211), .Z(n56212) );
  NOR U76403 ( .A(n56213), .B(n56212), .Z(n62704) );
  IV U76404 ( .A(n56214), .Z(n56216) );
  NOR U76405 ( .A(n56216), .B(n56215), .Z(n62711) );
  NOR U76406 ( .A(n62704), .B(n62711), .Z(n57558) );
  IV U76407 ( .A(n56217), .Z(n56220) );
  IV U76408 ( .A(n56219), .Z(n56218) );
  NOR U76409 ( .A(n56220), .B(n56218), .Z(n68158) );
  XOR U76410 ( .A(n56220), .B(n56219), .Z(n56221) );
  NOR U76411 ( .A(n56222), .B(n56221), .Z(n56223) );
  IV U76412 ( .A(n56223), .Z(n56224) );
  NOR U76413 ( .A(n56225), .B(n56224), .Z(n68164) );
  NOR U76414 ( .A(n68158), .B(n68164), .Z(n62703) );
  IV U76415 ( .A(n56226), .Z(n56227) );
  NOR U76416 ( .A(n57557), .B(n56227), .Z(n61331) );
  IV U76417 ( .A(n56228), .Z(n56229) );
  NOR U76418 ( .A(n57557), .B(n56229), .Z(n61338) );
  IV U76419 ( .A(n56230), .Z(n56233) );
  IV U76420 ( .A(n56231), .Z(n56232) );
  NOR U76421 ( .A(n56233), .B(n56232), .Z(n62699) );
  NOR U76422 ( .A(n61338), .B(n62699), .Z(n57553) );
  IV U76423 ( .A(n56234), .Z(n56236) );
  XOR U76424 ( .A(n56242), .B(n56243), .Z(n56235) );
  NOR U76425 ( .A(n56236), .B(n56235), .Z(n62695) );
  IV U76426 ( .A(n56237), .Z(n56238) );
  NOR U76427 ( .A(n56238), .B(n56243), .Z(n62692) );
  IV U76428 ( .A(n56239), .Z(n56241) );
  NOR U76429 ( .A(n56241), .B(n56240), .Z(n68138) );
  IV U76430 ( .A(n56242), .Z(n56244) );
  NOR U76431 ( .A(n56244), .B(n56243), .Z(n66901) );
  NOR U76432 ( .A(n68138), .B(n66901), .Z(n62681) );
  IV U76433 ( .A(n56245), .Z(n56246) );
  NOR U76434 ( .A(n56247), .B(n56246), .Z(n62685) );
  IV U76435 ( .A(n56248), .Z(n56250) );
  NOR U76436 ( .A(n56250), .B(n56249), .Z(n62683) );
  NOR U76437 ( .A(n62685), .B(n62683), .Z(n57552) );
  IV U76438 ( .A(n56251), .Z(n56252) );
  NOR U76439 ( .A(n56252), .B(n62659), .Z(n62673) );
  NOR U76440 ( .A(n62659), .B(n56253), .Z(n56254) );
  IV U76441 ( .A(n56254), .Z(n57551) );
  IV U76442 ( .A(n56255), .Z(n56257) );
  NOR U76443 ( .A(n56257), .B(n56256), .Z(n62642) );
  IV U76444 ( .A(n56258), .Z(n56259) );
  NOR U76445 ( .A(n57517), .B(n56259), .Z(n62644) );
  NOR U76446 ( .A(n62642), .B(n62644), .Z(n57519) );
  IV U76447 ( .A(n68093), .Z(n56260) );
  NOR U76448 ( .A(n56260), .B(n68092), .Z(n62633) );
  IV U76449 ( .A(n56261), .Z(n56262) );
  NOR U76450 ( .A(n56263), .B(n56262), .Z(n68083) );
  NOR U76451 ( .A(n66921), .B(n68083), .Z(n62627) );
  IV U76452 ( .A(n56264), .Z(n56265) );
  NOR U76453 ( .A(n56271), .B(n56265), .Z(n56266) );
  IV U76454 ( .A(n56266), .Z(n62626) );
  IV U76455 ( .A(n56267), .Z(n56269) );
  NOR U76456 ( .A(n56269), .B(n56268), .Z(n62616) );
  IV U76457 ( .A(n56270), .Z(n56272) );
  NOR U76458 ( .A(n56272), .B(n56271), .Z(n61358) );
  NOR U76459 ( .A(n62616), .B(n61358), .Z(n57509) );
  IV U76460 ( .A(n56273), .Z(n61368) );
  NOR U76461 ( .A(n57504), .B(n61368), .Z(n56277) );
  IV U76462 ( .A(n56274), .Z(n56276) );
  NOR U76463 ( .A(n56276), .B(n56275), .Z(n62619) );
  NOR U76464 ( .A(n56277), .B(n62619), .Z(n57508) );
  IV U76465 ( .A(n56278), .Z(n56280) );
  IV U76466 ( .A(n56279), .Z(n61377) );
  NOR U76467 ( .A(n56280), .B(n61377), .Z(n56281) );
  IV U76468 ( .A(n56281), .Z(n61370) );
  IV U76469 ( .A(n56283), .Z(n56290) );
  XOR U76470 ( .A(n56291), .B(n56290), .Z(n56285) );
  IV U76471 ( .A(n56282), .Z(n56288) );
  NOR U76472 ( .A(n56283), .B(n56288), .Z(n56284) );
  NOR U76473 ( .A(n56285), .B(n56284), .Z(n56287) );
  NOR U76474 ( .A(n56287), .B(n56286), .Z(n56289) );
  NOR U76475 ( .A(n56291), .B(n56288), .Z(n62607) );
  NOR U76476 ( .A(n56289), .B(n62607), .Z(n57502) );
  NOR U76477 ( .A(n56291), .B(n56290), .Z(n56292) );
  IV U76478 ( .A(n56292), .Z(n62606) );
  IV U76479 ( .A(n56293), .Z(n56294) );
  NOR U76480 ( .A(n56295), .B(n56294), .Z(n57498) );
  IV U76481 ( .A(n56296), .Z(n56297) );
  NOR U76482 ( .A(n56298), .B(n56297), .Z(n62592) );
  IV U76483 ( .A(n56299), .Z(n56300) );
  NOR U76484 ( .A(n56300), .B(n57489), .Z(n56301) );
  IV U76485 ( .A(n56301), .Z(n62583) );
  IV U76486 ( .A(n56302), .Z(n56304) );
  IV U76487 ( .A(n56303), .Z(n57456) );
  NOR U76488 ( .A(n56304), .B(n57456), .Z(n56305) );
  IV U76489 ( .A(n56305), .Z(n57462) );
  IV U76490 ( .A(n56306), .Z(n56307) );
  NOR U76491 ( .A(n56308), .B(n56307), .Z(n56309) );
  IV U76492 ( .A(n56309), .Z(n62548) );
  IV U76493 ( .A(n56310), .Z(n56311) );
  NOR U76494 ( .A(n56311), .B(n56313), .Z(n67994) );
  IV U76495 ( .A(n56312), .Z(n56314) );
  NOR U76496 ( .A(n56314), .B(n56313), .Z(n68002) );
  NOR U76497 ( .A(n67994), .B(n68002), .Z(n62532) );
  IV U76498 ( .A(n56315), .Z(n56317) );
  NOR U76499 ( .A(n56317), .B(n56316), .Z(n61402) );
  IV U76500 ( .A(n56318), .Z(n56319) );
  NOR U76501 ( .A(n56320), .B(n56319), .Z(n61396) );
  NOR U76502 ( .A(n61402), .B(n61396), .Z(n57424) );
  IV U76503 ( .A(n56321), .Z(n56323) );
  NOR U76504 ( .A(n56323), .B(n56322), .Z(n57420) );
  IV U76505 ( .A(n56324), .Z(n61415) );
  IV U76506 ( .A(n56325), .Z(n56326) );
  NOR U76507 ( .A(n61415), .B(n56326), .Z(n61411) );
  IV U76508 ( .A(n56327), .Z(n56329) );
  NOR U76509 ( .A(n56329), .B(n56328), .Z(n61408) );
  NOR U76510 ( .A(n61411), .B(n61408), .Z(n57397) );
  NOR U76511 ( .A(n56330), .B(n61415), .Z(n57396) );
  IV U76512 ( .A(n56331), .Z(n56333) );
  NOR U76513 ( .A(n56333), .B(n56332), .Z(n61418) );
  IV U76514 ( .A(n56334), .Z(n56335) );
  NOR U76515 ( .A(n56336), .B(n56335), .Z(n66995) );
  IV U76516 ( .A(n56337), .Z(n56338) );
  NOR U76517 ( .A(n56339), .B(n56338), .Z(n66987) );
  NOR U76518 ( .A(n66995), .B(n66987), .Z(n62510) );
  IV U76519 ( .A(n56340), .Z(n56342) );
  IV U76520 ( .A(n56341), .Z(n56344) );
  NOR U76521 ( .A(n56342), .B(n56344), .Z(n62507) );
  IV U76522 ( .A(n56343), .Z(n56347) );
  NOR U76523 ( .A(n56345), .B(n56344), .Z(n56346) );
  IV U76524 ( .A(n56346), .Z(n56349) );
  NOR U76525 ( .A(n56347), .B(n56349), .Z(n61425) );
  IV U76526 ( .A(n56348), .Z(n56350) );
  NOR U76527 ( .A(n56350), .B(n56349), .Z(n62500) );
  IV U76528 ( .A(n56351), .Z(n56352) );
  NOR U76529 ( .A(n56355), .B(n56352), .Z(n61428) );
  IV U76530 ( .A(n56353), .Z(n56354) );
  NOR U76531 ( .A(n56355), .B(n56354), .Z(n62483) );
  IV U76532 ( .A(n56356), .Z(n56363) );
  XOR U76533 ( .A(n56364), .B(n56365), .Z(n56357) );
  NOR U76534 ( .A(n56358), .B(n56357), .Z(n56359) );
  IV U76535 ( .A(n56359), .Z(n56360) );
  NOR U76536 ( .A(n56361), .B(n56360), .Z(n56362) );
  IV U76537 ( .A(n56362), .Z(n56368) );
  NOR U76538 ( .A(n56363), .B(n56368), .Z(n62480) );
  IV U76539 ( .A(n56364), .Z(n56366) );
  NOR U76540 ( .A(n56366), .B(n56365), .Z(n67932) );
  IV U76541 ( .A(n56367), .Z(n56369) );
  NOR U76542 ( .A(n56369), .B(n56368), .Z(n67937) );
  NOR U76543 ( .A(n67932), .B(n67937), .Z(n61432) );
  IV U76544 ( .A(n56370), .Z(n56372) );
  NOR U76545 ( .A(n56372), .B(n56371), .Z(n61438) );
  IV U76546 ( .A(n56373), .Z(n56374) );
  NOR U76547 ( .A(n56375), .B(n56374), .Z(n61433) );
  NOR U76548 ( .A(n61438), .B(n61433), .Z(n57391) );
  IV U76549 ( .A(n56376), .Z(n56378) );
  NOR U76550 ( .A(n56378), .B(n56377), .Z(n61436) );
  IV U76551 ( .A(n56379), .Z(n56380) );
  NOR U76552 ( .A(n56381), .B(n56380), .Z(n61445) );
  IV U76553 ( .A(n56382), .Z(n56384) );
  NOR U76554 ( .A(n56384), .B(n56383), .Z(n62469) );
  NOR U76555 ( .A(n61445), .B(n62469), .Z(n57383) );
  IV U76556 ( .A(n56385), .Z(n67014) );
  NOR U76557 ( .A(n67014), .B(n56386), .Z(n56387) );
  IV U76558 ( .A(n56387), .Z(n57371) );
  IV U76559 ( .A(n56388), .Z(n56389) );
  NOR U76560 ( .A(n56393), .B(n56389), .Z(n56390) );
  IV U76561 ( .A(n56390), .Z(n61469) );
  IV U76562 ( .A(n56391), .Z(n56392) );
  NOR U76563 ( .A(n56393), .B(n56392), .Z(n61471) );
  IV U76564 ( .A(n56394), .Z(n56396) );
  IV U76565 ( .A(n56395), .Z(n56398) );
  NOR U76566 ( .A(n56396), .B(n56398), .Z(n61474) );
  NOR U76567 ( .A(n61471), .B(n61474), .Z(n57352) );
  IV U76568 ( .A(n56397), .Z(n56399) );
  NOR U76569 ( .A(n56399), .B(n56398), .Z(n61480) );
  IV U76570 ( .A(n56400), .Z(n56401) );
  NOR U76571 ( .A(n56404), .B(n56401), .Z(n61477) );
  IV U76572 ( .A(n56402), .Z(n56403) );
  NOR U76573 ( .A(n56404), .B(n56403), .Z(n61484) );
  IV U76574 ( .A(n56405), .Z(n56409) );
  NOR U76575 ( .A(n56407), .B(n56406), .Z(n56408) );
  IV U76576 ( .A(n56408), .Z(n56414) );
  NOR U76577 ( .A(n56409), .B(n56414), .Z(n61486) );
  NOR U76578 ( .A(n61484), .B(n61486), .Z(n57351) );
  IV U76579 ( .A(n56410), .Z(n56411) );
  NOR U76580 ( .A(n56412), .B(n56411), .Z(n61498) );
  IV U76581 ( .A(n56413), .Z(n56415) );
  NOR U76582 ( .A(n56415), .B(n56414), .Z(n61489) );
  NOR U76583 ( .A(n61498), .B(n61489), .Z(n57350) );
  IV U76584 ( .A(n56416), .Z(n56418) );
  NOR U76585 ( .A(n56418), .B(n56417), .Z(n61492) );
  IV U76586 ( .A(n56419), .Z(n56421) );
  NOR U76587 ( .A(n56421), .B(n56420), .Z(n61494) );
  NOR U76588 ( .A(n61492), .B(n61494), .Z(n57349) );
  IV U76589 ( .A(n56422), .Z(n56423) );
  NOR U76590 ( .A(n56424), .B(n56423), .Z(n61502) );
  IV U76591 ( .A(n56425), .Z(n56432) );
  NOR U76592 ( .A(n56427), .B(n56426), .Z(n56428) );
  IV U76593 ( .A(n56428), .Z(n56429) );
  NOR U76594 ( .A(n56430), .B(n56429), .Z(n56431) );
  IV U76595 ( .A(n56431), .Z(n57346) );
  NOR U76596 ( .A(n56432), .B(n57346), .Z(n62446) );
  NOR U76597 ( .A(n61502), .B(n62446), .Z(n57348) );
  IV U76598 ( .A(n56433), .Z(n56434) );
  NOR U76599 ( .A(n56435), .B(n56434), .Z(n67879) );
  IV U76600 ( .A(n56436), .Z(n56437) );
  NOR U76601 ( .A(n56438), .B(n56437), .Z(n67884) );
  NOR U76602 ( .A(n67879), .B(n67884), .Z(n61511) );
  IV U76603 ( .A(n56439), .Z(n56440) );
  NOR U76604 ( .A(n56440), .B(n56446), .Z(n56441) );
  IV U76605 ( .A(n56441), .Z(n61509) );
  IV U76606 ( .A(n56442), .Z(n56444) );
  NOR U76607 ( .A(n56444), .B(n56443), .Z(n67872) );
  IV U76608 ( .A(n56445), .Z(n56447) );
  NOR U76609 ( .A(n56447), .B(n56446), .Z(n67876) );
  NOR U76610 ( .A(n67872), .B(n67876), .Z(n62422) );
  IV U76611 ( .A(n56448), .Z(n56450) );
  NOR U76612 ( .A(n56450), .B(n56449), .Z(n62403) );
  IV U76613 ( .A(n56451), .Z(n56453) );
  IV U76614 ( .A(n56452), .Z(n57324) );
  NOR U76615 ( .A(n56453), .B(n57324), .Z(n62401) );
  NOR U76616 ( .A(n62403), .B(n62401), .Z(n57321) );
  IV U76617 ( .A(n56454), .Z(n56456) );
  NOR U76618 ( .A(n56456), .B(n56455), .Z(n67848) );
  NOR U76619 ( .A(n67848), .B(n67856), .Z(n62400) );
  IV U76620 ( .A(n56457), .Z(n56464) );
  NOR U76621 ( .A(n56459), .B(n56458), .Z(n56460) );
  IV U76622 ( .A(n56460), .Z(n56461) );
  NOR U76623 ( .A(n56462), .B(n56461), .Z(n56463) );
  IV U76624 ( .A(n56463), .Z(n56466) );
  NOR U76625 ( .A(n56464), .B(n56466), .Z(n61522) );
  IV U76626 ( .A(n56465), .Z(n56467) );
  NOR U76627 ( .A(n56467), .B(n56466), .Z(n61523) );
  NOR U76628 ( .A(n61522), .B(n61523), .Z(n57320) );
  IV U76629 ( .A(n56468), .Z(n56469) );
  NOR U76630 ( .A(n56469), .B(n56478), .Z(n61529) );
  IV U76631 ( .A(n56470), .Z(n56472) );
  NOR U76632 ( .A(n56472), .B(n56471), .Z(n61527) );
  NOR U76633 ( .A(n61529), .B(n61527), .Z(n57319) );
  IV U76634 ( .A(n56473), .Z(n56474) );
  NOR U76635 ( .A(n56475), .B(n56474), .Z(n61534) );
  IV U76636 ( .A(n56476), .Z(n56477) );
  NOR U76637 ( .A(n56478), .B(n56477), .Z(n61532) );
  NOR U76638 ( .A(n61534), .B(n61532), .Z(n57318) );
  IV U76639 ( .A(n56479), .Z(n56480) );
  NOR U76640 ( .A(n56480), .B(n56482), .Z(n61541) );
  IV U76641 ( .A(n56481), .Z(n56483) );
  NOR U76642 ( .A(n56483), .B(n56482), .Z(n56484) );
  IV U76643 ( .A(n56484), .Z(n61539) );
  IV U76644 ( .A(n56485), .Z(n56492) );
  NOR U76645 ( .A(n56487), .B(n56486), .Z(n56488) );
  IV U76646 ( .A(n56488), .Z(n56489) );
  NOR U76647 ( .A(n56490), .B(n56489), .Z(n56491) );
  IV U76648 ( .A(n56491), .Z(n56494) );
  NOR U76649 ( .A(n56492), .B(n56494), .Z(n62391) );
  IV U76650 ( .A(n56493), .Z(n56495) );
  NOR U76651 ( .A(n56495), .B(n56494), .Z(n62389) );
  IV U76652 ( .A(n56496), .Z(n56497) );
  NOR U76653 ( .A(n56503), .B(n56497), .Z(n62384) );
  IV U76654 ( .A(n56498), .Z(n56500) );
  NOR U76655 ( .A(n56500), .B(n56499), .Z(n62386) );
  NOR U76656 ( .A(n62384), .B(n62386), .Z(n57310) );
  IV U76657 ( .A(n56501), .Z(n56502) );
  NOR U76658 ( .A(n56503), .B(n56502), .Z(n61547) );
  IV U76659 ( .A(n56504), .Z(n56509) );
  IV U76660 ( .A(n56505), .Z(n56506) );
  NOR U76661 ( .A(n56509), .B(n56506), .Z(n61549) );
  NOR U76662 ( .A(n61547), .B(n61549), .Z(n57309) );
  NOR U76663 ( .A(n56507), .B(n61556), .Z(n56511) );
  IV U76664 ( .A(n56508), .Z(n56510) );
  NOR U76665 ( .A(n56510), .B(n56509), .Z(n61552) );
  NOR U76666 ( .A(n56511), .B(n61552), .Z(n57308) );
  IV U76667 ( .A(n56512), .Z(n56514) );
  IV U76668 ( .A(n56513), .Z(n57305) );
  NOR U76669 ( .A(n56514), .B(n57305), .Z(n61562) );
  IV U76670 ( .A(n56515), .Z(n56516) );
  NOR U76671 ( .A(n56516), .B(n57302), .Z(n57299) );
  IV U76672 ( .A(n56517), .Z(n56519) );
  NOR U76673 ( .A(n56519), .B(n56518), .Z(n56520) );
  IV U76674 ( .A(n56520), .Z(n61569) );
  IV U76675 ( .A(n56521), .Z(n56523) );
  NOR U76676 ( .A(n56523), .B(n56522), .Z(n62374) );
  IV U76677 ( .A(n56524), .Z(n56526) );
  NOR U76678 ( .A(n56526), .B(n56525), .Z(n61571) );
  NOR U76679 ( .A(n62374), .B(n61571), .Z(n57296) );
  IV U76680 ( .A(n56527), .Z(n56528) );
  NOR U76681 ( .A(n56529), .B(n56528), .Z(n56530) );
  IV U76682 ( .A(n56530), .Z(n56536) );
  IV U76683 ( .A(n56531), .Z(n56533) );
  NOR U76684 ( .A(n56533), .B(n56532), .Z(n56534) );
  IV U76685 ( .A(n56534), .Z(n56535) );
  NOR U76686 ( .A(n56536), .B(n56535), .Z(n61573) );
  NOR U76687 ( .A(n56547), .B(n56537), .Z(n56538) );
  IV U76688 ( .A(n56538), .Z(n56544) );
  IV U76689 ( .A(n56539), .Z(n56541) );
  NOR U76690 ( .A(n56541), .B(n56540), .Z(n56542) );
  IV U76691 ( .A(n56542), .Z(n56543) );
  NOR U76692 ( .A(n56544), .B(n56543), .Z(n62366) );
  IV U76693 ( .A(n56545), .Z(n56546) );
  NOR U76694 ( .A(n56547), .B(n56546), .Z(n61576) );
  IV U76695 ( .A(n56548), .Z(n56549) );
  NOR U76696 ( .A(n56552), .B(n56549), .Z(n62350) );
  IV U76697 ( .A(n56550), .Z(n56551) );
  NOR U76698 ( .A(n56552), .B(n56551), .Z(n62347) );
  IV U76699 ( .A(n56553), .Z(n56555) );
  NOR U76700 ( .A(n56555), .B(n56554), .Z(n61580) );
  IV U76701 ( .A(n56556), .Z(n56557) );
  NOR U76702 ( .A(n56558), .B(n56557), .Z(n62344) );
  NOR U76703 ( .A(n61580), .B(n62344), .Z(n57295) );
  IV U76704 ( .A(n56559), .Z(n56560) );
  NOR U76705 ( .A(n56561), .B(n56560), .Z(n62341) );
  IV U76706 ( .A(n56562), .Z(n56563) );
  NOR U76707 ( .A(n56570), .B(n56563), .Z(n62339) );
  NOR U76708 ( .A(n62341), .B(n62339), .Z(n57294) );
  NOR U76709 ( .A(n56564), .B(n56572), .Z(n56565) );
  IV U76710 ( .A(n56565), .Z(n56568) );
  IV U76711 ( .A(n56566), .Z(n56567) );
  NOR U76712 ( .A(n56568), .B(n56567), .Z(n61585) );
  NOR U76713 ( .A(n56570), .B(n56569), .Z(n61582) );
  IV U76714 ( .A(n56571), .Z(n56575) );
  NOR U76715 ( .A(n56573), .B(n56572), .Z(n56574) );
  IV U76716 ( .A(n56574), .Z(n57291) );
  NOR U76717 ( .A(n56575), .B(n57291), .Z(n62335) );
  IV U76718 ( .A(n56576), .Z(n56577) );
  NOR U76719 ( .A(n56577), .B(n56583), .Z(n56578) );
  IV U76720 ( .A(n56578), .Z(n61592) );
  IV U76721 ( .A(n56579), .Z(n56580) );
  NOR U76722 ( .A(n62312), .B(n56580), .Z(n61596) );
  IV U76723 ( .A(n56581), .Z(n56582) );
  NOR U76724 ( .A(n56583), .B(n56582), .Z(n61594) );
  NOR U76725 ( .A(n61596), .B(n61594), .Z(n57278) );
  IV U76726 ( .A(n56584), .Z(n56585) );
  NOR U76727 ( .A(n56586), .B(n56585), .Z(n56587) );
  IV U76728 ( .A(n56587), .Z(n57276) );
  NOR U76729 ( .A(n56588), .B(n57276), .Z(n62309) );
  IV U76730 ( .A(n56589), .Z(n56591) );
  NOR U76731 ( .A(n56591), .B(n56590), .Z(n67136) );
  IV U76732 ( .A(n56592), .Z(n56598) );
  NOR U76733 ( .A(n56593), .B(n56600), .Z(n56594) );
  IV U76734 ( .A(n56594), .Z(n56595) );
  NOR U76735 ( .A(n56596), .B(n56595), .Z(n56597) );
  IV U76736 ( .A(n56597), .Z(n56603) );
  NOR U76737 ( .A(n56598), .B(n56603), .Z(n67140) );
  NOR U76738 ( .A(n67136), .B(n67140), .Z(n62302) );
  IV U76739 ( .A(n56599), .Z(n56601) );
  NOR U76740 ( .A(n56601), .B(n56600), .Z(n61603) );
  IV U76741 ( .A(n56602), .Z(n56604) );
  NOR U76742 ( .A(n56604), .B(n56603), .Z(n61601) );
  NOR U76743 ( .A(n61603), .B(n61601), .Z(n57273) );
  NOR U76744 ( .A(n56605), .B(n61610), .Z(n56608) );
  IV U76745 ( .A(n56606), .Z(n56607) );
  NOR U76746 ( .A(n56607), .B(n61610), .Z(n61606) );
  NOR U76747 ( .A(n56608), .B(n61606), .Z(n57272) );
  IV U76748 ( .A(n56609), .Z(n56613) );
  NOR U76749 ( .A(n56611), .B(n56610), .Z(n56612) );
  IV U76750 ( .A(n56612), .Z(n56619) );
  NOR U76751 ( .A(n56613), .B(n56619), .Z(n56614) );
  IV U76752 ( .A(n56614), .Z(n62293) );
  IV U76753 ( .A(n56615), .Z(n56616) );
  NOR U76754 ( .A(n56617), .B(n56616), .Z(n61613) );
  IV U76755 ( .A(n56618), .Z(n56620) );
  NOR U76756 ( .A(n56620), .B(n56619), .Z(n62289) );
  NOR U76757 ( .A(n61613), .B(n62289), .Z(n57271) );
  IV U76758 ( .A(n56621), .Z(n56623) );
  NOR U76759 ( .A(n56623), .B(n56622), .Z(n62284) );
  IV U76760 ( .A(n56624), .Z(n56625) );
  NOR U76761 ( .A(n56626), .B(n56625), .Z(n62286) );
  NOR U76762 ( .A(n62284), .B(n62286), .Z(n57270) );
  IV U76763 ( .A(n56627), .Z(n61618) );
  IV U76764 ( .A(n56628), .Z(n56632) );
  NOR U76765 ( .A(n56630), .B(n56629), .Z(n56631) );
  IV U76766 ( .A(n56631), .Z(n56634) );
  NOR U76767 ( .A(n56632), .B(n56634), .Z(n61615) );
  IV U76768 ( .A(n56633), .Z(n56635) );
  NOR U76769 ( .A(n56635), .B(n56634), .Z(n61620) );
  NOR U76770 ( .A(n61623), .B(n61620), .Z(n57267) );
  IV U76771 ( .A(n56636), .Z(n56638) );
  NOR U76772 ( .A(n56638), .B(n56637), .Z(n62272) );
  IV U76773 ( .A(n56639), .Z(n56643) );
  NOR U76774 ( .A(n56641), .B(n56640), .Z(n56642) );
  IV U76775 ( .A(n56642), .Z(n56648) );
  NOR U76776 ( .A(n56643), .B(n56648), .Z(n61626) );
  IV U76777 ( .A(n56644), .Z(n56646) );
  NOR U76778 ( .A(n56646), .B(n56645), .Z(n61634) );
  IV U76779 ( .A(n56647), .Z(n56649) );
  NOR U76780 ( .A(n56649), .B(n56648), .Z(n61632) );
  NOR U76781 ( .A(n61634), .B(n61632), .Z(n57259) );
  IV U76782 ( .A(n56650), .Z(n56652) );
  NOR U76783 ( .A(n56652), .B(n56651), .Z(n57255) );
  IV U76784 ( .A(n56653), .Z(n56655) );
  NOR U76785 ( .A(n56655), .B(n56654), .Z(n56656) );
  IV U76786 ( .A(n56656), .Z(n62247) );
  IV U76787 ( .A(n56657), .Z(n56658) );
  NOR U76788 ( .A(n56661), .B(n56658), .Z(n61652) );
  IV U76789 ( .A(n56659), .Z(n56660) );
  NOR U76790 ( .A(n56661), .B(n56660), .Z(n61649) );
  IV U76791 ( .A(n56662), .Z(n56669) );
  NOR U76792 ( .A(n56664), .B(n56663), .Z(n56665) );
  IV U76793 ( .A(n56665), .Z(n56666) );
  NOR U76794 ( .A(n56667), .B(n56666), .Z(n56668) );
  IV U76795 ( .A(n56668), .Z(n56671) );
  NOR U76796 ( .A(n56669), .B(n56671), .Z(n61655) );
  IV U76797 ( .A(n56670), .Z(n56672) );
  NOR U76798 ( .A(n56672), .B(n56671), .Z(n57219) );
  IV U76799 ( .A(n56673), .Z(n62235) );
  IV U76800 ( .A(n56674), .Z(n56676) );
  NOR U76801 ( .A(n56676), .B(n56675), .Z(n61666) );
  IV U76802 ( .A(n56677), .Z(n56678) );
  NOR U76803 ( .A(n56679), .B(n56678), .Z(n67187) );
  IV U76804 ( .A(n56680), .Z(n56683) );
  NOR U76805 ( .A(n56681), .B(n56691), .Z(n56682) );
  IV U76806 ( .A(n56682), .Z(n56685) );
  NOR U76807 ( .A(n56683), .B(n56685), .Z(n67667) );
  NOR U76808 ( .A(n67187), .B(n67667), .Z(n61673) );
  IV U76809 ( .A(n56684), .Z(n56686) );
  NOR U76810 ( .A(n56686), .B(n56685), .Z(n61670) );
  IV U76811 ( .A(n56687), .Z(n56689) );
  NOR U76812 ( .A(n56689), .B(n56688), .Z(n61677) );
  IV U76813 ( .A(n56690), .Z(n56692) );
  NOR U76814 ( .A(n56692), .B(n56691), .Z(n61675) );
  NOR U76815 ( .A(n61677), .B(n61675), .Z(n57203) );
  NOR U76816 ( .A(n56694), .B(n56693), .Z(n61680) );
  IV U76817 ( .A(n56695), .Z(n56696) );
  NOR U76818 ( .A(n56696), .B(n57193), .Z(n62224) );
  NOR U76819 ( .A(n61680), .B(n62224), .Z(n57202) );
  IV U76820 ( .A(n56697), .Z(n56699) );
  NOR U76821 ( .A(n56699), .B(n56698), .Z(n57177) );
  IV U76822 ( .A(n57177), .Z(n57170) );
  IV U76823 ( .A(n56700), .Z(n61692) );
  NOR U76824 ( .A(n61692), .B(n56701), .Z(n57174) );
  IV U76825 ( .A(n56702), .Z(n56703) );
  NOR U76826 ( .A(n56703), .B(n56707), .Z(n62200) );
  IV U76827 ( .A(n56704), .Z(n56706) );
  NOR U76828 ( .A(n56706), .B(n56705), .Z(n61696) );
  NOR U76829 ( .A(n56708), .B(n56707), .Z(n56709) );
  IV U76830 ( .A(n56709), .Z(n56710) );
  NOR U76831 ( .A(n56711), .B(n56710), .Z(n62197) );
  NOR U76832 ( .A(n61696), .B(n62197), .Z(n57168) );
  IV U76833 ( .A(n56712), .Z(n56713) );
  NOR U76834 ( .A(n56714), .B(n56713), .Z(n62187) );
  IV U76835 ( .A(n56715), .Z(n56717) );
  NOR U76836 ( .A(n56717), .B(n56716), .Z(n61698) );
  NOR U76837 ( .A(n62187), .B(n61698), .Z(n57167) );
  IV U76838 ( .A(n56718), .Z(n56719) );
  NOR U76839 ( .A(n56719), .B(n56722), .Z(n62184) );
  IV U76840 ( .A(n56720), .Z(n56721) );
  NOR U76841 ( .A(n56722), .B(n56721), .Z(n61700) );
  IV U76842 ( .A(n56723), .Z(n56725) );
  NOR U76843 ( .A(n56725), .B(n56724), .Z(n62193) );
  IV U76844 ( .A(n56726), .Z(n56727) );
  NOR U76845 ( .A(n56728), .B(n56727), .Z(n62191) );
  NOR U76846 ( .A(n62193), .B(n62191), .Z(n57166) );
  IV U76847 ( .A(n56729), .Z(n56730) );
  NOR U76848 ( .A(n56731), .B(n56730), .Z(n62180) );
  NOR U76849 ( .A(n62176), .B(n62180), .Z(n57165) );
  IV U76850 ( .A(n56732), .Z(n56733) );
  NOR U76851 ( .A(n57161), .B(n56733), .Z(n62173) );
  IV U76852 ( .A(n56734), .Z(n56736) );
  NOR U76853 ( .A(n56736), .B(n56735), .Z(n61709) );
  IV U76854 ( .A(n56737), .Z(n56744) );
  NOR U76855 ( .A(n56739), .B(n56738), .Z(n56740) );
  IV U76856 ( .A(n56740), .Z(n56741) );
  NOR U76857 ( .A(n56742), .B(n56741), .Z(n56743) );
  IV U76858 ( .A(n56743), .Z(n57155) );
  NOR U76859 ( .A(n56744), .B(n57155), .Z(n61712) );
  IV U76860 ( .A(n56745), .Z(n56748) );
  NOR U76861 ( .A(n57148), .B(n56754), .Z(n56746) );
  IV U76862 ( .A(n56746), .Z(n56747) );
  NOR U76863 ( .A(n56748), .B(n56747), .Z(n61715) );
  NOR U76864 ( .A(n56749), .B(n62153), .Z(n56756) );
  IV U76865 ( .A(n56750), .Z(n56752) );
  NOR U76866 ( .A(n56752), .B(n56751), .Z(n56753) );
  IV U76867 ( .A(n56753), .Z(n56755) );
  NOR U76868 ( .A(n56755), .B(n56754), .Z(n61719) );
  NOR U76869 ( .A(n56756), .B(n61719), .Z(n57145) );
  IV U76870 ( .A(n56757), .Z(n57138) );
  IV U76871 ( .A(n56758), .Z(n56759) );
  NOR U76872 ( .A(n57138), .B(n56759), .Z(n57143) );
  IV U76873 ( .A(n57143), .Z(n57136) );
  IV U76874 ( .A(n57139), .Z(n56760) );
  NOR U76875 ( .A(n57138), .B(n56760), .Z(n61724) );
  IV U76876 ( .A(n56761), .Z(n56762) );
  NOR U76877 ( .A(n57132), .B(n56762), .Z(n62142) );
  IV U76878 ( .A(n56763), .Z(n56764) );
  NOR U76879 ( .A(n56764), .B(n56771), .Z(n56765) );
  IV U76880 ( .A(n56765), .Z(n62134) );
  IV U76881 ( .A(n56766), .Z(n56767) );
  NOR U76882 ( .A(n56768), .B(n56767), .Z(n62128) );
  IV U76883 ( .A(n56769), .Z(n56770) );
  NOR U76884 ( .A(n56771), .B(n56770), .Z(n61733) );
  NOR U76885 ( .A(n62128), .B(n61733), .Z(n57124) );
  IV U76886 ( .A(n56772), .Z(n56773) );
  NOR U76887 ( .A(n56774), .B(n56773), .Z(n56775) );
  IV U76888 ( .A(n56775), .Z(n57115) );
  IV U76889 ( .A(n56776), .Z(n56777) );
  NOR U76890 ( .A(n57105), .B(n56777), .Z(n61735) );
  IV U76891 ( .A(n61735), .Z(n67252) );
  IV U76892 ( .A(n56778), .Z(n56780) );
  IV U76893 ( .A(n56779), .Z(n57107) );
  NOR U76894 ( .A(n56780), .B(n57107), .Z(n67265) );
  NOR U76895 ( .A(n67270), .B(n67265), .Z(n61745) );
  NOR U76896 ( .A(n56782), .B(n56781), .Z(n56783) );
  IV U76897 ( .A(n56783), .Z(n61751) );
  IV U76898 ( .A(n56784), .Z(n56785) );
  NOR U76899 ( .A(n56785), .B(n56791), .Z(n56786) );
  IV U76900 ( .A(n56786), .Z(n62112) );
  IV U76901 ( .A(n56787), .Z(n56788) );
  NOR U76902 ( .A(n56789), .B(n56788), .Z(n61760) );
  IV U76903 ( .A(n56790), .Z(n56792) );
  NOR U76904 ( .A(n56792), .B(n56791), .Z(n62108) );
  NOR U76905 ( .A(n61760), .B(n62108), .Z(n57094) );
  IV U76906 ( .A(n56793), .Z(n56794) );
  NOR U76907 ( .A(n56795), .B(n56794), .Z(n67291) );
  IV U76908 ( .A(n61767), .Z(n56796) );
  NOR U76909 ( .A(n56796), .B(n61766), .Z(n67286) );
  NOR U76910 ( .A(n67291), .B(n67286), .Z(n61771) );
  IV U76911 ( .A(n56797), .Z(n56799) );
  NOR U76912 ( .A(n56799), .B(n56798), .Z(n61772) );
  IV U76913 ( .A(n56800), .Z(n56801) );
  NOR U76914 ( .A(n56802), .B(n56801), .Z(n61780) );
  IV U76915 ( .A(n56803), .Z(n56804) );
  NOR U76916 ( .A(n56805), .B(n56804), .Z(n61775) );
  NOR U76917 ( .A(n61780), .B(n61775), .Z(n57084) );
  IV U76918 ( .A(n56806), .Z(n67306) );
  NOR U76919 ( .A(n67306), .B(n67309), .Z(n61783) );
  IV U76920 ( .A(n56807), .Z(n56808) );
  NOR U76921 ( .A(n56809), .B(n56808), .Z(n61777) );
  NOR U76922 ( .A(n61783), .B(n61777), .Z(n57083) );
  IV U76923 ( .A(n56810), .Z(n56811) );
  NOR U76924 ( .A(n56812), .B(n56811), .Z(n62086) );
  IV U76925 ( .A(n67310), .Z(n56813) );
  NOR U76926 ( .A(n56813), .B(n67309), .Z(n62079) );
  NOR U76927 ( .A(n62086), .B(n62079), .Z(n61785) );
  IV U76928 ( .A(n56814), .Z(n56820) );
  XOR U76929 ( .A(n56820), .B(n56819), .Z(n56817) );
  IV U76930 ( .A(n56815), .Z(n56816) );
  NOR U76931 ( .A(n56817), .B(n56816), .Z(n56818) );
  IV U76932 ( .A(n56818), .Z(n62075) );
  IV U76933 ( .A(n56819), .Z(n56821) );
  NOR U76934 ( .A(n56821), .B(n56820), .Z(n67318) );
  IV U76935 ( .A(n56822), .Z(n56823) );
  NOR U76936 ( .A(n56823), .B(n57080), .Z(n67323) );
  NOR U76937 ( .A(n67318), .B(n67323), .Z(n62072) );
  NOR U76938 ( .A(n61796), .B(n61790), .Z(n57074) );
  IV U76939 ( .A(n56824), .Z(n56826) );
  NOR U76940 ( .A(n56826), .B(n56825), .Z(n62041) );
  IV U76941 ( .A(n56827), .Z(n61801) );
  NOR U76942 ( .A(n56828), .B(n61801), .Z(n56829) );
  NOR U76943 ( .A(n62031), .B(n56829), .Z(n57060) );
  IV U76944 ( .A(n56830), .Z(n56831) );
  NOR U76945 ( .A(n56831), .B(n57058), .Z(n62018) );
  IV U76946 ( .A(n56832), .Z(n56833) );
  NOR U76947 ( .A(n56834), .B(n56833), .Z(n56835) );
  IV U76948 ( .A(n56835), .Z(n61807) );
  IV U76949 ( .A(n56836), .Z(n56837) );
  NOR U76950 ( .A(n56837), .B(n56839), .Z(n61810) );
  IV U76951 ( .A(n56838), .Z(n56840) );
  NOR U76952 ( .A(n56840), .B(n56839), .Z(n61808) );
  NOR U76953 ( .A(n61810), .B(n61808), .Z(n57052) );
  IV U76954 ( .A(n56841), .Z(n56843) );
  IV U76955 ( .A(n56842), .Z(n57050) );
  NOR U76956 ( .A(n56843), .B(n57050), .Z(n61816) );
  NOR U76957 ( .A(n56844), .B(n61838), .Z(n61827) );
  IV U76958 ( .A(n56845), .Z(n61833) );
  NOR U76959 ( .A(n56846), .B(n61833), .Z(n56847) );
  NOR U76960 ( .A(n61827), .B(n56847), .Z(n57013) );
  IV U76961 ( .A(n56848), .Z(n56849) );
  NOR U76962 ( .A(n56850), .B(n56849), .Z(n61850) );
  IV U76963 ( .A(n56851), .Z(n56852) );
  NOR U76964 ( .A(n56853), .B(n56852), .Z(n61845) );
  NOR U76965 ( .A(n61850), .B(n61845), .Z(n57012) );
  IV U76966 ( .A(n56854), .Z(n56855) );
  NOR U76967 ( .A(n56856), .B(n56855), .Z(n61847) );
  IV U76968 ( .A(n56857), .Z(n56858) );
  NOR U76969 ( .A(n56861), .B(n56858), .Z(n61969) );
  IV U76970 ( .A(n56859), .Z(n56860) );
  NOR U76971 ( .A(n56861), .B(n56860), .Z(n61966) );
  IV U76972 ( .A(n56862), .Z(n56863) );
  NOR U76973 ( .A(n56864), .B(n56863), .Z(n61856) );
  IV U76974 ( .A(n56865), .Z(n56867) );
  IV U76975 ( .A(n56866), .Z(n57010) );
  NOR U76976 ( .A(n56867), .B(n57010), .Z(n61853) );
  NOR U76977 ( .A(n56869), .B(n56868), .Z(n61862) );
  IV U76978 ( .A(n56870), .Z(n56871) );
  NOR U76979 ( .A(n56874), .B(n56871), .Z(n61870) );
  IV U76980 ( .A(n56872), .Z(n56873) );
  NOR U76981 ( .A(n56874), .B(n56873), .Z(n61868) );
  XOR U76982 ( .A(n61870), .B(n61868), .Z(n56875) );
  NOR U76983 ( .A(n61862), .B(n56875), .Z(n57007) );
  IV U76984 ( .A(n56876), .Z(n56877) );
  NOR U76985 ( .A(n56877), .B(n57005), .Z(n56878) );
  IV U76986 ( .A(n56878), .Z(n61874) );
  IV U76987 ( .A(n56879), .Z(n56883) );
  NOR U76988 ( .A(n56881), .B(n56880), .Z(n56882) );
  IV U76989 ( .A(n56882), .Z(n56889) );
  NOR U76990 ( .A(n56883), .B(n56889), .Z(n56884) );
  IV U76991 ( .A(n56884), .Z(n61957) );
  IV U76992 ( .A(n56885), .Z(n56886) );
  NOR U76993 ( .A(n56887), .B(n56886), .Z(n61883) );
  IV U76994 ( .A(n56888), .Z(n56890) );
  NOR U76995 ( .A(n56890), .B(n56889), .Z(n61878) );
  NOR U76996 ( .A(n61883), .B(n61878), .Z(n56999) );
  IV U76997 ( .A(n56891), .Z(n56892) );
  NOR U76998 ( .A(n56893), .B(n56892), .Z(n61880) );
  IV U76999 ( .A(n56894), .Z(n56895) );
  NOR U77000 ( .A(n56995), .B(n56895), .Z(n56896) );
  IV U77001 ( .A(n56896), .Z(n61953) );
  IV U77002 ( .A(n56897), .Z(n56899) );
  IV U77003 ( .A(n56898), .Z(n56997) );
  NOR U77004 ( .A(n56899), .B(n56997), .Z(n61886) );
  IV U77005 ( .A(n56900), .Z(n56902) );
  NOR U77006 ( .A(n56902), .B(n56901), .Z(n61943) );
  NOR U77007 ( .A(n56903), .B(n61891), .Z(n56904) );
  NOR U77008 ( .A(n61943), .B(n56904), .Z(n56992) );
  IV U77009 ( .A(n56905), .Z(n56907) );
  NOR U77010 ( .A(n56907), .B(n56906), .Z(n61894) );
  IV U77011 ( .A(n56908), .Z(n56909) );
  NOR U77012 ( .A(n56909), .B(n56911), .Z(n61897) );
  IV U77013 ( .A(n56910), .Z(n56912) );
  NOR U77014 ( .A(n56912), .B(n56911), .Z(n61899) );
  IV U77015 ( .A(n56913), .Z(n56914) );
  NOR U77016 ( .A(n56915), .B(n56914), .Z(n61905) );
  NOR U77017 ( .A(n61899), .B(n61905), .Z(n56916) );
  IV U77018 ( .A(n56916), .Z(n56917) );
  NOR U77019 ( .A(n61897), .B(n56917), .Z(n56918) );
  IV U77020 ( .A(n56918), .Z(n56985) );
  IV U77021 ( .A(n56919), .Z(n56921) );
  NOR U77022 ( .A(n56921), .B(n56920), .Z(n61902) );
  IV U77023 ( .A(n56924), .Z(n56922) );
  NOR U77024 ( .A(n56923), .B(n56922), .Z(n61939) );
  NOR U77025 ( .A(n56925), .B(n56924), .Z(n56928) );
  IV U77026 ( .A(n56926), .Z(n56927) );
  NOR U77027 ( .A(n56928), .B(n56927), .Z(n56929) );
  NOR U77028 ( .A(n61939), .B(n56929), .Z(n61935) );
  IV U77029 ( .A(n56930), .Z(n56931) );
  NOR U77030 ( .A(n56932), .B(n56931), .Z(n61908) );
  NOR U77031 ( .A(n56934), .B(n56933), .Z(n61928) );
  NOR U77032 ( .A(n61908), .B(n61928), .Z(n56984) );
  IV U77033 ( .A(n56935), .Z(n56936) );
  NOR U77034 ( .A(n56938), .B(n56936), .Z(n61913) );
  IV U77035 ( .A(n56937), .Z(n56939) );
  NOR U77036 ( .A(n56939), .B(n56938), .Z(n56940) );
  IV U77037 ( .A(n56940), .Z(n61911) );
  IV U77038 ( .A(n56941), .Z(n56942) );
  NOR U77039 ( .A(n56943), .B(n56942), .Z(n61920) );
  NOR U77040 ( .A(n56945), .B(n56944), .Z(n56968) );
  NOR U77041 ( .A(n56971), .B(n56968), .Z(n56961) );
  IV U77042 ( .A(n56946), .Z(n56948) );
  NOR U77043 ( .A(n56957), .B(n56948), .Z(n56955) );
  IV U77044 ( .A(n56947), .Z(n56953) );
  IV U77045 ( .A(n56949), .Z(n56956) );
  XOR U77046 ( .A(n56957), .B(n56956), .Z(n56951) );
  NOR U77047 ( .A(n56949), .B(n56948), .Z(n56950) );
  NOR U77048 ( .A(n56951), .B(n56950), .Z(n56952) );
  NOR U77049 ( .A(n56953), .B(n56952), .Z(n56954) );
  NOR U77050 ( .A(n56955), .B(n56954), .Z(n56967) );
  IV U77051 ( .A(n56967), .Z(n56958) );
  NOR U77052 ( .A(n56957), .B(n56956), .Z(n56964) );
  NOR U77053 ( .A(n56958), .B(n56964), .Z(n56959) );
  IV U77054 ( .A(n56959), .Z(n56960) );
  NOR U77055 ( .A(n56961), .B(n56960), .Z(n56973) );
  NOR U77056 ( .A(n56963), .B(n56962), .Z(n56966) );
  IV U77057 ( .A(n56964), .Z(n56965) );
  NOR U77058 ( .A(n56966), .B(n56965), .Z(n56970) );
  NOR U77059 ( .A(n56968), .B(n56967), .Z(n56969) );
  NOR U77060 ( .A(n56970), .B(n56969), .Z(n56972) );
  NOR U77061 ( .A(n56972), .B(n56971), .Z(n67454) );
  NOR U77062 ( .A(n56973), .B(n67454), .Z(n56974) );
  IV U77063 ( .A(n56974), .Z(n61921) );
  XOR U77064 ( .A(n61920), .B(n61921), .Z(n61918) );
  IV U77065 ( .A(n56977), .Z(n56976) );
  NOR U77066 ( .A(n56976), .B(n56975), .Z(n56983) );
  NOR U77067 ( .A(n56978), .B(n56977), .Z(n56981) );
  IV U77068 ( .A(n56979), .Z(n56980) );
  NOR U77069 ( .A(n56981), .B(n56980), .Z(n56982) );
  NOR U77070 ( .A(n56983), .B(n56982), .Z(n61919) );
  XOR U77071 ( .A(n61918), .B(n61919), .Z(n61910) );
  XOR U77072 ( .A(n61911), .B(n61910), .Z(n61914) );
  XOR U77073 ( .A(n61913), .B(n61914), .Z(n61929) );
  XOR U77074 ( .A(n56984), .B(n61929), .Z(n61931) );
  XOR U77075 ( .A(n61935), .B(n61931), .Z(n61903) );
  XOR U77076 ( .A(n61902), .B(n61903), .Z(n61906) );
  XOR U77077 ( .A(n56985), .B(n61906), .Z(n67440) );
  XOR U77078 ( .A(n61894), .B(n67440), .Z(n61941) );
  IV U77079 ( .A(n56986), .Z(n56988) );
  NOR U77080 ( .A(n56988), .B(n56987), .Z(n67438) );
  IV U77081 ( .A(n56989), .Z(n67437) );
  NOR U77082 ( .A(n56990), .B(n67437), .Z(n56991) );
  NOR U77083 ( .A(n67438), .B(n56991), .Z(n61942) );
  XOR U77084 ( .A(n61941), .B(n61942), .Z(n61890) );
  XOR U77085 ( .A(n56992), .B(n61890), .Z(n61888) );
  XOR U77086 ( .A(n61886), .B(n61888), .Z(n67424) );
  IV U77087 ( .A(n56993), .Z(n56994) );
  NOR U77088 ( .A(n56995), .B(n56994), .Z(n67422) );
  IV U77089 ( .A(n56996), .Z(n56998) );
  NOR U77090 ( .A(n56998), .B(n56997), .Z(n67428) );
  NOR U77091 ( .A(n67422), .B(n67428), .Z(n61950) );
  XOR U77092 ( .A(n67424), .B(n61950), .Z(n61951) );
  XOR U77093 ( .A(n61953), .B(n61951), .Z(n61881) );
  XOR U77094 ( .A(n61880), .B(n61881), .Z(n61884) );
  XOR U77095 ( .A(n56999), .B(n61884), .Z(n61956) );
  XOR U77096 ( .A(n61957), .B(n61956), .Z(n61960) );
  IV U77097 ( .A(n57000), .Z(n57002) );
  NOR U77098 ( .A(n57002), .B(n57001), .Z(n61959) );
  IV U77099 ( .A(n57003), .Z(n57004) );
  NOR U77100 ( .A(n57005), .B(n57004), .Z(n61876) );
  NOR U77101 ( .A(n61959), .B(n61876), .Z(n57006) );
  XOR U77102 ( .A(n61960), .B(n57006), .Z(n61873) );
  XOR U77103 ( .A(n61874), .B(n61873), .Z(n61869) );
  XOR U77104 ( .A(n57007), .B(n61869), .Z(n61860) );
  IV U77105 ( .A(n57008), .Z(n57009) );
  NOR U77106 ( .A(n57010), .B(n57009), .Z(n61859) );
  NOR U77107 ( .A(n61864), .B(n61859), .Z(n57011) );
  XOR U77108 ( .A(n61860), .B(n57011), .Z(n61854) );
  XOR U77109 ( .A(n61853), .B(n61854), .Z(n61857) );
  XOR U77110 ( .A(n61856), .B(n61857), .Z(n61967) );
  XOR U77111 ( .A(n61966), .B(n61967), .Z(n61970) );
  XOR U77112 ( .A(n61969), .B(n61970), .Z(n61849) );
  XOR U77113 ( .A(n61847), .B(n61849), .Z(n61851) );
  XOR U77114 ( .A(n57012), .B(n61851), .Z(n61826) );
  XOR U77115 ( .A(n57013), .B(n61826), .Z(n61987) );
  NOR U77116 ( .A(n57014), .B(n61828), .Z(n57018) );
  IV U77117 ( .A(n57015), .Z(n57017) );
  NOR U77118 ( .A(n57017), .B(n57016), .Z(n61985) );
  NOR U77119 ( .A(n57018), .B(n61985), .Z(n57019) );
  XOR U77120 ( .A(n61987), .B(n57019), .Z(n61983) );
  IV U77121 ( .A(n57022), .Z(n57020) );
  NOR U77122 ( .A(n57020), .B(n57021), .Z(n61982) );
  XOR U77123 ( .A(n57022), .B(n57021), .Z(n57023) );
  NOR U77124 ( .A(n57024), .B(n57023), .Z(n57025) );
  IV U77125 ( .A(n57025), .Z(n57026) );
  NOR U77126 ( .A(n57027), .B(n57026), .Z(n61991) );
  NOR U77127 ( .A(n61982), .B(n61991), .Z(n57028) );
  XOR U77128 ( .A(n61983), .B(n57028), .Z(n61997) );
  IV U77129 ( .A(n57029), .Z(n57031) );
  NOR U77130 ( .A(n57031), .B(n57030), .Z(n61989) );
  IV U77131 ( .A(n57032), .Z(n57034) );
  NOR U77132 ( .A(n57034), .B(n57033), .Z(n61995) );
  NOR U77133 ( .A(n61989), .B(n61995), .Z(n57035) );
  XOR U77134 ( .A(n61997), .B(n57035), .Z(n61823) );
  IV U77135 ( .A(n57036), .Z(n57038) );
  NOR U77136 ( .A(n57038), .B(n57037), .Z(n62001) );
  IV U77137 ( .A(n57039), .Z(n57041) );
  NOR U77138 ( .A(n57041), .B(n57040), .Z(n61822) );
  NOR U77139 ( .A(n62001), .B(n61822), .Z(n57042) );
  XOR U77140 ( .A(n61823), .B(n57042), .Z(n62000) );
  IV U77141 ( .A(n57043), .Z(n57044) );
  NOR U77142 ( .A(n57044), .B(n57046), .Z(n61820) );
  IV U77143 ( .A(n57045), .Z(n57047) );
  NOR U77144 ( .A(n57047), .B(n57046), .Z(n61998) );
  NOR U77145 ( .A(n61820), .B(n61998), .Z(n57048) );
  XOR U77146 ( .A(n62000), .B(n57048), .Z(n61814) );
  IV U77147 ( .A(n57049), .Z(n57051) );
  NOR U77148 ( .A(n57051), .B(n57050), .Z(n67352) );
  NOR U77149 ( .A(n67357), .B(n67352), .Z(n61815) );
  XOR U77150 ( .A(n61814), .B(n61815), .Z(n61817) );
  XOR U77151 ( .A(n61816), .B(n61817), .Z(n61811) );
  XOR U77152 ( .A(n57052), .B(n61811), .Z(n61805) );
  XOR U77153 ( .A(n61807), .B(n61805), .Z(n67343) );
  IV U77154 ( .A(n67343), .Z(n57059) );
  IV U77155 ( .A(n57053), .Z(n57055) );
  NOR U77156 ( .A(n57055), .B(n57054), .Z(n62012) );
  IV U77157 ( .A(n57056), .Z(n57057) );
  NOR U77158 ( .A(n57058), .B(n57057), .Z(n62009) );
  NOR U77159 ( .A(n62012), .B(n62009), .Z(n61804) );
  XOR U77160 ( .A(n57059), .B(n61804), .Z(n62019) );
  XOR U77161 ( .A(n62018), .B(n62019), .Z(n62032) );
  XOR U77162 ( .A(n57060), .B(n62032), .Z(n57061) );
  IV U77163 ( .A(n57061), .Z(n62043) );
  XOR U77164 ( .A(n62041), .B(n62043), .Z(n62046) );
  IV U77165 ( .A(n57062), .Z(n57066) );
  NOR U77166 ( .A(n57064), .B(n57063), .Z(n57065) );
  IV U77167 ( .A(n57065), .Z(n57071) );
  NOR U77168 ( .A(n57066), .B(n57071), .Z(n62044) );
  XOR U77169 ( .A(n62046), .B(n62044), .Z(n62056) );
  IV U77170 ( .A(n57067), .Z(n57069) );
  NOR U77171 ( .A(n57069), .B(n57068), .Z(n62050) );
  IV U77172 ( .A(n57070), .Z(n57072) );
  NOR U77173 ( .A(n57072), .B(n57071), .Z(n62052) );
  NOR U77174 ( .A(n62050), .B(n62052), .Z(n57073) );
  XOR U77175 ( .A(n62056), .B(n57073), .Z(n61791) );
  XOR U77176 ( .A(n57074), .B(n61791), .Z(n61794) );
  IV U77177 ( .A(n57075), .Z(n61787) );
  NOR U77178 ( .A(n57076), .B(n61787), .Z(n57077) );
  NOR U77179 ( .A(n61793), .B(n57077), .Z(n57078) );
  XOR U77180 ( .A(n61794), .B(n57078), .Z(n62065) );
  IV U77181 ( .A(n57079), .Z(n57081) );
  NOR U77182 ( .A(n57081), .B(n57080), .Z(n57082) );
  IV U77183 ( .A(n57082), .Z(n62066) );
  XOR U77184 ( .A(n62065), .B(n62066), .Z(n67319) );
  XOR U77185 ( .A(n62072), .B(n67319), .Z(n62073) );
  XOR U77186 ( .A(n62075), .B(n62073), .Z(n62082) );
  XOR U77187 ( .A(n61785), .B(n62082), .Z(n61778) );
  XOR U77188 ( .A(n57083), .B(n61778), .Z(n61782) );
  XOR U77189 ( .A(n57084), .B(n61782), .Z(n57085) );
  IV U77190 ( .A(n57085), .Z(n61773) );
  XOR U77191 ( .A(n61772), .B(n61773), .Z(n67288) );
  XOR U77192 ( .A(n61771), .B(n67288), .Z(n61762) );
  IV U77193 ( .A(n57086), .Z(n61769) );
  NOR U77194 ( .A(n61769), .B(n61766), .Z(n62101) );
  IV U77195 ( .A(n57087), .Z(n57089) );
  IV U77196 ( .A(n57088), .Z(n57092) );
  NOR U77197 ( .A(n57089), .B(n57092), .Z(n61763) );
  NOR U77198 ( .A(n62101), .B(n61763), .Z(n57090) );
  XOR U77199 ( .A(n61762), .B(n57090), .Z(n61759) );
  IV U77200 ( .A(n57091), .Z(n57093) );
  NOR U77201 ( .A(n57093), .B(n57092), .Z(n61757) );
  XOR U77202 ( .A(n61759), .B(n61757), .Z(n62109) );
  XOR U77203 ( .A(n57094), .B(n62109), .Z(n62111) );
  XOR U77204 ( .A(n62112), .B(n62111), .Z(n62115) );
  IV U77205 ( .A(n57095), .Z(n57097) );
  NOR U77206 ( .A(n57097), .B(n57096), .Z(n62114) );
  IV U77207 ( .A(n57098), .Z(n57099) );
  NOR U77208 ( .A(n57100), .B(n57099), .Z(n61755) );
  NOR U77209 ( .A(n62114), .B(n61755), .Z(n57101) );
  XOR U77210 ( .A(n62115), .B(n57101), .Z(n61750) );
  XOR U77211 ( .A(n61751), .B(n61750), .Z(n61753) );
  XOR U77212 ( .A(n57102), .B(n61753), .Z(n67266) );
  XOR U77213 ( .A(n61745), .B(n67266), .Z(n61746) );
  IV U77214 ( .A(n57103), .Z(n57104) );
  NOR U77215 ( .A(n57105), .B(n57104), .Z(n67256) );
  IV U77216 ( .A(n57106), .Z(n57108) );
  NOR U77217 ( .A(n57108), .B(n57107), .Z(n61747) );
  NOR U77218 ( .A(n67256), .B(n61747), .Z(n57109) );
  XOR U77219 ( .A(n61746), .B(n57109), .Z(n67253) );
  XOR U77220 ( .A(n67252), .B(n67253), .Z(n61736) );
  IV U77221 ( .A(n61736), .Z(n61739) );
  NOR U77222 ( .A(n57115), .B(n61739), .Z(n67245) );
  IV U77223 ( .A(n57110), .Z(n57111) );
  NOR U77224 ( .A(n57122), .B(n57111), .Z(n62122) );
  IV U77225 ( .A(n57112), .Z(n57114) );
  NOR U77226 ( .A(n57114), .B(n57113), .Z(n61738) );
  XOR U77227 ( .A(n61738), .B(n61739), .Z(n62123) );
  IV U77228 ( .A(n62123), .Z(n57116) );
  XOR U77229 ( .A(n62122), .B(n57116), .Z(n57118) );
  NOR U77230 ( .A(n57116), .B(n57115), .Z(n57117) );
  NOR U77231 ( .A(n57118), .B(n57117), .Z(n57119) );
  NOR U77232 ( .A(n67245), .B(n57119), .Z(n57120) );
  IV U77233 ( .A(n57120), .Z(n62126) );
  IV U77234 ( .A(n57121), .Z(n57123) );
  NOR U77235 ( .A(n57123), .B(n57122), .Z(n62125) );
  XOR U77236 ( .A(n62126), .B(n62125), .Z(n62129) );
  XOR U77237 ( .A(n57124), .B(n62129), .Z(n62133) );
  XOR U77238 ( .A(n62134), .B(n62133), .Z(n62138) );
  IV U77239 ( .A(n57125), .Z(n57127) );
  NOR U77240 ( .A(n57127), .B(n57126), .Z(n62136) );
  XOR U77241 ( .A(n62138), .B(n62136), .Z(n61730) );
  IV U77242 ( .A(n57128), .Z(n57129) );
  NOR U77243 ( .A(n57132), .B(n57129), .Z(n61729) );
  IV U77244 ( .A(n57130), .Z(n57131) );
  NOR U77245 ( .A(n57132), .B(n57131), .Z(n61727) );
  NOR U77246 ( .A(n61729), .B(n61727), .Z(n57133) );
  XOR U77247 ( .A(n61730), .B(n57133), .Z(n57134) );
  IV U77248 ( .A(n57134), .Z(n62144) );
  XOR U77249 ( .A(n62142), .B(n62144), .Z(n61725) );
  XOR U77250 ( .A(n61724), .B(n61725), .Z(n57135) );
  NOR U77251 ( .A(n57136), .B(n57135), .Z(n67601) );
  IV U77252 ( .A(n57137), .Z(n57141) );
  XOR U77253 ( .A(n57139), .B(n57138), .Z(n57140) );
  NOR U77254 ( .A(n57141), .B(n57140), .Z(n61722) );
  NOR U77255 ( .A(n61724), .B(n61722), .Z(n57142) );
  XOR U77256 ( .A(n57142), .B(n61725), .Z(n62151) );
  NOR U77257 ( .A(n57143), .B(n62151), .Z(n57144) );
  NOR U77258 ( .A(n67601), .B(n57144), .Z(n61718) );
  XOR U77259 ( .A(n57145), .B(n61718), .Z(n61717) );
  XOR U77260 ( .A(n61715), .B(n61717), .Z(n62163) );
  IV U77261 ( .A(n57146), .Z(n57150) );
  NOR U77262 ( .A(n57148), .B(n57147), .Z(n57149) );
  IV U77263 ( .A(n57149), .Z(n57152) );
  NOR U77264 ( .A(n57150), .B(n57152), .Z(n62161) );
  XOR U77265 ( .A(n62163), .B(n62161), .Z(n62166) );
  IV U77266 ( .A(n57151), .Z(n57153) );
  NOR U77267 ( .A(n57153), .B(n57152), .Z(n62164) );
  XOR U77268 ( .A(n62166), .B(n62164), .Z(n61713) );
  XOR U77269 ( .A(n61712), .B(n61713), .Z(n61708) );
  IV U77270 ( .A(n57154), .Z(n57156) );
  NOR U77271 ( .A(n57156), .B(n57155), .Z(n61706) );
  XOR U77272 ( .A(n61708), .B(n61706), .Z(n61710) );
  XOR U77273 ( .A(n61709), .B(n61710), .Z(n62171) );
  IV U77274 ( .A(n62171), .Z(n57164) );
  IV U77275 ( .A(n57157), .Z(n57158) );
  NOR U77276 ( .A(n57159), .B(n57158), .Z(n61704) );
  IV U77277 ( .A(n57160), .Z(n57162) );
  NOR U77278 ( .A(n57162), .B(n57161), .Z(n62170) );
  NOR U77279 ( .A(n61704), .B(n62170), .Z(n57163) );
  XOR U77280 ( .A(n57164), .B(n57163), .Z(n62175) );
  XOR U77281 ( .A(n62173), .B(n62175), .Z(n62181) );
  XOR U77282 ( .A(n57165), .B(n62181), .Z(n62190) );
  XOR U77283 ( .A(n57166), .B(n62190), .Z(n61701) );
  XOR U77284 ( .A(n61700), .B(n61701), .Z(n62185) );
  XOR U77285 ( .A(n62184), .B(n62185), .Z(n62188) );
  XOR U77286 ( .A(n57167), .B(n62188), .Z(n61695) );
  XOR U77287 ( .A(n57168), .B(n61695), .Z(n62202) );
  XOR U77288 ( .A(n62200), .B(n62202), .Z(n61689) );
  XOR U77289 ( .A(n57174), .B(n61689), .Z(n57169) );
  NOR U77290 ( .A(n57170), .B(n57169), .Z(n67638) );
  IV U77291 ( .A(n57171), .Z(n57173) );
  NOR U77292 ( .A(n57173), .B(n57172), .Z(n61688) );
  NOR U77293 ( .A(n57174), .B(n61688), .Z(n57175) );
  XOR U77294 ( .A(n61689), .B(n57175), .Z(n57176) );
  NOR U77295 ( .A(n57177), .B(n57176), .Z(n57178) );
  NOR U77296 ( .A(n67638), .B(n57178), .Z(n61684) );
  NOR U77297 ( .A(n57179), .B(n57188), .Z(n57180) );
  IV U77298 ( .A(n57180), .Z(n57181) );
  NOR U77299 ( .A(n57182), .B(n57181), .Z(n57183) );
  IV U77300 ( .A(n57183), .Z(n61685) );
  XOR U77301 ( .A(n61684), .B(n61685), .Z(n62219) );
  IV U77302 ( .A(n57184), .Z(n57198) );
  IV U77303 ( .A(n57185), .Z(n57186) );
  NOR U77304 ( .A(n57198), .B(n57186), .Z(n62217) );
  IV U77305 ( .A(n57187), .Z(n57189) );
  NOR U77306 ( .A(n57189), .B(n57188), .Z(n62207) );
  NOR U77307 ( .A(n62217), .B(n62207), .Z(n57190) );
  XOR U77308 ( .A(n62219), .B(n57190), .Z(n57191) );
  IV U77309 ( .A(n57191), .Z(n62216) );
  IV U77310 ( .A(n57192), .Z(n57194) );
  NOR U77311 ( .A(n57194), .B(n57193), .Z(n57200) );
  IV U77312 ( .A(n57200), .Z(n57195) );
  NOR U77313 ( .A(n62216), .B(n57195), .Z(n62222) );
  IV U77314 ( .A(n57196), .Z(n57197) );
  NOR U77315 ( .A(n57198), .B(n57197), .Z(n62214) );
  XOR U77316 ( .A(n62214), .B(n62216), .Z(n62226) );
  IV U77317 ( .A(n62226), .Z(n57199) );
  NOR U77318 ( .A(n57200), .B(n57199), .Z(n57201) );
  NOR U77319 ( .A(n62222), .B(n57201), .Z(n61681) );
  XOR U77320 ( .A(n57202), .B(n61681), .Z(n61679) );
  XOR U77321 ( .A(n57203), .B(n61679), .Z(n57204) );
  IV U77322 ( .A(n57204), .Z(n61671) );
  XOR U77323 ( .A(n61670), .B(n61671), .Z(n67189) );
  XOR U77324 ( .A(n61673), .B(n67189), .Z(n57205) );
  IV U77325 ( .A(n57205), .Z(n61664) );
  XOR U77326 ( .A(n61663), .B(n61664), .Z(n61667) );
  XOR U77327 ( .A(n61666), .B(n61667), .Z(n62232) );
  IV U77328 ( .A(n57206), .Z(n57209) );
  IV U77329 ( .A(n57207), .Z(n57208) );
  NOR U77330 ( .A(n57209), .B(n57208), .Z(n61661) );
  NOR U77331 ( .A(n61661), .B(n62231), .Z(n57210) );
  XOR U77332 ( .A(n62232), .B(n57210), .Z(n62234) );
  XOR U77333 ( .A(n62235), .B(n62234), .Z(n62238) );
  IV U77334 ( .A(n57211), .Z(n57212) );
  NOR U77335 ( .A(n57213), .B(n57212), .Z(n62237) );
  IV U77336 ( .A(n57214), .Z(n57216) );
  NOR U77337 ( .A(n57216), .B(n57215), .Z(n61658) );
  NOR U77338 ( .A(n62237), .B(n61658), .Z(n57217) );
  XOR U77339 ( .A(n62238), .B(n57217), .Z(n57218) );
  NOR U77340 ( .A(n57219), .B(n57218), .Z(n57222) );
  IV U77341 ( .A(n57219), .Z(n57221) );
  XOR U77342 ( .A(n62237), .B(n62238), .Z(n57220) );
  NOR U77343 ( .A(n57221), .B(n57220), .Z(n67672) );
  NOR U77344 ( .A(n57222), .B(n67672), .Z(n57223) );
  IV U77345 ( .A(n57223), .Z(n61656) );
  XOR U77346 ( .A(n61655), .B(n61656), .Z(n61650) );
  XOR U77347 ( .A(n61649), .B(n61650), .Z(n61653) );
  XOR U77348 ( .A(n61652), .B(n61653), .Z(n61646) );
  IV U77349 ( .A(n57224), .Z(n57226) );
  NOR U77350 ( .A(n57226), .B(n57225), .Z(n61645) );
  IV U77351 ( .A(n57227), .Z(n57228) );
  NOR U77352 ( .A(n57229), .B(n57228), .Z(n61643) );
  NOR U77353 ( .A(n61645), .B(n61643), .Z(n57230) );
  XOR U77354 ( .A(n61646), .B(n57230), .Z(n61637) );
  IV U77355 ( .A(n57231), .Z(n57233) );
  NOR U77356 ( .A(n57233), .B(n57232), .Z(n61640) );
  IV U77357 ( .A(n57234), .Z(n57235) );
  NOR U77358 ( .A(n57235), .B(n57238), .Z(n61638) );
  NOR U77359 ( .A(n61640), .B(n61638), .Z(n57236) );
  XOR U77360 ( .A(n61637), .B(n57236), .Z(n62245) );
  IV U77361 ( .A(n57237), .Z(n57239) );
  NOR U77362 ( .A(n57239), .B(n57238), .Z(n62243) );
  XOR U77363 ( .A(n62245), .B(n62243), .Z(n62246) );
  XOR U77364 ( .A(n62247), .B(n62246), .Z(n62257) );
  IV U77365 ( .A(n57240), .Z(n57241) );
  NOR U77366 ( .A(n57242), .B(n57241), .Z(n62256) );
  IV U77367 ( .A(n57243), .Z(n57245) );
  NOR U77368 ( .A(n57245), .B(n57244), .Z(n62261) );
  NOR U77369 ( .A(n62256), .B(n62261), .Z(n57246) );
  XOR U77370 ( .A(n62257), .B(n57246), .Z(n62254) );
  IV U77371 ( .A(n57247), .Z(n57248) );
  NOR U77372 ( .A(n57249), .B(n57248), .Z(n62249) );
  IV U77373 ( .A(n57250), .Z(n57252) );
  NOR U77374 ( .A(n57252), .B(n57251), .Z(n62252) );
  NOR U77375 ( .A(n62249), .B(n62252), .Z(n57253) );
  XOR U77376 ( .A(n62254), .B(n57253), .Z(n57254) );
  NOR U77377 ( .A(n57255), .B(n57254), .Z(n57258) );
  IV U77378 ( .A(n57255), .Z(n57257) );
  XOR U77379 ( .A(n62249), .B(n62254), .Z(n57256) );
  NOR U77380 ( .A(n57257), .B(n57256), .Z(n67709) );
  NOR U77381 ( .A(n57258), .B(n67709), .Z(n61631) );
  XOR U77382 ( .A(n57259), .B(n61631), .Z(n61628) );
  XOR U77383 ( .A(n61626), .B(n61628), .Z(n62271) );
  IV U77384 ( .A(n62271), .Z(n57266) );
  NOR U77385 ( .A(n57261), .B(n57260), .Z(n61629) );
  IV U77386 ( .A(n57262), .Z(n57264) );
  NOR U77387 ( .A(n57264), .B(n57263), .Z(n62269) );
  NOR U77388 ( .A(n61629), .B(n62269), .Z(n57265) );
  XOR U77389 ( .A(n57266), .B(n57265), .Z(n62274) );
  XOR U77390 ( .A(n62272), .B(n62274), .Z(n61624) );
  XOR U77391 ( .A(n57267), .B(n61624), .Z(n57268) );
  IV U77392 ( .A(n57268), .Z(n61617) );
  XOR U77393 ( .A(n61615), .B(n61617), .Z(n62287) );
  XOR U77394 ( .A(n61618), .B(n62287), .Z(n57269) );
  XOR U77395 ( .A(n57270), .B(n57269), .Z(n62291) );
  XOR U77396 ( .A(n57271), .B(n62291), .Z(n62292) );
  XOR U77397 ( .A(n62293), .B(n62292), .Z(n61609) );
  XOR U77398 ( .A(n57272), .B(n61609), .Z(n61600) );
  XOR U77399 ( .A(n57273), .B(n61600), .Z(n67137) );
  XOR U77400 ( .A(n62302), .B(n67137), .Z(n62303) );
  NOR U77401 ( .A(n57275), .B(n57274), .Z(n67127) );
  NOR U77402 ( .A(n57277), .B(n57276), .Z(n67132) );
  NOR U77403 ( .A(n67127), .B(n67132), .Z(n62304) );
  XOR U77404 ( .A(n62303), .B(n62304), .Z(n62310) );
  XOR U77405 ( .A(n62309), .B(n62310), .Z(n62317) );
  XOR U77406 ( .A(n57278), .B(n62317), .Z(n61591) );
  XOR U77407 ( .A(n61592), .B(n61591), .Z(n67759) );
  IV U77408 ( .A(n57279), .Z(n57280) );
  NOR U77409 ( .A(n57281), .B(n57280), .Z(n61588) );
  IV U77410 ( .A(n57282), .Z(n57283) );
  NOR U77411 ( .A(n57284), .B(n57283), .Z(n67758) );
  IV U77412 ( .A(n57285), .Z(n57286) );
  NOR U77413 ( .A(n57287), .B(n57286), .Z(n67767) );
  NOR U77414 ( .A(n67758), .B(n67767), .Z(n61590) );
  IV U77415 ( .A(n61590), .Z(n57288) );
  NOR U77416 ( .A(n61588), .B(n57288), .Z(n57289) );
  XOR U77417 ( .A(n67759), .B(n57289), .Z(n62332) );
  IV U77418 ( .A(n57290), .Z(n57292) );
  NOR U77419 ( .A(n57292), .B(n57291), .Z(n57293) );
  IV U77420 ( .A(n57293), .Z(n62333) );
  XOR U77421 ( .A(n62332), .B(n62333), .Z(n62337) );
  XOR U77422 ( .A(n62335), .B(n62337), .Z(n61583) );
  XOR U77423 ( .A(n61582), .B(n61583), .Z(n61587) );
  XOR U77424 ( .A(n61585), .B(n61587), .Z(n62342) );
  XOR U77425 ( .A(n57294), .B(n62342), .Z(n61579) );
  XOR U77426 ( .A(n57295), .B(n61579), .Z(n62349) );
  XOR U77427 ( .A(n62347), .B(n62349), .Z(n62352) );
  XOR U77428 ( .A(n62350), .B(n62352), .Z(n61577) );
  XOR U77429 ( .A(n61576), .B(n61577), .Z(n62368) );
  XOR U77430 ( .A(n62366), .B(n62368), .Z(n61574) );
  XOR U77431 ( .A(n61573), .B(n61574), .Z(n62375) );
  XOR U77432 ( .A(n57296), .B(n62375), .Z(n57297) );
  IV U77433 ( .A(n57297), .Z(n61570) );
  XOR U77434 ( .A(n61569), .B(n61570), .Z(n57298) );
  NOR U77435 ( .A(n57299), .B(n57298), .Z(n62380) );
  IV U77436 ( .A(n57299), .Z(n57300) );
  NOR U77437 ( .A(n61570), .B(n57300), .Z(n78166) );
  NOR U77438 ( .A(n62380), .B(n78166), .Z(n61566) );
  IV U77439 ( .A(n57301), .Z(n57303) );
  NOR U77440 ( .A(n57303), .B(n57302), .Z(n62378) );
  IV U77441 ( .A(n57304), .Z(n57306) );
  NOR U77442 ( .A(n57306), .B(n57305), .Z(n61565) );
  NOR U77443 ( .A(n62378), .B(n61565), .Z(n57307) );
  XOR U77444 ( .A(n61566), .B(n57307), .Z(n61564) );
  XOR U77445 ( .A(n61562), .B(n61564), .Z(n61554) );
  XOR U77446 ( .A(n57308), .B(n61554), .Z(n61546) );
  XOR U77447 ( .A(n57309), .B(n61546), .Z(n62387) );
  XOR U77448 ( .A(n57310), .B(n62387), .Z(n57311) );
  IV U77449 ( .A(n57311), .Z(n67829) );
  XOR U77450 ( .A(n62389), .B(n67829), .Z(n62392) );
  XOR U77451 ( .A(n62391), .B(n62392), .Z(n61544) );
  IV U77452 ( .A(n57312), .Z(n57313) );
  NOR U77453 ( .A(n57314), .B(n57313), .Z(n67827) );
  IV U77454 ( .A(n57315), .Z(n57317) );
  NOR U77455 ( .A(n57317), .B(n57316), .Z(n67078) );
  NOR U77456 ( .A(n67827), .B(n67078), .Z(n61545) );
  XOR U77457 ( .A(n61544), .B(n61545), .Z(n61538) );
  XOR U77458 ( .A(n61539), .B(n61538), .Z(n61543) );
  XOR U77459 ( .A(n61541), .B(n61543), .Z(n61535) );
  XOR U77460 ( .A(n57318), .B(n61535), .Z(n61526) );
  XOR U77461 ( .A(n57319), .B(n61526), .Z(n61521) );
  XOR U77462 ( .A(n57320), .B(n61521), .Z(n62399) );
  XOR U77463 ( .A(n62400), .B(n62399), .Z(n62404) );
  XOR U77464 ( .A(n57321), .B(n62404), .Z(n57322) );
  IV U77465 ( .A(n57322), .Z(n62412) );
  IV U77466 ( .A(n57323), .Z(n57325) );
  NOR U77467 ( .A(n57325), .B(n57324), .Z(n62410) );
  XOR U77468 ( .A(n62412), .B(n62410), .Z(n62420) );
  IV U77469 ( .A(n57326), .Z(n57327) );
  NOR U77470 ( .A(n57328), .B(n57327), .Z(n62413) );
  IV U77471 ( .A(n57329), .Z(n57330) );
  NOR U77472 ( .A(n57330), .B(n57335), .Z(n62418) );
  NOR U77473 ( .A(n62413), .B(n62418), .Z(n57331) );
  XOR U77474 ( .A(n62420), .B(n57331), .Z(n61514) );
  IV U77475 ( .A(n57332), .Z(n61515) );
  NOR U77476 ( .A(n61515), .B(n57333), .Z(n62423) );
  IV U77477 ( .A(n57334), .Z(n57336) );
  NOR U77478 ( .A(n57336), .B(n57335), .Z(n62416) );
  NOR U77479 ( .A(n62423), .B(n62416), .Z(n57337) );
  XOR U77480 ( .A(n61514), .B(n57337), .Z(n67873) );
  XOR U77481 ( .A(n62422), .B(n67873), .Z(n61508) );
  XOR U77482 ( .A(n61509), .B(n61508), .Z(n67880) );
  XOR U77483 ( .A(n61511), .B(n67880), .Z(n62433) );
  IV U77484 ( .A(n57338), .Z(n57340) );
  NOR U77485 ( .A(n57340), .B(n57339), .Z(n62432) );
  IV U77486 ( .A(n57341), .Z(n57343) );
  NOR U77487 ( .A(n57343), .B(n57342), .Z(n62437) );
  NOR U77488 ( .A(n62432), .B(n62437), .Z(n57344) );
  XOR U77489 ( .A(n62433), .B(n57344), .Z(n61506) );
  IV U77490 ( .A(n57345), .Z(n57347) );
  NOR U77491 ( .A(n57347), .B(n57346), .Z(n61504) );
  XOR U77492 ( .A(n61506), .B(n61504), .Z(n62448) );
  XOR U77493 ( .A(n57348), .B(n62448), .Z(n61491) );
  XOR U77494 ( .A(n57349), .B(n61491), .Z(n61499) );
  XOR U77495 ( .A(n57350), .B(n61499), .Z(n61483) );
  XOR U77496 ( .A(n57351), .B(n61483), .Z(n61478) );
  XOR U77497 ( .A(n61477), .B(n61478), .Z(n61481) );
  XOR U77498 ( .A(n61480), .B(n61481), .Z(n61472) );
  XOR U77499 ( .A(n57352), .B(n61472), .Z(n61464) );
  XOR U77500 ( .A(n61469), .B(n61464), .Z(n62465) );
  IV U77501 ( .A(n62465), .Z(n57361) );
  IV U77502 ( .A(n57353), .Z(n61466) );
  NOR U77503 ( .A(n57354), .B(n61466), .Z(n57359) );
  NOR U77504 ( .A(n57356), .B(n57355), .Z(n57357) );
  IV U77505 ( .A(n57357), .Z(n57362) );
  NOR U77506 ( .A(n57358), .B(n57362), .Z(n62463) );
  NOR U77507 ( .A(n57359), .B(n62463), .Z(n57360) );
  XOR U77508 ( .A(n57361), .B(n57360), .Z(n62462) );
  NOR U77509 ( .A(n57363), .B(n57362), .Z(n62460) );
  XOR U77510 ( .A(n62462), .B(n62460), .Z(n61458) );
  NOR U77511 ( .A(n57371), .B(n61458), .Z(n67008) );
  IV U77512 ( .A(n57364), .Z(n67012) );
  IV U77513 ( .A(n57365), .Z(n57366) );
  NOR U77514 ( .A(n67012), .B(n57366), .Z(n61455) );
  IV U77515 ( .A(n57367), .Z(n57368) );
  NOR U77516 ( .A(n67012), .B(n57368), .Z(n61457) );
  NOR U77517 ( .A(n61455), .B(n61457), .Z(n57369) );
  XOR U77518 ( .A(n57369), .B(n61458), .Z(n61451) );
  IV U77519 ( .A(n57377), .Z(n57370) );
  NOR U77520 ( .A(n57370), .B(n57376), .Z(n61452) );
  XOR U77521 ( .A(n61451), .B(n61452), .Z(n57373) );
  NOR U77522 ( .A(n61452), .B(n57371), .Z(n57372) );
  NOR U77523 ( .A(n57373), .B(n57372), .Z(n57374) );
  NOR U77524 ( .A(n67008), .B(n57374), .Z(n57375) );
  IV U77525 ( .A(n57375), .Z(n61450) );
  XOR U77526 ( .A(n57377), .B(n57376), .Z(n57378) );
  NOR U77527 ( .A(n57379), .B(n57378), .Z(n57380) );
  IV U77528 ( .A(n57380), .Z(n57381) );
  NOR U77529 ( .A(n57382), .B(n57381), .Z(n61448) );
  XOR U77530 ( .A(n61450), .B(n61448), .Z(n62470) );
  XOR U77531 ( .A(n57383), .B(n62470), .Z(n61443) );
  IV U77532 ( .A(n57384), .Z(n57386) );
  NOR U77533 ( .A(n57386), .B(n57385), .Z(n62472) );
  IV U77534 ( .A(n57387), .Z(n57388) );
  NOR U77535 ( .A(n57389), .B(n57388), .Z(n61442) );
  NOR U77536 ( .A(n62472), .B(n61442), .Z(n57390) );
  XOR U77537 ( .A(n61443), .B(n57390), .Z(n61439) );
  XOR U77538 ( .A(n61436), .B(n61439), .Z(n61434) );
  XOR U77539 ( .A(n57391), .B(n61434), .Z(n61431) );
  XOR U77540 ( .A(n61432), .B(n61431), .Z(n62481) );
  XOR U77541 ( .A(n62480), .B(n62481), .Z(n62485) );
  XOR U77542 ( .A(n62483), .B(n62485), .Z(n61430) );
  XOR U77543 ( .A(n61428), .B(n61430), .Z(n62501) );
  XOR U77544 ( .A(n62500), .B(n62501), .Z(n61427) );
  XOR U77545 ( .A(n61425), .B(n61427), .Z(n62509) );
  XOR U77546 ( .A(n62507), .B(n62509), .Z(n66989) );
  XOR U77547 ( .A(n62510), .B(n66989), .Z(n61423) );
  IV U77548 ( .A(n57392), .Z(n57394) );
  NOR U77549 ( .A(n57394), .B(n57393), .Z(n61422) );
  NOR U77550 ( .A(n61422), .B(n62513), .Z(n57395) );
  XOR U77551 ( .A(n61423), .B(n57395), .Z(n61419) );
  XOR U77552 ( .A(n61418), .B(n61419), .Z(n61409) );
  XOR U77553 ( .A(n57396), .B(n61409), .Z(n61412) );
  XOR U77554 ( .A(n57397), .B(n61412), .Z(n57398) );
  IV U77555 ( .A(n57398), .Z(n61407) );
  IV U77556 ( .A(n57399), .Z(n57400) );
  NOR U77557 ( .A(n57401), .B(n57400), .Z(n57407) );
  IV U77558 ( .A(n57402), .Z(n57403) );
  NOR U77559 ( .A(n57403), .B(n57409), .Z(n57404) );
  IV U77560 ( .A(n57404), .Z(n57405) );
  NOR U77561 ( .A(n57407), .B(n57405), .Z(n57417) );
  IV U77562 ( .A(n57417), .Z(n57406) );
  NOR U77563 ( .A(n61407), .B(n57406), .Z(n67964) );
  IV U77564 ( .A(n57407), .Z(n57408) );
  NOR U77565 ( .A(n57409), .B(n57408), .Z(n57410) );
  IV U77566 ( .A(n57410), .Z(n57415) );
  NOR U77567 ( .A(n57412), .B(n57411), .Z(n57413) );
  IV U77568 ( .A(n57413), .Z(n57414) );
  NOR U77569 ( .A(n57415), .B(n57414), .Z(n61405) );
  XOR U77570 ( .A(n61405), .B(n61407), .Z(n57421) );
  IV U77571 ( .A(n57421), .Z(n57416) );
  NOR U77572 ( .A(n57417), .B(n57416), .Z(n57418) );
  NOR U77573 ( .A(n67964), .B(n57418), .Z(n57419) );
  NOR U77574 ( .A(n57420), .B(n57419), .Z(n57423) );
  IV U77575 ( .A(n57420), .Z(n57422) );
  NOR U77576 ( .A(n57422), .B(n57421), .Z(n67967) );
  NOR U77577 ( .A(n57423), .B(n67967), .Z(n61397) );
  XOR U77578 ( .A(n57424), .B(n61397), .Z(n62531) );
  IV U77579 ( .A(n57425), .Z(n57427) );
  NOR U77580 ( .A(n57427), .B(n57426), .Z(n61399) );
  IV U77581 ( .A(n57428), .Z(n57441) );
  IV U77582 ( .A(n57429), .Z(n57430) );
  NOR U77583 ( .A(n57431), .B(n57430), .Z(n57439) );
  NOR U77584 ( .A(n57433), .B(n57432), .Z(n57434) );
  IV U77585 ( .A(n57434), .Z(n57436) );
  NOR U77586 ( .A(n57436), .B(n57435), .Z(n57437) );
  IV U77587 ( .A(n57437), .Z(n57438) );
  NOR U77588 ( .A(n57439), .B(n57438), .Z(n57440) );
  IV U77589 ( .A(n57440), .Z(n57445) );
  NOR U77590 ( .A(n57441), .B(n57445), .Z(n62529) );
  NOR U77591 ( .A(n61399), .B(n62529), .Z(n57442) );
  XOR U77592 ( .A(n62531), .B(n57442), .Z(n57443) );
  IV U77593 ( .A(n57443), .Z(n62536) );
  IV U77594 ( .A(n57444), .Z(n57446) );
  NOR U77595 ( .A(n57446), .B(n57445), .Z(n62534) );
  XOR U77596 ( .A(n62536), .B(n62534), .Z(n67996) );
  XOR U77597 ( .A(n62532), .B(n67996), .Z(n62546) );
  XOR U77598 ( .A(n62548), .B(n62546), .Z(n66976) );
  IV U77599 ( .A(n57447), .Z(n57449) );
  NOR U77600 ( .A(n57449), .B(n57448), .Z(n68006) );
  IV U77601 ( .A(n57450), .Z(n57452) );
  NOR U77602 ( .A(n57452), .B(n57451), .Z(n66975) );
  NOR U77603 ( .A(n68006), .B(n66975), .Z(n62549) );
  XOR U77604 ( .A(n66976), .B(n62549), .Z(n57458) );
  IV U77605 ( .A(n57458), .Z(n61392) );
  NOR U77606 ( .A(n57462), .B(n61392), .Z(n68018) );
  NOR U77607 ( .A(n57453), .B(n61393), .Z(n57457) );
  IV U77608 ( .A(n57454), .Z(n57455) );
  NOR U77609 ( .A(n57456), .B(n57455), .Z(n61389) );
  NOR U77610 ( .A(n57457), .B(n61389), .Z(n57459) );
  XOR U77611 ( .A(n57459), .B(n57458), .Z(n61388) );
  IV U77612 ( .A(n57460), .Z(n57461) );
  NOR U77613 ( .A(n57461), .B(n57468), .Z(n57463) );
  IV U77614 ( .A(n57463), .Z(n61387) );
  XOR U77615 ( .A(n61388), .B(n61387), .Z(n57465) );
  NOR U77616 ( .A(n57463), .B(n57462), .Z(n57464) );
  NOR U77617 ( .A(n57465), .B(n57464), .Z(n57466) );
  NOR U77618 ( .A(n68018), .B(n57466), .Z(n61385) );
  IV U77619 ( .A(n57467), .Z(n57469) );
  NOR U77620 ( .A(n57469), .B(n57468), .Z(n61384) );
  NOR U77621 ( .A(n62565), .B(n61384), .Z(n57470) );
  XOR U77622 ( .A(n61385), .B(n57470), .Z(n62564) );
  IV U77623 ( .A(n57471), .Z(n57474) );
  IV U77624 ( .A(n57472), .Z(n57473) );
  NOR U77625 ( .A(n57474), .B(n57473), .Z(n62562) );
  NOR U77626 ( .A(n57476), .B(n57475), .Z(n61382) );
  NOR U77627 ( .A(n62562), .B(n61382), .Z(n57477) );
  XOR U77628 ( .A(n62564), .B(n57477), .Z(n57478) );
  IV U77629 ( .A(n57478), .Z(n62576) );
  IV U77630 ( .A(n57479), .Z(n57480) );
  NOR U77631 ( .A(n57480), .B(n57482), .Z(n62574) );
  XOR U77632 ( .A(n62576), .B(n62574), .Z(n62579) );
  IV U77633 ( .A(n57481), .Z(n57483) );
  NOR U77634 ( .A(n57483), .B(n57482), .Z(n62577) );
  XOR U77635 ( .A(n62579), .B(n62577), .Z(n66952) );
  IV U77636 ( .A(n57484), .Z(n57486) );
  NOR U77637 ( .A(n57486), .B(n57485), .Z(n71775) );
  IV U77638 ( .A(n57487), .Z(n57488) );
  NOR U77639 ( .A(n57489), .B(n57488), .Z(n72907) );
  NOR U77640 ( .A(n71775), .B(n72907), .Z(n66955) );
  XOR U77641 ( .A(n66952), .B(n66955), .Z(n62581) );
  XOR U77642 ( .A(n62583), .B(n62581), .Z(n62593) );
  XOR U77643 ( .A(n62592), .B(n62593), .Z(n62590) );
  IV U77644 ( .A(n57490), .Z(n57491) );
  NOR U77645 ( .A(n57492), .B(n57491), .Z(n62589) );
  IV U77646 ( .A(n57493), .Z(n57495) );
  NOR U77647 ( .A(n57495), .B(n57494), .Z(n61380) );
  NOR U77648 ( .A(n62589), .B(n61380), .Z(n57496) );
  XOR U77649 ( .A(n62590), .B(n57496), .Z(n57497) );
  NOR U77650 ( .A(n57498), .B(n57497), .Z(n57501) );
  IV U77651 ( .A(n57498), .Z(n57500) );
  XOR U77652 ( .A(n62589), .B(n62590), .Z(n57499) );
  NOR U77653 ( .A(n57500), .B(n57499), .Z(n68057) );
  NOR U77654 ( .A(n57501), .B(n68057), .Z(n61376) );
  XOR U77655 ( .A(n62606), .B(n61376), .Z(n62608) );
  XOR U77656 ( .A(n57502), .B(n62608), .Z(n61369) );
  XOR U77657 ( .A(n61370), .B(n61369), .Z(n61373) );
  IV U77658 ( .A(n57505), .Z(n57503) );
  NOR U77659 ( .A(n57504), .B(n57503), .Z(n61372) );
  IV U77660 ( .A(n61363), .Z(n57506) );
  XOR U77661 ( .A(n57505), .B(n57504), .Z(n61362) );
  NOR U77662 ( .A(n57506), .B(n61362), .Z(n61360) );
  NOR U77663 ( .A(n61372), .B(n61360), .Z(n57507) );
  XOR U77664 ( .A(n61373), .B(n57507), .Z(n61364) );
  XOR U77665 ( .A(n57508), .B(n61364), .Z(n62618) );
  XOR U77666 ( .A(n57509), .B(n62618), .Z(n62624) );
  XOR U77667 ( .A(n62626), .B(n62624), .Z(n66922) );
  XOR U77668 ( .A(n62627), .B(n66922), .Z(n62632) );
  IV U77669 ( .A(n62632), .Z(n68089) );
  XOR U77670 ( .A(n62633), .B(n68089), .Z(n61356) );
  IV U77671 ( .A(n61356), .Z(n57515) );
  IV U77672 ( .A(n57510), .Z(n68095) );
  NOR U77673 ( .A(n68095), .B(n68092), .Z(n62631) );
  IV U77674 ( .A(n57511), .Z(n57513) );
  NOR U77675 ( .A(n57513), .B(n57512), .Z(n61355) );
  NOR U77676 ( .A(n62631), .B(n61355), .Z(n57514) );
  XOR U77677 ( .A(n57515), .B(n57514), .Z(n61354) );
  IV U77678 ( .A(n57516), .Z(n57518) );
  NOR U77679 ( .A(n57518), .B(n57517), .Z(n61352) );
  XOR U77680 ( .A(n61354), .B(n61352), .Z(n62646) );
  XOR U77681 ( .A(n57519), .B(n62646), .Z(n62639) );
  IV U77682 ( .A(n57520), .Z(n57521) );
  NOR U77683 ( .A(n57522), .B(n57521), .Z(n62638) );
  IV U77684 ( .A(n57523), .Z(n57524) );
  NOR U77685 ( .A(n57524), .B(n57529), .Z(n62654) );
  NOR U77686 ( .A(n62638), .B(n62654), .Z(n57525) );
  XOR U77687 ( .A(n62639), .B(n57525), .Z(n61351) );
  IV U77688 ( .A(n57526), .Z(n57527) );
  NOR U77689 ( .A(n57527), .B(n57529), .Z(n61347) );
  IV U77690 ( .A(n57528), .Z(n57530) );
  NOR U77691 ( .A(n57530), .B(n57529), .Z(n61349) );
  NOR U77692 ( .A(n61347), .B(n61349), .Z(n57531) );
  XOR U77693 ( .A(n61351), .B(n57531), .Z(n61341) );
  IV U77694 ( .A(n57534), .Z(n57545) );
  IV U77695 ( .A(n57532), .Z(n57535) );
  NOR U77696 ( .A(n57545), .B(n57535), .Z(n61344) );
  IV U77697 ( .A(n57533), .Z(n57537) );
  XOR U77698 ( .A(n57535), .B(n57534), .Z(n57536) );
  NOR U77699 ( .A(n57537), .B(n57536), .Z(n57538) );
  IV U77700 ( .A(n57538), .Z(n57539) );
  NOR U77701 ( .A(n57540), .B(n57539), .Z(n61340) );
  NOR U77702 ( .A(n61344), .B(n61340), .Z(n57541) );
  XOR U77703 ( .A(n61341), .B(n57541), .Z(n62665) );
  IV U77704 ( .A(n57542), .Z(n57548) );
  IV U77705 ( .A(n57543), .Z(n57544) );
  NOR U77706 ( .A(n57545), .B(n57544), .Z(n57546) );
  IV U77707 ( .A(n57546), .Z(n57547) );
  NOR U77708 ( .A(n57548), .B(n57547), .Z(n57549) );
  IV U77709 ( .A(n57549), .Z(n62664) );
  XOR U77710 ( .A(n62665), .B(n62664), .Z(n57550) );
  XOR U77711 ( .A(n57551), .B(n57550), .Z(n62674) );
  XOR U77712 ( .A(n62673), .B(n62674), .Z(n62686) );
  XOR U77713 ( .A(n57552), .B(n62686), .Z(n62680) );
  XOR U77714 ( .A(n62681), .B(n62680), .Z(n62693) );
  XOR U77715 ( .A(n62692), .B(n62693), .Z(n62696) );
  XOR U77716 ( .A(n62695), .B(n62696), .Z(n62701) );
  XOR U77717 ( .A(n57553), .B(n62701), .Z(n57554) );
  IV U77718 ( .A(n57554), .Z(n61333) );
  XOR U77719 ( .A(n61331), .B(n61333), .Z(n61336) );
  IV U77720 ( .A(n57555), .Z(n57556) );
  NOR U77721 ( .A(n57557), .B(n57556), .Z(n61334) );
  XOR U77722 ( .A(n61336), .B(n61334), .Z(n68160) );
  XOR U77723 ( .A(n62703), .B(n68160), .Z(n62705) );
  XOR U77724 ( .A(n57558), .B(n62705), .Z(n62717) );
  XOR U77725 ( .A(n57559), .B(n62717), .Z(n62719) );
  XOR U77726 ( .A(n62718), .B(n62719), .Z(n62723) );
  XOR U77727 ( .A(n62721), .B(n62723), .Z(n62726) );
  XOR U77728 ( .A(n62725), .B(n62726), .Z(n62730) );
  XOR U77729 ( .A(n62728), .B(n62730), .Z(n66867) );
  XOR U77730 ( .A(n62732), .B(n66867), .Z(n62737) );
  XOR U77731 ( .A(n57560), .B(n62737), .Z(n61326) );
  XOR U77732 ( .A(n57561), .B(n61326), .Z(n62740) );
  XOR U77733 ( .A(n62738), .B(n62740), .Z(n62742) );
  XOR U77734 ( .A(n62741), .B(n62742), .Z(n61320) );
  XOR U77735 ( .A(n61319), .B(n61320), .Z(n61323) );
  IV U77736 ( .A(n57562), .Z(n57566) );
  NOR U77737 ( .A(n57566), .B(n57563), .Z(n61322) );
  IV U77738 ( .A(n57564), .Z(n57568) );
  XOR U77739 ( .A(n57566), .B(n57565), .Z(n57567) );
  NOR U77740 ( .A(n57568), .B(n57567), .Z(n61317) );
  NOR U77741 ( .A(n61322), .B(n61317), .Z(n57569) );
  XOR U77742 ( .A(n61323), .B(n57569), .Z(n62746) );
  XOR U77743 ( .A(n62747), .B(n62746), .Z(n62748) );
  XOR U77744 ( .A(n62749), .B(n62748), .Z(n61307) );
  NOR U77745 ( .A(n57570), .B(n61311), .Z(n57574) );
  IV U77746 ( .A(n57571), .Z(n57573) );
  NOR U77747 ( .A(n57573), .B(n57572), .Z(n61306) );
  NOR U77748 ( .A(n57574), .B(n61306), .Z(n57575) );
  XOR U77749 ( .A(n61307), .B(n57575), .Z(n62765) );
  IV U77750 ( .A(n57576), .Z(n57578) );
  NOR U77751 ( .A(n57578), .B(n57577), .Z(n62758) );
  IV U77752 ( .A(n57579), .Z(n57583) );
  NOR U77753 ( .A(n57581), .B(n57580), .Z(n57582) );
  IV U77754 ( .A(n57582), .Z(n57593) );
  NOR U77755 ( .A(n57583), .B(n57593), .Z(n62763) );
  NOR U77756 ( .A(n62758), .B(n62763), .Z(n57584) );
  XOR U77757 ( .A(n62765), .B(n57584), .Z(n61304) );
  IV U77758 ( .A(n57585), .Z(n57586) );
  NOR U77759 ( .A(n57587), .B(n57586), .Z(n61303) );
  XOR U77760 ( .A(n57589), .B(n57588), .Z(n57590) );
  NOR U77761 ( .A(n57591), .B(n57590), .Z(n57592) );
  IV U77762 ( .A(n57592), .Z(n57594) );
  NOR U77763 ( .A(n57594), .B(n57593), .Z(n62760) );
  NOR U77764 ( .A(n61303), .B(n62760), .Z(n57595) );
  XOR U77765 ( .A(n61304), .B(n57595), .Z(n66824) );
  XOR U77766 ( .A(n61296), .B(n66824), .Z(n61294) );
  NOR U77767 ( .A(n57596), .B(n61299), .Z(n57600) );
  IV U77768 ( .A(n57597), .Z(n57599) );
  NOR U77769 ( .A(n57599), .B(n57598), .Z(n61293) );
  NOR U77770 ( .A(n57600), .B(n61293), .Z(n57601) );
  XOR U77771 ( .A(n61294), .B(n57601), .Z(n62780) );
  IV U77772 ( .A(n57602), .Z(n57603) );
  NOR U77773 ( .A(n57604), .B(n57603), .Z(n62778) );
  NOR U77774 ( .A(n57605), .B(n61290), .Z(n57606) );
  NOR U77775 ( .A(n62778), .B(n57606), .Z(n57607) );
  XOR U77776 ( .A(n62780), .B(n57607), .Z(n62790) );
  IV U77777 ( .A(n57608), .Z(n57610) );
  NOR U77778 ( .A(n57610), .B(n57609), .Z(n66811) );
  NOR U77779 ( .A(n57612), .B(n57611), .Z(n57613) );
  IV U77780 ( .A(n57613), .Z(n57614) );
  NOR U77781 ( .A(n57615), .B(n57614), .Z(n68207) );
  NOR U77782 ( .A(n66811), .B(n68207), .Z(n62791) );
  XOR U77783 ( .A(n62790), .B(n62791), .Z(n62800) );
  XOR U77784 ( .A(n62792), .B(n62800), .Z(n57616) );
  NOR U77785 ( .A(n57617), .B(n57616), .Z(n78589) );
  IV U77786 ( .A(n57618), .Z(n62786) );
  NOR U77787 ( .A(n57619), .B(n62786), .Z(n62799) );
  NOR U77788 ( .A(n62799), .B(n62792), .Z(n57620) );
  XOR U77789 ( .A(n62800), .B(n57620), .Z(n57621) );
  NOR U77790 ( .A(n57622), .B(n57621), .Z(n61287) );
  NOR U77791 ( .A(n78589), .B(n61287), .Z(n61281) );
  IV U77792 ( .A(n57623), .Z(n77143) );
  NOR U77793 ( .A(n77143), .B(n57628), .Z(n61285) );
  IV U77794 ( .A(n57624), .Z(n57626) );
  NOR U77795 ( .A(n57626), .B(n57625), .Z(n61280) );
  NOR U77796 ( .A(n61285), .B(n61280), .Z(n57627) );
  XOR U77797 ( .A(n61281), .B(n57627), .Z(n61279) );
  XOR U77798 ( .A(n57629), .B(n57628), .Z(n57632) );
  IV U77799 ( .A(n57630), .Z(n57631) );
  NOR U77800 ( .A(n57632), .B(n57631), .Z(n61277) );
  XOR U77801 ( .A(n61279), .B(n61277), .Z(n61273) );
  XOR U77802 ( .A(n61271), .B(n61273), .Z(n61275) );
  XOR U77803 ( .A(n57633), .B(n61275), .Z(n57634) );
  IV U77804 ( .A(n57634), .Z(n61268) );
  XOR U77805 ( .A(n61266), .B(n61268), .Z(n61261) );
  IV U77806 ( .A(n57635), .Z(n57637) );
  NOR U77807 ( .A(n57637), .B(n57636), .Z(n61259) );
  XOR U77808 ( .A(n61261), .B(n61259), .Z(n61263) );
  IV U77809 ( .A(n57638), .Z(n57639) );
  NOR U77810 ( .A(n57640), .B(n57639), .Z(n61262) );
  IV U77811 ( .A(n57641), .Z(n57643) );
  NOR U77812 ( .A(n57643), .B(n57642), .Z(n61257) );
  NOR U77813 ( .A(n61262), .B(n61257), .Z(n57644) );
  XOR U77814 ( .A(n61263), .B(n57644), .Z(n57645) );
  IV U77815 ( .A(n57645), .Z(n61256) );
  NOR U77816 ( .A(n57647), .B(n57646), .Z(n57648) );
  IV U77817 ( .A(n57648), .Z(n57656) );
  IV U77818 ( .A(n57649), .Z(n57653) );
  XOR U77819 ( .A(n57651), .B(n57650), .Z(n57652) );
  NOR U77820 ( .A(n57653), .B(n57652), .Z(n57654) );
  IV U77821 ( .A(n57654), .Z(n57655) );
  NOR U77822 ( .A(n57656), .B(n57655), .Z(n61254) );
  XOR U77823 ( .A(n61256), .B(n61254), .Z(n62810) );
  XOR U77824 ( .A(n62809), .B(n62810), .Z(n66774) );
  XOR U77825 ( .A(n62812), .B(n66774), .Z(n61246) );
  IV U77826 ( .A(n57657), .Z(n57658) );
  NOR U77827 ( .A(n57659), .B(n57658), .Z(n61245) );
  IV U77828 ( .A(n57660), .Z(n57662) );
  NOR U77829 ( .A(n57662), .B(n57661), .Z(n61251) );
  NOR U77830 ( .A(n61245), .B(n61251), .Z(n57663) );
  XOR U77831 ( .A(n61246), .B(n57663), .Z(n61249) );
  XOR U77832 ( .A(n61248), .B(n61249), .Z(n61242) );
  XOR U77833 ( .A(n61241), .B(n61242), .Z(n62817) );
  XOR U77834 ( .A(n62816), .B(n62817), .Z(n62820) );
  XOR U77835 ( .A(n62819), .B(n62820), .Z(n62825) );
  XOR U77836 ( .A(n57664), .B(n62825), .Z(n61233) );
  XOR U77837 ( .A(n61234), .B(n61233), .Z(n61237) );
  XOR U77838 ( .A(n61236), .B(n61237), .Z(n66756) );
  IV U77839 ( .A(n57665), .Z(n57666) );
  NOR U77840 ( .A(n57667), .B(n57666), .Z(n66755) );
  IV U77841 ( .A(n57668), .Z(n57670) );
  NOR U77842 ( .A(n57670), .B(n57669), .Z(n68248) );
  NOR U77843 ( .A(n66755), .B(n68248), .Z(n61228) );
  XOR U77844 ( .A(n66756), .B(n61228), .Z(n61230) );
  XOR U77845 ( .A(n57671), .B(n61230), .Z(n61226) );
  XOR U77846 ( .A(n61224), .B(n61226), .Z(n62830) );
  IV U77847 ( .A(n57672), .Z(n57673) );
  NOR U77848 ( .A(n57674), .B(n57673), .Z(n62829) );
  IV U77849 ( .A(n57675), .Z(n57676) );
  NOR U77850 ( .A(n57677), .B(n57676), .Z(n61219) );
  NOR U77851 ( .A(n62829), .B(n61219), .Z(n57678) );
  XOR U77852 ( .A(n62830), .B(n57678), .Z(n61221) );
  XOR U77853 ( .A(n61222), .B(n61221), .Z(n61214) );
  XOR U77854 ( .A(n61213), .B(n61214), .Z(n61208) );
  XOR U77855 ( .A(n57679), .B(n61208), .Z(n66741) );
  IV U77856 ( .A(n57680), .Z(n57682) );
  IV U77857 ( .A(n57681), .Z(n57686) );
  NOR U77858 ( .A(n57682), .B(n57686), .Z(n61204) );
  NOR U77859 ( .A(n57684), .B(n57683), .Z(n68271) );
  IV U77860 ( .A(n57685), .Z(n57687) );
  NOR U77861 ( .A(n57687), .B(n57686), .Z(n66739) );
  NOR U77862 ( .A(n68271), .B(n66739), .Z(n61206) );
  IV U77863 ( .A(n61206), .Z(n57691) );
  NOR U77864 ( .A(n61204), .B(n57691), .Z(n57688) );
  XOR U77865 ( .A(n66741), .B(n57688), .Z(n57689) );
  NOR U77866 ( .A(n57690), .B(n57689), .Z(n57694) );
  IV U77867 ( .A(n57690), .Z(n57693) );
  XOR U77868 ( .A(n66741), .B(n57691), .Z(n57692) );
  NOR U77869 ( .A(n57693), .B(n57692), .Z(n66735) );
  NOR U77870 ( .A(n57694), .B(n66735), .Z(n57695) );
  IV U77871 ( .A(n57695), .Z(n62844) );
  XOR U77872 ( .A(n62843), .B(n62844), .Z(n68278) );
  IV U77873 ( .A(n57696), .Z(n68283) );
  NOR U77874 ( .A(n68283), .B(n68275), .Z(n57700) );
  IV U77875 ( .A(n57697), .Z(n57699) );
  NOR U77876 ( .A(n57699), .B(n57698), .Z(n68284) );
  NOR U77877 ( .A(n57700), .B(n68284), .Z(n62847) );
  XOR U77878 ( .A(n68278), .B(n62847), .Z(n62849) );
  XOR U77879 ( .A(n57701), .B(n62849), .Z(n68295) );
  XOR U77880 ( .A(n62864), .B(n68295), .Z(n62866) );
  XOR U77881 ( .A(n57702), .B(n62866), .Z(n62874) );
  XOR U77882 ( .A(n62873), .B(n62874), .Z(n62877) );
  XOR U77883 ( .A(n62878), .B(n62877), .Z(n62880) );
  IV U77884 ( .A(n57703), .Z(n62887) );
  NOR U77885 ( .A(n62887), .B(n66706), .Z(n57705) );
  IV U77886 ( .A(n66707), .Z(n57704) );
  NOR U77887 ( .A(n57704), .B(n66706), .Z(n62879) );
  NOR U77888 ( .A(n57705), .B(n62879), .Z(n57706) );
  XOR U77889 ( .A(n62880), .B(n57706), .Z(n62885) );
  IV U77890 ( .A(n57707), .Z(n57709) );
  NOR U77891 ( .A(n57709), .B(n57708), .Z(n62883) );
  XOR U77892 ( .A(n62885), .B(n62883), .Z(n62894) );
  XOR U77893 ( .A(n62891), .B(n62894), .Z(n61199) );
  XOR U77894 ( .A(n57710), .B(n61199), .Z(n61197) );
  IV U77895 ( .A(n57711), .Z(n57713) );
  NOR U77896 ( .A(n57713), .B(n57712), .Z(n61195) );
  XOR U77897 ( .A(n61197), .B(n61195), .Z(n61189) );
  XOR U77898 ( .A(n61188), .B(n61189), .Z(n68307) );
  XOR U77899 ( .A(n61191), .B(n68307), .Z(n61182) );
  XOR U77900 ( .A(n57714), .B(n61182), .Z(n61181) );
  XOR U77901 ( .A(n61179), .B(n61181), .Z(n62904) );
  IV U77902 ( .A(n57715), .Z(n57716) );
  NOR U77903 ( .A(n57717), .B(n57716), .Z(n61176) );
  IV U77904 ( .A(n57718), .Z(n57720) );
  NOR U77905 ( .A(n57720), .B(n57719), .Z(n62903) );
  NOR U77906 ( .A(n61176), .B(n62903), .Z(n57721) );
  XOR U77907 ( .A(n62904), .B(n57721), .Z(n62907) );
  XOR U77908 ( .A(n57722), .B(n62907), .Z(n62912) );
  XOR U77909 ( .A(n62910), .B(n62912), .Z(n62924) );
  IV U77910 ( .A(n57723), .Z(n57724) );
  NOR U77911 ( .A(n57725), .B(n57724), .Z(n62917) );
  IV U77912 ( .A(n57726), .Z(n57727) );
  NOR U77913 ( .A(n57728), .B(n57727), .Z(n62922) );
  NOR U77914 ( .A(n62917), .B(n62922), .Z(n57729) );
  XOR U77915 ( .A(n62924), .B(n57729), .Z(n62919) );
  XOR U77916 ( .A(n62920), .B(n62919), .Z(n61172) );
  XOR U77917 ( .A(n61170), .B(n61172), .Z(n61175) );
  XOR U77918 ( .A(n57730), .B(n61175), .Z(n57731) );
  IV U77919 ( .A(n57731), .Z(n61167) );
  XOR U77920 ( .A(n61165), .B(n61167), .Z(n61163) );
  XOR U77921 ( .A(n61160), .B(n61163), .Z(n61158) );
  IV U77922 ( .A(n61158), .Z(n57738) );
  NOR U77923 ( .A(n57733), .B(n57732), .Z(n61162) );
  IV U77924 ( .A(n57734), .Z(n57736) );
  NOR U77925 ( .A(n57736), .B(n57735), .Z(n61157) );
  NOR U77926 ( .A(n61162), .B(n61157), .Z(n57737) );
  XOR U77927 ( .A(n57738), .B(n57737), .Z(n61156) );
  XOR U77928 ( .A(n61154), .B(n61156), .Z(n61151) );
  XOR U77929 ( .A(n57739), .B(n61151), .Z(n61143) );
  IV U77930 ( .A(n57740), .Z(n57742) );
  NOR U77931 ( .A(n57742), .B(n57741), .Z(n61145) );
  IV U77932 ( .A(n57743), .Z(n57745) );
  NOR U77933 ( .A(n57745), .B(n57744), .Z(n61142) );
  NOR U77934 ( .A(n61145), .B(n61142), .Z(n57746) );
  XOR U77935 ( .A(n61143), .B(n57746), .Z(n62932) );
  XOR U77936 ( .A(n62931), .B(n62932), .Z(n62935) );
  XOR U77937 ( .A(n57747), .B(n62935), .Z(n57748) );
  IV U77938 ( .A(n57748), .Z(n61135) );
  XOR U77939 ( .A(n61134), .B(n61135), .Z(n61139) );
  IV U77940 ( .A(n57749), .Z(n57751) );
  NOR U77941 ( .A(n57751), .B(n57750), .Z(n61137) );
  XOR U77942 ( .A(n61139), .B(n61137), .Z(n66642) );
  IV U77943 ( .A(n57753), .Z(n57752) );
  NOR U77944 ( .A(n57754), .B(n57752), .Z(n66640) );
  XOR U77945 ( .A(n57754), .B(n57753), .Z(n57757) );
  IV U77946 ( .A(n57755), .Z(n57756) );
  NOR U77947 ( .A(n57757), .B(n57756), .Z(n68375) );
  NOR U77948 ( .A(n66640), .B(n68375), .Z(n61130) );
  XOR U77949 ( .A(n66642), .B(n61130), .Z(n66632) );
  XOR U77950 ( .A(n57758), .B(n66632), .Z(n61126) );
  XOR U77951 ( .A(n61125), .B(n61126), .Z(n66619) );
  XOR U77952 ( .A(n57759), .B(n66619), .Z(n61122) );
  IV U77953 ( .A(n57760), .Z(n57761) );
  NOR U77954 ( .A(n57762), .B(n57761), .Z(n61120) );
  XOR U77955 ( .A(n61122), .B(n61120), .Z(n62946) );
  XOR U77956 ( .A(n62943), .B(n62946), .Z(n61118) );
  IV U77957 ( .A(n57763), .Z(n57765) );
  NOR U77958 ( .A(n57765), .B(n57764), .Z(n62945) );
  IV U77959 ( .A(n57766), .Z(n57770) );
  NOR U77960 ( .A(n57768), .B(n57767), .Z(n57769) );
  IV U77961 ( .A(n57769), .Z(n57773) );
  NOR U77962 ( .A(n57770), .B(n57773), .Z(n61116) );
  NOR U77963 ( .A(n62945), .B(n61116), .Z(n57771) );
  XOR U77964 ( .A(n61118), .B(n57771), .Z(n61113) );
  IV U77965 ( .A(n57772), .Z(n57774) );
  NOR U77966 ( .A(n57774), .B(n57773), .Z(n57775) );
  IV U77967 ( .A(n57775), .Z(n61114) );
  XOR U77968 ( .A(n61113), .B(n61114), .Z(n61111) );
  XOR U77969 ( .A(n57776), .B(n61111), .Z(n61100) );
  IV U77970 ( .A(n57777), .Z(n57778) );
  NOR U77971 ( .A(n57779), .B(n57778), .Z(n61107) );
  IV U77972 ( .A(n57780), .Z(n57782) );
  NOR U77973 ( .A(n57782), .B(n57781), .Z(n61099) );
  NOR U77974 ( .A(n61107), .B(n61099), .Z(n57783) );
  XOR U77975 ( .A(n61100), .B(n57783), .Z(n61103) );
  NOR U77976 ( .A(n57790), .B(n61103), .Z(n66596) );
  IV U77977 ( .A(n57784), .Z(n57785) );
  NOR U77978 ( .A(n57786), .B(n57785), .Z(n62956) );
  IV U77979 ( .A(n57787), .Z(n57789) );
  NOR U77980 ( .A(n57789), .B(n57788), .Z(n61102) );
  XOR U77981 ( .A(n61102), .B(n61103), .Z(n62957) );
  IV U77982 ( .A(n62957), .Z(n57791) );
  XOR U77983 ( .A(n62956), .B(n57791), .Z(n57793) );
  NOR U77984 ( .A(n57791), .B(n57790), .Z(n57792) );
  NOR U77985 ( .A(n57793), .B(n57792), .Z(n57794) );
  NOR U77986 ( .A(n66596), .B(n57794), .Z(n61097) );
  IV U77987 ( .A(n57795), .Z(n57797) );
  NOR U77988 ( .A(n57797), .B(n57796), .Z(n62952) );
  IV U77989 ( .A(n57798), .Z(n57800) );
  NOR U77990 ( .A(n57800), .B(n57799), .Z(n61096) );
  NOR U77991 ( .A(n62952), .B(n61096), .Z(n57801) );
  XOR U77992 ( .A(n61097), .B(n57801), .Z(n61095) );
  XOR U77993 ( .A(n61093), .B(n61095), .Z(n61088) );
  XOR U77994 ( .A(n61087), .B(n61088), .Z(n66579) );
  XOR U77995 ( .A(n61090), .B(n66579), .Z(n57802) );
  IV U77996 ( .A(n57802), .Z(n61084) );
  NOR U77997 ( .A(n57803), .B(n57812), .Z(n57804) );
  IV U77998 ( .A(n57804), .Z(n57805) );
  NOR U77999 ( .A(n57806), .B(n57805), .Z(n61082) );
  XOR U78000 ( .A(n61084), .B(n61082), .Z(n62968) );
  IV U78001 ( .A(n57807), .Z(n57809) );
  NOR U78002 ( .A(n57809), .B(n57808), .Z(n62967) );
  IV U78003 ( .A(n57810), .Z(n57811) );
  NOR U78004 ( .A(n57812), .B(n57811), .Z(n61085) );
  NOR U78005 ( .A(n62967), .B(n61085), .Z(n57813) );
  XOR U78006 ( .A(n62968), .B(n57813), .Z(n61080) );
  XOR U78007 ( .A(n57814), .B(n61080), .Z(n61078) );
  XOR U78008 ( .A(n57815), .B(n61078), .Z(n61071) );
  XOR U78009 ( .A(n61073), .B(n61071), .Z(n62979) );
  XOR U78010 ( .A(n62978), .B(n62979), .Z(n62990) );
  XOR U78011 ( .A(n57816), .B(n62990), .Z(n62987) );
  XOR U78012 ( .A(n62985), .B(n62987), .Z(n62994) );
  IV U78013 ( .A(n57817), .Z(n57818) );
  NOR U78014 ( .A(n57824), .B(n57818), .Z(n62992) );
  XOR U78015 ( .A(n62994), .B(n62992), .Z(n62997) );
  IV U78016 ( .A(n57819), .Z(n57821) );
  NOR U78017 ( .A(n57821), .B(n57820), .Z(n61069) );
  IV U78018 ( .A(n57822), .Z(n57823) );
  NOR U78019 ( .A(n57824), .B(n57823), .Z(n62995) );
  NOR U78020 ( .A(n61069), .B(n62995), .Z(n57825) );
  XOR U78021 ( .A(n62997), .B(n57825), .Z(n63000) );
  XOR U78022 ( .A(n57826), .B(n63000), .Z(n63008) );
  XOR U78023 ( .A(n61065), .B(n63008), .Z(n61054) );
  XOR U78024 ( .A(n57827), .B(n61054), .Z(n61052) );
  XOR U78025 ( .A(n57828), .B(n61052), .Z(n61041) );
  XOR U78026 ( .A(n57829), .B(n61041), .Z(n63023) );
  XOR U78027 ( .A(n63021), .B(n63023), .Z(n61038) );
  XOR U78028 ( .A(n61037), .B(n61038), .Z(n66533) );
  IV U78029 ( .A(n66533), .Z(n57836) );
  IV U78030 ( .A(n57830), .Z(n57832) );
  NOR U78031 ( .A(n57832), .B(n57831), .Z(n66536) );
  IV U78032 ( .A(n57833), .Z(n57835) );
  NOR U78033 ( .A(n57835), .B(n57834), .Z(n66531) );
  NOR U78034 ( .A(n66536), .B(n66531), .Z(n61036) );
  XOR U78035 ( .A(n57836), .B(n61036), .Z(n61032) );
  XOR U78036 ( .A(n61031), .B(n61032), .Z(n66522) );
  XOR U78037 ( .A(n61034), .B(n66522), .Z(n61027) );
  IV U78038 ( .A(n57837), .Z(n57838) );
  NOR U78039 ( .A(n57839), .B(n57838), .Z(n61026) );
  IV U78040 ( .A(n61026), .Z(n61024) );
  XOR U78041 ( .A(n61027), .B(n61024), .Z(n61021) );
  IV U78042 ( .A(n61021), .Z(n57847) );
  IV U78043 ( .A(n57840), .Z(n57842) );
  NOR U78044 ( .A(n57842), .B(n57841), .Z(n61028) );
  IV U78045 ( .A(n57843), .Z(n57845) );
  NOR U78046 ( .A(n57845), .B(n57844), .Z(n61020) );
  NOR U78047 ( .A(n61028), .B(n61020), .Z(n57846) );
  XOR U78048 ( .A(n57847), .B(n57846), .Z(n63036) );
  XOR U78049 ( .A(n63034), .B(n63036), .Z(n63038) );
  XOR U78050 ( .A(n57848), .B(n63038), .Z(n61010) );
  XOR U78051 ( .A(n57849), .B(n61010), .Z(n61009) );
  XOR U78052 ( .A(n61007), .B(n61009), .Z(n61002) );
  XOR U78053 ( .A(n61001), .B(n61002), .Z(n61006) );
  XOR U78054 ( .A(n61004), .B(n61006), .Z(n60994) );
  XOR U78055 ( .A(n57850), .B(n60994), .Z(n63047) );
  XOR U78056 ( .A(n57851), .B(n63047), .Z(n63058) );
  XOR U78057 ( .A(n63059), .B(n63058), .Z(n63065) );
  XOR U78058 ( .A(n63066), .B(n63065), .Z(n57852) );
  IV U78059 ( .A(n57852), .Z(n63068) );
  XOR U78060 ( .A(n63067), .B(n63068), .Z(n63074) );
  XOR U78061 ( .A(n63073), .B(n63074), .Z(n60988) );
  XOR U78062 ( .A(n60986), .B(n60988), .Z(n68493) );
  XOR U78063 ( .A(n57853), .B(n68493), .Z(n60984) );
  IV U78064 ( .A(n57854), .Z(n57856) );
  NOR U78065 ( .A(n57856), .B(n57855), .Z(n60982) );
  XOR U78066 ( .A(n60984), .B(n60982), .Z(n60980) );
  IV U78067 ( .A(n57857), .Z(n57858) );
  NOR U78068 ( .A(n57859), .B(n57858), .Z(n60976) );
  IV U78069 ( .A(n57860), .Z(n57862) );
  NOR U78070 ( .A(n57862), .B(n57861), .Z(n60978) );
  NOR U78071 ( .A(n60976), .B(n60978), .Z(n57863) );
  XOR U78072 ( .A(n60980), .B(n57863), .Z(n57864) );
  IV U78073 ( .A(n57864), .Z(n60975) );
  IV U78074 ( .A(n57865), .Z(n57867) );
  NOR U78075 ( .A(n57867), .B(n57866), .Z(n57868) );
  IV U78076 ( .A(n57868), .Z(n57874) );
  NOR U78077 ( .A(n60975), .B(n57874), .Z(n66478) );
  IV U78078 ( .A(n57869), .Z(n57871) );
  NOR U78079 ( .A(n57871), .B(n57870), .Z(n60973) );
  XOR U78080 ( .A(n60973), .B(n60975), .Z(n60972) );
  IV U78081 ( .A(n57872), .Z(n57873) );
  NOR U78082 ( .A(n57873), .B(n57883), .Z(n57875) );
  IV U78083 ( .A(n57875), .Z(n60971) );
  XOR U78084 ( .A(n60972), .B(n60971), .Z(n57877) );
  NOR U78085 ( .A(n57875), .B(n57874), .Z(n57876) );
  NOR U78086 ( .A(n57877), .B(n57876), .Z(n57878) );
  NOR U78087 ( .A(n66478), .B(n57878), .Z(n63087) );
  IV U78088 ( .A(n57879), .Z(n57881) );
  NOR U78089 ( .A(n57881), .B(n57880), .Z(n73454) );
  IV U78090 ( .A(n57882), .Z(n57884) );
  NOR U78091 ( .A(n57884), .B(n57883), .Z(n71412) );
  NOR U78092 ( .A(n73454), .B(n71412), .Z(n63088) );
  XOR U78093 ( .A(n63087), .B(n63088), .Z(n63096) );
  IV U78094 ( .A(n57885), .Z(n57887) );
  NOR U78095 ( .A(n57887), .B(n57886), .Z(n63089) );
  IV U78096 ( .A(n57888), .Z(n57889) );
  NOR U78097 ( .A(n57889), .B(n57892), .Z(n63095) );
  IV U78098 ( .A(n57890), .Z(n57891) );
  NOR U78099 ( .A(n57892), .B(n57891), .Z(n63085) );
  NOR U78100 ( .A(n63095), .B(n63085), .Z(n57893) );
  IV U78101 ( .A(n57893), .Z(n57894) );
  NOR U78102 ( .A(n63089), .B(n57894), .Z(n57895) );
  XOR U78103 ( .A(n63096), .B(n57895), .Z(n57896) );
  IV U78104 ( .A(n57896), .Z(n66467) );
  XOR U78105 ( .A(n63098), .B(n66467), .Z(n73471) );
  IV U78106 ( .A(n57897), .Z(n57898) );
  NOR U78107 ( .A(n57899), .B(n57898), .Z(n76770) );
  IV U78108 ( .A(n57900), .Z(n57902) );
  IV U78109 ( .A(n57901), .Z(n76785) );
  NOR U78110 ( .A(n57902), .B(n76785), .Z(n76774) );
  NOR U78111 ( .A(n76770), .B(n76774), .Z(n73473) );
  XOR U78112 ( .A(n73471), .B(n73473), .Z(n63101) );
  XOR U78113 ( .A(n63102), .B(n63101), .Z(n63111) );
  XOR U78114 ( .A(n63110), .B(n63111), .Z(n63108) );
  XOR U78115 ( .A(n63107), .B(n63108), .Z(n63124) );
  XOR U78116 ( .A(n63123), .B(n63124), .Z(n63127) );
  IV U78117 ( .A(n63127), .Z(n57909) );
  IV U78118 ( .A(n57903), .Z(n57905) );
  NOR U78119 ( .A(n57905), .B(n57904), .Z(n63126) );
  NOR U78120 ( .A(n57907), .B(n57906), .Z(n60966) );
  NOR U78121 ( .A(n63126), .B(n60966), .Z(n57908) );
  XOR U78122 ( .A(n57909), .B(n57908), .Z(n60969) );
  XOR U78123 ( .A(n60968), .B(n60969), .Z(n63134) );
  XOR U78124 ( .A(n57910), .B(n63134), .Z(n63137) );
  XOR U78125 ( .A(n63135), .B(n63137), .Z(n63139) );
  XOR U78126 ( .A(n63138), .B(n63139), .Z(n63144) );
  IV U78127 ( .A(n57911), .Z(n57912) );
  NOR U78128 ( .A(n57913), .B(n57912), .Z(n63142) );
  XOR U78129 ( .A(n63144), .B(n63142), .Z(n63151) );
  IV U78130 ( .A(n57914), .Z(n57916) );
  NOR U78131 ( .A(n57916), .B(n57915), .Z(n63150) );
  IV U78132 ( .A(n57917), .Z(n57919) );
  NOR U78133 ( .A(n57919), .B(n57918), .Z(n63145) );
  NOR U78134 ( .A(n63150), .B(n63145), .Z(n57920) );
  XOR U78135 ( .A(n63151), .B(n57920), .Z(n57921) );
  IV U78136 ( .A(n57921), .Z(n63149) );
  XOR U78137 ( .A(n63147), .B(n63149), .Z(n63165) );
  XOR U78138 ( .A(n63163), .B(n63165), .Z(n63162) );
  XOR U78139 ( .A(n57922), .B(n63162), .Z(n57923) );
  IV U78140 ( .A(n57923), .Z(n63159) );
  XOR U78141 ( .A(n63157), .B(n63159), .Z(n60964) );
  XOR U78142 ( .A(n60963), .B(n60964), .Z(n71355) );
  XOR U78143 ( .A(n60962), .B(n71355), .Z(n63183) );
  XOR U78144 ( .A(n57924), .B(n63183), .Z(n60961) );
  IV U78145 ( .A(n57925), .Z(n57927) );
  NOR U78146 ( .A(n57927), .B(n57926), .Z(n60959) );
  XOR U78147 ( .A(n60961), .B(n60959), .Z(n60953) );
  IV U78148 ( .A(n57928), .Z(n57930) );
  NOR U78149 ( .A(n57930), .B(n57929), .Z(n60951) );
  XOR U78150 ( .A(n60953), .B(n60951), .Z(n60956) );
  NOR U78151 ( .A(n57932), .B(n57931), .Z(n60954) );
  XOR U78152 ( .A(n60956), .B(n60954), .Z(n60946) );
  XOR U78153 ( .A(n60945), .B(n60946), .Z(n60950) );
  IV U78154 ( .A(n57933), .Z(n57935) );
  NOR U78155 ( .A(n57935), .B(n57934), .Z(n57936) );
  IV U78156 ( .A(n57936), .Z(n57937) );
  NOR U78157 ( .A(n57938), .B(n57937), .Z(n60948) );
  XOR U78158 ( .A(n60950), .B(n60948), .Z(n63192) );
  XOR U78159 ( .A(n63191), .B(n63192), .Z(n63199) );
  IV U78160 ( .A(n57939), .Z(n57940) );
  NOR U78161 ( .A(n57941), .B(n57940), .Z(n63194) );
  NOR U78162 ( .A(n57943), .B(n57942), .Z(n63198) );
  NOR U78163 ( .A(n63194), .B(n63198), .Z(n57944) );
  XOR U78164 ( .A(n63199), .B(n57944), .Z(n57945) );
  IV U78165 ( .A(n57945), .Z(n66403) );
  IV U78166 ( .A(n57946), .Z(n57948) );
  IV U78167 ( .A(n57947), .Z(n57950) );
  NOR U78168 ( .A(n57948), .B(n57950), .Z(n66401) );
  NOR U78169 ( .A(n66406), .B(n66401), .Z(n63197) );
  XOR U78170 ( .A(n66403), .B(n63197), .Z(n60940) );
  IV U78171 ( .A(n57949), .Z(n57951) );
  NOR U78172 ( .A(n57951), .B(n57950), .Z(n60942) );
  IV U78173 ( .A(n57952), .Z(n57953) );
  NOR U78174 ( .A(n57954), .B(n57953), .Z(n60939) );
  NOR U78175 ( .A(n60942), .B(n60939), .Z(n57955) );
  XOR U78176 ( .A(n60940), .B(n57955), .Z(n60934) );
  XOR U78177 ( .A(n60933), .B(n60934), .Z(n60937) );
  XOR U78178 ( .A(n60936), .B(n60937), .Z(n60929) );
  XOR U78179 ( .A(n57956), .B(n60929), .Z(n57957) );
  IV U78180 ( .A(n57957), .Z(n60925) );
  XOR U78181 ( .A(n60924), .B(n60925), .Z(n63207) );
  XOR U78182 ( .A(n63206), .B(n63207), .Z(n63213) );
  IV U78183 ( .A(n57958), .Z(n57960) );
  NOR U78184 ( .A(n57960), .B(n57959), .Z(n63209) );
  IV U78185 ( .A(n57961), .Z(n57962) );
  NOR U78186 ( .A(n57963), .B(n57962), .Z(n63212) );
  NOR U78187 ( .A(n63209), .B(n63212), .Z(n57964) );
  XOR U78188 ( .A(n63213), .B(n57964), .Z(n63216) );
  XOR U78189 ( .A(n57965), .B(n63216), .Z(n66375) );
  XOR U78190 ( .A(n57966), .B(n66375), .Z(n63224) );
  XOR U78191 ( .A(n63223), .B(n63224), .Z(n57967) );
  NOR U78192 ( .A(n57968), .B(n57967), .Z(n66369) );
  IV U78193 ( .A(n57969), .Z(n57971) );
  NOR U78194 ( .A(n57971), .B(n57970), .Z(n60920) );
  NOR U78195 ( .A(n63223), .B(n60920), .Z(n57972) );
  XOR U78196 ( .A(n63224), .B(n57972), .Z(n57973) );
  NOR U78197 ( .A(n57974), .B(n57973), .Z(n57975) );
  NOR U78198 ( .A(n66369), .B(n57975), .Z(n57976) );
  IV U78199 ( .A(n57976), .Z(n60919) );
  IV U78200 ( .A(n57977), .Z(n57978) );
  NOR U78201 ( .A(n57979), .B(n57978), .Z(n60917) );
  XOR U78202 ( .A(n60919), .B(n60917), .Z(n63232) );
  IV U78203 ( .A(n57980), .Z(n57981) );
  NOR U78204 ( .A(n57982), .B(n57981), .Z(n63230) );
  XOR U78205 ( .A(n63232), .B(n63230), .Z(n66363) );
  IV U78206 ( .A(n57983), .Z(n57984) );
  NOR U78207 ( .A(n57985), .B(n57984), .Z(n68600) );
  IV U78208 ( .A(n57986), .Z(n57988) );
  NOR U78209 ( .A(n57988), .B(n57987), .Z(n66361) );
  NOR U78210 ( .A(n68600), .B(n66361), .Z(n63233) );
  XOR U78211 ( .A(n66363), .B(n63233), .Z(n60908) );
  XOR U78212 ( .A(n57989), .B(n60908), .Z(n60911) );
  IV U78213 ( .A(n57990), .Z(n57991) );
  NOR U78214 ( .A(n57991), .B(n57993), .Z(n60910) );
  IV U78215 ( .A(n57992), .Z(n57994) );
  NOR U78216 ( .A(n57994), .B(n57993), .Z(n60905) );
  NOR U78217 ( .A(n60910), .B(n60905), .Z(n57995) );
  XOR U78218 ( .A(n60911), .B(n57995), .Z(n60903) );
  XOR U78219 ( .A(n57996), .B(n60903), .Z(n63242) );
  XOR U78220 ( .A(n63240), .B(n63242), .Z(n63244) );
  IV U78221 ( .A(n57999), .Z(n57997) );
  NOR U78222 ( .A(n57997), .B(n57998), .Z(n63243) );
  XOR U78223 ( .A(n57999), .B(n57998), .Z(n58002) );
  IV U78224 ( .A(n58000), .Z(n58001) );
  NOR U78225 ( .A(n58002), .B(n58001), .Z(n60899) );
  NOR U78226 ( .A(n63243), .B(n60899), .Z(n58003) );
  XOR U78227 ( .A(n63244), .B(n58003), .Z(n60893) );
  IV U78228 ( .A(n58004), .Z(n58006) );
  NOR U78229 ( .A(n58006), .B(n58005), .Z(n60896) );
  IV U78230 ( .A(n58007), .Z(n58008) );
  NOR U78231 ( .A(n58011), .B(n58008), .Z(n60894) );
  NOR U78232 ( .A(n60896), .B(n60894), .Z(n58009) );
  XOR U78233 ( .A(n60893), .B(n58009), .Z(n60891) );
  IV U78234 ( .A(n58010), .Z(n58012) );
  NOR U78235 ( .A(n58012), .B(n58011), .Z(n60890) );
  IV U78236 ( .A(n58013), .Z(n58014) );
  NOR U78237 ( .A(n58015), .B(n58014), .Z(n60885) );
  NOR U78238 ( .A(n60890), .B(n60885), .Z(n58016) );
  XOR U78239 ( .A(n60891), .B(n58016), .Z(n60881) );
  XOR U78240 ( .A(n58017), .B(n60881), .Z(n63249) );
  XOR U78241 ( .A(n63248), .B(n63249), .Z(n63252) );
  XOR U78242 ( .A(n63251), .B(n63252), .Z(n60879) );
  XOR U78243 ( .A(n60878), .B(n60879), .Z(n66328) );
  XOR U78244 ( .A(n58023), .B(n66328), .Z(n58018) );
  NOR U78245 ( .A(n58019), .B(n58018), .Z(n60877) );
  IV U78246 ( .A(n58020), .Z(n58022) );
  NOR U78247 ( .A(n58022), .B(n58021), .Z(n63256) );
  NOR U78248 ( .A(n63256), .B(n58023), .Z(n58024) );
  XOR U78249 ( .A(n66328), .B(n58024), .Z(n58025) );
  NOR U78250 ( .A(n58026), .B(n58025), .Z(n58027) );
  NOR U78251 ( .A(n60877), .B(n58027), .Z(n58028) );
  IV U78252 ( .A(n58028), .Z(n63269) );
  XOR U78253 ( .A(n63269), .B(n63268), .Z(n63272) );
  IV U78254 ( .A(n58029), .Z(n58031) );
  NOR U78255 ( .A(n58031), .B(n58030), .Z(n63266) );
  NOR U78256 ( .A(n63271), .B(n63266), .Z(n58032) );
  XOR U78257 ( .A(n63272), .B(n58032), .Z(n58033) );
  NOR U78258 ( .A(n58034), .B(n58033), .Z(n58037) );
  IV U78259 ( .A(n58034), .Z(n58036) );
  XOR U78260 ( .A(n63271), .B(n63272), .Z(n58035) );
  NOR U78261 ( .A(n58036), .B(n58035), .Z(n76634) );
  NOR U78262 ( .A(n58037), .B(n76634), .Z(n58038) );
  IV U78263 ( .A(n58038), .Z(n63278) );
  XOR U78264 ( .A(n63277), .B(n63278), .Z(n63283) );
  IV U78265 ( .A(n58039), .Z(n58040) );
  NOR U78266 ( .A(n58041), .B(n58040), .Z(n60875) );
  IV U78267 ( .A(n58042), .Z(n58043) );
  NOR U78268 ( .A(n58044), .B(n58043), .Z(n63281) );
  NOR U78269 ( .A(n60875), .B(n63281), .Z(n58045) );
  XOR U78270 ( .A(n63283), .B(n58045), .Z(n60872) );
  XOR U78271 ( .A(n58046), .B(n60872), .Z(n60871) );
  XOR U78272 ( .A(n60869), .B(n60871), .Z(n63294) );
  IV U78273 ( .A(n58047), .Z(n58048) );
  NOR U78274 ( .A(n58049), .B(n58048), .Z(n63293) );
  IV U78275 ( .A(n58050), .Z(n58052) );
  NOR U78276 ( .A(n58052), .B(n58051), .Z(n63290) );
  NOR U78277 ( .A(n63293), .B(n63290), .Z(n58053) );
  XOR U78278 ( .A(n63294), .B(n58053), .Z(n60865) );
  NOR U78279 ( .A(n58054), .B(n60866), .Z(n58058) );
  IV U78280 ( .A(n58055), .Z(n58057) );
  NOR U78281 ( .A(n58057), .B(n58056), .Z(n63301) );
  NOR U78282 ( .A(n58058), .B(n63301), .Z(n58059) );
  XOR U78283 ( .A(n60865), .B(n58059), .Z(n63310) );
  XOR U78284 ( .A(n63308), .B(n63310), .Z(n63312) );
  XOR U78285 ( .A(n63311), .B(n63312), .Z(n71251) );
  IV U78286 ( .A(n58060), .Z(n58062) );
  NOR U78287 ( .A(n58062), .B(n58061), .Z(n71247) );
  NOR U78288 ( .A(n73646), .B(n71247), .Z(n60860) );
  XOR U78289 ( .A(n71251), .B(n60860), .Z(n60861) );
  XOR U78290 ( .A(n60863), .B(n60861), .Z(n60856) );
  XOR U78291 ( .A(n60855), .B(n60856), .Z(n63318) );
  XOR U78292 ( .A(n58063), .B(n63318), .Z(n60852) );
  XOR U78293 ( .A(n58064), .B(n60852), .Z(n60851) );
  XOR U78294 ( .A(n60849), .B(n60851), .Z(n60844) );
  XOR U78295 ( .A(n60843), .B(n60844), .Z(n60847) );
  XOR U78296 ( .A(n60846), .B(n60847), .Z(n60838) );
  XOR U78297 ( .A(n60837), .B(n60838), .Z(n60841) );
  XOR U78298 ( .A(n60840), .B(n60841), .Z(n60833) );
  XOR U78299 ( .A(n58065), .B(n60833), .Z(n68703) );
  NOR U78300 ( .A(n58066), .B(n68703), .Z(n58069) );
  IV U78301 ( .A(n58066), .Z(n58068) );
  XOR U78302 ( .A(n60830), .B(n60833), .Z(n58067) );
  NOR U78303 ( .A(n58068), .B(n58067), .Z(n68708) );
  NOR U78304 ( .A(n58069), .B(n68708), .Z(n60826) );
  IV U78305 ( .A(n58070), .Z(n58072) );
  NOR U78306 ( .A(n58072), .B(n58071), .Z(n58073) );
  IV U78307 ( .A(n58073), .Z(n68707) );
  XOR U78308 ( .A(n60826), .B(n68707), .Z(n66263) );
  XOR U78309 ( .A(n58074), .B(n66263), .Z(n60824) );
  XOR U78310 ( .A(n60823), .B(n60824), .Z(n60819) );
  IV U78311 ( .A(n58075), .Z(n58076) );
  NOR U78312 ( .A(n58077), .B(n58076), .Z(n63343) );
  IV U78313 ( .A(n58078), .Z(n58080) );
  NOR U78314 ( .A(n58080), .B(n58079), .Z(n60820) );
  NOR U78315 ( .A(n63343), .B(n60820), .Z(n58081) );
  XOR U78316 ( .A(n60819), .B(n58081), .Z(n60818) );
  XOR U78317 ( .A(n60816), .B(n60818), .Z(n60814) );
  XOR U78318 ( .A(n60813), .B(n60814), .Z(n63350) );
  XOR U78319 ( .A(n63349), .B(n63350), .Z(n63362) );
  IV U78320 ( .A(n58082), .Z(n58083) );
  NOR U78321 ( .A(n58084), .B(n58083), .Z(n60811) );
  IV U78322 ( .A(n58085), .Z(n58087) );
  NOR U78323 ( .A(n58087), .B(n58086), .Z(n63361) );
  NOR U78324 ( .A(n60811), .B(n63361), .Z(n58088) );
  XOR U78325 ( .A(n63362), .B(n58088), .Z(n58089) );
  IV U78326 ( .A(n58089), .Z(n60809) );
  XOR U78327 ( .A(n60807), .B(n60809), .Z(n63359) );
  XOR U78328 ( .A(n63360), .B(n63359), .Z(n63372) );
  XOR U78329 ( .A(n63371), .B(n63372), .Z(n60805) );
  XOR U78330 ( .A(n58090), .B(n60805), .Z(n60798) );
  XOR U78331 ( .A(n60799), .B(n60798), .Z(n66250) );
  IV U78332 ( .A(n58091), .Z(n58092) );
  NOR U78333 ( .A(n58093), .B(n58092), .Z(n68740) );
  IV U78334 ( .A(n58094), .Z(n58095) );
  NOR U78335 ( .A(n58096), .B(n58095), .Z(n66249) );
  NOR U78336 ( .A(n68740), .B(n66249), .Z(n60801) );
  XOR U78337 ( .A(n66250), .B(n60801), .Z(n60792) );
  XOR U78338 ( .A(n58097), .B(n60792), .Z(n71173) );
  IV U78339 ( .A(n71173), .Z(n58104) );
  IV U78340 ( .A(n58098), .Z(n58099) );
  NOR U78341 ( .A(n58100), .B(n58099), .Z(n71182) );
  IV U78342 ( .A(n58101), .Z(n58102) );
  NOR U78343 ( .A(n58103), .B(n58102), .Z(n71168) );
  NOR U78344 ( .A(n71182), .B(n71168), .Z(n60790) );
  XOR U78345 ( .A(n58104), .B(n60790), .Z(n60786) );
  XOR U78346 ( .A(n60784), .B(n60786), .Z(n60789) );
  XOR U78347 ( .A(n60787), .B(n60789), .Z(n63383) );
  XOR U78348 ( .A(n63381), .B(n63383), .Z(n68753) );
  XOR U78349 ( .A(n63384), .B(n68753), .Z(n63387) );
  IV U78350 ( .A(n58105), .Z(n58107) );
  NOR U78351 ( .A(n58107), .B(n58106), .Z(n68759) );
  IV U78352 ( .A(n58108), .Z(n58110) );
  NOR U78353 ( .A(n58110), .B(n58109), .Z(n68763) );
  NOR U78354 ( .A(n68759), .B(n68763), .Z(n63388) );
  XOR U78355 ( .A(n63387), .B(n63388), .Z(n63390) );
  XOR U78356 ( .A(n63389), .B(n63390), .Z(n68768) );
  XOR U78357 ( .A(n63394), .B(n68768), .Z(n63395) );
  XOR U78358 ( .A(n63397), .B(n63395), .Z(n63406) );
  IV U78359 ( .A(n58111), .Z(n58113) );
  NOR U78360 ( .A(n58113), .B(n58112), .Z(n63405) );
  IV U78361 ( .A(n58114), .Z(n58116) );
  NOR U78362 ( .A(n58116), .B(n58115), .Z(n63403) );
  NOR U78363 ( .A(n63405), .B(n63403), .Z(n58117) );
  XOR U78364 ( .A(n63406), .B(n58117), .Z(n63400) );
  IV U78365 ( .A(n58118), .Z(n58120) );
  NOR U78366 ( .A(n58120), .B(n58119), .Z(n63401) );
  IV U78367 ( .A(n58121), .Z(n58122) );
  NOR U78368 ( .A(n58122), .B(n58125), .Z(n63414) );
  NOR U78369 ( .A(n63401), .B(n63414), .Z(n58123) );
  XOR U78370 ( .A(n63400), .B(n58123), .Z(n63413) );
  IV U78371 ( .A(n58124), .Z(n58126) );
  NOR U78372 ( .A(n58126), .B(n58125), .Z(n63411) );
  XOR U78373 ( .A(n63413), .B(n63411), .Z(n63419) );
  NOR U78374 ( .A(n58127), .B(n63419), .Z(n66224) );
  IV U78375 ( .A(n58128), .Z(n58133) );
  IV U78376 ( .A(n58129), .Z(n58130) );
  NOR U78377 ( .A(n58133), .B(n58130), .Z(n63421) );
  IV U78378 ( .A(n58131), .Z(n58132) );
  NOR U78379 ( .A(n58133), .B(n58132), .Z(n63418) );
  XOR U78380 ( .A(n63418), .B(n63419), .Z(n63422) );
  XOR U78381 ( .A(n63421), .B(n63422), .Z(n58139) );
  IV U78382 ( .A(n58139), .Z(n58134) );
  NOR U78383 ( .A(n58135), .B(n58134), .Z(n58136) );
  NOR U78384 ( .A(n66224), .B(n58136), .Z(n58137) );
  NOR U78385 ( .A(n58138), .B(n58137), .Z(n58141) );
  IV U78386 ( .A(n58138), .Z(n58140) );
  NOR U78387 ( .A(n58140), .B(n58139), .Z(n68788) );
  NOR U78388 ( .A(n58141), .B(n68788), .Z(n63425) );
  XOR U78389 ( .A(n63427), .B(n63425), .Z(n66218) );
  XOR U78390 ( .A(n63429), .B(n66218), .Z(n60782) );
  XOR U78391 ( .A(n58142), .B(n60782), .Z(n60780) );
  XOR U78392 ( .A(n60778), .B(n60780), .Z(n66204) );
  XOR U78393 ( .A(n60777), .B(n66204), .Z(n58143) );
  IV U78394 ( .A(n58143), .Z(n63438) );
  XOR U78395 ( .A(n63437), .B(n63438), .Z(n66195) );
  XOR U78396 ( .A(n58144), .B(n66195), .Z(n66187) );
  XOR U78397 ( .A(n58145), .B(n66187), .Z(n63455) );
  IV U78398 ( .A(n58146), .Z(n66190) );
  NOR U78399 ( .A(n58147), .B(n66190), .Z(n63450) );
  IV U78400 ( .A(n58148), .Z(n58149) );
  NOR U78401 ( .A(n58150), .B(n58149), .Z(n63454) );
  NOR U78402 ( .A(n63450), .B(n63454), .Z(n58151) );
  XOR U78403 ( .A(n63455), .B(n58151), .Z(n60772) );
  XOR U78404 ( .A(n60773), .B(n60772), .Z(n60775) );
  NOR U78405 ( .A(n58152), .B(n60775), .Z(n68822) );
  IV U78406 ( .A(n58153), .Z(n58154) );
  NOR U78407 ( .A(n58155), .B(n58154), .Z(n58156) );
  IV U78408 ( .A(n58156), .Z(n60776) );
  XOR U78409 ( .A(n60776), .B(n60775), .Z(n58157) );
  NOR U78410 ( .A(n58158), .B(n58157), .Z(n60767) );
  IV U78411 ( .A(n58159), .Z(n58160) );
  NOR U78412 ( .A(n58161), .B(n58160), .Z(n60765) );
  XOR U78413 ( .A(n60767), .B(n60765), .Z(n58162) );
  NOR U78414 ( .A(n68822), .B(n58162), .Z(n60761) );
  NOR U78415 ( .A(n58164), .B(n58163), .Z(n60769) );
  NOR U78416 ( .A(n60769), .B(n60762), .Z(n58165) );
  XOR U78417 ( .A(n60761), .B(n58165), .Z(n63465) );
  XOR U78418 ( .A(n60760), .B(n63465), .Z(n60758) );
  NOR U78419 ( .A(n58171), .B(n60758), .Z(n68833) );
  IV U78420 ( .A(n58166), .Z(n58167) );
  NOR U78421 ( .A(n58168), .B(n58167), .Z(n60757) );
  XOR U78422 ( .A(n60757), .B(n60758), .Z(n63472) );
  IV U78423 ( .A(n58169), .Z(n58170) );
  NOR U78424 ( .A(n58170), .B(n58177), .Z(n58172) );
  IV U78425 ( .A(n58172), .Z(n63471) );
  XOR U78426 ( .A(n63472), .B(n63471), .Z(n58174) );
  NOR U78427 ( .A(n58172), .B(n58171), .Z(n58173) );
  NOR U78428 ( .A(n58174), .B(n58173), .Z(n58175) );
  NOR U78429 ( .A(n68833), .B(n58175), .Z(n60755) );
  IV U78430 ( .A(n58176), .Z(n58178) );
  NOR U78431 ( .A(n58178), .B(n58177), .Z(n60754) );
  IV U78432 ( .A(n58179), .Z(n58180) );
  NOR U78433 ( .A(n58187), .B(n58180), .Z(n63481) );
  NOR U78434 ( .A(n60754), .B(n63481), .Z(n58181) );
  XOR U78435 ( .A(n60755), .B(n58181), .Z(n63480) );
  IV U78436 ( .A(n58182), .Z(n58184) );
  NOR U78437 ( .A(n58184), .B(n58183), .Z(n58185) );
  IV U78438 ( .A(n58185), .Z(n58186) );
  NOR U78439 ( .A(n58187), .B(n58186), .Z(n63478) );
  XOR U78440 ( .A(n63480), .B(n63478), .Z(n63486) );
  XOR U78441 ( .A(n63485), .B(n63486), .Z(n63490) );
  IV U78442 ( .A(n58188), .Z(n58190) );
  IV U78443 ( .A(n58189), .Z(n58204) );
  NOR U78444 ( .A(n58190), .B(n58204), .Z(n58191) );
  IV U78445 ( .A(n58191), .Z(n58197) );
  NOR U78446 ( .A(n63490), .B(n58197), .Z(n68857) );
  IV U78447 ( .A(n58192), .Z(n58193) );
  NOR U78448 ( .A(n58196), .B(n58193), .Z(n63488) );
  XOR U78449 ( .A(n63490), .B(n63488), .Z(n60753) );
  IV U78450 ( .A(n58194), .Z(n58195) );
  NOR U78451 ( .A(n58196), .B(n58195), .Z(n58198) );
  IV U78452 ( .A(n58198), .Z(n60752) );
  XOR U78453 ( .A(n60753), .B(n60752), .Z(n58200) );
  NOR U78454 ( .A(n58198), .B(n58197), .Z(n58199) );
  NOR U78455 ( .A(n58200), .B(n58199), .Z(n58201) );
  NOR U78456 ( .A(n68857), .B(n58201), .Z(n58202) );
  IV U78457 ( .A(n58202), .Z(n63495) );
  IV U78458 ( .A(n58203), .Z(n58205) );
  NOR U78459 ( .A(n58205), .B(n58204), .Z(n63493) );
  XOR U78460 ( .A(n63495), .B(n63493), .Z(n60748) );
  IV U78461 ( .A(n58206), .Z(n58207) );
  NOR U78462 ( .A(n58210), .B(n58207), .Z(n60746) );
  XOR U78463 ( .A(n60748), .B(n60746), .Z(n60751) );
  IV U78464 ( .A(n58208), .Z(n58209) );
  NOR U78465 ( .A(n58210), .B(n58209), .Z(n60749) );
  XOR U78466 ( .A(n60751), .B(n60749), .Z(n63501) );
  IV U78467 ( .A(n58211), .Z(n58213) );
  NOR U78468 ( .A(n58213), .B(n58212), .Z(n60744) );
  IV U78469 ( .A(n58214), .Z(n58216) );
  NOR U78470 ( .A(n58216), .B(n58215), .Z(n63500) );
  NOR U78471 ( .A(n60744), .B(n63500), .Z(n58217) );
  XOR U78472 ( .A(n63501), .B(n58217), .Z(n58218) );
  IV U78473 ( .A(n58218), .Z(n71105) );
  IV U78474 ( .A(n58219), .Z(n58221) );
  NOR U78475 ( .A(n58221), .B(n58220), .Z(n63498) );
  XOR U78476 ( .A(n71105), .B(n63498), .Z(n63505) );
  XOR U78477 ( .A(n60739), .B(n63505), .Z(n63507) );
  XOR U78478 ( .A(n58222), .B(n63507), .Z(n60735) );
  IV U78479 ( .A(n58223), .Z(n58225) );
  NOR U78480 ( .A(n58225), .B(n58224), .Z(n60733) );
  XOR U78481 ( .A(n60735), .B(n60733), .Z(n60738) );
  IV U78482 ( .A(n58226), .Z(n58227) );
  NOR U78483 ( .A(n58230), .B(n58227), .Z(n60736) );
  XOR U78484 ( .A(n60738), .B(n60736), .Z(n60732) );
  IV U78485 ( .A(n58228), .Z(n58229) );
  NOR U78486 ( .A(n58230), .B(n58229), .Z(n60730) );
  XOR U78487 ( .A(n60732), .B(n60730), .Z(n60726) );
  XOR U78488 ( .A(n60725), .B(n60726), .Z(n66150) );
  IV U78489 ( .A(n66150), .Z(n58234) );
  IV U78490 ( .A(n58231), .Z(n58233) );
  NOR U78491 ( .A(n58233), .B(n58232), .Z(n66148) );
  NOR U78492 ( .A(n66153), .B(n66148), .Z(n60728) );
  XOR U78493 ( .A(n58234), .B(n60728), .Z(n60720) );
  XOR U78494 ( .A(n60719), .B(n60720), .Z(n60723) );
  XOR U78495 ( .A(n58235), .B(n60723), .Z(n60712) );
  IV U78496 ( .A(n58236), .Z(n58238) );
  NOR U78497 ( .A(n58238), .B(n58237), .Z(n60716) );
  IV U78498 ( .A(n58239), .Z(n58241) );
  NOR U78499 ( .A(n58241), .B(n58240), .Z(n60711) );
  NOR U78500 ( .A(n60716), .B(n60711), .Z(n58242) );
  XOR U78501 ( .A(n60712), .B(n58242), .Z(n60710) );
  XOR U78502 ( .A(n60708), .B(n60710), .Z(n63518) );
  NOR U78503 ( .A(n58248), .B(n63518), .Z(n66133) );
  IV U78504 ( .A(n58243), .Z(n58244) );
  NOR U78505 ( .A(n58245), .B(n58244), .Z(n60699) );
  IV U78506 ( .A(n58246), .Z(n63519) );
  NOR U78507 ( .A(n63519), .B(n58247), .Z(n60703) );
  XOR U78508 ( .A(n60703), .B(n63518), .Z(n60700) );
  IV U78509 ( .A(n60700), .Z(n58249) );
  XOR U78510 ( .A(n60699), .B(n58249), .Z(n58251) );
  NOR U78511 ( .A(n58249), .B(n58248), .Z(n58250) );
  NOR U78512 ( .A(n58251), .B(n58250), .Z(n58252) );
  NOR U78513 ( .A(n66133), .B(n58252), .Z(n63523) );
  IV U78514 ( .A(n58253), .Z(n58255) );
  NOR U78515 ( .A(n58255), .B(n58254), .Z(n68893) );
  IV U78516 ( .A(n58256), .Z(n58257) );
  NOR U78517 ( .A(n58257), .B(n58260), .Z(n68899) );
  NOR U78518 ( .A(n68893), .B(n68899), .Z(n63524) );
  XOR U78519 ( .A(n63523), .B(n63524), .Z(n63526) );
  NOR U78520 ( .A(n58264), .B(n63526), .Z(n66124) );
  IV U78521 ( .A(n58258), .Z(n58259) );
  NOR U78522 ( .A(n58260), .B(n58259), .Z(n63525) );
  XOR U78523 ( .A(n63525), .B(n63526), .Z(n63536) );
  IV U78524 ( .A(n58261), .Z(n58263) );
  NOR U78525 ( .A(n58263), .B(n58262), .Z(n58265) );
  IV U78526 ( .A(n58265), .Z(n63535) );
  XOR U78527 ( .A(n63536), .B(n63535), .Z(n58267) );
  NOR U78528 ( .A(n58265), .B(n58264), .Z(n58266) );
  NOR U78529 ( .A(n58267), .B(n58266), .Z(n58268) );
  NOR U78530 ( .A(n66124), .B(n58268), .Z(n60691) );
  XOR U78531 ( .A(n58269), .B(n60691), .Z(n60698) );
  IV U78532 ( .A(n58270), .Z(n58278) );
  NOR U78533 ( .A(n58278), .B(n58271), .Z(n60690) );
  IV U78534 ( .A(n58272), .Z(n58274) );
  NOR U78535 ( .A(n58274), .B(n58273), .Z(n60696) );
  NOR U78536 ( .A(n60690), .B(n60696), .Z(n58275) );
  XOR U78537 ( .A(n60698), .B(n58275), .Z(n60687) );
  IV U78538 ( .A(n58276), .Z(n58277) );
  NOR U78539 ( .A(n58278), .B(n58277), .Z(n58279) );
  IV U78540 ( .A(n58279), .Z(n60688) );
  XOR U78541 ( .A(n60687), .B(n60688), .Z(n60685) );
  XOR U78542 ( .A(n58280), .B(n60685), .Z(n60678) );
  XOR U78543 ( .A(n60679), .B(n60678), .Z(n60676) );
  XOR U78544 ( .A(n60672), .B(n60676), .Z(n68916) );
  XOR U78545 ( .A(n58281), .B(n68916), .Z(n63556) );
  IV U78546 ( .A(n58282), .Z(n58284) );
  NOR U78547 ( .A(n58284), .B(n58283), .Z(n63554) );
  XOR U78548 ( .A(n63556), .B(n63554), .Z(n60670) );
  XOR U78549 ( .A(n60669), .B(n60670), .Z(n63563) );
  IV U78550 ( .A(n58285), .Z(n58287) );
  NOR U78551 ( .A(n58287), .B(n58286), .Z(n63561) );
  XOR U78552 ( .A(n63563), .B(n63561), .Z(n63566) );
  IV U78553 ( .A(n58288), .Z(n58289) );
  NOR U78554 ( .A(n58290), .B(n58289), .Z(n63564) );
  XOR U78555 ( .A(n63566), .B(n63564), .Z(n60664) );
  XOR U78556 ( .A(n60663), .B(n60664), .Z(n60657) );
  NOR U78557 ( .A(n58291), .B(n60660), .Z(n58295) );
  IV U78558 ( .A(n58292), .Z(n58294) );
  NOR U78559 ( .A(n58294), .B(n58293), .Z(n60656) );
  NOR U78560 ( .A(n58295), .B(n60656), .Z(n58296) );
  XOR U78561 ( .A(n60657), .B(n58296), .Z(n68922) );
  IV U78562 ( .A(n58297), .Z(n58301) );
  NOR U78563 ( .A(n58299), .B(n58298), .Z(n58300) );
  IV U78564 ( .A(n58300), .Z(n58303) );
  NOR U78565 ( .A(n58301), .B(n58303), .Z(n63570) );
  IV U78566 ( .A(n58302), .Z(n58304) );
  NOR U78567 ( .A(n58304), .B(n58303), .Z(n60655) );
  NOR U78568 ( .A(n63570), .B(n60655), .Z(n58305) );
  XOR U78569 ( .A(n68922), .B(n58305), .Z(n63577) );
  IV U78570 ( .A(n63577), .Z(n58310) );
  IV U78571 ( .A(n58306), .Z(n58307) );
  NOR U78572 ( .A(n58308), .B(n58307), .Z(n63572) );
  NOR U78573 ( .A(n63572), .B(n63576), .Z(n58309) );
  XOR U78574 ( .A(n58310), .B(n58309), .Z(n63584) );
  XOR U78575 ( .A(n63582), .B(n63584), .Z(n60652) );
  XOR U78576 ( .A(n60651), .B(n60652), .Z(n63580) );
  XOR U78577 ( .A(n63579), .B(n63580), .Z(n60648) );
  XOR U78578 ( .A(n58311), .B(n60648), .Z(n60645) );
  XOR U78579 ( .A(n60644), .B(n60645), .Z(n66077) );
  XOR U78580 ( .A(n63593), .B(n66077), .Z(n63594) );
  XOR U78581 ( .A(n63595), .B(n63594), .Z(n63600) );
  IV U78582 ( .A(n58312), .Z(n58313) );
  NOR U78583 ( .A(n58313), .B(n58316), .Z(n63598) );
  XOR U78584 ( .A(n63600), .B(n63598), .Z(n63603) );
  IV U78585 ( .A(n58314), .Z(n58315) );
  NOR U78586 ( .A(n58316), .B(n58315), .Z(n63601) );
  XOR U78587 ( .A(n63603), .B(n63601), .Z(n66054) );
  XOR U78588 ( .A(n60641), .B(n66054), .Z(n60636) );
  XOR U78589 ( .A(n60637), .B(n60636), .Z(n60639) );
  XOR U78590 ( .A(n60638), .B(n60639), .Z(n63612) );
  IV U78591 ( .A(n58317), .Z(n58319) );
  NOR U78592 ( .A(n58319), .B(n58318), .Z(n63610) );
  XOR U78593 ( .A(n63612), .B(n63610), .Z(n63625) );
  NOR U78594 ( .A(n60634), .B(n63624), .Z(n58320) );
  XOR U78595 ( .A(n63625), .B(n58320), .Z(n63621) );
  IV U78596 ( .A(n58321), .Z(n58324) );
  IV U78597 ( .A(n58322), .Z(n58323) );
  NOR U78598 ( .A(n58324), .B(n58323), .Z(n58325) );
  IV U78599 ( .A(n58325), .Z(n63622) );
  XOR U78600 ( .A(n63621), .B(n63622), .Z(n60630) );
  XOR U78601 ( .A(n60628), .B(n60630), .Z(n60632) );
  XOR U78602 ( .A(n60631), .B(n60632), .Z(n63630) );
  XOR U78603 ( .A(n58326), .B(n63630), .Z(n63634) );
  IV U78604 ( .A(n58327), .Z(n58328) );
  NOR U78605 ( .A(n58329), .B(n58328), .Z(n63632) );
  XOR U78606 ( .A(n63634), .B(n63632), .Z(n90897) );
  NOR U78607 ( .A(n58331), .B(n58330), .Z(n90898) );
  NOR U78608 ( .A(n90898), .B(n63646), .Z(n58332) );
  XOR U78609 ( .A(n90897), .B(n58332), .Z(n60623) );
  XOR U78610 ( .A(n60624), .B(n60623), .Z(n60619) );
  IV U78611 ( .A(n58333), .Z(n58335) );
  NOR U78612 ( .A(n58335), .B(n58334), .Z(n60617) );
  XOR U78613 ( .A(n60619), .B(n60617), .Z(n60622) );
  IV U78614 ( .A(n58336), .Z(n58337) );
  NOR U78615 ( .A(n58340), .B(n58337), .Z(n60620) );
  XOR U78616 ( .A(n60622), .B(n60620), .Z(n66019) );
  IV U78617 ( .A(n58338), .Z(n58339) );
  NOR U78618 ( .A(n58340), .B(n58339), .Z(n66023) );
  IV U78619 ( .A(n58341), .Z(n58343) );
  NOR U78620 ( .A(n58343), .B(n58342), .Z(n66018) );
  NOR U78621 ( .A(n66023), .B(n66018), .Z(n60613) );
  XOR U78622 ( .A(n66019), .B(n60613), .Z(n58344) );
  IV U78623 ( .A(n58344), .Z(n60616) );
  XOR U78624 ( .A(n60614), .B(n60616), .Z(n63657) );
  XOR U78625 ( .A(n58345), .B(n63657), .Z(n60608) );
  XOR U78626 ( .A(n58346), .B(n60608), .Z(n60604) );
  XOR U78627 ( .A(n60602), .B(n60604), .Z(n60606) );
  NOR U78628 ( .A(n58353), .B(n60606), .Z(n60601) );
  IV U78629 ( .A(n58347), .Z(n58348) );
  NOR U78630 ( .A(n58349), .B(n58348), .Z(n60598) );
  IV U78631 ( .A(n58350), .Z(n58352) );
  NOR U78632 ( .A(n58352), .B(n58351), .Z(n60605) );
  XOR U78633 ( .A(n60605), .B(n60606), .Z(n60599) );
  IV U78634 ( .A(n60599), .Z(n58354) );
  XOR U78635 ( .A(n60598), .B(n58354), .Z(n58356) );
  NOR U78636 ( .A(n58354), .B(n58353), .Z(n58355) );
  NOR U78637 ( .A(n58356), .B(n58355), .Z(n58357) );
  NOR U78638 ( .A(n60601), .B(n58357), .Z(n58358) );
  IV U78639 ( .A(n58358), .Z(n63677) );
  IV U78640 ( .A(n58359), .Z(n58361) );
  NOR U78641 ( .A(n58361), .B(n58360), .Z(n63676) );
  XOR U78642 ( .A(n63677), .B(n63676), .Z(n63680) );
  XOR U78643 ( .A(n58362), .B(n63680), .Z(n60591) );
  XOR U78644 ( .A(n60590), .B(n60591), .Z(n60594) );
  XOR U78645 ( .A(n60593), .B(n60594), .Z(n63687) );
  IV U78646 ( .A(n58363), .Z(n58364) );
  NOR U78647 ( .A(n58365), .B(n58364), .Z(n63685) );
  XOR U78648 ( .A(n63687), .B(n63685), .Z(n63690) );
  IV U78649 ( .A(n58366), .Z(n58367) );
  NOR U78650 ( .A(n58367), .B(n58372), .Z(n63688) );
  XOR U78651 ( .A(n63690), .B(n63688), .Z(n60585) );
  XOR U78652 ( .A(n60584), .B(n60585), .Z(n60589) );
  IV U78653 ( .A(n60589), .Z(n58375) );
  IV U78654 ( .A(n58368), .Z(n58369) );
  NOR U78655 ( .A(n58370), .B(n58369), .Z(n60582) );
  IV U78656 ( .A(n58371), .Z(n58373) );
  NOR U78657 ( .A(n58373), .B(n58372), .Z(n60587) );
  NOR U78658 ( .A(n60582), .B(n60587), .Z(n58374) );
  XOR U78659 ( .A(n58375), .B(n58374), .Z(n63695) );
  XOR U78660 ( .A(n63692), .B(n63695), .Z(n65987) );
  XOR U78661 ( .A(n58376), .B(n65987), .Z(n60578) );
  XOR U78662 ( .A(n58377), .B(n60578), .Z(n60577) );
  XOR U78663 ( .A(n60575), .B(n60577), .Z(n63703) );
  XOR U78664 ( .A(n63701), .B(n63703), .Z(n63706) );
  IV U78665 ( .A(n58378), .Z(n58386) );
  IV U78666 ( .A(n58379), .Z(n58380) );
  NOR U78667 ( .A(n58386), .B(n58380), .Z(n58381) );
  IV U78668 ( .A(n58381), .Z(n58400) );
  NOR U78669 ( .A(n63706), .B(n58400), .Z(n65966) );
  IV U78670 ( .A(n58382), .Z(n58383) );
  NOR U78671 ( .A(n58383), .B(n58388), .Z(n69010) );
  IV U78672 ( .A(n58384), .Z(n58385) );
  NOR U78673 ( .A(n58386), .B(n58385), .Z(n65969) );
  NOR U78674 ( .A(n69010), .B(n65969), .Z(n60574) );
  IV U78675 ( .A(n58387), .Z(n58389) );
  NOR U78676 ( .A(n58389), .B(n58388), .Z(n63704) );
  XOR U78677 ( .A(n63704), .B(n63706), .Z(n65971) );
  XOR U78678 ( .A(n60574), .B(n65971), .Z(n58390) );
  IV U78679 ( .A(n58390), .Z(n60572) );
  IV U78680 ( .A(n58391), .Z(n58392) );
  NOR U78681 ( .A(n58393), .B(n58392), .Z(n58394) );
  IV U78682 ( .A(n58394), .Z(n58399) );
  NOR U78683 ( .A(n58396), .B(n58395), .Z(n58397) );
  IV U78684 ( .A(n58397), .Z(n58398) );
  NOR U78685 ( .A(n58399), .B(n58398), .Z(n58401) );
  IV U78686 ( .A(n58401), .Z(n60571) );
  XOR U78687 ( .A(n60572), .B(n60571), .Z(n58403) );
  NOR U78688 ( .A(n58401), .B(n58400), .Z(n58402) );
  NOR U78689 ( .A(n58403), .B(n58402), .Z(n58404) );
  NOR U78690 ( .A(n65966), .B(n58404), .Z(n60569) );
  XOR U78691 ( .A(n58405), .B(n60569), .Z(n63713) );
  IV U78692 ( .A(n58406), .Z(n58407) );
  NOR U78693 ( .A(n58408), .B(n58407), .Z(n63712) );
  XOR U78694 ( .A(n63713), .B(n63712), .Z(n63717) );
  IV U78695 ( .A(n58409), .Z(n58414) );
  IV U78696 ( .A(n58410), .Z(n58411) );
  NOR U78697 ( .A(n58414), .B(n58411), .Z(n63715) );
  XOR U78698 ( .A(n63717), .B(n63715), .Z(n63720) );
  IV U78699 ( .A(n58412), .Z(n58413) );
  NOR U78700 ( .A(n58414), .B(n58413), .Z(n63718) );
  XOR U78701 ( .A(n63720), .B(n63718), .Z(n60567) );
  IV U78702 ( .A(n58415), .Z(n58416) );
  NOR U78703 ( .A(n58417), .B(n58416), .Z(n60566) );
  NOR U78704 ( .A(n58418), .B(n60563), .Z(n58419) );
  NOR U78705 ( .A(n60566), .B(n58419), .Z(n58420) );
  XOR U78706 ( .A(n60567), .B(n58420), .Z(n60558) );
  IV U78707 ( .A(n58421), .Z(n58423) );
  NOR U78708 ( .A(n58423), .B(n58422), .Z(n58424) );
  IV U78709 ( .A(n58424), .Z(n60559) );
  XOR U78710 ( .A(n60558), .B(n60559), .Z(n65941) );
  XOR U78711 ( .A(n63731), .B(n65941), .Z(n58425) );
  IV U78712 ( .A(n58425), .Z(n63734) );
  IV U78713 ( .A(n58426), .Z(n58428) );
  NOR U78714 ( .A(n58428), .B(n58427), .Z(n63732) );
  XOR U78715 ( .A(n63734), .B(n63732), .Z(n60556) );
  IV U78716 ( .A(n60556), .Z(n58436) );
  IV U78717 ( .A(n58429), .Z(n58431) );
  NOR U78718 ( .A(n58431), .B(n58430), .Z(n60555) );
  IV U78719 ( .A(n58432), .Z(n58433) );
  NOR U78720 ( .A(n58434), .B(n58433), .Z(n60553) );
  NOR U78721 ( .A(n60555), .B(n60553), .Z(n58435) );
  XOR U78722 ( .A(n58436), .B(n58435), .Z(n65932) );
  XOR U78723 ( .A(n63739), .B(n65932), .Z(n63738) );
  XOR U78724 ( .A(n58437), .B(n63738), .Z(n63750) );
  XOR U78725 ( .A(n58438), .B(n63750), .Z(n58446) );
  IV U78726 ( .A(n58446), .Z(n58439) );
  NOR U78727 ( .A(n58440), .B(n58439), .Z(n69030) );
  IV U78728 ( .A(n58441), .Z(n58443) );
  NOR U78729 ( .A(n58443), .B(n58442), .Z(n58447) );
  IV U78730 ( .A(n58447), .Z(n58445) );
  XOR U78731 ( .A(n63750), .B(n63746), .Z(n58444) );
  NOR U78732 ( .A(n58445), .B(n58444), .Z(n65920) );
  NOR U78733 ( .A(n58447), .B(n58446), .Z(n58448) );
  NOR U78734 ( .A(n65920), .B(n58448), .Z(n58449) );
  NOR U78735 ( .A(n58450), .B(n58449), .Z(n58451) );
  NOR U78736 ( .A(n69030), .B(n58451), .Z(n58452) );
  IV U78737 ( .A(n58452), .Z(n63754) );
  IV U78738 ( .A(n58453), .Z(n58455) );
  NOR U78739 ( .A(n58455), .B(n58454), .Z(n63752) );
  XOR U78740 ( .A(n63754), .B(n63752), .Z(n63757) );
  XOR U78741 ( .A(n63755), .B(n63757), .Z(n63760) );
  IV U78742 ( .A(n58456), .Z(n58458) );
  NOR U78743 ( .A(n58458), .B(n58457), .Z(n58459) );
  IV U78744 ( .A(n58459), .Z(n58465) );
  NOR U78745 ( .A(n63760), .B(n58465), .Z(n65906) );
  IV U78746 ( .A(n58460), .Z(n58461) );
  NOR U78747 ( .A(n58464), .B(n58461), .Z(n63762) );
  IV U78748 ( .A(n58462), .Z(n58463) );
  NOR U78749 ( .A(n58464), .B(n58463), .Z(n63759) );
  XOR U78750 ( .A(n63759), .B(n63760), .Z(n63763) );
  IV U78751 ( .A(n63763), .Z(n58466) );
  XOR U78752 ( .A(n63762), .B(n58466), .Z(n58468) );
  NOR U78753 ( .A(n58466), .B(n58465), .Z(n58467) );
  NOR U78754 ( .A(n58468), .B(n58467), .Z(n58469) );
  NOR U78755 ( .A(n65906), .B(n58469), .Z(n58470) );
  IV U78756 ( .A(n58470), .Z(n63767) );
  XOR U78757 ( .A(n63766), .B(n63767), .Z(n63770) );
  IV U78758 ( .A(n63770), .Z(n58477) );
  IV U78759 ( .A(n58471), .Z(n58472) );
  NOR U78760 ( .A(n58473), .B(n58472), .Z(n63769) );
  IV U78761 ( .A(n58474), .Z(n58475) );
  NOR U78762 ( .A(n58475), .B(n58478), .Z(n60551) );
  NOR U78763 ( .A(n63769), .B(n60551), .Z(n58476) );
  XOR U78764 ( .A(n58477), .B(n58476), .Z(n60550) );
  NOR U78765 ( .A(n58479), .B(n58478), .Z(n58480) );
  IV U78766 ( .A(n58480), .Z(n58481) );
  NOR U78767 ( .A(n58482), .B(n58481), .Z(n60548) );
  XOR U78768 ( .A(n60550), .B(n60548), .Z(n60544) );
  XOR U78769 ( .A(n60542), .B(n60544), .Z(n60547) );
  XOR U78770 ( .A(n58483), .B(n60547), .Z(n60539) );
  IV U78771 ( .A(n58484), .Z(n58488) );
  NOR U78772 ( .A(n58486), .B(n58485), .Z(n58487) );
  IV U78773 ( .A(n58487), .Z(n58491) );
  NOR U78774 ( .A(n58488), .B(n58491), .Z(n58489) );
  IV U78775 ( .A(n58489), .Z(n60540) );
  XOR U78776 ( .A(n60539), .B(n60540), .Z(n63778) );
  IV U78777 ( .A(n58490), .Z(n58492) );
  NOR U78778 ( .A(n58492), .B(n58491), .Z(n63776) );
  XOR U78779 ( .A(n63778), .B(n63776), .Z(n63781) );
  IV U78780 ( .A(n58493), .Z(n58494) );
  NOR U78781 ( .A(n58495), .B(n58494), .Z(n63779) );
  XOR U78782 ( .A(n63781), .B(n63779), .Z(n60532) );
  XOR U78783 ( .A(n60531), .B(n60532), .Z(n60535) );
  XOR U78784 ( .A(n60534), .B(n60535), .Z(n60530) );
  IV U78785 ( .A(n58496), .Z(n58498) );
  NOR U78786 ( .A(n58498), .B(n58497), .Z(n60523) );
  IV U78787 ( .A(n58499), .Z(n58501) );
  NOR U78788 ( .A(n58501), .B(n58500), .Z(n60528) );
  NOR U78789 ( .A(n60523), .B(n60528), .Z(n58502) );
  XOR U78790 ( .A(n60530), .B(n58502), .Z(n58508) );
  XOR U78791 ( .A(n60525), .B(n58508), .Z(n58514) );
  IV U78792 ( .A(n58514), .Z(n58503) );
  NOR U78793 ( .A(n58504), .B(n58503), .Z(n65879) );
  IV U78794 ( .A(n58505), .Z(n58507) );
  NOR U78795 ( .A(n58507), .B(n58506), .Z(n58511) );
  IV U78796 ( .A(n58511), .Z(n58509) );
  IV U78797 ( .A(n58508), .Z(n60526) );
  NOR U78798 ( .A(n58509), .B(n60526), .Z(n65876) );
  NOR U78799 ( .A(n58511), .B(n58510), .Z(n58512) );
  IV U78800 ( .A(n58512), .Z(n58513) );
  NOR U78801 ( .A(n58514), .B(n58513), .Z(n58515) );
  NOR U78802 ( .A(n65876), .B(n58515), .Z(n58516) );
  IV U78803 ( .A(n58516), .Z(n60520) );
  NOR U78804 ( .A(n65879), .B(n60520), .Z(n63787) );
  IV U78805 ( .A(n58517), .Z(n65873) );
  NOR U78806 ( .A(n65873), .B(n65875), .Z(n60519) );
  IV U78807 ( .A(n58518), .Z(n58520) );
  NOR U78808 ( .A(n58520), .B(n58519), .Z(n63786) );
  NOR U78809 ( .A(n60519), .B(n63786), .Z(n58521) );
  XOR U78810 ( .A(n63787), .B(n58521), .Z(n65860) );
  XOR U78811 ( .A(n58522), .B(n65860), .Z(n60511) );
  XOR U78812 ( .A(n58523), .B(n60511), .Z(n60509) );
  XOR U78813 ( .A(n58524), .B(n60509), .Z(n60504) );
  XOR U78814 ( .A(n58525), .B(n60504), .Z(n60493) );
  IV U78815 ( .A(n58526), .Z(n58528) );
  NOR U78816 ( .A(n58528), .B(n58527), .Z(n60497) );
  IV U78817 ( .A(n58529), .Z(n58531) );
  NOR U78818 ( .A(n58531), .B(n58530), .Z(n60494) );
  NOR U78819 ( .A(n60497), .B(n60494), .Z(n58532) );
  XOR U78820 ( .A(n60493), .B(n58532), .Z(n60492) );
  XOR U78821 ( .A(n60490), .B(n60492), .Z(n65837) );
  XOR U78822 ( .A(n60489), .B(n65837), .Z(n58533) );
  IV U78823 ( .A(n58533), .Z(n60484) );
  XOR U78824 ( .A(n65836), .B(n60484), .Z(n60487) );
  XOR U78825 ( .A(n60486), .B(n60487), .Z(n60482) );
  XOR U78826 ( .A(n60481), .B(n60482), .Z(n65833) );
  XOR U78827 ( .A(n63800), .B(n65833), .Z(n60478) );
  XOR U78828 ( .A(n58534), .B(n60478), .Z(n65826) );
  XOR U78829 ( .A(n60476), .B(n65826), .Z(n60474) );
  XOR U78830 ( .A(n58535), .B(n60474), .Z(n63812) );
  XOR U78831 ( .A(n63810), .B(n63812), .Z(n63815) );
  IV U78832 ( .A(n58536), .Z(n58542) );
  XOR U78833 ( .A(n58537), .B(n58544), .Z(n58538) );
  NOR U78834 ( .A(n58539), .B(n58538), .Z(n58540) );
  IV U78835 ( .A(n58540), .Z(n58541) );
  NOR U78836 ( .A(n58542), .B(n58541), .Z(n60471) );
  IV U78837 ( .A(n58543), .Z(n58548) );
  NOR U78838 ( .A(n58545), .B(n58544), .Z(n58546) );
  IV U78839 ( .A(n58546), .Z(n58547) );
  NOR U78840 ( .A(n58548), .B(n58547), .Z(n63813) );
  NOR U78841 ( .A(n60471), .B(n63813), .Z(n58549) );
  XOR U78842 ( .A(n63815), .B(n58549), .Z(n60468) );
  IV U78843 ( .A(n58550), .Z(n58551) );
  NOR U78844 ( .A(n58554), .B(n58551), .Z(n60469) );
  IV U78845 ( .A(n58552), .Z(n58553) );
  NOR U78846 ( .A(n58554), .B(n58553), .Z(n63818) );
  NOR U78847 ( .A(n60469), .B(n63818), .Z(n58555) );
  XOR U78848 ( .A(n60468), .B(n58555), .Z(n63822) );
  XOR U78849 ( .A(n63821), .B(n63822), .Z(n63827) );
  XOR U78850 ( .A(n60464), .B(n63827), .Z(n63830) );
  NOR U78851 ( .A(n58556), .B(n58561), .Z(n60466) );
  IV U78852 ( .A(n58557), .Z(n58558) );
  NOR U78853 ( .A(n58559), .B(n58558), .Z(n63828) );
  IV U78854 ( .A(n58560), .Z(n58562) );
  NOR U78855 ( .A(n58562), .B(n58561), .Z(n63825) );
  NOR U78856 ( .A(n63828), .B(n63825), .Z(n58563) );
  IV U78857 ( .A(n58563), .Z(n58564) );
  NOR U78858 ( .A(n60466), .B(n58564), .Z(n58565) );
  XOR U78859 ( .A(n63830), .B(n58565), .Z(n60461) );
  IV U78860 ( .A(n58566), .Z(n58567) );
  NOR U78861 ( .A(n58568), .B(n58567), .Z(n60462) );
  IV U78862 ( .A(n58569), .Z(n58571) );
  NOR U78863 ( .A(n58571), .B(n58570), .Z(n63831) );
  NOR U78864 ( .A(n60462), .B(n63831), .Z(n58572) );
  XOR U78865 ( .A(n60461), .B(n58572), .Z(n60456) );
  XOR U78866 ( .A(n60455), .B(n60456), .Z(n60459) );
  IV U78867 ( .A(n58573), .Z(n58575) );
  NOR U78868 ( .A(n58575), .B(n58574), .Z(n60458) );
  IV U78869 ( .A(n58576), .Z(n58583) );
  NOR U78870 ( .A(n58578), .B(n58577), .Z(n58579) );
  IV U78871 ( .A(n58579), .Z(n58580) );
  NOR U78872 ( .A(n58581), .B(n58580), .Z(n58582) );
  IV U78873 ( .A(n58582), .Z(n58587) );
  NOR U78874 ( .A(n58583), .B(n58587), .Z(n60453) );
  NOR U78875 ( .A(n60458), .B(n60453), .Z(n58584) );
  XOR U78876 ( .A(n60459), .B(n58584), .Z(n58585) );
  IV U78877 ( .A(n58585), .Z(n60452) );
  IV U78878 ( .A(n58586), .Z(n58588) );
  NOR U78879 ( .A(n58588), .B(n58587), .Z(n60450) );
  XOR U78880 ( .A(n60452), .B(n60450), .Z(n58590) );
  NOR U78881 ( .A(n58595), .B(n58590), .Z(n69115) );
  NOR U78882 ( .A(n58589), .B(n60444), .Z(n58591) );
  XOR U78883 ( .A(n58591), .B(n58590), .Z(n60439) );
  IV U78884 ( .A(n58592), .Z(n58594) );
  NOR U78885 ( .A(n58594), .B(n58593), .Z(n58596) );
  IV U78886 ( .A(n58596), .Z(n60438) );
  XOR U78887 ( .A(n60439), .B(n60438), .Z(n58598) );
  NOR U78888 ( .A(n58596), .B(n58595), .Z(n58597) );
  NOR U78889 ( .A(n58598), .B(n58597), .Z(n58599) );
  NOR U78890 ( .A(n69115), .B(n58599), .Z(n60441) );
  XOR U78891 ( .A(n58600), .B(n60441), .Z(n63843) );
  XOR U78892 ( .A(n58601), .B(n63843), .Z(n60436) );
  XOR U78893 ( .A(n60435), .B(n60436), .Z(n60431) );
  XOR U78894 ( .A(n60429), .B(n60431), .Z(n60434) );
  XOR U78895 ( .A(n60432), .B(n60434), .Z(n60427) );
  NOR U78896 ( .A(n58608), .B(n60427), .Z(n65786) );
  IV U78897 ( .A(n58602), .Z(n58604) );
  NOR U78898 ( .A(n58604), .B(n58603), .Z(n60423) );
  IV U78899 ( .A(n58605), .Z(n58606) );
  NOR U78900 ( .A(n58607), .B(n58606), .Z(n60426) );
  XOR U78901 ( .A(n60426), .B(n60427), .Z(n60424) );
  IV U78902 ( .A(n60424), .Z(n58609) );
  XOR U78903 ( .A(n60423), .B(n58609), .Z(n58611) );
  NOR U78904 ( .A(n58609), .B(n58608), .Z(n58610) );
  NOR U78905 ( .A(n58611), .B(n58610), .Z(n58612) );
  NOR U78906 ( .A(n65786), .B(n58612), .Z(n58613) );
  IV U78907 ( .A(n58613), .Z(n63848) );
  IV U78908 ( .A(n58614), .Z(n58616) );
  NOR U78909 ( .A(n58616), .B(n58615), .Z(n63846) );
  XOR U78910 ( .A(n63848), .B(n63846), .Z(n63851) );
  XOR U78911 ( .A(n63849), .B(n63851), .Z(n63854) );
  NOR U78912 ( .A(n58623), .B(n63854), .Z(n74199) );
  IV U78913 ( .A(n58617), .Z(n58619) );
  NOR U78914 ( .A(n58619), .B(n58618), .Z(n63856) );
  IV U78915 ( .A(n58620), .Z(n58621) );
  NOR U78916 ( .A(n58622), .B(n58621), .Z(n63853) );
  XOR U78917 ( .A(n63853), .B(n63854), .Z(n63857) );
  IV U78918 ( .A(n63857), .Z(n58624) );
  XOR U78919 ( .A(n63856), .B(n58624), .Z(n58626) );
  NOR U78920 ( .A(n58624), .B(n58623), .Z(n58625) );
  NOR U78921 ( .A(n58626), .B(n58625), .Z(n58627) );
  NOR U78922 ( .A(n74199), .B(n58627), .Z(n63859) );
  XOR U78923 ( .A(n63860), .B(n63859), .Z(n60419) );
  XOR U78924 ( .A(n60417), .B(n60419), .Z(n60421) );
  XOR U78925 ( .A(n60420), .B(n60421), .Z(n74230) );
  XOR U78926 ( .A(n60416), .B(n74230), .Z(n63864) );
  IV U78927 ( .A(n58628), .Z(n58630) );
  NOR U78928 ( .A(n58630), .B(n58629), .Z(n58631) );
  IV U78929 ( .A(n58631), .Z(n63865) );
  XOR U78930 ( .A(n63864), .B(n63865), .Z(n63872) );
  IV U78931 ( .A(n58632), .Z(n58633) );
  NOR U78932 ( .A(n58634), .B(n58633), .Z(n63867) );
  IV U78933 ( .A(n58635), .Z(n58637) );
  NOR U78934 ( .A(n58637), .B(n58636), .Z(n63871) );
  NOR U78935 ( .A(n63867), .B(n63871), .Z(n58638) );
  XOR U78936 ( .A(n63872), .B(n58638), .Z(n60410) );
  XOR U78937 ( .A(n60411), .B(n60410), .Z(n60414) );
  XOR U78938 ( .A(n60413), .B(n60414), .Z(n60407) );
  XOR U78939 ( .A(n58639), .B(n60407), .Z(n58640) );
  IV U78940 ( .A(n58640), .Z(n60402) );
  IV U78941 ( .A(n58641), .Z(n58642) );
  NOR U78942 ( .A(n58642), .B(n58645), .Z(n60401) );
  IV U78943 ( .A(n58643), .Z(n58644) );
  NOR U78944 ( .A(n58645), .B(n58644), .Z(n60399) );
  NOR U78945 ( .A(n60401), .B(n60399), .Z(n58646) );
  XOR U78946 ( .A(n60402), .B(n58646), .Z(n60393) );
  IV U78947 ( .A(n58647), .Z(n58648) );
  NOR U78948 ( .A(n58649), .B(n58648), .Z(n60396) );
  IV U78949 ( .A(n58650), .Z(n58651) );
  NOR U78950 ( .A(n58655), .B(n58651), .Z(n60394) );
  NOR U78951 ( .A(n60396), .B(n60394), .Z(n58652) );
  XOR U78952 ( .A(n60393), .B(n58652), .Z(n60392) );
  IV U78953 ( .A(n58653), .Z(n58654) );
  NOR U78954 ( .A(n58655), .B(n58654), .Z(n60390) );
  XOR U78955 ( .A(n60392), .B(n60390), .Z(n63878) );
  XOR U78956 ( .A(n63877), .B(n63878), .Z(n63881) );
  XOR U78957 ( .A(n63880), .B(n63881), .Z(n63890) );
  IV U78958 ( .A(n58656), .Z(n58658) );
  NOR U78959 ( .A(n58658), .B(n58657), .Z(n63875) );
  IV U78960 ( .A(n58659), .Z(n58661) );
  NOR U78961 ( .A(n58661), .B(n58660), .Z(n63889) );
  NOR U78962 ( .A(n63875), .B(n63889), .Z(n58662) );
  XOR U78963 ( .A(n63890), .B(n58662), .Z(n58663) );
  IV U78964 ( .A(n58663), .Z(n63888) );
  IV U78965 ( .A(n58664), .Z(n58665) );
  NOR U78966 ( .A(n58666), .B(n58665), .Z(n58667) );
  IV U78967 ( .A(n58667), .Z(n58674) );
  NOR U78968 ( .A(n63888), .B(n58674), .Z(n65733) );
  IV U78969 ( .A(n58668), .Z(n58670) );
  NOR U78970 ( .A(n58670), .B(n58669), .Z(n63886) );
  XOR U78971 ( .A(n63886), .B(n63888), .Z(n63894) );
  IV U78972 ( .A(n58671), .Z(n58672) );
  NOR U78973 ( .A(n58673), .B(n58672), .Z(n58675) );
  IV U78974 ( .A(n58675), .Z(n63893) );
  XOR U78975 ( .A(n63894), .B(n63893), .Z(n58677) );
  NOR U78976 ( .A(n58675), .B(n58674), .Z(n58676) );
  NOR U78977 ( .A(n58677), .B(n58676), .Z(n65731) );
  NOR U78978 ( .A(n65733), .B(n65731), .Z(n60387) );
  XOR U78979 ( .A(n58678), .B(n60387), .Z(n63901) );
  XOR U78980 ( .A(n63899), .B(n63901), .Z(n63904) );
  IV U78981 ( .A(n58679), .Z(n58681) );
  NOR U78982 ( .A(n58681), .B(n58680), .Z(n63902) );
  XOR U78983 ( .A(n63904), .B(n63902), .Z(n60384) );
  IV U78984 ( .A(n58682), .Z(n58684) );
  NOR U78985 ( .A(n58684), .B(n58683), .Z(n60383) );
  IV U78986 ( .A(n58685), .Z(n58686) );
  NOR U78987 ( .A(n58687), .B(n58686), .Z(n60381) );
  NOR U78988 ( .A(n60383), .B(n60381), .Z(n58688) );
  XOR U78989 ( .A(n60384), .B(n58688), .Z(n63912) );
  XOR U78990 ( .A(n63914), .B(n63912), .Z(n63917) );
  XOR U78991 ( .A(n63915), .B(n63917), .Z(n60380) );
  XOR U78992 ( .A(n60378), .B(n60380), .Z(n58689) );
  NOR U78993 ( .A(n58690), .B(n58689), .Z(n65711) );
  NOR U78994 ( .A(n58691), .B(n60370), .Z(n58692) );
  NOR U78995 ( .A(n58692), .B(n60378), .Z(n58693) );
  XOR U78996 ( .A(n58693), .B(n60380), .Z(n58703) );
  NOR U78997 ( .A(n58694), .B(n58703), .Z(n58695) );
  NOR U78998 ( .A(n65711), .B(n58695), .Z(n58706) );
  IV U78999 ( .A(n58706), .Z(n58696) );
  NOR U79000 ( .A(n58709), .B(n58696), .Z(n65704) );
  IV U79001 ( .A(n58697), .Z(n58699) );
  NOR U79002 ( .A(n58699), .B(n58698), .Z(n60362) );
  IV U79003 ( .A(n58700), .Z(n58702) );
  NOR U79004 ( .A(n58702), .B(n58701), .Z(n58707) );
  IV U79005 ( .A(n58707), .Z(n58705) );
  IV U79006 ( .A(n58703), .Z(n58704) );
  NOR U79007 ( .A(n58705), .B(n58704), .Z(n65709) );
  NOR U79008 ( .A(n58707), .B(n58706), .Z(n58708) );
  NOR U79009 ( .A(n65709), .B(n58708), .Z(n60363) );
  XOR U79010 ( .A(n60362), .B(n60363), .Z(n58711) );
  NOR U79011 ( .A(n60363), .B(n58709), .Z(n58710) );
  NOR U79012 ( .A(n58711), .B(n58710), .Z(n58712) );
  NOR U79013 ( .A(n65704), .B(n58712), .Z(n58713) );
  IV U79014 ( .A(n58713), .Z(n60367) );
  XOR U79015 ( .A(n60366), .B(n60367), .Z(n63925) );
  IV U79016 ( .A(n58714), .Z(n58715) );
  NOR U79017 ( .A(n58716), .B(n58715), .Z(n63923) );
  XOR U79018 ( .A(n63925), .B(n63923), .Z(n63928) );
  IV U79019 ( .A(n58717), .Z(n58718) );
  NOR U79020 ( .A(n58719), .B(n58718), .Z(n60360) );
  IV U79021 ( .A(n58720), .Z(n58721) );
  NOR U79022 ( .A(n58722), .B(n58721), .Z(n63926) );
  NOR U79023 ( .A(n60360), .B(n63926), .Z(n58723) );
  XOR U79024 ( .A(n63928), .B(n58723), .Z(n60353) );
  XOR U79025 ( .A(n58724), .B(n60353), .Z(n63947) );
  XOR U79026 ( .A(n58725), .B(n63947), .Z(n60350) );
  XOR U79027 ( .A(n60351), .B(n60350), .Z(n60347) );
  IV U79028 ( .A(n58726), .Z(n58728) );
  NOR U79029 ( .A(n58728), .B(n58727), .Z(n60345) );
  XOR U79030 ( .A(n60347), .B(n60345), .Z(n63965) );
  XOR U79031 ( .A(n58729), .B(n63965), .Z(n60344) );
  IV U79032 ( .A(n58730), .Z(n58731) );
  NOR U79033 ( .A(n58732), .B(n58731), .Z(n63964) );
  IV U79034 ( .A(n58733), .Z(n58737) );
  NOR U79035 ( .A(n58735), .B(n58734), .Z(n58736) );
  IV U79036 ( .A(n58736), .Z(n58741) );
  NOR U79037 ( .A(n58737), .B(n58741), .Z(n60342) );
  NOR U79038 ( .A(n63964), .B(n60342), .Z(n58738) );
  XOR U79039 ( .A(n60344), .B(n58738), .Z(n58739) );
  IV U79040 ( .A(n58739), .Z(n63969) );
  IV U79041 ( .A(n58740), .Z(n58742) );
  NOR U79042 ( .A(n58742), .B(n58741), .Z(n63967) );
  XOR U79043 ( .A(n63969), .B(n63967), .Z(n63971) );
  XOR U79044 ( .A(n63970), .B(n63971), .Z(n60340) );
  IV U79045 ( .A(n58743), .Z(n58745) );
  NOR U79046 ( .A(n58745), .B(n58744), .Z(n58746) );
  NOR U79047 ( .A(n60339), .B(n58746), .Z(n58747) );
  XOR U79048 ( .A(n60340), .B(n58747), .Z(n63974) );
  XOR U79049 ( .A(n58748), .B(n63974), .Z(n63990) );
  XOR U79050 ( .A(n63988), .B(n63990), .Z(n60329) );
  XOR U79051 ( .A(n60328), .B(n60329), .Z(n63987) );
  XOR U79052 ( .A(n63985), .B(n63987), .Z(n60324) );
  XOR U79053 ( .A(n60322), .B(n60324), .Z(n60326) );
  XOR U79054 ( .A(n60325), .B(n60326), .Z(n60320) );
  XOR U79055 ( .A(n58749), .B(n60320), .Z(n60310) );
  IV U79056 ( .A(n58750), .Z(n58751) );
  NOR U79057 ( .A(n58752), .B(n58751), .Z(n60313) );
  IV U79058 ( .A(n58753), .Z(n58754) );
  NOR U79059 ( .A(n58755), .B(n58754), .Z(n60309) );
  NOR U79060 ( .A(n60313), .B(n60309), .Z(n58756) );
  XOR U79061 ( .A(n60310), .B(n58756), .Z(n60306) );
  IV U79062 ( .A(n58757), .Z(n58758) );
  NOR U79063 ( .A(n58758), .B(n58761), .Z(n58768) );
  IV U79064 ( .A(n58768), .Z(n79790) );
  NOR U79065 ( .A(n60306), .B(n79790), .Z(n65646) );
  IV U79066 ( .A(n58762), .Z(n58759) );
  NOR U79067 ( .A(n58759), .B(n58761), .Z(n65652) );
  IV U79068 ( .A(n58760), .Z(n58764) );
  XOR U79069 ( .A(n58762), .B(n58761), .Z(n58763) );
  NOR U79070 ( .A(n58764), .B(n58763), .Z(n65648) );
  NOR U79071 ( .A(n65652), .B(n65648), .Z(n60307) );
  IV U79072 ( .A(n58765), .Z(n58767) );
  NOR U79073 ( .A(n58767), .B(n58766), .Z(n60304) );
  XOR U79074 ( .A(n60304), .B(n60306), .Z(n65649) );
  XOR U79075 ( .A(n60307), .B(n65649), .Z(n79792) );
  NOR U79076 ( .A(n58768), .B(n79792), .Z(n58769) );
  NOR U79077 ( .A(n65646), .B(n58769), .Z(n60302) );
  IV U79078 ( .A(n58770), .Z(n58771) );
  NOR U79079 ( .A(n58772), .B(n58771), .Z(n60301) );
  NOR U79080 ( .A(n58773), .B(n64002), .Z(n58774) );
  NOR U79081 ( .A(n60301), .B(n58774), .Z(n58775) );
  XOR U79082 ( .A(n60302), .B(n58775), .Z(n60300) );
  IV U79083 ( .A(n58776), .Z(n58778) );
  NOR U79084 ( .A(n58778), .B(n58777), .Z(n58779) );
  IV U79085 ( .A(n58779), .Z(n58785) );
  NOR U79086 ( .A(n60300), .B(n58785), .Z(n69253) );
  IV U79087 ( .A(n58780), .Z(n58781) );
  NOR U79088 ( .A(n58782), .B(n58781), .Z(n60298) );
  XOR U79089 ( .A(n60298), .B(n60300), .Z(n64013) );
  IV U79090 ( .A(n58783), .Z(n58784) );
  NOR U79091 ( .A(n69271), .B(n58784), .Z(n58786) );
  IV U79092 ( .A(n58786), .Z(n64012) );
  XOR U79093 ( .A(n64013), .B(n64012), .Z(n58788) );
  NOR U79094 ( .A(n58786), .B(n58785), .Z(n58787) );
  NOR U79095 ( .A(n58788), .B(n58787), .Z(n58789) );
  NOR U79096 ( .A(n69253), .B(n58789), .Z(n64014) );
  IV U79097 ( .A(n58790), .Z(n58791) );
  NOR U79098 ( .A(n58792), .B(n58791), .Z(n64019) );
  IV U79099 ( .A(n58793), .Z(n58794) );
  NOR U79100 ( .A(n69271), .B(n58794), .Z(n64015) );
  NOR U79101 ( .A(n64019), .B(n64015), .Z(n58795) );
  XOR U79102 ( .A(n64014), .B(n58795), .Z(n64023) );
  XOR U79103 ( .A(n64021), .B(n64023), .Z(n64025) );
  NOR U79104 ( .A(n58802), .B(n64025), .Z(n65634) );
  IV U79105 ( .A(n58796), .Z(n58798) );
  NOR U79106 ( .A(n58798), .B(n58797), .Z(n64028) );
  IV U79107 ( .A(n58799), .Z(n58800) );
  NOR U79108 ( .A(n58801), .B(n58800), .Z(n64024) );
  XOR U79109 ( .A(n64024), .B(n64025), .Z(n64029) );
  IV U79110 ( .A(n64029), .Z(n58803) );
  XOR U79111 ( .A(n64028), .B(n58803), .Z(n58805) );
  NOR U79112 ( .A(n58803), .B(n58802), .Z(n58804) );
  NOR U79113 ( .A(n58805), .B(n58804), .Z(n58806) );
  NOR U79114 ( .A(n65634), .B(n58806), .Z(n64031) );
  XOR U79115 ( .A(n64032), .B(n64031), .Z(n64035) );
  NOR U79116 ( .A(n58811), .B(n64035), .Z(n69274) );
  IV U79117 ( .A(n58807), .Z(n65625) );
  NOR U79118 ( .A(n65622), .B(n65625), .Z(n64034) );
  XOR U79119 ( .A(n64034), .B(n64035), .Z(n60297) );
  IV U79120 ( .A(n58808), .Z(n58809) );
  NOR U79121 ( .A(n58810), .B(n58809), .Z(n58812) );
  IV U79122 ( .A(n58812), .Z(n60296) );
  XOR U79123 ( .A(n60297), .B(n60296), .Z(n58814) );
  NOR U79124 ( .A(n58812), .B(n58811), .Z(n58813) );
  NOR U79125 ( .A(n58814), .B(n58813), .Z(n58815) );
  NOR U79126 ( .A(n69274), .B(n58815), .Z(n60290) );
  XOR U79127 ( .A(n60292), .B(n60290), .Z(n60293) );
  NOR U79128 ( .A(n58816), .B(n60293), .Z(n65609) );
  IV U79129 ( .A(n58817), .Z(n58818) );
  NOR U79130 ( .A(n58819), .B(n58818), .Z(n58820) );
  IV U79131 ( .A(n58820), .Z(n60294) );
  XOR U79132 ( .A(n60294), .B(n60293), .Z(n58821) );
  NOR U79133 ( .A(n58822), .B(n58821), .Z(n64042) );
  NOR U79134 ( .A(n65609), .B(n64042), .Z(n60288) );
  IV U79135 ( .A(n58823), .Z(n58829) );
  IV U79136 ( .A(n58824), .Z(n58825) );
  NOR U79137 ( .A(n58829), .B(n58825), .Z(n60287) );
  NOR U79138 ( .A(n64040), .B(n60287), .Z(n58826) );
  XOR U79139 ( .A(n60288), .B(n58826), .Z(n60286) );
  IV U79140 ( .A(n58827), .Z(n58828) );
  NOR U79141 ( .A(n58829), .B(n58828), .Z(n60284) );
  IV U79142 ( .A(n58830), .Z(n58831) );
  NOR U79143 ( .A(n58832), .B(n58831), .Z(n60282) );
  NOR U79144 ( .A(n60284), .B(n60282), .Z(n58833) );
  XOR U79145 ( .A(n60286), .B(n58833), .Z(n60280) );
  IV U79146 ( .A(n58834), .Z(n58836) );
  NOR U79147 ( .A(n58836), .B(n58835), .Z(n60279) );
  IV U79148 ( .A(n58837), .Z(n58838) );
  NOR U79149 ( .A(n58839), .B(n58838), .Z(n64045) );
  NOR U79150 ( .A(n60279), .B(n64045), .Z(n58840) );
  XOR U79151 ( .A(n60280), .B(n58840), .Z(n64050) );
  XOR U79152 ( .A(n64048), .B(n64050), .Z(n60274) );
  XOR U79153 ( .A(n60273), .B(n60274), .Z(n60277) );
  XOR U79154 ( .A(n60276), .B(n60277), .Z(n60271) );
  XOR U79155 ( .A(n58841), .B(n60271), .Z(n60265) );
  XOR U79156 ( .A(n60266), .B(n60265), .Z(n70621) );
  IV U79157 ( .A(n58842), .Z(n58843) );
  NOR U79158 ( .A(n58844), .B(n58843), .Z(n70616) );
  IV U79159 ( .A(n58845), .Z(n58847) );
  NOR U79160 ( .A(n58847), .B(n58846), .Z(n70624) );
  NOR U79161 ( .A(n70616), .B(n70624), .Z(n64053) );
  XOR U79162 ( .A(n70621), .B(n64053), .Z(n64054) );
  XOR U79163 ( .A(n64056), .B(n64054), .Z(n60263) );
  XOR U79164 ( .A(n60262), .B(n60263), .Z(n60252) );
  IV U79165 ( .A(n58848), .Z(n58849) );
  NOR U79166 ( .A(n58850), .B(n58849), .Z(n58851) );
  IV U79167 ( .A(n58851), .Z(n58857) );
  NOR U79168 ( .A(n60252), .B(n58857), .Z(n69299) );
  NOR U79169 ( .A(n60253), .B(n58852), .Z(n58853) );
  XOR U79170 ( .A(n60252), .B(n58853), .Z(n60247) );
  IV U79171 ( .A(n58854), .Z(n58856) );
  NOR U79172 ( .A(n58856), .B(n58855), .Z(n58858) );
  IV U79173 ( .A(n58858), .Z(n60246) );
  XOR U79174 ( .A(n60247), .B(n60246), .Z(n58860) );
  NOR U79175 ( .A(n58858), .B(n58857), .Z(n58859) );
  NOR U79176 ( .A(n58860), .B(n58859), .Z(n58861) );
  NOR U79177 ( .A(n69299), .B(n58861), .Z(n60243) );
  XOR U79178 ( .A(n58862), .B(n60243), .Z(n64062) );
  XOR U79179 ( .A(n64060), .B(n64062), .Z(n64064) );
  XOR U79180 ( .A(n64063), .B(n64064), .Z(n64068) );
  XOR U79181 ( .A(n64067), .B(n64068), .Z(n64071) );
  XOR U79182 ( .A(n64070), .B(n64071), .Z(n60240) );
  IV U79183 ( .A(n58863), .Z(n58864) );
  NOR U79184 ( .A(n58865), .B(n58864), .Z(n60238) );
  XOR U79185 ( .A(n60240), .B(n60238), .Z(n64075) );
  XOR U79186 ( .A(n64074), .B(n64075), .Z(n64078) );
  IV U79187 ( .A(n58866), .Z(n58867) );
  NOR U79188 ( .A(n58868), .B(n58867), .Z(n64077) );
  IV U79189 ( .A(n58869), .Z(n58871) );
  NOR U79190 ( .A(n58871), .B(n58870), .Z(n60236) );
  NOR U79191 ( .A(n64077), .B(n60236), .Z(n58872) );
  XOR U79192 ( .A(n64078), .B(n58872), .Z(n58873) );
  IV U79193 ( .A(n58873), .Z(n64116) );
  XOR U79194 ( .A(n58874), .B(n64116), .Z(n64113) );
  XOR U79195 ( .A(n58875), .B(n64113), .Z(n60228) );
  XOR U79196 ( .A(n58876), .B(n60228), .Z(n60227) );
  XOR U79197 ( .A(n60225), .B(n60227), .Z(n60224) );
  XOR U79198 ( .A(n58877), .B(n60224), .Z(n58878) );
  IV U79199 ( .A(n58878), .Z(n64122) );
  XOR U79200 ( .A(n64121), .B(n64122), .Z(n64125) );
  XOR U79201 ( .A(n64124), .B(n64125), .Z(n60218) );
  IV U79202 ( .A(n60218), .Z(n58886) );
  IV U79203 ( .A(n58879), .Z(n58881) );
  NOR U79204 ( .A(n58881), .B(n58880), .Z(n60214) );
  IV U79205 ( .A(n58882), .Z(n58884) );
  NOR U79206 ( .A(n58884), .B(n58883), .Z(n60216) );
  NOR U79207 ( .A(n60214), .B(n60216), .Z(n58885) );
  XOR U79208 ( .A(n58886), .B(n58885), .Z(n60210) );
  NOR U79209 ( .A(n58888), .B(n58887), .Z(n58889) );
  IV U79210 ( .A(n58889), .Z(n58890) );
  NOR U79211 ( .A(n58891), .B(n58890), .Z(n60208) );
  XOR U79212 ( .A(n60210), .B(n60208), .Z(n60212) );
  XOR U79213 ( .A(n58892), .B(n60212), .Z(n64128) );
  XOR U79214 ( .A(n64129), .B(n64128), .Z(n60202) );
  IV U79215 ( .A(n60202), .Z(n58900) );
  IV U79216 ( .A(n58893), .Z(n58895) );
  NOR U79217 ( .A(n58895), .B(n58894), .Z(n64130) );
  IV U79218 ( .A(n58896), .Z(n58898) );
  NOR U79219 ( .A(n58898), .B(n58897), .Z(n60201) );
  NOR U79220 ( .A(n64130), .B(n60201), .Z(n58899) );
  XOR U79221 ( .A(n58900), .B(n58899), .Z(n60200) );
  XOR U79222 ( .A(n60198), .B(n60200), .Z(n65509) );
  XOR U79223 ( .A(n64133), .B(n65509), .Z(n60195) );
  NOR U79224 ( .A(n58902), .B(n58901), .Z(n64134) );
  IV U79225 ( .A(n58903), .Z(n58905) );
  IV U79226 ( .A(n58904), .Z(n58908) );
  NOR U79227 ( .A(n58905), .B(n58908), .Z(n60196) );
  NOR U79228 ( .A(n64134), .B(n60196), .Z(n58906) );
  XOR U79229 ( .A(n60195), .B(n58906), .Z(n60194) );
  IV U79230 ( .A(n58907), .Z(n58909) );
  NOR U79231 ( .A(n58909), .B(n58908), .Z(n60192) );
  XOR U79232 ( .A(n60194), .B(n60192), .Z(n65492) );
  XOR U79233 ( .A(n60191), .B(n65492), .Z(n64142) );
  XOR U79234 ( .A(n64144), .B(n64142), .Z(n75894) );
  IV U79235 ( .A(n58910), .Z(n58911) );
  NOR U79236 ( .A(n75892), .B(n58911), .Z(n75895) );
  NOR U79237 ( .A(n65487), .B(n65485), .Z(n58912) );
  NOR U79238 ( .A(n75895), .B(n58912), .Z(n58913) );
  XOR U79239 ( .A(n75894), .B(n58913), .Z(n64154) );
  XOR U79240 ( .A(n58914), .B(n64154), .Z(n64166) );
  IV U79241 ( .A(n58915), .Z(n58917) );
  NOR U79242 ( .A(n58917), .B(n58916), .Z(n64164) );
  XOR U79243 ( .A(n64166), .B(n64164), .Z(n64170) );
  IV U79244 ( .A(n58918), .Z(n58920) );
  NOR U79245 ( .A(n58920), .B(n58919), .Z(n64168) );
  XOR U79246 ( .A(n64170), .B(n64168), .Z(n64176) );
  IV U79247 ( .A(n58921), .Z(n58922) );
  NOR U79248 ( .A(n58923), .B(n58922), .Z(n64171) );
  IV U79249 ( .A(n58924), .Z(n58925) );
  NOR U79250 ( .A(n58926), .B(n58925), .Z(n64175) );
  NOR U79251 ( .A(n64171), .B(n64175), .Z(n58927) );
  XOR U79252 ( .A(n64176), .B(n58927), .Z(n60184) );
  XOR U79253 ( .A(n60185), .B(n60184), .Z(n60188) );
  XOR U79254 ( .A(n60187), .B(n60188), .Z(n60179) );
  XOR U79255 ( .A(n60178), .B(n60179), .Z(n60182) );
  XOR U79256 ( .A(n58928), .B(n60182), .Z(n58929) );
  IV U79257 ( .A(n58929), .Z(n60174) );
  XOR U79258 ( .A(n60172), .B(n60174), .Z(n60165) );
  NOR U79259 ( .A(n60164), .B(n60169), .Z(n58930) );
  NOR U79260 ( .A(n58930), .B(n60166), .Z(n58931) );
  XOR U79261 ( .A(n60165), .B(n58931), .Z(n64181) );
  XOR U79262 ( .A(n64180), .B(n64181), .Z(n64184) );
  XOR U79263 ( .A(n64183), .B(n64184), .Z(n60160) );
  XOR U79264 ( .A(n60159), .B(n60160), .Z(n64192) );
  IV U79265 ( .A(n58932), .Z(n58933) );
  NOR U79266 ( .A(n58934), .B(n58933), .Z(n60162) );
  IV U79267 ( .A(n58935), .Z(n58936) );
  NOR U79268 ( .A(n58940), .B(n58936), .Z(n64190) );
  NOR U79269 ( .A(n60162), .B(n64190), .Z(n58937) );
  XOR U79270 ( .A(n64192), .B(n58937), .Z(n58938) );
  IV U79271 ( .A(n58938), .Z(n64195) );
  IV U79272 ( .A(n58939), .Z(n58941) );
  NOR U79273 ( .A(n58941), .B(n58940), .Z(n64188) );
  XOR U79274 ( .A(n64195), .B(n64188), .Z(n64198) );
  XOR U79275 ( .A(n58942), .B(n64198), .Z(n64204) );
  IV U79276 ( .A(n58943), .Z(n58952) );
  IV U79277 ( .A(n58944), .Z(n58945) );
  NOR U79278 ( .A(n58952), .B(n58945), .Z(n64210) );
  NOR U79279 ( .A(n64203), .B(n64210), .Z(n58946) );
  XOR U79280 ( .A(n64204), .B(n58946), .Z(n64209) );
  IV U79281 ( .A(n58947), .Z(n58948) );
  NOR U79282 ( .A(n58949), .B(n58948), .Z(n60153) );
  IV U79283 ( .A(n58950), .Z(n58951) );
  NOR U79284 ( .A(n58952), .B(n58951), .Z(n64207) );
  NOR U79285 ( .A(n60153), .B(n64207), .Z(n58953) );
  XOR U79286 ( .A(n64209), .B(n58953), .Z(n60137) );
  IV U79287 ( .A(n58954), .Z(n58955) );
  NOR U79288 ( .A(n60152), .B(n58955), .Z(n58958) );
  IV U79289 ( .A(n58956), .Z(n58957) );
  NOR U79290 ( .A(n58957), .B(n58961), .Z(n64219) );
  NOR U79291 ( .A(n58958), .B(n64219), .Z(n58959) );
  XOR U79292 ( .A(n60137), .B(n58959), .Z(n64218) );
  IV U79293 ( .A(n58960), .Z(n58962) );
  NOR U79294 ( .A(n58962), .B(n58961), .Z(n64216) );
  XOR U79295 ( .A(n64218), .B(n64216), .Z(n60135) );
  XOR U79296 ( .A(n60134), .B(n60135), .Z(n60129) );
  XOR U79297 ( .A(n60128), .B(n60129), .Z(n60132) );
  XOR U79298 ( .A(n60131), .B(n60132), .Z(n58963) );
  NOR U79299 ( .A(n58964), .B(n58963), .Z(n65427) );
  IV U79300 ( .A(n58965), .Z(n58967) );
  NOR U79301 ( .A(n58967), .B(n58966), .Z(n60125) );
  NOR U79302 ( .A(n60131), .B(n60125), .Z(n58968) );
  XOR U79303 ( .A(n60132), .B(n58968), .Z(n58969) );
  NOR U79304 ( .A(n58970), .B(n58969), .Z(n64225) );
  NOR U79305 ( .A(n65427), .B(n64225), .Z(n60121) );
  IV U79306 ( .A(n58971), .Z(n58972) );
  NOR U79307 ( .A(n58973), .B(n58972), .Z(n64224) );
  NOR U79308 ( .A(n58974), .B(n60122), .Z(n58975) );
  NOR U79309 ( .A(n64224), .B(n58975), .Z(n58976) );
  XOR U79310 ( .A(n60121), .B(n58976), .Z(n60119) );
  IV U79311 ( .A(n58977), .Z(n58978) );
  NOR U79312 ( .A(n58979), .B(n58978), .Z(n58980) );
  IV U79313 ( .A(n58980), .Z(n58987) );
  NOR U79314 ( .A(n60119), .B(n58987), .Z(n69402) );
  IV U79315 ( .A(n58981), .Z(n58983) );
  NOR U79316 ( .A(n58983), .B(n58982), .Z(n60111) );
  IV U79317 ( .A(n58984), .Z(n58986) );
  NOR U79318 ( .A(n58986), .B(n58985), .Z(n60117) );
  XOR U79319 ( .A(n60117), .B(n60119), .Z(n60112) );
  IV U79320 ( .A(n60112), .Z(n58988) );
  XOR U79321 ( .A(n60111), .B(n58988), .Z(n58990) );
  NOR U79322 ( .A(n58988), .B(n58987), .Z(n58989) );
  NOR U79323 ( .A(n58990), .B(n58989), .Z(n58991) );
  NOR U79324 ( .A(n69402), .B(n58991), .Z(n58992) );
  IV U79325 ( .A(n58992), .Z(n60115) );
  XOR U79326 ( .A(n60114), .B(n60115), .Z(n60106) );
  XOR U79327 ( .A(n60105), .B(n60106), .Z(n60109) );
  IV U79328 ( .A(n58993), .Z(n58994) );
  NOR U79329 ( .A(n58995), .B(n58994), .Z(n60108) );
  IV U79330 ( .A(n58996), .Z(n58997) );
  NOR U79331 ( .A(n58998), .B(n58997), .Z(n60103) );
  NOR U79332 ( .A(n60108), .B(n60103), .Z(n58999) );
  XOR U79333 ( .A(n60109), .B(n58999), .Z(n60097) );
  IV U79334 ( .A(n59000), .Z(n59002) );
  NOR U79335 ( .A(n59002), .B(n59001), .Z(n60100) );
  IV U79336 ( .A(n59003), .Z(n59005) );
  NOR U79337 ( .A(n59005), .B(n59004), .Z(n60098) );
  NOR U79338 ( .A(n60100), .B(n60098), .Z(n59006) );
  XOR U79339 ( .A(n60097), .B(n59006), .Z(n65395) );
  IV U79340 ( .A(n59007), .Z(n59011) );
  NOR U79341 ( .A(n59009), .B(n59008), .Z(n59010) );
  IV U79342 ( .A(n59010), .Z(n59013) );
  NOR U79343 ( .A(n59011), .B(n59013), .Z(n60091) );
  IV U79344 ( .A(n59012), .Z(n59014) );
  NOR U79345 ( .A(n59014), .B(n59013), .Z(n65396) );
  NOR U79346 ( .A(n60091), .B(n65396), .Z(n59015) );
  XOR U79347 ( .A(n65395), .B(n59015), .Z(n59016) );
  IV U79348 ( .A(n59016), .Z(n60093) );
  XOR U79349 ( .A(n59017), .B(n60093), .Z(n60086) );
  IV U79350 ( .A(n59018), .Z(n59020) );
  NOR U79351 ( .A(n59020), .B(n59019), .Z(n60087) );
  NOR U79352 ( .A(n64238), .B(n60087), .Z(n59021) );
  XOR U79353 ( .A(n60086), .B(n59021), .Z(n64248) );
  XOR U79354 ( .A(n59022), .B(n64248), .Z(n60083) );
  IV U79355 ( .A(n59023), .Z(n59025) );
  NOR U79356 ( .A(n59025), .B(n59024), .Z(n64243) );
  NOR U79357 ( .A(n59027), .B(n59026), .Z(n60082) );
  NOR U79358 ( .A(n64243), .B(n60082), .Z(n59028) );
  XOR U79359 ( .A(n60083), .B(n59028), .Z(n60079) );
  NOR U79360 ( .A(n60081), .B(n60078), .Z(n59029) );
  XOR U79361 ( .A(n60079), .B(n59029), .Z(n60075) );
  XOR U79362 ( .A(n60072), .B(n60075), .Z(n69434) );
  XOR U79363 ( .A(n69435), .B(n69434), .Z(n59030) );
  IV U79364 ( .A(n59030), .Z(n60070) );
  IV U79365 ( .A(n59031), .Z(n65357) );
  NOR U79366 ( .A(n65357), .B(n59032), .Z(n64252) );
  IV U79367 ( .A(n59033), .Z(n59035) );
  NOR U79368 ( .A(n59035), .B(n59034), .Z(n60069) );
  NOR U79369 ( .A(n64252), .B(n60069), .Z(n59036) );
  XOR U79370 ( .A(n60070), .B(n59036), .Z(n60059) );
  NOR U79371 ( .A(n59037), .B(n60059), .Z(n59045) );
  IV U79372 ( .A(n59037), .Z(n59043) );
  IV U79373 ( .A(n59038), .Z(n59040) );
  NOR U79374 ( .A(n59040), .B(n59039), .Z(n60066) );
  IV U79375 ( .A(n59041), .Z(n60064) );
  XOR U79376 ( .A(n60064), .B(n60059), .Z(n60067) );
  XOR U79377 ( .A(n60066), .B(n60067), .Z(n59042) );
  NOR U79378 ( .A(n59043), .B(n59042), .Z(n59044) );
  NOR U79379 ( .A(n59045), .B(n59044), .Z(n64258) );
  XOR U79380 ( .A(n64256), .B(n64258), .Z(n64260) );
  NOR U79381 ( .A(n59052), .B(n64260), .Z(n65341) );
  IV U79382 ( .A(n59046), .Z(n59047) );
  NOR U79383 ( .A(n59048), .B(n59047), .Z(n60056) );
  IV U79384 ( .A(n59049), .Z(n59050) );
  NOR U79385 ( .A(n59051), .B(n59050), .Z(n64259) );
  XOR U79386 ( .A(n64259), .B(n64260), .Z(n60057) );
  IV U79387 ( .A(n60057), .Z(n59053) );
  XOR U79388 ( .A(n60056), .B(n59053), .Z(n59055) );
  NOR U79389 ( .A(n59053), .B(n59052), .Z(n59054) );
  NOR U79390 ( .A(n59055), .B(n59054), .Z(n59056) );
  NOR U79391 ( .A(n65341), .B(n59056), .Z(n59057) );
  IV U79392 ( .A(n59057), .Z(n60051) );
  XOR U79393 ( .A(n60050), .B(n60051), .Z(n60054) );
  IV U79394 ( .A(n59058), .Z(n59059) );
  NOR U79395 ( .A(n59059), .B(n59062), .Z(n60047) );
  NOR U79396 ( .A(n60053), .B(n60047), .Z(n59060) );
  XOR U79397 ( .A(n60054), .B(n59060), .Z(n59061) );
  IV U79398 ( .A(n59061), .Z(n60038) );
  NOR U79399 ( .A(n59063), .B(n59062), .Z(n59064) );
  IV U79400 ( .A(n59064), .Z(n60037) );
  IV U79401 ( .A(n59065), .Z(n59066) );
  NOR U79402 ( .A(n60037), .B(n59066), .Z(n59067) );
  XOR U79403 ( .A(n60038), .B(n59067), .Z(n60035) );
  XOR U79404 ( .A(n60034), .B(n60035), .Z(n60029) );
  IV U79405 ( .A(n60029), .Z(n60027) );
  XOR U79406 ( .A(n60028), .B(n60027), .Z(n65334) );
  XOR U79407 ( .A(n59068), .B(n65334), .Z(n60020) );
  XOR U79408 ( .A(n59069), .B(n60020), .Z(n60018) );
  XOR U79409 ( .A(n59070), .B(n60018), .Z(n60009) );
  NOR U79410 ( .A(n59072), .B(n59071), .Z(n60012) );
  NOR U79411 ( .A(n59074), .B(n59073), .Z(n59075) );
  IV U79412 ( .A(n59075), .Z(n59081) );
  IV U79413 ( .A(n59076), .Z(n59078) );
  NOR U79414 ( .A(n59078), .B(n59077), .Z(n59079) );
  IV U79415 ( .A(n59079), .Z(n59080) );
  NOR U79416 ( .A(n59081), .B(n59080), .Z(n60010) );
  NOR U79417 ( .A(n60012), .B(n60010), .Z(n59082) );
  XOR U79418 ( .A(n60009), .B(n59082), .Z(n64277) );
  XOR U79419 ( .A(n64275), .B(n64277), .Z(n69482) );
  XOR U79420 ( .A(n59083), .B(n69482), .Z(n59084) );
  IV U79421 ( .A(n59084), .Z(n64282) );
  XOR U79422 ( .A(n64281), .B(n64282), .Z(n64287) );
  XOR U79423 ( .A(n64286), .B(n64287), .Z(n64290) );
  XOR U79424 ( .A(n64289), .B(n64290), .Z(n65291) );
  IV U79425 ( .A(n59085), .Z(n59086) );
  NOR U79426 ( .A(n59086), .B(n59088), .Z(n65295) );
  IV U79427 ( .A(n59087), .Z(n59089) );
  NOR U79428 ( .A(n59089), .B(n59088), .Z(n65290) );
  NOR U79429 ( .A(n65295), .B(n65290), .Z(n64296) );
  XOR U79430 ( .A(n65291), .B(n64296), .Z(n64297) );
  XOR U79431 ( .A(n64299), .B(n64297), .Z(n64295) );
  XOR U79432 ( .A(n64293), .B(n64295), .Z(n60008) );
  XOR U79433 ( .A(n59090), .B(n60008), .Z(n64304) );
  XOR U79434 ( .A(n64306), .B(n64304), .Z(n64308) );
  IV U79435 ( .A(n59091), .Z(n59093) );
  NOR U79436 ( .A(n59093), .B(n59092), .Z(n64307) );
  IV U79437 ( .A(n59094), .Z(n59096) );
  NOR U79438 ( .A(n59096), .B(n59095), .Z(n60001) );
  NOR U79439 ( .A(n64307), .B(n60001), .Z(n59097) );
  XOR U79440 ( .A(n64308), .B(n59097), .Z(n59998) );
  XOR U79441 ( .A(n60000), .B(n59998), .Z(n64316) );
  XOR U79442 ( .A(n64315), .B(n64316), .Z(n64325) );
  XOR U79443 ( .A(n59098), .B(n64325), .Z(n59995) );
  XOR U79444 ( .A(n59099), .B(n59995), .Z(n59994) );
  XOR U79445 ( .A(n59992), .B(n59994), .Z(n64339) );
  XOR U79446 ( .A(n59100), .B(n64339), .Z(n59989) );
  XOR U79447 ( .A(n59101), .B(n59989), .Z(n64351) );
  XOR U79448 ( .A(n59102), .B(n64351), .Z(n59988) );
  IV U79449 ( .A(n59103), .Z(n59104) );
  NOR U79450 ( .A(n59105), .B(n59104), .Z(n59986) );
  XOR U79451 ( .A(n59988), .B(n59986), .Z(n59979) );
  XOR U79452 ( .A(n59978), .B(n59979), .Z(n59982) );
  XOR U79453 ( .A(n59981), .B(n59982), .Z(n59976) );
  IV U79454 ( .A(n59106), .Z(n59107) );
  NOR U79455 ( .A(n59108), .B(n59107), .Z(n59969) );
  IV U79456 ( .A(n59109), .Z(n59111) );
  NOR U79457 ( .A(n59111), .B(n59110), .Z(n59974) );
  NOR U79458 ( .A(n59969), .B(n59974), .Z(n59112) );
  XOR U79459 ( .A(n59976), .B(n59112), .Z(n59972) );
  IV U79460 ( .A(n59113), .Z(n59115) );
  NOR U79461 ( .A(n59115), .B(n59114), .Z(n59971) );
  IV U79462 ( .A(n59116), .Z(n59118) );
  NOR U79463 ( .A(n59118), .B(n59117), .Z(n64358) );
  NOR U79464 ( .A(n59971), .B(n64358), .Z(n59119) );
  XOR U79465 ( .A(n59972), .B(n59119), .Z(n64357) );
  XOR U79466 ( .A(n64355), .B(n64357), .Z(n64363) );
  IV U79467 ( .A(n59120), .Z(n59121) );
  NOR U79468 ( .A(n59122), .B(n59121), .Z(n64362) );
  IV U79469 ( .A(n59123), .Z(n59124) );
  NOR U79470 ( .A(n59125), .B(n59124), .Z(n59967) );
  NOR U79471 ( .A(n64362), .B(n59967), .Z(n59126) );
  XOR U79472 ( .A(n64363), .B(n59126), .Z(n59960) );
  IV U79473 ( .A(n59127), .Z(n59129) );
  NOR U79474 ( .A(n59129), .B(n59128), .Z(n59963) );
  IV U79475 ( .A(n59130), .Z(n59132) );
  NOR U79476 ( .A(n59132), .B(n59131), .Z(n59961) );
  NOR U79477 ( .A(n59963), .B(n59961), .Z(n59133) );
  XOR U79478 ( .A(n59960), .B(n59133), .Z(n59958) );
  XOR U79479 ( .A(n59957), .B(n59958), .Z(n59951) );
  XOR U79480 ( .A(n59950), .B(n59951), .Z(n59944) );
  NOR U79481 ( .A(n59134), .B(n59947), .Z(n59137) );
  NOR U79482 ( .A(n59136), .B(n59135), .Z(n59943) );
  NOR U79483 ( .A(n59137), .B(n59943), .Z(n59138) );
  XOR U79484 ( .A(n59944), .B(n59138), .Z(n59139) );
  IV U79485 ( .A(n59139), .Z(n59942) );
  IV U79486 ( .A(n59140), .Z(n59142) );
  NOR U79487 ( .A(n59142), .B(n59141), .Z(n59143) );
  IV U79488 ( .A(n59143), .Z(n59146) );
  NOR U79489 ( .A(n59942), .B(n59146), .Z(n69552) );
  IV U79490 ( .A(n59144), .Z(n59145) );
  NOR U79491 ( .A(n59145), .B(n59153), .Z(n59937) );
  XOR U79492 ( .A(n59940), .B(n59942), .Z(n59938) );
  IV U79493 ( .A(n59938), .Z(n59147) );
  XOR U79494 ( .A(n59937), .B(n59147), .Z(n59149) );
  NOR U79495 ( .A(n59147), .B(n59146), .Z(n59148) );
  NOR U79496 ( .A(n59149), .B(n59148), .Z(n59150) );
  NOR U79497 ( .A(n69552), .B(n59150), .Z(n64371) );
  IV U79498 ( .A(n59151), .Z(n59152) );
  NOR U79499 ( .A(n59153), .B(n59152), .Z(n64370) );
  IV U79500 ( .A(n59154), .Z(n59155) );
  NOR U79501 ( .A(n59156), .B(n59155), .Z(n69560) );
  NOR U79502 ( .A(n64370), .B(n69560), .Z(n59157) );
  XOR U79503 ( .A(n64371), .B(n59157), .Z(n64378) );
  IV U79504 ( .A(n59158), .Z(n59160) );
  NOR U79505 ( .A(n59160), .B(n59159), .Z(n64376) );
  XOR U79506 ( .A(n64378), .B(n64376), .Z(n64380) );
  XOR U79507 ( .A(n64379), .B(n64380), .Z(n59932) );
  XOR U79508 ( .A(n59931), .B(n59932), .Z(n59936) );
  XOR U79509 ( .A(n59934), .B(n59936), .Z(n59926) );
  XOR U79510 ( .A(n59925), .B(n59926), .Z(n59929) );
  XOR U79511 ( .A(n59928), .B(n59929), .Z(n64390) );
  XOR U79512 ( .A(n59161), .B(n64390), .Z(n59162) );
  IV U79513 ( .A(n59162), .Z(n59923) );
  XOR U79514 ( .A(n59921), .B(n59923), .Z(n64397) );
  IV U79515 ( .A(n59163), .Z(n59165) );
  NOR U79516 ( .A(n59165), .B(n59164), .Z(n64396) );
  IV U79517 ( .A(n59166), .Z(n59168) );
  NOR U79518 ( .A(n59168), .B(n59167), .Z(n59919) );
  NOR U79519 ( .A(n64396), .B(n59919), .Z(n59169) );
  XOR U79520 ( .A(n64397), .B(n59169), .Z(n59914) );
  XOR U79521 ( .A(n59170), .B(n59914), .Z(n59911) );
  IV U79522 ( .A(n59911), .Z(n59177) );
  IV U79523 ( .A(n59171), .Z(n59173) );
  NOR U79524 ( .A(n59173), .B(n59172), .Z(n59910) );
  NOR U79525 ( .A(n59174), .B(n59904), .Z(n59175) );
  NOR U79526 ( .A(n59910), .B(n59175), .Z(n59176) );
  XOR U79527 ( .A(n59177), .B(n59176), .Z(n64402) );
  IV U79528 ( .A(n59178), .Z(n59179) );
  NOR U79529 ( .A(n59179), .B(n59188), .Z(n59186) );
  IV U79530 ( .A(n59186), .Z(n64415) );
  NOR U79531 ( .A(n64402), .B(n64415), .Z(n64404) );
  IV U79532 ( .A(n59180), .Z(n59182) );
  NOR U79533 ( .A(n59182), .B(n59181), .Z(n59901) );
  IV U79534 ( .A(n59183), .Z(n59184) );
  NOR U79535 ( .A(n59184), .B(n59188), .Z(n64400) );
  NOR U79536 ( .A(n59901), .B(n64400), .Z(n59185) );
  XOR U79537 ( .A(n64402), .B(n59185), .Z(n64410) );
  NOR U79538 ( .A(n59186), .B(n64410), .Z(n64406) );
  NOR U79539 ( .A(n64404), .B(n64406), .Z(n64420) );
  IV U79540 ( .A(n59187), .Z(n59189) );
  NOR U79541 ( .A(n59189), .B(n59188), .Z(n64409) );
  IV U79542 ( .A(n59190), .Z(n59196) );
  IV U79543 ( .A(n59191), .Z(n59192) );
  NOR U79544 ( .A(n59196), .B(n59192), .Z(n64421) );
  NOR U79545 ( .A(n64409), .B(n64421), .Z(n59193) );
  XOR U79546 ( .A(n64420), .B(n59193), .Z(n69598) );
  IV U79547 ( .A(n59194), .Z(n59195) );
  NOR U79548 ( .A(n59196), .B(n59195), .Z(n65191) );
  IV U79549 ( .A(n59197), .Z(n59201) );
  NOR U79550 ( .A(n59199), .B(n59198), .Z(n59200) );
  IV U79551 ( .A(n59200), .Z(n59209) );
  NOR U79552 ( .A(n59201), .B(n59209), .Z(n69594) );
  NOR U79553 ( .A(n65191), .B(n69594), .Z(n64424) );
  XOR U79554 ( .A(n69598), .B(n64424), .Z(n64425) );
  IV U79555 ( .A(n59202), .Z(n59204) );
  NOR U79556 ( .A(n59204), .B(n59203), .Z(n69604) );
  IV U79557 ( .A(n59205), .Z(n59207) );
  NOR U79558 ( .A(n59207), .B(n59206), .Z(n59208) );
  IV U79559 ( .A(n59208), .Z(n59210) );
  NOR U79560 ( .A(n59210), .B(n59209), .Z(n69599) );
  NOR U79561 ( .A(n69604), .B(n69599), .Z(n64426) );
  XOR U79562 ( .A(n64425), .B(n64426), .Z(n64431) );
  XOR U79563 ( .A(n64430), .B(n64431), .Z(n64434) );
  XOR U79564 ( .A(n64433), .B(n64434), .Z(n59899) );
  XOR U79565 ( .A(n59211), .B(n59899), .Z(n59212) );
  IV U79566 ( .A(n59212), .Z(n64438) );
  XOR U79567 ( .A(n64437), .B(n64438), .Z(n64440) );
  XOR U79568 ( .A(n64441), .B(n64440), .Z(n59892) );
  IV U79569 ( .A(n59213), .Z(n59214) );
  NOR U79570 ( .A(n59215), .B(n59214), .Z(n64443) );
  IV U79571 ( .A(n59216), .Z(n59217) );
  NOR U79572 ( .A(n59217), .B(n59220), .Z(n59893) );
  NOR U79573 ( .A(n64443), .B(n59893), .Z(n59218) );
  XOR U79574 ( .A(n59892), .B(n59218), .Z(n64451) );
  IV U79575 ( .A(n59219), .Z(n59221) );
  NOR U79576 ( .A(n59221), .B(n59220), .Z(n59222) );
  IV U79577 ( .A(n59222), .Z(n64450) );
  XOR U79578 ( .A(n64451), .B(n64450), .Z(n59225) );
  IV U79579 ( .A(n59225), .Z(n59223) );
  NOR U79580 ( .A(n59224), .B(n59223), .Z(n69623) );
  NOR U79581 ( .A(n59226), .B(n59225), .Z(n64459) );
  IV U79582 ( .A(n59227), .Z(n59228) );
  NOR U79583 ( .A(n59229), .B(n59228), .Z(n64457) );
  XOR U79584 ( .A(n64459), .B(n64457), .Z(n59230) );
  NOR U79585 ( .A(n69623), .B(n59230), .Z(n59231) );
  IV U79586 ( .A(n59231), .Z(n64464) );
  IV U79587 ( .A(n59232), .Z(n59234) );
  NOR U79588 ( .A(n59234), .B(n59233), .Z(n64455) );
  IV U79589 ( .A(n59235), .Z(n59237) );
  NOR U79590 ( .A(n59237), .B(n59236), .Z(n64463) );
  NOR U79591 ( .A(n64455), .B(n64463), .Z(n59238) );
  XOR U79592 ( .A(n64464), .B(n59238), .Z(n59881) );
  IV U79593 ( .A(n59239), .Z(n59241) );
  NOR U79594 ( .A(n59241), .B(n59240), .Z(n59884) );
  IV U79595 ( .A(n59242), .Z(n59243) );
  NOR U79596 ( .A(n59244), .B(n59243), .Z(n59882) );
  NOR U79597 ( .A(n59884), .B(n59882), .Z(n59245) );
  XOR U79598 ( .A(n59881), .B(n59245), .Z(n59889) );
  IV U79599 ( .A(n59246), .Z(n59247) );
  NOR U79600 ( .A(n59248), .B(n59247), .Z(n59888) );
  IV U79601 ( .A(n59249), .Z(n59251) );
  NOR U79602 ( .A(n59251), .B(n59250), .Z(n59878) );
  NOR U79603 ( .A(n59888), .B(n59878), .Z(n59252) );
  XOR U79604 ( .A(n59889), .B(n59252), .Z(n64469) );
  IV U79605 ( .A(n59253), .Z(n59255) );
  NOR U79606 ( .A(n59255), .B(n59254), .Z(n64472) );
  IV U79607 ( .A(n59256), .Z(n59258) );
  NOR U79608 ( .A(n59258), .B(n59257), .Z(n64470) );
  NOR U79609 ( .A(n64472), .B(n64470), .Z(n59259) );
  XOR U79610 ( .A(n64469), .B(n59259), .Z(n65165) );
  IV U79611 ( .A(n59260), .Z(n59262) );
  NOR U79612 ( .A(n59262), .B(n59261), .Z(n64467) );
  NOR U79613 ( .A(n64467), .B(n59263), .Z(n59264) );
  XOR U79614 ( .A(n65165), .B(n59264), .Z(n59875) );
  IV U79615 ( .A(n59265), .Z(n59267) );
  NOR U79616 ( .A(n59267), .B(n59266), .Z(n59268) );
  IV U79617 ( .A(n59268), .Z(n59876) );
  XOR U79618 ( .A(n69650), .B(n59876), .Z(n59269) );
  XOR U79619 ( .A(n59875), .B(n59269), .Z(n65159) );
  IV U79620 ( .A(n59270), .Z(n59271) );
  NOR U79621 ( .A(n59271), .B(n59277), .Z(n59272) );
  IV U79622 ( .A(n59272), .Z(n59873) );
  IV U79623 ( .A(n59273), .Z(n59274) );
  NOR U79624 ( .A(n59275), .B(n59274), .Z(n69656) );
  IV U79625 ( .A(n59276), .Z(n59278) );
  NOR U79626 ( .A(n59278), .B(n59277), .Z(n65157) );
  NOR U79627 ( .A(n69656), .B(n65157), .Z(n59874) );
  XOR U79628 ( .A(n59873), .B(n59874), .Z(n59279) );
  XOR U79629 ( .A(n65159), .B(n59279), .Z(n59872) );
  IV U79630 ( .A(n59280), .Z(n59281) );
  NOR U79631 ( .A(n59282), .B(n59281), .Z(n59868) );
  NOR U79632 ( .A(n59870), .B(n59868), .Z(n59283) );
  XOR U79633 ( .A(n59872), .B(n59283), .Z(n59862) );
  XOR U79634 ( .A(n59863), .B(n59862), .Z(n59865) );
  XOR U79635 ( .A(n59284), .B(n59865), .Z(n64483) );
  XOR U79636 ( .A(n59285), .B(n64483), .Z(n64491) );
  XOR U79637 ( .A(n64489), .B(n64491), .Z(n64496) );
  XOR U79638 ( .A(n59286), .B(n64496), .Z(n59851) );
  XOR U79639 ( .A(n59287), .B(n59851), .Z(n59849) );
  XOR U79640 ( .A(n59848), .B(n59849), .Z(n65121) );
  XOR U79641 ( .A(n65120), .B(n65121), .Z(n59845) );
  XOR U79642 ( .A(n59288), .B(n59845), .Z(n59289) );
  IV U79643 ( .A(n59289), .Z(n59841) );
  XOR U79644 ( .A(n59290), .B(n59841), .Z(n59301) );
  IV U79645 ( .A(n59301), .Z(n59294) );
  IV U79646 ( .A(n59291), .Z(n59292) );
  NOR U79647 ( .A(n59293), .B(n59292), .Z(n59297) );
  NOR U79648 ( .A(n59294), .B(n59297), .Z(n59295) );
  IV U79649 ( .A(n59295), .Z(n59296) );
  NOR U79650 ( .A(n59299), .B(n59296), .Z(n59303) );
  IV U79651 ( .A(n59297), .Z(n59298) );
  NOR U79652 ( .A(n59841), .B(n59298), .Z(n69703) );
  IV U79653 ( .A(n59299), .Z(n59300) );
  NOR U79654 ( .A(n59301), .B(n59300), .Z(n65109) );
  NOR U79655 ( .A(n69703), .B(n65109), .Z(n59302) );
  IV U79656 ( .A(n59302), .Z(n64508) );
  NOR U79657 ( .A(n59303), .B(n64508), .Z(n64506) );
  IV U79658 ( .A(n59304), .Z(n59305) );
  NOR U79659 ( .A(n59306), .B(n59305), .Z(n64505) );
  IV U79660 ( .A(n59307), .Z(n59309) );
  NOR U79661 ( .A(n59309), .B(n59308), .Z(n64510) );
  NOR U79662 ( .A(n64505), .B(n64510), .Z(n59310) );
  XOR U79663 ( .A(n64506), .B(n59310), .Z(n59833) );
  XOR U79664 ( .A(n59311), .B(n59833), .Z(n59312) );
  IV U79665 ( .A(n59312), .Z(n59824) );
  NOR U79666 ( .A(n59321), .B(n59824), .Z(n65096) );
  IV U79667 ( .A(n59313), .Z(n59314) );
  NOR U79668 ( .A(n59314), .B(n59327), .Z(n59818) );
  NOR U79669 ( .A(n59316), .B(n59315), .Z(n59317) );
  IV U79670 ( .A(n59317), .Z(n59825) );
  IV U79671 ( .A(n59318), .Z(n59319) );
  NOR U79672 ( .A(n59825), .B(n59319), .Z(n59320) );
  XOR U79673 ( .A(n59824), .B(n59320), .Z(n59819) );
  IV U79674 ( .A(n59819), .Z(n59322) );
  XOR U79675 ( .A(n59818), .B(n59322), .Z(n59324) );
  NOR U79676 ( .A(n59322), .B(n59321), .Z(n59323) );
  NOR U79677 ( .A(n59324), .B(n59323), .Z(n59325) );
  NOR U79678 ( .A(n65096), .B(n59325), .Z(n59815) );
  IV U79679 ( .A(n59326), .Z(n59328) );
  NOR U79680 ( .A(n59328), .B(n59327), .Z(n59329) );
  IV U79681 ( .A(n59329), .Z(n59816) );
  XOR U79682 ( .A(n59815), .B(n59816), .Z(n69717) );
  IV U79683 ( .A(n69717), .Z(n59336) );
  IV U79684 ( .A(n59330), .Z(n59331) );
  NOR U79685 ( .A(n59332), .B(n59331), .Z(n69721) );
  IV U79686 ( .A(n59333), .Z(n59334) );
  NOR U79687 ( .A(n59335), .B(n59334), .Z(n69715) );
  NOR U79688 ( .A(n69721), .B(n69715), .Z(n59811) );
  XOR U79689 ( .A(n59336), .B(n59811), .Z(n59809) );
  XOR U79690 ( .A(n59808), .B(n59809), .Z(n59805) );
  XOR U79691 ( .A(n59337), .B(n59805), .Z(n59800) );
  XOR U79692 ( .A(n59338), .B(n59800), .Z(n64525) );
  XOR U79693 ( .A(n59339), .B(n64525), .Z(n59797) );
  IV U79694 ( .A(n59340), .Z(n59342) );
  NOR U79695 ( .A(n59342), .B(n59341), .Z(n59343) );
  IV U79696 ( .A(n59343), .Z(n59798) );
  XOR U79697 ( .A(n59797), .B(n59798), .Z(n64532) );
  XOR U79698 ( .A(n64531), .B(n64532), .Z(n64541) );
  IV U79699 ( .A(n59344), .Z(n59345) );
  NOR U79700 ( .A(n59346), .B(n59345), .Z(n64534) );
  IV U79701 ( .A(n59347), .Z(n59348) );
  NOR U79702 ( .A(n59351), .B(n59348), .Z(n64540) );
  NOR U79703 ( .A(n64534), .B(n64540), .Z(n59349) );
  XOR U79704 ( .A(n64541), .B(n59349), .Z(n59350) );
  IV U79705 ( .A(n59350), .Z(n64539) );
  NOR U79706 ( .A(n59352), .B(n59351), .Z(n64537) );
  XOR U79707 ( .A(n64539), .B(n64537), .Z(n64544) );
  XOR U79708 ( .A(n64543), .B(n64544), .Z(n64547) );
  XOR U79709 ( .A(n64546), .B(n64547), .Z(n59791) );
  XOR U79710 ( .A(n59353), .B(n59791), .Z(n59783) );
  XOR U79711 ( .A(n59354), .B(n59783), .Z(n64554) );
  XOR U79712 ( .A(n64551), .B(n64554), .Z(n59781) );
  XOR U79713 ( .A(n59355), .B(n59781), .Z(n59771) );
  XOR U79714 ( .A(n59356), .B(n59771), .Z(n64560) );
  XOR U79715 ( .A(n59357), .B(n64560), .Z(n59768) );
  XOR U79716 ( .A(n59358), .B(n59768), .Z(n64566) );
  XOR U79717 ( .A(n64564), .B(n64566), .Z(n59765) );
  XOR U79718 ( .A(n59764), .B(n59765), .Z(n64578) );
  XOR U79719 ( .A(n59359), .B(n64578), .Z(n59757) );
  XOR U79720 ( .A(n59360), .B(n59757), .Z(n59750) );
  XOR U79721 ( .A(n59361), .B(n59750), .Z(n59362) );
  IV U79722 ( .A(n59362), .Z(n59744) );
  XOR U79723 ( .A(n59743), .B(n59744), .Z(n59739) );
  XOR U79724 ( .A(n59738), .B(n59739), .Z(n69819) );
  XOR U79725 ( .A(n59741), .B(n69819), .Z(n64595) );
  IV U79726 ( .A(n59363), .Z(n65052) );
  NOR U79727 ( .A(n65052), .B(n59365), .Z(n59367) );
  IV U79728 ( .A(n59364), .Z(n59366) );
  NOR U79729 ( .A(n59366), .B(n59365), .Z(n69817) );
  NOR U79730 ( .A(n59367), .B(n69817), .Z(n64596) );
  IV U79731 ( .A(n64596), .Z(n59368) );
  NOR U79732 ( .A(n64593), .B(n59368), .Z(n59369) );
  XOR U79733 ( .A(n64595), .B(n59369), .Z(n59370) );
  IV U79734 ( .A(n59370), .Z(n59736) );
  XOR U79735 ( .A(n59735), .B(n59736), .Z(n69826) );
  IV U79736 ( .A(n59371), .Z(n59373) );
  NOR U79737 ( .A(n59373), .B(n59372), .Z(n69824) );
  IV U79738 ( .A(n59374), .Z(n59376) );
  NOR U79739 ( .A(n59376), .B(n59375), .Z(n69829) );
  NOR U79740 ( .A(n69824), .B(n69829), .Z(n64600) );
  XOR U79741 ( .A(n69826), .B(n64600), .Z(n64601) );
  XOR U79742 ( .A(n64603), .B(n64601), .Z(n64607) );
  XOR U79743 ( .A(n64606), .B(n64607), .Z(n65037) );
  XOR U79744 ( .A(n64609), .B(n65037), .Z(n59732) );
  IV U79745 ( .A(n59377), .Z(n59378) );
  NOR U79746 ( .A(n59379), .B(n59378), .Z(n64613) );
  IV U79747 ( .A(n59380), .Z(n59382) );
  NOR U79748 ( .A(n59382), .B(n59381), .Z(n59733) );
  NOR U79749 ( .A(n64613), .B(n59733), .Z(n59383) );
  XOR U79750 ( .A(n59732), .B(n59383), .Z(n64617) );
  XOR U79751 ( .A(n64616), .B(n64617), .Z(n59722) );
  NOR U79752 ( .A(n59384), .B(n59726), .Z(n59391) );
  IV U79753 ( .A(n59385), .Z(n59387) );
  NOR U79754 ( .A(n59387), .B(n59386), .Z(n59721) );
  NOR U79755 ( .A(n59391), .B(n59721), .Z(n59388) );
  XOR U79756 ( .A(n59722), .B(n59388), .Z(n59389) );
  NOR U79757 ( .A(n59390), .B(n59389), .Z(n59394) );
  IV U79758 ( .A(n59390), .Z(n59393) );
  XOR U79759 ( .A(n59391), .B(n59722), .Z(n59392) );
  NOR U79760 ( .A(n59393), .B(n59392), .Z(n69852) );
  NOR U79761 ( .A(n59394), .B(n69852), .Z(n59719) );
  XOR U79762 ( .A(n59395), .B(n59719), .Z(n64626) );
  XOR U79763 ( .A(n64625), .B(n64626), .Z(n64633) );
  IV U79764 ( .A(n59396), .Z(n59398) );
  NOR U79765 ( .A(n59398), .B(n59397), .Z(n64628) );
  IV U79766 ( .A(n59399), .Z(n59400) );
  NOR U79767 ( .A(n59400), .B(n59404), .Z(n64632) );
  NOR U79768 ( .A(n64628), .B(n64632), .Z(n59401) );
  XOR U79769 ( .A(n64633), .B(n59401), .Z(n59402) );
  IV U79770 ( .A(n59402), .Z(n59714) );
  IV U79771 ( .A(n59403), .Z(n59405) );
  NOR U79772 ( .A(n59405), .B(n59404), .Z(n59712) );
  XOR U79773 ( .A(n59714), .B(n59712), .Z(n59717) );
  XOR U79774 ( .A(n59715), .B(n59717), .Z(n64639) );
  XOR U79775 ( .A(n64638), .B(n64639), .Z(n59711) );
  NOR U79776 ( .A(n59412), .B(n59711), .Z(n64649) );
  IV U79777 ( .A(n59406), .Z(n59407) );
  NOR U79778 ( .A(n59408), .B(n59407), .Z(n64655) );
  IV U79779 ( .A(n59409), .Z(n59410) );
  NOR U79780 ( .A(n59411), .B(n59410), .Z(n59709) );
  XOR U79781 ( .A(n59711), .B(n59709), .Z(n64656) );
  IV U79782 ( .A(n64656), .Z(n59413) );
  XOR U79783 ( .A(n64655), .B(n59413), .Z(n59415) );
  NOR U79784 ( .A(n59413), .B(n59412), .Z(n59414) );
  NOR U79785 ( .A(n59415), .B(n59414), .Z(n59416) );
  NOR U79786 ( .A(n64649), .B(n59416), .Z(n59703) );
  XOR U79787 ( .A(n59417), .B(n59703), .Z(n69890) );
  XOR U79788 ( .A(n64662), .B(n69890), .Z(n69895) );
  XOR U79789 ( .A(n64665), .B(n69895), .Z(n59418) );
  IV U79790 ( .A(n59418), .Z(n65001) );
  XOR U79791 ( .A(n64666), .B(n65001), .Z(n64672) );
  XOR U79792 ( .A(n64671), .B(n64672), .Z(n64675) );
  XOR U79793 ( .A(n64674), .B(n64675), .Z(n64679) );
  XOR U79794 ( .A(n64678), .B(n64679), .Z(n64684) );
  IV U79795 ( .A(n59419), .Z(n59420) );
  NOR U79796 ( .A(n59421), .B(n59420), .Z(n64681) );
  IV U79797 ( .A(n59422), .Z(n59423) );
  NOR U79798 ( .A(n59424), .B(n59423), .Z(n64683) );
  NOR U79799 ( .A(n64681), .B(n64683), .Z(n59425) );
  XOR U79800 ( .A(n64684), .B(n59425), .Z(n59426) );
  IV U79801 ( .A(n59426), .Z(n64687) );
  XOR U79802 ( .A(n64686), .B(n64687), .Z(n64694) );
  XOR U79803 ( .A(n64693), .B(n64694), .Z(n59700) );
  XOR U79804 ( .A(n59699), .B(n59700), .Z(n64691) );
  XOR U79805 ( .A(n64690), .B(n64691), .Z(n59697) );
  XOR U79806 ( .A(n59696), .B(n59697), .Z(n64704) );
  XOR U79807 ( .A(n64702), .B(n64704), .Z(n64706) );
  NOR U79808 ( .A(n59433), .B(n64706), .Z(n70097) );
  IV U79809 ( .A(n59427), .Z(n59429) );
  NOR U79810 ( .A(n59429), .B(n59428), .Z(n59692) );
  IV U79811 ( .A(n59430), .Z(n59431) );
  NOR U79812 ( .A(n59432), .B(n59431), .Z(n64705) );
  XOR U79813 ( .A(n64705), .B(n64706), .Z(n59693) );
  IV U79814 ( .A(n59693), .Z(n59434) );
  XOR U79815 ( .A(n59692), .B(n59434), .Z(n59436) );
  NOR U79816 ( .A(n59434), .B(n59433), .Z(n59435) );
  NOR U79817 ( .A(n59436), .B(n59435), .Z(n59437) );
  NOR U79818 ( .A(n70097), .B(n59437), .Z(n64715) );
  IV U79819 ( .A(n59438), .Z(n59440) );
  NOR U79820 ( .A(n59440), .B(n59439), .Z(n64717) );
  IV U79821 ( .A(n59441), .Z(n59443) );
  NOR U79822 ( .A(n59443), .B(n59442), .Z(n64714) );
  NOR U79823 ( .A(n64717), .B(n64714), .Z(n59444) );
  XOR U79824 ( .A(n64715), .B(n59444), .Z(n64712) );
  XOR U79825 ( .A(n64711), .B(n64712), .Z(n59445) );
  NOR U79826 ( .A(n59446), .B(n59445), .Z(n69926) );
  IV U79827 ( .A(n59447), .Z(n59449) );
  NOR U79828 ( .A(n59449), .B(n59448), .Z(n59690) );
  NOR U79829 ( .A(n64711), .B(n59690), .Z(n59450) );
  XOR U79830 ( .A(n59450), .B(n64712), .Z(n69924) );
  NOR U79831 ( .A(n59451), .B(n69924), .Z(n59452) );
  NOR U79832 ( .A(n69926), .B(n59452), .Z(n64723) );
  XOR U79833 ( .A(n64725), .B(n64723), .Z(n64733) );
  IV U79834 ( .A(n59453), .Z(n59454) );
  NOR U79835 ( .A(n59454), .B(n69941), .Z(n59455) );
  IV U79836 ( .A(n59455), .Z(n59456) );
  NOR U79837 ( .A(n59457), .B(n59456), .Z(n64731) );
  XOR U79838 ( .A(n64733), .B(n64731), .Z(n59687) );
  XOR U79839 ( .A(n59686), .B(n59687), .Z(n64729) );
  XOR U79840 ( .A(n64728), .B(n64729), .Z(n59683) );
  IV U79841 ( .A(n59458), .Z(n59462) );
  XOR U79842 ( .A(n59460), .B(n59459), .Z(n59461) );
  NOR U79843 ( .A(n59462), .B(n59461), .Z(n59681) );
  XOR U79844 ( .A(n59683), .B(n59681), .Z(n64744) );
  IV U79845 ( .A(n59463), .Z(n59464) );
  NOR U79846 ( .A(n59465), .B(n59464), .Z(n64743) );
  IV U79847 ( .A(n59466), .Z(n59469) );
  IV U79848 ( .A(n59467), .Z(n59468) );
  NOR U79849 ( .A(n59469), .B(n59468), .Z(n59684) );
  NOR U79850 ( .A(n64743), .B(n59684), .Z(n59470) );
  XOR U79851 ( .A(n64744), .B(n59470), .Z(n59471) );
  IV U79852 ( .A(n59471), .Z(n64742) );
  IV U79853 ( .A(n59472), .Z(n59473) );
  NOR U79854 ( .A(n59474), .B(n59473), .Z(n59475) );
  IV U79855 ( .A(n59475), .Z(n59487) );
  NOR U79856 ( .A(n64742), .B(n59487), .Z(n64950) );
  IV U79857 ( .A(n59476), .Z(n59478) );
  NOR U79858 ( .A(n59478), .B(n59477), .Z(n64750) );
  IV U79859 ( .A(n59479), .Z(n59483) );
  NOR U79860 ( .A(n59481), .B(n59480), .Z(n59482) );
  IV U79861 ( .A(n59482), .Z(n59485) );
  NOR U79862 ( .A(n59483), .B(n59485), .Z(n64740) );
  XOR U79863 ( .A(n64740), .B(n64742), .Z(n59679) );
  IV U79864 ( .A(n59484), .Z(n59486) );
  NOR U79865 ( .A(n59486), .B(n59485), .Z(n59677) );
  XOR U79866 ( .A(n59679), .B(n59677), .Z(n64751) );
  IV U79867 ( .A(n64751), .Z(n59488) );
  XOR U79868 ( .A(n64750), .B(n59488), .Z(n59490) );
  NOR U79869 ( .A(n59488), .B(n59487), .Z(n59489) );
  NOR U79870 ( .A(n59490), .B(n59489), .Z(n59491) );
  NOR U79871 ( .A(n64950), .B(n59491), .Z(n64748) );
  XOR U79872 ( .A(n64754), .B(n64748), .Z(n64760) );
  IV U79873 ( .A(n59492), .Z(n59494) );
  NOR U79874 ( .A(n59494), .B(n59493), .Z(n64747) );
  IV U79875 ( .A(n59495), .Z(n59496) );
  NOR U79876 ( .A(n59497), .B(n59496), .Z(n64759) );
  NOR U79877 ( .A(n64747), .B(n64759), .Z(n59498) );
  XOR U79878 ( .A(n64760), .B(n59498), .Z(n59499) );
  IV U79879 ( .A(n59499), .Z(n64764) );
  IV U79880 ( .A(n59500), .Z(n59502) );
  NOR U79881 ( .A(n59502), .B(n59501), .Z(n64762) );
  XOR U79882 ( .A(n64764), .B(n64762), .Z(n64766) );
  XOR U79883 ( .A(n64765), .B(n64766), .Z(n64772) );
  XOR U79884 ( .A(n64769), .B(n64772), .Z(n59507) );
  IV U79885 ( .A(n59503), .Z(n59505) );
  NOR U79886 ( .A(n59505), .B(n59504), .Z(n59513) );
  IV U79887 ( .A(n59513), .Z(n59506) );
  NOR U79888 ( .A(n59507), .B(n59506), .Z(n64935) );
  IV U79889 ( .A(n59508), .Z(n59509) );
  NOR U79890 ( .A(n59510), .B(n59509), .Z(n64771) );
  NOR U79891 ( .A(n64769), .B(n64771), .Z(n59511) );
  XOR U79892 ( .A(n64772), .B(n59511), .Z(n59512) );
  NOR U79893 ( .A(n59513), .B(n59512), .Z(n59514) );
  NOR U79894 ( .A(n64935), .B(n59514), .Z(n59515) );
  IV U79895 ( .A(n59515), .Z(n64776) );
  XOR U79896 ( .A(n64775), .B(n64776), .Z(n64923) );
  IV U79897 ( .A(n64923), .Z(n59522) );
  IV U79898 ( .A(n59516), .Z(n59518) );
  NOR U79899 ( .A(n59518), .B(n59517), .Z(n64927) );
  IV U79900 ( .A(n59519), .Z(n59521) );
  NOR U79901 ( .A(n59521), .B(n59520), .Z(n64922) );
  NOR U79902 ( .A(n64927), .B(n64922), .Z(n64779) );
  XOR U79903 ( .A(n59522), .B(n64779), .Z(n64782) );
  XOR U79904 ( .A(n64780), .B(n64782), .Z(n64913) );
  XOR U79905 ( .A(n59523), .B(n64913), .Z(n64791) );
  IV U79906 ( .A(n59524), .Z(n59525) );
  NOR U79907 ( .A(n59526), .B(n59525), .Z(n64785) );
  IV U79908 ( .A(n59527), .Z(n59528) );
  NOR U79909 ( .A(n59529), .B(n59528), .Z(n64790) );
  NOR U79910 ( .A(n64785), .B(n64790), .Z(n59530) );
  XOR U79911 ( .A(n64791), .B(n59530), .Z(n59674) );
  IV U79912 ( .A(n59531), .Z(n59533) );
  NOR U79913 ( .A(n59533), .B(n59532), .Z(n59675) );
  IV U79914 ( .A(n59534), .Z(n59535) );
  NOR U79915 ( .A(n59536), .B(n59535), .Z(n64796) );
  NOR U79916 ( .A(n59675), .B(n64796), .Z(n59537) );
  XOR U79917 ( .A(n59674), .B(n59537), .Z(n59671) );
  XOR U79918 ( .A(n59670), .B(n59671), .Z(n64794) );
  IV U79919 ( .A(n59538), .Z(n59540) );
  NOR U79920 ( .A(n59540), .B(n59539), .Z(n64793) );
  NOR U79921 ( .A(n64793), .B(n59668), .Z(n59541) );
  XOR U79922 ( .A(n64794), .B(n59541), .Z(n59542) );
  IV U79923 ( .A(n59542), .Z(n64806) );
  XOR U79924 ( .A(n64805), .B(n64806), .Z(n64810) );
  XOR U79925 ( .A(n64808), .B(n64810), .Z(n64821) );
  XOR U79926 ( .A(n64820), .B(n64821), .Z(n64814) );
  XOR U79927 ( .A(n64813), .B(n64814), .Z(n64818) );
  XOR U79928 ( .A(n64817), .B(n64818), .Z(n59666) );
  NOR U79929 ( .A(n59550), .B(n59666), .Z(n64883) );
  IV U79930 ( .A(n59574), .Z(n59543) );
  NOR U79931 ( .A(n59544), .B(n59543), .Z(n59558) );
  IV U79932 ( .A(n59558), .Z(n59545) );
  NOR U79933 ( .A(n59546), .B(n59545), .Z(n64829) );
  IV U79934 ( .A(n59547), .Z(n59548) );
  NOR U79935 ( .A(n59549), .B(n59548), .Z(n59665) );
  XOR U79936 ( .A(n59665), .B(n59666), .Z(n64830) );
  IV U79937 ( .A(n64830), .Z(n59551) );
  XOR U79938 ( .A(n64829), .B(n59551), .Z(n59553) );
  NOR U79939 ( .A(n59551), .B(n59550), .Z(n59552) );
  NOR U79940 ( .A(n59553), .B(n59552), .Z(n59554) );
  NOR U79941 ( .A(n64883), .B(n59554), .Z(n59555) );
  IV U79942 ( .A(n59555), .Z(n64833) );
  XOR U79943 ( .A(n64832), .B(n64833), .Z(n59591) );
  IV U79944 ( .A(n59591), .Z(n59589) );
  IV U79945 ( .A(n59556), .Z(n59560) );
  NOR U79946 ( .A(n59558), .B(n59557), .Z(n59559) );
  XOR U79947 ( .A(n59560), .B(n59559), .Z(n59593) );
  IV U79948 ( .A(n59561), .Z(n59563) );
  NOR U79949 ( .A(n59563), .B(n59562), .Z(n69991) );
  NOR U79950 ( .A(n59565), .B(n59564), .Z(n59566) );
  NOR U79951 ( .A(n69991), .B(n59566), .Z(n59578) );
  XOR U79952 ( .A(n59568), .B(n59567), .Z(n59572) );
  NOR U79953 ( .A(n59570), .B(n59569), .Z(n59571) );
  NOR U79954 ( .A(n59572), .B(n59571), .Z(n59573) );
  NOR U79955 ( .A(n59574), .B(n59573), .Z(n59577) );
  IV U79956 ( .A(n59577), .Z(n69999) );
  NOR U79957 ( .A(n59578), .B(n69999), .Z(n59598) );
  IV U79958 ( .A(n59598), .Z(n59575) );
  NOR U79959 ( .A(n69988), .B(n59575), .Z(n59576) );
  IV U79960 ( .A(n59576), .Z(n59595) );
  NOR U79961 ( .A(n59593), .B(n59595), .Z(n59586) );
  XOR U79962 ( .A(n59593), .B(n59576), .Z(n59612) );
  XOR U79963 ( .A(n59578), .B(n59577), .Z(n59616) );
  IV U79964 ( .A(n59579), .Z(n59580) );
  NOR U79965 ( .A(n59581), .B(n59580), .Z(n59614) );
  IV U79966 ( .A(n59614), .Z(n59582) );
  NOR U79967 ( .A(n59616), .B(n59582), .Z(n59602) );
  IV U79968 ( .A(n59602), .Z(n59584) );
  XOR U79969 ( .A(n59599), .B(n69988), .Z(n59583) );
  NOR U79970 ( .A(n59584), .B(n59583), .Z(n59610) );
  IV U79971 ( .A(n59610), .Z(n59585) );
  NOR U79972 ( .A(n59612), .B(n59585), .Z(n59590) );
  NOR U79973 ( .A(n59586), .B(n59590), .Z(n59587) );
  IV U79974 ( .A(n59587), .Z(n59588) );
  NOR U79975 ( .A(n59589), .B(n59588), .Z(n59597) );
  IV U79976 ( .A(n59590), .Z(n59592) );
  NOR U79977 ( .A(n59592), .B(n59591), .Z(n64876) );
  NOR U79978 ( .A(n59593), .B(n64833), .Z(n59594) );
  IV U79979 ( .A(n59594), .Z(n69993) );
  NOR U79980 ( .A(n59595), .B(n69993), .Z(n64879) );
  NOR U79981 ( .A(n64876), .B(n64879), .Z(n59596) );
  IV U79982 ( .A(n59596), .Z(n59664) );
  NOR U79983 ( .A(n59597), .B(n59664), .Z(n59659) );
  NOR U79984 ( .A(n59599), .B(n59598), .Z(n59600) );
  XOR U79985 ( .A(n59600), .B(n69988), .Z(n59601) );
  NOR U79986 ( .A(n59602), .B(n59601), .Z(n59603) );
  NOR U79987 ( .A(n59610), .B(n59603), .Z(n59637) );
  IV U79988 ( .A(n59637), .Z(n59622) );
  IV U79989 ( .A(n59604), .Z(n59606) );
  NOR U79990 ( .A(n59606), .B(n59605), .Z(n59613) );
  IV U79991 ( .A(n59613), .Z(n59607) );
  NOR U79992 ( .A(n59616), .B(n59607), .Z(n59635) );
  IV U79993 ( .A(n59635), .Z(n59629) );
  NOR U79994 ( .A(n59622), .B(n59629), .Z(n59609) );
  IV U79995 ( .A(n59609), .Z(n59608) );
  NOR U79996 ( .A(n59612), .B(n59608), .Z(n59661) );
  NOR U79997 ( .A(n59610), .B(n59609), .Z(n59611) );
  XOR U79998 ( .A(n59612), .B(n59611), .Z(n59642) );
  IV U79999 ( .A(n59642), .Z(n59633) );
  NOR U80000 ( .A(n59614), .B(n59613), .Z(n59615) );
  XOR U80001 ( .A(n59616), .B(n59615), .Z(n59646) );
  IV U80002 ( .A(n59646), .Z(n59628) );
  IV U80003 ( .A(n59617), .Z(n59619) );
  NOR U80004 ( .A(n59619), .B(n59618), .Z(n59644) );
  IV U80005 ( .A(n59644), .Z(n59620) );
  NOR U80006 ( .A(n59628), .B(n59620), .Z(n59634) );
  IV U80007 ( .A(n59634), .Z(n59621) );
  NOR U80008 ( .A(n59622), .B(n59621), .Z(n59640) );
  IV U80009 ( .A(n59640), .Z(n59623) );
  NOR U80010 ( .A(n59633), .B(n59623), .Z(n59658) );
  NOR U80011 ( .A(n59661), .B(n59658), .Z(n59624) );
  XOR U80012 ( .A(n59659), .B(n59624), .Z(n59657) );
  NOR U80013 ( .A(n59626), .B(n59625), .Z(n59643) );
  IV U80014 ( .A(n59643), .Z(n59627) );
  NOR U80015 ( .A(n59628), .B(n59627), .Z(n70010) );
  IV U80016 ( .A(n70010), .Z(n59638) );
  XOR U80017 ( .A(n59637), .B(n59629), .Z(n59630) );
  NOR U80018 ( .A(n59638), .B(n59630), .Z(n59631) );
  IV U80019 ( .A(n59631), .Z(n59632) );
  NOR U80020 ( .A(n59633), .B(n59632), .Z(n59655) );
  XOR U80021 ( .A(n59657), .B(n59655), .Z(n64856) );
  NOR U80022 ( .A(n59635), .B(n59634), .Z(n59636) );
  XOR U80023 ( .A(n59637), .B(n59636), .Z(n70012) );
  NOR U80024 ( .A(n59638), .B(n70012), .Z(n59639) );
  NOR U80025 ( .A(n59640), .B(n59639), .Z(n59641) );
  XOR U80026 ( .A(n59642), .B(n59641), .Z(n64847) );
  NOR U80027 ( .A(n59644), .B(n59643), .Z(n59645) );
  XOR U80028 ( .A(n59646), .B(n59645), .Z(n64838) );
  IV U80029 ( .A(n59647), .Z(n59648) );
  NOR U80030 ( .A(n59649), .B(n59648), .Z(n64839) );
  IV U80031 ( .A(n64839), .Z(n59650) );
  NOR U80032 ( .A(n64838), .B(n59650), .Z(n70009) );
  IV U80033 ( .A(n70009), .Z(n59651) );
  NOR U80034 ( .A(n70012), .B(n59651), .Z(n64846) );
  IV U80035 ( .A(n64846), .Z(n59652) );
  NOR U80036 ( .A(n64847), .B(n59652), .Z(n64854) );
  IV U80037 ( .A(n64854), .Z(n59653) );
  NOR U80038 ( .A(n64856), .B(n59653), .Z(n59654) );
  IV U80039 ( .A(n59654), .Z(n64868) );
  IV U80040 ( .A(n59655), .Z(n59656) );
  NOR U80041 ( .A(n59657), .B(n59656), .Z(n70001) );
  IV U80042 ( .A(n59658), .Z(n59660) );
  IV U80043 ( .A(n59659), .Z(n59662) );
  NOR U80044 ( .A(n59660), .B(n59662), .Z(n64870) );
  NOR U80045 ( .A(n70001), .B(n64870), .Z(n64837) );
  IV U80046 ( .A(n59661), .Z(n59663) );
  NOR U80047 ( .A(n59663), .B(n59662), .Z(n64873) );
  NOR U80048 ( .A(n59664), .B(n64873), .Z(n64836) );
  IV U80049 ( .A(n59665), .Z(n59667) );
  NOR U80050 ( .A(n59667), .B(n59666), .Z(n69977) );
  IV U80051 ( .A(n59668), .Z(n59669) );
  NOR U80052 ( .A(n59669), .B(n64794), .Z(n64890) );
  IV U80053 ( .A(n59670), .Z(n59672) );
  NOR U80054 ( .A(n59672), .B(n59671), .Z(n59673) );
  IV U80055 ( .A(n59673), .Z(n64799) );
  IV U80056 ( .A(n59674), .Z(n64798) );
  IV U80057 ( .A(n59675), .Z(n59676) );
  NOR U80058 ( .A(n64798), .B(n59676), .Z(n64898) );
  IV U80059 ( .A(n59677), .Z(n59678) );
  NOR U80060 ( .A(n59679), .B(n59678), .Z(n59680) );
  IV U80061 ( .A(n59680), .Z(n64949) );
  IV U80062 ( .A(n59681), .Z(n59682) );
  NOR U80063 ( .A(n59683), .B(n59682), .Z(n69943) );
  IV U80064 ( .A(n59684), .Z(n59685) );
  NOR U80065 ( .A(n64744), .B(n59685), .Z(n69950) );
  NOR U80066 ( .A(n69943), .B(n69950), .Z(n64739) );
  IV U80067 ( .A(n59686), .Z(n59688) );
  NOR U80068 ( .A(n59688), .B(n59687), .Z(n59689) );
  IV U80069 ( .A(n59689), .Z(n64734) );
  IV U80070 ( .A(n59690), .Z(n59691) );
  NOR U80071 ( .A(n59691), .B(n64712), .Z(n69912) );
  IV U80072 ( .A(n59692), .Z(n59694) );
  NOR U80073 ( .A(n59694), .B(n59693), .Z(n59695) );
  IV U80074 ( .A(n59695), .Z(n64971) );
  IV U80075 ( .A(n59696), .Z(n59698) );
  NOR U80076 ( .A(n59698), .B(n59697), .Z(n64976) );
  IV U80077 ( .A(n59699), .Z(n59701) );
  NOR U80078 ( .A(n59701), .B(n59700), .Z(n59702) );
  IV U80079 ( .A(n59702), .Z(n64696) );
  IV U80080 ( .A(n59706), .Z(n59704) );
  IV U80081 ( .A(n59703), .Z(n64660) );
  NOR U80082 ( .A(n59704), .B(n64660), .Z(n69877) );
  IV U80083 ( .A(n59705), .Z(n59708) );
  XOR U80084 ( .A(n59706), .B(n64660), .Z(n59707) );
  NOR U80085 ( .A(n59708), .B(n59707), .Z(n65013) );
  NOR U80086 ( .A(n69877), .B(n65013), .Z(n64658) );
  IV U80087 ( .A(n59709), .Z(n59710) );
  NOR U80088 ( .A(n59711), .B(n59710), .Z(n64646) );
  IV U80089 ( .A(n64646), .Z(n64637) );
  IV U80090 ( .A(n59712), .Z(n59713) );
  NOR U80091 ( .A(n59714), .B(n59713), .Z(n69860) );
  IV U80092 ( .A(n59715), .Z(n59716) );
  NOR U80093 ( .A(n59717), .B(n59716), .Z(n69865) );
  NOR U80094 ( .A(n69860), .B(n69865), .Z(n64635) );
  IV U80095 ( .A(n59718), .Z(n59720) );
  IV U80096 ( .A(n59719), .Z(n64623) );
  NOR U80097 ( .A(n59720), .B(n64623), .Z(n65019) );
  IV U80098 ( .A(n59721), .Z(n59723) );
  NOR U80099 ( .A(n59723), .B(n59722), .Z(n59724) );
  IV U80100 ( .A(n59724), .Z(n69851) );
  IV U80101 ( .A(n59725), .Z(n59728) );
  NOR U80102 ( .A(n59726), .B(n64617), .Z(n59727) );
  IV U80103 ( .A(n59727), .Z(n59730) );
  NOR U80104 ( .A(n59728), .B(n59730), .Z(n69839) );
  IV U80105 ( .A(n59729), .Z(n59731) );
  NOR U80106 ( .A(n59731), .B(n59730), .Z(n65027) );
  IV U80107 ( .A(n59732), .Z(n64614) );
  IV U80108 ( .A(n59733), .Z(n59734) );
  NOR U80109 ( .A(n64614), .B(n59734), .Z(n65033) );
  IV U80110 ( .A(n59735), .Z(n59737) );
  NOR U80111 ( .A(n59737), .B(n59736), .Z(n64598) );
  IV U80112 ( .A(n64598), .Z(n64592) );
  IV U80113 ( .A(n59738), .Z(n59740) );
  NOR U80114 ( .A(n59740), .B(n59739), .Z(n69805) );
  IV U80115 ( .A(n59741), .Z(n59742) );
  NOR U80116 ( .A(n59742), .B(n69819), .Z(n69814) );
  NOR U80117 ( .A(n69805), .B(n69814), .Z(n64591) );
  IV U80118 ( .A(n59743), .Z(n59745) );
  NOR U80119 ( .A(n59745), .B(n59744), .Z(n69809) );
  IV U80120 ( .A(n59746), .Z(n59747) );
  NOR U80121 ( .A(n59750), .B(n59747), .Z(n69807) );
  NOR U80122 ( .A(n69809), .B(n69807), .Z(n64590) );
  IV U80123 ( .A(n59748), .Z(n59755) );
  NOR U80124 ( .A(n59750), .B(n59749), .Z(n59751) );
  IV U80125 ( .A(n59751), .Z(n59752) );
  NOR U80126 ( .A(n59753), .B(n59752), .Z(n59754) );
  IV U80127 ( .A(n59754), .Z(n59762) );
  NOR U80128 ( .A(n59755), .B(n59762), .Z(n69799) );
  IV U80129 ( .A(n59756), .Z(n59760) );
  IV U80130 ( .A(n59757), .Z(n64582) );
  NOR U80131 ( .A(n64582), .B(n59758), .Z(n59759) );
  IV U80132 ( .A(n59759), .Z(n64587) );
  NOR U80133 ( .A(n59760), .B(n64587), .Z(n70147) );
  IV U80134 ( .A(n59761), .Z(n59763) );
  NOR U80135 ( .A(n59763), .B(n59762), .Z(n75053) );
  NOR U80136 ( .A(n70147), .B(n75053), .Z(n69798) );
  IV U80137 ( .A(n59764), .Z(n59766) );
  NOR U80138 ( .A(n59766), .B(n59765), .Z(n59767) );
  IV U80139 ( .A(n59767), .Z(n64571) );
  IV U80140 ( .A(n59768), .Z(n70178) );
  IV U80141 ( .A(n59769), .Z(n59770) );
  NOR U80142 ( .A(n70178), .B(n59770), .Z(n65067) );
  IV U80143 ( .A(n59771), .Z(n59778) );
  IV U80144 ( .A(n59772), .Z(n59773) );
  NOR U80145 ( .A(n59778), .B(n59773), .Z(n75020) );
  IV U80146 ( .A(n59774), .Z(n59775) );
  NOR U80147 ( .A(n59775), .B(n64560), .Z(n70179) );
  NOR U80148 ( .A(n75020), .B(n70179), .Z(n65069) );
  IV U80149 ( .A(n59776), .Z(n59777) );
  NOR U80150 ( .A(n59778), .B(n59777), .Z(n69774) );
  IV U80151 ( .A(n59779), .Z(n59780) );
  NOR U80152 ( .A(n59781), .B(n59780), .Z(n59782) );
  IV U80153 ( .A(n59782), .Z(n69772) );
  IV U80154 ( .A(n59783), .Z(n59789) );
  IV U80155 ( .A(n59784), .Z(n59785) );
  NOR U80156 ( .A(n59789), .B(n59785), .Z(n59786) );
  IV U80157 ( .A(n59786), .Z(n65073) );
  IV U80158 ( .A(n59787), .Z(n59788) );
  NOR U80159 ( .A(n59789), .B(n59788), .Z(n65078) );
  IV U80160 ( .A(n59790), .Z(n59792) );
  NOR U80161 ( .A(n59792), .B(n59791), .Z(n69766) );
  NOR U80162 ( .A(n65078), .B(n69766), .Z(n64550) );
  IV U80163 ( .A(n59793), .Z(n59794) );
  NOR U80164 ( .A(n59794), .B(n64547), .Z(n69762) );
  IV U80165 ( .A(n59795), .Z(n59796) );
  NOR U80166 ( .A(n64525), .B(n59796), .Z(n69731) );
  IV U80167 ( .A(n59797), .Z(n59799) );
  NOR U80168 ( .A(n59799), .B(n59798), .Z(n65082) );
  NOR U80169 ( .A(n69731), .B(n65082), .Z(n64530) );
  IV U80170 ( .A(n59800), .Z(n64528) );
  IV U80171 ( .A(n59801), .Z(n59802) );
  NOR U80172 ( .A(n64528), .B(n59802), .Z(n69727) );
  IV U80173 ( .A(n59803), .Z(n59804) );
  NOR U80174 ( .A(n59805), .B(n59804), .Z(n69724) );
  IV U80175 ( .A(n59806), .Z(n59807) );
  NOR U80176 ( .A(n59807), .B(n59809), .Z(n65085) );
  IV U80177 ( .A(n59808), .Z(n59810) );
  NOR U80178 ( .A(n59810), .B(n59809), .Z(n65087) );
  NOR U80179 ( .A(n59811), .B(n69717), .Z(n59812) );
  NOR U80180 ( .A(n65087), .B(n59812), .Z(n59813) );
  IV U80181 ( .A(n59813), .Z(n59814) );
  NOR U80182 ( .A(n65085), .B(n59814), .Z(n64521) );
  IV U80183 ( .A(n59815), .Z(n59817) );
  NOR U80184 ( .A(n59817), .B(n59816), .Z(n65093) );
  IV U80185 ( .A(n59818), .Z(n59820) );
  NOR U80186 ( .A(n59820), .B(n59819), .Z(n65090) );
  IV U80187 ( .A(n59821), .Z(n59822) );
  NOR U80188 ( .A(n59833), .B(n59822), .Z(n65106) );
  IV U80189 ( .A(n59823), .Z(n59830) );
  NOR U80190 ( .A(n59825), .B(n59824), .Z(n59826) );
  IV U80191 ( .A(n59826), .Z(n59827) );
  NOR U80192 ( .A(n59828), .B(n59827), .Z(n59829) );
  IV U80193 ( .A(n59829), .Z(n64518) );
  NOR U80194 ( .A(n59830), .B(n64518), .Z(n65098) );
  NOR U80195 ( .A(n65106), .B(n65098), .Z(n64514) );
  IV U80196 ( .A(n59831), .Z(n59835) );
  NOR U80197 ( .A(n59833), .B(n59832), .Z(n59834) );
  IV U80198 ( .A(n59834), .Z(n59837) );
  NOR U80199 ( .A(n59835), .B(n59837), .Z(n65103) );
  IV U80200 ( .A(n59836), .Z(n59838) );
  NOR U80201 ( .A(n59838), .B(n59837), .Z(n69709) );
  IV U80202 ( .A(n59839), .Z(n59843) );
  NOR U80203 ( .A(n59841), .B(n59840), .Z(n59842) );
  IV U80204 ( .A(n59842), .Z(n64503) );
  NOR U80205 ( .A(n59843), .B(n64503), .Z(n69693) );
  IV U80206 ( .A(n59844), .Z(n59846) );
  NOR U80207 ( .A(n59846), .B(n59845), .Z(n69690) );
  NOR U80208 ( .A(n65116), .B(n65120), .Z(n59847) );
  NOR U80209 ( .A(n65121), .B(n59847), .Z(n64501) );
  IV U80210 ( .A(n59848), .Z(n59850) );
  NOR U80211 ( .A(n59850), .B(n59849), .Z(n65126) );
  IV U80212 ( .A(n59851), .Z(n59858) );
  IV U80213 ( .A(n59852), .Z(n59853) );
  NOR U80214 ( .A(n59858), .B(n59853), .Z(n65129) );
  NOR U80215 ( .A(n65126), .B(n65129), .Z(n64499) );
  IV U80216 ( .A(n59854), .Z(n59855) );
  NOR U80217 ( .A(n59858), .B(n59855), .Z(n65131) );
  IV U80218 ( .A(n59856), .Z(n59857) );
  NOR U80219 ( .A(n59858), .B(n59857), .Z(n65134) );
  IV U80220 ( .A(n59859), .Z(n59860) );
  NOR U80221 ( .A(n59860), .B(n59865), .Z(n59861) );
  IV U80222 ( .A(n59861), .Z(n65142) );
  IV U80223 ( .A(n59862), .Z(n65148) );
  NOR U80224 ( .A(n59863), .B(n65148), .Z(n59867) );
  IV U80225 ( .A(n59864), .Z(n59866) );
  NOR U80226 ( .A(n59866), .B(n59865), .Z(n65144) );
  NOR U80227 ( .A(n59867), .B(n65144), .Z(n64482) );
  IV U80228 ( .A(n59868), .Z(n59869) );
  NOR U80229 ( .A(n59872), .B(n59869), .Z(n69661) );
  IV U80230 ( .A(n59870), .Z(n59871) );
  NOR U80231 ( .A(n59872), .B(n59871), .Z(n65154) );
  NOR U80232 ( .A(n59873), .B(n65159), .Z(n65151) );
  NOR U80233 ( .A(n65159), .B(n59874), .Z(n64481) );
  IV U80234 ( .A(n59875), .Z(n59877) );
  NOR U80235 ( .A(n59877), .B(n59876), .Z(n69653) );
  IV U80236 ( .A(n59878), .Z(n59879) );
  NOR U80237 ( .A(n59879), .B(n59889), .Z(n59880) );
  IV U80238 ( .A(n59880), .Z(n69637) );
  IV U80239 ( .A(n59881), .Z(n59886) );
  IV U80240 ( .A(n59882), .Z(n59883) );
  NOR U80241 ( .A(n59886), .B(n59883), .Z(n69629) );
  IV U80242 ( .A(n59884), .Z(n59885) );
  NOR U80243 ( .A(n59886), .B(n59885), .Z(n65176) );
  NOR U80244 ( .A(n69629), .B(n65176), .Z(n59887) );
  IV U80245 ( .A(n59887), .Z(n59891) );
  IV U80246 ( .A(n59888), .Z(n59890) );
  NOR U80247 ( .A(n59890), .B(n59889), .Z(n69627) );
  NOR U80248 ( .A(n59891), .B(n69627), .Z(n64466) );
  IV U80249 ( .A(n59892), .Z(n64449) );
  IV U80250 ( .A(n59893), .Z(n59894) );
  NOR U80251 ( .A(n59894), .B(n64449), .Z(n59895) );
  IV U80252 ( .A(n59895), .Z(n65186) );
  IV U80253 ( .A(n59896), .Z(n59897) );
  NOR U80254 ( .A(n59897), .B(n59899), .Z(n69613) );
  IV U80255 ( .A(n59898), .Z(n59900) );
  NOR U80256 ( .A(n59900), .B(n59899), .Z(n65188) );
  IV U80257 ( .A(n59901), .Z(n59902) );
  NOR U80258 ( .A(n64402), .B(n59902), .Z(n65198) );
  IV U80259 ( .A(n59903), .Z(n59906) );
  NOR U80260 ( .A(n59904), .B(n59911), .Z(n59905) );
  IV U80261 ( .A(n59905), .Z(n59908) );
  NOR U80262 ( .A(n59906), .B(n59908), .Z(n65204) );
  IV U80263 ( .A(n59907), .Z(n59909) );
  NOR U80264 ( .A(n59909), .B(n59908), .Z(n65201) );
  IV U80265 ( .A(n59910), .Z(n59912) );
  NOR U80266 ( .A(n59912), .B(n59911), .Z(n65211) );
  IV U80267 ( .A(n59913), .Z(n59915) );
  IV U80268 ( .A(n59914), .Z(n59917) );
  NOR U80269 ( .A(n59915), .B(n59917), .Z(n65208) );
  IV U80270 ( .A(n59916), .Z(n59918) );
  NOR U80271 ( .A(n59918), .B(n59917), .Z(n65217) );
  IV U80272 ( .A(n59919), .Z(n59920) );
  NOR U80273 ( .A(n59920), .B(n64397), .Z(n65214) );
  IV U80274 ( .A(n59921), .Z(n59922) );
  NOR U80275 ( .A(n59923), .B(n59922), .Z(n59924) );
  IV U80276 ( .A(n59924), .Z(n64391) );
  IV U80277 ( .A(n59925), .Z(n59927) );
  NOR U80278 ( .A(n59927), .B(n59926), .Z(n65225) );
  IV U80279 ( .A(n59928), .Z(n59930) );
  NOR U80280 ( .A(n59930), .B(n59929), .Z(n65220) );
  NOR U80281 ( .A(n65225), .B(n65220), .Z(n64383) );
  IV U80282 ( .A(n59931), .Z(n59933) );
  NOR U80283 ( .A(n59933), .B(n59932), .Z(n69570) );
  IV U80284 ( .A(n59934), .Z(n59935) );
  NOR U80285 ( .A(n59936), .B(n59935), .Z(n65222) );
  NOR U80286 ( .A(n69570), .B(n65222), .Z(n64382) );
  IV U80287 ( .A(n59937), .Z(n59939) );
  NOR U80288 ( .A(n59939), .B(n59938), .Z(n69555) );
  IV U80289 ( .A(n59940), .Z(n59941) );
  NOR U80290 ( .A(n59942), .B(n59941), .Z(n69549) );
  IV U80291 ( .A(n59943), .Z(n59945) );
  NOR U80292 ( .A(n59945), .B(n59944), .Z(n65233) );
  NOR U80293 ( .A(n69549), .B(n65233), .Z(n64368) );
  IV U80294 ( .A(n59946), .Z(n59949) );
  NOR U80295 ( .A(n59947), .B(n59951), .Z(n59948) );
  IV U80296 ( .A(n59948), .Z(n59954) );
  NOR U80297 ( .A(n59949), .B(n59954), .Z(n65230) );
  IV U80298 ( .A(n59950), .Z(n59952) );
  NOR U80299 ( .A(n59952), .B(n59951), .Z(n65237) );
  IV U80300 ( .A(n59953), .Z(n59955) );
  NOR U80301 ( .A(n59955), .B(n59954), .Z(n65235) );
  NOR U80302 ( .A(n65237), .B(n65235), .Z(n59956) );
  IV U80303 ( .A(n59956), .Z(n64367) );
  IV U80304 ( .A(n59957), .Z(n59959) );
  NOR U80305 ( .A(n59959), .B(n59958), .Z(n65240) );
  IV U80306 ( .A(n59960), .Z(n59965) );
  IV U80307 ( .A(n59961), .Z(n59962) );
  NOR U80308 ( .A(n59965), .B(n59962), .Z(n65242) );
  NOR U80309 ( .A(n65240), .B(n65242), .Z(n64366) );
  IV U80310 ( .A(n59963), .Z(n59964) );
  NOR U80311 ( .A(n59965), .B(n59964), .Z(n59966) );
  IV U80312 ( .A(n59966), .Z(n65245) );
  IV U80313 ( .A(n59967), .Z(n59968) );
  NOR U80314 ( .A(n59968), .B(n64363), .Z(n69545) );
  IV U80315 ( .A(n59969), .Z(n59970) );
  NOR U80316 ( .A(n59970), .B(n59976), .Z(n70361) );
  IV U80317 ( .A(n59971), .Z(n59973) );
  IV U80318 ( .A(n59972), .Z(n64359) );
  NOR U80319 ( .A(n59973), .B(n64359), .Z(n70356) );
  NOR U80320 ( .A(n70361), .B(n70356), .Z(n65251) );
  IV U80321 ( .A(n59974), .Z(n59975) );
  NOR U80322 ( .A(n59976), .B(n59975), .Z(n59977) );
  IV U80323 ( .A(n59977), .Z(n65256) );
  IV U80324 ( .A(n59978), .Z(n59980) );
  NOR U80325 ( .A(n59980), .B(n59979), .Z(n65258) );
  IV U80326 ( .A(n59981), .Z(n59983) );
  NOR U80327 ( .A(n59983), .B(n59982), .Z(n65252) );
  NOR U80328 ( .A(n65258), .B(n65252), .Z(n64354) );
  IV U80329 ( .A(n59984), .Z(n59985) );
  NOR U80330 ( .A(n59985), .B(n64351), .Z(n69530) );
  IV U80331 ( .A(n59986), .Z(n59987) );
  NOR U80332 ( .A(n59988), .B(n59987), .Z(n69534) );
  NOR U80333 ( .A(n69530), .B(n69534), .Z(n64353) );
  IV U80334 ( .A(n59989), .Z(n64348) );
  IV U80335 ( .A(n59990), .Z(n59991) );
  NOR U80336 ( .A(n64348), .B(n59991), .Z(n65263) );
  IV U80337 ( .A(n59992), .Z(n59993) );
  NOR U80338 ( .A(n59994), .B(n59993), .Z(n64333) );
  IV U80339 ( .A(n64333), .Z(n64327) );
  IV U80340 ( .A(n59995), .Z(n64330) );
  IV U80341 ( .A(n59996), .Z(n59997) );
  NOR U80342 ( .A(n64330), .B(n59997), .Z(n65268) );
  IV U80343 ( .A(n59998), .Z(n59999) );
  NOR U80344 ( .A(n60000), .B(n59999), .Z(n69502) );
  IV U80345 ( .A(n60001), .Z(n60002) );
  NOR U80346 ( .A(n60002), .B(n64308), .Z(n60003) );
  IV U80347 ( .A(n60003), .Z(n69500) );
  IV U80348 ( .A(n60004), .Z(n60005) );
  NOR U80349 ( .A(n60008), .B(n60005), .Z(n65282) );
  IV U80350 ( .A(n60006), .Z(n60007) );
  NOR U80351 ( .A(n60008), .B(n60007), .Z(n65279) );
  IV U80352 ( .A(n60009), .Z(n60013) );
  IV U80353 ( .A(n60010), .Z(n60011) );
  NOR U80354 ( .A(n60013), .B(n60011), .Z(n65312) );
  IV U80355 ( .A(n60012), .Z(n60014) );
  NOR U80356 ( .A(n60014), .B(n60013), .Z(n65309) );
  IV U80357 ( .A(n60015), .Z(n60016) );
  NOR U80358 ( .A(n60016), .B(n60018), .Z(n65318) );
  IV U80359 ( .A(n60017), .Z(n60019) );
  NOR U80360 ( .A(n60019), .B(n60018), .Z(n65315) );
  IV U80361 ( .A(n60020), .Z(n60025) );
  IV U80362 ( .A(n60021), .Z(n60022) );
  NOR U80363 ( .A(n60025), .B(n60022), .Z(n65324) );
  IV U80364 ( .A(n60023), .Z(n60024) );
  NOR U80365 ( .A(n60025), .B(n60024), .Z(n65321) );
  IV U80366 ( .A(n60028), .Z(n60026) );
  NOR U80367 ( .A(n60027), .B(n60026), .Z(n69475) );
  NOR U80368 ( .A(n60029), .B(n60028), .Z(n60032) );
  IV U80369 ( .A(n60030), .Z(n60031) );
  NOR U80370 ( .A(n60032), .B(n60031), .Z(n60033) );
  NOR U80371 ( .A(n69475), .B(n60033), .Z(n65331) );
  NOR U80372 ( .A(n60035), .B(n60034), .Z(n69473) );
  IV U80373 ( .A(n60036), .Z(n60043) );
  NOR U80374 ( .A(n60038), .B(n60037), .Z(n60039) );
  IV U80375 ( .A(n60039), .Z(n60040) );
  NOR U80376 ( .A(n60041), .B(n60040), .Z(n60042) );
  IV U80377 ( .A(n60042), .Z(n60045) );
  NOR U80378 ( .A(n60043), .B(n60045), .Z(n65335) );
  IV U80379 ( .A(n60044), .Z(n60046) );
  NOR U80380 ( .A(n60046), .B(n60045), .Z(n64267) );
  IV U80381 ( .A(n60047), .Z(n60048) );
  NOR U80382 ( .A(n60054), .B(n60048), .Z(n60049) );
  IV U80383 ( .A(n60049), .Z(n69469) );
  IV U80384 ( .A(n60050), .Z(n60052) );
  NOR U80385 ( .A(n60052), .B(n60051), .Z(n65338) );
  IV U80386 ( .A(n60053), .Z(n60055) );
  NOR U80387 ( .A(n60055), .B(n60054), .Z(n69465) );
  NOR U80388 ( .A(n65338), .B(n69465), .Z(n64264) );
  IV U80389 ( .A(n60056), .Z(n60058) );
  NOR U80390 ( .A(n60058), .B(n60057), .Z(n65344) );
  IV U80391 ( .A(n60059), .Z(n60065) );
  IV U80392 ( .A(n60060), .Z(n60061) );
  NOR U80393 ( .A(n60065), .B(n60061), .Z(n65349) );
  IV U80394 ( .A(n60062), .Z(n60063) );
  NOR U80395 ( .A(n60065), .B(n60063), .Z(n69451) );
  NOR U80396 ( .A(n60065), .B(n60064), .Z(n69445) );
  IV U80397 ( .A(n60066), .Z(n60068) );
  NOR U80398 ( .A(n60068), .B(n60067), .Z(n69448) );
  NOR U80399 ( .A(n69445), .B(n69448), .Z(n64254) );
  IV U80400 ( .A(n60069), .Z(n60071) );
  NOR U80401 ( .A(n60071), .B(n60070), .Z(n69442) );
  IV U80402 ( .A(n60072), .Z(n60073) );
  NOR U80403 ( .A(n60073), .B(n60075), .Z(n65361) );
  IV U80404 ( .A(n60074), .Z(n60076) );
  NOR U80405 ( .A(n60076), .B(n60075), .Z(n65359) );
  NOR U80406 ( .A(n65361), .B(n65359), .Z(n60077) );
  IV U80407 ( .A(n60077), .Z(n69437) );
  NOR U80408 ( .A(n60079), .B(n60078), .Z(n60080) );
  IV U80409 ( .A(n60080), .Z(n65371) );
  NOR U80410 ( .A(n60081), .B(n65371), .Z(n60085) );
  IV U80411 ( .A(n60082), .Z(n60084) );
  IV U80412 ( .A(n60083), .Z(n64244) );
  NOR U80413 ( .A(n60084), .B(n64244), .Z(n69430) );
  NOR U80414 ( .A(n60085), .B(n69430), .Z(n64250) );
  IV U80415 ( .A(n60086), .Z(n65385) );
  IV U80416 ( .A(n60087), .Z(n60088) );
  NOR U80417 ( .A(n65385), .B(n60088), .Z(n65377) );
  IV U80418 ( .A(n60089), .Z(n60090) );
  NOR U80419 ( .A(n60090), .B(n60093), .Z(n65389) );
  IV U80420 ( .A(n60091), .Z(n65400) );
  NOR U80421 ( .A(n65395), .B(n65400), .Z(n60095) );
  IV U80422 ( .A(n60092), .Z(n60094) );
  NOR U80423 ( .A(n60094), .B(n60093), .Z(n65392) );
  NOR U80424 ( .A(n60095), .B(n65392), .Z(n64236) );
  IV U80425 ( .A(n65396), .Z(n60096) );
  NOR U80426 ( .A(n65395), .B(n60096), .Z(n65401) );
  IV U80427 ( .A(n60097), .Z(n60102) );
  IV U80428 ( .A(n60098), .Z(n60099) );
  NOR U80429 ( .A(n60102), .B(n60099), .Z(n65404) );
  IV U80430 ( .A(n60100), .Z(n60101) );
  NOR U80431 ( .A(n60102), .B(n60101), .Z(n65410) );
  IV U80432 ( .A(n60103), .Z(n60104) );
  NOR U80433 ( .A(n60104), .B(n60109), .Z(n65412) );
  NOR U80434 ( .A(n65410), .B(n65412), .Z(n64235) );
  IV U80435 ( .A(n60105), .Z(n60107) );
  NOR U80436 ( .A(n60107), .B(n60106), .Z(n69409) );
  IV U80437 ( .A(n60108), .Z(n60110) );
  NOR U80438 ( .A(n60110), .B(n60109), .Z(n65415) );
  NOR U80439 ( .A(n69409), .B(n65415), .Z(n64234) );
  IV U80440 ( .A(n60111), .Z(n60113) );
  NOR U80441 ( .A(n60113), .B(n60112), .Z(n69401) );
  IV U80442 ( .A(n60114), .Z(n60116) );
  NOR U80443 ( .A(n60116), .B(n60115), .Z(n69406) );
  NOR U80444 ( .A(n69401), .B(n69406), .Z(n64233) );
  IV U80445 ( .A(n60117), .Z(n60118) );
  NOR U80446 ( .A(n60119), .B(n60118), .Z(n69398) );
  NOR U80447 ( .A(n69398), .B(n69402), .Z(n64232) );
  IV U80448 ( .A(n60120), .Z(n60124) );
  IV U80449 ( .A(n60121), .Z(n65421) );
  NOR U80450 ( .A(n60122), .B(n65421), .Z(n60123) );
  IV U80451 ( .A(n60123), .Z(n64229) );
  NOR U80452 ( .A(n60124), .B(n64229), .Z(n69395) );
  IV U80453 ( .A(n60125), .Z(n60126) );
  NOR U80454 ( .A(n60126), .B(n60132), .Z(n60127) );
  IV U80455 ( .A(n60127), .Z(n65425) );
  IV U80456 ( .A(n60128), .Z(n60130) );
  NOR U80457 ( .A(n60130), .B(n60129), .Z(n69385) );
  IV U80458 ( .A(n60131), .Z(n60133) );
  NOR U80459 ( .A(n60133), .B(n60132), .Z(n69390) );
  NOR U80460 ( .A(n69385), .B(n69390), .Z(n64223) );
  IV U80461 ( .A(n60134), .Z(n60136) );
  NOR U80462 ( .A(n60136), .B(n60135), .Z(n69384) );
  IV U80463 ( .A(n69384), .Z(n69381) );
  IV U80464 ( .A(n60137), .Z(n64220) );
  IV U80465 ( .A(n60138), .Z(n60139) );
  NOR U80466 ( .A(n60139), .B(n60152), .Z(n60144) );
  IV U80467 ( .A(n60144), .Z(n60140) );
  NOR U80468 ( .A(n64220), .B(n60140), .Z(n60141) );
  IV U80469 ( .A(n60141), .Z(n60142) );
  NOR U80470 ( .A(n60146), .B(n60142), .Z(n65434) );
  IV U80471 ( .A(n60143), .Z(n60149) );
  XOR U80472 ( .A(n64220), .B(n60144), .Z(n60145) );
  NOR U80473 ( .A(n60146), .B(n60145), .Z(n60147) );
  IV U80474 ( .A(n60147), .Z(n60148) );
  NOR U80475 ( .A(n60149), .B(n60148), .Z(n60150) );
  IV U80476 ( .A(n60150), .Z(n60151) );
  NOR U80477 ( .A(n60152), .B(n60151), .Z(n65432) );
  NOR U80478 ( .A(n65434), .B(n65432), .Z(n64214) );
  IV U80479 ( .A(n60153), .Z(n60154) );
  NOR U80480 ( .A(n64209), .B(n60154), .Z(n65438) );
  IV U80481 ( .A(n60155), .Z(n60156) );
  NOR U80482 ( .A(n60156), .B(n64198), .Z(n60157) );
  IV U80483 ( .A(n60157), .Z(n65453) );
  IV U80484 ( .A(n60158), .Z(n64199) );
  IV U80485 ( .A(n60159), .Z(n60161) );
  NOR U80486 ( .A(n60161), .B(n60160), .Z(n65462) );
  IV U80487 ( .A(n60162), .Z(n60163) );
  NOR U80488 ( .A(n60163), .B(n64192), .Z(n65460) );
  NOR U80489 ( .A(n65462), .B(n65460), .Z(n64187) );
  IV U80490 ( .A(n60164), .Z(n60168) );
  NOR U80491 ( .A(n60166), .B(n60165), .Z(n60167) );
  IV U80492 ( .A(n60167), .Z(n60170) );
  NOR U80493 ( .A(n60168), .B(n60170), .Z(n69368) );
  IV U80494 ( .A(n60169), .Z(n60171) );
  NOR U80495 ( .A(n60171), .B(n60170), .Z(n69365) );
  IV U80496 ( .A(n60172), .Z(n60173) );
  NOR U80497 ( .A(n60174), .B(n60173), .Z(n65467) );
  IV U80498 ( .A(n60175), .Z(n60176) );
  NOR U80499 ( .A(n60182), .B(n60176), .Z(n65472) );
  NOR U80500 ( .A(n65467), .B(n65472), .Z(n60177) );
  IV U80501 ( .A(n60177), .Z(n64179) );
  IV U80502 ( .A(n60178), .Z(n60180) );
  NOR U80503 ( .A(n60180), .B(n60179), .Z(n75889) );
  IV U80504 ( .A(n60181), .Z(n60183) );
  NOR U80505 ( .A(n60183), .B(n60182), .Z(n75881) );
  NOR U80506 ( .A(n75889), .B(n75881), .Z(n65471) );
  IV U80507 ( .A(n60184), .Z(n60186) );
  NOR U80508 ( .A(n60186), .B(n60185), .Z(n69357) );
  IV U80509 ( .A(n60187), .Z(n60189) );
  NOR U80510 ( .A(n60189), .B(n60188), .Z(n69361) );
  NOR U80511 ( .A(n69357), .B(n69361), .Z(n64178) );
  IV U80512 ( .A(n75895), .Z(n60190) );
  NOR U80513 ( .A(n60190), .B(n75894), .Z(n64148) );
  IV U80514 ( .A(n64148), .Z(n64141) );
  NOR U80515 ( .A(n60191), .B(n65492), .Z(n64145) );
  IV U80516 ( .A(n60192), .Z(n60193) );
  NOR U80517 ( .A(n60194), .B(n60193), .Z(n65497) );
  IV U80518 ( .A(n60195), .Z(n64135) );
  IV U80519 ( .A(n60196), .Z(n60197) );
  NOR U80520 ( .A(n64135), .B(n60197), .Z(n65502) );
  NOR U80521 ( .A(n65497), .B(n65502), .Z(n64139) );
  IV U80522 ( .A(n60198), .Z(n60199) );
  NOR U80523 ( .A(n60200), .B(n60199), .Z(n65518) );
  IV U80524 ( .A(n60201), .Z(n60203) );
  NOR U80525 ( .A(n60203), .B(n60202), .Z(n60204) );
  IV U80526 ( .A(n60204), .Z(n65517) );
  IV U80527 ( .A(n60205), .Z(n60206) );
  NOR U80528 ( .A(n60206), .B(n60212), .Z(n60207) );
  IV U80529 ( .A(n60207), .Z(n65522) );
  IV U80530 ( .A(n60208), .Z(n60209) );
  NOR U80531 ( .A(n60210), .B(n60209), .Z(n65532) );
  IV U80532 ( .A(n60211), .Z(n60213) );
  NOR U80533 ( .A(n60213), .B(n60212), .Z(n65526) );
  NOR U80534 ( .A(n65532), .B(n65526), .Z(n64127) );
  IV U80535 ( .A(n60214), .Z(n60215) );
  NOR U80536 ( .A(n60215), .B(n60218), .Z(n65529) );
  IV U80537 ( .A(n60216), .Z(n60217) );
  NOR U80538 ( .A(n60218), .B(n60217), .Z(n60219) );
  IV U80539 ( .A(n60219), .Z(n65537) );
  IV U80540 ( .A(n60220), .Z(n60221) );
  NOR U80541 ( .A(n60221), .B(n60224), .Z(n69339) );
  IV U80542 ( .A(n60222), .Z(n60223) );
  NOR U80543 ( .A(n60224), .B(n60223), .Z(n69336) );
  IV U80544 ( .A(n60225), .Z(n60226) );
  NOR U80545 ( .A(n60227), .B(n60226), .Z(n65540) );
  IV U80546 ( .A(n60228), .Z(n60233) );
  IV U80547 ( .A(n60229), .Z(n60230) );
  NOR U80548 ( .A(n60233), .B(n60230), .Z(n65545) );
  NOR U80549 ( .A(n65540), .B(n65545), .Z(n64119) );
  IV U80550 ( .A(n60231), .Z(n60232) );
  NOR U80551 ( .A(n60233), .B(n60232), .Z(n65542) );
  IV U80552 ( .A(n60234), .Z(n60235) );
  NOR U80553 ( .A(n60235), .B(n64113), .Z(n65548) );
  IV U80554 ( .A(n60236), .Z(n60237) );
  NOR U80555 ( .A(n60237), .B(n64078), .Z(n65559) );
  IV U80556 ( .A(n60238), .Z(n60239) );
  NOR U80557 ( .A(n60240), .B(n60239), .Z(n60241) );
  IV U80558 ( .A(n60241), .Z(n69318) );
  IV U80559 ( .A(n60242), .Z(n60244) );
  IV U80560 ( .A(n60243), .Z(n60249) );
  NOR U80561 ( .A(n60244), .B(n60249), .Z(n60245) );
  IV U80562 ( .A(n60245), .Z(n65565) );
  NOR U80563 ( .A(n60247), .B(n60246), .Z(n69302) );
  IV U80564 ( .A(n60248), .Z(n60250) );
  NOR U80565 ( .A(n60250), .B(n60249), .Z(n65567) );
  NOR U80566 ( .A(n69302), .B(n65567), .Z(n64059) );
  IV U80567 ( .A(n60251), .Z(n60258) );
  NOR U80568 ( .A(n60253), .B(n60252), .Z(n60254) );
  IV U80569 ( .A(n60254), .Z(n60255) );
  NOR U80570 ( .A(n60256), .B(n60255), .Z(n60257) );
  IV U80571 ( .A(n60257), .Z(n60260) );
  NOR U80572 ( .A(n60258), .B(n60260), .Z(n65572) );
  IV U80573 ( .A(n60259), .Z(n60261) );
  NOR U80574 ( .A(n60261), .B(n60260), .Z(n65569) );
  IV U80575 ( .A(n60262), .Z(n60264) );
  NOR U80576 ( .A(n60264), .B(n60263), .Z(n65575) );
  IV U80577 ( .A(n60265), .Z(n60267) );
  NOR U80578 ( .A(n60267), .B(n60266), .Z(n65586) );
  IV U80579 ( .A(n60268), .Z(n60269) );
  NOR U80580 ( .A(n60269), .B(n60271), .Z(n65583) );
  IV U80581 ( .A(n60270), .Z(n60272) );
  NOR U80582 ( .A(n60272), .B(n60271), .Z(n65589) );
  IV U80583 ( .A(n60273), .Z(n60275) );
  NOR U80584 ( .A(n60275), .B(n60274), .Z(n65596) );
  IV U80585 ( .A(n60276), .Z(n60278) );
  NOR U80586 ( .A(n60278), .B(n60277), .Z(n65592) );
  NOR U80587 ( .A(n65596), .B(n65592), .Z(n64052) );
  IV U80588 ( .A(n60279), .Z(n60281) );
  IV U80589 ( .A(n60280), .Z(n64046) );
  NOR U80590 ( .A(n60281), .B(n64046), .Z(n65599) );
  IV U80591 ( .A(n60282), .Z(n60283) );
  NOR U80592 ( .A(n60286), .B(n60283), .Z(n69279) );
  IV U80593 ( .A(n69279), .Z(n79826) );
  IV U80594 ( .A(n60284), .Z(n60285) );
  NOR U80595 ( .A(n60286), .B(n60285), .Z(n75998) );
  IV U80596 ( .A(n60287), .Z(n60289) );
  IV U80597 ( .A(n60288), .Z(n65605) );
  NOR U80598 ( .A(n60289), .B(n65605), .Z(n69283) );
  NOR U80599 ( .A(n75998), .B(n69283), .Z(n64044) );
  IV U80600 ( .A(n60290), .Z(n60291) );
  NOR U80601 ( .A(n60292), .B(n60291), .Z(n65617) );
  NOR U80602 ( .A(n60294), .B(n60293), .Z(n65612) );
  NOR U80603 ( .A(n65617), .B(n65612), .Z(n60295) );
  IV U80604 ( .A(n60295), .Z(n64039) );
  NOR U80605 ( .A(n60297), .B(n60296), .Z(n65614) );
  IV U80606 ( .A(n60298), .Z(n60299) );
  NOR U80607 ( .A(n60300), .B(n60299), .Z(n65642) );
  NOR U80608 ( .A(n65642), .B(n69253), .Z(n64011) );
  IV U80609 ( .A(n60301), .Z(n60303) );
  IV U80610 ( .A(n60302), .Z(n64001) );
  NOR U80611 ( .A(n60303), .B(n64001), .Z(n69248) );
  NOR U80612 ( .A(n65646), .B(n69248), .Z(n63999) );
  IV U80613 ( .A(n60304), .Z(n60305) );
  NOR U80614 ( .A(n60306), .B(n60305), .Z(n65658) );
  NOR U80615 ( .A(n60307), .B(n65649), .Z(n60308) );
  NOR U80616 ( .A(n65658), .B(n60308), .Z(n63998) );
  IV U80617 ( .A(n60309), .Z(n60312) );
  IV U80618 ( .A(n60310), .Z(n60311) );
  NOR U80619 ( .A(n60312), .B(n60311), .Z(n65655) );
  IV U80620 ( .A(n60313), .Z(n60315) );
  XOR U80621 ( .A(n60317), .B(n60320), .Z(n60314) );
  NOR U80622 ( .A(n60315), .B(n60314), .Z(n60316) );
  IV U80623 ( .A(n60316), .Z(n65662) );
  IV U80624 ( .A(n60317), .Z(n60318) );
  NOR U80625 ( .A(n60318), .B(n60320), .Z(n69240) );
  IV U80626 ( .A(n60319), .Z(n60321) );
  NOR U80627 ( .A(n60321), .B(n60320), .Z(n69243) );
  NOR U80628 ( .A(n69240), .B(n69243), .Z(n63997) );
  IV U80629 ( .A(n60322), .Z(n60323) );
  NOR U80630 ( .A(n60324), .B(n60323), .Z(n65667) );
  IV U80631 ( .A(n60325), .Z(n60327) );
  NOR U80632 ( .A(n60327), .B(n60326), .Z(n69237) );
  NOR U80633 ( .A(n65667), .B(n69237), .Z(n63996) );
  IV U80634 ( .A(n60328), .Z(n60330) );
  NOR U80635 ( .A(n60330), .B(n60329), .Z(n60331) );
  IV U80636 ( .A(n60331), .Z(n63991) );
  IV U80637 ( .A(n60332), .Z(n60338) );
  NOR U80638 ( .A(n60333), .B(n60340), .Z(n60334) );
  IV U80639 ( .A(n60334), .Z(n60335) );
  NOR U80640 ( .A(n60336), .B(n60335), .Z(n60337) );
  IV U80641 ( .A(n60337), .Z(n63978) );
  NOR U80642 ( .A(n60338), .B(n63978), .Z(n65674) );
  IV U80643 ( .A(n60339), .Z(n60341) );
  NOR U80644 ( .A(n60341), .B(n60340), .Z(n65679) );
  NOR U80645 ( .A(n65674), .B(n65679), .Z(n63973) );
  IV U80646 ( .A(n60342), .Z(n60343) );
  NOR U80647 ( .A(n60344), .B(n60343), .Z(n69221) );
  IV U80648 ( .A(n60345), .Z(n60346) );
  NOR U80649 ( .A(n60347), .B(n60346), .Z(n69215) );
  IV U80650 ( .A(n60348), .Z(n60349) );
  NOR U80651 ( .A(n60349), .B(n63965), .Z(n65688) );
  NOR U80652 ( .A(n69215), .B(n65688), .Z(n63961) );
  IV U80653 ( .A(n60350), .Z(n63945) );
  NOR U80654 ( .A(n60351), .B(n63945), .Z(n63942) );
  IV U80655 ( .A(n60352), .Z(n60355) );
  IV U80656 ( .A(n60353), .Z(n60354) );
  NOR U80657 ( .A(n60355), .B(n60354), .Z(n60356) );
  IV U80658 ( .A(n60356), .Z(n69201) );
  XOR U80659 ( .A(n63926), .B(n63928), .Z(n60359) );
  IV U80660 ( .A(n60357), .Z(n60358) );
  NOR U80661 ( .A(n60359), .B(n60358), .Z(n65691) );
  IV U80662 ( .A(n60360), .Z(n60361) );
  NOR U80663 ( .A(n60361), .B(n63928), .Z(n69203) );
  IV U80664 ( .A(n60362), .Z(n60365) );
  IV U80665 ( .A(n60363), .Z(n60364) );
  NOR U80666 ( .A(n60365), .B(n60364), .Z(n65705) );
  IV U80667 ( .A(n60366), .Z(n60368) );
  NOR U80668 ( .A(n60368), .B(n60367), .Z(n65701) );
  NOR U80669 ( .A(n65705), .B(n65701), .Z(n63922) );
  IV U80670 ( .A(n60369), .Z(n60372) );
  NOR U80671 ( .A(n60370), .B(n63917), .Z(n60371) );
  IV U80672 ( .A(n60371), .Z(n60376) );
  NOR U80673 ( .A(n60372), .B(n60376), .Z(n65716) );
  NOR U80674 ( .A(n65711), .B(n65716), .Z(n63920) );
  IV U80675 ( .A(n60373), .Z(n60374) );
  NOR U80676 ( .A(n60374), .B(n60376), .Z(n65713) );
  IV U80677 ( .A(n60375), .Z(n60377) );
  NOR U80678 ( .A(n60377), .B(n60376), .Z(n65719) );
  IV U80679 ( .A(n60378), .Z(n60379) );
  NOR U80680 ( .A(n60380), .B(n60379), .Z(n69192) );
  IV U80681 ( .A(n60381), .Z(n60382) );
  NOR U80682 ( .A(n60382), .B(n60384), .Z(n65722) );
  IV U80683 ( .A(n60383), .Z(n60385) );
  NOR U80684 ( .A(n60385), .B(n60384), .Z(n63907) );
  IV U80685 ( .A(n60386), .Z(n60388) );
  IV U80686 ( .A(n60387), .Z(n63897) );
  NOR U80687 ( .A(n60388), .B(n63897), .Z(n60389) );
  IV U80688 ( .A(n60389), .Z(n69178) );
  IV U80689 ( .A(n60390), .Z(n60391) );
  NOR U80690 ( .A(n60392), .B(n60391), .Z(n65747) );
  IV U80691 ( .A(n60393), .Z(n60398) );
  IV U80692 ( .A(n60394), .Z(n60395) );
  NOR U80693 ( .A(n60398), .B(n60395), .Z(n65744) );
  IV U80694 ( .A(n60396), .Z(n60397) );
  NOR U80695 ( .A(n60398), .B(n60397), .Z(n65749) );
  IV U80696 ( .A(n60399), .Z(n60400) );
  NOR U80697 ( .A(n60400), .B(n60402), .Z(n69161) );
  IV U80698 ( .A(n60401), .Z(n60403) );
  NOR U80699 ( .A(n60403), .B(n60402), .Z(n69158) );
  IV U80700 ( .A(n60404), .Z(n60405) );
  NOR U80701 ( .A(n60405), .B(n60407), .Z(n65755) );
  IV U80702 ( .A(n60406), .Z(n60408) );
  NOR U80703 ( .A(n60408), .B(n60407), .Z(n60409) );
  IV U80704 ( .A(n60409), .Z(n65754) );
  IV U80705 ( .A(n60410), .Z(n60412) );
  NOR U80706 ( .A(n60412), .B(n60411), .Z(n69154) );
  IV U80707 ( .A(n60413), .Z(n60415) );
  NOR U80708 ( .A(n60415), .B(n60414), .Z(n65758) );
  NOR U80709 ( .A(n69154), .B(n65758), .Z(n63874) );
  NOR U80710 ( .A(n60416), .B(n74230), .Z(n65764) );
  IV U80711 ( .A(n60417), .Z(n60418) );
  NOR U80712 ( .A(n60419), .B(n60418), .Z(n65773) );
  IV U80713 ( .A(n60420), .Z(n60422) );
  NOR U80714 ( .A(n60422), .B(n60421), .Z(n65769) );
  NOR U80715 ( .A(n65773), .B(n65769), .Z(n63863) );
  IV U80716 ( .A(n60423), .Z(n60425) );
  NOR U80717 ( .A(n60425), .B(n60424), .Z(n65780) );
  IV U80718 ( .A(n60426), .Z(n60428) );
  NOR U80719 ( .A(n60428), .B(n60427), .Z(n65783) );
  IV U80720 ( .A(n60429), .Z(n60430) );
  NOR U80721 ( .A(n60431), .B(n60430), .Z(n65792) );
  IV U80722 ( .A(n60432), .Z(n60433) );
  NOR U80723 ( .A(n60434), .B(n60433), .Z(n65789) );
  NOR U80724 ( .A(n65792), .B(n65789), .Z(n63844) );
  IV U80725 ( .A(n60435), .Z(n60437) );
  NOR U80726 ( .A(n60437), .B(n60436), .Z(n69126) );
  NOR U80727 ( .A(n60439), .B(n60438), .Z(n70743) );
  IV U80728 ( .A(n60440), .Z(n60442) );
  IV U80729 ( .A(n60441), .Z(n63836) );
  NOR U80730 ( .A(n60442), .B(n63836), .Z(n74158) );
  NOR U80731 ( .A(n70743), .B(n74158), .Z(n69118) );
  IV U80732 ( .A(n60443), .Z(n60446) );
  NOR U80733 ( .A(n60452), .B(n60444), .Z(n60445) );
  IV U80734 ( .A(n60445), .Z(n60448) );
  NOR U80735 ( .A(n60446), .B(n60448), .Z(n69111) );
  IV U80736 ( .A(n60447), .Z(n60449) );
  NOR U80737 ( .A(n60449), .B(n60448), .Z(n69108) );
  IV U80738 ( .A(n60450), .Z(n60451) );
  NOR U80739 ( .A(n60452), .B(n60451), .Z(n65802) );
  IV U80740 ( .A(n60453), .Z(n60454) );
  NOR U80741 ( .A(n60459), .B(n60454), .Z(n65799) );
  IV U80742 ( .A(n60455), .Z(n60457) );
  NOR U80743 ( .A(n60457), .B(n60456), .Z(n70757) );
  IV U80744 ( .A(n60458), .Z(n60460) );
  NOR U80745 ( .A(n60460), .B(n60459), .Z(n70752) );
  NOR U80746 ( .A(n70757), .B(n70752), .Z(n69104) );
  IV U80747 ( .A(n69104), .Z(n63834) );
  IV U80748 ( .A(n60461), .Z(n63833) );
  IV U80749 ( .A(n60462), .Z(n60463) );
  NOR U80750 ( .A(n63833), .B(n60463), .Z(n65807) );
  IV U80751 ( .A(n60464), .Z(n60465) );
  NOR U80752 ( .A(n60465), .B(n63827), .Z(n65817) );
  IV U80753 ( .A(n60466), .Z(n60467) );
  NOR U80754 ( .A(n60467), .B(n63827), .Z(n65811) );
  NOR U80755 ( .A(n65817), .B(n65811), .Z(n63824) );
  IV U80756 ( .A(n60468), .Z(n63820) );
  IV U80757 ( .A(n60469), .Z(n60470) );
  NOR U80758 ( .A(n63820), .B(n60470), .Z(n65821) );
  IV U80759 ( .A(n60471), .Z(n60472) );
  NOR U80760 ( .A(n63815), .B(n60472), .Z(n69096) );
  NOR U80761 ( .A(n65821), .B(n69096), .Z(n63817) );
  IV U80762 ( .A(n60473), .Z(n60475) );
  IV U80763 ( .A(n60474), .Z(n63808) );
  NOR U80764 ( .A(n60475), .B(n63808), .Z(n69081) );
  NOR U80765 ( .A(n60476), .B(n65826), .Z(n60480) );
  IV U80766 ( .A(n60477), .Z(n60479) );
  IV U80767 ( .A(n60478), .Z(n63796) );
  NOR U80768 ( .A(n60479), .B(n63796), .Z(n65829) );
  NOR U80769 ( .A(n60480), .B(n65829), .Z(n63806) );
  IV U80770 ( .A(n60481), .Z(n60483) );
  NOR U80771 ( .A(n60483), .B(n60482), .Z(n69071) );
  IV U80772 ( .A(n65836), .Z(n60485) );
  NOR U80773 ( .A(n60485), .B(n60484), .Z(n70808) );
  IV U80774 ( .A(n60486), .Z(n60488) );
  NOR U80775 ( .A(n60488), .B(n60487), .Z(n69068) );
  NOR U80776 ( .A(n70808), .B(n69068), .Z(n63793) );
  NOR U80777 ( .A(n60489), .B(n65837), .Z(n63792) );
  IV U80778 ( .A(n60490), .Z(n60491) );
  NOR U80779 ( .A(n60492), .B(n60491), .Z(n65842) );
  IV U80780 ( .A(n60493), .Z(n60499) );
  IV U80781 ( .A(n60494), .Z(n60495) );
  NOR U80782 ( .A(n60499), .B(n60495), .Z(n65849) );
  NOR U80783 ( .A(n65842), .B(n65849), .Z(n60496) );
  IV U80784 ( .A(n60496), .Z(n63791) );
  IV U80785 ( .A(n60497), .Z(n60498) );
  NOR U80786 ( .A(n60499), .B(n60498), .Z(n65846) );
  IV U80787 ( .A(n60500), .Z(n60501) );
  NOR U80788 ( .A(n60501), .B(n60504), .Z(n65855) );
  IV U80789 ( .A(n60502), .Z(n60503) );
  NOR U80790 ( .A(n60504), .B(n60503), .Z(n65852) );
  IV U80791 ( .A(n60505), .Z(n60506) );
  NOR U80792 ( .A(n60509), .B(n60506), .Z(n69063) );
  IV U80793 ( .A(n69063), .Z(n74103) );
  IV U80794 ( .A(n60507), .Z(n60508) );
  NOR U80795 ( .A(n60509), .B(n60508), .Z(n76271) );
  IV U80796 ( .A(n60510), .Z(n60512) );
  IV U80797 ( .A(n60511), .Z(n60516) );
  NOR U80798 ( .A(n60512), .B(n60516), .Z(n65858) );
  NOR U80799 ( .A(n76271), .B(n65858), .Z(n70832) );
  IV U80800 ( .A(n60513), .Z(n60514) );
  NOR U80801 ( .A(n65860), .B(n60514), .Z(n69058) );
  IV U80802 ( .A(n60515), .Z(n65866) );
  NOR U80803 ( .A(n65866), .B(n60516), .Z(n60517) );
  NOR U80804 ( .A(n69058), .B(n60517), .Z(n63790) );
  IV U80805 ( .A(n65861), .Z(n60518) );
  NOR U80806 ( .A(n65860), .B(n60518), .Z(n69055) );
  IV U80807 ( .A(n60519), .Z(n60521) );
  NOR U80808 ( .A(n60521), .B(n60520), .Z(n60522) );
  NOR U80809 ( .A(n60522), .B(n65879), .Z(n63785) );
  IV U80810 ( .A(n60523), .Z(n60524) );
  NOR U80811 ( .A(n60524), .B(n60530), .Z(n70853) );
  IV U80812 ( .A(n60525), .Z(n60527) );
  NOR U80813 ( .A(n60527), .B(n60526), .Z(n70847) );
  NOR U80814 ( .A(n70853), .B(n70847), .Z(n65885) );
  IV U80815 ( .A(n65885), .Z(n63784) );
  IV U80816 ( .A(n60528), .Z(n60529) );
  NOR U80817 ( .A(n60530), .B(n60529), .Z(n65882) );
  IV U80818 ( .A(n60531), .Z(n60533) );
  NOR U80819 ( .A(n60533), .B(n60532), .Z(n65890) );
  IV U80820 ( .A(n60534), .Z(n60536) );
  NOR U80821 ( .A(n60536), .B(n60535), .Z(n65887) );
  NOR U80822 ( .A(n65890), .B(n65887), .Z(n63783) );
  IV U80823 ( .A(n60537), .Z(n60538) );
  NOR U80824 ( .A(n60538), .B(n60547), .Z(n65897) );
  IV U80825 ( .A(n60539), .Z(n60541) );
  NOR U80826 ( .A(n60541), .B(n60540), .Z(n69047) );
  NOR U80827 ( .A(n65897), .B(n69047), .Z(n63775) );
  IV U80828 ( .A(n60542), .Z(n60543) );
  NOR U80829 ( .A(n60544), .B(n60543), .Z(n65900) );
  IV U80830 ( .A(n60545), .Z(n60546) );
  NOR U80831 ( .A(n60547), .B(n60546), .Z(n65895) );
  NOR U80832 ( .A(n65900), .B(n65895), .Z(n63774) );
  IV U80833 ( .A(n60548), .Z(n60549) );
  NOR U80834 ( .A(n60550), .B(n60549), .Z(n65903) );
  IV U80835 ( .A(n60551), .Z(n60552) );
  NOR U80836 ( .A(n60552), .B(n63770), .Z(n69042) );
  NOR U80837 ( .A(n65903), .B(n69042), .Z(n63773) );
  IV U80838 ( .A(n60553), .Z(n60554) );
  NOR U80839 ( .A(n60554), .B(n60556), .Z(n69025) );
  IV U80840 ( .A(n60555), .Z(n60557) );
  NOR U80841 ( .A(n60557), .B(n60556), .Z(n69022) );
  IV U80842 ( .A(n60558), .Z(n60560) );
  NOR U80843 ( .A(n60560), .B(n60559), .Z(n60561) );
  IV U80844 ( .A(n60561), .Z(n65948) );
  IV U80845 ( .A(n60562), .Z(n60565) );
  NOR U80846 ( .A(n60563), .B(n60567), .Z(n60564) );
  IV U80847 ( .A(n60564), .Z(n63728) );
  NOR U80848 ( .A(n60565), .B(n63728), .Z(n65944) );
  IV U80849 ( .A(n60566), .Z(n60568) );
  NOR U80850 ( .A(n60568), .B(n60567), .Z(n63723) );
  IV U80851 ( .A(n60569), .Z(n79420) );
  IV U80852 ( .A(n79421), .Z(n60570) );
  NOR U80853 ( .A(n79420), .B(n60570), .Z(n65959) );
  NOR U80854 ( .A(n60572), .B(n60571), .Z(n65964) );
  XOR U80855 ( .A(n65966), .B(n65964), .Z(n60573) );
  NOR U80856 ( .A(n65959), .B(n60573), .Z(n63709) );
  NOR U80857 ( .A(n60574), .B(n65971), .Z(n63708) );
  IV U80858 ( .A(n60575), .Z(n60576) );
  NOR U80859 ( .A(n60577), .B(n60576), .Z(n65980) );
  IV U80860 ( .A(n60578), .Z(n60581) );
  IV U80861 ( .A(n60579), .Z(n60580) );
  NOR U80862 ( .A(n60581), .B(n60580), .Z(n65982) );
  NOR U80863 ( .A(n65980), .B(n65982), .Z(n63700) );
  IV U80864 ( .A(n60582), .Z(n60583) );
  NOR U80865 ( .A(n60583), .B(n60589), .Z(n65996) );
  IV U80866 ( .A(n60584), .Z(n60586) );
  NOR U80867 ( .A(n60586), .B(n60585), .Z(n70965) );
  IV U80868 ( .A(n60587), .Z(n60588) );
  NOR U80869 ( .A(n60589), .B(n60588), .Z(n70960) );
  NOR U80870 ( .A(n70965), .B(n70960), .Z(n69001) );
  IV U80871 ( .A(n60590), .Z(n60592) );
  NOR U80872 ( .A(n60592), .B(n60591), .Z(n68985) );
  IV U80873 ( .A(n60593), .Z(n60595) );
  NOR U80874 ( .A(n60595), .B(n60594), .Z(n68987) );
  NOR U80875 ( .A(n68985), .B(n68987), .Z(n63684) );
  IV U80876 ( .A(n60596), .Z(n60597) );
  NOR U80877 ( .A(n63680), .B(n60597), .Z(n66001) );
  IV U80878 ( .A(n60598), .Z(n60600) );
  NOR U80879 ( .A(n60600), .B(n60599), .Z(n68976) );
  IV U80880 ( .A(n60601), .Z(n68975) );
  IV U80881 ( .A(n60602), .Z(n60603) );
  NOR U80882 ( .A(n60604), .B(n60603), .Z(n66008) );
  IV U80883 ( .A(n60605), .Z(n60607) );
  NOR U80884 ( .A(n60607), .B(n60606), .Z(n68971) );
  NOR U80885 ( .A(n66008), .B(n68971), .Z(n63675) );
  IV U80886 ( .A(n60608), .Z(n63674) );
  IV U80887 ( .A(n60609), .Z(n60610) );
  NOR U80888 ( .A(n63674), .B(n60610), .Z(n63666) );
  IV U80889 ( .A(n60611), .Z(n60612) );
  NOR U80890 ( .A(n60612), .B(n63657), .Z(n63664) );
  IV U80891 ( .A(n63664), .Z(n63652) );
  NOR U80892 ( .A(n60613), .B(n66019), .Z(n63654) );
  IV U80893 ( .A(n60614), .Z(n60615) );
  NOR U80894 ( .A(n60616), .B(n60615), .Z(n66016) );
  NOR U80895 ( .A(n63654), .B(n66016), .Z(n63651) );
  IV U80896 ( .A(n60617), .Z(n60618) );
  NOR U80897 ( .A(n60619), .B(n60618), .Z(n68951) );
  IV U80898 ( .A(n60620), .Z(n60621) );
  NOR U80899 ( .A(n60622), .B(n60621), .Z(n66026) );
  NOR U80900 ( .A(n68951), .B(n66026), .Z(n63650) );
  IV U80901 ( .A(n60623), .Z(n68947) );
  NOR U80902 ( .A(n60624), .B(n68947), .Z(n68954) );
  IV U80903 ( .A(n60625), .Z(n60626) );
  NOR U80904 ( .A(n60626), .B(n63630), .Z(n60627) );
  IV U80905 ( .A(n60627), .Z(n66036) );
  IV U80906 ( .A(n60628), .Z(n60629) );
  NOR U80907 ( .A(n60630), .B(n60629), .Z(n68940) );
  IV U80908 ( .A(n60631), .Z(n60633) );
  NOR U80909 ( .A(n60633), .B(n60632), .Z(n66038) );
  NOR U80910 ( .A(n68940), .B(n66038), .Z(n63628) );
  IV U80911 ( .A(n60634), .Z(n60635) );
  NOR U80912 ( .A(n60635), .B(n63625), .Z(n63619) );
  IV U80913 ( .A(n63619), .Z(n63608) );
  IV U80914 ( .A(n60636), .Z(n66047) );
  NOR U80915 ( .A(n60637), .B(n66047), .Z(n63609) );
  IV U80916 ( .A(n60638), .Z(n60640) );
  NOR U80917 ( .A(n60640), .B(n60639), .Z(n66043) );
  NOR U80918 ( .A(n63609), .B(n66043), .Z(n63606) );
  NOR U80919 ( .A(n60641), .B(n66054), .Z(n63605) );
  IV U80920 ( .A(n60642), .Z(n60643) );
  NOR U80921 ( .A(n60643), .B(n60648), .Z(n66086) );
  IV U80922 ( .A(n60644), .Z(n60646) );
  NOR U80923 ( .A(n60646), .B(n60645), .Z(n66084) );
  NOR U80924 ( .A(n66086), .B(n66084), .Z(n63592) );
  IV U80925 ( .A(n60647), .Z(n60649) );
  NOR U80926 ( .A(n60649), .B(n60648), .Z(n60650) );
  IV U80927 ( .A(n60650), .Z(n66089) );
  IV U80928 ( .A(n60651), .Z(n60653) );
  NOR U80929 ( .A(n60653), .B(n60652), .Z(n60654) );
  IV U80930 ( .A(n60654), .Z(n63585) );
  IV U80931 ( .A(n68922), .Z(n63571) );
  IV U80932 ( .A(n60655), .Z(n68921) );
  NOR U80933 ( .A(n63571), .B(n68921), .Z(n66094) );
  IV U80934 ( .A(n60656), .Z(n60658) );
  NOR U80935 ( .A(n60658), .B(n60657), .Z(n66096) );
  NOR U80936 ( .A(n66094), .B(n66096), .Z(n63569) );
  IV U80937 ( .A(n60659), .Z(n60662) );
  NOR U80938 ( .A(n60660), .B(n63566), .Z(n60661) );
  IV U80939 ( .A(n60661), .Z(n60667) );
  NOR U80940 ( .A(n60662), .B(n60667), .Z(n66102) );
  IV U80941 ( .A(n60663), .Z(n60665) );
  NOR U80942 ( .A(n60665), .B(n60664), .Z(n66106) );
  IV U80943 ( .A(n60666), .Z(n60668) );
  NOR U80944 ( .A(n60668), .B(n60667), .Z(n66100) );
  NOR U80945 ( .A(n66106), .B(n66100), .Z(n63568) );
  IV U80946 ( .A(n60669), .Z(n60671) );
  NOR U80947 ( .A(n60671), .B(n60670), .Z(n66114) );
  IV U80948 ( .A(n60672), .Z(n60673) );
  NOR U80949 ( .A(n60673), .B(n60676), .Z(n68912) );
  IV U80950 ( .A(n60674), .Z(n60675) );
  NOR U80951 ( .A(n60676), .B(n60675), .Z(n60677) );
  NOR U80952 ( .A(n68912), .B(n60677), .Z(n73907) );
  IV U80953 ( .A(n60678), .Z(n63545) );
  NOR U80954 ( .A(n60679), .B(n63545), .Z(n63542) );
  IV U80955 ( .A(n60680), .Z(n60681) );
  NOR U80956 ( .A(n60681), .B(n60685), .Z(n60682) );
  IV U80957 ( .A(n60682), .Z(n66123) );
  IV U80958 ( .A(n60683), .Z(n60684) );
  NOR U80959 ( .A(n60685), .B(n60684), .Z(n60686) );
  IV U80960 ( .A(n60686), .Z(n66121) );
  IV U80961 ( .A(n60687), .Z(n60689) );
  NOR U80962 ( .A(n60689), .B(n60688), .Z(n82039) );
  IV U80963 ( .A(n60690), .Z(n60693) );
  IV U80964 ( .A(n60691), .Z(n63532) );
  XOR U80965 ( .A(n63531), .B(n63532), .Z(n60692) );
  NOR U80966 ( .A(n60693), .B(n60692), .Z(n82049) );
  NOR U80967 ( .A(n82039), .B(n82049), .Z(n68906) );
  IV U80968 ( .A(n60694), .Z(n60695) );
  NOR U80969 ( .A(n60695), .B(n63532), .Z(n68903) );
  IV U80970 ( .A(n60696), .Z(n60697) );
  NOR U80971 ( .A(n60698), .B(n60697), .Z(n68908) );
  NOR U80972 ( .A(n68903), .B(n68908), .Z(n63540) );
  IV U80973 ( .A(n60699), .Z(n60701) );
  NOR U80974 ( .A(n60701), .B(n60700), .Z(n68890) );
  IV U80975 ( .A(n60702), .Z(n60707) );
  IV U80976 ( .A(n60703), .Z(n60704) );
  NOR U80977 ( .A(n60704), .B(n63518), .Z(n60705) );
  IV U80978 ( .A(n60705), .Z(n60706) );
  NOR U80979 ( .A(n60707), .B(n60706), .Z(n68883) );
  IV U80980 ( .A(n60708), .Z(n60709) );
  NOR U80981 ( .A(n60710), .B(n60709), .Z(n66141) );
  IV U80982 ( .A(n60711), .Z(n60713) );
  IV U80983 ( .A(n60712), .Z(n60717) );
  NOR U80984 ( .A(n60713), .B(n60717), .Z(n66138) );
  IV U80985 ( .A(n60714), .Z(n60715) );
  NOR U80986 ( .A(n60715), .B(n60723), .Z(n79244) );
  IV U80987 ( .A(n60716), .Z(n60718) );
  NOR U80988 ( .A(n60718), .B(n60717), .Z(n79251) );
  NOR U80989 ( .A(n79244), .B(n79251), .Z(n73859) );
  IV U80990 ( .A(n60719), .Z(n60721) );
  NOR U80991 ( .A(n60721), .B(n60720), .Z(n73864) );
  IV U80992 ( .A(n60722), .Z(n60724) );
  NOR U80993 ( .A(n60724), .B(n60723), .Z(n73851) );
  NOR U80994 ( .A(n73864), .B(n73851), .Z(n66145) );
  IV U80995 ( .A(n60725), .Z(n60727) );
  NOR U80996 ( .A(n60727), .B(n60726), .Z(n68876) );
  NOR U80997 ( .A(n60728), .B(n66150), .Z(n60729) );
  NOR U80998 ( .A(n68876), .B(n60729), .Z(n63515) );
  IV U80999 ( .A(n60730), .Z(n60731) );
  NOR U81000 ( .A(n60732), .B(n60731), .Z(n68874) );
  IV U81001 ( .A(n60733), .Z(n60734) );
  NOR U81002 ( .A(n60735), .B(n60734), .Z(n68865) );
  IV U81003 ( .A(n60736), .Z(n60737) );
  NOR U81004 ( .A(n60738), .B(n60737), .Z(n66157) );
  NOR U81005 ( .A(n68865), .B(n66157), .Z(n63513) );
  IV U81006 ( .A(n60739), .Z(n66165) );
  NOR U81007 ( .A(n66165), .B(n63505), .Z(n60742) );
  IV U81008 ( .A(n60740), .Z(n60741) );
  NOR U81009 ( .A(n63507), .B(n60741), .Z(n66159) );
  NOR U81010 ( .A(n60742), .B(n66159), .Z(n63512) );
  IV U81011 ( .A(n60743), .Z(n63508) );
  IV U81012 ( .A(n60744), .Z(n60745) );
  NOR U81013 ( .A(n60745), .B(n63501), .Z(n66166) );
  IV U81014 ( .A(n60746), .Z(n60747) );
  NOR U81015 ( .A(n60748), .B(n60747), .Z(n68855) );
  IV U81016 ( .A(n60749), .Z(n60750) );
  NOR U81017 ( .A(n60751), .B(n60750), .Z(n68860) );
  NOR U81018 ( .A(n68855), .B(n68860), .Z(n63497) );
  NOR U81019 ( .A(n60753), .B(n60752), .Z(n68847) );
  IV U81020 ( .A(n60754), .Z(n60756) );
  IV U81021 ( .A(n60755), .Z(n63482) );
  NOR U81022 ( .A(n60756), .B(n63482), .Z(n63476) );
  IV U81023 ( .A(n63476), .Z(n63470) );
  IV U81024 ( .A(n60757), .Z(n60759) );
  NOR U81025 ( .A(n60759), .B(n60758), .Z(n68830) );
  IV U81026 ( .A(n60760), .Z(n63464) );
  IV U81027 ( .A(n60761), .Z(n63461) );
  IV U81028 ( .A(n60762), .Z(n60763) );
  NOR U81029 ( .A(n60763), .B(n63461), .Z(n60764) );
  IV U81030 ( .A(n60764), .Z(n66176) );
  IV U81031 ( .A(n60765), .Z(n60766) );
  NOR U81032 ( .A(n60767), .B(n60766), .Z(n68825) );
  NOR U81033 ( .A(n68822), .B(n68825), .Z(n60768) );
  IV U81034 ( .A(n60768), .Z(n60771) );
  IV U81035 ( .A(n60769), .Z(n60770) );
  NOR U81036 ( .A(n60770), .B(n63461), .Z(n66179) );
  NOR U81037 ( .A(n60771), .B(n66179), .Z(n63459) );
  IV U81038 ( .A(n60772), .Z(n60774) );
  NOR U81039 ( .A(n60774), .B(n60773), .Z(n66184) );
  NOR U81040 ( .A(n60776), .B(n60775), .Z(n68819) );
  NOR U81041 ( .A(n66184), .B(n68819), .Z(n63458) );
  NOR U81042 ( .A(n60777), .B(n66204), .Z(n63436) );
  IV U81043 ( .A(n60778), .Z(n60779) );
  NOR U81044 ( .A(n60780), .B(n60779), .Z(n66214) );
  IV U81045 ( .A(n60781), .Z(n60783) );
  IV U81046 ( .A(n60782), .Z(n63431) );
  NOR U81047 ( .A(n60783), .B(n63431), .Z(n68799) );
  NOR U81048 ( .A(n66214), .B(n68799), .Z(n63435) );
  IV U81049 ( .A(n60784), .Z(n60785) );
  NOR U81050 ( .A(n60786), .B(n60785), .Z(n73709) );
  IV U81051 ( .A(n60787), .Z(n60788) );
  NOR U81052 ( .A(n60789), .B(n60788), .Z(n73714) );
  NOR U81053 ( .A(n73709), .B(n73714), .Z(n66246) );
  NOR U81054 ( .A(n60790), .B(n71173), .Z(n66244) );
  IV U81055 ( .A(n60791), .Z(n60793) );
  IV U81056 ( .A(n60792), .Z(n60795) );
  NOR U81057 ( .A(n60793), .B(n60795), .Z(n68743) );
  IV U81058 ( .A(n60794), .Z(n60796) );
  NOR U81059 ( .A(n60796), .B(n60795), .Z(n68744) );
  XOR U81060 ( .A(n68743), .B(n68744), .Z(n60797) );
  NOR U81061 ( .A(n66244), .B(n60797), .Z(n63380) );
  IV U81062 ( .A(n60798), .Z(n60800) );
  NOR U81063 ( .A(n60800), .B(n60799), .Z(n68737) );
  NOR U81064 ( .A(n60801), .B(n66250), .Z(n60802) );
  NOR U81065 ( .A(n68737), .B(n60802), .Z(n63379) );
  IV U81066 ( .A(n60803), .Z(n60804) );
  NOR U81067 ( .A(n60805), .B(n60804), .Z(n60806) );
  IV U81068 ( .A(n60806), .Z(n66253) );
  IV U81069 ( .A(n60807), .Z(n60808) );
  NOR U81070 ( .A(n60809), .B(n60808), .Z(n60810) );
  IV U81071 ( .A(n60810), .Z(n63364) );
  IV U81072 ( .A(n60811), .Z(n60812) );
  NOR U81073 ( .A(n60812), .B(n63362), .Z(n63356) );
  IV U81074 ( .A(n63356), .Z(n63348) );
  IV U81075 ( .A(n60813), .Z(n60815) );
  NOR U81076 ( .A(n60815), .B(n60814), .Z(n63352) );
  IV U81077 ( .A(n63352), .Z(n68722) );
  IV U81078 ( .A(n60816), .Z(n60817) );
  NOR U81079 ( .A(n60818), .B(n60817), .Z(n71212) );
  IV U81080 ( .A(n60819), .Z(n60822) );
  IV U81081 ( .A(n60820), .Z(n60821) );
  NOR U81082 ( .A(n60822), .B(n60821), .Z(n71217) );
  NOR U81083 ( .A(n71212), .B(n71217), .Z(n68720) );
  IV U81084 ( .A(n60823), .Z(n60825) );
  IV U81085 ( .A(n60824), .Z(n63344) );
  NOR U81086 ( .A(n60825), .B(n63344), .Z(n63341) );
  IV U81087 ( .A(n63341), .Z(n63329) );
  IV U81088 ( .A(n60826), .Z(n60827) );
  NOR U81089 ( .A(n68707), .B(n60827), .Z(n60829) );
  IV U81090 ( .A(n66264), .Z(n60828) );
  NOR U81091 ( .A(n60828), .B(n66263), .Z(n68712) );
  NOR U81092 ( .A(n60829), .B(n68712), .Z(n63328) );
  IV U81093 ( .A(n60830), .Z(n60831) );
  NOR U81094 ( .A(n60831), .B(n60833), .Z(n66276) );
  IV U81095 ( .A(n60832), .Z(n60834) );
  NOR U81096 ( .A(n60834), .B(n60833), .Z(n66270) );
  NOR U81097 ( .A(n66276), .B(n66270), .Z(n60835) );
  IV U81098 ( .A(n60835), .Z(n60836) );
  NOR U81099 ( .A(n68708), .B(n60836), .Z(n63326) );
  IV U81100 ( .A(n60837), .Z(n60839) );
  NOR U81101 ( .A(n60839), .B(n60838), .Z(n66278) );
  IV U81102 ( .A(n60840), .Z(n60842) );
  NOR U81103 ( .A(n60842), .B(n60841), .Z(n66274) );
  NOR U81104 ( .A(n66278), .B(n66274), .Z(n63325) );
  IV U81105 ( .A(n60843), .Z(n60845) );
  NOR U81106 ( .A(n60845), .B(n60844), .Z(n66286) );
  IV U81107 ( .A(n60846), .Z(n60848) );
  NOR U81108 ( .A(n60848), .B(n60847), .Z(n66281) );
  NOR U81109 ( .A(n66286), .B(n66281), .Z(n63324) );
  IV U81110 ( .A(n60849), .Z(n60850) );
  NOR U81111 ( .A(n60851), .B(n60850), .Z(n66283) );
  IV U81112 ( .A(n60852), .Z(n63322) );
  IV U81113 ( .A(n60853), .Z(n60854) );
  NOR U81114 ( .A(n63322), .B(n60854), .Z(n66289) );
  IV U81115 ( .A(n60855), .Z(n60857) );
  NOR U81116 ( .A(n60857), .B(n60856), .Z(n68695) );
  IV U81117 ( .A(n60858), .Z(n60859) );
  NOR U81118 ( .A(n60859), .B(n63318), .Z(n66298) );
  NOR U81119 ( .A(n68695), .B(n66298), .Z(n63316) );
  NOR U81120 ( .A(n60860), .B(n71251), .Z(n68687) );
  IV U81121 ( .A(n60861), .Z(n60862) );
  NOR U81122 ( .A(n60863), .B(n60862), .Z(n68693) );
  NOR U81123 ( .A(n68687), .B(n68693), .Z(n63315) );
  IV U81124 ( .A(n60864), .Z(n60868) );
  IV U81125 ( .A(n60865), .Z(n63302) );
  NOR U81126 ( .A(n60866), .B(n63302), .Z(n60867) );
  IV U81127 ( .A(n60867), .Z(n63305) );
  NOR U81128 ( .A(n60868), .B(n63305), .Z(n63299) );
  IV U81129 ( .A(n63299), .Z(n63289) );
  IV U81130 ( .A(n60869), .Z(n60870) );
  NOR U81131 ( .A(n60871), .B(n60870), .Z(n66304) );
  IV U81132 ( .A(n60872), .Z(n63286) );
  IV U81133 ( .A(n60873), .Z(n60874) );
  NOR U81134 ( .A(n63286), .B(n60874), .Z(n66309) );
  IV U81135 ( .A(n60875), .Z(n60876) );
  NOR U81136 ( .A(n60876), .B(n63283), .Z(n68659) );
  IV U81137 ( .A(n60877), .Z(n63261) );
  IV U81138 ( .A(n60878), .Z(n60880) );
  NOR U81139 ( .A(n60880), .B(n60879), .Z(n66334) );
  IV U81140 ( .A(n60881), .Z(n60888) );
  IV U81141 ( .A(n60882), .Z(n60883) );
  NOR U81142 ( .A(n60888), .B(n60883), .Z(n60884) );
  IV U81143 ( .A(n60884), .Z(n66338) );
  IV U81144 ( .A(n60885), .Z(n60886) );
  NOR U81145 ( .A(n60886), .B(n60891), .Z(n68645) );
  IV U81146 ( .A(n60887), .Z(n60889) );
  NOR U81147 ( .A(n60889), .B(n60888), .Z(n66343) );
  NOR U81148 ( .A(n68645), .B(n66343), .Z(n63247) );
  IV U81149 ( .A(n60890), .Z(n60892) );
  NOR U81150 ( .A(n60892), .B(n60891), .Z(n68642) );
  IV U81151 ( .A(n60893), .Z(n60898) );
  IV U81152 ( .A(n60894), .Z(n60895) );
  NOR U81153 ( .A(n60898), .B(n60895), .Z(n66345) );
  IV U81154 ( .A(n60896), .Z(n60897) );
  NOR U81155 ( .A(n60898), .B(n60897), .Z(n68635) );
  IV U81156 ( .A(n60899), .Z(n60900) );
  NOR U81157 ( .A(n63244), .B(n60900), .Z(n60901) );
  IV U81158 ( .A(n60901), .Z(n66349) );
  IV U81159 ( .A(n60902), .Z(n60904) );
  IV U81160 ( .A(n60903), .Z(n63238) );
  NOR U81161 ( .A(n60904), .B(n63238), .Z(n68626) );
  IV U81162 ( .A(n60905), .Z(n60906) );
  NOR U81163 ( .A(n60911), .B(n60906), .Z(n66356) );
  IV U81164 ( .A(n60907), .Z(n60909) );
  IV U81165 ( .A(n60908), .Z(n60916) );
  NOR U81166 ( .A(n60909), .B(n60916), .Z(n66359) );
  IV U81167 ( .A(n60910), .Z(n60912) );
  NOR U81168 ( .A(n60912), .B(n60911), .Z(n68613) );
  NOR U81169 ( .A(n66359), .B(n68613), .Z(n60913) );
  IV U81170 ( .A(n60913), .Z(n63236) );
  IV U81171 ( .A(n60914), .Z(n60915) );
  NOR U81172 ( .A(n60916), .B(n60915), .Z(n68605) );
  IV U81173 ( .A(n60917), .Z(n60918) );
  NOR U81174 ( .A(n60919), .B(n60918), .Z(n68593) );
  NOR U81175 ( .A(n66369), .B(n68593), .Z(n63229) );
  IV U81176 ( .A(n60920), .Z(n60921) );
  NOR U81177 ( .A(n60921), .B(n63224), .Z(n66366) );
  IV U81178 ( .A(n60922), .Z(n60923) );
  NOR U81179 ( .A(n60923), .B(n60929), .Z(n66389) );
  IV U81180 ( .A(n60924), .Z(n60926) );
  NOR U81181 ( .A(n60926), .B(n60925), .Z(n66384) );
  NOR U81182 ( .A(n66389), .B(n66384), .Z(n63205) );
  IV U81183 ( .A(n60930), .Z(n60927) );
  NOR U81184 ( .A(n60927), .B(n60929), .Z(n66395) );
  IV U81185 ( .A(n60928), .Z(n60932) );
  XOR U81186 ( .A(n60930), .B(n60929), .Z(n60931) );
  NOR U81187 ( .A(n60932), .B(n60931), .Z(n66393) );
  NOR U81188 ( .A(n66395), .B(n66393), .Z(n63204) );
  IV U81189 ( .A(n60933), .Z(n60935) );
  NOR U81190 ( .A(n60935), .B(n60934), .Z(n68579) );
  IV U81191 ( .A(n60936), .Z(n60938) );
  NOR U81192 ( .A(n60938), .B(n60937), .Z(n68582) );
  NOR U81193 ( .A(n68579), .B(n68582), .Z(n63203) );
  IV U81194 ( .A(n60939), .Z(n60941) );
  IV U81195 ( .A(n60940), .Z(n60943) );
  NOR U81196 ( .A(n60941), .B(n60943), .Z(n68576) );
  IV U81197 ( .A(n60942), .Z(n60944) );
  NOR U81198 ( .A(n60944), .B(n60943), .Z(n66398) );
  IV U81199 ( .A(n60945), .Z(n60947) );
  NOR U81200 ( .A(n60947), .B(n60946), .Z(n66422) );
  IV U81201 ( .A(n60948), .Z(n60949) );
  NOR U81202 ( .A(n60950), .B(n60949), .Z(n66417) );
  NOR U81203 ( .A(n66422), .B(n66417), .Z(n63190) );
  IV U81204 ( .A(n60951), .Z(n60952) );
  NOR U81205 ( .A(n60953), .B(n60952), .Z(n66425) );
  IV U81206 ( .A(n60954), .Z(n60955) );
  NOR U81207 ( .A(n60956), .B(n60955), .Z(n66420) );
  NOR U81208 ( .A(n66425), .B(n66420), .Z(n63189) );
  IV U81209 ( .A(n60957), .Z(n60958) );
  IV U81210 ( .A(n63183), .Z(n63181) );
  NOR U81211 ( .A(n60958), .B(n63181), .Z(n68567) );
  IV U81212 ( .A(n60959), .Z(n60960) );
  NOR U81213 ( .A(n60961), .B(n60960), .Z(n66428) );
  NOR U81214 ( .A(n68567), .B(n66428), .Z(n63188) );
  NOR U81215 ( .A(n60962), .B(n71355), .Z(n68557) );
  IV U81216 ( .A(n60963), .Z(n60965) );
  NOR U81217 ( .A(n60965), .B(n60964), .Z(n71350) );
  IV U81218 ( .A(n60966), .Z(n60967) );
  NOR U81219 ( .A(n60967), .B(n63127), .Z(n71390) );
  IV U81220 ( .A(n60968), .Z(n60970) );
  NOR U81221 ( .A(n60970), .B(n60969), .Z(n71386) );
  NOR U81222 ( .A(n71390), .B(n71386), .Z(n68537) );
  NOR U81223 ( .A(n60972), .B(n60971), .Z(n66481) );
  IV U81224 ( .A(n60973), .Z(n60974) );
  NOR U81225 ( .A(n60975), .B(n60974), .Z(n68505) );
  IV U81226 ( .A(n60976), .Z(n60977) );
  NOR U81227 ( .A(n60977), .B(n60980), .Z(n68511) );
  NOR U81228 ( .A(n68505), .B(n68511), .Z(n66484) );
  IV U81229 ( .A(n60978), .Z(n60979) );
  NOR U81230 ( .A(n60980), .B(n60979), .Z(n66485) );
  NOR U81231 ( .A(n60981), .B(n68493), .Z(n60985) );
  IV U81232 ( .A(n60982), .Z(n60983) );
  NOR U81233 ( .A(n60984), .B(n60983), .Z(n68499) );
  NOR U81234 ( .A(n60985), .B(n68499), .Z(n63083) );
  IV U81235 ( .A(n60986), .Z(n60987) );
  NOR U81236 ( .A(n60988), .B(n60987), .Z(n63081) );
  IV U81237 ( .A(n63081), .Z(n63072) );
  IV U81238 ( .A(n60989), .Z(n60992) );
  NOR U81239 ( .A(n60990), .B(n60994), .Z(n60991) );
  IV U81240 ( .A(n60991), .Z(n63044) );
  NOR U81241 ( .A(n60992), .B(n63044), .Z(n66499) );
  IV U81242 ( .A(n60993), .Z(n60997) );
  NOR U81243 ( .A(n60995), .B(n60994), .Z(n60996) );
  IV U81244 ( .A(n60996), .Z(n60999) );
  NOR U81245 ( .A(n60997), .B(n60999), .Z(n68472) );
  NOR U81246 ( .A(n66499), .B(n68472), .Z(n63042) );
  IV U81247 ( .A(n60998), .Z(n61000) );
  NOR U81248 ( .A(n61000), .B(n60999), .Z(n68469) );
  IV U81249 ( .A(n61001), .Z(n61003) );
  NOR U81250 ( .A(n61003), .B(n61002), .Z(n71464) );
  IV U81251 ( .A(n61004), .Z(n61005) );
  NOR U81252 ( .A(n61006), .B(n61005), .Z(n71460) );
  NOR U81253 ( .A(n71464), .B(n71460), .Z(n68463) );
  IV U81254 ( .A(n61007), .Z(n61008) );
  NOR U81255 ( .A(n61009), .B(n61008), .Z(n68464) );
  IV U81256 ( .A(n61010), .Z(n61017) );
  IV U81257 ( .A(n61011), .Z(n61012) );
  NOR U81258 ( .A(n61017), .B(n61012), .Z(n66504) );
  NOR U81259 ( .A(n68464), .B(n66504), .Z(n63041) );
  IV U81260 ( .A(n61013), .Z(n61014) );
  NOR U81261 ( .A(n61017), .B(n61014), .Z(n66501) );
  IV U81262 ( .A(n61015), .Z(n61016) );
  NOR U81263 ( .A(n61017), .B(n61016), .Z(n68457) );
  IV U81264 ( .A(n61018), .Z(n61019) );
  NOR U81265 ( .A(n63038), .B(n61019), .Z(n68454) );
  IV U81266 ( .A(n61020), .Z(n61022) );
  NOR U81267 ( .A(n61022), .B(n61021), .Z(n61023) );
  IV U81268 ( .A(n61023), .Z(n66510) );
  IV U81269 ( .A(n61027), .Z(n61025) );
  NOR U81270 ( .A(n61025), .B(n61024), .Z(n66518) );
  NOR U81271 ( .A(n61027), .B(n61026), .Z(n61030) );
  IV U81272 ( .A(n61028), .Z(n61029) );
  NOR U81273 ( .A(n61030), .B(n61029), .Z(n66515) );
  NOR U81274 ( .A(n66518), .B(n66515), .Z(n63033) );
  IV U81275 ( .A(n61031), .Z(n61033) );
  NOR U81276 ( .A(n61033), .B(n61032), .Z(n66528) );
  NOR U81277 ( .A(n61034), .B(n66522), .Z(n61035) );
  NOR U81278 ( .A(n66528), .B(n61035), .Z(n63032) );
  NOR U81279 ( .A(n61036), .B(n66533), .Z(n63027) );
  IV U81280 ( .A(n61037), .Z(n61039) );
  NOR U81281 ( .A(n61039), .B(n61038), .Z(n63024) );
  IV U81282 ( .A(n63024), .Z(n63019) );
  IV U81283 ( .A(n61040), .Z(n61043) );
  IV U81284 ( .A(n61041), .Z(n61042) );
  NOR U81285 ( .A(n61043), .B(n61042), .Z(n68446) );
  IV U81286 ( .A(n61044), .Z(n61045) );
  NOR U81287 ( .A(n61052), .B(n61045), .Z(n61046) );
  IV U81288 ( .A(n61046), .Z(n66539) );
  IV U81289 ( .A(n61047), .Z(n61048) );
  NOR U81290 ( .A(n61052), .B(n61048), .Z(n61049) );
  IV U81291 ( .A(n61049), .Z(n68445) );
  IV U81292 ( .A(n61050), .Z(n61051) );
  NOR U81293 ( .A(n61052), .B(n61051), .Z(n68441) );
  IV U81294 ( .A(n61053), .Z(n61055) );
  IV U81295 ( .A(n61054), .Z(n63016) );
  NOR U81296 ( .A(n61055), .B(n63016), .Z(n66544) );
  IV U81297 ( .A(n61056), .Z(n61061) );
  NOR U81298 ( .A(n61068), .B(n63016), .Z(n61057) );
  IV U81299 ( .A(n61057), .Z(n61058) );
  NOR U81300 ( .A(n61059), .B(n61058), .Z(n61060) );
  IV U81301 ( .A(n61060), .Z(n61063) );
  NOR U81302 ( .A(n61061), .B(n61063), .Z(n66547) );
  IV U81303 ( .A(n61062), .Z(n61064) );
  NOR U81304 ( .A(n61064), .B(n61063), .Z(n66550) );
  NOR U81305 ( .A(n63008), .B(n61065), .Z(n61066) );
  IV U81306 ( .A(n61066), .Z(n61067) );
  NOR U81307 ( .A(n61068), .B(n61067), .Z(n66556) );
  NOR U81308 ( .A(n66550), .B(n66556), .Z(n63014) );
  IV U81309 ( .A(n61069), .Z(n61070) );
  NOR U81310 ( .A(n62997), .B(n61070), .Z(n66559) );
  IV U81311 ( .A(n61071), .Z(n61072) );
  NOR U81312 ( .A(n61073), .B(n61072), .Z(n66566) );
  IV U81313 ( .A(n61074), .Z(n61075) );
  NOR U81314 ( .A(n61078), .B(n61075), .Z(n68412) );
  IV U81315 ( .A(n61076), .Z(n61077) );
  NOR U81316 ( .A(n61078), .B(n61077), .Z(n68409) );
  IV U81317 ( .A(n61079), .Z(n61081) );
  IV U81318 ( .A(n61080), .Z(n62974) );
  NOR U81319 ( .A(n61081), .B(n62974), .Z(n68406) );
  NOR U81320 ( .A(n68409), .B(n68406), .Z(n62976) );
  IV U81321 ( .A(n61082), .Z(n61083) );
  NOR U81322 ( .A(n61084), .B(n61083), .Z(n66575) );
  IV U81323 ( .A(n61085), .Z(n61086) );
  NOR U81324 ( .A(n62968), .B(n61086), .Z(n66573) );
  NOR U81325 ( .A(n66575), .B(n66573), .Z(n62966) );
  IV U81326 ( .A(n61087), .Z(n61089) );
  NOR U81327 ( .A(n61089), .B(n61088), .Z(n68396) );
  NOR U81328 ( .A(n61090), .B(n66579), .Z(n61091) );
  NOR U81329 ( .A(n68396), .B(n61091), .Z(n61092) );
  IV U81330 ( .A(n61092), .Z(n62965) );
  IV U81331 ( .A(n61093), .Z(n61094) );
  NOR U81332 ( .A(n61095), .B(n61094), .Z(n66585) );
  IV U81333 ( .A(n61096), .Z(n61098) );
  IV U81334 ( .A(n61097), .Z(n62953) );
  NOR U81335 ( .A(n61098), .B(n62953), .Z(n66589) );
  NOR U81336 ( .A(n66585), .B(n66589), .Z(n62964) );
  IV U81337 ( .A(n61099), .Z(n61101) );
  IV U81338 ( .A(n61100), .Z(n61108) );
  NOR U81339 ( .A(n61101), .B(n61108), .Z(n68380) );
  IV U81340 ( .A(n61102), .Z(n61104) );
  NOR U81341 ( .A(n61104), .B(n61103), .Z(n68387) );
  NOR U81342 ( .A(n68380), .B(n68387), .Z(n62951) );
  IV U81343 ( .A(n61105), .Z(n61106) );
  NOR U81344 ( .A(n61106), .B(n61111), .Z(n66602) );
  IV U81345 ( .A(n61107), .Z(n61109) );
  NOR U81346 ( .A(n61109), .B(n61108), .Z(n68382) );
  NOR U81347 ( .A(n66602), .B(n68382), .Z(n62950) );
  IV U81348 ( .A(n61110), .Z(n61112) );
  NOR U81349 ( .A(n61112), .B(n61111), .Z(n66599) );
  IV U81350 ( .A(n61113), .Z(n61115) );
  NOR U81351 ( .A(n61115), .B(n61114), .Z(n66605) );
  IV U81352 ( .A(n61116), .Z(n61117) );
  NOR U81353 ( .A(n61118), .B(n61117), .Z(n66607) );
  NOR U81354 ( .A(n66605), .B(n66607), .Z(n62949) );
  NOR U81355 ( .A(n61119), .B(n66619), .Z(n61123) );
  IV U81356 ( .A(n61120), .Z(n61121) );
  NOR U81357 ( .A(n61122), .B(n61121), .Z(n66616) );
  NOR U81358 ( .A(n61123), .B(n66616), .Z(n62942) );
  IV U81359 ( .A(n61124), .Z(n66636) );
  IV U81360 ( .A(n66632), .Z(n61131) );
  NOR U81361 ( .A(n66636), .B(n61131), .Z(n61128) );
  IV U81362 ( .A(n61125), .Z(n61127) );
  NOR U81363 ( .A(n61127), .B(n61126), .Z(n66626) );
  NOR U81364 ( .A(n61128), .B(n66626), .Z(n62941) );
  IV U81365 ( .A(n66629), .Z(n61129) );
  NOR U81366 ( .A(n61129), .B(n61131), .Z(n66637) );
  NOR U81367 ( .A(n61130), .B(n66642), .Z(n61133) );
  IV U81368 ( .A(n66630), .Z(n61132) );
  NOR U81369 ( .A(n61132), .B(n61131), .Z(n68372) );
  NOR U81370 ( .A(n61133), .B(n68372), .Z(n62940) );
  IV U81371 ( .A(n61134), .Z(n61136) );
  NOR U81372 ( .A(n61136), .B(n61135), .Z(n66649) );
  IV U81373 ( .A(n61137), .Z(n61138) );
  NOR U81374 ( .A(n61139), .B(n61138), .Z(n68369) );
  NOR U81375 ( .A(n66649), .B(n68369), .Z(n62939) );
  IV U81376 ( .A(n61140), .Z(n61141) );
  NOR U81377 ( .A(n61141), .B(n62935), .Z(n66646) );
  IV U81378 ( .A(n61142), .Z(n61144) );
  IV U81379 ( .A(n61143), .Z(n61146) );
  NOR U81380 ( .A(n61144), .B(n61146), .Z(n66654) );
  IV U81381 ( .A(n61145), .Z(n61147) );
  NOR U81382 ( .A(n61147), .B(n61146), .Z(n66660) );
  IV U81383 ( .A(n61148), .Z(n61149) );
  NOR U81384 ( .A(n61149), .B(n61151), .Z(n66662) );
  IV U81385 ( .A(n61150), .Z(n61152) );
  NOR U81386 ( .A(n61152), .B(n61151), .Z(n68348) );
  XOR U81387 ( .A(n66662), .B(n68348), .Z(n61153) );
  NOR U81388 ( .A(n66660), .B(n61153), .Z(n62930) );
  IV U81389 ( .A(n61154), .Z(n61155) );
  NOR U81390 ( .A(n61156), .B(n61155), .Z(n68353) );
  IV U81391 ( .A(n61157), .Z(n61159) );
  NOR U81392 ( .A(n61159), .B(n61158), .Z(n66664) );
  NOR U81393 ( .A(n68353), .B(n66664), .Z(n62929) );
  IV U81394 ( .A(n61160), .Z(n61161) );
  NOR U81395 ( .A(n61161), .B(n61163), .Z(n66666) );
  IV U81396 ( .A(n61162), .Z(n61164) );
  NOR U81397 ( .A(n61164), .B(n61163), .Z(n68344) );
  NOR U81398 ( .A(n66666), .B(n68344), .Z(n62928) );
  IV U81399 ( .A(n61165), .Z(n61166) );
  NOR U81400 ( .A(n61167), .B(n61166), .Z(n66669) );
  IV U81401 ( .A(n61168), .Z(n61169) );
  NOR U81402 ( .A(n61175), .B(n61169), .Z(n66671) );
  NOR U81403 ( .A(n66669), .B(n66671), .Z(n62927) );
  IV U81404 ( .A(n61170), .Z(n61171) );
  NOR U81405 ( .A(n61172), .B(n61171), .Z(n68338) );
  IV U81406 ( .A(n61173), .Z(n61174) );
  NOR U81407 ( .A(n61175), .B(n61174), .Z(n68341) );
  NOR U81408 ( .A(n68338), .B(n68341), .Z(n62926) );
  IV U81409 ( .A(n61176), .Z(n61177) );
  NOR U81410 ( .A(n61177), .B(n62904), .Z(n61178) );
  IV U81411 ( .A(n61178), .Z(n68318) );
  IV U81412 ( .A(n61179), .Z(n61180) );
  NOR U81413 ( .A(n61181), .B(n61180), .Z(n66684) );
  IV U81414 ( .A(n61182), .Z(n61187) );
  IV U81415 ( .A(n61183), .Z(n61184) );
  NOR U81416 ( .A(n61187), .B(n61184), .Z(n66690) );
  NOR U81417 ( .A(n66684), .B(n66690), .Z(n62902) );
  IV U81418 ( .A(n61185), .Z(n61186) );
  NOR U81419 ( .A(n61187), .B(n61186), .Z(n66687) );
  IV U81420 ( .A(n61188), .Z(n61190) );
  NOR U81421 ( .A(n61190), .B(n61189), .Z(n68304) );
  NOR U81422 ( .A(n61191), .B(n68307), .Z(n61192) );
  NOR U81423 ( .A(n68304), .B(n61192), .Z(n62901) );
  IV U81424 ( .A(n61193), .Z(n61194) );
  NOR U81425 ( .A(n61194), .B(n61199), .Z(n66699) );
  IV U81426 ( .A(n61195), .Z(n61196) );
  NOR U81427 ( .A(n61197), .B(n61196), .Z(n66693) );
  NOR U81428 ( .A(n66699), .B(n66693), .Z(n62900) );
  IV U81429 ( .A(n61198), .Z(n61200) );
  NOR U81430 ( .A(n61200), .B(n61199), .Z(n61201) );
  IV U81431 ( .A(n61201), .Z(n61202) );
  NOR U81432 ( .A(n61203), .B(n61202), .Z(n66696) );
  IV U81433 ( .A(n61204), .Z(n61205) );
  NOR U81434 ( .A(n66741), .B(n61205), .Z(n66732) );
  NOR U81435 ( .A(n61206), .B(n66741), .Z(n61212) );
  IV U81436 ( .A(n61207), .Z(n61211) );
  NOR U81437 ( .A(n61209), .B(n61208), .Z(n61210) );
  IV U81438 ( .A(n61210), .Z(n61217) );
  NOR U81439 ( .A(n61211), .B(n61217), .Z(n68267) );
  NOR U81440 ( .A(n61212), .B(n68267), .Z(n62842) );
  IV U81441 ( .A(n61213), .Z(n61215) );
  NOR U81442 ( .A(n61215), .B(n61214), .Z(n66744) );
  IV U81443 ( .A(n61216), .Z(n61218) );
  NOR U81444 ( .A(n61218), .B(n61217), .Z(n68264) );
  NOR U81445 ( .A(n66744), .B(n68264), .Z(n62841) );
  IV U81446 ( .A(n61219), .Z(n61220) );
  NOR U81447 ( .A(n61220), .B(n62830), .Z(n68259) );
  IV U81448 ( .A(n61221), .Z(n61223) );
  NOR U81449 ( .A(n61223), .B(n61222), .Z(n66746) );
  NOR U81450 ( .A(n68259), .B(n66746), .Z(n62840) );
  IV U81451 ( .A(n61224), .Z(n61225) );
  NOR U81452 ( .A(n61226), .B(n61225), .Z(n61227) );
  IV U81453 ( .A(n61227), .Z(n62835) );
  NOR U81454 ( .A(n61228), .B(n66756), .Z(n61232) );
  IV U81455 ( .A(n61229), .Z(n61231) );
  IV U81456 ( .A(n61230), .Z(n62834) );
  NOR U81457 ( .A(n61231), .B(n62834), .Z(n66753) );
  NOR U81458 ( .A(n61232), .B(n66753), .Z(n62828) );
  IV U81459 ( .A(n61233), .Z(n61235) );
  NOR U81460 ( .A(n61235), .B(n61234), .Z(n68241) );
  IV U81461 ( .A(n61236), .Z(n61238) );
  NOR U81462 ( .A(n61238), .B(n61237), .Z(n68251) );
  NOR U81463 ( .A(n68241), .B(n68251), .Z(n62827) );
  IV U81464 ( .A(n61239), .Z(n61240) );
  NOR U81465 ( .A(n61240), .B(n62825), .Z(n66760) );
  IV U81466 ( .A(n61241), .Z(n61243) );
  NOR U81467 ( .A(n61243), .B(n61242), .Z(n61244) );
  IV U81468 ( .A(n61244), .Z(n68232) );
  IV U81469 ( .A(n61245), .Z(n61247) );
  IV U81470 ( .A(n61246), .Z(n61253) );
  NOR U81471 ( .A(n61247), .B(n61253), .Z(n66770) );
  IV U81472 ( .A(n61248), .Z(n61250) );
  NOR U81473 ( .A(n61250), .B(n61249), .Z(n68228) );
  NOR U81474 ( .A(n66770), .B(n68228), .Z(n62815) );
  IV U81475 ( .A(n61251), .Z(n61252) );
  NOR U81476 ( .A(n61253), .B(n61252), .Z(n66767) );
  IV U81477 ( .A(n61254), .Z(n61255) );
  NOR U81478 ( .A(n61256), .B(n61255), .Z(n68214) );
  IV U81479 ( .A(n61257), .Z(n61258) );
  NOR U81480 ( .A(n61258), .B(n61263), .Z(n66781) );
  NOR U81481 ( .A(n68214), .B(n66781), .Z(n62808) );
  IV U81482 ( .A(n61259), .Z(n61260) );
  NOR U81483 ( .A(n61261), .B(n61260), .Z(n66785) );
  IV U81484 ( .A(n61262), .Z(n61264) );
  NOR U81485 ( .A(n61264), .B(n61263), .Z(n66783) );
  NOR U81486 ( .A(n66785), .B(n66783), .Z(n61265) );
  IV U81487 ( .A(n61265), .Z(n62807) );
  IV U81488 ( .A(n61266), .Z(n61267) );
  NOR U81489 ( .A(n61268), .B(n61267), .Z(n66788) );
  IV U81490 ( .A(n61269), .Z(n61270) );
  NOR U81491 ( .A(n61275), .B(n61270), .Z(n66792) );
  NOR U81492 ( .A(n66788), .B(n66792), .Z(n62806) );
  IV U81493 ( .A(n61271), .Z(n61272) );
  NOR U81494 ( .A(n61273), .B(n61272), .Z(n71659) );
  IV U81495 ( .A(n61274), .Z(n61276) );
  NOR U81496 ( .A(n61276), .B(n61275), .Z(n73102) );
  NOR U81497 ( .A(n71659), .B(n73102), .Z(n66791) );
  IV U81498 ( .A(n61277), .Z(n61278) );
  NOR U81499 ( .A(n61279), .B(n61278), .Z(n66799) );
  IV U81500 ( .A(n61280), .Z(n61283) );
  IV U81501 ( .A(n61281), .Z(n61282) );
  NOR U81502 ( .A(n61283), .B(n61282), .Z(n61284) );
  IV U81503 ( .A(n61284), .Z(n66798) );
  IV U81504 ( .A(n61285), .Z(n61286) );
  NOR U81505 ( .A(n61287), .B(n61286), .Z(n61288) );
  NOR U81506 ( .A(n78589), .B(n61288), .Z(n71667) );
  IV U81507 ( .A(n61289), .Z(n61292) );
  NOR U81508 ( .A(n62780), .B(n61290), .Z(n61291) );
  IV U81509 ( .A(n61291), .Z(n62782) );
  NOR U81510 ( .A(n61292), .B(n62782), .Z(n66808) );
  IV U81511 ( .A(n61293), .Z(n61295) );
  IV U81512 ( .A(n61294), .Z(n61298) );
  NOR U81513 ( .A(n61295), .B(n61298), .Z(n62775) );
  NOR U81514 ( .A(n61296), .B(n66824), .Z(n61302) );
  IV U81515 ( .A(n61297), .Z(n61301) );
  NOR U81516 ( .A(n61299), .B(n61298), .Z(n61300) );
  IV U81517 ( .A(n61300), .Z(n62771) );
  NOR U81518 ( .A(n61301), .B(n62771), .Z(n66820) );
  NOR U81519 ( .A(n61302), .B(n66820), .Z(n62768) );
  IV U81520 ( .A(n61303), .Z(n61305) );
  IV U81521 ( .A(n61304), .Z(n62761) );
  NOR U81522 ( .A(n61305), .B(n62761), .Z(n66832) );
  IV U81523 ( .A(n61306), .Z(n61308) );
  IV U81524 ( .A(n61307), .Z(n61310) );
  NOR U81525 ( .A(n61308), .B(n61310), .Z(n66842) );
  IV U81526 ( .A(n61309), .Z(n61313) );
  NOR U81527 ( .A(n61311), .B(n61310), .Z(n61312) );
  IV U81528 ( .A(n61312), .Z(n61315) );
  NOR U81529 ( .A(n61313), .B(n61315), .Z(n68193) );
  NOR U81530 ( .A(n66842), .B(n68193), .Z(n62757) );
  IV U81531 ( .A(n61314), .Z(n61316) );
  NOR U81532 ( .A(n61316), .B(n61315), .Z(n62752) );
  IV U81533 ( .A(n61317), .Z(n61318) );
  NOR U81534 ( .A(n61318), .B(n61323), .Z(n66851) );
  IV U81535 ( .A(n61319), .Z(n61321) );
  NOR U81536 ( .A(n61321), .B(n61320), .Z(n66857) );
  IV U81537 ( .A(n61322), .Z(n61324) );
  NOR U81538 ( .A(n61324), .B(n61323), .Z(n66855) );
  NOR U81539 ( .A(n66857), .B(n66855), .Z(n62745) );
  IV U81540 ( .A(n61325), .Z(n61327) );
  IV U81541 ( .A(n61326), .Z(n61329) );
  NOR U81542 ( .A(n61327), .B(n61329), .Z(n66860) );
  IV U81543 ( .A(n61328), .Z(n61330) );
  NOR U81544 ( .A(n61330), .B(n61329), .Z(n68182) );
  IV U81545 ( .A(n61331), .Z(n61332) );
  NOR U81546 ( .A(n61333), .B(n61332), .Z(n68145) );
  IV U81547 ( .A(n61334), .Z(n61335) );
  NOR U81548 ( .A(n61336), .B(n61335), .Z(n68155) );
  NOR U81549 ( .A(n68145), .B(n68155), .Z(n61337) );
  IV U81550 ( .A(n61337), .Z(n62702) );
  IV U81551 ( .A(n61338), .Z(n61339) );
  NOR U81552 ( .A(n62701), .B(n61339), .Z(n66890) );
  IV U81553 ( .A(n61340), .Z(n61342) );
  IV U81554 ( .A(n61341), .Z(n61345) );
  NOR U81555 ( .A(n61342), .B(n61345), .Z(n61343) );
  IV U81556 ( .A(n61343), .Z(n68132) );
  IV U81557 ( .A(n61344), .Z(n61346) );
  NOR U81558 ( .A(n61346), .B(n61345), .Z(n66917) );
  IV U81559 ( .A(n61347), .Z(n61348) );
  NOR U81560 ( .A(n61351), .B(n61348), .Z(n68122) );
  IV U81561 ( .A(n61349), .Z(n61350) );
  NOR U81562 ( .A(n61351), .B(n61350), .Z(n68119) );
  IV U81563 ( .A(n61352), .Z(n61353) );
  NOR U81564 ( .A(n61354), .B(n61353), .Z(n72942) );
  IV U81565 ( .A(n61355), .Z(n61357) );
  NOR U81566 ( .A(n61357), .B(n61356), .Z(n72948) );
  NOR U81567 ( .A(n72942), .B(n72948), .Z(n66920) );
  IV U81568 ( .A(n61358), .Z(n61359) );
  NOR U81569 ( .A(n62618), .B(n61359), .Z(n66925) );
  IV U81570 ( .A(n61360), .Z(n61361) );
  NOR U81571 ( .A(n61361), .B(n61373), .Z(n66933) );
  XOR U81572 ( .A(n61363), .B(n61362), .Z(n61365) );
  IV U81573 ( .A(n61364), .Z(n62620) );
  NOR U81574 ( .A(n61365), .B(n62620), .Z(n61366) );
  IV U81575 ( .A(n61366), .Z(n61367) );
  NOR U81576 ( .A(n61368), .B(n61367), .Z(n68067) );
  NOR U81577 ( .A(n66933), .B(n68067), .Z(n62615) );
  IV U81578 ( .A(n61369), .Z(n61371) );
  NOR U81579 ( .A(n61371), .B(n61370), .Z(n66936) );
  IV U81580 ( .A(n61372), .Z(n61374) );
  NOR U81581 ( .A(n61374), .B(n61373), .Z(n68062) );
  NOR U81582 ( .A(n66936), .B(n68062), .Z(n62614) );
  IV U81583 ( .A(n61375), .Z(n61379) );
  IV U81584 ( .A(n61376), .Z(n62605) );
  NOR U81585 ( .A(n61377), .B(n62605), .Z(n61378) );
  IV U81586 ( .A(n61378), .Z(n62612) );
  NOR U81587 ( .A(n61379), .B(n62612), .Z(n66942) );
  IV U81588 ( .A(n61380), .Z(n61381) );
  NOR U81589 ( .A(n61381), .B(n62590), .Z(n68045) );
  NOR U81590 ( .A(n68045), .B(n68057), .Z(n62604) );
  IV U81591 ( .A(n61382), .Z(n61383) );
  NOR U81592 ( .A(n62564), .B(n61383), .Z(n62570) );
  IV U81593 ( .A(n61384), .Z(n61386) );
  IV U81594 ( .A(n61385), .Z(n62566) );
  NOR U81595 ( .A(n61386), .B(n62566), .Z(n62558) );
  NOR U81596 ( .A(n61388), .B(n61387), .Z(n68025) );
  IV U81597 ( .A(n61389), .Z(n61390) );
  NOR U81598 ( .A(n61390), .B(n61392), .Z(n68011) );
  NOR U81599 ( .A(n68018), .B(n68011), .Z(n62556) );
  IV U81600 ( .A(n61391), .Z(n61395) );
  NOR U81601 ( .A(n61393), .B(n61392), .Z(n61394) );
  IV U81602 ( .A(n61394), .Z(n66969) );
  NOR U81603 ( .A(n61395), .B(n66969), .Z(n62555) );
  IV U81604 ( .A(n61396), .Z(n61398) );
  IV U81605 ( .A(n61397), .Z(n61403) );
  NOR U81606 ( .A(n61398), .B(n61403), .Z(n67980) );
  IV U81607 ( .A(n61399), .Z(n61401) );
  XOR U81608 ( .A(n61402), .B(n61403), .Z(n61400) );
  NOR U81609 ( .A(n61401), .B(n61400), .Z(n67986) );
  NOR U81610 ( .A(n67980), .B(n67986), .Z(n62528) );
  IV U81611 ( .A(n61402), .Z(n61404) );
  NOR U81612 ( .A(n61404), .B(n61403), .Z(n67982) );
  NOR U81613 ( .A(n67967), .B(n67982), .Z(n62527) );
  IV U81614 ( .A(n61405), .Z(n61406) );
  NOR U81615 ( .A(n61407), .B(n61406), .Z(n67961) );
  IV U81616 ( .A(n61408), .Z(n61410) );
  NOR U81617 ( .A(n61410), .B(n61409), .Z(n67959) );
  NOR U81618 ( .A(n67961), .B(n67959), .Z(n62525) );
  IV U81619 ( .A(n61411), .Z(n61413) );
  NOR U81620 ( .A(n61413), .B(n61412), .Z(n67956) );
  IV U81621 ( .A(n61414), .Z(n61417) );
  NOR U81622 ( .A(n61415), .B(n61419), .Z(n61416) );
  IV U81623 ( .A(n61416), .Z(n62517) );
  NOR U81624 ( .A(n61417), .B(n62517), .Z(n67953) );
  NOR U81625 ( .A(n67956), .B(n67953), .Z(n62524) );
  IV U81626 ( .A(n61418), .Z(n61420) );
  NOR U81627 ( .A(n61420), .B(n61419), .Z(n61421) );
  IV U81628 ( .A(n61421), .Z(n62519) );
  IV U81629 ( .A(n61422), .Z(n61424) );
  IV U81630 ( .A(n61423), .Z(n62514) );
  NOR U81631 ( .A(n61424), .B(n62514), .Z(n66984) );
  IV U81632 ( .A(n61425), .Z(n61426) );
  NOR U81633 ( .A(n61427), .B(n61426), .Z(n62505) );
  IV U81634 ( .A(n62505), .Z(n62499) );
  IV U81635 ( .A(n61428), .Z(n61429) );
  NOR U81636 ( .A(n61430), .B(n61429), .Z(n67940) );
  IV U81637 ( .A(n61431), .Z(n67934) );
  NOR U81638 ( .A(n67934), .B(n61432), .Z(n62479) );
  IV U81639 ( .A(n61433), .Z(n61435) );
  NOR U81640 ( .A(n61435), .B(n61434), .Z(n66998) );
  IV U81641 ( .A(n61436), .Z(n61437) );
  NOR U81642 ( .A(n61437), .B(n61439), .Z(n67927) );
  IV U81643 ( .A(n61438), .Z(n61440) );
  NOR U81644 ( .A(n61440), .B(n61439), .Z(n67000) );
  NOR U81645 ( .A(n67927), .B(n67000), .Z(n61441) );
  IV U81646 ( .A(n61441), .Z(n62478) );
  IV U81647 ( .A(n61442), .Z(n61444) );
  IV U81648 ( .A(n61443), .Z(n62473) );
  NOR U81649 ( .A(n61444), .B(n62473), .Z(n67920) );
  IV U81650 ( .A(n61445), .Z(n61446) );
  NOR U81651 ( .A(n61446), .B(n62470), .Z(n61447) );
  IV U81652 ( .A(n61447), .Z(n67006) );
  IV U81653 ( .A(n61448), .Z(n61449) );
  NOR U81654 ( .A(n61450), .B(n61449), .Z(n67002) );
  IV U81655 ( .A(n61451), .Z(n67011) );
  IV U81656 ( .A(n61452), .Z(n61453) );
  NOR U81657 ( .A(n67011), .B(n61453), .Z(n67007) );
  XOR U81658 ( .A(n67008), .B(n67007), .Z(n61454) );
  NOR U81659 ( .A(n67002), .B(n61454), .Z(n62468) );
  IV U81660 ( .A(n61455), .Z(n61456) );
  NOR U81661 ( .A(n61456), .B(n61458), .Z(n67023) );
  IV U81662 ( .A(n61457), .Z(n61459) );
  NOR U81663 ( .A(n61459), .B(n61458), .Z(n67020) );
  IV U81664 ( .A(n61460), .Z(n61463) );
  NOR U81665 ( .A(n61466), .B(n62465), .Z(n61461) );
  IV U81666 ( .A(n61461), .Z(n61462) );
  NOR U81667 ( .A(n61463), .B(n61462), .Z(n67903) );
  IV U81668 ( .A(n61464), .Z(n62454) );
  IV U81669 ( .A(n61465), .Z(n61467) );
  NOR U81670 ( .A(n61467), .B(n61466), .Z(n61468) );
  IV U81671 ( .A(n61468), .Z(n62455) );
  NOR U81672 ( .A(n62454), .B(n61469), .Z(n61470) );
  IV U81673 ( .A(n61470), .Z(n67907) );
  IV U81674 ( .A(n61471), .Z(n61473) );
  NOR U81675 ( .A(n61473), .B(n61472), .Z(n67035) );
  IV U81676 ( .A(n61474), .Z(n61475) );
  NOR U81677 ( .A(n61475), .B(n61481), .Z(n61476) );
  IV U81678 ( .A(n61476), .Z(n67033) );
  IV U81679 ( .A(n61477), .Z(n61479) );
  NOR U81680 ( .A(n61479), .B(n61478), .Z(n71853) );
  IV U81681 ( .A(n61480), .Z(n61482) );
  NOR U81682 ( .A(n61482), .B(n61481), .Z(n72783) );
  NOR U81683 ( .A(n71853), .B(n72783), .Z(n67038) );
  IV U81684 ( .A(n61483), .Z(n61488) );
  IV U81685 ( .A(n61484), .Z(n61485) );
  NOR U81686 ( .A(n61488), .B(n61485), .Z(n67042) );
  IV U81687 ( .A(n61486), .Z(n61487) );
  NOR U81688 ( .A(n61488), .B(n61487), .Z(n67039) );
  IV U81689 ( .A(n61489), .Z(n61490) );
  NOR U81690 ( .A(n61499), .B(n61490), .Z(n67046) );
  IV U81691 ( .A(n61491), .Z(n61496) );
  IV U81692 ( .A(n61492), .Z(n61493) );
  NOR U81693 ( .A(n61496), .B(n61493), .Z(n67049) );
  IV U81694 ( .A(n61494), .Z(n61495) );
  NOR U81695 ( .A(n61496), .B(n61495), .Z(n67896) );
  NOR U81696 ( .A(n67049), .B(n67896), .Z(n61497) );
  IV U81697 ( .A(n61497), .Z(n61501) );
  IV U81698 ( .A(n61498), .Z(n61500) );
  NOR U81699 ( .A(n61500), .B(n61499), .Z(n67894) );
  NOR U81700 ( .A(n61501), .B(n67894), .Z(n62449) );
  IV U81701 ( .A(n61502), .Z(n61503) );
  NOR U81702 ( .A(n61503), .B(n62448), .Z(n67055) );
  IV U81703 ( .A(n61504), .Z(n61505) );
  NOR U81704 ( .A(n61506), .B(n61505), .Z(n61507) );
  IV U81705 ( .A(n61507), .Z(n62440) );
  IV U81706 ( .A(n61508), .Z(n61510) );
  NOR U81707 ( .A(n61510), .B(n61509), .Z(n67058) );
  NOR U81708 ( .A(n61511), .B(n67880), .Z(n61512) );
  NOR U81709 ( .A(n67058), .B(n61512), .Z(n62431) );
  IV U81710 ( .A(n61513), .Z(n61518) );
  IV U81711 ( .A(n61514), .Z(n62425) );
  NOR U81712 ( .A(n61515), .B(n62425), .Z(n61516) );
  IV U81713 ( .A(n61516), .Z(n61517) );
  NOR U81714 ( .A(n61518), .B(n61517), .Z(n61519) );
  IV U81715 ( .A(n61519), .Z(n78206) );
  IV U81716 ( .A(n61522), .Z(n61520) );
  NOR U81717 ( .A(n61521), .B(n61520), .Z(n67842) );
  XOR U81718 ( .A(n61522), .B(n61521), .Z(n61525) );
  IV U81719 ( .A(n61523), .Z(n61524) );
  NOR U81720 ( .A(n61525), .B(n61524), .Z(n67845) );
  NOR U81721 ( .A(n67842), .B(n67845), .Z(n62398) );
  IV U81722 ( .A(n61526), .Z(n61531) );
  IV U81723 ( .A(n61527), .Z(n61528) );
  NOR U81724 ( .A(n61531), .B(n61528), .Z(n67839) );
  IV U81725 ( .A(n61529), .Z(n61530) );
  NOR U81726 ( .A(n61531), .B(n61530), .Z(n67064) );
  IV U81727 ( .A(n61532), .Z(n61533) );
  NOR U81728 ( .A(n61533), .B(n61535), .Z(n67070) );
  IV U81729 ( .A(n61534), .Z(n61536) );
  NOR U81730 ( .A(n61536), .B(n61535), .Z(n67068) );
  XOR U81731 ( .A(n67070), .B(n67068), .Z(n61537) );
  NOR U81732 ( .A(n67064), .B(n61537), .Z(n62397) );
  IV U81733 ( .A(n61538), .Z(n61540) );
  NOR U81734 ( .A(n61540), .B(n61539), .Z(n67076) );
  IV U81735 ( .A(n61541), .Z(n61542) );
  NOR U81736 ( .A(n61543), .B(n61542), .Z(n67073) );
  NOR U81737 ( .A(n67076), .B(n67073), .Z(n62396) );
  NOR U81738 ( .A(n61545), .B(n61544), .Z(n67079) );
  IV U81739 ( .A(n61546), .Z(n61551) );
  IV U81740 ( .A(n61547), .Z(n61548) );
  NOR U81741 ( .A(n61551), .B(n61548), .Z(n67815) );
  IV U81742 ( .A(n61549), .Z(n61550) );
  NOR U81743 ( .A(n61551), .B(n61550), .Z(n67084) );
  IV U81744 ( .A(n61552), .Z(n61553) );
  NOR U81745 ( .A(n61554), .B(n61553), .Z(n67811) );
  NOR U81746 ( .A(n67084), .B(n67811), .Z(n62382) );
  IV U81747 ( .A(n61555), .Z(n61558) );
  NOR U81748 ( .A(n61564), .B(n61556), .Z(n61557) );
  IV U81749 ( .A(n61557), .Z(n61560) );
  NOR U81750 ( .A(n61558), .B(n61560), .Z(n67808) );
  IV U81751 ( .A(n61559), .Z(n61561) );
  NOR U81752 ( .A(n61561), .B(n61560), .Z(n67090) );
  IV U81753 ( .A(n61562), .Z(n61563) );
  NOR U81754 ( .A(n61564), .B(n61563), .Z(n67087) );
  IV U81755 ( .A(n61565), .Z(n61568) );
  IV U81756 ( .A(n61566), .Z(n61567) );
  NOR U81757 ( .A(n61568), .B(n61567), .Z(n67803) );
  NOR U81758 ( .A(n61570), .B(n61569), .Z(n67093) );
  IV U81759 ( .A(n61571), .Z(n61572) );
  NOR U81760 ( .A(n61572), .B(n62375), .Z(n67095) );
  NOR U81761 ( .A(n67093), .B(n67095), .Z(n62377) );
  IV U81762 ( .A(n61573), .Z(n61575) );
  NOR U81763 ( .A(n61575), .B(n61574), .Z(n62371) );
  IV U81764 ( .A(n62371), .Z(n62365) );
  IV U81765 ( .A(n61576), .Z(n61578) );
  NOR U81766 ( .A(n61578), .B(n61577), .Z(n67103) );
  IV U81767 ( .A(n61579), .Z(n62346) );
  IV U81768 ( .A(n61580), .Z(n61581) );
  NOR U81769 ( .A(n62346), .B(n61581), .Z(n67107) );
  IV U81770 ( .A(n61582), .Z(n61584) );
  NOR U81771 ( .A(n61584), .B(n61583), .Z(n67783) );
  IV U81772 ( .A(n61585), .Z(n61586) );
  NOR U81773 ( .A(n61587), .B(n61586), .Z(n67778) );
  NOR U81774 ( .A(n67783), .B(n67778), .Z(n67775) );
  IV U81775 ( .A(n61588), .Z(n61589) );
  NOR U81776 ( .A(n61589), .B(n67759), .Z(n67116) );
  NOR U81777 ( .A(n67759), .B(n61590), .Z(n62331) );
  IV U81778 ( .A(n61591), .Z(n61593) );
  NOR U81779 ( .A(n61593), .B(n61592), .Z(n67763) );
  IV U81780 ( .A(n61594), .Z(n61595) );
  NOR U81781 ( .A(n62317), .B(n61595), .Z(n67755) );
  NOR U81782 ( .A(n67763), .B(n67755), .Z(n62330) );
  IV U81783 ( .A(n61596), .Z(n61597) );
  NOR U81784 ( .A(n61597), .B(n62317), .Z(n61598) );
  IV U81785 ( .A(n61598), .Z(n61599) );
  NOR U81786 ( .A(n62315), .B(n61599), .Z(n62326) );
  IV U81787 ( .A(n61600), .Z(n61605) );
  IV U81788 ( .A(n61601), .Z(n61602) );
  NOR U81789 ( .A(n61605), .B(n61602), .Z(n67143) );
  IV U81790 ( .A(n61603), .Z(n61604) );
  NOR U81791 ( .A(n61605), .B(n61604), .Z(n67146) );
  IV U81792 ( .A(n61606), .Z(n61607) );
  NOR U81793 ( .A(n61607), .B(n61609), .Z(n67748) );
  NOR U81794 ( .A(n67146), .B(n67748), .Z(n62300) );
  IV U81795 ( .A(n61608), .Z(n61612) );
  NOR U81796 ( .A(n61610), .B(n61609), .Z(n61611) );
  IV U81797 ( .A(n61611), .Z(n62297) );
  NOR U81798 ( .A(n61612), .B(n62297), .Z(n67745) );
  IV U81799 ( .A(n61613), .Z(n61614) );
  NOR U81800 ( .A(n62291), .B(n61614), .Z(n67738) );
  IV U81801 ( .A(n61615), .Z(n61616) );
  NOR U81802 ( .A(n61617), .B(n61616), .Z(n67154) );
  NOR U81803 ( .A(n61618), .B(n62287), .Z(n67728) );
  NOR U81804 ( .A(n67154), .B(n67728), .Z(n61619) );
  IV U81805 ( .A(n61619), .Z(n62283) );
  IV U81806 ( .A(n61620), .Z(n61621) );
  NOR U81807 ( .A(n61624), .B(n61621), .Z(n61622) );
  IV U81808 ( .A(n61622), .Z(n67158) );
  IV U81809 ( .A(n61623), .Z(n61625) );
  NOR U81810 ( .A(n61625), .B(n61624), .Z(n62277) );
  IV U81811 ( .A(n61626), .Z(n61627) );
  NOR U81812 ( .A(n61628), .B(n61627), .Z(n71980) );
  IV U81813 ( .A(n61629), .Z(n61630) );
  NOR U81814 ( .A(n61630), .B(n62271), .Z(n71974) );
  NOR U81815 ( .A(n71980), .B(n71974), .Z(n67722) );
  IV U81816 ( .A(n61631), .Z(n61635) );
  IV U81817 ( .A(n61632), .Z(n61633) );
  NOR U81818 ( .A(n61635), .B(n61633), .Z(n67161) );
  IV U81819 ( .A(n61634), .Z(n61636) );
  NOR U81820 ( .A(n61636), .B(n61635), .Z(n67164) );
  NOR U81821 ( .A(n67709), .B(n67164), .Z(n62268) );
  IV U81822 ( .A(n61637), .Z(n61642) );
  IV U81823 ( .A(n61638), .Z(n61639) );
  NOR U81824 ( .A(n61642), .B(n61639), .Z(n67694) );
  IV U81825 ( .A(n61640), .Z(n61641) );
  NOR U81826 ( .A(n61642), .B(n61641), .Z(n67690) );
  IV U81827 ( .A(n61643), .Z(n61644) );
  NOR U81828 ( .A(n61644), .B(n61646), .Z(n67687) );
  IV U81829 ( .A(n61645), .Z(n61647) );
  NOR U81830 ( .A(n61647), .B(n61646), .Z(n61648) );
  IV U81831 ( .A(n61648), .Z(n67168) );
  IV U81832 ( .A(n61649), .Z(n61651) );
  NOR U81833 ( .A(n61651), .B(n61650), .Z(n67681) );
  IV U81834 ( .A(n61652), .Z(n61654) );
  NOR U81835 ( .A(n61654), .B(n61653), .Z(n67684) );
  NOR U81836 ( .A(n67681), .B(n67684), .Z(n62242) );
  IV U81837 ( .A(n61655), .Z(n61657) );
  NOR U81838 ( .A(n61657), .B(n61656), .Z(n67678) );
  IV U81839 ( .A(n61658), .Z(n61659) );
  NOR U81840 ( .A(n61659), .B(n62238), .Z(n67671) );
  XOR U81841 ( .A(n67672), .B(n67671), .Z(n61660) );
  NOR U81842 ( .A(n67678), .B(n61660), .Z(n62241) );
  IV U81843 ( .A(n61661), .Z(n61662) );
  NOR U81844 ( .A(n61662), .B(n62232), .Z(n67175) );
  IV U81845 ( .A(n61663), .Z(n61665) );
  NOR U81846 ( .A(n61665), .B(n61664), .Z(n67184) );
  IV U81847 ( .A(n61666), .Z(n61668) );
  NOR U81848 ( .A(n61668), .B(n61667), .Z(n67182) );
  NOR U81849 ( .A(n67184), .B(n67182), .Z(n61669) );
  IV U81850 ( .A(n61669), .Z(n62230) );
  IV U81851 ( .A(n61670), .Z(n61672) );
  NOR U81852 ( .A(n61672), .B(n61671), .Z(n67664) );
  NOR U81853 ( .A(n61673), .B(n67189), .Z(n61674) );
  NOR U81854 ( .A(n67664), .B(n61674), .Z(n62229) );
  IV U81855 ( .A(n61675), .Z(n61676) );
  NOR U81856 ( .A(n61679), .B(n61676), .Z(n67660) );
  IV U81857 ( .A(n61677), .Z(n61678) );
  NOR U81858 ( .A(n61679), .B(n61678), .Z(n67661) );
  NOR U81859 ( .A(n67660), .B(n67661), .Z(n62228) );
  IV U81860 ( .A(n61680), .Z(n61683) );
  IV U81861 ( .A(n61681), .Z(n61682) );
  NOR U81862 ( .A(n61683), .B(n61682), .Z(n67657) );
  IV U81863 ( .A(n62222), .Z(n77516) );
  IV U81864 ( .A(n61684), .Z(n61686) );
  NOR U81865 ( .A(n61686), .B(n61685), .Z(n61687) );
  IV U81866 ( .A(n61687), .Z(n62209) );
  IV U81867 ( .A(n61688), .Z(n61690) );
  NOR U81868 ( .A(n61690), .B(n61689), .Z(n67201) );
  IV U81869 ( .A(n61691), .Z(n61694) );
  NOR U81870 ( .A(n61692), .B(n62202), .Z(n61693) );
  IV U81871 ( .A(n61693), .Z(n62205) );
  NOR U81872 ( .A(n61694), .B(n62205), .Z(n67198) );
  IV U81873 ( .A(n61695), .Z(n62199) );
  IV U81874 ( .A(n61696), .Z(n61697) );
  NOR U81875 ( .A(n62199), .B(n61697), .Z(n67211) );
  IV U81876 ( .A(n61698), .Z(n61699) );
  NOR U81877 ( .A(n61699), .B(n62188), .Z(n67629) );
  NOR U81878 ( .A(n67211), .B(n67629), .Z(n62196) );
  IV U81879 ( .A(n61700), .Z(n61702) );
  NOR U81880 ( .A(n61702), .B(n61701), .Z(n61703) );
  IV U81881 ( .A(n61703), .Z(n62183) );
  IV U81882 ( .A(n61704), .Z(n61705) );
  NOR U81883 ( .A(n61705), .B(n61710), .Z(n67227) );
  IV U81884 ( .A(n61706), .Z(n61707) );
  NOR U81885 ( .A(n61708), .B(n61707), .Z(n67613) );
  IV U81886 ( .A(n61709), .Z(n61711) );
  NOR U81887 ( .A(n61711), .B(n61710), .Z(n67230) );
  NOR U81888 ( .A(n67613), .B(n67230), .Z(n62168) );
  IV U81889 ( .A(n61712), .Z(n61714) );
  NOR U81890 ( .A(n61714), .B(n61713), .Z(n67610) );
  IV U81891 ( .A(n61715), .Z(n61716) );
  NOR U81892 ( .A(n61717), .B(n61716), .Z(n72471) );
  IV U81893 ( .A(n61718), .Z(n61721) );
  IV U81894 ( .A(n61719), .Z(n61720) );
  NOR U81895 ( .A(n61721), .B(n61720), .Z(n72461) );
  NOR U81896 ( .A(n72471), .B(n72461), .Z(n67235) );
  IV U81897 ( .A(n61722), .Z(n61723) );
  NOR U81898 ( .A(n61723), .B(n61725), .Z(n67597) );
  IV U81899 ( .A(n61724), .Z(n61726) );
  NOR U81900 ( .A(n61726), .B(n61725), .Z(n62147) );
  IV U81901 ( .A(n62147), .Z(n62141) );
  IV U81902 ( .A(n61727), .Z(n61728) );
  NOR U81903 ( .A(n61730), .B(n61728), .Z(n67591) );
  IV U81904 ( .A(n61729), .Z(n61731) );
  NOR U81905 ( .A(n61731), .B(n61730), .Z(n61732) );
  IV U81906 ( .A(n61732), .Z(n67586) );
  IV U81907 ( .A(n61733), .Z(n61734) );
  NOR U81908 ( .A(n61734), .B(n62129), .Z(n67579) );
  NOR U81909 ( .A(n61735), .B(n67256), .Z(n61737) );
  NOR U81910 ( .A(n61737), .B(n61736), .Z(n61743) );
  IV U81911 ( .A(n61738), .Z(n61740) );
  NOR U81912 ( .A(n61740), .B(n61739), .Z(n67250) );
  NOR U81913 ( .A(n67250), .B(n67245), .Z(n61741) );
  IV U81914 ( .A(n61741), .Z(n61742) );
  NOR U81915 ( .A(n61743), .B(n61742), .Z(n61744) );
  IV U81916 ( .A(n61744), .Z(n62121) );
  NOR U81917 ( .A(n61745), .B(n67266), .Z(n61749) );
  IV U81918 ( .A(n61746), .Z(n67258) );
  IV U81919 ( .A(n61747), .Z(n61748) );
  NOR U81920 ( .A(n67258), .B(n61748), .Z(n67263) );
  NOR U81921 ( .A(n61749), .B(n67263), .Z(n62120) );
  IV U81922 ( .A(n61750), .Z(n61752) );
  NOR U81923 ( .A(n61752), .B(n61751), .Z(n67276) );
  NOR U81924 ( .A(n61754), .B(n61753), .Z(n67573) );
  NOR U81925 ( .A(n67276), .B(n67573), .Z(n62119) );
  IV U81926 ( .A(n61755), .Z(n61756) );
  NOR U81927 ( .A(n61756), .B(n62115), .Z(n67273) );
  IV U81928 ( .A(n61757), .Z(n61758) );
  NOR U81929 ( .A(n61759), .B(n61758), .Z(n72390) );
  IV U81930 ( .A(n61760), .Z(n61761) );
  NOR U81931 ( .A(n61761), .B(n62109), .Z(n72395) );
  NOR U81932 ( .A(n72390), .B(n72395), .Z(n67282) );
  IV U81933 ( .A(n61762), .Z(n62102) );
  IV U81934 ( .A(n61763), .Z(n61764) );
  NOR U81935 ( .A(n62102), .B(n61764), .Z(n61765) );
  IV U81936 ( .A(n61765), .Z(n67285) );
  XOR U81937 ( .A(n61767), .B(n61766), .Z(n61768) );
  NOR U81938 ( .A(n61769), .B(n61768), .Z(n61770) );
  IV U81939 ( .A(n61770), .Z(n62099) );
  NOR U81940 ( .A(n61771), .B(n67288), .Z(n62096) );
  IV U81941 ( .A(n61772), .Z(n61774) );
  NOR U81942 ( .A(n61774), .B(n61773), .Z(n67295) );
  IV U81943 ( .A(n61775), .Z(n61776) );
  NOR U81944 ( .A(n61782), .B(n61776), .Z(n67297) );
  NOR U81945 ( .A(n67295), .B(n67297), .Z(n62095) );
  IV U81946 ( .A(n61777), .Z(n61779) );
  IV U81947 ( .A(n61778), .Z(n67312) );
  NOR U81948 ( .A(n61779), .B(n67312), .Z(n67303) );
  IV U81949 ( .A(n61780), .Z(n61781) );
  NOR U81950 ( .A(n61782), .B(n61781), .Z(n67300) );
  NOR U81951 ( .A(n67303), .B(n67300), .Z(n62094) );
  IV U81952 ( .A(n61783), .Z(n61784) );
  NOR U81953 ( .A(n61784), .B(n67312), .Z(n62093) );
  NOR U81954 ( .A(n61785), .B(n62082), .Z(n62078) );
  IV U81955 ( .A(n61786), .Z(n61789) );
  NOR U81956 ( .A(n61787), .B(n61794), .Z(n61788) );
  IV U81957 ( .A(n61788), .Z(n62069) );
  NOR U81958 ( .A(n61789), .B(n62069), .Z(n67552) );
  IV U81959 ( .A(n61790), .Z(n61792) );
  IV U81960 ( .A(n61791), .Z(n61797) );
  NOR U81961 ( .A(n61792), .B(n61797), .Z(n67329) );
  IV U81962 ( .A(n61793), .Z(n61795) );
  NOR U81963 ( .A(n61795), .B(n61794), .Z(n67327) );
  NOR U81964 ( .A(n67329), .B(n67327), .Z(n62064) );
  IV U81965 ( .A(n61796), .Z(n61798) );
  NOR U81966 ( .A(n61798), .B(n61797), .Z(n62062) );
  IV U81967 ( .A(n62062), .Z(n62049) );
  IV U81968 ( .A(n62052), .Z(n61799) );
  NOR U81969 ( .A(n62056), .B(n61799), .Z(n67547) );
  IV U81970 ( .A(n61800), .Z(n61803) );
  NOR U81971 ( .A(n61801), .B(n62032), .Z(n61802) );
  IV U81972 ( .A(n61802), .Z(n62026) );
  NOR U81973 ( .A(n61803), .B(n62026), .Z(n67339) );
  NOR U81974 ( .A(n61804), .B(n67343), .Z(n62008) );
  IV U81975 ( .A(n61805), .Z(n61806) );
  NOR U81976 ( .A(n61807), .B(n61806), .Z(n67541) );
  IV U81977 ( .A(n61808), .Z(n61809) );
  NOR U81978 ( .A(n61809), .B(n61811), .Z(n67538) );
  IV U81979 ( .A(n61810), .Z(n61812) );
  NOR U81980 ( .A(n61812), .B(n61811), .Z(n61813) );
  IV U81981 ( .A(n61813), .Z(n67349) );
  IV U81982 ( .A(n61814), .Z(n67353) );
  NOR U81983 ( .A(n61815), .B(n67353), .Z(n61819) );
  IV U81984 ( .A(n61816), .Z(n61818) );
  NOR U81985 ( .A(n61818), .B(n61817), .Z(n67350) );
  NOR U81986 ( .A(n61819), .B(n67350), .Z(n62006) );
  IV U81987 ( .A(n61820), .Z(n61821) );
  NOR U81988 ( .A(n62000), .B(n61821), .Z(n72113) );
  IV U81989 ( .A(n61822), .Z(n61824) );
  IV U81990 ( .A(n61823), .Z(n62002) );
  NOR U81991 ( .A(n61824), .B(n62002), .Z(n72277) );
  NOR U81992 ( .A(n72113), .B(n72277), .Z(n67362) );
  IV U81993 ( .A(n61825), .Z(n61831) );
  IV U81994 ( .A(n61826), .Z(n61839) );
  XOR U81995 ( .A(n61827), .B(n61839), .Z(n61829) );
  NOR U81996 ( .A(n61829), .B(n61828), .Z(n61830) );
  IV U81997 ( .A(n61830), .Z(n61979) );
  NOR U81998 ( .A(n61831), .B(n61979), .Z(n67525) );
  IV U81999 ( .A(n61832), .Z(n61835) );
  NOR U82000 ( .A(n61839), .B(n61833), .Z(n61834) );
  IV U82001 ( .A(n61834), .Z(n61976) );
  NOR U82002 ( .A(n61835), .B(n61976), .Z(n61836) );
  IV U82003 ( .A(n61836), .Z(n67375) );
  IV U82004 ( .A(n61837), .Z(n61841) );
  NOR U82005 ( .A(n61839), .B(n61838), .Z(n61840) );
  IV U82006 ( .A(n61840), .Z(n61843) );
  NOR U82007 ( .A(n61841), .B(n61843), .Z(n67518) );
  IV U82008 ( .A(n61842), .Z(n61844) );
  NOR U82009 ( .A(n61844), .B(n61843), .Z(n67515) );
  IV U82010 ( .A(n61845), .Z(n61846) );
  NOR U82011 ( .A(n61846), .B(n61851), .Z(n67380) );
  NOR U82012 ( .A(n67515), .B(n67380), .Z(n61974) );
  IV U82013 ( .A(n61847), .Z(n61848) );
  NOR U82014 ( .A(n61849), .B(n61848), .Z(n67510) );
  IV U82015 ( .A(n61850), .Z(n61852) );
  NOR U82016 ( .A(n61852), .B(n61851), .Z(n67382) );
  NOR U82017 ( .A(n67510), .B(n67382), .Z(n61973) );
  IV U82018 ( .A(n61853), .Z(n61855) );
  NOR U82019 ( .A(n61855), .B(n61854), .Z(n67392) );
  IV U82020 ( .A(n61856), .Z(n61858) );
  NOR U82021 ( .A(n61858), .B(n61857), .Z(n67389) );
  NOR U82022 ( .A(n67392), .B(n67389), .Z(n61965) );
  IV U82023 ( .A(n61859), .Z(n61861) );
  IV U82024 ( .A(n61860), .Z(n61865) );
  NOR U82025 ( .A(n61861), .B(n61865), .Z(n67402) );
  IV U82026 ( .A(n61862), .Z(n61863) );
  NOR U82027 ( .A(n61863), .B(n61869), .Z(n67396) );
  IV U82028 ( .A(n61864), .Z(n61866) );
  NOR U82029 ( .A(n61866), .B(n61865), .Z(n67398) );
  NOR U82030 ( .A(n67396), .B(n67398), .Z(n61964) );
  IV U82031 ( .A(n61870), .Z(n61867) );
  NOR U82032 ( .A(n61867), .B(n61869), .Z(n67499) );
  IV U82033 ( .A(n61868), .Z(n61872) );
  XOR U82034 ( .A(n61870), .B(n61869), .Z(n61871) );
  NOR U82035 ( .A(n61872), .B(n61871), .Z(n67503) );
  NOR U82036 ( .A(n67499), .B(n67503), .Z(n61963) );
  IV U82037 ( .A(n61873), .Z(n61875) );
  NOR U82038 ( .A(n61875), .B(n61874), .Z(n67497) );
  IV U82039 ( .A(n61876), .Z(n61877) );
  NOR U82040 ( .A(n61960), .B(n61877), .Z(n67409) );
  IV U82041 ( .A(n61878), .Z(n61879) );
  NOR U82042 ( .A(n61884), .B(n61879), .Z(n67488) );
  IV U82043 ( .A(n61880), .Z(n61882) );
  NOR U82044 ( .A(n61882), .B(n61881), .Z(n67415) );
  IV U82045 ( .A(n61883), .Z(n61885) );
  NOR U82046 ( .A(n61885), .B(n61884), .Z(n67491) );
  NOR U82047 ( .A(n67415), .B(n67491), .Z(n61955) );
  IV U82048 ( .A(n61886), .Z(n61887) );
  NOR U82049 ( .A(n61888), .B(n61887), .Z(n72231) );
  IV U82050 ( .A(n61889), .Z(n61893) );
  IV U82051 ( .A(n61890), .Z(n61944) );
  NOR U82052 ( .A(n61891), .B(n61944), .Z(n61892) );
  IV U82053 ( .A(n61892), .Z(n61948) );
  NOR U82054 ( .A(n61893), .B(n61948), .Z(n72226) );
  NOR U82055 ( .A(n72231), .B(n72226), .Z(n67427) );
  IV U82056 ( .A(n61894), .Z(n61895) );
  NOR U82057 ( .A(n67440), .B(n61895), .Z(n61896) );
  IV U82058 ( .A(n61896), .Z(n67443) );
  IV U82059 ( .A(n61897), .Z(n61898) );
  NOR U82060 ( .A(n61906), .B(n61898), .Z(n67448) );
  IV U82061 ( .A(n61899), .Z(n61900) );
  NOR U82062 ( .A(n61900), .B(n61906), .Z(n61901) );
  IV U82063 ( .A(n61901), .Z(n67446) );
  IV U82064 ( .A(n61902), .Z(n61904) );
  NOR U82065 ( .A(n61904), .B(n61903), .Z(n67472) );
  IV U82066 ( .A(n61905), .Z(n61907) );
  NOR U82067 ( .A(n61907), .B(n61906), .Z(n67476) );
  NOR U82068 ( .A(n67472), .B(n67476), .Z(n61940) );
  IV U82069 ( .A(n61908), .Z(n61909) );
  NOR U82070 ( .A(n61909), .B(n61929), .Z(n67458) );
  IV U82071 ( .A(n61910), .Z(n61912) );
  NOR U82072 ( .A(n61912), .B(n61911), .Z(n61917) );
  IV U82073 ( .A(n61913), .Z(n61915) );
  NOR U82074 ( .A(n61915), .B(n61914), .Z(n61916) );
  NOR U82075 ( .A(n61917), .B(n61916), .Z(n67461) );
  IV U82076 ( .A(n67461), .Z(n61927) );
  NOR U82077 ( .A(n61919), .B(n61918), .Z(n67455) );
  XOR U82078 ( .A(n67454), .B(n67455), .Z(n61926) );
  IV U82079 ( .A(n61920), .Z(n61922) );
  NOR U82080 ( .A(n61922), .B(n61921), .Z(n61923) );
  IV U82081 ( .A(n61923), .Z(n61924) );
  NOR U82082 ( .A(n67455), .B(n61924), .Z(n61925) );
  NOR U82083 ( .A(n61926), .B(n61925), .Z(n67460) );
  XOR U82084 ( .A(n61927), .B(n67460), .Z(n67468) );
  XOR U82085 ( .A(n67458), .B(n67468), .Z(n67453) );
  IV U82086 ( .A(n67453), .Z(n61934) );
  IV U82087 ( .A(n61928), .Z(n61930) );
  NOR U82088 ( .A(n61930), .B(n61929), .Z(n67466) );
  IV U82089 ( .A(n61931), .Z(n61936) );
  IV U82090 ( .A(n61939), .Z(n61932) );
  NOR U82091 ( .A(n61936), .B(n61932), .Z(n67451) );
  NOR U82092 ( .A(n67466), .B(n67451), .Z(n61933) );
  XOR U82093 ( .A(n61934), .B(n61933), .Z(n67471) );
  NOR U82094 ( .A(n61936), .B(n61935), .Z(n61937) );
  IV U82095 ( .A(n61937), .Z(n61938) );
  NOR U82096 ( .A(n61939), .B(n61938), .Z(n67469) );
  XOR U82097 ( .A(n67471), .B(n67469), .Z(n67478) );
  XOR U82098 ( .A(n61940), .B(n67478), .Z(n67445) );
  XOR U82099 ( .A(n67446), .B(n67445), .Z(n67449) );
  XOR U82100 ( .A(n67448), .B(n67449), .Z(n67442) );
  XOR U82101 ( .A(n67443), .B(n67442), .Z(n67433) );
  NOR U82102 ( .A(n61942), .B(n61941), .Z(n67432) );
  IV U82103 ( .A(n61943), .Z(n61945) );
  NOR U82104 ( .A(n61945), .B(n61944), .Z(n67483) );
  NOR U82105 ( .A(n67432), .B(n67483), .Z(n61946) );
  XOR U82106 ( .A(n67433), .B(n61946), .Z(n67482) );
  IV U82107 ( .A(n61947), .Z(n61949) );
  NOR U82108 ( .A(n61949), .B(n61948), .Z(n67480) );
  XOR U82109 ( .A(n67482), .B(n67480), .Z(n72228) );
  XOR U82110 ( .A(n67427), .B(n72228), .Z(n67416) );
  NOR U82111 ( .A(n61950), .B(n67424), .Z(n67417) );
  IV U82112 ( .A(n61951), .Z(n61952) );
  NOR U82113 ( .A(n61953), .B(n61952), .Z(n67420) );
  NOR U82114 ( .A(n67417), .B(n67420), .Z(n61954) );
  XOR U82115 ( .A(n67416), .B(n61954), .Z(n67492) );
  XOR U82116 ( .A(n61955), .B(n67492), .Z(n67487) );
  XOR U82117 ( .A(n67488), .B(n67487), .Z(n67407) );
  IV U82118 ( .A(n61956), .Z(n61958) );
  NOR U82119 ( .A(n61958), .B(n61957), .Z(n67412) );
  IV U82120 ( .A(n61959), .Z(n61961) );
  NOR U82121 ( .A(n61961), .B(n61960), .Z(n67406) );
  NOR U82122 ( .A(n67412), .B(n67406), .Z(n61962) );
  XOR U82123 ( .A(n67407), .B(n61962), .Z(n67410) );
  XOR U82124 ( .A(n67409), .B(n67410), .Z(n67500) );
  XOR U82125 ( .A(n67497), .B(n67500), .Z(n67504) );
  XOR U82126 ( .A(n61963), .B(n67504), .Z(n67395) );
  XOR U82127 ( .A(n61964), .B(n67395), .Z(n67403) );
  XOR U82128 ( .A(n67402), .B(n67403), .Z(n67393) );
  XOR U82129 ( .A(n61965), .B(n67393), .Z(n67511) );
  IV U82130 ( .A(n61966), .Z(n61968) );
  NOR U82131 ( .A(n61968), .B(n61967), .Z(n67385) );
  IV U82132 ( .A(n61969), .Z(n61971) );
  NOR U82133 ( .A(n61971), .B(n61970), .Z(n67386) );
  NOR U82134 ( .A(n67385), .B(n67386), .Z(n61972) );
  XOR U82135 ( .A(n67511), .B(n61972), .Z(n67384) );
  XOR U82136 ( .A(n61973), .B(n67384), .Z(n67379) );
  XOR U82137 ( .A(n61974), .B(n67379), .Z(n67520) );
  XOR U82138 ( .A(n67518), .B(n67520), .Z(n67374) );
  XOR U82139 ( .A(n67375), .B(n67374), .Z(n67376) );
  IV U82140 ( .A(n61975), .Z(n61977) );
  NOR U82141 ( .A(n61977), .B(n61976), .Z(n67377) );
  IV U82142 ( .A(n61978), .Z(n61980) );
  NOR U82143 ( .A(n61980), .B(n61979), .Z(n67522) );
  NOR U82144 ( .A(n67377), .B(n67522), .Z(n61981) );
  XOR U82145 ( .A(n67376), .B(n61981), .Z(n67527) );
  XOR U82146 ( .A(n67525), .B(n67527), .Z(n67534) );
  IV U82147 ( .A(n61982), .Z(n61984) );
  IV U82148 ( .A(n61983), .Z(n61992) );
  NOR U82149 ( .A(n61984), .B(n61992), .Z(n67532) );
  IV U82150 ( .A(n61985), .Z(n61986) );
  NOR U82151 ( .A(n61987), .B(n61986), .Z(n67528) );
  NOR U82152 ( .A(n67532), .B(n67528), .Z(n61988) );
  XOR U82153 ( .A(n67534), .B(n61988), .Z(n67368) );
  IV U82154 ( .A(n61989), .Z(n61990) );
  NOR U82155 ( .A(n61997), .B(n61990), .Z(n67369) );
  IV U82156 ( .A(n61991), .Z(n61993) );
  NOR U82157 ( .A(n61993), .B(n61992), .Z(n67371) );
  NOR U82158 ( .A(n67369), .B(n67371), .Z(n61994) );
  XOR U82159 ( .A(n67368), .B(n61994), .Z(n67366) );
  IV U82160 ( .A(n61995), .Z(n61996) );
  NOR U82161 ( .A(n61997), .B(n61996), .Z(n67363) );
  XOR U82162 ( .A(n67366), .B(n67363), .Z(n72115) );
  XOR U82163 ( .A(n67362), .B(n72115), .Z(n62005) );
  IV U82164 ( .A(n61998), .Z(n61999) );
  NOR U82165 ( .A(n62000), .B(n61999), .Z(n67360) );
  IV U82166 ( .A(n62001), .Z(n62003) );
  NOR U82167 ( .A(n62003), .B(n62002), .Z(n67365) );
  NOR U82168 ( .A(n67360), .B(n67365), .Z(n62004) );
  XOR U82169 ( .A(n62005), .B(n62004), .Z(n67354) );
  XOR U82170 ( .A(n62006), .B(n67354), .Z(n67347) );
  XOR U82171 ( .A(n67349), .B(n67347), .Z(n67539) );
  XOR U82172 ( .A(n67538), .B(n67539), .Z(n67542) );
  XOR U82173 ( .A(n67541), .B(n67542), .Z(n62021) );
  IV U82174 ( .A(n62021), .Z(n62007) );
  NOR U82175 ( .A(n62008), .B(n62007), .Z(n62017) );
  IV U82176 ( .A(n62009), .Z(n62011) );
  NOR U82177 ( .A(n67343), .B(n67542), .Z(n62010) );
  IV U82178 ( .A(n62010), .Z(n62013) );
  NOR U82179 ( .A(n62011), .B(n62013), .Z(n72306) );
  IV U82180 ( .A(n62012), .Z(n62014) );
  NOR U82181 ( .A(n62014), .B(n62013), .Z(n72303) );
  NOR U82182 ( .A(n72306), .B(n72303), .Z(n62015) );
  IV U82183 ( .A(n62015), .Z(n62016) );
  NOR U82184 ( .A(n62017), .B(n62016), .Z(n62030) );
  IV U82185 ( .A(n62018), .Z(n67346) );
  NOR U82186 ( .A(n67346), .B(n62019), .Z(n62020) );
  NOR U82187 ( .A(n62030), .B(n62020), .Z(n62024) );
  IV U82188 ( .A(n62020), .Z(n62022) );
  NOR U82189 ( .A(n62022), .B(n62021), .Z(n62023) );
  NOR U82190 ( .A(n62024), .B(n62023), .Z(n62035) );
  IV U82191 ( .A(n62035), .Z(n62029) );
  IV U82192 ( .A(n62025), .Z(n62027) );
  NOR U82193 ( .A(n62027), .B(n62026), .Z(n62038) );
  IV U82194 ( .A(n62038), .Z(n62028) );
  NOR U82195 ( .A(n62029), .B(n62028), .Z(n72108) );
  IV U82196 ( .A(n62030), .Z(n67342) );
  IV U82197 ( .A(n62031), .Z(n62033) );
  NOR U82198 ( .A(n62033), .B(n62032), .Z(n62036) );
  IV U82199 ( .A(n62036), .Z(n62034) );
  NOR U82200 ( .A(n67342), .B(n62034), .Z(n72313) );
  NOR U82201 ( .A(n62036), .B(n62035), .Z(n62037) );
  NOR U82202 ( .A(n72313), .B(n62037), .Z(n67336) );
  NOR U82203 ( .A(n62038), .B(n67336), .Z(n62039) );
  NOR U82204 ( .A(n72108), .B(n62039), .Z(n62040) );
  IV U82205 ( .A(n62040), .Z(n67340) );
  XOR U82206 ( .A(n67339), .B(n67340), .Z(n67333) );
  IV U82207 ( .A(n62041), .Z(n62042) );
  NOR U82208 ( .A(n62043), .B(n62042), .Z(n67335) );
  IV U82209 ( .A(n62044), .Z(n62045) );
  NOR U82210 ( .A(n62046), .B(n62045), .Z(n67332) );
  NOR U82211 ( .A(n67335), .B(n67332), .Z(n62047) );
  XOR U82212 ( .A(n67333), .B(n62047), .Z(n62051) );
  XOR U82213 ( .A(n67547), .B(n62051), .Z(n62058) );
  IV U82214 ( .A(n62058), .Z(n62048) );
  NOR U82215 ( .A(n62049), .B(n62048), .Z(n72103) );
  IV U82216 ( .A(n62050), .Z(n62057) );
  IV U82217 ( .A(n62051), .Z(n67549) );
  XOR U82218 ( .A(n62052), .B(n62056), .Z(n62053) );
  NOR U82219 ( .A(n67549), .B(n62053), .Z(n62054) );
  IV U82220 ( .A(n62054), .Z(n62055) );
  NOR U82221 ( .A(n62057), .B(n62055), .Z(n72325) );
  NOR U82222 ( .A(n62057), .B(n62056), .Z(n62059) );
  NOR U82223 ( .A(n62059), .B(n62058), .Z(n62060) );
  NOR U82224 ( .A(n72325), .B(n62060), .Z(n62061) );
  NOR U82225 ( .A(n62062), .B(n62061), .Z(n62063) );
  NOR U82226 ( .A(n72103), .B(n62063), .Z(n67326) );
  XOR U82227 ( .A(n62064), .B(n67326), .Z(n67554) );
  XOR U82228 ( .A(n67552), .B(n67554), .Z(n67560) );
  IV U82229 ( .A(n62065), .Z(n62067) );
  NOR U82230 ( .A(n62067), .B(n62066), .Z(n67559) );
  IV U82231 ( .A(n62068), .Z(n62070) );
  NOR U82232 ( .A(n62070), .B(n62069), .Z(n67555) );
  NOR U82233 ( .A(n67559), .B(n67555), .Z(n62071) );
  XOR U82234 ( .A(n67560), .B(n62071), .Z(n62080) );
  NOR U82235 ( .A(n62072), .B(n67319), .Z(n62081) );
  IV U82236 ( .A(n62073), .Z(n62074) );
  NOR U82237 ( .A(n62075), .B(n62074), .Z(n67316) );
  NOR U82238 ( .A(n62081), .B(n67316), .Z(n62076) );
  XOR U82239 ( .A(n62080), .B(n62076), .Z(n67307) );
  IV U82240 ( .A(n67307), .Z(n62077) );
  NOR U82241 ( .A(n62078), .B(n62077), .Z(n62091) );
  IV U82242 ( .A(n62079), .Z(n62085) );
  IV U82243 ( .A(n62080), .Z(n67320) );
  XOR U82244 ( .A(n62081), .B(n67320), .Z(n62083) );
  NOR U82245 ( .A(n62083), .B(n62082), .Z(n62084) );
  IV U82246 ( .A(n62084), .Z(n62087) );
  NOR U82247 ( .A(n62085), .B(n62087), .Z(n72083) );
  IV U82248 ( .A(n62086), .Z(n62088) );
  NOR U82249 ( .A(n62088), .B(n62087), .Z(n72089) );
  NOR U82250 ( .A(n72083), .B(n72089), .Z(n62089) );
  IV U82251 ( .A(n62089), .Z(n62090) );
  NOR U82252 ( .A(n62091), .B(n62090), .Z(n62092) );
  IV U82253 ( .A(n62092), .Z(n67304) );
  XOR U82254 ( .A(n62093), .B(n67304), .Z(n67301) );
  XOR U82255 ( .A(n62094), .B(n67301), .Z(n67294) );
  XOR U82256 ( .A(n62095), .B(n67294), .Z(n67287) );
  XOR U82257 ( .A(n62096), .B(n67287), .Z(n62100) );
  NOR U82258 ( .A(n62100), .B(n62102), .Z(n62097) );
  IV U82259 ( .A(n62097), .Z(n62098) );
  NOR U82260 ( .A(n62099), .B(n62098), .Z(n72384) );
  IV U82261 ( .A(n62100), .Z(n62105) );
  IV U82262 ( .A(n62101), .Z(n62103) );
  NOR U82263 ( .A(n62103), .B(n62102), .Z(n62104) );
  NOR U82264 ( .A(n62105), .B(n62104), .Z(n62106) );
  NOR U82265 ( .A(n72384), .B(n62106), .Z(n67283) );
  XOR U82266 ( .A(n67285), .B(n67283), .Z(n72391) );
  XOR U82267 ( .A(n67282), .B(n72391), .Z(n62107) );
  IV U82268 ( .A(n62107), .Z(n67567) );
  IV U82269 ( .A(n62108), .Z(n62110) );
  NOR U82270 ( .A(n62110), .B(n62109), .Z(n67565) );
  XOR U82271 ( .A(n67567), .B(n67565), .Z(n67569) );
  IV U82272 ( .A(n67569), .Z(n62118) );
  IV U82273 ( .A(n62111), .Z(n62113) );
  NOR U82274 ( .A(n62113), .B(n62112), .Z(n67568) );
  IV U82275 ( .A(n62114), .Z(n62116) );
  NOR U82276 ( .A(n62116), .B(n62115), .Z(n67279) );
  NOR U82277 ( .A(n67568), .B(n67279), .Z(n62117) );
  XOR U82278 ( .A(n62118), .B(n62117), .Z(n67275) );
  XOR U82279 ( .A(n67273), .B(n67275), .Z(n67574) );
  XOR U82280 ( .A(n62119), .B(n67574), .Z(n67262) );
  XOR U82281 ( .A(n62120), .B(n67262), .Z(n67257) );
  XOR U82282 ( .A(n62121), .B(n67257), .Z(n67248) );
  IV U82283 ( .A(n62122), .Z(n62124) );
  NOR U82284 ( .A(n62124), .B(n62123), .Z(n67247) );
  XOR U82285 ( .A(n67248), .B(n67247), .Z(n67243) );
  IV U82286 ( .A(n62125), .Z(n62127) );
  NOR U82287 ( .A(n62127), .B(n62126), .Z(n67242) );
  IV U82288 ( .A(n62128), .Z(n62130) );
  NOR U82289 ( .A(n62130), .B(n62129), .Z(n67240) );
  NOR U82290 ( .A(n67242), .B(n67240), .Z(n62131) );
  XOR U82291 ( .A(n67243), .B(n62131), .Z(n62132) );
  IV U82292 ( .A(n62132), .Z(n67581) );
  XOR U82293 ( .A(n67579), .B(n67581), .Z(n67589) );
  IV U82294 ( .A(n62133), .Z(n62135) );
  NOR U82295 ( .A(n62135), .B(n62134), .Z(n67582) );
  IV U82296 ( .A(n62136), .Z(n62137) );
  NOR U82297 ( .A(n62138), .B(n62137), .Z(n67588) );
  NOR U82298 ( .A(n67582), .B(n67588), .Z(n62139) );
  XOR U82299 ( .A(n67589), .B(n62139), .Z(n67585) );
  XOR U82300 ( .A(n67586), .B(n67585), .Z(n67594) );
  XOR U82301 ( .A(n67591), .B(n67594), .Z(n62140) );
  NOR U82302 ( .A(n62141), .B(n62140), .Z(n72451) );
  IV U82303 ( .A(n62142), .Z(n62143) );
  NOR U82304 ( .A(n62144), .B(n62143), .Z(n67593) );
  NOR U82305 ( .A(n67591), .B(n67593), .Z(n62145) );
  XOR U82306 ( .A(n67594), .B(n62145), .Z(n62146) );
  NOR U82307 ( .A(n62147), .B(n62146), .Z(n62148) );
  NOR U82308 ( .A(n72451), .B(n62148), .Z(n62149) );
  IV U82309 ( .A(n62149), .Z(n67598) );
  XOR U82310 ( .A(n67597), .B(n67598), .Z(n67608) );
  IV U82311 ( .A(n62150), .Z(n62155) );
  IV U82312 ( .A(n62151), .Z(n62152) );
  NOR U82313 ( .A(n62153), .B(n62152), .Z(n62154) );
  IV U82314 ( .A(n62154), .Z(n62158) );
  NOR U82315 ( .A(n62155), .B(n62158), .Z(n67606) );
  NOR U82316 ( .A(n67601), .B(n67606), .Z(n62156) );
  XOR U82317 ( .A(n67608), .B(n62156), .Z(n67603) );
  IV U82318 ( .A(n62157), .Z(n62159) );
  NOR U82319 ( .A(n62159), .B(n62158), .Z(n62160) );
  IV U82320 ( .A(n62160), .Z(n67604) );
  XOR U82321 ( .A(n67603), .B(n67604), .Z(n72463) );
  XOR U82322 ( .A(n67235), .B(n72463), .Z(n67233) );
  IV U82323 ( .A(n62161), .Z(n62162) );
  NOR U82324 ( .A(n62163), .B(n62162), .Z(n67236) );
  IV U82325 ( .A(n62164), .Z(n62165) );
  NOR U82326 ( .A(n62166), .B(n62165), .Z(n67232) );
  NOR U82327 ( .A(n67236), .B(n67232), .Z(n62167) );
  XOR U82328 ( .A(n67233), .B(n62167), .Z(n67612) );
  XOR U82329 ( .A(n67610), .B(n67612), .Z(n67614) );
  XOR U82330 ( .A(n62168), .B(n67614), .Z(n62169) );
  IV U82331 ( .A(n62169), .Z(n67228) );
  XOR U82332 ( .A(n67227), .B(n67228), .Z(n67223) );
  IV U82333 ( .A(n62170), .Z(n62172) );
  NOR U82334 ( .A(n62172), .B(n62171), .Z(n67221) );
  XOR U82335 ( .A(n67223), .B(n67221), .Z(n67225) );
  IV U82336 ( .A(n62173), .Z(n62174) );
  NOR U82337 ( .A(n62175), .B(n62174), .Z(n67224) );
  IV U82338 ( .A(n62176), .Z(n62177) );
  NOR U82339 ( .A(n62177), .B(n62181), .Z(n67218) );
  NOR U82340 ( .A(n67224), .B(n67218), .Z(n62178) );
  XOR U82341 ( .A(n67225), .B(n62178), .Z(n62179) );
  IV U82342 ( .A(n62179), .Z(n67620) );
  IV U82343 ( .A(n62180), .Z(n62182) );
  NOR U82344 ( .A(n62182), .B(n62181), .Z(n67618) );
  XOR U82345 ( .A(n67620), .B(n67618), .Z(n67623) );
  NOR U82346 ( .A(n62183), .B(n67623), .Z(n72049) );
  IV U82347 ( .A(n62184), .Z(n62186) );
  NOR U82348 ( .A(n62186), .B(n62185), .Z(n67216) );
  IV U82349 ( .A(n62187), .Z(n62189) );
  NOR U82350 ( .A(n62189), .B(n62188), .Z(n67632) );
  IV U82351 ( .A(n62190), .Z(n62195) );
  IV U82352 ( .A(n62191), .Z(n62192) );
  NOR U82353 ( .A(n62195), .B(n62192), .Z(n67625) );
  IV U82354 ( .A(n62193), .Z(n62194) );
  NOR U82355 ( .A(n62195), .B(n62194), .Z(n67621) );
  XOR U82356 ( .A(n67623), .B(n67621), .Z(n67626) );
  XOR U82357 ( .A(n67625), .B(n67626), .Z(n67634) );
  XOR U82358 ( .A(n62196), .B(n67631), .Z(n67208) );
  IV U82359 ( .A(n62197), .Z(n62198) );
  NOR U82360 ( .A(n62199), .B(n62198), .Z(n67213) );
  IV U82361 ( .A(n62200), .Z(n62201) );
  NOR U82362 ( .A(n62202), .B(n62201), .Z(n67207) );
  NOR U82363 ( .A(n67213), .B(n67207), .Z(n62203) );
  XOR U82364 ( .A(n67208), .B(n62203), .Z(n67206) );
  IV U82365 ( .A(n62204), .Z(n62206) );
  NOR U82366 ( .A(n62206), .B(n62205), .Z(n67204) );
  XOR U82367 ( .A(n67206), .B(n67204), .Z(n67199) );
  XOR U82368 ( .A(n67198), .B(n67199), .Z(n67202) );
  XOR U82369 ( .A(n67201), .B(n67202), .Z(n67639) );
  NOR U82370 ( .A(n62209), .B(n67639), .Z(n77523) );
  IV U82371 ( .A(n62207), .Z(n62208) );
  NOR U82372 ( .A(n62219), .B(n62208), .Z(n67195) );
  XOR U82373 ( .A(n67638), .B(n67639), .Z(n67196) );
  IV U82374 ( .A(n67196), .Z(n62210) );
  XOR U82375 ( .A(n67195), .B(n62210), .Z(n62212) );
  NOR U82376 ( .A(n62210), .B(n62209), .Z(n62211) );
  NOR U82377 ( .A(n62212), .B(n62211), .Z(n62213) );
  NOR U82378 ( .A(n77523), .B(n62213), .Z(n62220) );
  IV U82379 ( .A(n62220), .Z(n67644) );
  NOR U82380 ( .A(n77516), .B(n67644), .Z(n72034) );
  IV U82381 ( .A(n62214), .Z(n62215) );
  NOR U82382 ( .A(n62216), .B(n62215), .Z(n67643) );
  IV U82383 ( .A(n62217), .Z(n62218) );
  NOR U82384 ( .A(n62219), .B(n62218), .Z(n67647) );
  NOR U82385 ( .A(n67643), .B(n67647), .Z(n67194) );
  XOR U82386 ( .A(n67194), .B(n62220), .Z(n77518) );
  IV U82387 ( .A(n77518), .Z(n62221) );
  NOR U82388 ( .A(n62222), .B(n62221), .Z(n62223) );
  NOR U82389 ( .A(n72034), .B(n62223), .Z(n67654) );
  IV U82390 ( .A(n62224), .Z(n62225) );
  NOR U82391 ( .A(n62226), .B(n62225), .Z(n62227) );
  IV U82392 ( .A(n62227), .Z(n67655) );
  XOR U82393 ( .A(n67654), .B(n67655), .Z(n78031) );
  XOR U82394 ( .A(n67657), .B(n78031), .Z(n67665) );
  XOR U82395 ( .A(n62228), .B(n67665), .Z(n67188) );
  XOR U82396 ( .A(n62229), .B(n67188), .Z(n67185) );
  XOR U82397 ( .A(n62230), .B(n67185), .Z(n67177) );
  XOR U82398 ( .A(n67175), .B(n67177), .Z(n67180) );
  IV U82399 ( .A(n62231), .Z(n62233) );
  NOR U82400 ( .A(n62233), .B(n62232), .Z(n67178) );
  XOR U82401 ( .A(n67180), .B(n67178), .Z(n67173) );
  IV U82402 ( .A(n62234), .Z(n62236) );
  NOR U82403 ( .A(n62236), .B(n62235), .Z(n67172) );
  IV U82404 ( .A(n62237), .Z(n62239) );
  NOR U82405 ( .A(n62239), .B(n62238), .Z(n67170) );
  NOR U82406 ( .A(n67172), .B(n67170), .Z(n62240) );
  XOR U82407 ( .A(n67173), .B(n62240), .Z(n67673) );
  XOR U82408 ( .A(n62241), .B(n67673), .Z(n67685) );
  XOR U82409 ( .A(n62242), .B(n67685), .Z(n67167) );
  XOR U82410 ( .A(n67168), .B(n67167), .Z(n67688) );
  XOR U82411 ( .A(n67687), .B(n67688), .Z(n67691) );
  XOR U82412 ( .A(n67690), .B(n67691), .Z(n67695) );
  XOR U82413 ( .A(n67694), .B(n67695), .Z(n67701) );
  IV U82414 ( .A(n62243), .Z(n62244) );
  NOR U82415 ( .A(n62245), .B(n62244), .Z(n67697) );
  NOR U82416 ( .A(n62247), .B(n62246), .Z(n67700) );
  NOR U82417 ( .A(n67697), .B(n67700), .Z(n62248) );
  XOR U82418 ( .A(n67701), .B(n62248), .Z(n62260) );
  IV U82419 ( .A(n62260), .Z(n67704) );
  IV U82420 ( .A(n62249), .Z(n62250) );
  NOR U82421 ( .A(n62254), .B(n62250), .Z(n62251) );
  IV U82422 ( .A(n62251), .Z(n62255) );
  NOR U82423 ( .A(n67704), .B(n62255), .Z(n71985) );
  IV U82424 ( .A(n62252), .Z(n62253) );
  NOR U82425 ( .A(n62254), .B(n62253), .Z(n67713) );
  NOR U82426 ( .A(n67713), .B(n62255), .Z(n62266) );
  IV U82427 ( .A(n62256), .Z(n62258) );
  IV U82428 ( .A(n62257), .Z(n62262) );
  NOR U82429 ( .A(n62258), .B(n62262), .Z(n62259) );
  IV U82430 ( .A(n62259), .Z(n67703) );
  XOR U82431 ( .A(n62260), .B(n67703), .Z(n67714) );
  IV U82432 ( .A(n62261), .Z(n62263) );
  NOR U82433 ( .A(n62263), .B(n62262), .Z(n67705) );
  NOR U82434 ( .A(n67713), .B(n67705), .Z(n62264) );
  XOR U82435 ( .A(n67714), .B(n62264), .Z(n62265) );
  NOR U82436 ( .A(n62266), .B(n62265), .Z(n62267) );
  NOR U82437 ( .A(n71985), .B(n62267), .Z(n67165) );
  XOR U82438 ( .A(n62268), .B(n67165), .Z(n67163) );
  XOR U82439 ( .A(n67161), .B(n67163), .Z(n71976) );
  XOR U82440 ( .A(n67722), .B(n71976), .Z(n62279) );
  IV U82441 ( .A(n62279), .Z(n67723) );
  IV U82442 ( .A(n62269), .Z(n62270) );
  NOR U82443 ( .A(n62271), .B(n62270), .Z(n62278) );
  IV U82444 ( .A(n62272), .Z(n62273) );
  NOR U82445 ( .A(n62274), .B(n62273), .Z(n67159) );
  NOR U82446 ( .A(n62278), .B(n67159), .Z(n62275) );
  XOR U82447 ( .A(n67723), .B(n62275), .Z(n62276) );
  NOR U82448 ( .A(n62277), .B(n62276), .Z(n62282) );
  IV U82449 ( .A(n62277), .Z(n62281) );
  IV U82450 ( .A(n62278), .Z(n67724) );
  XOR U82451 ( .A(n67724), .B(n62279), .Z(n62280) );
  NOR U82452 ( .A(n62281), .B(n62280), .Z(n71970) );
  NOR U82453 ( .A(n62282), .B(n71970), .Z(n67156) );
  XOR U82454 ( .A(n67158), .B(n67156), .Z(n67729) );
  XOR U82455 ( .A(n62283), .B(n67729), .Z(n67733) );
  IV U82456 ( .A(n62284), .Z(n62285) );
  NOR U82457 ( .A(n62285), .B(n62287), .Z(n67731) );
  XOR U82458 ( .A(n67733), .B(n67731), .Z(n67737) );
  IV U82459 ( .A(n62286), .Z(n62288) );
  NOR U82460 ( .A(n62288), .B(n62287), .Z(n67735) );
  XOR U82461 ( .A(n67737), .B(n67735), .Z(n67739) );
  XOR U82462 ( .A(n67738), .B(n67739), .Z(n67743) );
  IV U82463 ( .A(n62289), .Z(n62290) );
  NOR U82464 ( .A(n62291), .B(n62290), .Z(n67152) );
  IV U82465 ( .A(n62292), .Z(n62294) );
  NOR U82466 ( .A(n62294), .B(n62293), .Z(n67742) );
  NOR U82467 ( .A(n67152), .B(n67742), .Z(n62295) );
  XOR U82468 ( .A(n67743), .B(n62295), .Z(n67148) );
  IV U82469 ( .A(n62296), .Z(n62298) );
  NOR U82470 ( .A(n62298), .B(n62297), .Z(n62299) );
  IV U82471 ( .A(n62299), .Z(n67149) );
  XOR U82472 ( .A(n67148), .B(n67149), .Z(n67746) );
  XOR U82473 ( .A(n67745), .B(n67746), .Z(n67750) );
  XOR U82474 ( .A(n62300), .B(n67750), .Z(n62301) );
  IV U82475 ( .A(n62301), .Z(n67144) );
  XOR U82476 ( .A(n67143), .B(n67144), .Z(n67128) );
  NOR U82477 ( .A(n62302), .B(n67137), .Z(n62306) );
  IV U82478 ( .A(n62303), .Z(n67129) );
  NOR U82479 ( .A(n62304), .B(n67129), .Z(n62305) );
  NOR U82480 ( .A(n62306), .B(n62305), .Z(n62307) );
  XOR U82481 ( .A(n67128), .B(n62307), .Z(n62308) );
  IV U82482 ( .A(n62308), .Z(n67126) );
  IV U82483 ( .A(n62309), .Z(n62311) );
  NOR U82484 ( .A(n62311), .B(n62310), .Z(n67124) );
  NOR U82485 ( .A(n62313), .B(n62312), .Z(n62314) );
  IV U82486 ( .A(n62314), .Z(n62320) );
  IV U82487 ( .A(n62315), .Z(n62316) );
  NOR U82488 ( .A(n62317), .B(n62316), .Z(n62318) );
  IV U82489 ( .A(n62318), .Z(n62319) );
  NOR U82490 ( .A(n62320), .B(n62319), .Z(n62321) );
  IV U82491 ( .A(n62321), .Z(n62322) );
  NOR U82492 ( .A(n62323), .B(n62322), .Z(n67122) );
  NOR U82493 ( .A(n67124), .B(n67122), .Z(n62324) );
  XOR U82494 ( .A(n67126), .B(n62324), .Z(n62325) );
  NOR U82495 ( .A(n62326), .B(n62325), .Z(n62329) );
  IV U82496 ( .A(n62326), .Z(n62328) );
  XOR U82497 ( .A(n67124), .B(n67126), .Z(n62327) );
  NOR U82498 ( .A(n62328), .B(n62327), .Z(n72637) );
  NOR U82499 ( .A(n62329), .B(n72637), .Z(n67754) );
  XOR U82500 ( .A(n62330), .B(n67754), .Z(n67760) );
  XOR U82501 ( .A(n62331), .B(n67760), .Z(n67118) );
  XOR U82502 ( .A(n67116), .B(n67118), .Z(n67120) );
  IV U82503 ( .A(n62332), .Z(n62334) );
  NOR U82504 ( .A(n62334), .B(n62333), .Z(n67119) );
  IV U82505 ( .A(n62335), .Z(n62336) );
  NOR U82506 ( .A(n62337), .B(n62336), .Z(n67114) );
  NOR U82507 ( .A(n67119), .B(n67114), .Z(n62338) );
  XOR U82508 ( .A(n67120), .B(n62338), .Z(n67774) );
  XOR U82509 ( .A(n67775), .B(n67774), .Z(n67112) );
  IV U82510 ( .A(n62339), .Z(n62340) );
  NOR U82511 ( .A(n62342), .B(n62340), .Z(n67110) );
  XOR U82512 ( .A(n67112), .B(n67110), .Z(n67773) );
  IV U82513 ( .A(n62341), .Z(n62343) );
  NOR U82514 ( .A(n62343), .B(n62342), .Z(n67771) );
  XOR U82515 ( .A(n67773), .B(n67771), .Z(n67108) );
  XOR U82516 ( .A(n67107), .B(n67108), .Z(n67796) );
  IV U82517 ( .A(n62344), .Z(n62345) );
  NOR U82518 ( .A(n62346), .B(n62345), .Z(n67794) );
  XOR U82519 ( .A(n67796), .B(n67794), .Z(n62357) );
  IV U82520 ( .A(n62357), .Z(n62355) );
  IV U82521 ( .A(n62347), .Z(n62348) );
  NOR U82522 ( .A(n62349), .B(n62348), .Z(n62359) );
  IV U82523 ( .A(n62350), .Z(n62351) );
  NOR U82524 ( .A(n62352), .B(n62351), .Z(n62356) );
  NOR U82525 ( .A(n62359), .B(n62356), .Z(n62353) );
  IV U82526 ( .A(n62353), .Z(n62354) );
  NOR U82527 ( .A(n62355), .B(n62354), .Z(n62362) );
  IV U82528 ( .A(n62356), .Z(n62358) );
  NOR U82529 ( .A(n62358), .B(n62357), .Z(n71929) );
  IV U82530 ( .A(n62359), .Z(n62360) );
  NOR U82531 ( .A(n62360), .B(n67796), .Z(n71927) );
  NOR U82532 ( .A(n71929), .B(n71927), .Z(n62361) );
  IV U82533 ( .A(n62361), .Z(n67797) );
  NOR U82534 ( .A(n62362), .B(n67797), .Z(n62363) );
  IV U82535 ( .A(n62363), .Z(n67104) );
  XOR U82536 ( .A(n67103), .B(n67104), .Z(n62364) );
  NOR U82537 ( .A(n62365), .B(n62364), .Z(n72663) );
  IV U82538 ( .A(n62366), .Z(n62367) );
  NOR U82539 ( .A(n62368), .B(n62367), .Z(n67101) );
  NOR U82540 ( .A(n67103), .B(n67101), .Z(n62369) );
  XOR U82541 ( .A(n67104), .B(n62369), .Z(n62370) );
  NOR U82542 ( .A(n62371), .B(n62370), .Z(n62372) );
  NOR U82543 ( .A(n72663), .B(n62372), .Z(n62373) );
  IV U82544 ( .A(n62373), .Z(n67100) );
  IV U82545 ( .A(n62374), .Z(n62376) );
  NOR U82546 ( .A(n62376), .B(n62375), .Z(n67098) );
  XOR U82547 ( .A(n67100), .B(n67098), .Z(n67097) );
  XOR U82548 ( .A(n62377), .B(n67097), .Z(n67801) );
  IV U82549 ( .A(n62378), .Z(n62379) );
  NOR U82550 ( .A(n62380), .B(n62379), .Z(n62381) );
  NOR U82551 ( .A(n78166), .B(n62381), .Z(n67802) );
  XOR U82552 ( .A(n67801), .B(n67802), .Z(n67805) );
  XOR U82553 ( .A(n67803), .B(n67805), .Z(n67088) );
  XOR U82554 ( .A(n67087), .B(n67088), .Z(n67091) );
  XOR U82555 ( .A(n67090), .B(n67091), .Z(n67809) );
  XOR U82556 ( .A(n67808), .B(n67809), .Z(n67813) );
  XOR U82557 ( .A(n62382), .B(n67813), .Z(n62383) );
  IV U82558 ( .A(n62383), .Z(n67816) );
  XOR U82559 ( .A(n67815), .B(n67816), .Z(n67820) );
  IV U82560 ( .A(n62384), .Z(n62385) );
  NOR U82561 ( .A(n62385), .B(n62387), .Z(n67818) );
  XOR U82562 ( .A(n67820), .B(n67818), .Z(n67824) );
  IV U82563 ( .A(n62386), .Z(n62388) );
  NOR U82564 ( .A(n62388), .B(n62387), .Z(n67822) );
  XOR U82565 ( .A(n67824), .B(n67822), .Z(n67834) );
  IV U82566 ( .A(n67834), .Z(n62395) );
  IV U82567 ( .A(n62389), .Z(n62390) );
  NOR U82568 ( .A(n67829), .B(n62390), .Z(n67825) );
  IV U82569 ( .A(n62391), .Z(n62393) );
  NOR U82570 ( .A(n62393), .B(n62392), .Z(n67833) );
  NOR U82571 ( .A(n67825), .B(n67833), .Z(n62394) );
  XOR U82572 ( .A(n62395), .B(n62394), .Z(n67828) );
  XOR U82573 ( .A(n67079), .B(n67828), .Z(n67074) );
  XOR U82574 ( .A(n62396), .B(n67074), .Z(n67063) );
  XOR U82575 ( .A(n62397), .B(n67063), .Z(n67840) );
  XOR U82576 ( .A(n67839), .B(n67840), .Z(n67847) );
  XOR U82577 ( .A(n62398), .B(n67847), .Z(n67849) );
  IV U82578 ( .A(n62399), .Z(n67850) );
  NOR U82579 ( .A(n62400), .B(n67850), .Z(n62408) );
  IV U82580 ( .A(n62401), .Z(n62402) );
  NOR U82581 ( .A(n62402), .B(n62404), .Z(n67860) );
  IV U82582 ( .A(n62403), .Z(n62405) );
  NOR U82583 ( .A(n62405), .B(n62404), .Z(n67854) );
  NOR U82584 ( .A(n67860), .B(n67854), .Z(n62406) );
  IV U82585 ( .A(n62406), .Z(n62407) );
  NOR U82586 ( .A(n62408), .B(n62407), .Z(n62409) );
  XOR U82587 ( .A(n67849), .B(n62409), .Z(n67867) );
  IV U82588 ( .A(n62410), .Z(n62411) );
  NOR U82589 ( .A(n62412), .B(n62411), .Z(n67863) );
  IV U82590 ( .A(n62413), .Z(n62414) );
  NOR U82591 ( .A(n62414), .B(n62420), .Z(n67865) );
  NOR U82592 ( .A(n67863), .B(n67865), .Z(n62415) );
  XOR U82593 ( .A(n67867), .B(n62415), .Z(n67869) );
  IV U82594 ( .A(n62416), .Z(n62417) );
  NOR U82595 ( .A(n62425), .B(n62417), .Z(n67868) );
  IV U82596 ( .A(n62418), .Z(n62419) );
  NOR U82597 ( .A(n62420), .B(n62419), .Z(n67061) );
  NOR U82598 ( .A(n67868), .B(n67061), .Z(n62421) );
  XOR U82599 ( .A(n67869), .B(n62421), .Z(n78221) );
  XOR U82600 ( .A(n78206), .B(n78221), .Z(n62430) );
  NOR U82601 ( .A(n62422), .B(n67873), .Z(n62428) );
  IV U82602 ( .A(n62423), .Z(n62424) );
  NOR U82603 ( .A(n62425), .B(n62424), .Z(n62426) );
  IV U82604 ( .A(n62426), .Z(n67060) );
  NOR U82605 ( .A(n62427), .B(n67060), .Z(n78219) );
  NOR U82606 ( .A(n62428), .B(n78219), .Z(n62429) );
  XOR U82607 ( .A(n62430), .B(n62429), .Z(n67881) );
  XOR U82608 ( .A(n62431), .B(n67881), .Z(n62436) );
  IV U82609 ( .A(n62436), .Z(n67888) );
  NOR U82610 ( .A(n62440), .B(n67888), .Z(n72752) );
  IV U82611 ( .A(n62432), .Z(n62434) );
  IV U82612 ( .A(n62433), .Z(n62438) );
  NOR U82613 ( .A(n62434), .B(n62438), .Z(n62435) );
  IV U82614 ( .A(n62435), .Z(n67887) );
  XOR U82615 ( .A(n62436), .B(n67887), .Z(n67890) );
  IV U82616 ( .A(n62437), .Z(n62439) );
  NOR U82617 ( .A(n62439), .B(n62438), .Z(n62441) );
  IV U82618 ( .A(n62441), .Z(n67889) );
  XOR U82619 ( .A(n67890), .B(n67889), .Z(n62443) );
  NOR U82620 ( .A(n62441), .B(n62440), .Z(n62442) );
  NOR U82621 ( .A(n62443), .B(n62442), .Z(n62444) );
  NOR U82622 ( .A(n72752), .B(n62444), .Z(n62445) );
  IV U82623 ( .A(n62445), .Z(n67054) );
  IV U82624 ( .A(n62446), .Z(n62447) );
  NOR U82625 ( .A(n62448), .B(n62447), .Z(n67052) );
  XOR U82626 ( .A(n67054), .B(n67052), .Z(n67057) );
  XOR U82627 ( .A(n67055), .B(n67057), .Z(n67897) );
  XOR U82628 ( .A(n62449), .B(n67897), .Z(n62450) );
  IV U82629 ( .A(n62450), .Z(n67048) );
  XOR U82630 ( .A(n67046), .B(n67048), .Z(n67040) );
  XOR U82631 ( .A(n67039), .B(n67040), .Z(n67043) );
  XOR U82632 ( .A(n67042), .B(n67043), .Z(n71854) );
  XOR U82633 ( .A(n67038), .B(n71854), .Z(n67032) );
  XOR U82634 ( .A(n67033), .B(n67032), .Z(n67036) );
  XOR U82635 ( .A(n67035), .B(n67036), .Z(n67906) );
  XOR U82636 ( .A(n67907), .B(n67906), .Z(n62457) );
  IV U82637 ( .A(n62457), .Z(n62451) );
  NOR U82638 ( .A(n62455), .B(n62451), .Z(n62452) );
  IV U82639 ( .A(n62452), .Z(n62453) );
  NOR U82640 ( .A(n62454), .B(n62453), .Z(n67031) );
  NOR U82641 ( .A(n62465), .B(n62455), .Z(n62456) );
  NOR U82642 ( .A(n62457), .B(n62456), .Z(n62458) );
  NOR U82643 ( .A(n67031), .B(n62458), .Z(n62459) );
  IV U82644 ( .A(n62459), .Z(n67904) );
  XOR U82645 ( .A(n67903), .B(n67904), .Z(n67029) );
  IV U82646 ( .A(n67029), .Z(n62467) );
  IV U82647 ( .A(n62460), .Z(n62461) );
  NOR U82648 ( .A(n62462), .B(n62461), .Z(n67026) );
  IV U82649 ( .A(n62463), .Z(n62464) );
  NOR U82650 ( .A(n62465), .B(n62464), .Z(n67028) );
  NOR U82651 ( .A(n67026), .B(n67028), .Z(n62466) );
  XOR U82652 ( .A(n62467), .B(n62466), .Z(n67021) );
  XOR U82653 ( .A(n67020), .B(n67021), .Z(n67025) );
  XOR U82654 ( .A(n67023), .B(n67025), .Z(n67015) );
  XOR U82655 ( .A(n62468), .B(n67015), .Z(n67004) );
  XOR U82656 ( .A(n67006), .B(n67004), .Z(n67923) );
  IV U82657 ( .A(n67923), .Z(n62476) );
  IV U82658 ( .A(n62469), .Z(n62471) );
  NOR U82659 ( .A(n62471), .B(n62470), .Z(n67918) );
  IV U82660 ( .A(n62472), .Z(n62474) );
  NOR U82661 ( .A(n62474), .B(n62473), .Z(n67922) );
  NOR U82662 ( .A(n67918), .B(n67922), .Z(n62475) );
  XOR U82663 ( .A(n62476), .B(n62475), .Z(n67929) );
  XOR U82664 ( .A(n67920), .B(n67929), .Z(n62477) );
  XOR U82665 ( .A(n62478), .B(n62477), .Z(n67933) );
  XOR U82666 ( .A(n66998), .B(n67933), .Z(n62493) );
  XOR U82667 ( .A(n62479), .B(n62493), .Z(n62490) );
  IV U82668 ( .A(n62490), .Z(n62488) );
  IV U82669 ( .A(n62480), .Z(n62482) );
  NOR U82670 ( .A(n62482), .B(n62481), .Z(n62492) );
  IV U82671 ( .A(n62483), .Z(n62484) );
  NOR U82672 ( .A(n62485), .B(n62484), .Z(n62489) );
  NOR U82673 ( .A(n62492), .B(n62489), .Z(n62486) );
  IV U82674 ( .A(n62486), .Z(n62487) );
  NOR U82675 ( .A(n62488), .B(n62487), .Z(n62496) );
  IV U82676 ( .A(n62489), .Z(n62491) );
  NOR U82677 ( .A(n62491), .B(n62490), .Z(n72840) );
  IV U82678 ( .A(n62492), .Z(n62494) );
  NOR U82679 ( .A(n62494), .B(n62493), .Z(n72838) );
  NOR U82680 ( .A(n72840), .B(n72838), .Z(n62495) );
  IV U82681 ( .A(n62495), .Z(n67947) );
  NOR U82682 ( .A(n62496), .B(n67947), .Z(n62497) );
  IV U82683 ( .A(n62497), .Z(n67943) );
  XOR U82684 ( .A(n67940), .B(n67943), .Z(n62498) );
  NOR U82685 ( .A(n62499), .B(n62498), .Z(n72842) );
  IV U82686 ( .A(n62500), .Z(n62502) );
  NOR U82687 ( .A(n62502), .B(n62501), .Z(n67942) );
  NOR U82688 ( .A(n67940), .B(n67942), .Z(n62503) );
  XOR U82689 ( .A(n62503), .B(n67943), .Z(n62504) );
  NOR U82690 ( .A(n62505), .B(n62504), .Z(n62506) );
  NOR U82691 ( .A(n72842), .B(n62506), .Z(n66988) );
  IV U82692 ( .A(n62507), .Z(n62508) );
  NOR U82693 ( .A(n62509), .B(n62508), .Z(n66992) );
  NOR U82694 ( .A(n62510), .B(n66989), .Z(n62511) );
  NOR U82695 ( .A(n66992), .B(n62511), .Z(n62512) );
  XOR U82696 ( .A(n66988), .B(n62512), .Z(n66986) );
  XOR U82697 ( .A(n66984), .B(n66986), .Z(n66982) );
  NOR U82698 ( .A(n62519), .B(n66982), .Z(n77291) );
  IV U82699 ( .A(n62513), .Z(n62515) );
  NOR U82700 ( .A(n62515), .B(n62514), .Z(n66981) );
  XOR U82701 ( .A(n66981), .B(n66982), .Z(n66980) );
  IV U82702 ( .A(n62516), .Z(n62518) );
  NOR U82703 ( .A(n62518), .B(n62517), .Z(n62520) );
  IV U82704 ( .A(n62520), .Z(n66979) );
  XOR U82705 ( .A(n66980), .B(n66979), .Z(n62522) );
  NOR U82706 ( .A(n62520), .B(n62519), .Z(n62521) );
  NOR U82707 ( .A(n62522), .B(n62521), .Z(n62523) );
  NOR U82708 ( .A(n77291), .B(n62523), .Z(n67954) );
  XOR U82709 ( .A(n62524), .B(n67954), .Z(n67963) );
  XOR U82710 ( .A(n62525), .B(n67963), .Z(n62526) );
  IV U82711 ( .A(n62526), .Z(n67965) );
  XOR U82712 ( .A(n67964), .B(n67965), .Z(n67983) );
  XOR U82713 ( .A(n62527), .B(n67983), .Z(n67979) );
  XOR U82714 ( .A(n62528), .B(n67979), .Z(n67991) );
  IV U82715 ( .A(n62529), .Z(n62530) );
  NOR U82716 ( .A(n62531), .B(n62530), .Z(n67989) );
  XOR U82717 ( .A(n67991), .B(n67989), .Z(n67995) );
  IV U82718 ( .A(n67995), .Z(n62539) );
  NOR U82719 ( .A(n62532), .B(n67996), .Z(n62543) );
  IV U82720 ( .A(n62543), .Z(n62533) );
  NOR U82721 ( .A(n62539), .B(n62533), .Z(n62545) );
  IV U82722 ( .A(n62534), .Z(n62535) );
  NOR U82723 ( .A(n62536), .B(n62535), .Z(n62538) );
  IV U82724 ( .A(n62538), .Z(n62537) );
  NOR U82725 ( .A(n62537), .B(n67991), .Z(n71818) );
  NOR U82726 ( .A(n62539), .B(n62538), .Z(n62540) );
  NOR U82727 ( .A(n71818), .B(n62540), .Z(n62541) );
  IV U82728 ( .A(n62541), .Z(n62542) );
  NOR U82729 ( .A(n62543), .B(n62542), .Z(n62544) );
  NOR U82730 ( .A(n62545), .B(n62544), .Z(n68000) );
  IV U82731 ( .A(n62546), .Z(n62547) );
  NOR U82732 ( .A(n62548), .B(n62547), .Z(n67999) );
  NOR U82733 ( .A(n62549), .B(n66976), .Z(n62550) );
  NOR U82734 ( .A(n67999), .B(n62550), .Z(n62551) );
  XOR U82735 ( .A(n68000), .B(n62551), .Z(n66961) );
  IV U82736 ( .A(n62552), .Z(n62553) );
  NOR U82737 ( .A(n62553), .B(n66969), .Z(n62554) );
  IV U82738 ( .A(n62554), .Z(n66962) );
  XOR U82739 ( .A(n66961), .B(n66962), .Z(n66965) );
  XOR U82740 ( .A(n62555), .B(n66965), .Z(n68013) );
  XOR U82741 ( .A(n62556), .B(n68013), .Z(n68024) );
  XOR U82742 ( .A(n68025), .B(n68024), .Z(n62557) );
  NOR U82743 ( .A(n62558), .B(n62557), .Z(n62560) );
  IV U82744 ( .A(n62558), .Z(n62559) );
  XOR U82745 ( .A(n68011), .B(n68013), .Z(n68019) );
  NOR U82746 ( .A(n62559), .B(n68019), .Z(n66960) );
  NOR U82747 ( .A(n62560), .B(n66960), .Z(n62561) );
  IV U82748 ( .A(n62561), .Z(n68023) );
  IV U82749 ( .A(n62562), .Z(n62563) );
  NOR U82750 ( .A(n62564), .B(n62563), .Z(n66957) );
  IV U82751 ( .A(n62565), .Z(n62567) );
  NOR U82752 ( .A(n62567), .B(n62566), .Z(n68021) );
  NOR U82753 ( .A(n66957), .B(n68021), .Z(n62568) );
  XOR U82754 ( .A(n68023), .B(n62568), .Z(n62569) );
  NOR U82755 ( .A(n62570), .B(n62569), .Z(n62573) );
  IV U82756 ( .A(n62570), .Z(n62572) );
  XOR U82757 ( .A(n68021), .B(n68023), .Z(n62571) );
  NOR U82758 ( .A(n62572), .B(n62571), .Z(n71787) );
  NOR U82759 ( .A(n62573), .B(n71787), .Z(n68034) );
  IV U82760 ( .A(n62574), .Z(n62575) );
  NOR U82761 ( .A(n62576), .B(n62575), .Z(n68033) );
  IV U82762 ( .A(n62577), .Z(n62578) );
  NOR U82763 ( .A(n62579), .B(n62578), .Z(n68037) );
  NOR U82764 ( .A(n68033), .B(n68037), .Z(n62580) );
  XOR U82765 ( .A(n68034), .B(n62580), .Z(n66953) );
  IV U82766 ( .A(n62581), .Z(n62582) );
  NOR U82767 ( .A(n62583), .B(n62582), .Z(n62587) );
  IV U82768 ( .A(n62587), .Z(n62584) );
  NOR U82769 ( .A(n66953), .B(n62584), .Z(n72910) );
  NOR U82770 ( .A(n66955), .B(n66952), .Z(n62585) );
  XOR U82771 ( .A(n66953), .B(n62585), .Z(n62595) );
  IV U82772 ( .A(n62595), .Z(n62586) );
  NOR U82773 ( .A(n62587), .B(n62586), .Z(n62588) );
  NOR U82774 ( .A(n72910), .B(n62588), .Z(n68042) );
  IV U82775 ( .A(n62589), .Z(n62591) );
  NOR U82776 ( .A(n62591), .B(n62590), .Z(n62601) );
  IV U82777 ( .A(n62601), .Z(n68044) );
  NOR U82778 ( .A(n68042), .B(n68044), .Z(n62603) );
  IV U82779 ( .A(n62592), .Z(n62594) );
  NOR U82780 ( .A(n62594), .B(n62593), .Z(n62597) );
  IV U82781 ( .A(n62597), .Z(n62596) );
  NOR U82782 ( .A(n62596), .B(n62595), .Z(n71772) );
  NOR U82783 ( .A(n68042), .B(n62597), .Z(n62598) );
  NOR U82784 ( .A(n71772), .B(n62598), .Z(n62599) );
  IV U82785 ( .A(n62599), .Z(n62600) );
  NOR U82786 ( .A(n62601), .B(n62600), .Z(n62602) );
  NOR U82787 ( .A(n62603), .B(n62602), .Z(n68058) );
  XOR U82788 ( .A(n62604), .B(n68058), .Z(n66945) );
  NOR U82789 ( .A(n62606), .B(n62605), .Z(n66949) );
  IV U82790 ( .A(n62607), .Z(n62609) );
  NOR U82791 ( .A(n62609), .B(n62608), .Z(n66946) );
  NOR U82792 ( .A(n66949), .B(n66946), .Z(n62610) );
  XOR U82793 ( .A(n66945), .B(n62610), .Z(n66941) );
  IV U82794 ( .A(n62611), .Z(n62613) );
  NOR U82795 ( .A(n62613), .B(n62612), .Z(n66939) );
  XOR U82796 ( .A(n66941), .B(n66939), .Z(n66944) );
  XOR U82797 ( .A(n66942), .B(n66944), .Z(n68063) );
  XOR U82798 ( .A(n62614), .B(n68063), .Z(n66934) );
  XOR U82799 ( .A(n62615), .B(n66934), .Z(n68080) );
  IV U82800 ( .A(n68080), .Z(n62623) );
  IV U82801 ( .A(n62616), .Z(n62617) );
  NOR U82802 ( .A(n62618), .B(n62617), .Z(n66931) );
  IV U82803 ( .A(n62619), .Z(n62621) );
  NOR U82804 ( .A(n62621), .B(n62620), .Z(n68078) );
  NOR U82805 ( .A(n66931), .B(n68078), .Z(n62622) );
  XOR U82806 ( .A(n62623), .B(n62622), .Z(n66926) );
  XOR U82807 ( .A(n66925), .B(n66926), .Z(n66929) );
  IV U82808 ( .A(n62624), .Z(n62625) );
  NOR U82809 ( .A(n62626), .B(n62625), .Z(n66928) );
  NOR U82810 ( .A(n62627), .B(n66922), .Z(n62628) );
  NOR U82811 ( .A(n66928), .B(n62628), .Z(n62629) );
  XOR U82812 ( .A(n66929), .B(n62629), .Z(n68086) );
  IV U82813 ( .A(n62633), .Z(n62630) );
  NOR U82814 ( .A(n62630), .B(n68089), .Z(n68087) );
  IV U82815 ( .A(n62631), .Z(n62635) );
  NOR U82816 ( .A(n62633), .B(n62632), .Z(n62634) );
  NOR U82817 ( .A(n62635), .B(n62634), .Z(n62636) );
  NOR U82818 ( .A(n68087), .B(n62636), .Z(n62637) );
  XOR U82819 ( .A(n68086), .B(n62637), .Z(n72944) );
  XOR U82820 ( .A(n66920), .B(n72944), .Z(n62648) );
  IV U82821 ( .A(n62648), .Z(n68100) );
  IV U82822 ( .A(n62638), .Z(n62640) );
  IV U82823 ( .A(n62639), .Z(n62655) );
  NOR U82824 ( .A(n62640), .B(n62655), .Z(n62641) );
  IV U82825 ( .A(n62641), .Z(n62649) );
  NOR U82826 ( .A(n68100), .B(n62649), .Z(n71751) );
  IV U82827 ( .A(n62642), .Z(n62643) );
  NOR U82828 ( .A(n62643), .B(n62646), .Z(n68102) );
  IV U82829 ( .A(n62644), .Z(n62645) );
  NOR U82830 ( .A(n62646), .B(n62645), .Z(n62647) );
  IV U82831 ( .A(n62647), .Z(n68101) );
  XOR U82832 ( .A(n68101), .B(n62648), .Z(n68103) );
  IV U82833 ( .A(n68103), .Z(n62650) );
  XOR U82834 ( .A(n68102), .B(n62650), .Z(n62652) );
  NOR U82835 ( .A(n62650), .B(n62649), .Z(n62651) );
  NOR U82836 ( .A(n62652), .B(n62651), .Z(n62653) );
  NOR U82837 ( .A(n71751), .B(n62653), .Z(n68115) );
  IV U82838 ( .A(n62654), .Z(n62656) );
  NOR U82839 ( .A(n62656), .B(n62655), .Z(n62657) );
  IV U82840 ( .A(n62657), .Z(n68116) );
  XOR U82841 ( .A(n68115), .B(n68116), .Z(n68120) );
  XOR U82842 ( .A(n68119), .B(n68120), .Z(n68123) );
  XOR U82843 ( .A(n68122), .B(n68123), .Z(n66919) );
  XOR U82844 ( .A(n66917), .B(n66919), .Z(n68133) );
  XOR U82845 ( .A(n68132), .B(n68133), .Z(n62667) );
  IV U82846 ( .A(n62667), .Z(n62663) );
  IV U82847 ( .A(n62658), .Z(n62661) );
  NOR U82848 ( .A(n62665), .B(n62659), .Z(n62660) );
  IV U82849 ( .A(n62660), .Z(n62677) );
  NOR U82850 ( .A(n62661), .B(n62677), .Z(n62670) );
  IV U82851 ( .A(n62670), .Z(n62662) );
  NOR U82852 ( .A(n62663), .B(n62662), .Z(n71740) );
  NOR U82853 ( .A(n62665), .B(n62664), .Z(n62668) );
  IV U82854 ( .A(n62668), .Z(n62666) );
  NOR U82855 ( .A(n62666), .B(n66919), .Z(n72961) );
  NOR U82856 ( .A(n62668), .B(n62667), .Z(n62669) );
  NOR U82857 ( .A(n72961), .B(n62669), .Z(n66910) );
  NOR U82858 ( .A(n62670), .B(n66910), .Z(n62671) );
  NOR U82859 ( .A(n71740), .B(n62671), .Z(n62672) );
  IV U82860 ( .A(n62672), .Z(n66916) );
  IV U82861 ( .A(n62673), .Z(n62675) );
  NOR U82862 ( .A(n62675), .B(n62674), .Z(n66909) );
  IV U82863 ( .A(n62676), .Z(n62678) );
  NOR U82864 ( .A(n62678), .B(n62677), .Z(n66914) );
  NOR U82865 ( .A(n66909), .B(n66914), .Z(n62679) );
  XOR U82866 ( .A(n66916), .B(n62679), .Z(n68137) );
  IV U82867 ( .A(n68137), .Z(n66908) );
  IV U82868 ( .A(n62680), .Z(n68139) );
  NOR U82869 ( .A(n62681), .B(n68139), .Z(n62690) );
  IV U82870 ( .A(n62690), .Z(n62682) );
  NOR U82871 ( .A(n66908), .B(n62682), .Z(n66902) );
  IV U82872 ( .A(n62683), .Z(n62684) );
  NOR U82873 ( .A(n62684), .B(n62686), .Z(n66906) );
  IV U82874 ( .A(n62685), .Z(n62687) );
  NOR U82875 ( .A(n62687), .B(n62686), .Z(n68136) );
  NOR U82876 ( .A(n66906), .B(n68136), .Z(n62688) );
  XOR U82877 ( .A(n68137), .B(n62688), .Z(n66899) );
  IV U82878 ( .A(n66899), .Z(n62689) );
  NOR U82879 ( .A(n62690), .B(n62689), .Z(n62691) );
  NOR U82880 ( .A(n66902), .B(n62691), .Z(n66895) );
  IV U82881 ( .A(n62692), .Z(n62694) );
  NOR U82882 ( .A(n62694), .B(n62693), .Z(n66898) );
  IV U82883 ( .A(n62695), .Z(n62697) );
  NOR U82884 ( .A(n62697), .B(n62696), .Z(n66894) );
  NOR U82885 ( .A(n66898), .B(n66894), .Z(n62698) );
  XOR U82886 ( .A(n66895), .B(n62698), .Z(n68149) );
  IV U82887 ( .A(n62699), .Z(n62700) );
  NOR U82888 ( .A(n62701), .B(n62700), .Z(n68147) );
  XOR U82889 ( .A(n68149), .B(n68147), .Z(n66892) );
  XOR U82890 ( .A(n66890), .B(n66892), .Z(n68156) );
  XOR U82891 ( .A(n62702), .B(n68156), .Z(n68159) );
  NOR U82892 ( .A(n62703), .B(n68160), .Z(n62707) );
  IV U82893 ( .A(n62704), .Z(n62706) );
  IV U82894 ( .A(n62705), .Z(n62712) );
  NOR U82895 ( .A(n62706), .B(n62712), .Z(n66888) );
  NOR U82896 ( .A(n62707), .B(n66888), .Z(n62708) );
  XOR U82897 ( .A(n68159), .B(n62708), .Z(n66881) );
  IV U82898 ( .A(n62709), .Z(n62710) );
  NOR U82899 ( .A(n62717), .B(n62710), .Z(n66882) );
  IV U82900 ( .A(n62711), .Z(n62713) );
  NOR U82901 ( .A(n62713), .B(n62712), .Z(n66885) );
  NOR U82902 ( .A(n66882), .B(n66885), .Z(n62714) );
  XOR U82903 ( .A(n66881), .B(n62714), .Z(n68170) );
  IV U82904 ( .A(n62715), .Z(n62716) );
  NOR U82905 ( .A(n62717), .B(n62716), .Z(n68168) );
  XOR U82906 ( .A(n68170), .B(n68168), .Z(n68176) );
  IV U82907 ( .A(n62718), .Z(n62720) );
  NOR U82908 ( .A(n62720), .B(n62719), .Z(n68171) );
  IV U82909 ( .A(n62721), .Z(n62722) );
  NOR U82910 ( .A(n62723), .B(n62722), .Z(n68175) );
  NOR U82911 ( .A(n68171), .B(n68175), .Z(n62724) );
  XOR U82912 ( .A(n68176), .B(n62724), .Z(n66875) );
  IV U82913 ( .A(n62725), .Z(n62727) );
  NOR U82914 ( .A(n62727), .B(n62726), .Z(n66878) );
  IV U82915 ( .A(n62728), .Z(n62729) );
  NOR U82916 ( .A(n62730), .B(n62729), .Z(n66876) );
  NOR U82917 ( .A(n66878), .B(n66876), .Z(n62731) );
  XOR U82918 ( .A(n66875), .B(n62731), .Z(n66866) );
  NOR U82919 ( .A(n62732), .B(n66865), .Z(n62733) );
  NOR U82920 ( .A(n62733), .B(n66867), .Z(n62734) );
  XOR U82921 ( .A(n66866), .B(n62734), .Z(n68181) );
  IV U82922 ( .A(n62735), .Z(n62736) );
  NOR U82923 ( .A(n62737), .B(n62736), .Z(n68179) );
  XOR U82924 ( .A(n68181), .B(n68179), .Z(n68184) );
  XOR U82925 ( .A(n68182), .B(n68184), .Z(n66862) );
  XOR U82926 ( .A(n66860), .B(n66862), .Z(n68187) );
  IV U82927 ( .A(n62738), .Z(n62739) );
  NOR U82928 ( .A(n62740), .B(n62739), .Z(n66863) );
  IV U82929 ( .A(n62741), .Z(n62743) );
  NOR U82930 ( .A(n62743), .B(n62742), .Z(n68186) );
  NOR U82931 ( .A(n66863), .B(n68186), .Z(n62744) );
  XOR U82932 ( .A(n68187), .B(n62744), .Z(n66854) );
  XOR U82933 ( .A(n62745), .B(n66854), .Z(n66852) );
  XOR U82934 ( .A(n66851), .B(n66852), .Z(n66845) );
  IV U82935 ( .A(n62746), .Z(n66848) );
  NOR U82936 ( .A(n62747), .B(n66848), .Z(n62753) );
  NOR U82937 ( .A(n62749), .B(n62748), .Z(n66844) );
  NOR U82938 ( .A(n62753), .B(n66844), .Z(n62750) );
  XOR U82939 ( .A(n66845), .B(n62750), .Z(n62751) );
  NOR U82940 ( .A(n62752), .B(n62751), .Z(n62756) );
  IV U82941 ( .A(n62752), .Z(n62755) );
  XOR U82942 ( .A(n62753), .B(n66845), .Z(n62754) );
  NOR U82943 ( .A(n62755), .B(n62754), .Z(n73055) );
  NOR U82944 ( .A(n62756), .B(n73055), .Z(n66841) );
  XOR U82945 ( .A(n62757), .B(n66841), .Z(n66837) );
  IV U82946 ( .A(n62758), .Z(n62759) );
  NOR U82947 ( .A(n62765), .B(n62759), .Z(n66835) );
  XOR U82948 ( .A(n66837), .B(n66835), .Z(n66839) );
  IV U82949 ( .A(n62760), .Z(n62762) );
  NOR U82950 ( .A(n62762), .B(n62761), .Z(n66830) );
  IV U82951 ( .A(n62763), .Z(n62764) );
  NOR U82952 ( .A(n62765), .B(n62764), .Z(n66838) );
  NOR U82953 ( .A(n66830), .B(n66838), .Z(n62766) );
  XOR U82954 ( .A(n66839), .B(n62766), .Z(n62767) );
  IV U82955 ( .A(n62767), .Z(n78562) );
  XOR U82956 ( .A(n66832), .B(n78562), .Z(n66822) );
  XOR U82957 ( .A(n62768), .B(n66822), .Z(n62769) );
  IV U82958 ( .A(n62769), .Z(n66819) );
  IV U82959 ( .A(n62770), .Z(n62772) );
  NOR U82960 ( .A(n62772), .B(n62771), .Z(n62773) );
  IV U82961 ( .A(n62773), .Z(n66818) );
  XOR U82962 ( .A(n66819), .B(n66818), .Z(n62774) );
  NOR U82963 ( .A(n62775), .B(n62774), .Z(n62777) );
  IV U82964 ( .A(n62775), .Z(n62776) );
  NOR U82965 ( .A(n62776), .B(n66822), .Z(n71676) );
  NOR U82966 ( .A(n62777), .B(n71676), .Z(n66815) );
  IV U82967 ( .A(n62778), .Z(n62779) );
  NOR U82968 ( .A(n62780), .B(n62779), .Z(n68200) );
  IV U82969 ( .A(n62781), .Z(n62783) );
  NOR U82970 ( .A(n62783), .B(n62782), .Z(n66816) );
  NOR U82971 ( .A(n68200), .B(n66816), .Z(n62784) );
  XOR U82972 ( .A(n66815), .B(n62784), .Z(n66810) );
  XOR U82973 ( .A(n66808), .B(n66810), .Z(n68205) );
  IV U82974 ( .A(n62785), .Z(n62789) );
  NOR U82975 ( .A(n62786), .B(n62800), .Z(n62787) );
  IV U82976 ( .A(n62787), .Z(n62788) );
  NOR U82977 ( .A(n62789), .B(n62788), .Z(n66806) );
  IV U82978 ( .A(n62790), .Z(n66812) );
  NOR U82979 ( .A(n62791), .B(n66812), .Z(n62794) );
  IV U82980 ( .A(n62792), .Z(n62793) );
  NOR U82981 ( .A(n62800), .B(n62793), .Z(n68204) );
  NOR U82982 ( .A(n62794), .B(n68204), .Z(n62795) );
  IV U82983 ( .A(n62795), .Z(n62796) );
  NOR U82984 ( .A(n66806), .B(n62796), .Z(n62797) );
  XOR U82985 ( .A(n68205), .B(n62797), .Z(n66802) );
  IV U82986 ( .A(n62798), .Z(n62804) );
  IV U82987 ( .A(n62799), .Z(n62801) );
  NOR U82988 ( .A(n62801), .B(n62800), .Z(n62802) );
  IV U82989 ( .A(n62802), .Z(n62803) );
  NOR U82990 ( .A(n62804), .B(n62803), .Z(n62805) );
  IV U82991 ( .A(n62805), .Z(n66803) );
  XOR U82992 ( .A(n66802), .B(n66803), .Z(n71665) );
  XOR U82993 ( .A(n71667), .B(n71665), .Z(n66796) );
  XOR U82994 ( .A(n66798), .B(n66796), .Z(n66800) );
  XOR U82995 ( .A(n66799), .B(n66800), .Z(n71660) );
  XOR U82996 ( .A(n66791), .B(n71660), .Z(n66789) );
  XOR U82997 ( .A(n62806), .B(n66789), .Z(n66787) );
  XOR U82998 ( .A(n62807), .B(n66787), .Z(n68215) );
  XOR U82999 ( .A(n62808), .B(n68215), .Z(n66773) );
  IV U83000 ( .A(n62809), .Z(n62811) );
  NOR U83001 ( .A(n62811), .B(n62810), .Z(n68217) );
  NOR U83002 ( .A(n62812), .B(n66774), .Z(n62813) );
  NOR U83003 ( .A(n68217), .B(n62813), .Z(n62814) );
  XOR U83004 ( .A(n66773), .B(n62814), .Z(n66769) );
  XOR U83005 ( .A(n66767), .B(n66769), .Z(n68229) );
  XOR U83006 ( .A(n62815), .B(n68229), .Z(n68231) );
  XOR U83007 ( .A(n68232), .B(n68231), .Z(n66765) );
  IV U83008 ( .A(n62816), .Z(n62818) );
  NOR U83009 ( .A(n62818), .B(n62817), .Z(n68233) );
  IV U83010 ( .A(n62819), .Z(n62821) );
  NOR U83011 ( .A(n62821), .B(n62820), .Z(n66764) );
  NOR U83012 ( .A(n68233), .B(n66764), .Z(n62822) );
  XOR U83013 ( .A(n66765), .B(n62822), .Z(n68238) );
  IV U83014 ( .A(n62823), .Z(n62824) );
  NOR U83015 ( .A(n62825), .B(n62824), .Z(n62826) );
  IV U83016 ( .A(n62826), .Z(n68239) );
  XOR U83017 ( .A(n68238), .B(n68239), .Z(n66762) );
  XOR U83018 ( .A(n66760), .B(n66762), .Z(n68252) );
  XOR U83019 ( .A(n62827), .B(n68252), .Z(n66752) );
  XOR U83020 ( .A(n62828), .B(n66752), .Z(n66751) );
  NOR U83021 ( .A(n62835), .B(n66751), .Z(n71632) );
  IV U83022 ( .A(n62829), .Z(n62831) );
  NOR U83023 ( .A(n62831), .B(n62830), .Z(n68256) );
  IV U83024 ( .A(n62832), .Z(n62833) );
  NOR U83025 ( .A(n62834), .B(n62833), .Z(n66749) );
  XOR U83026 ( .A(n66751), .B(n66749), .Z(n68257) );
  IV U83027 ( .A(n68257), .Z(n62836) );
  XOR U83028 ( .A(n68256), .B(n62836), .Z(n62838) );
  NOR U83029 ( .A(n62836), .B(n62835), .Z(n62837) );
  NOR U83030 ( .A(n62838), .B(n62837), .Z(n62839) );
  NOR U83031 ( .A(n71632), .B(n62839), .Z(n66747) );
  XOR U83032 ( .A(n62840), .B(n66747), .Z(n68266) );
  XOR U83033 ( .A(n62841), .B(n68266), .Z(n66740) );
  XOR U83034 ( .A(n62842), .B(n66740), .Z(n66734) );
  XOR U83035 ( .A(n66732), .B(n66734), .Z(n66736) );
  IV U83036 ( .A(n62843), .Z(n62845) );
  NOR U83037 ( .A(n62845), .B(n62844), .Z(n66730) );
  NOR U83038 ( .A(n66735), .B(n66730), .Z(n62846) );
  XOR U83039 ( .A(n66736), .B(n62846), .Z(n68277) );
  NOR U83040 ( .A(n62847), .B(n68278), .Z(n62851) );
  IV U83041 ( .A(n62848), .Z(n62850) );
  IV U83042 ( .A(n62849), .Z(n62854) );
  NOR U83043 ( .A(n62850), .B(n62854), .Z(n68287) );
  NOR U83044 ( .A(n62851), .B(n68287), .Z(n62852) );
  XOR U83045 ( .A(n68277), .B(n62852), .Z(n66728) );
  IV U83046 ( .A(n62853), .Z(n62860) );
  NOR U83047 ( .A(n62855), .B(n62854), .Z(n62856) );
  IV U83048 ( .A(n62856), .Z(n62857) );
  NOR U83049 ( .A(n62858), .B(n62857), .Z(n62859) );
  IV U83050 ( .A(n62859), .Z(n62862) );
  NOR U83051 ( .A(n62860), .B(n62862), .Z(n66726) );
  XOR U83052 ( .A(n66728), .B(n66726), .Z(n68292) );
  IV U83053 ( .A(n62861), .Z(n62863) );
  NOR U83054 ( .A(n62863), .B(n62862), .Z(n68290) );
  XOR U83055 ( .A(n68292), .B(n68290), .Z(n68294) );
  NOR U83056 ( .A(n62864), .B(n68295), .Z(n62868) );
  IV U83057 ( .A(n62865), .Z(n62867) );
  IV U83058 ( .A(n62866), .Z(n62871) );
  NOR U83059 ( .A(n62867), .B(n62871), .Z(n66724) );
  NOR U83060 ( .A(n62868), .B(n66724), .Z(n62869) );
  XOR U83061 ( .A(n68294), .B(n62869), .Z(n66718) );
  IV U83062 ( .A(n62870), .Z(n62872) );
  NOR U83063 ( .A(n62872), .B(n62871), .Z(n66722) );
  IV U83064 ( .A(n62873), .Z(n62875) );
  NOR U83065 ( .A(n62875), .B(n62874), .Z(n66719) );
  NOR U83066 ( .A(n66722), .B(n66719), .Z(n62876) );
  XOR U83067 ( .A(n66718), .B(n62876), .Z(n66716) );
  NOR U83068 ( .A(n62878), .B(n62877), .Z(n66715) );
  IV U83069 ( .A(n62879), .Z(n62881) );
  IV U83070 ( .A(n62880), .Z(n62886) );
  NOR U83071 ( .A(n62881), .B(n62886), .Z(n66713) );
  NOR U83072 ( .A(n66715), .B(n66713), .Z(n62882) );
  XOR U83073 ( .A(n66716), .B(n62882), .Z(n66703) );
  IV U83074 ( .A(n62883), .Z(n62884) );
  NOR U83075 ( .A(n62885), .B(n62884), .Z(n66704) );
  NOR U83076 ( .A(n62887), .B(n62886), .Z(n62888) );
  IV U83077 ( .A(n62888), .Z(n66708) );
  NOR U83078 ( .A(n66706), .B(n66708), .Z(n62889) );
  NOR U83079 ( .A(n66704), .B(n62889), .Z(n62890) );
  XOR U83080 ( .A(n66703), .B(n62890), .Z(n73226) );
  IV U83081 ( .A(n62891), .Z(n62892) );
  NOR U83082 ( .A(n62894), .B(n62892), .Z(n73225) );
  IV U83083 ( .A(n62893), .Z(n62898) );
  NOR U83084 ( .A(n62895), .B(n62894), .Z(n62896) );
  IV U83085 ( .A(n62896), .Z(n62897) );
  NOR U83086 ( .A(n62898), .B(n62897), .Z(n73231) );
  NOR U83087 ( .A(n73225), .B(n73231), .Z(n66702) );
  XOR U83088 ( .A(n73226), .B(n66702), .Z(n62899) );
  IV U83089 ( .A(n62899), .Z(n66697) );
  XOR U83090 ( .A(n66696), .B(n66697), .Z(n66700) );
  XOR U83091 ( .A(n62900), .B(n66700), .Z(n68303) );
  XOR U83092 ( .A(n62901), .B(n68303), .Z(n66689) );
  XOR U83093 ( .A(n66687), .B(n66689), .Z(n66692) );
  XOR U83094 ( .A(n62902), .B(n66692), .Z(n68317) );
  XOR U83095 ( .A(n68318), .B(n68317), .Z(n68320) );
  IV U83096 ( .A(n62903), .Z(n62905) );
  NOR U83097 ( .A(n62905), .B(n62904), .Z(n68319) );
  IV U83098 ( .A(n62906), .Z(n62908) );
  IV U83099 ( .A(n62907), .Z(n62914) );
  NOR U83100 ( .A(n62908), .B(n62914), .Z(n68323) );
  NOR U83101 ( .A(n68319), .B(n68323), .Z(n62909) );
  XOR U83102 ( .A(n68320), .B(n62909), .Z(n66681) );
  IV U83103 ( .A(n62910), .Z(n62911) );
  NOR U83104 ( .A(n62912), .B(n62911), .Z(n68330) );
  IV U83105 ( .A(n62913), .Z(n62915) );
  NOR U83106 ( .A(n62915), .B(n62914), .Z(n66682) );
  NOR U83107 ( .A(n68330), .B(n66682), .Z(n62916) );
  XOR U83108 ( .A(n66681), .B(n62916), .Z(n66679) );
  IV U83109 ( .A(n62917), .Z(n62918) );
  NOR U83110 ( .A(n62918), .B(n62924), .Z(n66677) );
  XOR U83111 ( .A(n66679), .B(n66677), .Z(n68329) );
  IV U83112 ( .A(n62919), .Z(n62921) );
  NOR U83113 ( .A(n62921), .B(n62920), .Z(n66674) );
  IV U83114 ( .A(n62922), .Z(n62923) );
  NOR U83115 ( .A(n62924), .B(n62923), .Z(n68327) );
  NOR U83116 ( .A(n66674), .B(n68327), .Z(n62925) );
  XOR U83117 ( .A(n68329), .B(n62925), .Z(n68339) );
  XOR U83118 ( .A(n62926), .B(n68339), .Z(n66673) );
  XOR U83119 ( .A(n62927), .B(n66673), .Z(n66667) );
  XOR U83120 ( .A(n62928), .B(n66667), .Z(n68355) );
  XOR U83121 ( .A(n62929), .B(n68355), .Z(n68349) );
  XOR U83122 ( .A(n62930), .B(n68349), .Z(n66656) );
  XOR U83123 ( .A(n66654), .B(n66656), .Z(n66658) );
  IV U83124 ( .A(n66658), .Z(n62938) );
  IV U83125 ( .A(n62931), .Z(n62933) );
  NOR U83126 ( .A(n62933), .B(n62932), .Z(n66657) );
  IV U83127 ( .A(n62934), .Z(n62936) );
  NOR U83128 ( .A(n62936), .B(n62935), .Z(n66651) );
  NOR U83129 ( .A(n66657), .B(n66651), .Z(n62937) );
  XOR U83130 ( .A(n62938), .B(n62937), .Z(n66648) );
  XOR U83131 ( .A(n66646), .B(n66648), .Z(n68370) );
  XOR U83132 ( .A(n62939), .B(n68370), .Z(n66641) );
  XOR U83133 ( .A(n62940), .B(n66641), .Z(n66638) );
  XOR U83134 ( .A(n66637), .B(n66638), .Z(n66627) );
  XOR U83135 ( .A(n62941), .B(n66627), .Z(n66615) );
  XOR U83136 ( .A(n62942), .B(n66615), .Z(n66613) );
  IV U83137 ( .A(n62943), .Z(n62944) );
  NOR U83138 ( .A(n62944), .B(n62946), .Z(n66612) );
  IV U83139 ( .A(n62945), .Z(n62947) );
  NOR U83140 ( .A(n62947), .B(n62946), .Z(n66610) );
  NOR U83141 ( .A(n66612), .B(n66610), .Z(n62948) );
  XOR U83142 ( .A(n66613), .B(n62948), .Z(n66604) );
  XOR U83143 ( .A(n62949), .B(n66604), .Z(n66600) );
  XOR U83144 ( .A(n66599), .B(n66600), .Z(n68383) );
  XOR U83145 ( .A(n62950), .B(n68383), .Z(n68379) );
  XOR U83146 ( .A(n62951), .B(n68379), .Z(n66597) );
  IV U83147 ( .A(n62952), .Z(n62954) );
  NOR U83148 ( .A(n62954), .B(n62953), .Z(n62955) );
  IV U83149 ( .A(n62955), .Z(n62959) );
  NOR U83150 ( .A(n66597), .B(n62959), .Z(n73313) );
  IV U83151 ( .A(n62956), .Z(n62958) );
  NOR U83152 ( .A(n62958), .B(n62957), .Z(n66592) );
  XOR U83153 ( .A(n66596), .B(n66597), .Z(n66593) );
  IV U83154 ( .A(n66593), .Z(n62960) );
  XOR U83155 ( .A(n66592), .B(n62960), .Z(n62962) );
  NOR U83156 ( .A(n62960), .B(n62959), .Z(n62961) );
  NOR U83157 ( .A(n62962), .B(n62961), .Z(n62963) );
  NOR U83158 ( .A(n73313), .B(n62963), .Z(n66586) );
  XOR U83159 ( .A(n62964), .B(n66586), .Z(n68398) );
  XOR U83160 ( .A(n62965), .B(n68398), .Z(n66576) );
  XOR U83161 ( .A(n62966), .B(n66576), .Z(n68400) );
  IV U83162 ( .A(n62967), .Z(n62969) );
  NOR U83163 ( .A(n62969), .B(n62968), .Z(n66571) );
  IV U83164 ( .A(n62970), .Z(n62971) );
  NOR U83165 ( .A(n62971), .B(n62974), .Z(n68399) );
  NOR U83166 ( .A(n66571), .B(n68399), .Z(n62972) );
  XOR U83167 ( .A(n68400), .B(n62972), .Z(n68405) );
  IV U83168 ( .A(n62973), .Z(n62975) );
  NOR U83169 ( .A(n62975), .B(n62974), .Z(n68403) );
  XOR U83170 ( .A(n68405), .B(n68403), .Z(n68410) );
  XOR U83171 ( .A(n62976), .B(n68410), .Z(n62977) );
  IV U83172 ( .A(n62977), .Z(n68413) );
  XOR U83173 ( .A(n68412), .B(n68413), .Z(n66569) );
  XOR U83174 ( .A(n66566), .B(n66569), .Z(n68421) );
  IV U83175 ( .A(n62978), .Z(n62980) );
  NOR U83176 ( .A(n62980), .B(n62979), .Z(n66568) );
  IV U83177 ( .A(n62981), .Z(n62982) );
  NOR U83178 ( .A(n62982), .B(n62990), .Z(n68419) );
  NOR U83179 ( .A(n66568), .B(n68419), .Z(n62983) );
  XOR U83180 ( .A(n68421), .B(n62983), .Z(n62984) );
  IV U83181 ( .A(n62984), .Z(n68425) );
  IV U83182 ( .A(n62985), .Z(n62986) );
  NOR U83183 ( .A(n62987), .B(n62986), .Z(n68423) );
  IV U83184 ( .A(n62988), .Z(n62989) );
  NOR U83185 ( .A(n62990), .B(n62989), .Z(n68417) );
  NOR U83186 ( .A(n68423), .B(n68417), .Z(n62991) );
  XOR U83187 ( .A(n68425), .B(n62991), .Z(n66564) );
  IV U83188 ( .A(n62992), .Z(n62993) );
  NOR U83189 ( .A(n62994), .B(n62993), .Z(n66563) );
  IV U83190 ( .A(n62995), .Z(n62996) );
  NOR U83191 ( .A(n62997), .B(n62996), .Z(n68429) );
  NOR U83192 ( .A(n66563), .B(n68429), .Z(n62998) );
  XOR U83193 ( .A(n66564), .B(n62998), .Z(n66560) );
  XOR U83194 ( .A(n66559), .B(n66560), .Z(n68428) );
  IV U83195 ( .A(n62999), .Z(n63001) );
  IV U83196 ( .A(n63000), .Z(n63004) );
  NOR U83197 ( .A(n63001), .B(n63004), .Z(n63002) );
  IV U83198 ( .A(n63002), .Z(n63009) );
  NOR U83199 ( .A(n68428), .B(n63009), .Z(n71490) );
  IV U83200 ( .A(n63003), .Z(n63005) );
  NOR U83201 ( .A(n63005), .B(n63004), .Z(n68426) );
  XOR U83202 ( .A(n68428), .B(n68426), .Z(n66555) );
  IV U83203 ( .A(n63006), .Z(n63007) );
  NOR U83204 ( .A(n63008), .B(n63007), .Z(n63010) );
  IV U83205 ( .A(n63010), .Z(n66554) );
  XOR U83206 ( .A(n66555), .B(n66554), .Z(n63012) );
  NOR U83207 ( .A(n63010), .B(n63009), .Z(n63011) );
  NOR U83208 ( .A(n63012), .B(n63011), .Z(n63013) );
  NOR U83209 ( .A(n71490), .B(n63013), .Z(n66551) );
  XOR U83210 ( .A(n63014), .B(n66551), .Z(n66549) );
  XOR U83211 ( .A(n66547), .B(n66549), .Z(n66543) );
  IV U83212 ( .A(n63015), .Z(n63017) );
  NOR U83213 ( .A(n63017), .B(n63016), .Z(n66541) );
  XOR U83214 ( .A(n66543), .B(n66541), .Z(n66545) );
  XOR U83215 ( .A(n66544), .B(n66545), .Z(n68442) );
  XOR U83216 ( .A(n68441), .B(n68442), .Z(n68444) );
  XOR U83217 ( .A(n68445), .B(n68444), .Z(n63018) );
  XOR U83218 ( .A(n66539), .B(n63018), .Z(n68447) );
  XOR U83219 ( .A(n68446), .B(n68447), .Z(n68450) );
  NOR U83220 ( .A(n63019), .B(n68450), .Z(n71467) );
  NOR U83221 ( .A(n63027), .B(n71467), .Z(n63020) );
  IV U83222 ( .A(n63020), .Z(n63026) );
  IV U83223 ( .A(n63021), .Z(n63022) );
  NOR U83224 ( .A(n63023), .B(n63022), .Z(n68449) );
  XOR U83225 ( .A(n68449), .B(n68450), .Z(n66532) );
  IV U83226 ( .A(n66532), .Z(n63029) );
  NOR U83227 ( .A(n63024), .B(n63029), .Z(n63025) );
  NOR U83228 ( .A(n63026), .B(n63025), .Z(n63031) );
  IV U83229 ( .A(n63027), .Z(n63028) );
  NOR U83230 ( .A(n63029), .B(n63028), .Z(n63030) );
  NOR U83231 ( .A(n63031), .B(n63030), .Z(n66530) );
  XOR U83232 ( .A(n63032), .B(n66530), .Z(n66516) );
  XOR U83233 ( .A(n63033), .B(n66516), .Z(n66511) );
  XOR U83234 ( .A(n66510), .B(n66511), .Z(n66506) );
  IV U83235 ( .A(n63034), .Z(n63035) );
  NOR U83236 ( .A(n63036), .B(n63035), .Z(n66512) );
  IV U83237 ( .A(n63037), .Z(n63039) );
  NOR U83238 ( .A(n63039), .B(n63038), .Z(n66507) );
  NOR U83239 ( .A(n66512), .B(n66507), .Z(n63040) );
  XOR U83240 ( .A(n66506), .B(n63040), .Z(n68456) );
  XOR U83241 ( .A(n68454), .B(n68456), .Z(n68458) );
  XOR U83242 ( .A(n68457), .B(n68458), .Z(n66503) );
  XOR U83243 ( .A(n66501), .B(n66503), .Z(n68465) );
  XOR U83244 ( .A(n63041), .B(n68465), .Z(n68462) );
  XOR U83245 ( .A(n68463), .B(n68462), .Z(n68471) );
  XOR U83246 ( .A(n68469), .B(n68471), .Z(n68474) );
  XOR U83247 ( .A(n63042), .B(n68474), .Z(n68477) );
  IV U83248 ( .A(n63043), .Z(n63045) );
  NOR U83249 ( .A(n63045), .B(n63044), .Z(n66497) );
  IV U83250 ( .A(n63046), .Z(n63056) );
  NOR U83251 ( .A(n63048), .B(n63047), .Z(n63049) );
  IV U83252 ( .A(n63049), .Z(n63054) );
  NOR U83253 ( .A(n63051), .B(n63050), .Z(n63052) );
  IV U83254 ( .A(n63052), .Z(n63053) );
  NOR U83255 ( .A(n63054), .B(n63053), .Z(n63055) );
  IV U83256 ( .A(n63055), .Z(n63061) );
  NOR U83257 ( .A(n63056), .B(n63061), .Z(n68476) );
  NOR U83258 ( .A(n66497), .B(n68476), .Z(n63057) );
  XOR U83259 ( .A(n68477), .B(n63057), .Z(n68482) );
  IV U83260 ( .A(n68482), .Z(n63064) );
  IV U83261 ( .A(n63058), .Z(n66491) );
  NOR U83262 ( .A(n66491), .B(n63059), .Z(n66495) );
  IV U83263 ( .A(n63060), .Z(n63062) );
  NOR U83264 ( .A(n63062), .B(n63061), .Z(n68480) );
  NOR U83265 ( .A(n66495), .B(n68480), .Z(n63063) );
  XOR U83266 ( .A(n63064), .B(n63063), .Z(n68485) );
  NOR U83267 ( .A(n63066), .B(n63065), .Z(n68484) );
  IV U83268 ( .A(n63067), .Z(n63069) );
  NOR U83269 ( .A(n63069), .B(n63068), .Z(n66488) );
  NOR U83270 ( .A(n68484), .B(n66488), .Z(n63070) );
  XOR U83271 ( .A(n68485), .B(n63070), .Z(n63076) );
  IV U83272 ( .A(n63076), .Z(n63071) );
  NOR U83273 ( .A(n63072), .B(n63071), .Z(n71444) );
  IV U83274 ( .A(n63073), .Z(n63075) );
  NOR U83275 ( .A(n63075), .B(n63074), .Z(n63077) );
  NOR U83276 ( .A(n63077), .B(n63076), .Z(n63080) );
  IV U83277 ( .A(n63077), .Z(n63079) );
  XOR U83278 ( .A(n68484), .B(n68485), .Z(n63078) );
  NOR U83279 ( .A(n63079), .B(n63078), .Z(n71441) );
  NOR U83280 ( .A(n63080), .B(n71441), .Z(n68491) );
  NOR U83281 ( .A(n63081), .B(n68491), .Z(n63082) );
  NOR U83282 ( .A(n71444), .B(n63082), .Z(n68500) );
  XOR U83283 ( .A(n63083), .B(n68500), .Z(n66487) );
  XOR U83284 ( .A(n66485), .B(n66487), .Z(n68507) );
  XOR U83285 ( .A(n66484), .B(n68507), .Z(n63084) );
  IV U83286 ( .A(n63084), .Z(n66479) );
  XOR U83287 ( .A(n66478), .B(n66479), .Z(n66482) );
  XOR U83288 ( .A(n66481), .B(n66482), .Z(n71413) );
  IV U83289 ( .A(n63085), .Z(n63086) );
  NOR U83290 ( .A(n63086), .B(n63096), .Z(n66472) );
  IV U83291 ( .A(n63087), .Z(n71416) );
  NOR U83292 ( .A(n63088), .B(n71416), .Z(n63091) );
  IV U83293 ( .A(n63089), .Z(n63090) );
  NOR U83294 ( .A(n63090), .B(n63096), .Z(n73460) );
  NOR U83295 ( .A(n63091), .B(n73460), .Z(n66477) );
  IV U83296 ( .A(n66477), .Z(n63092) );
  NOR U83297 ( .A(n66472), .B(n63092), .Z(n63093) );
  XOR U83298 ( .A(n71413), .B(n63093), .Z(n63094) );
  IV U83299 ( .A(n63094), .Z(n66476) );
  IV U83300 ( .A(n63095), .Z(n63097) );
  NOR U83301 ( .A(n63097), .B(n63096), .Z(n66474) );
  XOR U83302 ( .A(n66476), .B(n66474), .Z(n73468) );
  IV U83303 ( .A(n63098), .Z(n63099) );
  NOR U83304 ( .A(n66467), .B(n63099), .Z(n66459) );
  NOR U83305 ( .A(n73473), .B(n73471), .Z(n66462) );
  NOR U83306 ( .A(n66459), .B(n66462), .Z(n63100) );
  XOR U83307 ( .A(n73468), .B(n63100), .Z(n63113) );
  IV U83308 ( .A(n63101), .Z(n66456) );
  NOR U83309 ( .A(n63102), .B(n66456), .Z(n63103) );
  NOR U83310 ( .A(n63113), .B(n63103), .Z(n63106) );
  IV U83311 ( .A(n63103), .Z(n63104) );
  XOR U83312 ( .A(n66459), .B(n73468), .Z(n66455) );
  NOR U83313 ( .A(n63104), .B(n66455), .Z(n63105) );
  NOR U83314 ( .A(n63106), .B(n63105), .Z(n68525) );
  IV U83315 ( .A(n63107), .Z(n63109) );
  NOR U83316 ( .A(n63109), .B(n63108), .Z(n63120) );
  IV U83317 ( .A(n63120), .Z(n68526) );
  NOR U83318 ( .A(n68525), .B(n68526), .Z(n63122) );
  IV U83319 ( .A(n63110), .Z(n63112) );
  NOR U83320 ( .A(n63112), .B(n63111), .Z(n63116) );
  IV U83321 ( .A(n63116), .Z(n63115) );
  IV U83322 ( .A(n63113), .Z(n63114) );
  NOR U83323 ( .A(n63115), .B(n63114), .Z(n71398) );
  NOR U83324 ( .A(n68525), .B(n63116), .Z(n63117) );
  NOR U83325 ( .A(n71398), .B(n63117), .Z(n63118) );
  IV U83326 ( .A(n63118), .Z(n63119) );
  NOR U83327 ( .A(n63120), .B(n63119), .Z(n63121) );
  NOR U83328 ( .A(n63122), .B(n63121), .Z(n68529) );
  IV U83329 ( .A(n63123), .Z(n63125) );
  NOR U83330 ( .A(n63125), .B(n63124), .Z(n68528) );
  IV U83331 ( .A(n63126), .Z(n63128) );
  NOR U83332 ( .A(n63128), .B(n63127), .Z(n66452) );
  NOR U83333 ( .A(n68528), .B(n66452), .Z(n63129) );
  XOR U83334 ( .A(n68529), .B(n63129), .Z(n68536) );
  XOR U83335 ( .A(n68537), .B(n68536), .Z(n66450) );
  IV U83336 ( .A(n63130), .Z(n63131) );
  NOR U83337 ( .A(n63134), .B(n63131), .Z(n66448) );
  XOR U83338 ( .A(n66450), .B(n66448), .Z(n68535) );
  IV U83339 ( .A(n63132), .Z(n63133) );
  NOR U83340 ( .A(n63134), .B(n63133), .Z(n68533) );
  XOR U83341 ( .A(n68535), .B(n68533), .Z(n66442) );
  IV U83342 ( .A(n63135), .Z(n63136) );
  NOR U83343 ( .A(n63137), .B(n63136), .Z(n66445) );
  IV U83344 ( .A(n63138), .Z(n63140) );
  NOR U83345 ( .A(n63140), .B(n63139), .Z(n66441) );
  NOR U83346 ( .A(n66445), .B(n66441), .Z(n63141) );
  XOR U83347 ( .A(n66442), .B(n63141), .Z(n66439) );
  IV U83348 ( .A(n63142), .Z(n63143) );
  NOR U83349 ( .A(n63144), .B(n63143), .Z(n71379) );
  IV U83350 ( .A(n63145), .Z(n63146) );
  NOR U83351 ( .A(n63151), .B(n63146), .Z(n71372) );
  NOR U83352 ( .A(n71379), .B(n71372), .Z(n66440) );
  XOR U83353 ( .A(n66439), .B(n66440), .Z(n66437) );
  IV U83354 ( .A(n63147), .Z(n63148) );
  NOR U83355 ( .A(n63149), .B(n63148), .Z(n66436) );
  IV U83356 ( .A(n63150), .Z(n63152) );
  NOR U83357 ( .A(n63152), .B(n63151), .Z(n66434) );
  NOR U83358 ( .A(n66436), .B(n66434), .Z(n63153) );
  XOR U83359 ( .A(n66437), .B(n63153), .Z(n63168) );
  IV U83360 ( .A(n63168), .Z(n63173) );
  IV U83361 ( .A(n63154), .Z(n63155) );
  NOR U83362 ( .A(n63155), .B(n63162), .Z(n63156) );
  IV U83363 ( .A(n63156), .Z(n63176) );
  NOR U83364 ( .A(n63173), .B(n63176), .Z(n73488) );
  IV U83365 ( .A(n63157), .Z(n63158) );
  NOR U83366 ( .A(n63159), .B(n63158), .Z(n68548) );
  IV U83367 ( .A(n63160), .Z(n63161) );
  NOR U83368 ( .A(n63162), .B(n63161), .Z(n63172) );
  IV U83369 ( .A(n63163), .Z(n63164) );
  NOR U83370 ( .A(n63165), .B(n63164), .Z(n63169) );
  IV U83371 ( .A(n63169), .Z(n63167) );
  XOR U83372 ( .A(n66434), .B(n66437), .Z(n63166) );
  NOR U83373 ( .A(n63167), .B(n63166), .Z(n71364) );
  NOR U83374 ( .A(n63169), .B(n63168), .Z(n63170) );
  NOR U83375 ( .A(n71364), .B(n63170), .Z(n63171) );
  NOR U83376 ( .A(n63172), .B(n63171), .Z(n63175) );
  IV U83377 ( .A(n63172), .Z(n63174) );
  NOR U83378 ( .A(n63174), .B(n63173), .Z(n71361) );
  NOR U83379 ( .A(n63175), .B(n71361), .Z(n68549) );
  XOR U83380 ( .A(n68548), .B(n68549), .Z(n63178) );
  NOR U83381 ( .A(n68549), .B(n63176), .Z(n63177) );
  NOR U83382 ( .A(n63178), .B(n63177), .Z(n63179) );
  NOR U83383 ( .A(n73488), .B(n63179), .Z(n71349) );
  IV U83384 ( .A(n71349), .Z(n66431) );
  XOR U83385 ( .A(n71350), .B(n66431), .Z(n68558) );
  XOR U83386 ( .A(n68557), .B(n68558), .Z(n68565) );
  IV U83387 ( .A(n63180), .Z(n63184) );
  NOR U83388 ( .A(n63184), .B(n63181), .Z(n68560) );
  IV U83389 ( .A(n63182), .Z(n63186) );
  XOR U83390 ( .A(n63184), .B(n63183), .Z(n63185) );
  NOR U83391 ( .A(n63186), .B(n63185), .Z(n68564) );
  NOR U83392 ( .A(n68560), .B(n68564), .Z(n63187) );
  XOR U83393 ( .A(n68565), .B(n63187), .Z(n66429) );
  XOR U83394 ( .A(n63188), .B(n66429), .Z(n66427) );
  XOR U83395 ( .A(n63189), .B(n66427), .Z(n66418) );
  XOR U83396 ( .A(n63190), .B(n66418), .Z(n66416) );
  IV U83397 ( .A(n63191), .Z(n63193) );
  NOR U83398 ( .A(n63193), .B(n63192), .Z(n66414) );
  IV U83399 ( .A(n63194), .Z(n63195) );
  NOR U83400 ( .A(n63195), .B(n63199), .Z(n66409) );
  NOR U83401 ( .A(n66414), .B(n66409), .Z(n63196) );
  XOR U83402 ( .A(n66416), .B(n63196), .Z(n66402) );
  NOR U83403 ( .A(n66403), .B(n63197), .Z(n63201) );
  IV U83404 ( .A(n63198), .Z(n63200) );
  NOR U83405 ( .A(n63200), .B(n63199), .Z(n66411) );
  NOR U83406 ( .A(n63201), .B(n66411), .Z(n63202) );
  XOR U83407 ( .A(n66402), .B(n63202), .Z(n66400) );
  XOR U83408 ( .A(n66398), .B(n66400), .Z(n68577) );
  XOR U83409 ( .A(n68576), .B(n68577), .Z(n68583) );
  XOR U83410 ( .A(n63203), .B(n68583), .Z(n66392) );
  XOR U83411 ( .A(n63204), .B(n66392), .Z(n66390) );
  XOR U83412 ( .A(n63205), .B(n66390), .Z(n66387) );
  IV U83413 ( .A(n63206), .Z(n63208) );
  NOR U83414 ( .A(n63208), .B(n63207), .Z(n66386) );
  IV U83415 ( .A(n63209), .Z(n63210) );
  NOR U83416 ( .A(n63210), .B(n63213), .Z(n68588) );
  NOR U83417 ( .A(n66386), .B(n68588), .Z(n63211) );
  XOR U83418 ( .A(n66387), .B(n63211), .Z(n73545) );
  IV U83419 ( .A(n63212), .Z(n63214) );
  NOR U83420 ( .A(n63214), .B(n63213), .Z(n73541) );
  IV U83421 ( .A(n63215), .Z(n63217) );
  IV U83422 ( .A(n63216), .Z(n63220) );
  NOR U83423 ( .A(n63217), .B(n63220), .Z(n73551) );
  NOR U83424 ( .A(n73541), .B(n73551), .Z(n68587) );
  XOR U83425 ( .A(n73545), .B(n68587), .Z(n63218) );
  IV U83426 ( .A(n63218), .Z(n66383) );
  IV U83427 ( .A(n63219), .Z(n63221) );
  NOR U83428 ( .A(n63221), .B(n63220), .Z(n66381) );
  XOR U83429 ( .A(n66383), .B(n66381), .Z(n66372) );
  NOR U83430 ( .A(n66375), .B(n63222), .Z(n63226) );
  IV U83431 ( .A(n63223), .Z(n63225) );
  NOR U83432 ( .A(n63225), .B(n63224), .Z(n66371) );
  NOR U83433 ( .A(n63226), .B(n66371), .Z(n63227) );
  XOR U83434 ( .A(n66372), .B(n63227), .Z(n63228) );
  IV U83435 ( .A(n63228), .Z(n66368) );
  XOR U83436 ( .A(n66366), .B(n66368), .Z(n68594) );
  XOR U83437 ( .A(n63229), .B(n68594), .Z(n66362) );
  IV U83438 ( .A(n63230), .Z(n63231) );
  NOR U83439 ( .A(n63232), .B(n63231), .Z(n68596) );
  NOR U83440 ( .A(n63233), .B(n66363), .Z(n63234) );
  NOR U83441 ( .A(n68596), .B(n63234), .Z(n63235) );
  XOR U83442 ( .A(n66362), .B(n63235), .Z(n68607) );
  XOR U83443 ( .A(n68605), .B(n68607), .Z(n68614) );
  XOR U83444 ( .A(n63236), .B(n68614), .Z(n66357) );
  XOR U83445 ( .A(n66356), .B(n66357), .Z(n68627) );
  XOR U83446 ( .A(n68626), .B(n68627), .Z(n68631) );
  IV U83447 ( .A(n63237), .Z(n63239) );
  NOR U83448 ( .A(n63239), .B(n63238), .Z(n68629) );
  XOR U83449 ( .A(n68631), .B(n68629), .Z(n66354) );
  IV U83450 ( .A(n63240), .Z(n63241) );
  NOR U83451 ( .A(n63242), .B(n63241), .Z(n66353) );
  IV U83452 ( .A(n63243), .Z(n63245) );
  NOR U83453 ( .A(n63245), .B(n63244), .Z(n66351) );
  NOR U83454 ( .A(n66353), .B(n66351), .Z(n63246) );
  XOR U83455 ( .A(n66354), .B(n63246), .Z(n66348) );
  XOR U83456 ( .A(n66349), .B(n66348), .Z(n68636) );
  XOR U83457 ( .A(n68635), .B(n68636), .Z(n66347) );
  XOR U83458 ( .A(n66345), .B(n66347), .Z(n68643) );
  XOR U83459 ( .A(n68642), .B(n68643), .Z(n68646) );
  XOR U83460 ( .A(n63247), .B(n68646), .Z(n66337) );
  XOR U83461 ( .A(n66338), .B(n66337), .Z(n66341) );
  IV U83462 ( .A(n63248), .Z(n63250) );
  NOR U83463 ( .A(n63250), .B(n63249), .Z(n66340) );
  IV U83464 ( .A(n63251), .Z(n63253) );
  NOR U83465 ( .A(n63253), .B(n63252), .Z(n66332) );
  NOR U83466 ( .A(n66340), .B(n66332), .Z(n63254) );
  XOR U83467 ( .A(n66341), .B(n63254), .Z(n63259) );
  IV U83468 ( .A(n63259), .Z(n66335) );
  XOR U83469 ( .A(n66334), .B(n66335), .Z(n63255) );
  NOR U83470 ( .A(n63261), .B(n63255), .Z(n73605) );
  IV U83471 ( .A(n63256), .Z(n63257) );
  NOR U83472 ( .A(n63257), .B(n66328), .Z(n66318) );
  NOR U83473 ( .A(n63258), .B(n66328), .Z(n66322) );
  NOR U83474 ( .A(n66334), .B(n66322), .Z(n63260) );
  XOR U83475 ( .A(n63260), .B(n63259), .Z(n66319) );
  IV U83476 ( .A(n66319), .Z(n63262) );
  XOR U83477 ( .A(n66318), .B(n63262), .Z(n63264) );
  NOR U83478 ( .A(n63262), .B(n63261), .Z(n63263) );
  NOR U83479 ( .A(n63264), .B(n63263), .Z(n63265) );
  NOR U83480 ( .A(n73605), .B(n63265), .Z(n66316) );
  IV U83481 ( .A(n63266), .Z(n63267) );
  NOR U83482 ( .A(n63267), .B(n63272), .Z(n68655) );
  IV U83483 ( .A(n63268), .Z(n63270) );
  NOR U83484 ( .A(n63270), .B(n63269), .Z(n66315) );
  IV U83485 ( .A(n63271), .Z(n63273) );
  NOR U83486 ( .A(n63273), .B(n63272), .Z(n68652) );
  NOR U83487 ( .A(n66315), .B(n68652), .Z(n63274) );
  IV U83488 ( .A(n63274), .Z(n63275) );
  NOR U83489 ( .A(n68655), .B(n63275), .Z(n63276) );
  XOR U83490 ( .A(n66316), .B(n63276), .Z(n76636) );
  IV U83491 ( .A(n63277), .Z(n63279) );
  NOR U83492 ( .A(n63279), .B(n63278), .Z(n76642) );
  NOR U83493 ( .A(n76634), .B(n76642), .Z(n68658) );
  XOR U83494 ( .A(n76636), .B(n68658), .Z(n63280) );
  IV U83495 ( .A(n63280), .Z(n68660) );
  XOR U83496 ( .A(n68659), .B(n68660), .Z(n66313) );
  IV U83497 ( .A(n63281), .Z(n63282) );
  NOR U83498 ( .A(n63283), .B(n63282), .Z(n66312) );
  IV U83499 ( .A(n63284), .Z(n63285) );
  NOR U83500 ( .A(n63286), .B(n63285), .Z(n66306) );
  NOR U83501 ( .A(n66312), .B(n66306), .Z(n63287) );
  XOR U83502 ( .A(n66313), .B(n63287), .Z(n66308) );
  XOR U83503 ( .A(n66309), .B(n66308), .Z(n63296) );
  IV U83504 ( .A(n63296), .Z(n68666) );
  XOR U83505 ( .A(n66304), .B(n68666), .Z(n63288) );
  NOR U83506 ( .A(n63289), .B(n63288), .Z(n71258) );
  IV U83507 ( .A(n63290), .Z(n63291) );
  NOR U83508 ( .A(n63291), .B(n63294), .Z(n63292) );
  IV U83509 ( .A(n63292), .Z(n68669) );
  IV U83510 ( .A(n63293), .Z(n63295) );
  NOR U83511 ( .A(n63295), .B(n63294), .Z(n68665) );
  NOR U83512 ( .A(n66304), .B(n68665), .Z(n63297) );
  XOR U83513 ( .A(n63297), .B(n63296), .Z(n68668) );
  XOR U83514 ( .A(n68669), .B(n68668), .Z(n63298) );
  NOR U83515 ( .A(n63299), .B(n63298), .Z(n63300) );
  NOR U83516 ( .A(n71258), .B(n63300), .Z(n66302) );
  IV U83517 ( .A(n63301), .Z(n63303) );
  NOR U83518 ( .A(n63303), .B(n63302), .Z(n66303) );
  IV U83519 ( .A(n63304), .Z(n63306) );
  NOR U83520 ( .A(n63306), .B(n63305), .Z(n68677) );
  NOR U83521 ( .A(n66303), .B(n68677), .Z(n63307) );
  XOR U83522 ( .A(n66302), .B(n63307), .Z(n68689) );
  IV U83523 ( .A(n63308), .Z(n63309) );
  NOR U83524 ( .A(n63310), .B(n63309), .Z(n68685) );
  IV U83525 ( .A(n63311), .Z(n63313) );
  NOR U83526 ( .A(n63313), .B(n63312), .Z(n68688) );
  NOR U83527 ( .A(n68685), .B(n68688), .Z(n63314) );
  XOR U83528 ( .A(n68689), .B(n63314), .Z(n68696) );
  XOR U83529 ( .A(n63315), .B(n68696), .Z(n66300) );
  XOR U83530 ( .A(n63316), .B(n66300), .Z(n66292) );
  IV U83531 ( .A(n63317), .Z(n63319) );
  NOR U83532 ( .A(n63319), .B(n63318), .Z(n66295) );
  IV U83533 ( .A(n63320), .Z(n63321) );
  NOR U83534 ( .A(n63322), .B(n63321), .Z(n66293) );
  NOR U83535 ( .A(n66295), .B(n66293), .Z(n63323) );
  XOR U83536 ( .A(n66292), .B(n63323), .Z(n66291) );
  XOR U83537 ( .A(n66289), .B(n66291), .Z(n66284) );
  XOR U83538 ( .A(n66283), .B(n66284), .Z(n66287) );
  XOR U83539 ( .A(n63324), .B(n66287), .Z(n66273) );
  XOR U83540 ( .A(n63325), .B(n66273), .Z(n68709) );
  XOR U83541 ( .A(n63326), .B(n68709), .Z(n63327) );
  IV U83542 ( .A(n63327), .Z(n68714) );
  XOR U83543 ( .A(n63328), .B(n68714), .Z(n63334) );
  IV U83544 ( .A(n63334), .Z(n66261) );
  NOR U83545 ( .A(n63329), .B(n66261), .Z(n73679) );
  IV U83546 ( .A(n63330), .Z(n63331) );
  NOR U83547 ( .A(n63331), .B(n66263), .Z(n63339) );
  IV U83548 ( .A(n63332), .Z(n63333) );
  NOR U83549 ( .A(n63333), .B(n66263), .Z(n63335) );
  NOR U83550 ( .A(n63335), .B(n63334), .Z(n63337) );
  IV U83551 ( .A(n63335), .Z(n63336) );
  NOR U83552 ( .A(n68714), .B(n63336), .Z(n73671) );
  NOR U83553 ( .A(n63337), .B(n73671), .Z(n63338) );
  XOR U83554 ( .A(n63339), .B(n63338), .Z(n63340) );
  NOR U83555 ( .A(n63341), .B(n63340), .Z(n63342) );
  NOR U83556 ( .A(n73679), .B(n63342), .Z(n68716) );
  IV U83557 ( .A(n63343), .Z(n63345) );
  NOR U83558 ( .A(n63345), .B(n63344), .Z(n63346) );
  IV U83559 ( .A(n63346), .Z(n68717) );
  XOR U83560 ( .A(n68716), .B(n68717), .Z(n71213) );
  XOR U83561 ( .A(n68720), .B(n71213), .Z(n63353) );
  XOR U83562 ( .A(n68722), .B(n63353), .Z(n63347) );
  NOR U83563 ( .A(n63348), .B(n63347), .Z(n71203) );
  IV U83564 ( .A(n63349), .Z(n63351) );
  NOR U83565 ( .A(n63351), .B(n63350), .Z(n66258) );
  NOR U83566 ( .A(n63352), .B(n66258), .Z(n63354) );
  IV U83567 ( .A(n63353), .Z(n68721) );
  XOR U83568 ( .A(n63354), .B(n68721), .Z(n63355) );
  NOR U83569 ( .A(n63356), .B(n63355), .Z(n63357) );
  NOR U83570 ( .A(n71203), .B(n63357), .Z(n63358) );
  IV U83571 ( .A(n63358), .Z(n68726) );
  NOR U83572 ( .A(n63364), .B(n68726), .Z(n71198) );
  NOR U83573 ( .A(n63360), .B(n63359), .Z(n66254) );
  IV U83574 ( .A(n63361), .Z(n63363) );
  NOR U83575 ( .A(n63363), .B(n63362), .Z(n68725) );
  XOR U83576 ( .A(n68725), .B(n68726), .Z(n66255) );
  IV U83577 ( .A(n66255), .Z(n63365) );
  XOR U83578 ( .A(n66254), .B(n63365), .Z(n63367) );
  NOR U83579 ( .A(n63365), .B(n63364), .Z(n63366) );
  NOR U83580 ( .A(n63367), .B(n63366), .Z(n63368) );
  NOR U83581 ( .A(n71198), .B(n63368), .Z(n63369) );
  IV U83582 ( .A(n63369), .Z(n68732) );
  XOR U83583 ( .A(n66253), .B(n68732), .Z(n63378) );
  IV U83584 ( .A(n63372), .Z(n63370) );
  NOR U83585 ( .A(n63371), .B(n63370), .Z(n68735) );
  NOR U83586 ( .A(n63373), .B(n63372), .Z(n63376) );
  IV U83587 ( .A(n63374), .Z(n63375) );
  NOR U83588 ( .A(n63376), .B(n63375), .Z(n68730) );
  NOR U83589 ( .A(n68735), .B(n68730), .Z(n63377) );
  XOR U83590 ( .A(n63378), .B(n63377), .Z(n68739) );
  XOR U83591 ( .A(n63379), .B(n68739), .Z(n68745) );
  XOR U83592 ( .A(n63380), .B(n68745), .Z(n73711) );
  XOR U83593 ( .A(n66246), .B(n73711), .Z(n66242) );
  IV U83594 ( .A(n63381), .Z(n63382) );
  NOR U83595 ( .A(n63383), .B(n63382), .Z(n66241) );
  NOR U83596 ( .A(n63384), .B(n68753), .Z(n63385) );
  NOR U83597 ( .A(n66241), .B(n63385), .Z(n63386) );
  XOR U83598 ( .A(n66242), .B(n63386), .Z(n68773) );
  IV U83599 ( .A(n63387), .Z(n68760) );
  NOR U83600 ( .A(n63388), .B(n68760), .Z(n63392) );
  IV U83601 ( .A(n63389), .Z(n63391) );
  NOR U83602 ( .A(n63391), .B(n63390), .Z(n68771) );
  NOR U83603 ( .A(n63392), .B(n68771), .Z(n63393) );
  XOR U83604 ( .A(n68773), .B(n63393), .Z(n66239) );
  NOR U83605 ( .A(n63394), .B(n68768), .Z(n63398) );
  IV U83606 ( .A(n63395), .Z(n63396) );
  NOR U83607 ( .A(n63397), .B(n63396), .Z(n66238) );
  NOR U83608 ( .A(n63398), .B(n66238), .Z(n63399) );
  XOR U83609 ( .A(n66239), .B(n63399), .Z(n68781) );
  IV U83610 ( .A(n68781), .Z(n63410) );
  IV U83611 ( .A(n63400), .Z(n63416) );
  IV U83612 ( .A(n63401), .Z(n63402) );
  NOR U83613 ( .A(n63416), .B(n63402), .Z(n68779) );
  IV U83614 ( .A(n63403), .Z(n63404) );
  NOR U83615 ( .A(n63404), .B(n63406), .Z(n66234) );
  IV U83616 ( .A(n63405), .Z(n63407) );
  NOR U83617 ( .A(n63407), .B(n63406), .Z(n66235) );
  XOR U83618 ( .A(n66234), .B(n66235), .Z(n63408) );
  NOR U83619 ( .A(n68779), .B(n63408), .Z(n63409) );
  XOR U83620 ( .A(n63410), .B(n63409), .Z(n68784) );
  IV U83621 ( .A(n63411), .Z(n63412) );
  NOR U83622 ( .A(n63413), .B(n63412), .Z(n66231) );
  IV U83623 ( .A(n63414), .Z(n63415) );
  NOR U83624 ( .A(n63416), .B(n63415), .Z(n68782) );
  NOR U83625 ( .A(n66231), .B(n68782), .Z(n63417) );
  XOR U83626 ( .A(n68784), .B(n63417), .Z(n66228) );
  IV U83627 ( .A(n63418), .Z(n63420) );
  NOR U83628 ( .A(n63420), .B(n63419), .Z(n66229) );
  IV U83629 ( .A(n63421), .Z(n63423) );
  NOR U83630 ( .A(n63423), .B(n63422), .Z(n68785) );
  NOR U83631 ( .A(n66229), .B(n68785), .Z(n63424) );
  XOR U83632 ( .A(n66228), .B(n63424), .Z(n66225) );
  XOR U83633 ( .A(n66224), .B(n66225), .Z(n68789) );
  IV U83634 ( .A(n63425), .Z(n63426) );
  NOR U83635 ( .A(n63427), .B(n63426), .Z(n66221) );
  NOR U83636 ( .A(n68788), .B(n66221), .Z(n63428) );
  XOR U83637 ( .A(n68789), .B(n63428), .Z(n66217) );
  NOR U83638 ( .A(n63429), .B(n66218), .Z(n63433) );
  IV U83639 ( .A(n63430), .Z(n63432) );
  NOR U83640 ( .A(n63432), .B(n63431), .Z(n68802) );
  NOR U83641 ( .A(n63433), .B(n68802), .Z(n63434) );
  XOR U83642 ( .A(n66217), .B(n63434), .Z(n68800) );
  XOR U83643 ( .A(n63435), .B(n68800), .Z(n66203) );
  XOR U83644 ( .A(n63436), .B(n66203), .Z(n66194) );
  IV U83645 ( .A(n63437), .Z(n63439) );
  NOR U83646 ( .A(n63439), .B(n63438), .Z(n66207) );
  NOR U83647 ( .A(n63440), .B(n66195), .Z(n63441) );
  NOR U83648 ( .A(n66207), .B(n63441), .Z(n63442) );
  XOR U83649 ( .A(n66194), .B(n63442), .Z(n68809) );
  IV U83650 ( .A(n63443), .Z(n63446) );
  NOR U83651 ( .A(n63444), .B(n66187), .Z(n63445) );
  IV U83652 ( .A(n63445), .Z(n63448) );
  NOR U83653 ( .A(n63446), .B(n63448), .Z(n68807) );
  XOR U83654 ( .A(n68809), .B(n68807), .Z(n68812) );
  IV U83655 ( .A(n63447), .Z(n63449) );
  NOR U83656 ( .A(n63449), .B(n63448), .Z(n68810) );
  IV U83657 ( .A(n63450), .Z(n63451) );
  NOR U83658 ( .A(n66187), .B(n63451), .Z(n63452) );
  NOR U83659 ( .A(n68810), .B(n63452), .Z(n63453) );
  XOR U83660 ( .A(n68812), .B(n63453), .Z(n66181) );
  IV U83661 ( .A(n63454), .Z(n63456) );
  NOR U83662 ( .A(n63456), .B(n63455), .Z(n63457) );
  IV U83663 ( .A(n63457), .Z(n66182) );
  XOR U83664 ( .A(n66181), .B(n66182), .Z(n68820) );
  XOR U83665 ( .A(n63458), .B(n68820), .Z(n66178) );
  XOR U83666 ( .A(n63459), .B(n66178), .Z(n66177) );
  XOR U83667 ( .A(n66176), .B(n66177), .Z(n63466) );
  IV U83668 ( .A(n63466), .Z(n63460) );
  NOR U83669 ( .A(n63461), .B(n63460), .Z(n63462) );
  IV U83670 ( .A(n63462), .Z(n63463) );
  NOR U83671 ( .A(n63464), .B(n63463), .Z(n73794) );
  NOR U83672 ( .A(n63465), .B(n63464), .Z(n63467) );
  NOR U83673 ( .A(n63467), .B(n63466), .Z(n63468) );
  NOR U83674 ( .A(n73794), .B(n63468), .Z(n63473) );
  IV U83675 ( .A(n63473), .Z(n68834) );
  XOR U83676 ( .A(n68830), .B(n68834), .Z(n63469) );
  NOR U83677 ( .A(n63470), .B(n63469), .Z(n73802) );
  NOR U83678 ( .A(n63472), .B(n63471), .Z(n68836) );
  NOR U83679 ( .A(n68830), .B(n68833), .Z(n63474) );
  XOR U83680 ( .A(n63474), .B(n63473), .Z(n68837) );
  XOR U83681 ( .A(n68836), .B(n68837), .Z(n66174) );
  IV U83682 ( .A(n66174), .Z(n63475) );
  NOR U83683 ( .A(n63476), .B(n63475), .Z(n63477) );
  NOR U83684 ( .A(n73802), .B(n63477), .Z(n68841) );
  IV U83685 ( .A(n63478), .Z(n63479) );
  NOR U83686 ( .A(n63480), .B(n63479), .Z(n68840) );
  IV U83687 ( .A(n63481), .Z(n63483) );
  NOR U83688 ( .A(n63483), .B(n63482), .Z(n66173) );
  NOR U83689 ( .A(n68840), .B(n66173), .Z(n63484) );
  XOR U83690 ( .A(n68841), .B(n63484), .Z(n68846) );
  IV U83691 ( .A(n63485), .Z(n63487) );
  NOR U83692 ( .A(n63487), .B(n63486), .Z(n66171) );
  IV U83693 ( .A(n63488), .Z(n63489) );
  NOR U83694 ( .A(n63490), .B(n63489), .Z(n68844) );
  NOR U83695 ( .A(n66171), .B(n68844), .Z(n63491) );
  XOR U83696 ( .A(n68846), .B(n63491), .Z(n63492) );
  IV U83697 ( .A(n63492), .Z(n68848) );
  XOR U83698 ( .A(n68847), .B(n68848), .Z(n68856) );
  IV U83699 ( .A(n63493), .Z(n63494) );
  NOR U83700 ( .A(n63495), .B(n63494), .Z(n68851) );
  NOR U83701 ( .A(n68857), .B(n68851), .Z(n63496) );
  XOR U83702 ( .A(n68856), .B(n63496), .Z(n68861) );
  XOR U83703 ( .A(n63497), .B(n68861), .Z(n73837) );
  XOR U83704 ( .A(n66166), .B(n73837), .Z(n66168) );
  IV U83705 ( .A(n63498), .Z(n63499) );
  NOR U83706 ( .A(n71105), .B(n63499), .Z(n63503) );
  IV U83707 ( .A(n63500), .Z(n63502) );
  NOR U83708 ( .A(n63502), .B(n63501), .Z(n73832) );
  NOR U83709 ( .A(n63503), .B(n73832), .Z(n66169) );
  XOR U83710 ( .A(n66168), .B(n66169), .Z(n63509) );
  IV U83711 ( .A(n63509), .Z(n63504) );
  NOR U83712 ( .A(n63505), .B(n63504), .Z(n63506) );
  IV U83713 ( .A(n63506), .Z(n66164) );
  NOR U83714 ( .A(n63508), .B(n66164), .Z(n73840) );
  NOR U83715 ( .A(n63508), .B(n63507), .Z(n63510) );
  NOR U83716 ( .A(n63510), .B(n63509), .Z(n63511) );
  NOR U83717 ( .A(n73840), .B(n63511), .Z(n66160) );
  XOR U83718 ( .A(n63512), .B(n66160), .Z(n68867) );
  XOR U83719 ( .A(n63513), .B(n68867), .Z(n63514) );
  IV U83720 ( .A(n63514), .Z(n68877) );
  XOR U83721 ( .A(n68874), .B(n68877), .Z(n66149) );
  XOR U83722 ( .A(n63515), .B(n66149), .Z(n66144) );
  XOR U83723 ( .A(n66145), .B(n66144), .Z(n73857) );
  XOR U83724 ( .A(n73859), .B(n73857), .Z(n63516) );
  IV U83725 ( .A(n63516), .Z(n66139) );
  XOR U83726 ( .A(n66138), .B(n66139), .Z(n66142) );
  XOR U83727 ( .A(n66141), .B(n66142), .Z(n66137) );
  IV U83728 ( .A(n63517), .Z(n63522) );
  NOR U83729 ( .A(n63519), .B(n63518), .Z(n63520) );
  IV U83730 ( .A(n63520), .Z(n63521) );
  NOR U83731 ( .A(n63522), .B(n63521), .Z(n66135) );
  XOR U83732 ( .A(n66137), .B(n66135), .Z(n68884) );
  XOR U83733 ( .A(n68883), .B(n68884), .Z(n68894) );
  XOR U83734 ( .A(n66133), .B(n68894), .Z(n68891) );
  XOR U83735 ( .A(n68890), .B(n68891), .Z(n66131) );
  IV U83736 ( .A(n63523), .Z(n68895) );
  NOR U83737 ( .A(n63524), .B(n68895), .Z(n63528) );
  IV U83738 ( .A(n63525), .Z(n63527) );
  NOR U83739 ( .A(n63527), .B(n63526), .Z(n66130) );
  NOR U83740 ( .A(n63528), .B(n66130), .Z(n63529) );
  XOR U83741 ( .A(n66131), .B(n63529), .Z(n63530) );
  IV U83742 ( .A(n63530), .Z(n66126) );
  IV U83743 ( .A(n63531), .Z(n63533) );
  NOR U83744 ( .A(n63533), .B(n63532), .Z(n63538) );
  IV U83745 ( .A(n63538), .Z(n63534) );
  NOR U83746 ( .A(n66126), .B(n63534), .Z(n73893) );
  NOR U83747 ( .A(n63536), .B(n63535), .Z(n66127) );
  XOR U83748 ( .A(n66124), .B(n66126), .Z(n66128) );
  XOR U83749 ( .A(n66127), .B(n66128), .Z(n68904) );
  IV U83750 ( .A(n68904), .Z(n63537) );
  NOR U83751 ( .A(n63538), .B(n63537), .Z(n63539) );
  NOR U83752 ( .A(n73893), .B(n63539), .Z(n68907) );
  XOR U83753 ( .A(n63540), .B(n68907), .Z(n82040) );
  XOR U83754 ( .A(n68906), .B(n82040), .Z(n63544) );
  XOR U83755 ( .A(n66121), .B(n63544), .Z(n66122) );
  XOR U83756 ( .A(n66123), .B(n66122), .Z(n63541) );
  NOR U83757 ( .A(n63542), .B(n63541), .Z(n63553) );
  IV U83758 ( .A(n63543), .Z(n63547) );
  IV U83759 ( .A(n63544), .Z(n66120) );
  NOR U83760 ( .A(n63545), .B(n66120), .Z(n63546) );
  IV U83761 ( .A(n63546), .Z(n63549) );
  NOR U83762 ( .A(n63547), .B(n63549), .Z(n82026) );
  IV U83763 ( .A(n63548), .Z(n63550) );
  NOR U83764 ( .A(n63550), .B(n63549), .Z(n73901) );
  NOR U83765 ( .A(n82026), .B(n73901), .Z(n63551) );
  IV U83766 ( .A(n63551), .Z(n63552) );
  NOR U83767 ( .A(n63553), .B(n63552), .Z(n68913) );
  XOR U83768 ( .A(n73907), .B(n68913), .Z(n66118) );
  IV U83769 ( .A(n63554), .Z(n63555) );
  NOR U83770 ( .A(n63556), .B(n63555), .Z(n66117) );
  IV U83771 ( .A(n63557), .Z(n71076) );
  NOR U83772 ( .A(n71076), .B(n68916), .Z(n63558) );
  NOR U83773 ( .A(n66117), .B(n63558), .Z(n63559) );
  XOR U83774 ( .A(n66118), .B(n63559), .Z(n63560) );
  IV U83775 ( .A(n63560), .Z(n66116) );
  XOR U83776 ( .A(n66114), .B(n66116), .Z(n66110) );
  IV U83777 ( .A(n63561), .Z(n63562) );
  NOR U83778 ( .A(n63563), .B(n63562), .Z(n66112) );
  IV U83779 ( .A(n63564), .Z(n63565) );
  NOR U83780 ( .A(n63566), .B(n63565), .Z(n66109) );
  NOR U83781 ( .A(n66112), .B(n66109), .Z(n63567) );
  XOR U83782 ( .A(n66110), .B(n63567), .Z(n66099) );
  XOR U83783 ( .A(n63568), .B(n66099), .Z(n66103) );
  XOR U83784 ( .A(n66102), .B(n66103), .Z(n66098) );
  XOR U83785 ( .A(n63569), .B(n66098), .Z(n68923) );
  IV U83786 ( .A(n63570), .Z(n68927) );
  NOR U83787 ( .A(n63571), .B(n68927), .Z(n63574) );
  IV U83788 ( .A(n63572), .Z(n63573) );
  NOR U83789 ( .A(n63573), .B(n63577), .Z(n68928) );
  NOR U83790 ( .A(n63574), .B(n68928), .Z(n63575) );
  XOR U83791 ( .A(n68923), .B(n63575), .Z(n68933) );
  IV U83792 ( .A(n63576), .Z(n63578) );
  NOR U83793 ( .A(n63578), .B(n63577), .Z(n68931) );
  XOR U83794 ( .A(n68933), .B(n68931), .Z(n68935) );
  NOR U83795 ( .A(n63585), .B(n68935), .Z(n66093) );
  IV U83796 ( .A(n63579), .Z(n63581) );
  NOR U83797 ( .A(n63581), .B(n63580), .Z(n66090) );
  IV U83798 ( .A(n63582), .Z(n63583) );
  NOR U83799 ( .A(n63584), .B(n63583), .Z(n68934) );
  XOR U83800 ( .A(n68934), .B(n68935), .Z(n66091) );
  IV U83801 ( .A(n66091), .Z(n63586) );
  XOR U83802 ( .A(n66090), .B(n63586), .Z(n63588) );
  NOR U83803 ( .A(n63586), .B(n63585), .Z(n63587) );
  NOR U83804 ( .A(n63588), .B(n63587), .Z(n63589) );
  NOR U83805 ( .A(n66093), .B(n63589), .Z(n63590) );
  IV U83806 ( .A(n63590), .Z(n66088) );
  XOR U83807 ( .A(n66089), .B(n66088), .Z(n63591) );
  XOR U83808 ( .A(n63592), .B(n63591), .Z(n66078) );
  NOR U83809 ( .A(n63593), .B(n66077), .Z(n66065) );
  IV U83810 ( .A(n63594), .Z(n66070) );
  NOR U83811 ( .A(n63595), .B(n66070), .Z(n63596) );
  NOR U83812 ( .A(n66065), .B(n63596), .Z(n63597) );
  XOR U83813 ( .A(n66078), .B(n63597), .Z(n66062) );
  IV U83814 ( .A(n63598), .Z(n63599) );
  NOR U83815 ( .A(n63600), .B(n63599), .Z(n66066) );
  IV U83816 ( .A(n63601), .Z(n63602) );
  NOR U83817 ( .A(n63603), .B(n63602), .Z(n66061) );
  NOR U83818 ( .A(n66066), .B(n66061), .Z(n63604) );
  XOR U83819 ( .A(n66062), .B(n63604), .Z(n66055) );
  XOR U83820 ( .A(n63605), .B(n66055), .Z(n66045) );
  XOR U83821 ( .A(n63606), .B(n66045), .Z(n63615) );
  IV U83822 ( .A(n63615), .Z(n63607) );
  NOR U83823 ( .A(n63608), .B(n63607), .Z(n81943) );
  XOR U83824 ( .A(n63609), .B(n66045), .Z(n63614) );
  IV U83825 ( .A(n63610), .Z(n63611) );
  NOR U83826 ( .A(n63612), .B(n63611), .Z(n63616) );
  IV U83827 ( .A(n63616), .Z(n63613) );
  NOR U83828 ( .A(n63614), .B(n63613), .Z(n73968) );
  NOR U83829 ( .A(n63616), .B(n63615), .Z(n63617) );
  NOR U83830 ( .A(n73968), .B(n63617), .Z(n63618) );
  NOR U83831 ( .A(n63619), .B(n63618), .Z(n63620) );
  NOR U83832 ( .A(n81943), .B(n63620), .Z(n66040) );
  IV U83833 ( .A(n63621), .Z(n63623) );
  NOR U83834 ( .A(n63623), .B(n63622), .Z(n68937) );
  IV U83835 ( .A(n63624), .Z(n63626) );
  NOR U83836 ( .A(n63626), .B(n63625), .Z(n66041) );
  NOR U83837 ( .A(n68937), .B(n66041), .Z(n63627) );
  XOR U83838 ( .A(n66040), .B(n63627), .Z(n68941) );
  XOR U83839 ( .A(n63628), .B(n68941), .Z(n63641) );
  XOR U83840 ( .A(n66036), .B(n63641), .Z(n63639) );
  IV U83841 ( .A(n63639), .Z(n63637) );
  IV U83842 ( .A(n63629), .Z(n63631) );
  NOR U83843 ( .A(n63631), .B(n63630), .Z(n63638) );
  IV U83844 ( .A(n63632), .Z(n63633) );
  NOR U83845 ( .A(n63634), .B(n63633), .Z(n63642) );
  NOR U83846 ( .A(n63638), .B(n63642), .Z(n63635) );
  IV U83847 ( .A(n63635), .Z(n63636) );
  NOR U83848 ( .A(n63637), .B(n63636), .Z(n63645) );
  IV U83849 ( .A(n63638), .Z(n63640) );
  NOR U83850 ( .A(n63640), .B(n63639), .Z(n73988) );
  IV U83851 ( .A(n63641), .Z(n66037) );
  IV U83852 ( .A(n63642), .Z(n63643) );
  NOR U83853 ( .A(n66037), .B(n63643), .Z(n71011) );
  NOR U83854 ( .A(n73988), .B(n71011), .Z(n63644) );
  IV U83855 ( .A(n63644), .Z(n66035) );
  NOR U83856 ( .A(n63645), .B(n66035), .Z(n66029) );
  IV U83857 ( .A(n63646), .Z(n66030) );
  NOR U83858 ( .A(n66030), .B(n90897), .Z(n63648) );
  IV U83859 ( .A(n90898), .Z(n63647) );
  NOR U83860 ( .A(n63647), .B(n90897), .Z(n66032) );
  NOR U83861 ( .A(n63648), .B(n66032), .Z(n63649) );
  XOR U83862 ( .A(n66029), .B(n63649), .Z(n68956) );
  XOR U83863 ( .A(n68954), .B(n68956), .Z(n66027) );
  XOR U83864 ( .A(n63650), .B(n66027), .Z(n63653) );
  XOR U83865 ( .A(n63651), .B(n63653), .Z(n63660) );
  NOR U83866 ( .A(n63652), .B(n63660), .Z(n70998) );
  IV U83867 ( .A(n63653), .Z(n66020) );
  XOR U83868 ( .A(n63654), .B(n66020), .Z(n63659) );
  IV U83869 ( .A(n63655), .Z(n63656) );
  NOR U83870 ( .A(n63657), .B(n63656), .Z(n63662) );
  IV U83871 ( .A(n63662), .Z(n63658) );
  NOR U83872 ( .A(n63659), .B(n63658), .Z(n74019) );
  IV U83873 ( .A(n63660), .Z(n63661) );
  NOR U83874 ( .A(n63662), .B(n63661), .Z(n63663) );
  NOR U83875 ( .A(n74019), .B(n63663), .Z(n63667) );
  NOR U83876 ( .A(n63664), .B(n63667), .Z(n63665) );
  NOR U83877 ( .A(n70998), .B(n63665), .Z(n66009) );
  NOR U83878 ( .A(n63666), .B(n66009), .Z(n63670) );
  IV U83879 ( .A(n63666), .Z(n63669) );
  IV U83880 ( .A(n63667), .Z(n63668) );
  NOR U83881 ( .A(n63669), .B(n63668), .Z(n71001) );
  NOR U83882 ( .A(n63670), .B(n71001), .Z(n63671) );
  IV U83883 ( .A(n63671), .Z(n66015) );
  IV U83884 ( .A(n63672), .Z(n63673) );
  NOR U83885 ( .A(n63674), .B(n63673), .Z(n66013) );
  XOR U83886 ( .A(n66015), .B(n66013), .Z(n68972) );
  XOR U83887 ( .A(n63675), .B(n68972), .Z(n68974) );
  XOR U83888 ( .A(n68975), .B(n68974), .Z(n68977) );
  XOR U83889 ( .A(n68976), .B(n68977), .Z(n66005) );
  IV U83890 ( .A(n66005), .Z(n63683) );
  IV U83891 ( .A(n63676), .Z(n63678) );
  NOR U83892 ( .A(n63678), .B(n63677), .Z(n68980) );
  IV U83893 ( .A(n63679), .Z(n63681) );
  NOR U83894 ( .A(n63681), .B(n63680), .Z(n66004) );
  NOR U83895 ( .A(n68980), .B(n66004), .Z(n63682) );
  XOR U83896 ( .A(n63683), .B(n63682), .Z(n66003) );
  XOR U83897 ( .A(n66001), .B(n66003), .Z(n68988) );
  XOR U83898 ( .A(n63684), .B(n68988), .Z(n68990) );
  IV U83899 ( .A(n63685), .Z(n63686) );
  NOR U83900 ( .A(n63687), .B(n63686), .Z(n68991) );
  IV U83901 ( .A(n63688), .Z(n63689) );
  NOR U83902 ( .A(n63690), .B(n63689), .Z(n68994) );
  NOR U83903 ( .A(n68991), .B(n68994), .Z(n63691) );
  XOR U83904 ( .A(n68990), .B(n63691), .Z(n70962) );
  XOR U83905 ( .A(n69001), .B(n70962), .Z(n65997) );
  XOR U83906 ( .A(n65996), .B(n65997), .Z(n65993) );
  IV U83907 ( .A(n63692), .Z(n63693) );
  NOR U83908 ( .A(n63693), .B(n63695), .Z(n68998) );
  IV U83909 ( .A(n63694), .Z(n63696) );
  NOR U83910 ( .A(n63696), .B(n63695), .Z(n65994) );
  NOR U83911 ( .A(n68998), .B(n65994), .Z(n63697) );
  XOR U83912 ( .A(n65993), .B(n63697), .Z(n65986) );
  NOR U83913 ( .A(n63698), .B(n65987), .Z(n63699) );
  XOR U83914 ( .A(n65986), .B(n63699), .Z(n65984) );
  XOR U83915 ( .A(n63700), .B(n65984), .Z(n65975) );
  IV U83916 ( .A(n63701), .Z(n63702) );
  NOR U83917 ( .A(n63703), .B(n63702), .Z(n65977) );
  IV U83918 ( .A(n63704), .Z(n63705) );
  NOR U83919 ( .A(n63706), .B(n63705), .Z(n65974) );
  NOR U83920 ( .A(n65977), .B(n65974), .Z(n63707) );
  XOR U83921 ( .A(n65975), .B(n63707), .Z(n65970) );
  XOR U83922 ( .A(n63708), .B(n65970), .Z(n65965) );
  XOR U83923 ( .A(n63709), .B(n65965), .Z(n79418) );
  IV U83924 ( .A(n63710), .Z(n63711) );
  NOR U83925 ( .A(n79420), .B(n63711), .Z(n65961) );
  IV U83926 ( .A(n63712), .Z(n79427) );
  NOR U83927 ( .A(n63713), .B(n79427), .Z(n65957) );
  NOR U83928 ( .A(n65961), .B(n65957), .Z(n63714) );
  XOR U83929 ( .A(n79418), .B(n63714), .Z(n65955) );
  IV U83930 ( .A(n63715), .Z(n63716) );
  NOR U83931 ( .A(n63717), .B(n63716), .Z(n65954) );
  IV U83932 ( .A(n63718), .Z(n63719) );
  NOR U83933 ( .A(n63720), .B(n63719), .Z(n65952) );
  NOR U83934 ( .A(n65954), .B(n65952), .Z(n63721) );
  XOR U83935 ( .A(n65955), .B(n63721), .Z(n63722) );
  NOR U83936 ( .A(n63723), .B(n63722), .Z(n63726) );
  IV U83937 ( .A(n63723), .Z(n63725) );
  XOR U83938 ( .A(n65954), .B(n65955), .Z(n63724) );
  NOR U83939 ( .A(n63725), .B(n63724), .Z(n70930) );
  NOR U83940 ( .A(n63726), .B(n70930), .Z(n65949) );
  IV U83941 ( .A(n63727), .Z(n63729) );
  NOR U83942 ( .A(n63729), .B(n63728), .Z(n63730) );
  IV U83943 ( .A(n63730), .Z(n65950) );
  XOR U83944 ( .A(n65949), .B(n65950), .Z(n65945) );
  XOR U83945 ( .A(n65944), .B(n65945), .Z(n65947) );
  XOR U83946 ( .A(n65948), .B(n65947), .Z(n65936) );
  NOR U83947 ( .A(n63731), .B(n65941), .Z(n63735) );
  IV U83948 ( .A(n63732), .Z(n63733) );
  NOR U83949 ( .A(n63734), .B(n63733), .Z(n65935) );
  NOR U83950 ( .A(n63735), .B(n65935), .Z(n63736) );
  XOR U83951 ( .A(n65936), .B(n63736), .Z(n69024) );
  XOR U83952 ( .A(n69022), .B(n69024), .Z(n69026) );
  XOR U83953 ( .A(n69025), .B(n69026), .Z(n65927) );
  IV U83954 ( .A(n63737), .Z(n65929) );
  NOR U83955 ( .A(n63738), .B(n65929), .Z(n63744) );
  IV U83956 ( .A(n63739), .Z(n63740) );
  NOR U83957 ( .A(n65932), .B(n63740), .Z(n65933) );
  IV U83958 ( .A(n63741), .Z(n63742) );
  NOR U83959 ( .A(n65932), .B(n63742), .Z(n65926) );
  NOR U83960 ( .A(n65933), .B(n65926), .Z(n63743) );
  XOR U83961 ( .A(n63744), .B(n63743), .Z(n63745) );
  XOR U83962 ( .A(n65927), .B(n63745), .Z(n65917) );
  IV U83963 ( .A(n63746), .Z(n63747) );
  NOR U83964 ( .A(n63750), .B(n63747), .Z(n65923) );
  IV U83965 ( .A(n63748), .Z(n63749) );
  NOR U83966 ( .A(n63750), .B(n63749), .Z(n65918) );
  NOR U83967 ( .A(n65923), .B(n65918), .Z(n63751) );
  XOR U83968 ( .A(n65917), .B(n63751), .Z(n65921) );
  XOR U83969 ( .A(n65920), .B(n65921), .Z(n69033) );
  XOR U83970 ( .A(n69030), .B(n69033), .Z(n69037) );
  IV U83971 ( .A(n63752), .Z(n63753) );
  NOR U83972 ( .A(n63754), .B(n63753), .Z(n69032) );
  IV U83973 ( .A(n63755), .Z(n63756) );
  NOR U83974 ( .A(n63757), .B(n63756), .Z(n69036) );
  NOR U83975 ( .A(n69032), .B(n69036), .Z(n63758) );
  XOR U83976 ( .A(n69037), .B(n63758), .Z(n65911) );
  IV U83977 ( .A(n63759), .Z(n63761) );
  NOR U83978 ( .A(n63761), .B(n63760), .Z(n65914) );
  IV U83979 ( .A(n63762), .Z(n63764) );
  NOR U83980 ( .A(n63764), .B(n63763), .Z(n65912) );
  NOR U83981 ( .A(n65914), .B(n65912), .Z(n63765) );
  XOR U83982 ( .A(n65911), .B(n63765), .Z(n65907) );
  XOR U83983 ( .A(n65906), .B(n65907), .Z(n69041) );
  IV U83984 ( .A(n63766), .Z(n63768) );
  NOR U83985 ( .A(n63768), .B(n63767), .Z(n65909) );
  IV U83986 ( .A(n63769), .Z(n63771) );
  NOR U83987 ( .A(n63771), .B(n63770), .Z(n69039) );
  NOR U83988 ( .A(n65909), .B(n69039), .Z(n63772) );
  XOR U83989 ( .A(n69041), .B(n63772), .Z(n69043) );
  XOR U83990 ( .A(n63773), .B(n69043), .Z(n65902) );
  XOR U83991 ( .A(n63774), .B(n65902), .Z(n65898) );
  XOR U83992 ( .A(n63775), .B(n65898), .Z(n69052) );
  IV U83993 ( .A(n63776), .Z(n63777) );
  NOR U83994 ( .A(n63778), .B(n63777), .Z(n69050) );
  IV U83995 ( .A(n63779), .Z(n63780) );
  NOR U83996 ( .A(n63781), .B(n63780), .Z(n65893) );
  NOR U83997 ( .A(n69050), .B(n65893), .Z(n63782) );
  XOR U83998 ( .A(n69052), .B(n63782), .Z(n65888) );
  XOR U83999 ( .A(n63783), .B(n65888), .Z(n65884) );
  XOR U84000 ( .A(n65882), .B(n65884), .Z(n70848) );
  XOR U84001 ( .A(n63784), .B(n70848), .Z(n65877) );
  XOR U84002 ( .A(n65876), .B(n65877), .Z(n65880) );
  XOR U84003 ( .A(n63785), .B(n65880), .Z(n65867) );
  IV U84004 ( .A(n63786), .Z(n63788) );
  IV U84005 ( .A(n63787), .Z(n65870) );
  NOR U84006 ( .A(n63788), .B(n65870), .Z(n63789) );
  IV U84007 ( .A(n63789), .Z(n65868) );
  XOR U84008 ( .A(n65867), .B(n65868), .Z(n69056) );
  XOR U84009 ( .A(n69055), .B(n69056), .Z(n69059) );
  XOR U84010 ( .A(n63790), .B(n69059), .Z(n65859) );
  XOR U84011 ( .A(n70832), .B(n65859), .Z(n74102) );
  XOR U84012 ( .A(n74103), .B(n74102), .Z(n69064) );
  IV U84013 ( .A(n69064), .Z(n65853) );
  XOR U84014 ( .A(n65852), .B(n65853), .Z(n65857) );
  XOR U84015 ( .A(n65855), .B(n65857), .Z(n65848) );
  XOR U84016 ( .A(n65846), .B(n65848), .Z(n65851) );
  XOR U84017 ( .A(n63791), .B(n65851), .Z(n65838) );
  XOR U84018 ( .A(n63792), .B(n65838), .Z(n69070) );
  XOR U84019 ( .A(n63793), .B(n69070), .Z(n63794) );
  IV U84020 ( .A(n63794), .Z(n69072) );
  XOR U84021 ( .A(n69071), .B(n69072), .Z(n63799) );
  IV U84022 ( .A(n63795), .Z(n63797) );
  NOR U84023 ( .A(n63797), .B(n63796), .Z(n63804) );
  IV U84024 ( .A(n63804), .Z(n63798) );
  NOR U84025 ( .A(n63799), .B(n63798), .Z(n74120) );
  NOR U84026 ( .A(n63800), .B(n65833), .Z(n63801) );
  NOR U84027 ( .A(n69071), .B(n63801), .Z(n63802) );
  XOR U84028 ( .A(n69072), .B(n63802), .Z(n63803) );
  NOR U84029 ( .A(n63804), .B(n63803), .Z(n63805) );
  NOR U84030 ( .A(n74120), .B(n63805), .Z(n65825) );
  XOR U84031 ( .A(n63806), .B(n65825), .Z(n69083) );
  XOR U84032 ( .A(n69081), .B(n69083), .Z(n69089) );
  IV U84033 ( .A(n63807), .Z(n63809) );
  NOR U84034 ( .A(n63809), .B(n63808), .Z(n69087) );
  XOR U84035 ( .A(n69089), .B(n69087), .Z(n69095) );
  IV U84036 ( .A(n63810), .Z(n63811) );
  NOR U84037 ( .A(n63812), .B(n63811), .Z(n69090) );
  IV U84038 ( .A(n63813), .Z(n63814) );
  NOR U84039 ( .A(n63815), .B(n63814), .Z(n69093) );
  NOR U84040 ( .A(n69090), .B(n69093), .Z(n63816) );
  XOR U84041 ( .A(n69095), .B(n63816), .Z(n65822) );
  XOR U84042 ( .A(n63817), .B(n65822), .Z(n70781) );
  IV U84043 ( .A(n63818), .Z(n63819) );
  NOR U84044 ( .A(n63820), .B(n63819), .Z(n70779) );
  IV U84045 ( .A(n63821), .Z(n63823) );
  NOR U84046 ( .A(n63823), .B(n63822), .Z(n70774) );
  NOR U84047 ( .A(n70779), .B(n70774), .Z(n65816) );
  XOR U84048 ( .A(n70781), .B(n65816), .Z(n65812) );
  XOR U84049 ( .A(n63824), .B(n65812), .Z(n79610) );
  IV U84050 ( .A(n63825), .Z(n63826) );
  NOR U84051 ( .A(n63827), .B(n63826), .Z(n65814) );
  XOR U84052 ( .A(n79610), .B(n65814), .Z(n65806) );
  IV U84053 ( .A(n63828), .Z(n63829) );
  NOR U84054 ( .A(n63830), .B(n63829), .Z(n65805) );
  XOR U84055 ( .A(n65806), .B(n65805), .Z(n65808) );
  XOR U84056 ( .A(n65807), .B(n65808), .Z(n69103) );
  IV U84057 ( .A(n63831), .Z(n63832) );
  NOR U84058 ( .A(n63833), .B(n63832), .Z(n69101) );
  XOR U84059 ( .A(n69103), .B(n69101), .Z(n70754) );
  XOR U84060 ( .A(n63834), .B(n70754), .Z(n65801) );
  XOR U84061 ( .A(n65799), .B(n65801), .Z(n65803) );
  XOR U84062 ( .A(n65802), .B(n65803), .Z(n69109) );
  XOR U84063 ( .A(n69108), .B(n69109), .Z(n69112) );
  XOR U84064 ( .A(n69111), .B(n69112), .Z(n69116) );
  XOR U84065 ( .A(n69115), .B(n69116), .Z(n70745) );
  XOR U84066 ( .A(n69118), .B(n70745), .Z(n65795) );
  IV U84067 ( .A(n63835), .Z(n63837) );
  NOR U84068 ( .A(n63837), .B(n63836), .Z(n69121) );
  IV U84069 ( .A(n63838), .Z(n63839) );
  NOR U84070 ( .A(n63843), .B(n63839), .Z(n65794) );
  NOR U84071 ( .A(n69121), .B(n65794), .Z(n63840) );
  XOR U84072 ( .A(n65795), .B(n63840), .Z(n69125) );
  IV U84073 ( .A(n63841), .Z(n63842) );
  NOR U84074 ( .A(n63843), .B(n63842), .Z(n69123) );
  XOR U84075 ( .A(n69125), .B(n69123), .Z(n69127) );
  XOR U84076 ( .A(n69126), .B(n69127), .Z(n65790) );
  XOR U84077 ( .A(n63844), .B(n65790), .Z(n63845) );
  IV U84078 ( .A(n63845), .Z(n65785) );
  XOR U84079 ( .A(n65783), .B(n65785), .Z(n69132) );
  XOR U84080 ( .A(n65786), .B(n69132), .Z(n65781) );
  XOR U84081 ( .A(n65780), .B(n65781), .Z(n69135) );
  IV U84082 ( .A(n63846), .Z(n63847) );
  NOR U84083 ( .A(n63848), .B(n63847), .Z(n69131) );
  IV U84084 ( .A(n63849), .Z(n63850) );
  NOR U84085 ( .A(n63851), .B(n63850), .Z(n69134) );
  NOR U84086 ( .A(n69131), .B(n69134), .Z(n63852) );
  XOR U84087 ( .A(n69135), .B(n63852), .Z(n69137) );
  IV U84088 ( .A(n63853), .Z(n63855) );
  NOR U84089 ( .A(n63855), .B(n63854), .Z(n70725) );
  NOR U84090 ( .A(n70725), .B(n74199), .Z(n69138) );
  XOR U84091 ( .A(n69137), .B(n69138), .Z(n69140) );
  IV U84092 ( .A(n63856), .Z(n63858) );
  NOR U84093 ( .A(n63858), .B(n63857), .Z(n69139) );
  IV U84094 ( .A(n63859), .Z(n65777) );
  NOR U84095 ( .A(n63860), .B(n65777), .Z(n63861) );
  NOR U84096 ( .A(n69139), .B(n63861), .Z(n63862) );
  XOR U84097 ( .A(n69140), .B(n63862), .Z(n65770) );
  XOR U84098 ( .A(n63863), .B(n65770), .Z(n74227) );
  XOR U84099 ( .A(n65764), .B(n74227), .Z(n65762) );
  IV U84100 ( .A(n65762), .Z(n63870) );
  IV U84101 ( .A(n63864), .Z(n63866) );
  NOR U84102 ( .A(n63866), .B(n63865), .Z(n65766) );
  IV U84103 ( .A(n63867), .Z(n63868) );
  NOR U84104 ( .A(n63868), .B(n63872), .Z(n65760) );
  NOR U84105 ( .A(n65766), .B(n65760), .Z(n63869) );
  XOR U84106 ( .A(n63870), .B(n63869), .Z(n69153) );
  IV U84107 ( .A(n63871), .Z(n63873) );
  NOR U84108 ( .A(n63873), .B(n63872), .Z(n69151) );
  XOR U84109 ( .A(n69153), .B(n69151), .Z(n69155) );
  XOR U84110 ( .A(n63874), .B(n69155), .Z(n65752) );
  XOR U84111 ( .A(n65754), .B(n65752), .Z(n65756) );
  XOR U84112 ( .A(n65755), .B(n65756), .Z(n69159) );
  XOR U84113 ( .A(n69158), .B(n69159), .Z(n69162) );
  XOR U84114 ( .A(n69161), .B(n69162), .Z(n65750) );
  XOR U84115 ( .A(n65749), .B(n65750), .Z(n65745) );
  XOR U84116 ( .A(n65744), .B(n65745), .Z(n69167) );
  XOR U84117 ( .A(n65747), .B(n69167), .Z(n69174) );
  IV U84118 ( .A(n63875), .Z(n63876) );
  NOR U84119 ( .A(n63876), .B(n63881), .Z(n69172) );
  IV U84120 ( .A(n63877), .Z(n63879) );
  NOR U84121 ( .A(n63879), .B(n63878), .Z(n69166) );
  IV U84122 ( .A(n63880), .Z(n63882) );
  NOR U84123 ( .A(n63882), .B(n63881), .Z(n65742) );
  NOR U84124 ( .A(n69166), .B(n65742), .Z(n63883) );
  IV U84125 ( .A(n63883), .Z(n63884) );
  NOR U84126 ( .A(n69172), .B(n63884), .Z(n63885) );
  XOR U84127 ( .A(n69174), .B(n63885), .Z(n65739) );
  IV U84128 ( .A(n63886), .Z(n63887) );
  NOR U84129 ( .A(n63888), .B(n63887), .Z(n65740) );
  IV U84130 ( .A(n63889), .Z(n63891) );
  NOR U84131 ( .A(n63891), .B(n63890), .Z(n69169) );
  NOR U84132 ( .A(n65740), .B(n69169), .Z(n63892) );
  XOR U84133 ( .A(n65739), .B(n63892), .Z(n65734) );
  XOR U84134 ( .A(n65733), .B(n65734), .Z(n65737) );
  NOR U84135 ( .A(n63894), .B(n63893), .Z(n65736) );
  IV U84136 ( .A(n63895), .Z(n63896) );
  NOR U84137 ( .A(n63897), .B(n63896), .Z(n63898) );
  NOR U84138 ( .A(n65736), .B(n63898), .Z(n65728) );
  XOR U84139 ( .A(n65737), .B(n65728), .Z(n69177) );
  XOR U84140 ( .A(n69178), .B(n69177), .Z(n69181) );
  IV U84141 ( .A(n63899), .Z(n63900) );
  NOR U84142 ( .A(n63901), .B(n63900), .Z(n69180) );
  IV U84143 ( .A(n63902), .Z(n63903) );
  NOR U84144 ( .A(n63904), .B(n63903), .Z(n65726) );
  NOR U84145 ( .A(n69180), .B(n65726), .Z(n63905) );
  XOR U84146 ( .A(n69181), .B(n63905), .Z(n63906) );
  NOR U84147 ( .A(n63907), .B(n63906), .Z(n63910) );
  IV U84148 ( .A(n63907), .Z(n63909) );
  XOR U84149 ( .A(n69180), .B(n69181), .Z(n63908) );
  NOR U84150 ( .A(n63909), .B(n63908), .Z(n74279) );
  NOR U84151 ( .A(n63910), .B(n74279), .Z(n63911) );
  IV U84152 ( .A(n63911), .Z(n65723) );
  XOR U84153 ( .A(n65722), .B(n65723), .Z(n69196) );
  IV U84154 ( .A(n63912), .Z(n63913) );
  NOR U84155 ( .A(n63914), .B(n63913), .Z(n69185) );
  IV U84156 ( .A(n63915), .Z(n63916) );
  NOR U84157 ( .A(n63917), .B(n63916), .Z(n69195) );
  NOR U84158 ( .A(n69185), .B(n69195), .Z(n63918) );
  XOR U84159 ( .A(n69196), .B(n63918), .Z(n63919) );
  IV U84160 ( .A(n63919), .Z(n69194) );
  XOR U84161 ( .A(n69192), .B(n69194), .Z(n65720) );
  XOR U84162 ( .A(n65719), .B(n65720), .Z(n65715) );
  XOR U84163 ( .A(n65713), .B(n65715), .Z(n65718) );
  XOR U84164 ( .A(n63920), .B(n65718), .Z(n79724) );
  NOR U84165 ( .A(n65709), .B(n65704), .Z(n63921) );
  XOR U84166 ( .A(n79724), .B(n63921), .Z(n65706) );
  XOR U84167 ( .A(n63922), .B(n65706), .Z(n65696) );
  IV U84168 ( .A(n63923), .Z(n63924) );
  NOR U84169 ( .A(n63925), .B(n63924), .Z(n65698) );
  IV U84170 ( .A(n63926), .Z(n63927) );
  NOR U84171 ( .A(n63928), .B(n63927), .Z(n65695) );
  NOR U84172 ( .A(n65698), .B(n65695), .Z(n63929) );
  XOR U84173 ( .A(n65696), .B(n63929), .Z(n69205) );
  XOR U84174 ( .A(n69203), .B(n69205), .Z(n65692) );
  XOR U84175 ( .A(n65691), .B(n65692), .Z(n69202) );
  XOR U84176 ( .A(n69201), .B(n69202), .Z(n63949) );
  IV U84177 ( .A(n63930), .Z(n69213) );
  NOR U84178 ( .A(n63947), .B(n69213), .Z(n63938) );
  IV U84179 ( .A(n63938), .Z(n63931) );
  NOR U84180 ( .A(n63949), .B(n63931), .Z(n63940) );
  IV U84181 ( .A(n63948), .Z(n63932) );
  NOR U84182 ( .A(n63947), .B(n63932), .Z(n63934) );
  IV U84183 ( .A(n63934), .Z(n63933) );
  NOR U84184 ( .A(n63933), .B(n69202), .Z(n70692) );
  NOR U84185 ( .A(n63949), .B(n63934), .Z(n63935) );
  NOR U84186 ( .A(n70692), .B(n63935), .Z(n63936) );
  IV U84187 ( .A(n63936), .Z(n63937) );
  NOR U84188 ( .A(n63938), .B(n63937), .Z(n63939) );
  NOR U84189 ( .A(n63940), .B(n63939), .Z(n63956) );
  IV U84190 ( .A(n63956), .Z(n63941) );
  NOR U84191 ( .A(n63942), .B(n63941), .Z(n63960) );
  IV U84192 ( .A(n63943), .Z(n63944) );
  NOR U84193 ( .A(n63945), .B(n63944), .Z(n63954) );
  IV U84194 ( .A(n63946), .Z(n63953) );
  XOR U84195 ( .A(n63948), .B(n63947), .Z(n63951) );
  IV U84196 ( .A(n63949), .Z(n63950) );
  NOR U84197 ( .A(n63951), .B(n63950), .Z(n63952) );
  IV U84198 ( .A(n63952), .Z(n69212) );
  NOR U84199 ( .A(n63953), .B(n69212), .Z(n69214) );
  IV U84200 ( .A(n69214), .Z(n70691) );
  NOR U84201 ( .A(n63954), .B(n70691), .Z(n63957) );
  IV U84202 ( .A(n63954), .Z(n63955) );
  NOR U84203 ( .A(n63956), .B(n63955), .Z(n70688) );
  NOR U84204 ( .A(n63957), .B(n70688), .Z(n63958) );
  IV U84205 ( .A(n63958), .Z(n63959) );
  NOR U84206 ( .A(n63960), .B(n63959), .Z(n65689) );
  XOR U84207 ( .A(n63961), .B(n65689), .Z(n65684) );
  IV U84208 ( .A(n63962), .Z(n63963) );
  NOR U84209 ( .A(n63963), .B(n63965), .Z(n65682) );
  XOR U84210 ( .A(n65684), .B(n65682), .Z(n65687) );
  IV U84211 ( .A(n63964), .Z(n63966) );
  NOR U84212 ( .A(n63966), .B(n63965), .Z(n65685) );
  XOR U84213 ( .A(n65687), .B(n65685), .Z(n69222) );
  XOR U84214 ( .A(n69221), .B(n69222), .Z(n74353) );
  IV U84215 ( .A(n63967), .Z(n63968) );
  NOR U84216 ( .A(n63969), .B(n63968), .Z(n69224) );
  IV U84217 ( .A(n63970), .Z(n63972) );
  NOR U84218 ( .A(n63972), .B(n63971), .Z(n69227) );
  NOR U84219 ( .A(n69224), .B(n69227), .Z(n74354) );
  XOR U84220 ( .A(n74353), .B(n74354), .Z(n65673) );
  XOR U84221 ( .A(n63973), .B(n65673), .Z(n65677) );
  IV U84222 ( .A(n65677), .Z(n63981) );
  IV U84223 ( .A(n63974), .Z(n63984) );
  IV U84224 ( .A(n63975), .Z(n63976) );
  NOR U84225 ( .A(n63984), .B(n63976), .Z(n65670) );
  IV U84226 ( .A(n63977), .Z(n63979) );
  NOR U84227 ( .A(n63979), .B(n63978), .Z(n65676) );
  NOR U84228 ( .A(n65670), .B(n65676), .Z(n63980) );
  XOR U84229 ( .A(n63981), .B(n63980), .Z(n69232) );
  IV U84230 ( .A(n63982), .Z(n63983) );
  NOR U84231 ( .A(n63984), .B(n63983), .Z(n69230) );
  XOR U84232 ( .A(n69232), .B(n69230), .Z(n69234) );
  NOR U84233 ( .A(n63991), .B(n69234), .Z(n70669) );
  IV U84234 ( .A(n63985), .Z(n63986) );
  NOR U84235 ( .A(n63987), .B(n63986), .Z(n65664) );
  IV U84236 ( .A(n63988), .Z(n63989) );
  NOR U84237 ( .A(n63990), .B(n63989), .Z(n69233) );
  XOR U84238 ( .A(n69233), .B(n69234), .Z(n65665) );
  IV U84239 ( .A(n65665), .Z(n63992) );
  XOR U84240 ( .A(n65664), .B(n63992), .Z(n63994) );
  NOR U84241 ( .A(n63992), .B(n63991), .Z(n63993) );
  NOR U84242 ( .A(n63994), .B(n63993), .Z(n63995) );
  NOR U84243 ( .A(n70669), .B(n63995), .Z(n65668) );
  XOR U84244 ( .A(n63996), .B(n65668), .Z(n69245) );
  XOR U84245 ( .A(n63997), .B(n69245), .Z(n65661) );
  XOR U84246 ( .A(n65662), .B(n65661), .Z(n65657) );
  XOR U84247 ( .A(n65655), .B(n65657), .Z(n65659) );
  XOR U84248 ( .A(n63998), .B(n65659), .Z(n65645) );
  XOR U84249 ( .A(n63999), .B(n65645), .Z(n69251) );
  IV U84250 ( .A(n64000), .Z(n64004) );
  NOR U84251 ( .A(n64002), .B(n64001), .Z(n64003) );
  IV U84252 ( .A(n64003), .Z(n64006) );
  NOR U84253 ( .A(n64004), .B(n64006), .Z(n69250) );
  IV U84254 ( .A(n64005), .Z(n64007) );
  NOR U84255 ( .A(n64007), .B(n64006), .Z(n64008) );
  IV U84256 ( .A(n64008), .Z(n65644) );
  XOR U84257 ( .A(n69250), .B(n65644), .Z(n64009) );
  XOR U84258 ( .A(n69251), .B(n64009), .Z(n64010) );
  IV U84259 ( .A(n64010), .Z(n69254) );
  XOR U84260 ( .A(n64011), .B(n69254), .Z(n69257) );
  NOR U84261 ( .A(n64013), .B(n64012), .Z(n69256) );
  IV U84262 ( .A(n64014), .Z(n69265) );
  IV U84263 ( .A(n64015), .Z(n64016) );
  NOR U84264 ( .A(n69265), .B(n64016), .Z(n64017) );
  NOR U84265 ( .A(n69256), .B(n64017), .Z(n64018) );
  XOR U84266 ( .A(n69257), .B(n64018), .Z(n70649) );
  IV U84267 ( .A(n64019), .Z(n64020) );
  NOR U84268 ( .A(n64020), .B(n69265), .Z(n74423) );
  IV U84269 ( .A(n64021), .Z(n64022) );
  NOR U84270 ( .A(n64023), .B(n64022), .Z(n70648) );
  NOR U84271 ( .A(n74423), .B(n70648), .Z(n65637) );
  XOR U84272 ( .A(n70649), .B(n65637), .Z(n65635) );
  IV U84273 ( .A(n64024), .Z(n64026) );
  NOR U84274 ( .A(n64026), .B(n64025), .Z(n65638) );
  NOR U84275 ( .A(n65638), .B(n65634), .Z(n64027) );
  XOR U84276 ( .A(n65635), .B(n64027), .Z(n65633) );
  IV U84277 ( .A(n64028), .Z(n64030) );
  NOR U84278 ( .A(n64030), .B(n64029), .Z(n65631) );
  IV U84279 ( .A(n64031), .Z(n65620) );
  NOR U84280 ( .A(n64032), .B(n65620), .Z(n65629) );
  NOR U84281 ( .A(n65631), .B(n65629), .Z(n64033) );
  XOR U84282 ( .A(n65633), .B(n64033), .Z(n69275) );
  IV U84283 ( .A(n64034), .Z(n64036) );
  NOR U84284 ( .A(n64036), .B(n64035), .Z(n64037) );
  NOR U84285 ( .A(n64037), .B(n69274), .Z(n64038) );
  XOR U84286 ( .A(n69275), .B(n64038), .Z(n65616) );
  XOR U84287 ( .A(n65614), .B(n65616), .Z(n65618) );
  XOR U84288 ( .A(n64039), .B(n65618), .Z(n65610) );
  NOR U84289 ( .A(n64040), .B(n65609), .Z(n64041) );
  NOR U84290 ( .A(n64042), .B(n64041), .Z(n64043) );
  XOR U84291 ( .A(n65610), .B(n64043), .Z(n76001) );
  XOR U84292 ( .A(n64044), .B(n76001), .Z(n79825) );
  XOR U84293 ( .A(n79826), .B(n79825), .Z(n69280) );
  XOR U84294 ( .A(n65599), .B(n69280), .Z(n69293) );
  IV U84295 ( .A(n64045), .Z(n64047) );
  NOR U84296 ( .A(n64047), .B(n64046), .Z(n69292) );
  IV U84297 ( .A(n64048), .Z(n64049) );
  NOR U84298 ( .A(n64050), .B(n64049), .Z(n69290) );
  NOR U84299 ( .A(n69292), .B(n69290), .Z(n64051) );
  XOR U84300 ( .A(n69293), .B(n64051), .Z(n65593) );
  XOR U84301 ( .A(n64052), .B(n65593), .Z(n65591) );
  XOR U84302 ( .A(n65589), .B(n65591), .Z(n65584) );
  XOR U84303 ( .A(n65583), .B(n65584), .Z(n70617) );
  XOR U84304 ( .A(n65586), .B(n70617), .Z(n65579) );
  NOR U84305 ( .A(n64053), .B(n70621), .Z(n65581) );
  IV U84306 ( .A(n64054), .Z(n64055) );
  NOR U84307 ( .A(n64056), .B(n64055), .Z(n65578) );
  NOR U84308 ( .A(n65581), .B(n65578), .Z(n64057) );
  XOR U84309 ( .A(n65579), .B(n64057), .Z(n64058) );
  IV U84310 ( .A(n64058), .Z(n65577) );
  XOR U84311 ( .A(n65575), .B(n65577), .Z(n65571) );
  XOR U84312 ( .A(n65569), .B(n65571), .Z(n65574) );
  XOR U84313 ( .A(n65572), .B(n65574), .Z(n69300) );
  XOR U84314 ( .A(n69299), .B(n69300), .Z(n69303) );
  XOR U84315 ( .A(n64059), .B(n69303), .Z(n65564) );
  XOR U84316 ( .A(n65565), .B(n65564), .Z(n69311) );
  IV U84317 ( .A(n64060), .Z(n64061) );
  NOR U84318 ( .A(n64062), .B(n64061), .Z(n65562) );
  IV U84319 ( .A(n64063), .Z(n64065) );
  NOR U84320 ( .A(n64065), .B(n64064), .Z(n69310) );
  NOR U84321 ( .A(n65562), .B(n69310), .Z(n64066) );
  XOR U84322 ( .A(n69311), .B(n64066), .Z(n69307) );
  IV U84323 ( .A(n64067), .Z(n64069) );
  NOR U84324 ( .A(n64069), .B(n64068), .Z(n69308) );
  IV U84325 ( .A(n64070), .Z(n64072) );
  NOR U84326 ( .A(n64072), .B(n64071), .Z(n69319) );
  NOR U84327 ( .A(n69308), .B(n69319), .Z(n64073) );
  XOR U84328 ( .A(n69307), .B(n64073), .Z(n69317) );
  XOR U84329 ( .A(n69318), .B(n69317), .Z(n69330) );
  IV U84330 ( .A(n64074), .Z(n64076) );
  NOR U84331 ( .A(n64076), .B(n64075), .Z(n69314) );
  IV U84332 ( .A(n64077), .Z(n64079) );
  NOR U84333 ( .A(n64079), .B(n64078), .Z(n69329) );
  NOR U84334 ( .A(n69314), .B(n69329), .Z(n64080) );
  XOR U84335 ( .A(n69330), .B(n64080), .Z(n65561) );
  XOR U84336 ( .A(n65559), .B(n65561), .Z(n64093) );
  XOR U84337 ( .A(n64082), .B(n64081), .Z(n64083) );
  NOR U84338 ( .A(n64084), .B(n64083), .Z(n64085) );
  IV U84339 ( .A(n64085), .Z(n64091) );
  NOR U84340 ( .A(n64086), .B(n64116), .Z(n64087) );
  IV U84341 ( .A(n64087), .Z(n64088) );
  NOR U84342 ( .A(n64089), .B(n64088), .Z(n64090) );
  IV U84343 ( .A(n64090), .Z(n64101) );
  NOR U84344 ( .A(n64091), .B(n64101), .Z(n64108) );
  IV U84345 ( .A(n64108), .Z(n64092) );
  NOR U84346 ( .A(n64093), .B(n64092), .Z(n70587) );
  IV U84347 ( .A(n64094), .Z(n64096) );
  NOR U84348 ( .A(n64096), .B(n64095), .Z(n64097) );
  IV U84349 ( .A(n64097), .Z(n64098) );
  NOR U84350 ( .A(n64098), .B(n64116), .Z(n64105) );
  IV U84351 ( .A(n64105), .Z(n64099) );
  NOR U84352 ( .A(n65561), .B(n64099), .Z(n70581) );
  IV U84353 ( .A(n64100), .Z(n64102) );
  NOR U84354 ( .A(n64102), .B(n64101), .Z(n65557) );
  NOR U84355 ( .A(n65559), .B(n65557), .Z(n64103) );
  XOR U84356 ( .A(n65561), .B(n64103), .Z(n64104) );
  NOR U84357 ( .A(n64105), .B(n64104), .Z(n64106) );
  IV U84358 ( .A(n64106), .Z(n64107) );
  NOR U84359 ( .A(n64108), .B(n64107), .Z(n64109) );
  NOR U84360 ( .A(n70581), .B(n64109), .Z(n64110) );
  IV U84361 ( .A(n64110), .Z(n64111) );
  NOR U84362 ( .A(n70587), .B(n64111), .Z(n65552) );
  IV U84363 ( .A(n64112), .Z(n64114) );
  NOR U84364 ( .A(n64114), .B(n64113), .Z(n65551) );
  IV U84365 ( .A(n64115), .Z(n64117) );
  NOR U84366 ( .A(n64117), .B(n64116), .Z(n65554) );
  NOR U84367 ( .A(n65551), .B(n65554), .Z(n64118) );
  XOR U84368 ( .A(n65552), .B(n64118), .Z(n65549) );
  XOR U84369 ( .A(n65548), .B(n65549), .Z(n65544) );
  XOR U84370 ( .A(n65542), .B(n65544), .Z(n65547) );
  XOR U84371 ( .A(n64119), .B(n65547), .Z(n64120) );
  IV U84372 ( .A(n64120), .Z(n69338) );
  XOR U84373 ( .A(n69336), .B(n69338), .Z(n69340) );
  XOR U84374 ( .A(n69339), .B(n69340), .Z(n70560) );
  IV U84375 ( .A(n64121), .Z(n64123) );
  NOR U84376 ( .A(n64123), .B(n64122), .Z(n70558) );
  IV U84377 ( .A(n64124), .Z(n64126) );
  NOR U84378 ( .A(n64126), .B(n64125), .Z(n74495) );
  NOR U84379 ( .A(n70558), .B(n74495), .Z(n65535) );
  XOR U84380 ( .A(n70560), .B(n65535), .Z(n65536) );
  XOR U84381 ( .A(n65537), .B(n65536), .Z(n65531) );
  XOR U84382 ( .A(n65529), .B(n65531), .Z(n65533) );
  XOR U84383 ( .A(n64127), .B(n65533), .Z(n65521) );
  XOR U84384 ( .A(n65522), .B(n65521), .Z(n70553) );
  IV U84385 ( .A(n64128), .Z(n64132) );
  NOR U84386 ( .A(n64132), .B(n64129), .Z(n74509) );
  IV U84387 ( .A(n64130), .Z(n64131) );
  NOR U84388 ( .A(n64132), .B(n64131), .Z(n70552) );
  NOR U84389 ( .A(n74509), .B(n70552), .Z(n65524) );
  XOR U84390 ( .A(n70553), .B(n65524), .Z(n65515) );
  XOR U84391 ( .A(n65517), .B(n65515), .Z(n65519) );
  XOR U84392 ( .A(n65518), .B(n65519), .Z(n65507) );
  NOR U84393 ( .A(n64133), .B(n65509), .Z(n64137) );
  IV U84394 ( .A(n64134), .Z(n64136) );
  NOR U84395 ( .A(n64136), .B(n64135), .Z(n65505) );
  NOR U84396 ( .A(n64137), .B(n65505), .Z(n64138) );
  XOR U84397 ( .A(n65507), .B(n64138), .Z(n65496) );
  XOR U84398 ( .A(n64139), .B(n65496), .Z(n65491) );
  XOR U84399 ( .A(n64145), .B(n65491), .Z(n64140) );
  NOR U84400 ( .A(n64141), .B(n64140), .Z(n79949) );
  IV U84401 ( .A(n64142), .Z(n64143) );
  NOR U84402 ( .A(n64144), .B(n64143), .Z(n65488) );
  NOR U84403 ( .A(n64145), .B(n65488), .Z(n64146) );
  XOR U84404 ( .A(n65491), .B(n64146), .Z(n64147) );
  NOR U84405 ( .A(n64148), .B(n64147), .Z(n64149) );
  NOR U84406 ( .A(n79949), .B(n64149), .Z(n64150) );
  IV U84407 ( .A(n64150), .Z(n75905) );
  NOR U84408 ( .A(n65487), .B(n75894), .Z(n64151) );
  IV U84409 ( .A(n64151), .Z(n64152) );
  NOR U84410 ( .A(n65485), .B(n64152), .Z(n64153) );
  XOR U84411 ( .A(n75905), .B(n64153), .Z(n69348) );
  IV U84412 ( .A(n64154), .Z(n64162) );
  IV U84413 ( .A(n64157), .Z(n64155) );
  NOR U84414 ( .A(n64162), .B(n64155), .Z(n65481) );
  IV U84415 ( .A(n64156), .Z(n64159) );
  XOR U84416 ( .A(n64157), .B(n64162), .Z(n64158) );
  NOR U84417 ( .A(n64159), .B(n64158), .Z(n69347) );
  NOR U84418 ( .A(n65481), .B(n69347), .Z(n64160) );
  XOR U84419 ( .A(n69348), .B(n64160), .Z(n65475) );
  IV U84420 ( .A(n64161), .Z(n64163) );
  NOR U84421 ( .A(n64163), .B(n64162), .Z(n65478) );
  IV U84422 ( .A(n64164), .Z(n64165) );
  NOR U84423 ( .A(n64166), .B(n64165), .Z(n65476) );
  NOR U84424 ( .A(n65478), .B(n65476), .Z(n64167) );
  XOR U84425 ( .A(n65475), .B(n64167), .Z(n69353) );
  IV U84426 ( .A(n69353), .Z(n64174) );
  IV U84427 ( .A(n64168), .Z(n64169) );
  NOR U84428 ( .A(n64170), .B(n64169), .Z(n69350) );
  IV U84429 ( .A(n64171), .Z(n64172) );
  NOR U84430 ( .A(n64172), .B(n64176), .Z(n69352) );
  NOR U84431 ( .A(n69350), .B(n69352), .Z(n64173) );
  XOR U84432 ( .A(n64174), .B(n64173), .Z(n69359) );
  IV U84433 ( .A(n64175), .Z(n64177) );
  NOR U84434 ( .A(n64177), .B(n64176), .Z(n69355) );
  XOR U84435 ( .A(n69359), .B(n69355), .Z(n69362) );
  XOR U84436 ( .A(n64178), .B(n69362), .Z(n65470) );
  XOR U84437 ( .A(n65471), .B(n65470), .Z(n65474) );
  XOR U84438 ( .A(n64179), .B(n65474), .Z(n69367) );
  XOR U84439 ( .A(n69365), .B(n69367), .Z(n69369) );
  XOR U84440 ( .A(n69368), .B(n69369), .Z(n69373) );
  IV U84441 ( .A(n64180), .Z(n64182) );
  NOR U84442 ( .A(n64182), .B(n64181), .Z(n69372) );
  IV U84443 ( .A(n64183), .Z(n64185) );
  NOR U84444 ( .A(n64185), .B(n64184), .Z(n65465) );
  NOR U84445 ( .A(n69372), .B(n65465), .Z(n64186) );
  XOR U84446 ( .A(n69373), .B(n64186), .Z(n65459) );
  XOR U84447 ( .A(n64187), .B(n65459), .Z(n65457) );
  IV U84448 ( .A(n64188), .Z(n64189) );
  NOR U84449 ( .A(n64195), .B(n64189), .Z(n65454) );
  IV U84450 ( .A(n64190), .Z(n64191) );
  NOR U84451 ( .A(n64192), .B(n64191), .Z(n65456) );
  NOR U84452 ( .A(n65454), .B(n65456), .Z(n64193) );
  XOR U84453 ( .A(n65457), .B(n64193), .Z(n64200) );
  IV U84454 ( .A(n64200), .Z(n64194) );
  NOR U84455 ( .A(n64195), .B(n64194), .Z(n64196) );
  IV U84456 ( .A(n64196), .Z(n64197) );
  NOR U84457 ( .A(n64199), .B(n64197), .Z(n74571) );
  NOR U84458 ( .A(n64199), .B(n64198), .Z(n64201) );
  NOR U84459 ( .A(n64201), .B(n64200), .Z(n64202) );
  NOR U84460 ( .A(n74571), .B(n64202), .Z(n65451) );
  XOR U84461 ( .A(n65453), .B(n65451), .Z(n65447) );
  IV U84462 ( .A(n64203), .Z(n64205) );
  IV U84463 ( .A(n64204), .Z(n64212) );
  NOR U84464 ( .A(n64205), .B(n64212), .Z(n64206) );
  IV U84465 ( .A(n64206), .Z(n65446) );
  XOR U84466 ( .A(n65447), .B(n65446), .Z(n65444) );
  IV U84467 ( .A(n64207), .Z(n64208) );
  NOR U84468 ( .A(n64209), .B(n64208), .Z(n65443) );
  IV U84469 ( .A(n64210), .Z(n64211) );
  NOR U84470 ( .A(n64212), .B(n64211), .Z(n65448) );
  NOR U84471 ( .A(n65443), .B(n65448), .Z(n64213) );
  XOR U84472 ( .A(n65444), .B(n64213), .Z(n65440) );
  XOR U84473 ( .A(n65438), .B(n65440), .Z(n65435) );
  XOR U84474 ( .A(n64214), .B(n65435), .Z(n64215) );
  IV U84475 ( .A(n64215), .Z(n69379) );
  IV U84476 ( .A(n64216), .Z(n64217) );
  NOR U84477 ( .A(n64218), .B(n64217), .Z(n69378) );
  IV U84478 ( .A(n64219), .Z(n64221) );
  NOR U84479 ( .A(n64221), .B(n64220), .Z(n65430) );
  NOR U84480 ( .A(n69378), .B(n65430), .Z(n64222) );
  XOR U84481 ( .A(n69379), .B(n64222), .Z(n69383) );
  XOR U84482 ( .A(n69381), .B(n69383), .Z(n69391) );
  XOR U84483 ( .A(n64223), .B(n69391), .Z(n65424) );
  XOR U84484 ( .A(n65425), .B(n65424), .Z(n65428) );
  IV U84485 ( .A(n64224), .Z(n65423) );
  NOR U84486 ( .A(n65423), .B(n64225), .Z(n64226) );
  NOR U84487 ( .A(n65427), .B(n64226), .Z(n64227) );
  XOR U84488 ( .A(n65428), .B(n64227), .Z(n65418) );
  IV U84489 ( .A(n64228), .Z(n64230) );
  NOR U84490 ( .A(n64230), .B(n64229), .Z(n64231) );
  IV U84491 ( .A(n64231), .Z(n65419) );
  XOR U84492 ( .A(n65418), .B(n65419), .Z(n69396) );
  XOR U84493 ( .A(n69395), .B(n69396), .Z(n69403) );
  XOR U84494 ( .A(n64232), .B(n69403), .Z(n69410) );
  XOR U84495 ( .A(n64233), .B(n69410), .Z(n65417) );
  XOR U84496 ( .A(n64234), .B(n65417), .Z(n65409) );
  XOR U84497 ( .A(n64235), .B(n65409), .Z(n65406) );
  XOR U84498 ( .A(n65404), .B(n65406), .Z(n65402) );
  XOR U84499 ( .A(n65401), .B(n65402), .Z(n65393) );
  XOR U84500 ( .A(n64236), .B(n65393), .Z(n64237) );
  IV U84501 ( .A(n64237), .Z(n65391) );
  XOR U84502 ( .A(n65389), .B(n65391), .Z(n65381) );
  IV U84503 ( .A(n64238), .Z(n64239) );
  NOR U84504 ( .A(n65385), .B(n64239), .Z(n64240) );
  XOR U84505 ( .A(n65381), .B(n64240), .Z(n65378) );
  XOR U84506 ( .A(n65377), .B(n65378), .Z(n69422) );
  IV U84507 ( .A(n64241), .Z(n64242) );
  NOR U84508 ( .A(n64248), .B(n64242), .Z(n69420) );
  XOR U84509 ( .A(n69422), .B(n69420), .Z(n69429) );
  IV U84510 ( .A(n64243), .Z(n64245) );
  NOR U84511 ( .A(n64245), .B(n64244), .Z(n69427) );
  IV U84512 ( .A(n64246), .Z(n64247) );
  NOR U84513 ( .A(n64248), .B(n64247), .Z(n65375) );
  NOR U84514 ( .A(n69427), .B(n65375), .Z(n64249) );
  XOR U84515 ( .A(n69429), .B(n64249), .Z(n65370) );
  XOR U84516 ( .A(n64250), .B(n65370), .Z(n69438) );
  XOR U84517 ( .A(n69437), .B(n69438), .Z(n65354) );
  NOR U84518 ( .A(n64252), .B(n64251), .Z(n64253) );
  NOR U84519 ( .A(n64253), .B(n69434), .Z(n65352) );
  XOR U84520 ( .A(n65354), .B(n65352), .Z(n69444) );
  XOR U84521 ( .A(n69442), .B(n69444), .Z(n69449) );
  XOR U84522 ( .A(n64254), .B(n69449), .Z(n64255) );
  IV U84523 ( .A(n64255), .Z(n69452) );
  XOR U84524 ( .A(n69451), .B(n69452), .Z(n65350) );
  XOR U84525 ( .A(n65349), .B(n65350), .Z(n69462) );
  IV U84526 ( .A(n64256), .Z(n64257) );
  NOR U84527 ( .A(n64258), .B(n64257), .Z(n69461) );
  IV U84528 ( .A(n64259), .Z(n64261) );
  NOR U84529 ( .A(n64261), .B(n64260), .Z(n65347) );
  NOR U84530 ( .A(n69461), .B(n65347), .Z(n64262) );
  XOR U84531 ( .A(n69462), .B(n64262), .Z(n64263) );
  IV U84532 ( .A(n64263), .Z(n65343) );
  XOR U84533 ( .A(n65341), .B(n65343), .Z(n65345) );
  XOR U84534 ( .A(n65344), .B(n65345), .Z(n69466) );
  XOR U84535 ( .A(n64264), .B(n69466), .Z(n64265) );
  IV U84536 ( .A(n64265), .Z(n69468) );
  XOR U84537 ( .A(n69469), .B(n69468), .Z(n64266) );
  NOR U84538 ( .A(n64267), .B(n64266), .Z(n64270) );
  IV U84539 ( .A(n64267), .Z(n64269) );
  XOR U84540 ( .A(n65338), .B(n69466), .Z(n64268) );
  NOR U84541 ( .A(n64269), .B(n64268), .Z(n70419) );
  NOR U84542 ( .A(n64270), .B(n70419), .Z(n64271) );
  IV U84543 ( .A(n64271), .Z(n65336) );
  XOR U84544 ( .A(n65335), .B(n65336), .Z(n69476) );
  XOR U84545 ( .A(n69473), .B(n69476), .Z(n65330) );
  XOR U84546 ( .A(n65331), .B(n65330), .Z(n65327) );
  IV U84547 ( .A(n64272), .Z(n64273) );
  NOR U84548 ( .A(n64273), .B(n65334), .Z(n64274) );
  IV U84549 ( .A(n64274), .Z(n65328) );
  XOR U84550 ( .A(n65327), .B(n65328), .Z(n65322) );
  XOR U84551 ( .A(n65321), .B(n65322), .Z(n65325) );
  XOR U84552 ( .A(n65324), .B(n65325), .Z(n65316) );
  XOR U84553 ( .A(n65315), .B(n65316), .Z(n65319) );
  XOR U84554 ( .A(n65318), .B(n65319), .Z(n65310) );
  XOR U84555 ( .A(n65309), .B(n65310), .Z(n65313) );
  XOR U84556 ( .A(n65312), .B(n65313), .Z(n69490) );
  IV U84557 ( .A(n64275), .Z(n64276) );
  NOR U84558 ( .A(n64277), .B(n64276), .Z(n65306) );
  IV U84559 ( .A(n69483), .Z(n64278) );
  NOR U84560 ( .A(n64278), .B(n69482), .Z(n69489) );
  NOR U84561 ( .A(n65306), .B(n69489), .Z(n64279) );
  XOR U84562 ( .A(n69490), .B(n64279), .Z(n65303) );
  IV U84563 ( .A(n64280), .Z(n69488) );
  NOR U84564 ( .A(n69488), .B(n69482), .Z(n64284) );
  IV U84565 ( .A(n64281), .Z(n64283) );
  NOR U84566 ( .A(n64283), .B(n64282), .Z(n65304) );
  NOR U84567 ( .A(n64284), .B(n65304), .Z(n64285) );
  XOR U84568 ( .A(n65303), .B(n64285), .Z(n65301) );
  IV U84569 ( .A(n64286), .Z(n64288) );
  NOR U84570 ( .A(n64288), .B(n64287), .Z(n65300) );
  IV U84571 ( .A(n64289), .Z(n64291) );
  NOR U84572 ( .A(n64291), .B(n64290), .Z(n65298) );
  NOR U84573 ( .A(n65300), .B(n65298), .Z(n64292) );
  XOR U84574 ( .A(n65301), .B(n64292), .Z(n65285) );
  IV U84575 ( .A(n64293), .Z(n64294) );
  NOR U84576 ( .A(n64295), .B(n64294), .Z(n65286) );
  NOR U84577 ( .A(n64296), .B(n65291), .Z(n64300) );
  IV U84578 ( .A(n64297), .Z(n64298) );
  NOR U84579 ( .A(n64299), .B(n64298), .Z(n65288) );
  NOR U84580 ( .A(n64300), .B(n65288), .Z(n64301) );
  IV U84581 ( .A(n64301), .Z(n64302) );
  NOR U84582 ( .A(n65286), .B(n64302), .Z(n64303) );
  XOR U84583 ( .A(n65285), .B(n64303), .Z(n65280) );
  XOR U84584 ( .A(n65279), .B(n65280), .Z(n65283) );
  XOR U84585 ( .A(n65282), .B(n65283), .Z(n69496) );
  IV U84586 ( .A(n64304), .Z(n64305) );
  NOR U84587 ( .A(n64306), .B(n64305), .Z(n65276) );
  IV U84588 ( .A(n64307), .Z(n64309) );
  NOR U84589 ( .A(n64309), .B(n64308), .Z(n69495) );
  NOR U84590 ( .A(n65276), .B(n69495), .Z(n64310) );
  XOR U84591 ( .A(n69496), .B(n64310), .Z(n69499) );
  XOR U84592 ( .A(n69500), .B(n69499), .Z(n69503) );
  XOR U84593 ( .A(n69502), .B(n69503), .Z(n64314) );
  IV U84594 ( .A(n64311), .Z(n64312) );
  NOR U84595 ( .A(n64312), .B(n64325), .Z(n64320) );
  IV U84596 ( .A(n64320), .Z(n64313) );
  NOR U84597 ( .A(n64314), .B(n64313), .Z(n75739) );
  IV U84598 ( .A(n64315), .Z(n64317) );
  NOR U84599 ( .A(n64317), .B(n64316), .Z(n65274) );
  NOR U84600 ( .A(n69502), .B(n65274), .Z(n64318) );
  XOR U84601 ( .A(n69503), .B(n64318), .Z(n64319) );
  NOR U84602 ( .A(n64320), .B(n64319), .Z(n64321) );
  NOR U84603 ( .A(n75739), .B(n64321), .Z(n64322) );
  IV U84604 ( .A(n64322), .Z(n65273) );
  IV U84605 ( .A(n64323), .Z(n64324) );
  NOR U84606 ( .A(n64325), .B(n64324), .Z(n65271) );
  XOR U84607 ( .A(n65273), .B(n65271), .Z(n65270) );
  XOR U84608 ( .A(n65268), .B(n65270), .Z(n64326) );
  NOR U84609 ( .A(n64327), .B(n64326), .Z(n70378) );
  IV U84610 ( .A(n64328), .Z(n64329) );
  NOR U84611 ( .A(n64330), .B(n64329), .Z(n65266) );
  NOR U84612 ( .A(n65268), .B(n65266), .Z(n64331) );
  XOR U84613 ( .A(n65270), .B(n64331), .Z(n64332) );
  NOR U84614 ( .A(n64333), .B(n64332), .Z(n64334) );
  NOR U84615 ( .A(n70378), .B(n64334), .Z(n69507) );
  IV U84616 ( .A(n64335), .Z(n64336) );
  NOR U84617 ( .A(n64336), .B(n64339), .Z(n64337) );
  IV U84618 ( .A(n64337), .Z(n69508) );
  XOR U84619 ( .A(n69507), .B(n69508), .Z(n69518) );
  IV U84620 ( .A(n64338), .Z(n64342) );
  NOR U84621 ( .A(n64340), .B(n64339), .Z(n64341) );
  IV U84622 ( .A(n64341), .Z(n64344) );
  NOR U84623 ( .A(n64342), .B(n64344), .Z(n69516) );
  XOR U84624 ( .A(n69518), .B(n69516), .Z(n69515) );
  IV U84625 ( .A(n64343), .Z(n64345) );
  NOR U84626 ( .A(n64345), .B(n64344), .Z(n69513) );
  XOR U84627 ( .A(n69515), .B(n69513), .Z(n65264) );
  XOR U84628 ( .A(n65263), .B(n65264), .Z(n69528) );
  IV U84629 ( .A(n64346), .Z(n64347) );
  NOR U84630 ( .A(n64348), .B(n64347), .Z(n65261) );
  IV U84631 ( .A(n64349), .Z(n64350) );
  NOR U84632 ( .A(n64351), .B(n64350), .Z(n69527) );
  NOR U84633 ( .A(n65261), .B(n69527), .Z(n64352) );
  XOR U84634 ( .A(n69528), .B(n64352), .Z(n69531) );
  XOR U84635 ( .A(n64353), .B(n69531), .Z(n65260) );
  XOR U84636 ( .A(n64354), .B(n65260), .Z(n65254) );
  XOR U84637 ( .A(n65256), .B(n65254), .Z(n70358) );
  XOR U84638 ( .A(n65251), .B(n70358), .Z(n65247) );
  IV U84639 ( .A(n64355), .Z(n64356) );
  NOR U84640 ( .A(n64357), .B(n64356), .Z(n65246) );
  IV U84641 ( .A(n64358), .Z(n64360) );
  NOR U84642 ( .A(n64360), .B(n64359), .Z(n69540) );
  NOR U84643 ( .A(n65246), .B(n69540), .Z(n64361) );
  XOR U84644 ( .A(n65247), .B(n64361), .Z(n69544) );
  IV U84645 ( .A(n64362), .Z(n64364) );
  NOR U84646 ( .A(n64364), .B(n64363), .Z(n69542) );
  XOR U84647 ( .A(n69544), .B(n69542), .Z(n69546) );
  XOR U84648 ( .A(n69545), .B(n69546), .Z(n65244) );
  XOR U84649 ( .A(n65245), .B(n65244), .Z(n64365) );
  XOR U84650 ( .A(n64366), .B(n64365), .Z(n65239) );
  XOR U84651 ( .A(n64367), .B(n65239), .Z(n65232) );
  XOR U84652 ( .A(n65230), .B(n65232), .Z(n69550) );
  XOR U84653 ( .A(n64368), .B(n69550), .Z(n64369) );
  IV U84654 ( .A(n64369), .Z(n69554) );
  XOR U84655 ( .A(n69552), .B(n69554), .Z(n69556) );
  XOR U84656 ( .A(n69555), .B(n69556), .Z(n69563) );
  NOR U84657 ( .A(n64370), .B(n64371), .Z(n64375) );
  IV U84658 ( .A(n64370), .Z(n64373) );
  IV U84659 ( .A(n64371), .Z(n64372) );
  NOR U84660 ( .A(n64373), .B(n64372), .Z(n65228) );
  NOR U84661 ( .A(n69560), .B(n65228), .Z(n64374) );
  NOR U84662 ( .A(n64375), .B(n64374), .Z(n69561) );
  XOR U84663 ( .A(n69563), .B(n69561), .Z(n70334) );
  IV U84664 ( .A(n64376), .Z(n64377) );
  NOR U84665 ( .A(n64378), .B(n64377), .Z(n80222) );
  IV U84666 ( .A(n64379), .Z(n64381) );
  NOR U84667 ( .A(n64381), .B(n64380), .Z(n80229) );
  NOR U84668 ( .A(n80222), .B(n80229), .Z(n70336) );
  XOR U84669 ( .A(n70334), .B(n70336), .Z(n65223) );
  XOR U84670 ( .A(n64382), .B(n65223), .Z(n65227) );
  XOR U84671 ( .A(n64383), .B(n65227), .Z(n64387) );
  IV U84672 ( .A(n64387), .Z(n69575) );
  NOR U84673 ( .A(n64391), .B(n69575), .Z(n70323) );
  IV U84674 ( .A(n64384), .Z(n64385) );
  NOR U84675 ( .A(n64385), .B(n64390), .Z(n64386) );
  IV U84676 ( .A(n64386), .Z(n69574) );
  XOR U84677 ( .A(n64387), .B(n69574), .Z(n69577) );
  IV U84678 ( .A(n64388), .Z(n64389) );
  NOR U84679 ( .A(n64390), .B(n64389), .Z(n64392) );
  IV U84680 ( .A(n64392), .Z(n69576) );
  XOR U84681 ( .A(n69577), .B(n69576), .Z(n64394) );
  NOR U84682 ( .A(n64392), .B(n64391), .Z(n64393) );
  NOR U84683 ( .A(n64394), .B(n64393), .Z(n64395) );
  NOR U84684 ( .A(n70323), .B(n64395), .Z(n69579) );
  IV U84685 ( .A(n64396), .Z(n64398) );
  NOR U84686 ( .A(n64398), .B(n64397), .Z(n64399) );
  IV U84687 ( .A(n64399), .Z(n69581) );
  XOR U84688 ( .A(n69579), .B(n69581), .Z(n65215) );
  XOR U84689 ( .A(n65214), .B(n65215), .Z(n65218) );
  XOR U84690 ( .A(n65217), .B(n65218), .Z(n65209) );
  XOR U84691 ( .A(n65208), .B(n65209), .Z(n65213) );
  XOR U84692 ( .A(n65211), .B(n65213), .Z(n65202) );
  XOR U84693 ( .A(n65201), .B(n65202), .Z(n65205) );
  XOR U84694 ( .A(n65204), .B(n65205), .Z(n65199) );
  XOR U84695 ( .A(n65198), .B(n65199), .Z(n69588) );
  IV U84696 ( .A(n64400), .Z(n64401) );
  NOR U84697 ( .A(n64402), .B(n64401), .Z(n64403) );
  IV U84698 ( .A(n64403), .Z(n69587) );
  XOR U84699 ( .A(n69588), .B(n69587), .Z(n64408) );
  NOR U84700 ( .A(n64404), .B(n64409), .Z(n64405) );
  NOR U84701 ( .A(n64406), .B(n64405), .Z(n64407) );
  NOR U84702 ( .A(n64408), .B(n64407), .Z(n64418) );
  IV U84703 ( .A(n64409), .Z(n64413) );
  IV U84704 ( .A(n64410), .Z(n64411) );
  NOR U84705 ( .A(n64411), .B(n65199), .Z(n64412) );
  IV U84706 ( .A(n64412), .Z(n64414) );
  NOR U84707 ( .A(n64413), .B(n64414), .Z(n74882) );
  NOR U84708 ( .A(n64415), .B(n64414), .Z(n69591) );
  NOR U84709 ( .A(n74882), .B(n69591), .Z(n64416) );
  IV U84710 ( .A(n64416), .Z(n64417) );
  NOR U84711 ( .A(n64418), .B(n64417), .Z(n64419) );
  IV U84712 ( .A(n64419), .Z(n65197) );
  IV U84713 ( .A(n64420), .Z(n64423) );
  IV U84714 ( .A(n64421), .Z(n64422) );
  NOR U84715 ( .A(n64423), .B(n64422), .Z(n65195) );
  XOR U84716 ( .A(n65197), .B(n65195), .Z(n69600) );
  NOR U84717 ( .A(n69598), .B(n64424), .Z(n64428) );
  IV U84718 ( .A(n64425), .Z(n69601) );
  NOR U84719 ( .A(n64426), .B(n69601), .Z(n64427) );
  NOR U84720 ( .A(n64428), .B(n64427), .Z(n64429) );
  XOR U84721 ( .A(n69600), .B(n64429), .Z(n69607) );
  IV U84722 ( .A(n64430), .Z(n64432) );
  NOR U84723 ( .A(n64432), .B(n64431), .Z(n69608) );
  IV U84724 ( .A(n64433), .Z(n64435) );
  NOR U84725 ( .A(n64435), .B(n64434), .Z(n69610) );
  NOR U84726 ( .A(n69608), .B(n69610), .Z(n64436) );
  XOR U84727 ( .A(n69607), .B(n64436), .Z(n65189) );
  XOR U84728 ( .A(n65188), .B(n65189), .Z(n69614) );
  XOR U84729 ( .A(n69613), .B(n69614), .Z(n69621) );
  IV U84730 ( .A(n64437), .Z(n64439) );
  NOR U84731 ( .A(n64439), .B(n64438), .Z(n69616) );
  NOR U84732 ( .A(n64441), .B(n64440), .Z(n69620) );
  NOR U84733 ( .A(n69616), .B(n69620), .Z(n64442) );
  XOR U84734 ( .A(n69621), .B(n64442), .Z(n65183) );
  IV U84735 ( .A(n64443), .Z(n64444) );
  NOR U84736 ( .A(n64444), .B(n64449), .Z(n64445) );
  IV U84737 ( .A(n64445), .Z(n65184) );
  XOR U84738 ( .A(n65183), .B(n65184), .Z(n65187) );
  XOR U84739 ( .A(n65186), .B(n65187), .Z(n64452) );
  IV U84740 ( .A(n64452), .Z(n64446) );
  NOR U84741 ( .A(n64450), .B(n64446), .Z(n64447) );
  IV U84742 ( .A(n64447), .Z(n64448) );
  NOR U84743 ( .A(n64449), .B(n64448), .Z(n75624) );
  NOR U84744 ( .A(n64451), .B(n64450), .Z(n64453) );
  NOR U84745 ( .A(n64453), .B(n64452), .Z(n64454) );
  NOR U84746 ( .A(n75624), .B(n64454), .Z(n65178) );
  IV U84747 ( .A(n64455), .Z(n64456) );
  NOR U84748 ( .A(n64456), .B(n64464), .Z(n65179) );
  IV U84749 ( .A(n64457), .Z(n64458) );
  NOR U84750 ( .A(n64459), .B(n64458), .Z(n65181) );
  NOR U84751 ( .A(n69623), .B(n65181), .Z(n64460) );
  IV U84752 ( .A(n64460), .Z(n64461) );
  NOR U84753 ( .A(n65179), .B(n64461), .Z(n64462) );
  XOR U84754 ( .A(n65178), .B(n64462), .Z(n65175) );
  IV U84755 ( .A(n64463), .Z(n64465) );
  NOR U84756 ( .A(n64465), .B(n64464), .Z(n65173) );
  XOR U84757 ( .A(n65175), .B(n65173), .Z(n69630) );
  XOR U84758 ( .A(n64466), .B(n69630), .Z(n69636) );
  XOR U84759 ( .A(n69637), .B(n69636), .Z(n69644) );
  IV U84760 ( .A(n64467), .Z(n64468) );
  NOR U84761 ( .A(n64468), .B(n65165), .Z(n69633) );
  IV U84762 ( .A(n64469), .Z(n64474) );
  IV U84763 ( .A(n64470), .Z(n64471) );
  NOR U84764 ( .A(n64474), .B(n64471), .Z(n69643) );
  IV U84765 ( .A(n64472), .Z(n64473) );
  NOR U84766 ( .A(n64474), .B(n64473), .Z(n69639) );
  NOR U84767 ( .A(n69643), .B(n69639), .Z(n64475) );
  IV U84768 ( .A(n64475), .Z(n64476) );
  NOR U84769 ( .A(n69633), .B(n64476), .Z(n64477) );
  XOR U84770 ( .A(n69644), .B(n64477), .Z(n64478) );
  IV U84771 ( .A(n64478), .Z(n65166) );
  NOR U84772 ( .A(n64479), .B(n65165), .Z(n64480) );
  XOR U84773 ( .A(n65166), .B(n64480), .Z(n69655) );
  XOR U84774 ( .A(n69653), .B(n69655), .Z(n65158) );
  XOR U84775 ( .A(n64481), .B(n65158), .Z(n65152) );
  XOR U84776 ( .A(n65151), .B(n65152), .Z(n65155) );
  XOR U84777 ( .A(n65154), .B(n65155), .Z(n69662) );
  XOR U84778 ( .A(n69661), .B(n69662), .Z(n65146) );
  XOR U84779 ( .A(n64482), .B(n65146), .Z(n65141) );
  XOR U84780 ( .A(n65142), .B(n65141), .Z(n65139) );
  IV U84781 ( .A(n64483), .Z(n64488) );
  IV U84782 ( .A(n64484), .Z(n64485) );
  NOR U84783 ( .A(n64488), .B(n64485), .Z(n65137) );
  XOR U84784 ( .A(n65139), .B(n65137), .Z(n69671) );
  IV U84785 ( .A(n64486), .Z(n64487) );
  NOR U84786 ( .A(n64488), .B(n64487), .Z(n69669) );
  XOR U84787 ( .A(n69671), .B(n69669), .Z(n69678) );
  IV U84788 ( .A(n64489), .Z(n64490) );
  NOR U84789 ( .A(n64491), .B(n64490), .Z(n69672) );
  IV U84790 ( .A(n64492), .Z(n64493) );
  NOR U84791 ( .A(n64493), .B(n64496), .Z(n69676) );
  NOR U84792 ( .A(n69672), .B(n69676), .Z(n64494) );
  XOR U84793 ( .A(n69678), .B(n64494), .Z(n69681) );
  IV U84794 ( .A(n64495), .Z(n64497) );
  NOR U84795 ( .A(n64497), .B(n64496), .Z(n64498) );
  IV U84796 ( .A(n64498), .Z(n69682) );
  XOR U84797 ( .A(n69681), .B(n69682), .Z(n65136) );
  XOR U84798 ( .A(n65134), .B(n65136), .Z(n65132) );
  XOR U84799 ( .A(n65131), .B(n65132), .Z(n65127) );
  XOR U84800 ( .A(n64499), .B(n65127), .Z(n64500) );
  IV U84801 ( .A(n64500), .Z(n65125) );
  XOR U84802 ( .A(n64501), .B(n65125), .Z(n69692) );
  XOR U84803 ( .A(n69690), .B(n69692), .Z(n69694) );
  XOR U84804 ( .A(n69693), .B(n69694), .Z(n65115) );
  IV U84805 ( .A(n64502), .Z(n64504) );
  NOR U84806 ( .A(n64504), .B(n64503), .Z(n65113) );
  XOR U84807 ( .A(n65115), .B(n65113), .Z(n69704) );
  IV U84808 ( .A(n64505), .Z(n64507) );
  IV U84809 ( .A(n64506), .Z(n64511) );
  NOR U84810 ( .A(n64507), .B(n64511), .Z(n65111) );
  NOR U84811 ( .A(n65111), .B(n64508), .Z(n64509) );
  XOR U84812 ( .A(n69704), .B(n64509), .Z(n69706) );
  IV U84813 ( .A(n64510), .Z(n64512) );
  NOR U84814 ( .A(n64512), .B(n64511), .Z(n64513) );
  IV U84815 ( .A(n64513), .Z(n69707) );
  XOR U84816 ( .A(n69706), .B(n69707), .Z(n69711) );
  XOR U84817 ( .A(n69709), .B(n69711), .Z(n65105) );
  XOR U84818 ( .A(n65103), .B(n65105), .Z(n65108) );
  XOR U84819 ( .A(n64514), .B(n65108), .Z(n65095) );
  NOR U84820 ( .A(n64516), .B(n64515), .Z(n64517) );
  IV U84821 ( .A(n64517), .Z(n64519) );
  NOR U84822 ( .A(n64519), .B(n64518), .Z(n65100) );
  NOR U84823 ( .A(n65096), .B(n65100), .Z(n64520) );
  XOR U84824 ( .A(n65095), .B(n64520), .Z(n65091) );
  XOR U84825 ( .A(n65090), .B(n65091), .Z(n69716) );
  XOR U84826 ( .A(n65093), .B(n69716), .Z(n65088) );
  XOR U84827 ( .A(n64521), .B(n65088), .Z(n64522) );
  IV U84828 ( .A(n64522), .Z(n69726) );
  XOR U84829 ( .A(n69724), .B(n69726), .Z(n69728) );
  XOR U84830 ( .A(n69727), .B(n69728), .Z(n69737) );
  IV U84831 ( .A(n64523), .Z(n64524) );
  NOR U84832 ( .A(n64525), .B(n64524), .Z(n69736) );
  IV U84833 ( .A(n64526), .Z(n64527) );
  NOR U84834 ( .A(n64528), .B(n64527), .Z(n69734) );
  NOR U84835 ( .A(n69736), .B(n69734), .Z(n64529) );
  XOR U84836 ( .A(n69737), .B(n64529), .Z(n65083) );
  XOR U84837 ( .A(n64530), .B(n65083), .Z(n69745) );
  IV U84838 ( .A(n64531), .Z(n64533) );
  NOR U84839 ( .A(n64533), .B(n64532), .Z(n69742) );
  IV U84840 ( .A(n64534), .Z(n64535) );
  NOR U84841 ( .A(n64535), .B(n64541), .Z(n69744) );
  NOR U84842 ( .A(n69742), .B(n69744), .Z(n64536) );
  XOR U84843 ( .A(n69745), .B(n64536), .Z(n65080) );
  IV U84844 ( .A(n64537), .Z(n64538) );
  NOR U84845 ( .A(n64539), .B(n64538), .Z(n69753) );
  IV U84846 ( .A(n64540), .Z(n64542) );
  NOR U84847 ( .A(n64542), .B(n64541), .Z(n69752) );
  NOR U84848 ( .A(n69753), .B(n69752), .Z(n65081) );
  XOR U84849 ( .A(n65080), .B(n65081), .Z(n75496) );
  IV U84850 ( .A(n64543), .Z(n64545) );
  NOR U84851 ( .A(n64545), .B(n64544), .Z(n75492) );
  IV U84852 ( .A(n64546), .Z(n64548) );
  NOR U84853 ( .A(n64548), .B(n64547), .Z(n80385) );
  NOR U84854 ( .A(n75492), .B(n80385), .Z(n69761) );
  XOR U84855 ( .A(n75496), .B(n69761), .Z(n64549) );
  IV U84856 ( .A(n64549), .Z(n69764) );
  XOR U84857 ( .A(n69762), .B(n69764), .Z(n69768) );
  XOR U84858 ( .A(n64550), .B(n69768), .Z(n65072) );
  XOR U84859 ( .A(n65073), .B(n65072), .Z(n65076) );
  IV U84860 ( .A(n64551), .Z(n64552) );
  NOR U84861 ( .A(n64552), .B(n64554), .Z(n65075) );
  IV U84862 ( .A(n64553), .Z(n64555) );
  NOR U84863 ( .A(n64555), .B(n64554), .Z(n65070) );
  NOR U84864 ( .A(n65075), .B(n65070), .Z(n64556) );
  XOR U84865 ( .A(n65076), .B(n64556), .Z(n69771) );
  XOR U84866 ( .A(n69772), .B(n69771), .Z(n69775) );
  XOR U84867 ( .A(n69774), .B(n69775), .Z(n75022) );
  XOR U84868 ( .A(n65069), .B(n75022), .Z(n69781) );
  IV U84869 ( .A(n64557), .Z(n64558) );
  NOR U84870 ( .A(n70178), .B(n64558), .Z(n69780) );
  IV U84871 ( .A(n64559), .Z(n64561) );
  NOR U84872 ( .A(n64561), .B(n64560), .Z(n69783) );
  NOR U84873 ( .A(n69780), .B(n69783), .Z(n64562) );
  XOR U84874 ( .A(n69781), .B(n64562), .Z(n69792) );
  XOR U84875 ( .A(n65067), .B(n69792), .Z(n64563) );
  NOR U84876 ( .A(n64571), .B(n64563), .Z(n70159) );
  IV U84877 ( .A(n64564), .Z(n64565) );
  NOR U84878 ( .A(n64566), .B(n64565), .Z(n69791) );
  NOR U84879 ( .A(n65067), .B(n69791), .Z(n64567) );
  XOR U84880 ( .A(n64567), .B(n69792), .Z(n64568) );
  IV U84881 ( .A(n64568), .Z(n65066) );
  IV U84882 ( .A(n64569), .Z(n64570) );
  NOR U84883 ( .A(n64578), .B(n64570), .Z(n64572) );
  IV U84884 ( .A(n64572), .Z(n65065) );
  XOR U84885 ( .A(n65066), .B(n65065), .Z(n64574) );
  NOR U84886 ( .A(n64572), .B(n64571), .Z(n64573) );
  NOR U84887 ( .A(n64574), .B(n64573), .Z(n64575) );
  NOR U84888 ( .A(n70159), .B(n64575), .Z(n65058) );
  IV U84889 ( .A(n64583), .Z(n64576) );
  NOR U84890 ( .A(n64582), .B(n64576), .Z(n65060) );
  IV U84891 ( .A(n64577), .Z(n64579) );
  NOR U84892 ( .A(n64579), .B(n64578), .Z(n65062) );
  NOR U84893 ( .A(n65060), .B(n65062), .Z(n64580) );
  XOR U84894 ( .A(n65058), .B(n64580), .Z(n65057) );
  IV U84895 ( .A(n64581), .Z(n64585) );
  XOR U84896 ( .A(n64583), .B(n64582), .Z(n64584) );
  NOR U84897 ( .A(n64585), .B(n64584), .Z(n65055) );
  IV U84898 ( .A(n64586), .Z(n64588) );
  NOR U84899 ( .A(n64588), .B(n64587), .Z(n65053) );
  NOR U84900 ( .A(n65055), .B(n65053), .Z(n64589) );
  XOR U84901 ( .A(n65057), .B(n64589), .Z(n69797) );
  XOR U84902 ( .A(n69798), .B(n69797), .Z(n69800) );
  XOR U84903 ( .A(n69799), .B(n69800), .Z(n69810) );
  XOR U84904 ( .A(n64590), .B(n69810), .Z(n69804) );
  XOR U84905 ( .A(n64591), .B(n69804), .Z(n69818) );
  NOR U84906 ( .A(n64592), .B(n69818), .Z(n70135) );
  IV U84907 ( .A(n64593), .Z(n64594) );
  NOR U84908 ( .A(n64594), .B(n64595), .Z(n65045) );
  NOR U84909 ( .A(n64596), .B(n64595), .Z(n65048) );
  XOR U84910 ( .A(n65048), .B(n69818), .Z(n65046) );
  XOR U84911 ( .A(n65045), .B(n65046), .Z(n69825) );
  IV U84912 ( .A(n69825), .Z(n64597) );
  NOR U84913 ( .A(n64598), .B(n64597), .Z(n64599) );
  NOR U84914 ( .A(n70135), .B(n64599), .Z(n65041) );
  NOR U84915 ( .A(n64600), .B(n69826), .Z(n64604) );
  IV U84916 ( .A(n64601), .Z(n64602) );
  NOR U84917 ( .A(n64603), .B(n64602), .Z(n65040) );
  NOR U84918 ( .A(n64604), .B(n65040), .Z(n64605) );
  XOR U84919 ( .A(n65041), .B(n64605), .Z(n69837) );
  IV U84920 ( .A(n64606), .Z(n64608) );
  NOR U84921 ( .A(n64608), .B(n64607), .Z(n69835) );
  NOR U84922 ( .A(n64609), .B(n65037), .Z(n64610) );
  NOR U84923 ( .A(n69835), .B(n64610), .Z(n64611) );
  XOR U84924 ( .A(n69837), .B(n64611), .Z(n64612) );
  IV U84925 ( .A(n64612), .Z(n65034) );
  XOR U84926 ( .A(n65033), .B(n65034), .Z(n69843) );
  IV U84927 ( .A(n64613), .Z(n64615) );
  NOR U84928 ( .A(n64615), .B(n64614), .Z(n65031) );
  IV U84929 ( .A(n64616), .Z(n64618) );
  NOR U84930 ( .A(n64618), .B(n64617), .Z(n69842) );
  NOR U84931 ( .A(n65031), .B(n69842), .Z(n64619) );
  XOR U84932 ( .A(n69843), .B(n64619), .Z(n64620) );
  IV U84933 ( .A(n64620), .Z(n65028) );
  XOR U84934 ( .A(n65027), .B(n65028), .Z(n69840) );
  XOR U84935 ( .A(n69839), .B(n69840), .Z(n69850) );
  XOR U84936 ( .A(n69851), .B(n69850), .Z(n65025) );
  IV U84937 ( .A(n64621), .Z(n64622) );
  NOR U84938 ( .A(n64623), .B(n64622), .Z(n65024) );
  NOR U84939 ( .A(n69852), .B(n65024), .Z(n64624) );
  XOR U84940 ( .A(n65025), .B(n64624), .Z(n65021) );
  XOR U84941 ( .A(n65019), .B(n65021), .Z(n69858) );
  IV U84942 ( .A(n64625), .Z(n64627) );
  NOR U84943 ( .A(n64627), .B(n64626), .Z(n65022) );
  IV U84944 ( .A(n64628), .Z(n64629) );
  NOR U84945 ( .A(n64629), .B(n64633), .Z(n69856) );
  NOR U84946 ( .A(n65022), .B(n69856), .Z(n64630) );
  XOR U84947 ( .A(n69858), .B(n64630), .Z(n64631) );
  IV U84948 ( .A(n64631), .Z(n69864) );
  IV U84949 ( .A(n64632), .Z(n64634) );
  NOR U84950 ( .A(n64634), .B(n64633), .Z(n69862) );
  XOR U84951 ( .A(n69864), .B(n69862), .Z(n69866) );
  XOR U84952 ( .A(n64635), .B(n69866), .Z(n64643) );
  IV U84953 ( .A(n64643), .Z(n64636) );
  NOR U84954 ( .A(n64637), .B(n64636), .Z(n70110) );
  IV U84955 ( .A(n64638), .Z(n64640) );
  NOR U84956 ( .A(n64640), .B(n64639), .Z(n64644) );
  IV U84957 ( .A(n64644), .Z(n64642) );
  XOR U84958 ( .A(n69860), .B(n69866), .Z(n64641) );
  NOR U84959 ( .A(n64642), .B(n64641), .Z(n69874) );
  NOR U84960 ( .A(n64644), .B(n64643), .Z(n64645) );
  NOR U84961 ( .A(n69874), .B(n64645), .Z(n64650) );
  NOR U84962 ( .A(n64646), .B(n64650), .Z(n64647) );
  NOR U84963 ( .A(n70110), .B(n64647), .Z(n64648) );
  NOR U84964 ( .A(n64649), .B(n64648), .Z(n64653) );
  IV U84965 ( .A(n64649), .Z(n64652) );
  IV U84966 ( .A(n64650), .Z(n64651) );
  NOR U84967 ( .A(n64652), .B(n64651), .Z(n75140) );
  NOR U84968 ( .A(n64653), .B(n75140), .Z(n64654) );
  IV U84969 ( .A(n64654), .Z(n65016) );
  IV U84970 ( .A(n64655), .Z(n64657) );
  NOR U84971 ( .A(n64657), .B(n64656), .Z(n65015) );
  XOR U84972 ( .A(n65016), .B(n65015), .Z(n69878) );
  XOR U84973 ( .A(n64658), .B(n69878), .Z(n65011) );
  IV U84974 ( .A(n64659), .Z(n64661) );
  NOR U84975 ( .A(n64661), .B(n64660), .Z(n65010) );
  IV U84976 ( .A(n64662), .Z(n64663) );
  NOR U84977 ( .A(n64663), .B(n69890), .Z(n69886) );
  NOR U84978 ( .A(n65010), .B(n69886), .Z(n64664) );
  XOR U84979 ( .A(n65011), .B(n64664), .Z(n69896) );
  NOR U84980 ( .A(n64665), .B(n69895), .Z(n64669) );
  IV U84981 ( .A(n64666), .Z(n64667) );
  NOR U84982 ( .A(n64667), .B(n65001), .Z(n64668) );
  NOR U84983 ( .A(n64669), .B(n64668), .Z(n64670) );
  XOR U84984 ( .A(n69896), .B(n64670), .Z(n64998) );
  IV U84985 ( .A(n64671), .Z(n64673) );
  NOR U84986 ( .A(n64673), .B(n64672), .Z(n69900) );
  IV U84987 ( .A(n64674), .Z(n64676) );
  NOR U84988 ( .A(n64676), .B(n64675), .Z(n64997) );
  NOR U84989 ( .A(n69900), .B(n64997), .Z(n64677) );
  XOR U84990 ( .A(n64998), .B(n64677), .Z(n75180) );
  IV U84991 ( .A(n64678), .Z(n64680) );
  NOR U84992 ( .A(n64680), .B(n64679), .Z(n75178) );
  IV U84993 ( .A(n64681), .Z(n64682) );
  NOR U84994 ( .A(n64682), .B(n64684), .Z(n75184) );
  NOR U84995 ( .A(n75178), .B(n75184), .Z(n64992) );
  XOR U84996 ( .A(n75180), .B(n64992), .Z(n64986) );
  IV U84997 ( .A(n64683), .Z(n64685) );
  NOR U84998 ( .A(n64685), .B(n64684), .Z(n64993) );
  IV U84999 ( .A(n64686), .Z(n64688) );
  NOR U85000 ( .A(n64688), .B(n64687), .Z(n64985) );
  NOR U85001 ( .A(n64993), .B(n64985), .Z(n64689) );
  XOR U85002 ( .A(n64986), .B(n64689), .Z(n64989) );
  NOR U85003 ( .A(n64696), .B(n64989), .Z(n75195) );
  IV U85004 ( .A(n64690), .Z(n64692) );
  NOR U85005 ( .A(n64692), .B(n64691), .Z(n64982) );
  IV U85006 ( .A(n64693), .Z(n64695) );
  NOR U85007 ( .A(n64695), .B(n64694), .Z(n64988) );
  XOR U85008 ( .A(n64988), .B(n64989), .Z(n64983) );
  IV U85009 ( .A(n64983), .Z(n64697) );
  XOR U85010 ( .A(n64982), .B(n64697), .Z(n64699) );
  NOR U85011 ( .A(n64697), .B(n64696), .Z(n64698) );
  NOR U85012 ( .A(n64699), .B(n64698), .Z(n64700) );
  NOR U85013 ( .A(n75195), .B(n64700), .Z(n64701) );
  IV U85014 ( .A(n64701), .Z(n64977) );
  XOR U85015 ( .A(n64976), .B(n64977), .Z(n70098) );
  IV U85016 ( .A(n70098), .Z(n64710) );
  IV U85017 ( .A(n64702), .Z(n64703) );
  NOR U85018 ( .A(n64704), .B(n64703), .Z(n64979) );
  IV U85019 ( .A(n64705), .Z(n64707) );
  NOR U85020 ( .A(n64707), .B(n64706), .Z(n70102) );
  NOR U85021 ( .A(n70102), .B(n70097), .Z(n64975) );
  IV U85022 ( .A(n64975), .Z(n64708) );
  NOR U85023 ( .A(n64979), .B(n64708), .Z(n64709) );
  XOR U85024 ( .A(n64710), .B(n64709), .Z(n64973) );
  XOR U85025 ( .A(n64971), .B(n64973), .Z(n64968) );
  IV U85026 ( .A(n64711), .Z(n64713) );
  NOR U85027 ( .A(n64713), .B(n64712), .Z(n69915) );
  IV U85028 ( .A(n64714), .Z(n64716) );
  IV U85029 ( .A(n64715), .Z(n64718) );
  NOR U85030 ( .A(n64716), .B(n64718), .Z(n64967) );
  IV U85031 ( .A(n64717), .Z(n64719) );
  NOR U85032 ( .A(n64719), .B(n64718), .Z(n64972) );
  NOR U85033 ( .A(n64967), .B(n64972), .Z(n64720) );
  IV U85034 ( .A(n64720), .Z(n64721) );
  NOR U85035 ( .A(n69915), .B(n64721), .Z(n64722) );
  XOR U85036 ( .A(n64968), .B(n64722), .Z(n69914) );
  XOR U85037 ( .A(n69912), .B(n69914), .Z(n69925) );
  IV U85038 ( .A(n64723), .Z(n64724) );
  NOR U85039 ( .A(n64725), .B(n64724), .Z(n64962) );
  NOR U85040 ( .A(n69926), .B(n64962), .Z(n64726) );
  XOR U85041 ( .A(n69925), .B(n64726), .Z(n64727) );
  IV U85042 ( .A(n64727), .Z(n64960) );
  NOR U85043 ( .A(n64734), .B(n64960), .Z(n70082) );
  IV U85044 ( .A(n64728), .Z(n64730) );
  NOR U85045 ( .A(n64730), .B(n64729), .Z(n64956) );
  IV U85046 ( .A(n64731), .Z(n64732) );
  NOR U85047 ( .A(n64733), .B(n64732), .Z(n64959) );
  XOR U85048 ( .A(n64959), .B(n64960), .Z(n64957) );
  IV U85049 ( .A(n64957), .Z(n64735) );
  XOR U85050 ( .A(n64956), .B(n64735), .Z(n64737) );
  NOR U85051 ( .A(n64735), .B(n64734), .Z(n64736) );
  NOR U85052 ( .A(n64737), .B(n64736), .Z(n64738) );
  NOR U85053 ( .A(n70082), .B(n64738), .Z(n69944) );
  XOR U85054 ( .A(n64739), .B(n69944), .Z(n69949) );
  IV U85055 ( .A(n64740), .Z(n64741) );
  NOR U85056 ( .A(n64742), .B(n64741), .Z(n64954) );
  IV U85057 ( .A(n64743), .Z(n64745) );
  NOR U85058 ( .A(n64745), .B(n64744), .Z(n69947) );
  NOR U85059 ( .A(n64954), .B(n69947), .Z(n64746) );
  XOR U85060 ( .A(n69949), .B(n64746), .Z(n64947) );
  XOR U85061 ( .A(n64949), .B(n64947), .Z(n64951) );
  XOR U85062 ( .A(n64950), .B(n64951), .Z(n69957) );
  IV U85063 ( .A(n69957), .Z(n64758) );
  IV U85064 ( .A(n64747), .Z(n64749) );
  IV U85065 ( .A(n64748), .Z(n64753) );
  NOR U85066 ( .A(n64749), .B(n64753), .Z(n69955) );
  IV U85067 ( .A(n64750), .Z(n64752) );
  NOR U85068 ( .A(n64752), .B(n64751), .Z(n64945) );
  NOR U85069 ( .A(n64754), .B(n64753), .Z(n64943) );
  NOR U85070 ( .A(n64945), .B(n64943), .Z(n64755) );
  IV U85071 ( .A(n64755), .Z(n64756) );
  NOR U85072 ( .A(n69955), .B(n64756), .Z(n64757) );
  XOR U85073 ( .A(n64758), .B(n64757), .Z(n69960) );
  IV U85074 ( .A(n64759), .Z(n64761) );
  NOR U85075 ( .A(n64761), .B(n64760), .Z(n69958) );
  XOR U85076 ( .A(n69960), .B(n69958), .Z(n69962) );
  IV U85077 ( .A(n64762), .Z(n64763) );
  NOR U85078 ( .A(n64764), .B(n64763), .Z(n69961) );
  IV U85079 ( .A(n64765), .Z(n64767) );
  NOR U85080 ( .A(n64767), .B(n64766), .Z(n64941) );
  NOR U85081 ( .A(n69961), .B(n64941), .Z(n64768) );
  XOR U85082 ( .A(n69962), .B(n64768), .Z(n64932) );
  IV U85083 ( .A(n64769), .Z(n64770) );
  NOR U85084 ( .A(n64770), .B(n64772), .Z(n64938) );
  IV U85085 ( .A(n64771), .Z(n64773) );
  NOR U85086 ( .A(n64773), .B(n64772), .Z(n64933) );
  NOR U85087 ( .A(n64938), .B(n64933), .Z(n64774) );
  XOR U85088 ( .A(n64932), .B(n64774), .Z(n64936) );
  IV U85089 ( .A(n64775), .Z(n64777) );
  NOR U85090 ( .A(n64777), .B(n64776), .Z(n64930) );
  NOR U85091 ( .A(n64935), .B(n64930), .Z(n64778) );
  XOR U85092 ( .A(n64936), .B(n64778), .Z(n64911) );
  NOR U85093 ( .A(n64779), .B(n64923), .Z(n64912) );
  IV U85094 ( .A(n64780), .Z(n64781) );
  NOR U85095 ( .A(n64782), .B(n64781), .Z(n64920) );
  NOR U85096 ( .A(n64912), .B(n64920), .Z(n64783) );
  XOR U85097 ( .A(n64911), .B(n64783), .Z(n64909) );
  NOR U85098 ( .A(n64784), .B(n64913), .Z(n64787) );
  IV U85099 ( .A(n64785), .Z(n64786) );
  NOR U85100 ( .A(n64786), .B(n64791), .Z(n64907) );
  NOR U85101 ( .A(n64787), .B(n64907), .Z(n64788) );
  XOR U85102 ( .A(n64909), .B(n64788), .Z(n64789) );
  IV U85103 ( .A(n64789), .Z(n64906) );
  IV U85104 ( .A(n64790), .Z(n64792) );
  NOR U85105 ( .A(n64792), .B(n64791), .Z(n64904) );
  XOR U85106 ( .A(n64906), .B(n64904), .Z(n64899) );
  XOR U85107 ( .A(n64898), .B(n64899), .Z(n64902) );
  NOR U85108 ( .A(n64799), .B(n64902), .Z(n70051) );
  IV U85109 ( .A(n64793), .Z(n64795) );
  NOR U85110 ( .A(n64795), .B(n64794), .Z(n64895) );
  IV U85111 ( .A(n64796), .Z(n64797) );
  NOR U85112 ( .A(n64798), .B(n64797), .Z(n64901) );
  XOR U85113 ( .A(n64901), .B(n64902), .Z(n64896) );
  IV U85114 ( .A(n64896), .Z(n64800) );
  XOR U85115 ( .A(n64895), .B(n64800), .Z(n64802) );
  NOR U85116 ( .A(n64800), .B(n64799), .Z(n64801) );
  NOR U85117 ( .A(n64802), .B(n64801), .Z(n64803) );
  NOR U85118 ( .A(n70051), .B(n64803), .Z(n64804) );
  IV U85119 ( .A(n64804), .Z(n64891) );
  XOR U85120 ( .A(n64890), .B(n64891), .Z(n69972) );
  IV U85121 ( .A(n64805), .Z(n64807) );
  NOR U85122 ( .A(n64807), .B(n64806), .Z(n64893) );
  IV U85123 ( .A(n64808), .Z(n64809) );
  NOR U85124 ( .A(n64810), .B(n64809), .Z(n69971) );
  NOR U85125 ( .A(n64893), .B(n69971), .Z(n64811) );
  XOR U85126 ( .A(n69972), .B(n64811), .Z(n64812) );
  IV U85127 ( .A(n64812), .Z(n69970) );
  IV U85128 ( .A(n64813), .Z(n64815) );
  NOR U85129 ( .A(n64815), .B(n64814), .Z(n64816) );
  IV U85130 ( .A(n64816), .Z(n64823) );
  NOR U85131 ( .A(n69970), .B(n64823), .Z(n75299) );
  IV U85132 ( .A(n64817), .Z(n64819) );
  NOR U85133 ( .A(n64819), .B(n64818), .Z(n64887) );
  IV U85134 ( .A(n64820), .Z(n64822) );
  NOR U85135 ( .A(n64822), .B(n64821), .Z(n69968) );
  XOR U85136 ( .A(n69968), .B(n69970), .Z(n64888) );
  IV U85137 ( .A(n64888), .Z(n64824) );
  XOR U85138 ( .A(n64887), .B(n64824), .Z(n64826) );
  NOR U85139 ( .A(n64824), .B(n64823), .Z(n64825) );
  NOR U85140 ( .A(n64826), .B(n64825), .Z(n64827) );
  NOR U85141 ( .A(n75299), .B(n64827), .Z(n64828) );
  IV U85142 ( .A(n64828), .Z(n69978) );
  XOR U85143 ( .A(n69977), .B(n69978), .Z(n64884) );
  XOR U85144 ( .A(n64883), .B(n64884), .Z(n69986) );
  IV U85145 ( .A(n64829), .Z(n64831) );
  NOR U85146 ( .A(n64831), .B(n64830), .Z(n69975) );
  IV U85147 ( .A(n64832), .Z(n64834) );
  NOR U85148 ( .A(n64834), .B(n64833), .Z(n69985) );
  NOR U85149 ( .A(n69975), .B(n69985), .Z(n64835) );
  XOR U85150 ( .A(n69986), .B(n64835), .Z(n64872) );
  XOR U85151 ( .A(n64836), .B(n64872), .Z(n70003) );
  XOR U85152 ( .A(n64837), .B(n70003), .Z(n64867) );
  XOR U85153 ( .A(n64868), .B(n64867), .Z(n64851) );
  XOR U85154 ( .A(n64839), .B(n64838), .Z(n80645) );
  XOR U85155 ( .A(n70010), .B(n70012), .Z(n64840) );
  NOR U85156 ( .A(n80645), .B(n64840), .Z(n64841) );
  IV U85157 ( .A(n64841), .Z(n64863) );
  IV U85158 ( .A(n64842), .Z(n64844) );
  NOR U85159 ( .A(n64844), .B(n64843), .Z(n70007) );
  IV U85160 ( .A(n70007), .Z(n64845) );
  NOR U85161 ( .A(n64863), .B(n64845), .Z(n64858) );
  IV U85162 ( .A(n64858), .Z(n64848) );
  XOR U85163 ( .A(n64847), .B(n64846), .Z(n64857) );
  NOR U85164 ( .A(n64848), .B(n64857), .Z(n64853) );
  IV U85165 ( .A(n64853), .Z(n64849) );
  NOR U85166 ( .A(n64856), .B(n64849), .Z(n64852) );
  IV U85167 ( .A(n64852), .Z(n64850) );
  NOR U85168 ( .A(n64851), .B(n64850), .Z(n80632) );
  XOR U85169 ( .A(n64852), .B(n64851), .Z(n70004) );
  NOR U85170 ( .A(n64854), .B(n64853), .Z(n64855) );
  XOR U85171 ( .A(n64856), .B(n64855), .Z(n75327) );
  IV U85172 ( .A(n75327), .Z(n70023) );
  XOR U85173 ( .A(n64858), .B(n64857), .Z(n70015) );
  IV U85174 ( .A(n64859), .Z(n64861) );
  NOR U85175 ( .A(n64861), .B(n64860), .Z(n70006) );
  IV U85176 ( .A(n70006), .Z(n64862) );
  NOR U85177 ( .A(n64863), .B(n64862), .Z(n70016) );
  IV U85178 ( .A(n70016), .Z(n64864) );
  NOR U85179 ( .A(n70015), .B(n64864), .Z(n75326) );
  IV U85180 ( .A(n75326), .Z(n64865) );
  NOR U85181 ( .A(n70023), .B(n64865), .Z(n70005) );
  IV U85182 ( .A(n70005), .Z(n64866) );
  NOR U85183 ( .A(n70004), .B(n64866), .Z(n75334) );
  NOR U85184 ( .A(n80632), .B(n75334), .Z(n70029) );
  IV U85185 ( .A(n64867), .Z(n64869) );
  NOR U85186 ( .A(n64869), .B(n64868), .Z(n70026) );
  IV U85187 ( .A(n64870), .Z(n64871) );
  NOR U85188 ( .A(n70003), .B(n64871), .Z(n70032) );
  IV U85189 ( .A(n64872), .Z(n64877) );
  IV U85190 ( .A(n64873), .Z(n64874) );
  NOR U85191 ( .A(n64877), .B(n64874), .Z(n64875) );
  IV U85192 ( .A(n64875), .Z(n70040) );
  IV U85193 ( .A(n64876), .Z(n64878) );
  NOR U85194 ( .A(n64878), .B(n64877), .Z(n75308) );
  IV U85195 ( .A(n64879), .Z(n64880) );
  XOR U85196 ( .A(n69975), .B(n69986), .Z(n69989) );
  NOR U85197 ( .A(n64880), .B(n69989), .Z(n64881) );
  IV U85198 ( .A(n64881), .Z(n64882) );
  NOR U85199 ( .A(n69991), .B(n64882), .Z(n75310) );
  NOR U85200 ( .A(n75308), .B(n75310), .Z(n70000) );
  IV U85201 ( .A(n64883), .Z(n64885) );
  NOR U85202 ( .A(n64885), .B(n64884), .Z(n64886) );
  IV U85203 ( .A(n64886), .Z(n69981) );
  IV U85204 ( .A(n64887), .Z(n64889) );
  NOR U85205 ( .A(n64889), .B(n64888), .Z(n75302) );
  IV U85206 ( .A(n64890), .Z(n64892) );
  NOR U85207 ( .A(n64892), .B(n64891), .Z(n80710) );
  IV U85208 ( .A(n64893), .Z(n64894) );
  NOR U85209 ( .A(n64894), .B(n69972), .Z(n80702) );
  NOR U85210 ( .A(n80710), .B(n80702), .Z(n70050) );
  IV U85211 ( .A(n64895), .Z(n64897) );
  NOR U85212 ( .A(n64897), .B(n64896), .Z(n75280) );
  IV U85213 ( .A(n64898), .Z(n64900) );
  NOR U85214 ( .A(n64900), .B(n64899), .Z(n75270) );
  IV U85215 ( .A(n64901), .Z(n64903) );
  NOR U85216 ( .A(n64903), .B(n64902), .Z(n75276) );
  NOR U85217 ( .A(n75270), .B(n75276), .Z(n69967) );
  IV U85218 ( .A(n64904), .Z(n64905) );
  NOR U85219 ( .A(n64906), .B(n64905), .Z(n75272) );
  IV U85220 ( .A(n64907), .Z(n64908) );
  NOR U85221 ( .A(n64909), .B(n64908), .Z(n70054) );
  NOR U85222 ( .A(n75272), .B(n70054), .Z(n69966) );
  IV U85223 ( .A(n64910), .Z(n64916) );
  IV U85224 ( .A(n64911), .Z(n64924) );
  XOR U85225 ( .A(n64912), .B(n64924), .Z(n64914) );
  NOR U85226 ( .A(n64914), .B(n64913), .Z(n64915) );
  IV U85227 ( .A(n64915), .Z(n64918) );
  NOR U85228 ( .A(n64916), .B(n64918), .Z(n75260) );
  IV U85229 ( .A(n64917), .Z(n64919) );
  NOR U85230 ( .A(n64919), .B(n64918), .Z(n75257) );
  IV U85231 ( .A(n64920), .Z(n64921) );
  NOR U85232 ( .A(n64924), .B(n64921), .Z(n75252) );
  IV U85233 ( .A(n64922), .Z(n64926) );
  NOR U85234 ( .A(n64924), .B(n64923), .Z(n64925) );
  IV U85235 ( .A(n64925), .Z(n64928) );
  NOR U85236 ( .A(n64926), .B(n64928), .Z(n75249) );
  IV U85237 ( .A(n64927), .Z(n64929) );
  NOR U85238 ( .A(n64929), .B(n64928), .Z(n70059) );
  IV U85239 ( .A(n64930), .Z(n64931) );
  NOR U85240 ( .A(n64931), .B(n64936), .Z(n70056) );
  IV U85241 ( .A(n64932), .Z(n64940) );
  IV U85242 ( .A(n64933), .Z(n64934) );
  NOR U85243 ( .A(n64940), .B(n64934), .Z(n75349) );
  IV U85244 ( .A(n64935), .Z(n64937) );
  NOR U85245 ( .A(n64937), .B(n64936), .Z(n80537) );
  NOR U85246 ( .A(n75349), .B(n80537), .Z(n70065) );
  IV U85247 ( .A(n70065), .Z(n69965) );
  IV U85248 ( .A(n64938), .Z(n64939) );
  NOR U85249 ( .A(n64940), .B(n64939), .Z(n70062) );
  IV U85250 ( .A(n64941), .Z(n64942) );
  NOR U85251 ( .A(n64942), .B(n69962), .Z(n75243) );
  NOR U85252 ( .A(n70062), .B(n75243), .Z(n69964) );
  IV U85253 ( .A(n64943), .Z(n64944) );
  NOR U85254 ( .A(n64944), .B(n69957), .Z(n75236) );
  IV U85255 ( .A(n64945), .Z(n64946) );
  NOR U85256 ( .A(n64946), .B(n69957), .Z(n70068) );
  IV U85257 ( .A(n64947), .Z(n64948) );
  NOR U85258 ( .A(n64949), .B(n64948), .Z(n70071) );
  IV U85259 ( .A(n64950), .Z(n64952) );
  NOR U85260 ( .A(n64952), .B(n64951), .Z(n70066) );
  NOR U85261 ( .A(n70071), .B(n70066), .Z(n64953) );
  IV U85262 ( .A(n64953), .Z(n69954) );
  IV U85263 ( .A(n64954), .Z(n64955) );
  NOR U85264 ( .A(n69949), .B(n64955), .Z(n70074) );
  IV U85265 ( .A(n64956), .Z(n64958) );
  NOR U85266 ( .A(n64958), .B(n64957), .Z(n70085) );
  IV U85267 ( .A(n64959), .Z(n64961) );
  NOR U85268 ( .A(n64961), .B(n64960), .Z(n75215) );
  IV U85269 ( .A(n64962), .Z(n64963) );
  NOR U85270 ( .A(n64963), .B(n69925), .Z(n64964) );
  IV U85271 ( .A(n64964), .Z(n64965) );
  NOR U85272 ( .A(n69930), .B(n64965), .Z(n75212) );
  IV U85273 ( .A(n69926), .Z(n64966) );
  NOR U85274 ( .A(n64966), .B(n69925), .Z(n69920) );
  IV U85275 ( .A(n64967), .Z(n64969) );
  IV U85276 ( .A(n64968), .Z(n69916) );
  NOR U85277 ( .A(n64969), .B(n69916), .Z(n64970) );
  IV U85278 ( .A(n64970), .Z(n70089) );
  NOR U85279 ( .A(n64971), .B(n64973), .Z(n70091) );
  IV U85280 ( .A(n64972), .Z(n64974) );
  NOR U85281 ( .A(n64974), .B(n64973), .Z(n70093) );
  NOR U85282 ( .A(n70091), .B(n70093), .Z(n69911) );
  NOR U85283 ( .A(n64975), .B(n70098), .Z(n69910) );
  IV U85284 ( .A(n64976), .Z(n64978) );
  NOR U85285 ( .A(n64978), .B(n64977), .Z(n75198) );
  IV U85286 ( .A(n64979), .Z(n64980) );
  NOR U85287 ( .A(n64980), .B(n70098), .Z(n70105) );
  NOR U85288 ( .A(n75198), .B(n70105), .Z(n64981) );
  IV U85289 ( .A(n64981), .Z(n69909) );
  IV U85290 ( .A(n64982), .Z(n64984) );
  NOR U85291 ( .A(n64984), .B(n64983), .Z(n75193) );
  IV U85292 ( .A(n64985), .Z(n64987) );
  IV U85293 ( .A(n64986), .Z(n64994) );
  NOR U85294 ( .A(n64987), .B(n64994), .Z(n80494) );
  IV U85295 ( .A(n64988), .Z(n64990) );
  NOR U85296 ( .A(n64990), .B(n64989), .Z(n80500) );
  NOR U85297 ( .A(n80494), .B(n80500), .Z(n70109) );
  IV U85298 ( .A(n70109), .Z(n64991) );
  NOR U85299 ( .A(n64991), .B(n75195), .Z(n69908) );
  NOR U85300 ( .A(n75180), .B(n64992), .Z(n64996) );
  IV U85301 ( .A(n64993), .Z(n64995) );
  NOR U85302 ( .A(n64995), .B(n64994), .Z(n75187) );
  NOR U85303 ( .A(n64996), .B(n75187), .Z(n69907) );
  IV U85304 ( .A(n64997), .Z(n64999) );
  IV U85305 ( .A(n64998), .Z(n69901) );
  NOR U85306 ( .A(n64999), .B(n69901), .Z(n75176) );
  IV U85307 ( .A(n65000), .Z(n65009) );
  NOR U85308 ( .A(n69896), .B(n65001), .Z(n65002) );
  IV U85309 ( .A(n65002), .Z(n65007) );
  NOR U85310 ( .A(n65004), .B(n65003), .Z(n65005) );
  IV U85311 ( .A(n65005), .Z(n65006) );
  NOR U85312 ( .A(n65007), .B(n65006), .Z(n65008) );
  IV U85313 ( .A(n65008), .Z(n69904) );
  NOR U85314 ( .A(n65009), .B(n69904), .Z(n75170) );
  IV U85315 ( .A(n65010), .Z(n65012) );
  IV U85316 ( .A(n65011), .Z(n69887) );
  NOR U85317 ( .A(n65012), .B(n69887), .Z(n75155) );
  IV U85318 ( .A(n65013), .Z(n65014) );
  NOR U85319 ( .A(n65014), .B(n69878), .Z(n75151) );
  IV U85320 ( .A(n65015), .Z(n65017) );
  NOR U85321 ( .A(n65017), .B(n65016), .Z(n65018) );
  IV U85322 ( .A(n65018), .Z(n69880) );
  IV U85323 ( .A(n65019), .Z(n65020) );
  NOR U85324 ( .A(n65021), .B(n65020), .Z(n75434) );
  IV U85325 ( .A(n65022), .Z(n65023) );
  NOR U85326 ( .A(n65023), .B(n69858), .Z(n75426) );
  NOR U85327 ( .A(n75434), .B(n75426), .Z(n70114) );
  IV U85328 ( .A(n65024), .Z(n65026) );
  IV U85329 ( .A(n65025), .Z(n69853) );
  NOR U85330 ( .A(n65026), .B(n69853), .Z(n75108) );
  IV U85331 ( .A(n65027), .Z(n65029) );
  NOR U85332 ( .A(n65029), .B(n65028), .Z(n65030) );
  IV U85333 ( .A(n65030), .Z(n69845) );
  IV U85334 ( .A(n65031), .Z(n65032) );
  NOR U85335 ( .A(n65032), .B(n69843), .Z(n75099) );
  IV U85336 ( .A(n65033), .Z(n65035) );
  NOR U85337 ( .A(n65035), .B(n65034), .Z(n75096) );
  IV U85338 ( .A(n65036), .Z(n65039) );
  NOR U85339 ( .A(n69837), .B(n65037), .Z(n65038) );
  IV U85340 ( .A(n65038), .Z(n69833) );
  NOR U85341 ( .A(n65039), .B(n69833), .Z(n70129) );
  IV U85342 ( .A(n65040), .Z(n65043) );
  IV U85343 ( .A(n65041), .Z(n65042) );
  NOR U85344 ( .A(n65043), .B(n65042), .Z(n65044) );
  IV U85345 ( .A(n65044), .Z(n75092) );
  IV U85346 ( .A(n65045), .Z(n65047) );
  NOR U85347 ( .A(n65047), .B(n65046), .Z(n75078) );
  IV U85348 ( .A(n65048), .Z(n65049) );
  NOR U85349 ( .A(n65049), .B(n69818), .Z(n65050) );
  IV U85350 ( .A(n65050), .Z(n65051) );
  NOR U85351 ( .A(n65052), .B(n65051), .Z(n75072) );
  NOR U85352 ( .A(n75078), .B(n75072), .Z(n70142) );
  IV U85353 ( .A(n65053), .Z(n65054) );
  NOR U85354 ( .A(n65057), .B(n65054), .Z(n70154) );
  IV U85355 ( .A(n65055), .Z(n65056) );
  NOR U85356 ( .A(n65057), .B(n65056), .Z(n70151) );
  IV U85357 ( .A(n65062), .Z(n65059) );
  IV U85358 ( .A(n65058), .Z(n65061) );
  NOR U85359 ( .A(n65059), .B(n65061), .Z(n75048) );
  IV U85360 ( .A(n65060), .Z(n65064) );
  XOR U85361 ( .A(n65062), .B(n65061), .Z(n65063) );
  NOR U85362 ( .A(n65064), .B(n65063), .Z(n70157) );
  NOR U85363 ( .A(n75048), .B(n70157), .Z(n69795) );
  NOR U85364 ( .A(n65066), .B(n65065), .Z(n75045) );
  IV U85365 ( .A(n65067), .Z(n65068) );
  NOR U85366 ( .A(n65068), .B(n69792), .Z(n69789) );
  IV U85367 ( .A(n69789), .Z(n69779) );
  NOR U85368 ( .A(n65069), .B(n75022), .Z(n69785) );
  IV U85369 ( .A(n65070), .Z(n65071) );
  NOR U85370 ( .A(n65076), .B(n65071), .Z(n75008) );
  IV U85371 ( .A(n65072), .Z(n65074) );
  NOR U85372 ( .A(n65074), .B(n65073), .Z(n74997) );
  IV U85373 ( .A(n65075), .Z(n65077) );
  NOR U85374 ( .A(n65077), .B(n65076), .Z(n70183) );
  NOR U85375 ( .A(n74997), .B(n70183), .Z(n69769) );
  IV U85376 ( .A(n65078), .Z(n65079) );
  NOR U85377 ( .A(n69768), .B(n65079), .Z(n70185) );
  IV U85378 ( .A(n65080), .Z(n69755) );
  NOR U85379 ( .A(n69755), .B(n65081), .Z(n69747) );
  IV U85380 ( .A(n65082), .Z(n65084) );
  IV U85381 ( .A(n65083), .Z(n69732) );
  NOR U85382 ( .A(n65084), .B(n69732), .Z(n70192) );
  IV U85383 ( .A(n65085), .Z(n65086) );
  NOR U85384 ( .A(n65088), .B(n65086), .Z(n74965) );
  IV U85385 ( .A(n65087), .Z(n65089) );
  NOR U85386 ( .A(n65089), .B(n65088), .Z(n70204) );
  IV U85387 ( .A(n65090), .Z(n65092) );
  NOR U85388 ( .A(n65092), .B(n65091), .Z(n75532) );
  IV U85389 ( .A(n65093), .Z(n65094) );
  NOR U85390 ( .A(n65094), .B(n69716), .Z(n75527) );
  NOR U85391 ( .A(n75532), .B(n75527), .Z(n70207) );
  IV U85392 ( .A(n65095), .Z(n65102) );
  IV U85393 ( .A(n65096), .Z(n65097) );
  NOR U85394 ( .A(n65102), .B(n65097), .Z(n70212) );
  IV U85395 ( .A(n65098), .Z(n65099) );
  NOR U85396 ( .A(n65108), .B(n65099), .Z(n70218) );
  IV U85397 ( .A(n65100), .Z(n65101) );
  NOR U85398 ( .A(n65102), .B(n65101), .Z(n70216) );
  NOR U85399 ( .A(n70218), .B(n70216), .Z(n69714) );
  IV U85400 ( .A(n65103), .Z(n65104) );
  NOR U85401 ( .A(n65105), .B(n65104), .Z(n74955) );
  IV U85402 ( .A(n65106), .Z(n65107) );
  NOR U85403 ( .A(n65108), .B(n65107), .Z(n74958) );
  NOR U85404 ( .A(n74955), .B(n74958), .Z(n69713) );
  IV U85405 ( .A(n65109), .Z(n65110) );
  NOR U85406 ( .A(n65110), .B(n69704), .Z(n75560) );
  IV U85407 ( .A(n65111), .Z(n65112) );
  NOR U85408 ( .A(n69704), .B(n65112), .Z(n75555) );
  NOR U85409 ( .A(n75560), .B(n75555), .Z(n74946) );
  IV U85410 ( .A(n65113), .Z(n65114) );
  NOR U85411 ( .A(n65115), .B(n65114), .Z(n69698) );
  IV U85412 ( .A(n65116), .Z(n65119) );
  NOR U85413 ( .A(n65125), .B(n65121), .Z(n65117) );
  IV U85414 ( .A(n65117), .Z(n65118) );
  NOR U85415 ( .A(n65119), .B(n65118), .Z(n70224) );
  IV U85416 ( .A(n65120), .Z(n65122) );
  NOR U85417 ( .A(n65122), .B(n65121), .Z(n65123) );
  IV U85418 ( .A(n65123), .Z(n65124) );
  NOR U85419 ( .A(n65125), .B(n65124), .Z(n75563) );
  IV U85420 ( .A(n65126), .Z(n65128) );
  NOR U85421 ( .A(n65128), .B(n65127), .Z(n75571) );
  NOR U85422 ( .A(n75563), .B(n75571), .Z(n70233) );
  IV U85423 ( .A(n70233), .Z(n69689) );
  IV U85424 ( .A(n65129), .Z(n65130) );
  NOR U85425 ( .A(n65130), .B(n65132), .Z(n70230) );
  IV U85426 ( .A(n65131), .Z(n65133) );
  NOR U85427 ( .A(n65133), .B(n65132), .Z(n74935) );
  IV U85428 ( .A(n65134), .Z(n65135) );
  NOR U85429 ( .A(n65136), .B(n65135), .Z(n69686) );
  IV U85430 ( .A(n69686), .Z(n69680) );
  IV U85431 ( .A(n65137), .Z(n65138) );
  NOR U85432 ( .A(n65139), .B(n65138), .Z(n65140) );
  IV U85433 ( .A(n65140), .Z(n70244) );
  IV U85434 ( .A(n65141), .Z(n65143) );
  NOR U85435 ( .A(n65143), .B(n65142), .Z(n70248) );
  IV U85436 ( .A(n65144), .Z(n65145) );
  NOR U85437 ( .A(n65146), .B(n65145), .Z(n74930) );
  NOR U85438 ( .A(n70248), .B(n74930), .Z(n69668) );
  IV U85439 ( .A(n65147), .Z(n65150) );
  NOR U85440 ( .A(n65148), .B(n65155), .Z(n65149) );
  IV U85441 ( .A(n65149), .Z(n69665) );
  NOR U85442 ( .A(n65150), .B(n69665), .Z(n74914) );
  IV U85443 ( .A(n65151), .Z(n65153) );
  NOR U85444 ( .A(n65153), .B(n65152), .Z(n80305) );
  IV U85445 ( .A(n65154), .Z(n65156) );
  NOR U85446 ( .A(n65156), .B(n65155), .Z(n75584) );
  NOR U85447 ( .A(n80305), .B(n75584), .Z(n74910) );
  IV U85448 ( .A(n65157), .Z(n65161) );
  NOR U85449 ( .A(n65159), .B(n65158), .Z(n65160) );
  IV U85450 ( .A(n65160), .Z(n69657) );
  NOR U85451 ( .A(n65161), .B(n69657), .Z(n74907) );
  XOR U85452 ( .A(n65163), .B(n65162), .Z(n65164) );
  IV U85453 ( .A(n65164), .Z(n65171) );
  NOR U85454 ( .A(n65166), .B(n65165), .Z(n65167) );
  IV U85455 ( .A(n65167), .Z(n69651) );
  NOR U85456 ( .A(n65168), .B(n69651), .Z(n65169) );
  IV U85457 ( .A(n65169), .Z(n65170) );
  NOR U85458 ( .A(n65171), .B(n65170), .Z(n65172) );
  IV U85459 ( .A(n65172), .Z(n70260) );
  IV U85460 ( .A(n65173), .Z(n65174) );
  NOR U85461 ( .A(n65175), .B(n65174), .Z(n70276) );
  IV U85462 ( .A(n65176), .Z(n65177) );
  NOR U85463 ( .A(n65177), .B(n69630), .Z(n70274) );
  NOR U85464 ( .A(n70276), .B(n70274), .Z(n69626) );
  IV U85465 ( .A(n65178), .Z(n69624) );
  IV U85466 ( .A(n65179), .Z(n65180) );
  NOR U85467 ( .A(n69624), .B(n65180), .Z(n70282) );
  IV U85468 ( .A(n65181), .Z(n65182) );
  NOR U85469 ( .A(n65182), .B(n69624), .Z(n70279) );
  IV U85470 ( .A(n65183), .Z(n65185) );
  NOR U85471 ( .A(n65185), .B(n65184), .Z(n75630) );
  NOR U85472 ( .A(n65187), .B(n65186), .Z(n75620) );
  NOR U85473 ( .A(n75630), .B(n75620), .Z(n74899) );
  IV U85474 ( .A(n65188), .Z(n65190) );
  NOR U85475 ( .A(n65190), .B(n65189), .Z(n70292) );
  IV U85476 ( .A(n65191), .Z(n65192) );
  NOR U85477 ( .A(n65192), .B(n65197), .Z(n65193) );
  IV U85478 ( .A(n65193), .Z(n65194) );
  NOR U85479 ( .A(n69598), .B(n65194), .Z(n70304) );
  IV U85480 ( .A(n65195), .Z(n65196) );
  NOR U85481 ( .A(n65197), .B(n65196), .Z(n70310) );
  NOR U85482 ( .A(n74882), .B(n70310), .Z(n69593) );
  IV U85483 ( .A(n69591), .Z(n69586) );
  IV U85484 ( .A(n65198), .Z(n65200) );
  NOR U85485 ( .A(n65200), .B(n65199), .Z(n70313) );
  IV U85486 ( .A(n65201), .Z(n65203) );
  NOR U85487 ( .A(n65203), .B(n65202), .Z(n70317) );
  IV U85488 ( .A(n65204), .Z(n65206) );
  NOR U85489 ( .A(n65206), .B(n65205), .Z(n70315) );
  NOR U85490 ( .A(n70317), .B(n70315), .Z(n65207) );
  IV U85491 ( .A(n65207), .Z(n69584) );
  IV U85492 ( .A(n65208), .Z(n65210) );
  NOR U85493 ( .A(n65210), .B(n65209), .Z(n74869) );
  IV U85494 ( .A(n65211), .Z(n65212) );
  NOR U85495 ( .A(n65213), .B(n65212), .Z(n74874) );
  NOR U85496 ( .A(n74869), .B(n74874), .Z(n69583) );
  IV U85497 ( .A(n65214), .Z(n65216) );
  NOR U85498 ( .A(n65216), .B(n65215), .Z(n75669) );
  IV U85499 ( .A(n65217), .Z(n65219) );
  NOR U85500 ( .A(n65219), .B(n65218), .Z(n80246) );
  NOR U85501 ( .A(n75669), .B(n80246), .Z(n74868) );
  IV U85502 ( .A(n65220), .Z(n65221) );
  NOR U85503 ( .A(n65227), .B(n65221), .Z(n74851) );
  IV U85504 ( .A(n74851), .Z(n74848) );
  IV U85505 ( .A(n65222), .Z(n65224) );
  IV U85506 ( .A(n65223), .Z(n69571) );
  NOR U85507 ( .A(n65224), .B(n69571), .Z(n70331) );
  IV U85508 ( .A(n65225), .Z(n65226) );
  NOR U85509 ( .A(n65227), .B(n65226), .Z(n70329) );
  NOR U85510 ( .A(n70331), .B(n70329), .Z(n69573) );
  IV U85511 ( .A(n65228), .Z(n65229) );
  NOR U85512 ( .A(n69554), .B(n65229), .Z(n74821) );
  IV U85513 ( .A(n65230), .Z(n65231) );
  NOR U85514 ( .A(n65232), .B(n65231), .Z(n75690) );
  IV U85515 ( .A(n65233), .Z(n65234) );
  NOR U85516 ( .A(n69550), .B(n65234), .Z(n75684) );
  NOR U85517 ( .A(n75690), .B(n75684), .Z(n74813) );
  IV U85518 ( .A(n74813), .Z(n69548) );
  IV U85519 ( .A(n65235), .Z(n65236) );
  NOR U85520 ( .A(n65239), .B(n65236), .Z(n70342) );
  IV U85521 ( .A(n65237), .Z(n65238) );
  NOR U85522 ( .A(n65239), .B(n65238), .Z(n74801) );
  IV U85523 ( .A(n65240), .Z(n65241) );
  NOR U85524 ( .A(n65241), .B(n65244), .Z(n70345) );
  IV U85525 ( .A(n65242), .Z(n65243) );
  NOR U85526 ( .A(n65243), .B(n69546), .Z(n74794) );
  NOR U85527 ( .A(n65245), .B(n65244), .Z(n74791) );
  IV U85528 ( .A(n65246), .Z(n65249) );
  IV U85529 ( .A(n65247), .Z(n65248) );
  NOR U85530 ( .A(n65249), .B(n65248), .Z(n65250) );
  IV U85531 ( .A(n65250), .Z(n70353) );
  NOR U85532 ( .A(n65251), .B(n70358), .Z(n69539) );
  IV U85533 ( .A(n65252), .Z(n65253) );
  NOR U85534 ( .A(n65260), .B(n65253), .Z(n74783) );
  IV U85535 ( .A(n65254), .Z(n65255) );
  NOR U85536 ( .A(n65256), .B(n65255), .Z(n70364) );
  NOR U85537 ( .A(n74783), .B(n70364), .Z(n65257) );
  IV U85538 ( .A(n65257), .Z(n69538) );
  IV U85539 ( .A(n65258), .Z(n65259) );
  NOR U85540 ( .A(n65260), .B(n65259), .Z(n74780) );
  IV U85541 ( .A(n65261), .Z(n65262) );
  NOR U85542 ( .A(n65262), .B(n69528), .Z(n70370) );
  IV U85543 ( .A(n65263), .Z(n65265) );
  NOR U85544 ( .A(n65265), .B(n65264), .Z(n69524) );
  IV U85545 ( .A(n69524), .Z(n69512) );
  IV U85546 ( .A(n65266), .Z(n65267) );
  NOR U85547 ( .A(n65270), .B(n65267), .Z(n70375) );
  IV U85548 ( .A(n65268), .Z(n65269) );
  NOR U85549 ( .A(n65270), .B(n65269), .Z(n70381) );
  IV U85550 ( .A(n65271), .Z(n65272) );
  NOR U85551 ( .A(n65273), .B(n65272), .Z(n75734) );
  NOR U85552 ( .A(n75739), .B(n75734), .Z(n74764) );
  IV U85553 ( .A(n65274), .Z(n65275) );
  NOR U85554 ( .A(n65275), .B(n69503), .Z(n74761) );
  IV U85555 ( .A(n65276), .Z(n65277) );
  NOR U85556 ( .A(n65277), .B(n65283), .Z(n65278) );
  IV U85557 ( .A(n65278), .Z(n74743) );
  IV U85558 ( .A(n65279), .Z(n65281) );
  NOR U85559 ( .A(n65281), .B(n65280), .Z(n74735) );
  IV U85560 ( .A(n65282), .Z(n65284) );
  NOR U85561 ( .A(n65284), .B(n65283), .Z(n74738) );
  NOR U85562 ( .A(n74735), .B(n74738), .Z(n69494) );
  IV U85563 ( .A(n65285), .Z(n65292) );
  IV U85564 ( .A(n65286), .Z(n65287) );
  NOR U85565 ( .A(n65292), .B(n65287), .Z(n74732) );
  IV U85566 ( .A(n65288), .Z(n65289) );
  NOR U85567 ( .A(n65292), .B(n65289), .Z(n74728) );
  IV U85568 ( .A(n65290), .Z(n65294) );
  NOR U85569 ( .A(n65292), .B(n65291), .Z(n65293) );
  IV U85570 ( .A(n65293), .Z(n65296) );
  NOR U85571 ( .A(n65294), .B(n65296), .Z(n74725) );
  IV U85572 ( .A(n65295), .Z(n65297) );
  NOR U85573 ( .A(n65297), .B(n65296), .Z(n70388) );
  IV U85574 ( .A(n65298), .Z(n65299) );
  NOR U85575 ( .A(n65299), .B(n65301), .Z(n74713) );
  IV U85576 ( .A(n65300), .Z(n65302) );
  NOR U85577 ( .A(n65302), .B(n65301), .Z(n70391) );
  IV U85578 ( .A(n65303), .Z(n69485) );
  IV U85579 ( .A(n65304), .Z(n65305) );
  NOR U85580 ( .A(n69485), .B(n65305), .Z(n74707) );
  IV U85581 ( .A(n65306), .Z(n65307) );
  NOR U85582 ( .A(n65307), .B(n69490), .Z(n65308) );
  IV U85583 ( .A(n65308), .Z(n70400) );
  IV U85584 ( .A(n65309), .Z(n65311) );
  NOR U85585 ( .A(n65311), .B(n65310), .Z(n74699) );
  IV U85586 ( .A(n65312), .Z(n65314) );
  NOR U85587 ( .A(n65314), .B(n65313), .Z(n70396) );
  NOR U85588 ( .A(n74699), .B(n70396), .Z(n69481) );
  IV U85589 ( .A(n65315), .Z(n65317) );
  NOR U85590 ( .A(n65317), .B(n65316), .Z(n70402) );
  IV U85591 ( .A(n65318), .Z(n65320) );
  NOR U85592 ( .A(n65320), .B(n65319), .Z(n74696) );
  NOR U85593 ( .A(n70402), .B(n74696), .Z(n69480) );
  IV U85594 ( .A(n65321), .Z(n65323) );
  NOR U85595 ( .A(n65323), .B(n65322), .Z(n70406) );
  IV U85596 ( .A(n65324), .Z(n65326) );
  NOR U85597 ( .A(n65326), .B(n65325), .Z(n74693) );
  NOR U85598 ( .A(n70406), .B(n74693), .Z(n69479) );
  IV U85599 ( .A(n65327), .Z(n65329) );
  NOR U85600 ( .A(n65329), .B(n65328), .Z(n70404) );
  NOR U85601 ( .A(n65331), .B(n65330), .Z(n65332) );
  IV U85602 ( .A(n65332), .Z(n65333) );
  NOR U85603 ( .A(n65334), .B(n65333), .Z(n70409) );
  IV U85604 ( .A(n65335), .Z(n65337) );
  NOR U85605 ( .A(n65337), .B(n65336), .Z(n70423) );
  NOR U85606 ( .A(n70419), .B(n70423), .Z(n69472) );
  IV U85607 ( .A(n65338), .Z(n65339) );
  NOR U85608 ( .A(n65339), .B(n69466), .Z(n65340) );
  IV U85609 ( .A(n65340), .Z(n74683) );
  IV U85610 ( .A(n65341), .Z(n65342) );
  NOR U85611 ( .A(n65343), .B(n65342), .Z(n74680) );
  IV U85612 ( .A(n65344), .Z(n65346) );
  NOR U85613 ( .A(n65346), .B(n65345), .Z(n74685) );
  NOR U85614 ( .A(n74680), .B(n74685), .Z(n69464) );
  IV U85615 ( .A(n65347), .Z(n65348) );
  NOR U85616 ( .A(n65348), .B(n69462), .Z(n70434) );
  IV U85617 ( .A(n65349), .Z(n65351) );
  NOR U85618 ( .A(n65351), .B(n65350), .Z(n69456) );
  IV U85619 ( .A(n65352), .Z(n65353) );
  NOR U85620 ( .A(n65354), .B(n65353), .Z(n65355) );
  IV U85621 ( .A(n65355), .Z(n65356) );
  NOR U85622 ( .A(n65357), .B(n65356), .Z(n65358) );
  IV U85623 ( .A(n65358), .Z(n70438) );
  IV U85624 ( .A(n65359), .Z(n65360) );
  NOR U85625 ( .A(n69438), .B(n65360), .Z(n74653) );
  IV U85626 ( .A(n65361), .Z(n65362) );
  NOR U85627 ( .A(n69438), .B(n65362), .Z(n74638) );
  IV U85628 ( .A(n65363), .Z(n65367) );
  IV U85629 ( .A(n69438), .Z(n65364) );
  NOR U85630 ( .A(n65371), .B(n65364), .Z(n65365) );
  IV U85631 ( .A(n65365), .Z(n65366) );
  NOR U85632 ( .A(n65367), .B(n65366), .Z(n74640) );
  NOR U85633 ( .A(n74638), .B(n74640), .Z(n65368) );
  IV U85634 ( .A(n65368), .Z(n69433) );
  IV U85635 ( .A(n65369), .Z(n65374) );
  IV U85636 ( .A(n65370), .Z(n69431) );
  NOR U85637 ( .A(n65371), .B(n69431), .Z(n65372) );
  IV U85638 ( .A(n65372), .Z(n65373) );
  NOR U85639 ( .A(n65374), .B(n65373), .Z(n70439) );
  IV U85640 ( .A(n65375), .Z(n65376) );
  NOR U85641 ( .A(n69429), .B(n65376), .Z(n69425) );
  IV U85642 ( .A(n69425), .Z(n69419) );
  IV U85643 ( .A(n65377), .Z(n65379) );
  NOR U85644 ( .A(n65379), .B(n65378), .Z(n70445) );
  NOR U85645 ( .A(n65381), .B(n65380), .Z(n65382) );
  IV U85646 ( .A(n65382), .Z(n65388) );
  IV U85647 ( .A(n65383), .Z(n65384) );
  NOR U85648 ( .A(n65385), .B(n65384), .Z(n65386) );
  IV U85649 ( .A(n65386), .Z(n65387) );
  NOR U85650 ( .A(n65388), .B(n65387), .Z(n70453) );
  IV U85651 ( .A(n65389), .Z(n65390) );
  NOR U85652 ( .A(n65391), .B(n65390), .Z(n70451) );
  IV U85653 ( .A(n65392), .Z(n65394) );
  NOR U85654 ( .A(n65394), .B(n65393), .Z(n74629) );
  NOR U85655 ( .A(n70451), .B(n74629), .Z(n69417) );
  XOR U85656 ( .A(n65396), .B(n65395), .Z(n65397) );
  NOR U85657 ( .A(n65397), .B(n65402), .Z(n65398) );
  IV U85658 ( .A(n65398), .Z(n65399) );
  NOR U85659 ( .A(n65400), .B(n65399), .Z(n74632) );
  IV U85660 ( .A(n65401), .Z(n65403) );
  NOR U85661 ( .A(n65403), .B(n65402), .Z(n74627) );
  IV U85662 ( .A(n65404), .Z(n65405) );
  NOR U85663 ( .A(n65406), .B(n65405), .Z(n74613) );
  NOR U85664 ( .A(n74627), .B(n74613), .Z(n65407) );
  IV U85665 ( .A(n65407), .Z(n65408) );
  NOR U85666 ( .A(n74632), .B(n65408), .Z(n69416) );
  IV U85667 ( .A(n65409), .Z(n65414) );
  IV U85668 ( .A(n65410), .Z(n65411) );
  NOR U85669 ( .A(n65414), .B(n65411), .Z(n74610) );
  IV U85670 ( .A(n65412), .Z(n65413) );
  NOR U85671 ( .A(n65414), .B(n65413), .Z(n70456) );
  IV U85672 ( .A(n65415), .Z(n65416) );
  NOR U85673 ( .A(n65417), .B(n65416), .Z(n70462) );
  IV U85674 ( .A(n65418), .Z(n65420) );
  NOR U85675 ( .A(n65420), .B(n65419), .Z(n70477) );
  NOR U85676 ( .A(n65421), .B(n65428), .Z(n65422) );
  IV U85677 ( .A(n65422), .Z(n75828) );
  NOR U85678 ( .A(n65423), .B(n75828), .Z(n70484) );
  IV U85679 ( .A(n65424), .Z(n65426) );
  NOR U85680 ( .A(n65426), .B(n65425), .Z(n70487) );
  IV U85681 ( .A(n65427), .Z(n65429) );
  NOR U85682 ( .A(n65429), .B(n65428), .Z(n70482) );
  NOR U85683 ( .A(n70487), .B(n70482), .Z(n69393) );
  IV U85684 ( .A(n65430), .Z(n65431) );
  NOR U85685 ( .A(n65431), .B(n69379), .Z(n70490) );
  IV U85686 ( .A(n65432), .Z(n65433) );
  NOR U85687 ( .A(n65433), .B(n65435), .Z(n70493) );
  IV U85688 ( .A(n65434), .Z(n65436) );
  NOR U85689 ( .A(n65436), .B(n65435), .Z(n74585) );
  NOR U85690 ( .A(n70493), .B(n74585), .Z(n65437) );
  IV U85691 ( .A(n65437), .Z(n65441) );
  IV U85692 ( .A(n65438), .Z(n65439) );
  NOR U85693 ( .A(n65440), .B(n65439), .Z(n74581) );
  NOR U85694 ( .A(n65441), .B(n74581), .Z(n65442) );
  IV U85695 ( .A(n65442), .Z(n69377) );
  IV U85696 ( .A(n65443), .Z(n65445) );
  IV U85697 ( .A(n65444), .Z(n65450) );
  NOR U85698 ( .A(n65445), .B(n65450), .Z(n74578) );
  NOR U85699 ( .A(n65447), .B(n65446), .Z(n75850) );
  IV U85700 ( .A(n65448), .Z(n65449) );
  NOR U85701 ( .A(n65450), .B(n65449), .Z(n75845) );
  NOR U85702 ( .A(n75850), .B(n75845), .Z(n70496) );
  IV U85703 ( .A(n65451), .Z(n65452) );
  NOR U85704 ( .A(n65453), .B(n65452), .Z(n74569) );
  NOR U85705 ( .A(n74571), .B(n74569), .Z(n69376) );
  IV U85706 ( .A(n65454), .Z(n65455) );
  NOR U85707 ( .A(n65455), .B(n65457), .Z(n74566) );
  IV U85708 ( .A(n65456), .Z(n65458) );
  NOR U85709 ( .A(n65458), .B(n65457), .Z(n74562) );
  IV U85710 ( .A(n65459), .Z(n65464) );
  IV U85711 ( .A(n65460), .Z(n65461) );
  NOR U85712 ( .A(n65464), .B(n65461), .Z(n74559) );
  IV U85713 ( .A(n65462), .Z(n65463) );
  NOR U85714 ( .A(n65464), .B(n65463), .Z(n74554) );
  IV U85715 ( .A(n65465), .Z(n65466) );
  NOR U85716 ( .A(n65466), .B(n69373), .Z(n74551) );
  IV U85717 ( .A(n65467), .Z(n65468) );
  NOR U85718 ( .A(n65468), .B(n65474), .Z(n65469) );
  IV U85719 ( .A(n65469), .Z(n74539) );
  IV U85720 ( .A(n65470), .Z(n75886) );
  NOR U85721 ( .A(n75886), .B(n65471), .Z(n74531) );
  IV U85722 ( .A(n65472), .Z(n65473) );
  NOR U85723 ( .A(n65474), .B(n65473), .Z(n74535) );
  NOR U85724 ( .A(n74531), .B(n74535), .Z(n69364) );
  IV U85725 ( .A(n65475), .Z(n65480) );
  IV U85726 ( .A(n65476), .Z(n65477) );
  NOR U85727 ( .A(n65480), .B(n65477), .Z(n70512) );
  IV U85728 ( .A(n65478), .Z(n65479) );
  NOR U85729 ( .A(n65480), .B(n65479), .Z(n70509) );
  IV U85730 ( .A(n65481), .Z(n65482) );
  NOR U85731 ( .A(n65482), .B(n75905), .Z(n70523) );
  NOR U85732 ( .A(n75894), .B(n75905), .Z(n65483) );
  IV U85733 ( .A(n65483), .Z(n65484) );
  NOR U85734 ( .A(n65485), .B(n65484), .Z(n65486) );
  IV U85735 ( .A(n65486), .Z(n70529) );
  NOR U85736 ( .A(n65487), .B(n70529), .Z(n69346) );
  IV U85737 ( .A(n65488), .Z(n65489) );
  NOR U85738 ( .A(n65489), .B(n65491), .Z(n74521) );
  IV U85739 ( .A(n65490), .Z(n65494) );
  NOR U85740 ( .A(n65492), .B(n65491), .Z(n65493) );
  IV U85741 ( .A(n65493), .Z(n65500) );
  NOR U85742 ( .A(n65494), .B(n65500), .Z(n65495) );
  IV U85743 ( .A(n65495), .Z(n74520) );
  IV U85744 ( .A(n65496), .Z(n65504) );
  IV U85745 ( .A(n65497), .Z(n65498) );
  NOR U85746 ( .A(n65504), .B(n65498), .Z(n70537) );
  IV U85747 ( .A(n65499), .Z(n65501) );
  NOR U85748 ( .A(n65501), .B(n65500), .Z(n70532) );
  NOR U85749 ( .A(n70537), .B(n70532), .Z(n69345) );
  IV U85750 ( .A(n65502), .Z(n65503) );
  NOR U85751 ( .A(n65504), .B(n65503), .Z(n70534) );
  IV U85752 ( .A(n65505), .Z(n65506) );
  NOR U85753 ( .A(n65507), .B(n65506), .Z(n70543) );
  IV U85754 ( .A(n65508), .Z(n65511) );
  NOR U85755 ( .A(n65509), .B(n65519), .Z(n65510) );
  IV U85756 ( .A(n65510), .Z(n65513) );
  NOR U85757 ( .A(n65511), .B(n65513), .Z(n70540) );
  IV U85758 ( .A(n65512), .Z(n65514) );
  NOR U85759 ( .A(n65514), .B(n65513), .Z(n70548) );
  IV U85760 ( .A(n65515), .Z(n65516) );
  NOR U85761 ( .A(n65517), .B(n65516), .Z(n75916) );
  IV U85762 ( .A(n65518), .Z(n65520) );
  NOR U85763 ( .A(n65520), .B(n65519), .Z(n75909) );
  NOR U85764 ( .A(n75916), .B(n75909), .Z(n70547) );
  IV U85765 ( .A(n65521), .Z(n65523) );
  NOR U85766 ( .A(n65523), .B(n65522), .Z(n74503) );
  NOR U85767 ( .A(n65524), .B(n70553), .Z(n65525) );
  NOR U85768 ( .A(n74503), .B(n65525), .Z(n69344) );
  IV U85769 ( .A(n65526), .Z(n65527) );
  NOR U85770 ( .A(n65533), .B(n65527), .Z(n65528) );
  IV U85771 ( .A(n65528), .Z(n74508) );
  IV U85772 ( .A(n65529), .Z(n65530) );
  NOR U85773 ( .A(n65531), .B(n65530), .Z(n79891) );
  IV U85774 ( .A(n65532), .Z(n65534) );
  NOR U85775 ( .A(n65534), .B(n65533), .Z(n79898) );
  NOR U85776 ( .A(n79891), .B(n79898), .Z(n70557) );
  NOR U85777 ( .A(n65535), .B(n70560), .Z(n65539) );
  IV U85778 ( .A(n65536), .Z(n65538) );
  NOR U85779 ( .A(n65538), .B(n65537), .Z(n74498) );
  NOR U85780 ( .A(n65539), .B(n74498), .Z(n69343) );
  IV U85781 ( .A(n65540), .Z(n65541) );
  NOR U85782 ( .A(n65541), .B(n65544), .Z(n70566) );
  IV U85783 ( .A(n65542), .Z(n65543) );
  NOR U85784 ( .A(n65544), .B(n65543), .Z(n74490) );
  IV U85785 ( .A(n65545), .Z(n65546) );
  NOR U85786 ( .A(n65547), .B(n65546), .Z(n70572) );
  NOR U85787 ( .A(n74490), .B(n70572), .Z(n69334) );
  IV U85788 ( .A(n65548), .Z(n65550) );
  NOR U85789 ( .A(n65550), .B(n65549), .Z(n74488) );
  IV U85790 ( .A(n65551), .Z(n65553) );
  IV U85791 ( .A(n65552), .Z(n65556) );
  NOR U85792 ( .A(n65553), .B(n65556), .Z(n70578) );
  IV U85793 ( .A(n65554), .Z(n65555) );
  NOR U85794 ( .A(n65556), .B(n65555), .Z(n70575) );
  IV U85795 ( .A(n65557), .Z(n65558) );
  NOR U85796 ( .A(n65561), .B(n65558), .Z(n70584) );
  IV U85797 ( .A(n65559), .Z(n65560) );
  NOR U85798 ( .A(n65561), .B(n65560), .Z(n70595) );
  IV U85799 ( .A(n65562), .Z(n65563) );
  NOR U85800 ( .A(n65563), .B(n69311), .Z(n70601) );
  IV U85801 ( .A(n65564), .Z(n65566) );
  NOR U85802 ( .A(n65566), .B(n65565), .Z(n70606) );
  IV U85803 ( .A(n65567), .Z(n65568) );
  NOR U85804 ( .A(n69300), .B(n65568), .Z(n74473) );
  NOR U85805 ( .A(n70606), .B(n74473), .Z(n69306) );
  IV U85806 ( .A(n65569), .Z(n65570) );
  NOR U85807 ( .A(n65571), .B(n65570), .Z(n79845) );
  IV U85808 ( .A(n65572), .Z(n65573) );
  NOR U85809 ( .A(n65574), .B(n65573), .Z(n79852) );
  NOR U85810 ( .A(n79845), .B(n79852), .Z(n74478) );
  IV U85811 ( .A(n65575), .Z(n65576) );
  NOR U85812 ( .A(n65577), .B(n65576), .Z(n70612) );
  IV U85813 ( .A(n65578), .Z(n65580) );
  NOR U85814 ( .A(n65580), .B(n65579), .Z(n70614) );
  NOR U85815 ( .A(n70612), .B(n70614), .Z(n69298) );
  IV U85816 ( .A(n65581), .Z(n65582) );
  NOR U85817 ( .A(n65582), .B(n70617), .Z(n69297) );
  IV U85818 ( .A(n65583), .Z(n65585) );
  NOR U85819 ( .A(n65585), .B(n65584), .Z(n70632) );
  IV U85820 ( .A(n65586), .Z(n65587) );
  NOR U85821 ( .A(n65587), .B(n70617), .Z(n70627) );
  NOR U85822 ( .A(n70632), .B(n70627), .Z(n65588) );
  IV U85823 ( .A(n65588), .Z(n69296) );
  IV U85824 ( .A(n65589), .Z(n65590) );
  NOR U85825 ( .A(n65591), .B(n65590), .Z(n70630) );
  IV U85826 ( .A(n65592), .Z(n65595) );
  IV U85827 ( .A(n65593), .Z(n65594) );
  NOR U85828 ( .A(n65595), .B(n65594), .Z(n70638) );
  IV U85829 ( .A(n65596), .Z(n65598) );
  XOR U85830 ( .A(n69292), .B(n69293), .Z(n65597) );
  NOR U85831 ( .A(n65598), .B(n65597), .Z(n70635) );
  IV U85832 ( .A(n65599), .Z(n65600) );
  NOR U85833 ( .A(n65600), .B(n69280), .Z(n65601) );
  IV U85834 ( .A(n65601), .Z(n69285) );
  NOR U85835 ( .A(n65610), .B(n65602), .Z(n65603) );
  IV U85836 ( .A(n65603), .Z(n65608) );
  NOR U85837 ( .A(n65605), .B(n65604), .Z(n65606) );
  IV U85838 ( .A(n65606), .Z(n65607) );
  NOR U85839 ( .A(n65608), .B(n65607), .Z(n74451) );
  IV U85840 ( .A(n65609), .Z(n65611) );
  NOR U85841 ( .A(n65611), .B(n65610), .Z(n74448) );
  IV U85842 ( .A(n65612), .Z(n65613) );
  NOR U85843 ( .A(n65613), .B(n65618), .Z(n70645) );
  IV U85844 ( .A(n65614), .Z(n65615) );
  NOR U85845 ( .A(n65616), .B(n65615), .Z(n85585) );
  IV U85846 ( .A(n65617), .Z(n65619) );
  NOR U85847 ( .A(n65619), .B(n65618), .Z(n85593) );
  NOR U85848 ( .A(n85585), .B(n85593), .Z(n70644) );
  IV U85849 ( .A(n70644), .Z(n69278) );
  NOR U85850 ( .A(n65633), .B(n65620), .Z(n65621) );
  IV U85851 ( .A(n65621), .Z(n65628) );
  XOR U85852 ( .A(n65623), .B(n65622), .Z(n65624) );
  NOR U85853 ( .A(n65625), .B(n65624), .Z(n65626) );
  IV U85854 ( .A(n65626), .Z(n65627) );
  NOR U85855 ( .A(n65628), .B(n65627), .Z(n74441) );
  IV U85856 ( .A(n65629), .Z(n65630) );
  NOR U85857 ( .A(n65633), .B(n65630), .Z(n74437) );
  IV U85858 ( .A(n65631), .Z(n65632) );
  NOR U85859 ( .A(n65633), .B(n65632), .Z(n74434) );
  IV U85860 ( .A(n65634), .Z(n65636) );
  IV U85861 ( .A(n65635), .Z(n65639) );
  NOR U85862 ( .A(n65636), .B(n65639), .Z(n74427) );
  NOR U85863 ( .A(n70649), .B(n65637), .Z(n65641) );
  IV U85864 ( .A(n65638), .Z(n65640) );
  NOR U85865 ( .A(n65640), .B(n65639), .Z(n74430) );
  NOR U85866 ( .A(n65641), .B(n74430), .Z(n69272) );
  IV U85867 ( .A(n65642), .Z(n65643) );
  NOR U85868 ( .A(n65643), .B(n69254), .Z(n85543) );
  NOR U85869 ( .A(n69251), .B(n65644), .Z(n70661) );
  IV U85870 ( .A(n65645), .Z(n79800) );
  IV U85871 ( .A(n65646), .Z(n65647) );
  NOR U85872 ( .A(n79800), .B(n65647), .Z(n74412) );
  IV U85873 ( .A(n65648), .Z(n65651) );
  NOR U85874 ( .A(n65649), .B(n65659), .Z(n65650) );
  IV U85875 ( .A(n65650), .Z(n65653) );
  NOR U85876 ( .A(n65651), .B(n65653), .Z(n74408) );
  IV U85877 ( .A(n65652), .Z(n65654) );
  NOR U85878 ( .A(n65654), .B(n65653), .Z(n74405) );
  IV U85879 ( .A(n65655), .Z(n65656) );
  NOR U85880 ( .A(n65657), .B(n65656), .Z(n74399) );
  IV U85881 ( .A(n65658), .Z(n65660) );
  NOR U85882 ( .A(n65660), .B(n65659), .Z(n74402) );
  NOR U85883 ( .A(n74399), .B(n74402), .Z(n69246) );
  IV U85884 ( .A(n65661), .Z(n65663) );
  NOR U85885 ( .A(n65663), .B(n65662), .Z(n74388) );
  IV U85886 ( .A(n65664), .Z(n65666) );
  NOR U85887 ( .A(n65666), .B(n65665), .Z(n76047) );
  IV U85888 ( .A(n65667), .Z(n65669) );
  IV U85889 ( .A(n65668), .Z(n69238) );
  NOR U85890 ( .A(n65669), .B(n69238), .Z(n79753) );
  NOR U85891 ( .A(n76047), .B(n79753), .Z(n70668) );
  IV U85892 ( .A(n65670), .Z(n65671) );
  NOR U85893 ( .A(n65671), .B(n65677), .Z(n65672) );
  IV U85894 ( .A(n65672), .Z(n74368) );
  IV U85895 ( .A(n65673), .Z(n65681) );
  IV U85896 ( .A(n65674), .Z(n65675) );
  NOR U85897 ( .A(n65681), .B(n65675), .Z(n70675) );
  IV U85898 ( .A(n65676), .Z(n65678) );
  NOR U85899 ( .A(n65678), .B(n65677), .Z(n74370) );
  NOR U85900 ( .A(n70675), .B(n74370), .Z(n69229) );
  IV U85901 ( .A(n65679), .Z(n65680) );
  NOR U85902 ( .A(n65681), .B(n65680), .Z(n70672) );
  IV U85903 ( .A(n65682), .Z(n65683) );
  NOR U85904 ( .A(n65684), .B(n65683), .Z(n70685) );
  IV U85905 ( .A(n65685), .Z(n65686) );
  NOR U85906 ( .A(n65687), .B(n65686), .Z(n70677) );
  NOR U85907 ( .A(n70685), .B(n70677), .Z(n69220) );
  IV U85908 ( .A(n65688), .Z(n65690) );
  IV U85909 ( .A(n65689), .Z(n69216) );
  NOR U85910 ( .A(n65690), .B(n69216), .Z(n70682) );
  IV U85911 ( .A(n65691), .Z(n65693) );
  NOR U85912 ( .A(n65693), .B(n65692), .Z(n65694) );
  IV U85913 ( .A(n65694), .Z(n69206) );
  IV U85914 ( .A(n65695), .Z(n65697) );
  IV U85915 ( .A(n65696), .Z(n65699) );
  NOR U85916 ( .A(n65697), .B(n65699), .Z(n74331) );
  IV U85917 ( .A(n65698), .Z(n65700) );
  NOR U85918 ( .A(n65700), .B(n65699), .Z(n74328) );
  IV U85919 ( .A(n65701), .Z(n65702) );
  NOR U85920 ( .A(n65702), .B(n65706), .Z(n65703) );
  IV U85921 ( .A(n65703), .Z(n74325) );
  IV U85922 ( .A(n65704), .Z(n79721) );
  IV U85923 ( .A(n79724), .Z(n65710) );
  NOR U85924 ( .A(n79721), .B(n65710), .Z(n65708) );
  IV U85925 ( .A(n65705), .Z(n65707) );
  NOR U85926 ( .A(n65707), .B(n65706), .Z(n76101) );
  NOR U85927 ( .A(n65708), .B(n76101), .Z(n74322) );
  IV U85928 ( .A(n65709), .Z(n79725) );
  NOR U85929 ( .A(n79725), .B(n65710), .Z(n74304) );
  IV U85930 ( .A(n65711), .Z(n65712) );
  NOR U85931 ( .A(n65712), .B(n65718), .Z(n74308) );
  IV U85932 ( .A(n65713), .Z(n65714) );
  NOR U85933 ( .A(n65715), .B(n65714), .Z(n74300) );
  IV U85934 ( .A(n65716), .Z(n65717) );
  NOR U85935 ( .A(n65718), .B(n65717), .Z(n74311) );
  NOR U85936 ( .A(n74300), .B(n74311), .Z(n69199) );
  IV U85937 ( .A(n65719), .Z(n65721) );
  NOR U85938 ( .A(n65721), .B(n65720), .Z(n74298) );
  IV U85939 ( .A(n65722), .Z(n65724) );
  NOR U85940 ( .A(n65724), .B(n65723), .Z(n65725) );
  IV U85941 ( .A(n65725), .Z(n69187) );
  IV U85942 ( .A(n65726), .Z(n65727) );
  NOR U85943 ( .A(n65727), .B(n69181), .Z(n74276) );
  NOR U85944 ( .A(n65728), .B(n65737), .Z(n65729) );
  IV U85945 ( .A(n65729), .Z(n65730) );
  NOR U85946 ( .A(n65731), .B(n65730), .Z(n65732) );
  IV U85947 ( .A(n65732), .Z(n74271) );
  IV U85948 ( .A(n65733), .Z(n65735) );
  NOR U85949 ( .A(n65735), .B(n65734), .Z(n74267) );
  IV U85950 ( .A(n65736), .Z(n65738) );
  NOR U85951 ( .A(n65738), .B(n65737), .Z(n74273) );
  NOR U85952 ( .A(n74267), .B(n74273), .Z(n69176) );
  IV U85953 ( .A(n65739), .Z(n69171) );
  IV U85954 ( .A(n65740), .Z(n65741) );
  NOR U85955 ( .A(n69171), .B(n65741), .Z(n74264) );
  IV U85956 ( .A(n65742), .Z(n65743) );
  NOR U85957 ( .A(n65743), .B(n69174), .Z(n74258) );
  IV U85958 ( .A(n65744), .Z(n65746) );
  NOR U85959 ( .A(n65746), .B(n65745), .Z(n76151) );
  IV U85960 ( .A(n65747), .Z(n65748) );
  NOR U85961 ( .A(n65748), .B(n69167), .Z(n76147) );
  NOR U85962 ( .A(n76151), .B(n76147), .Z(n74252) );
  IV U85963 ( .A(n74252), .Z(n69165) );
  IV U85964 ( .A(n65749), .Z(n65751) );
  NOR U85965 ( .A(n65751), .B(n65750), .Z(n70706) );
  IV U85966 ( .A(n65752), .Z(n65753) );
  NOR U85967 ( .A(n65754), .B(n65753), .Z(n85465) );
  IV U85968 ( .A(n65755), .Z(n65757) );
  NOR U85969 ( .A(n65757), .B(n65756), .Z(n85479) );
  NOR U85970 ( .A(n85465), .B(n85479), .Z(n70709) );
  IV U85971 ( .A(n65758), .Z(n65759) );
  NOR U85972 ( .A(n65759), .B(n69155), .Z(n70714) );
  IV U85973 ( .A(n65760), .Z(n65761) );
  NOR U85974 ( .A(n65762), .B(n65761), .Z(n65763) );
  IV U85975 ( .A(n65763), .Z(n70719) );
  IV U85976 ( .A(n65764), .Z(n65765) );
  NOR U85977 ( .A(n74227), .B(n65765), .Z(n65768) );
  IV U85978 ( .A(n65766), .Z(n65767) );
  NOR U85979 ( .A(n74227), .B(n65767), .Z(n74240) );
  NOR U85980 ( .A(n65768), .B(n74240), .Z(n69150) );
  IV U85981 ( .A(n65769), .Z(n65772) );
  IV U85982 ( .A(n65770), .Z(n65771) );
  NOR U85983 ( .A(n65772), .B(n65771), .Z(n74222) );
  IV U85984 ( .A(n65773), .Z(n65775) );
  XOR U85985 ( .A(n69139), .B(n69140), .Z(n65774) );
  NOR U85986 ( .A(n65775), .B(n65774), .Z(n74219) );
  IV U85987 ( .A(n65776), .Z(n65779) );
  NOR U85988 ( .A(n65777), .B(n69140), .Z(n65778) );
  IV U85989 ( .A(n65778), .Z(n69144) );
  NOR U85990 ( .A(n65779), .B(n69144), .Z(n74216) );
  IV U85991 ( .A(n65780), .Z(n65782) );
  NOR U85992 ( .A(n65782), .B(n65781), .Z(n70732) );
  IV U85993 ( .A(n65783), .Z(n65784) );
  NOR U85994 ( .A(n65785), .B(n65784), .Z(n70735) );
  IV U85995 ( .A(n65786), .Z(n65787) );
  NOR U85996 ( .A(n65787), .B(n69132), .Z(n74182) );
  NOR U85997 ( .A(n70735), .B(n74182), .Z(n65788) );
  IV U85998 ( .A(n65788), .Z(n69130) );
  IV U85999 ( .A(n65789), .Z(n65791) );
  NOR U86000 ( .A(n65791), .B(n65790), .Z(n74172) );
  IV U86001 ( .A(n65792), .Z(n65793) );
  NOR U86002 ( .A(n65793), .B(n69127), .Z(n74169) );
  IV U86003 ( .A(n65794), .Z(n65797) );
  IV U86004 ( .A(n65795), .Z(n65796) );
  NOR U86005 ( .A(n65797), .B(n65796), .Z(n65798) );
  IV U86006 ( .A(n65798), .Z(n74166) );
  IV U86007 ( .A(n65799), .Z(n65800) );
  NOR U86008 ( .A(n65801), .B(n65800), .Z(n79627) );
  IV U86009 ( .A(n65802), .Z(n65804) );
  NOR U86010 ( .A(n65804), .B(n65803), .Z(n76195) );
  NOR U86011 ( .A(n79627), .B(n76195), .Z(n70748) );
  IV U86012 ( .A(n70748), .Z(n69107) );
  IV U86013 ( .A(n65805), .Z(n79607) );
  NOR U86014 ( .A(n65806), .B(n79607), .Z(n65810) );
  IV U86015 ( .A(n65807), .Z(n65809) );
  NOR U86016 ( .A(n65809), .B(n65808), .Z(n79616) );
  NOR U86017 ( .A(n65810), .B(n79616), .Z(n70763) );
  IV U86018 ( .A(n65811), .Z(n65813) );
  IV U86019 ( .A(n65812), .Z(n65818) );
  NOR U86020 ( .A(n65813), .B(n65818), .Z(n70765) );
  IV U86021 ( .A(n65814), .Z(n65815) );
  NOR U86022 ( .A(n79610), .B(n65815), .Z(n70767) );
  NOR U86023 ( .A(n70765), .B(n70767), .Z(n69100) );
  NOR U86024 ( .A(n65816), .B(n70781), .Z(n65820) );
  IV U86025 ( .A(n65817), .Z(n65819) );
  NOR U86026 ( .A(n65819), .B(n65818), .Z(n70772) );
  NOR U86027 ( .A(n65820), .B(n70772), .Z(n69099) );
  IV U86028 ( .A(n65821), .Z(n65823) );
  IV U86029 ( .A(n65822), .Z(n81733) );
  NOR U86030 ( .A(n65823), .B(n81733), .Z(n65824) );
  IV U86031 ( .A(n65824), .Z(n70786) );
  IV U86032 ( .A(n65825), .Z(n65831) );
  NOR U86033 ( .A(n65826), .B(n65831), .Z(n65827) );
  IV U86034 ( .A(n65827), .Z(n74122) );
  NOR U86035 ( .A(n65828), .B(n74122), .Z(n70793) );
  IV U86036 ( .A(n65829), .Z(n65830) );
  NOR U86037 ( .A(n65831), .B(n65830), .Z(n70799) );
  NOR U86038 ( .A(n74120), .B(n70799), .Z(n69079) );
  IV U86039 ( .A(n65832), .Z(n65835) );
  NOR U86040 ( .A(n65833), .B(n69072), .Z(n65834) );
  IV U86041 ( .A(n65834), .Z(n69075) );
  NOR U86042 ( .A(n65835), .B(n69075), .Z(n70802) );
  NOR U86043 ( .A(n65836), .B(n70815), .Z(n65840) );
  NOR U86044 ( .A(n65838), .B(n65837), .Z(n65839) );
  IV U86045 ( .A(n65839), .Z(n70816) );
  NOR U86046 ( .A(n65840), .B(n70816), .Z(n65841) );
  IV U86047 ( .A(n65841), .Z(n70810) );
  IV U86048 ( .A(n65842), .Z(n65843) );
  NOR U86049 ( .A(n65843), .B(n65851), .Z(n70821) );
  IV U86050 ( .A(n65844), .Z(n70820) );
  NOR U86051 ( .A(n70820), .B(n70816), .Z(n65845) );
  NOR U86052 ( .A(n70821), .B(n65845), .Z(n69067) );
  IV U86053 ( .A(n65846), .Z(n65847) );
  NOR U86054 ( .A(n65848), .B(n65847), .Z(n76257) );
  IV U86055 ( .A(n65849), .Z(n65850) );
  NOR U86056 ( .A(n65851), .B(n65850), .Z(n76253) );
  NOR U86057 ( .A(n76257), .B(n76253), .Z(n70826) );
  IV U86058 ( .A(n65852), .Z(n65854) );
  NOR U86059 ( .A(n65854), .B(n65853), .Z(n76265) );
  IV U86060 ( .A(n65855), .Z(n65856) );
  NOR U86061 ( .A(n65857), .B(n65856), .Z(n76260) );
  NOR U86062 ( .A(n76265), .B(n76260), .Z(n70824) );
  IV U86063 ( .A(n65858), .Z(n76278) );
  IV U86064 ( .A(n65859), .Z(n70830) );
  NOR U86065 ( .A(n76278), .B(n70830), .Z(n69062) );
  XOR U86066 ( .A(n65861), .B(n65860), .Z(n65863) );
  XOR U86067 ( .A(n69058), .B(n69059), .Z(n65862) );
  NOR U86068 ( .A(n65863), .B(n65862), .Z(n65864) );
  IV U86069 ( .A(n65864), .Z(n65865) );
  NOR U86070 ( .A(n65866), .B(n65865), .Z(n70833) );
  IV U86071 ( .A(n65867), .Z(n65869) );
  NOR U86072 ( .A(n65869), .B(n65868), .Z(n70840) );
  NOR U86073 ( .A(n65870), .B(n65877), .Z(n65871) );
  IV U86074 ( .A(n65871), .Z(n65872) );
  NOR U86075 ( .A(n65873), .B(n65872), .Z(n65874) );
  IV U86076 ( .A(n65874), .Z(n79550) );
  NOR U86077 ( .A(n65875), .B(n79550), .Z(n70851) );
  NOR U86078 ( .A(n70840), .B(n70851), .Z(n69054) );
  IV U86079 ( .A(n65876), .Z(n65878) );
  NOR U86080 ( .A(n65878), .B(n65877), .Z(n85328) );
  IV U86081 ( .A(n65879), .Z(n65881) );
  NOR U86082 ( .A(n65881), .B(n65880), .Z(n85336) );
  NOR U86083 ( .A(n85328), .B(n85336), .Z(n70846) );
  IV U86084 ( .A(n65882), .Z(n65883) );
  NOR U86085 ( .A(n65884), .B(n65883), .Z(n70859) );
  NOR U86086 ( .A(n65885), .B(n70848), .Z(n65886) );
  NOR U86087 ( .A(n70859), .B(n65886), .Z(n69053) );
  IV U86088 ( .A(n65887), .Z(n65889) );
  IV U86089 ( .A(n65888), .Z(n65891) );
  NOR U86090 ( .A(n65889), .B(n65891), .Z(n70856) );
  IV U86091 ( .A(n65890), .Z(n65892) );
  NOR U86092 ( .A(n65892), .B(n65891), .Z(n70865) );
  IV U86093 ( .A(n65893), .Z(n65894) );
  NOR U86094 ( .A(n69052), .B(n65894), .Z(n70862) );
  IV U86095 ( .A(n65895), .Z(n65896) );
  NOR U86096 ( .A(n65902), .B(n65896), .Z(n76294) );
  IV U86097 ( .A(n65897), .Z(n65899) );
  IV U86098 ( .A(n65898), .Z(n69048) );
  NOR U86099 ( .A(n65899), .B(n69048), .Z(n79513) );
  NOR U86100 ( .A(n76294), .B(n79513), .Z(n70873) );
  IV U86101 ( .A(n65900), .Z(n65901) );
  NOR U86102 ( .A(n65902), .B(n65901), .Z(n70870) );
  IV U86103 ( .A(n65903), .Z(n65905) );
  XOR U86104 ( .A(n65909), .B(n69041), .Z(n65904) );
  NOR U86105 ( .A(n65905), .B(n65904), .Z(n70878) );
  IV U86106 ( .A(n65906), .Z(n65908) );
  NOR U86107 ( .A(n65908), .B(n65907), .Z(n79505) );
  IV U86108 ( .A(n65909), .Z(n65910) );
  NOR U86109 ( .A(n65910), .B(n69041), .Z(n76302) );
  NOR U86110 ( .A(n79505), .B(n76302), .Z(n70887) );
  IV U86111 ( .A(n65911), .Z(n65916) );
  IV U86112 ( .A(n65912), .Z(n65913) );
  NOR U86113 ( .A(n65916), .B(n65913), .Z(n70884) );
  IV U86114 ( .A(n65914), .Z(n65915) );
  NOR U86115 ( .A(n65916), .B(n65915), .Z(n74086) );
  IV U86116 ( .A(n65917), .Z(n65925) );
  IV U86117 ( .A(n65918), .Z(n65919) );
  NOR U86118 ( .A(n65925), .B(n65919), .Z(n70897) );
  IV U86119 ( .A(n65920), .Z(n65922) );
  NOR U86120 ( .A(n65922), .B(n65921), .Z(n70892) );
  NOR U86121 ( .A(n70897), .B(n70892), .Z(n69029) );
  IV U86122 ( .A(n65923), .Z(n65924) );
  NOR U86123 ( .A(n65925), .B(n65924), .Z(n70903) );
  IV U86124 ( .A(n65926), .Z(n65928) );
  NOR U86125 ( .A(n65928), .B(n65927), .Z(n70900) );
  NOR U86126 ( .A(n69024), .B(n65929), .Z(n65930) );
  IV U86127 ( .A(n65930), .Z(n65931) );
  NOR U86128 ( .A(n65932), .B(n65931), .Z(n70909) );
  IV U86129 ( .A(n65933), .Z(n65934) );
  NOR U86130 ( .A(n69024), .B(n65934), .Z(n70906) );
  IV U86131 ( .A(n65935), .Z(n65938) );
  IV U86132 ( .A(n65936), .Z(n65937) );
  NOR U86133 ( .A(n65938), .B(n65937), .Z(n65939) );
  IV U86134 ( .A(n65939), .Z(n74077) );
  IV U86135 ( .A(n65940), .Z(n65943) );
  NOR U86136 ( .A(n65941), .B(n65947), .Z(n65942) );
  IV U86137 ( .A(n65942), .Z(n69020) );
  NOR U86138 ( .A(n65943), .B(n69020), .Z(n70919) );
  IV U86139 ( .A(n65944), .Z(n65946) );
  NOR U86140 ( .A(n65946), .B(n65945), .Z(n70927) );
  NOR U86141 ( .A(n65948), .B(n65947), .Z(n70922) );
  NOR U86142 ( .A(n70927), .B(n70922), .Z(n69017) );
  IV U86143 ( .A(n65949), .Z(n65951) );
  NOR U86144 ( .A(n65951), .B(n65950), .Z(n70925) );
  NOR U86145 ( .A(n70930), .B(n70925), .Z(n69016) );
  IV U86146 ( .A(n65952), .Z(n65953) );
  NOR U86147 ( .A(n65953), .B(n65955), .Z(n74068) );
  IV U86148 ( .A(n65954), .Z(n65956) );
  NOR U86149 ( .A(n65956), .B(n65955), .Z(n74064) );
  NOR U86150 ( .A(n74068), .B(n74064), .Z(n69015) );
  IV U86151 ( .A(n65957), .Z(n65958) );
  IV U86152 ( .A(n79418), .Z(n65962) );
  NOR U86153 ( .A(n65958), .B(n65962), .Z(n74062) );
  IV U86154 ( .A(n65959), .Z(n65960) );
  NOR U86155 ( .A(n65960), .B(n65965), .Z(n74059) );
  IV U86156 ( .A(n65961), .Z(n79419) );
  NOR U86157 ( .A(n79419), .B(n65962), .Z(n74057) );
  NOR U86158 ( .A(n74059), .B(n74057), .Z(n69013) );
  IV U86159 ( .A(n65966), .Z(n65963) );
  NOR U86160 ( .A(n65963), .B(n65965), .Z(n76327) );
  IV U86161 ( .A(n65964), .Z(n65968) );
  XOR U86162 ( .A(n65966), .B(n65965), .Z(n65967) );
  NOR U86163 ( .A(n65968), .B(n65967), .Z(n76323) );
  NOR U86164 ( .A(n76327), .B(n76323), .Z(n70936) );
  IV U86165 ( .A(n65969), .Z(n65973) );
  NOR U86166 ( .A(n65971), .B(n65970), .Z(n65972) );
  IV U86167 ( .A(n65972), .Z(n69011) );
  NOR U86168 ( .A(n65973), .B(n69011), .Z(n70933) );
  IV U86169 ( .A(n65974), .Z(n65976) );
  IV U86170 ( .A(n65975), .Z(n65978) );
  NOR U86171 ( .A(n65976), .B(n65978), .Z(n70939) );
  IV U86172 ( .A(n65977), .Z(n65979) );
  NOR U86173 ( .A(n65979), .B(n65978), .Z(n74051) );
  IV U86174 ( .A(n65980), .Z(n65981) );
  NOR U86175 ( .A(n65981), .B(n65984), .Z(n74048) );
  IV U86176 ( .A(n65982), .Z(n65983) );
  NOR U86177 ( .A(n65984), .B(n65983), .Z(n70945) );
  IV U86178 ( .A(n65985), .Z(n65989) );
  NOR U86179 ( .A(n65987), .B(n65986), .Z(n65988) );
  IV U86180 ( .A(n65988), .Z(n65991) );
  NOR U86181 ( .A(n65989), .B(n65991), .Z(n70951) );
  IV U86182 ( .A(n65990), .Z(n65992) );
  NOR U86183 ( .A(n65992), .B(n65991), .Z(n70948) );
  IV U86184 ( .A(n65993), .Z(n68999) );
  IV U86185 ( .A(n65994), .Z(n65995) );
  NOR U86186 ( .A(n68999), .B(n65995), .Z(n70957) );
  IV U86187 ( .A(n65996), .Z(n65999) );
  IV U86188 ( .A(n65997), .Z(n65998) );
  NOR U86189 ( .A(n65999), .B(n65998), .Z(n66000) );
  IV U86190 ( .A(n66000), .Z(n69004) );
  IV U86191 ( .A(n66001), .Z(n66002) );
  NOR U86192 ( .A(n66003), .B(n66002), .Z(n70978) );
  IV U86193 ( .A(n66004), .Z(n66006) );
  NOR U86194 ( .A(n66006), .B(n66005), .Z(n70980) );
  NOR U86195 ( .A(n70978), .B(n70980), .Z(n66007) );
  IV U86196 ( .A(n66007), .Z(n68984) );
  IV U86197 ( .A(n66008), .Z(n66011) );
  IV U86198 ( .A(n66009), .Z(n66010) );
  NOR U86199 ( .A(n66011), .B(n66010), .Z(n66012) );
  IV U86200 ( .A(n66012), .Z(n70993) );
  IV U86201 ( .A(n66013), .Z(n66014) );
  NOR U86202 ( .A(n66015), .B(n66014), .Z(n70995) );
  NOR U86203 ( .A(n71001), .B(n70995), .Z(n68970) );
  IV U86204 ( .A(n66016), .Z(n66017) );
  NOR U86205 ( .A(n66020), .B(n66017), .Z(n71004) );
  IV U86206 ( .A(n66018), .Z(n66022) );
  NOR U86207 ( .A(n66020), .B(n66019), .Z(n66021) );
  IV U86208 ( .A(n66021), .Z(n66024) );
  NOR U86209 ( .A(n66022), .B(n66024), .Z(n74022) );
  IV U86210 ( .A(n66023), .Z(n66025) );
  NOR U86211 ( .A(n66025), .B(n66024), .Z(n74004) );
  IV U86212 ( .A(n66026), .Z(n66028) );
  NOR U86213 ( .A(n66028), .B(n66027), .Z(n74010) );
  IV U86214 ( .A(n66029), .Z(n66033) );
  NOR U86215 ( .A(n66030), .B(n66033), .Z(n66031) );
  IV U86216 ( .A(n66031), .Z(n90900) );
  NOR U86217 ( .A(n90897), .B(n90900), .Z(n71008) );
  IV U86218 ( .A(n66032), .Z(n66034) );
  NOR U86219 ( .A(n66034), .B(n66033), .Z(n73995) );
  NOR U86220 ( .A(n66035), .B(n73995), .Z(n68944) );
  NOR U86221 ( .A(n66037), .B(n66036), .Z(n71013) );
  IV U86222 ( .A(n66038), .Z(n66039) );
  NOR U86223 ( .A(n66039), .B(n68941), .Z(n73976) );
  IV U86224 ( .A(n66040), .Z(n68938) );
  IV U86225 ( .A(n66041), .Z(n66042) );
  NOR U86226 ( .A(n68938), .B(n66042), .Z(n85171) );
  NOR U86227 ( .A(n81943), .B(n85171), .Z(n73971) );
  IV U86228 ( .A(n66043), .Z(n66044) );
  NOR U86229 ( .A(n66045), .B(n66044), .Z(n71025) );
  IV U86230 ( .A(n66046), .Z(n66049) );
  NOR U86231 ( .A(n66055), .B(n66047), .Z(n66048) );
  IV U86232 ( .A(n66048), .Z(n66051) );
  NOR U86233 ( .A(n66049), .B(n66051), .Z(n71022) );
  IV U86234 ( .A(n66050), .Z(n66052) );
  NOR U86235 ( .A(n66052), .B(n66051), .Z(n73964) );
  IV U86236 ( .A(n66053), .Z(n66057) );
  NOR U86237 ( .A(n66055), .B(n66054), .Z(n66056) );
  IV U86238 ( .A(n66056), .Z(n66059) );
  NOR U86239 ( .A(n66057), .B(n66059), .Z(n73961) );
  IV U86240 ( .A(n66058), .Z(n66060) );
  NOR U86241 ( .A(n66060), .B(n66059), .Z(n71031) );
  IV U86242 ( .A(n66061), .Z(n66064) );
  IV U86243 ( .A(n66062), .Z(n66063) );
  NOR U86244 ( .A(n66064), .B(n66063), .Z(n71028) );
  XOR U86245 ( .A(n66065), .B(n66078), .Z(n66068) );
  IV U86246 ( .A(n66066), .Z(n66067) );
  NOR U86247 ( .A(n66068), .B(n66067), .Z(n73958) );
  IV U86248 ( .A(n66069), .Z(n66072) );
  NOR U86249 ( .A(n66078), .B(n66070), .Z(n66071) );
  IV U86250 ( .A(n66071), .Z(n66074) );
  NOR U86251 ( .A(n66072), .B(n66074), .Z(n73955) );
  IV U86252 ( .A(n66073), .Z(n66075) );
  NOR U86253 ( .A(n66075), .B(n66074), .Z(n71034) );
  IV U86254 ( .A(n66076), .Z(n66080) );
  NOR U86255 ( .A(n66078), .B(n66077), .Z(n66079) );
  IV U86256 ( .A(n66079), .Z(n66082) );
  NOR U86257 ( .A(n66080), .B(n66082), .Z(n71037) );
  IV U86258 ( .A(n66081), .Z(n66083) );
  NOR U86259 ( .A(n66083), .B(n66082), .Z(n73943) );
  IV U86260 ( .A(n66084), .Z(n66085) );
  NOR U86261 ( .A(n66085), .B(n66088), .Z(n71043) );
  IV U86262 ( .A(n66086), .Z(n66087) );
  NOR U86263 ( .A(n66087), .B(n66088), .Z(n71040) );
  NOR U86264 ( .A(n66089), .B(n66088), .Z(n73936) );
  IV U86265 ( .A(n66090), .Z(n66092) );
  NOR U86266 ( .A(n66092), .B(n66091), .Z(n73933) );
  IV U86267 ( .A(n66093), .Z(n71048) );
  IV U86268 ( .A(n66094), .Z(n66095) );
  NOR U86269 ( .A(n66095), .B(n66098), .Z(n71055) );
  IV U86270 ( .A(n66096), .Z(n66097) );
  NOR U86271 ( .A(n66098), .B(n66097), .Z(n71061) );
  IV U86272 ( .A(n66099), .Z(n66108) );
  IV U86273 ( .A(n66100), .Z(n66101) );
  NOR U86274 ( .A(n66108), .B(n66101), .Z(n79303) );
  IV U86275 ( .A(n66102), .Z(n66104) );
  NOR U86276 ( .A(n66104), .B(n66103), .Z(n73921) );
  NOR U86277 ( .A(n79303), .B(n73921), .Z(n66105) );
  IV U86278 ( .A(n66105), .Z(n68920) );
  IV U86279 ( .A(n66106), .Z(n66107) );
  NOR U86280 ( .A(n66108), .B(n66107), .Z(n79297) );
  IV U86281 ( .A(n66109), .Z(n66111) );
  NOR U86282 ( .A(n66111), .B(n66110), .Z(n73915) );
  IV U86283 ( .A(n66112), .Z(n66113) );
  NOR U86284 ( .A(n66116), .B(n66113), .Z(n73912) );
  IV U86285 ( .A(n66114), .Z(n66115) );
  NOR U86286 ( .A(n66116), .B(n66115), .Z(n71068) );
  IV U86287 ( .A(n66117), .Z(n66119) );
  NOR U86288 ( .A(n66119), .B(n66118), .Z(n71065) );
  NOR U86289 ( .A(n66121), .B(n66120), .Z(n76436) );
  NOR U86290 ( .A(n66123), .B(n66122), .Z(n76432) );
  NOR U86291 ( .A(n76436), .B(n76432), .Z(n73900) );
  IV U86292 ( .A(n66124), .Z(n66125) );
  NOR U86293 ( .A(n66126), .B(n66125), .Z(n76453) );
  IV U86294 ( .A(n66127), .Z(n66129) );
  NOR U86295 ( .A(n66129), .B(n66128), .Z(n76447) );
  NOR U86296 ( .A(n76453), .B(n76447), .Z(n73890) );
  IV U86297 ( .A(n66130), .Z(n66132) );
  NOR U86298 ( .A(n66132), .B(n66131), .Z(n73887) );
  IV U86299 ( .A(n66133), .Z(n66134) );
  NOR U86300 ( .A(n66134), .B(n68894), .Z(n68888) );
  IV U86301 ( .A(n68888), .Z(n68882) );
  IV U86302 ( .A(n66135), .Z(n66136) );
  NOR U86303 ( .A(n66137), .B(n66136), .Z(n73877) );
  IV U86304 ( .A(n66138), .Z(n66140) );
  NOR U86305 ( .A(n66140), .B(n66139), .Z(n79254) );
  IV U86306 ( .A(n66141), .Z(n66143) );
  NOR U86307 ( .A(n66143), .B(n66142), .Z(n79259) );
  NOR U86308 ( .A(n79254), .B(n79259), .Z(n73876) );
  IV U86309 ( .A(n66144), .Z(n73852) );
  NOR U86310 ( .A(n66145), .B(n73852), .Z(n66147) );
  NOR U86311 ( .A(n73859), .B(n73857), .Z(n66146) );
  NOR U86312 ( .A(n66147), .B(n66146), .Z(n68880) );
  IV U86313 ( .A(n66148), .Z(n66152) );
  NOR U86314 ( .A(n66150), .B(n66149), .Z(n66151) );
  IV U86315 ( .A(n66151), .Z(n66154) );
  NOR U86316 ( .A(n66152), .B(n66154), .Z(n73861) );
  IV U86317 ( .A(n66153), .Z(n66155) );
  NOR U86318 ( .A(n66155), .B(n66154), .Z(n66156) );
  IV U86319 ( .A(n66156), .Z(n73848) );
  IV U86320 ( .A(n66157), .Z(n66158) );
  NOR U86321 ( .A(n68867), .B(n66158), .Z(n71090) );
  IV U86322 ( .A(n66159), .Z(n66162) );
  IV U86323 ( .A(n66160), .Z(n66161) );
  NOR U86324 ( .A(n66162), .B(n66161), .Z(n66163) );
  IV U86325 ( .A(n66163), .Z(n68868) );
  NOR U86326 ( .A(n66165), .B(n66164), .Z(n71098) );
  IV U86327 ( .A(n66166), .Z(n66167) );
  NOR U86328 ( .A(n73837), .B(n66167), .Z(n73818) );
  NOR U86329 ( .A(n66169), .B(n66168), .Z(n66170) );
  NOR U86330 ( .A(n73818), .B(n66170), .Z(n71102) );
  IV U86331 ( .A(n66171), .Z(n66172) );
  NOR U86332 ( .A(n68846), .B(n66172), .Z(n71111) );
  IV U86333 ( .A(n66173), .Z(n66175) );
  NOR U86334 ( .A(n66175), .B(n66174), .Z(n73805) );
  NOR U86335 ( .A(n66177), .B(n66176), .Z(n73791) );
  IV U86336 ( .A(n66178), .Z(n68827) );
  IV U86337 ( .A(n66179), .Z(n66180) );
  NOR U86338 ( .A(n68827), .B(n66180), .Z(n71125) );
  NOR U86339 ( .A(n73791), .B(n71125), .Z(n68828) );
  IV U86340 ( .A(n66181), .Z(n66183) );
  NOR U86341 ( .A(n66183), .B(n66182), .Z(n71127) );
  IV U86342 ( .A(n66184), .Z(n66185) );
  NOR U86343 ( .A(n66185), .B(n68820), .Z(n73777) );
  NOR U86344 ( .A(n71127), .B(n73777), .Z(n68818) );
  IV U86345 ( .A(n66186), .Z(n66192) );
  NOR U86346 ( .A(n66187), .B(n68809), .Z(n66188) );
  IV U86347 ( .A(n66188), .Z(n66189) );
  NOR U86348 ( .A(n66190), .B(n66189), .Z(n66191) );
  IV U86349 ( .A(n66191), .Z(n68815) );
  NOR U86350 ( .A(n66192), .B(n68815), .Z(n71129) );
  IV U86351 ( .A(n66193), .Z(n66198) );
  IV U86352 ( .A(n66194), .Z(n66196) );
  NOR U86353 ( .A(n66196), .B(n66195), .Z(n66197) );
  IV U86354 ( .A(n66197), .Z(n66200) );
  NOR U86355 ( .A(n66198), .B(n66200), .Z(n73758) );
  IV U86356 ( .A(n66199), .Z(n66201) );
  NOR U86357 ( .A(n66201), .B(n66200), .Z(n71132) );
  IV U86358 ( .A(n66202), .Z(n66206) );
  IV U86359 ( .A(n66203), .Z(n66209) );
  NOR U86360 ( .A(n66209), .B(n66204), .Z(n66205) );
  IV U86361 ( .A(n66205), .Z(n66212) );
  NOR U86362 ( .A(n66206), .B(n66212), .Z(n71137) );
  IV U86363 ( .A(n66207), .Z(n66208) );
  NOR U86364 ( .A(n66209), .B(n66208), .Z(n71135) );
  NOR U86365 ( .A(n71137), .B(n71135), .Z(n66210) );
  IV U86366 ( .A(n66210), .Z(n68806) );
  IV U86367 ( .A(n66211), .Z(n66213) );
  NOR U86368 ( .A(n66213), .B(n66212), .Z(n73754) );
  IV U86369 ( .A(n66214), .Z(n66215) );
  NOR U86370 ( .A(n66215), .B(n68800), .Z(n73751) );
  IV U86371 ( .A(n66216), .Z(n66220) );
  IV U86372 ( .A(n66217), .Z(n68804) );
  NOR U86373 ( .A(n68804), .B(n66218), .Z(n66219) );
  IV U86374 ( .A(n66219), .Z(n68797) );
  NOR U86375 ( .A(n66220), .B(n68797), .Z(n73740) );
  IV U86376 ( .A(n66221), .Z(n66222) );
  NOR U86377 ( .A(n66222), .B(n68789), .Z(n66223) );
  IV U86378 ( .A(n66223), .Z(n73739) );
  IV U86379 ( .A(n66224), .Z(n66226) );
  NOR U86380 ( .A(n66226), .B(n66225), .Z(n66227) );
  IV U86381 ( .A(n66227), .Z(n68791) );
  IV U86382 ( .A(n66228), .Z(n68787) );
  IV U86383 ( .A(n66229), .Z(n66230) );
  NOR U86384 ( .A(n68787), .B(n66230), .Z(n71142) );
  IV U86385 ( .A(n66231), .Z(n66232) );
  NOR U86386 ( .A(n66232), .B(n68784), .Z(n71150) );
  IV U86387 ( .A(n66235), .Z(n66233) );
  NOR U86388 ( .A(n68781), .B(n66233), .Z(n79139) );
  IV U86389 ( .A(n66234), .Z(n66237) );
  XOR U86390 ( .A(n66235), .B(n68781), .Z(n66236) );
  NOR U86391 ( .A(n66237), .B(n66236), .Z(n79148) );
  NOR U86392 ( .A(n79139), .B(n79148), .Z(n71154) );
  IV U86393 ( .A(n66238), .Z(n66240) );
  IV U86394 ( .A(n66239), .Z(n68767) );
  NOR U86395 ( .A(n66240), .B(n68767), .Z(n71158) );
  IV U86396 ( .A(n66241), .Z(n66243) );
  IV U86397 ( .A(n66242), .Z(n68752) );
  NOR U86398 ( .A(n66243), .B(n68752), .Z(n73717) );
  IV U86399 ( .A(n66244), .Z(n66245) );
  IV U86400 ( .A(n68745), .Z(n71170) );
  NOR U86401 ( .A(n66245), .B(n71170), .Z(n66248) );
  NOR U86402 ( .A(n66246), .B(n73711), .Z(n66247) );
  NOR U86403 ( .A(n66248), .B(n66247), .Z(n68750) );
  IV U86404 ( .A(n66249), .Z(n66252) );
  NOR U86405 ( .A(n68739), .B(n66250), .Z(n66251) );
  IV U86406 ( .A(n66251), .Z(n68741) );
  NOR U86407 ( .A(n66252), .B(n68741), .Z(n71187) );
  NOR U86408 ( .A(n66253), .B(n68732), .Z(n73700) );
  IV U86409 ( .A(n66254), .Z(n66256) );
  NOR U86410 ( .A(n66256), .B(n66255), .Z(n84888) );
  IV U86411 ( .A(n68735), .Z(n66257) );
  NOR U86412 ( .A(n66257), .B(n68732), .Z(n84896) );
  NOR U86413 ( .A(n84888), .B(n84896), .Z(n73686) );
  IV U86414 ( .A(n66258), .Z(n66259) );
  NOR U86415 ( .A(n66259), .B(n68721), .Z(n71206) );
  NOR U86416 ( .A(n66261), .B(n66260), .Z(n66262) );
  IV U86417 ( .A(n66262), .Z(n66269) );
  XOR U86418 ( .A(n66264), .B(n66263), .Z(n66266) );
  NOR U86419 ( .A(n66266), .B(n66265), .Z(n66267) );
  IV U86420 ( .A(n66267), .Z(n66268) );
  NOR U86421 ( .A(n66269), .B(n66268), .Z(n73674) );
  IV U86422 ( .A(n66270), .Z(n66271) );
  NOR U86423 ( .A(n66271), .B(n68709), .Z(n66272) );
  IV U86424 ( .A(n66272), .Z(n71228) );
  IV U86425 ( .A(n66273), .Z(n66280) );
  IV U86426 ( .A(n66274), .Z(n66275) );
  NOR U86427 ( .A(n66280), .B(n66275), .Z(n71236) );
  IV U86428 ( .A(n66276), .Z(n66277) );
  NOR U86429 ( .A(n66277), .B(n68709), .Z(n71234) );
  NOR U86430 ( .A(n71236), .B(n71234), .Z(n68702) );
  IV U86431 ( .A(n66278), .Z(n66279) );
  NOR U86432 ( .A(n66280), .B(n66279), .Z(n73665) );
  IV U86433 ( .A(n66281), .Z(n66282) );
  NOR U86434 ( .A(n66282), .B(n66287), .Z(n73662) );
  IV U86435 ( .A(n66283), .Z(n66285) );
  NOR U86436 ( .A(n66285), .B(n66284), .Z(n71242) );
  IV U86437 ( .A(n66286), .Z(n66288) );
  NOR U86438 ( .A(n66288), .B(n66287), .Z(n71240) );
  NOR U86439 ( .A(n71242), .B(n71240), .Z(n68701) );
  IV U86440 ( .A(n66289), .Z(n66290) );
  NOR U86441 ( .A(n66291), .B(n66290), .Z(n71245) );
  IV U86442 ( .A(n66292), .Z(n66297) );
  IV U86443 ( .A(n66293), .Z(n66294) );
  NOR U86444 ( .A(n66297), .B(n66294), .Z(n73659) );
  NOR U86445 ( .A(n71245), .B(n73659), .Z(n68700) );
  IV U86446 ( .A(n66295), .Z(n66296) );
  NOR U86447 ( .A(n66297), .B(n66296), .Z(n73656) );
  IV U86448 ( .A(n66298), .Z(n66299) );
  NOR U86449 ( .A(n66300), .B(n66299), .Z(n66301) );
  IV U86450 ( .A(n66301), .Z(n73652) );
  IV U86451 ( .A(n66302), .Z(n68676) );
  IV U86452 ( .A(n66303), .Z(n68682) );
  NOR U86453 ( .A(n68676), .B(n68682), .Z(n68675) );
  IV U86454 ( .A(n66304), .Z(n66305) );
  NOR U86455 ( .A(n66305), .B(n68666), .Z(n73630) );
  IV U86456 ( .A(n66306), .Z(n66307) );
  NOR U86457 ( .A(n66307), .B(n66313), .Z(n79020) );
  IV U86458 ( .A(n66308), .Z(n66311) );
  IV U86459 ( .A(n66309), .Z(n66310) );
  NOR U86460 ( .A(n66311), .B(n66310), .Z(n76623) );
  NOR U86461 ( .A(n79020), .B(n76623), .Z(n73629) );
  IV U86462 ( .A(n66312), .Z(n66314) );
  NOR U86463 ( .A(n66314), .B(n66313), .Z(n73621) );
  IV U86464 ( .A(n66315), .Z(n66317) );
  IV U86465 ( .A(n66316), .Z(n68656) );
  NOR U86466 ( .A(n66317), .B(n68656), .Z(n73607) );
  NOR U86467 ( .A(n73605), .B(n73607), .Z(n68651) );
  IV U86468 ( .A(n66318), .Z(n66320) );
  NOR U86469 ( .A(n66320), .B(n66319), .Z(n73602) );
  IV U86470 ( .A(n66321), .Z(n66326) );
  IV U86471 ( .A(n66322), .Z(n66323) );
  NOR U86472 ( .A(n66323), .B(n66335), .Z(n66324) );
  IV U86473 ( .A(n66324), .Z(n66325) );
  NOR U86474 ( .A(n66326), .B(n66325), .Z(n71267) );
  IV U86475 ( .A(n66327), .Z(n66331) );
  NOR U86476 ( .A(n66328), .B(n66335), .Z(n66329) );
  IV U86477 ( .A(n66329), .Z(n66330) );
  NOR U86478 ( .A(n66331), .B(n66330), .Z(n71264) );
  IV U86479 ( .A(n66332), .Z(n66333) );
  NOR U86480 ( .A(n66333), .B(n66341), .Z(n73594) );
  IV U86481 ( .A(n66334), .Z(n66336) );
  NOR U86482 ( .A(n66336), .B(n66335), .Z(n71271) );
  NOR U86483 ( .A(n73594), .B(n71271), .Z(n68650) );
  IV U86484 ( .A(n66337), .Z(n66339) );
  NOR U86485 ( .A(n66339), .B(n66338), .Z(n71276) );
  IV U86486 ( .A(n66340), .Z(n66342) );
  NOR U86487 ( .A(n66342), .B(n66341), .Z(n73597) );
  NOR U86488 ( .A(n71276), .B(n73597), .Z(n68649) );
  IV U86489 ( .A(n66343), .Z(n66344) );
  NOR U86490 ( .A(n66344), .B(n68643), .Z(n71273) );
  IV U86491 ( .A(n66345), .Z(n66346) );
  NOR U86492 ( .A(n66347), .B(n66346), .Z(n68640) );
  IV U86493 ( .A(n68640), .Z(n68634) );
  IV U86494 ( .A(n66348), .Z(n66350) );
  NOR U86495 ( .A(n66350), .B(n66349), .Z(n71285) );
  IV U86496 ( .A(n66351), .Z(n66352) );
  NOR U86497 ( .A(n66354), .B(n66352), .Z(n73578) );
  IV U86498 ( .A(n66353), .Z(n66355) );
  NOR U86499 ( .A(n66355), .B(n66354), .Z(n73575) );
  IV U86500 ( .A(n66356), .Z(n66358) );
  NOR U86501 ( .A(n66358), .B(n66357), .Z(n68619) );
  IV U86502 ( .A(n68619), .Z(n68612) );
  IV U86503 ( .A(n66359), .Z(n66360) );
  NOR U86504 ( .A(n66360), .B(n68614), .Z(n68609) );
  IV U86505 ( .A(n68609), .Z(n68604) );
  IV U86506 ( .A(n66361), .Z(n66365) );
  IV U86507 ( .A(n66362), .Z(n68597) );
  NOR U86508 ( .A(n66363), .B(n68597), .Z(n66364) );
  IV U86509 ( .A(n66364), .Z(n68601) );
  NOR U86510 ( .A(n66365), .B(n68601), .Z(n71294) );
  IV U86511 ( .A(n66366), .Z(n66367) );
  NOR U86512 ( .A(n66368), .B(n66367), .Z(n78982) );
  IV U86513 ( .A(n66369), .Z(n66370) );
  NOR U86514 ( .A(n66370), .B(n68594), .Z(n76695) );
  NOR U86515 ( .A(n78982), .B(n76695), .Z(n71299) );
  IV U86516 ( .A(n66371), .Z(n66373) );
  NOR U86517 ( .A(n66373), .B(n66372), .Z(n71307) );
  IV U86518 ( .A(n66374), .Z(n66377) );
  NOR U86519 ( .A(n66375), .B(n66383), .Z(n66376) );
  IV U86520 ( .A(n66376), .Z(n66379) );
  NOR U86521 ( .A(n66377), .B(n66379), .Z(n71304) );
  IV U86522 ( .A(n66378), .Z(n66380) );
  NOR U86523 ( .A(n66380), .B(n66379), .Z(n71310) );
  IV U86524 ( .A(n66381), .Z(n66382) );
  NOR U86525 ( .A(n66383), .B(n66382), .Z(n73548) );
  IV U86526 ( .A(n66384), .Z(n66385) );
  NOR U86527 ( .A(n66385), .B(n66390), .Z(n73543) );
  IV U86528 ( .A(n66386), .Z(n66388) );
  IV U86529 ( .A(n66387), .Z(n68589) );
  NOR U86530 ( .A(n66388), .B(n68589), .Z(n73534) );
  NOR U86531 ( .A(n73543), .B(n73534), .Z(n68586) );
  IV U86532 ( .A(n66389), .Z(n66391) );
  NOR U86533 ( .A(n66391), .B(n66390), .Z(n73529) );
  IV U86534 ( .A(n66392), .Z(n66397) );
  IV U86535 ( .A(n66393), .Z(n66394) );
  NOR U86536 ( .A(n66397), .B(n66394), .Z(n71313) );
  IV U86537 ( .A(n66395), .Z(n66396) );
  NOR U86538 ( .A(n66397), .B(n66396), .Z(n71320) );
  IV U86539 ( .A(n66398), .Z(n66399) );
  NOR U86540 ( .A(n66400), .B(n66399), .Z(n71327) );
  IV U86541 ( .A(n66401), .Z(n66405) );
  IV U86542 ( .A(n66402), .Z(n66412) );
  NOR U86543 ( .A(n66403), .B(n66412), .Z(n66404) );
  IV U86544 ( .A(n66404), .Z(n66407) );
  NOR U86545 ( .A(n66405), .B(n66407), .Z(n71335) );
  IV U86546 ( .A(n66406), .Z(n66408) );
  NOR U86547 ( .A(n66408), .B(n66407), .Z(n71332) );
  IV U86548 ( .A(n66409), .Z(n66410) );
  NOR U86549 ( .A(n66416), .B(n66410), .Z(n73517) );
  IV U86550 ( .A(n66411), .Z(n66413) );
  NOR U86551 ( .A(n66413), .B(n66412), .Z(n73512) );
  NOR U86552 ( .A(n73517), .B(n73512), .Z(n68574) );
  IV U86553 ( .A(n66414), .Z(n66415) );
  NOR U86554 ( .A(n66416), .B(n66415), .Z(n73508) );
  IV U86555 ( .A(n66417), .Z(n66419) );
  IV U86556 ( .A(n66418), .Z(n66423) );
  NOR U86557 ( .A(n66419), .B(n66423), .Z(n73506) );
  IV U86558 ( .A(n66420), .Z(n66421) );
  NOR U86559 ( .A(n66427), .B(n66421), .Z(n73503) );
  IV U86560 ( .A(n66422), .Z(n66424) );
  NOR U86561 ( .A(n66424), .B(n66423), .Z(n71338) );
  NOR U86562 ( .A(n73503), .B(n71338), .Z(n68572) );
  IV U86563 ( .A(n66425), .Z(n66426) );
  NOR U86564 ( .A(n66427), .B(n66426), .Z(n73500) );
  IV U86565 ( .A(n66428), .Z(n66430) );
  IV U86566 ( .A(n66429), .Z(n68568) );
  NOR U86567 ( .A(n66430), .B(n68568), .Z(n71340) );
  NOR U86568 ( .A(n73500), .B(n71340), .Z(n68571) );
  IV U86569 ( .A(n71350), .Z(n66432) );
  NOR U86570 ( .A(n66432), .B(n66431), .Z(n66433) );
  IV U86571 ( .A(n66433), .Z(n68552) );
  IV U86572 ( .A(n66434), .Z(n66435) );
  NOR U86573 ( .A(n66435), .B(n66437), .Z(n71369) );
  IV U86574 ( .A(n66436), .Z(n66438) );
  NOR U86575 ( .A(n66438), .B(n66437), .Z(n71367) );
  NOR U86576 ( .A(n71369), .B(n71367), .Z(n68547) );
  IV U86577 ( .A(n66439), .Z(n71373) );
  NOR U86578 ( .A(n71373), .B(n66440), .Z(n66444) );
  IV U86579 ( .A(n66441), .Z(n66443) );
  NOR U86580 ( .A(n66443), .B(n66442), .Z(n71376) );
  NOR U86581 ( .A(n66444), .B(n71376), .Z(n68545) );
  IV U86582 ( .A(n66445), .Z(n66446) );
  NOR U86583 ( .A(n66446), .B(n68535), .Z(n66447) );
  IV U86584 ( .A(n66447), .Z(n71384) );
  IV U86585 ( .A(n66448), .Z(n66449) );
  NOR U86586 ( .A(n66450), .B(n66449), .Z(n66451) );
  IV U86587 ( .A(n66451), .Z(n68540) );
  IV U86588 ( .A(n66452), .Z(n66453) );
  NOR U86589 ( .A(n66453), .B(n68529), .Z(n71393) );
  IV U86590 ( .A(n66454), .Z(n66458) );
  NOR U86591 ( .A(n66456), .B(n66455), .Z(n66457) );
  IV U86592 ( .A(n66457), .Z(n68523) );
  NOR U86593 ( .A(n66458), .B(n68523), .Z(n71404) );
  IV U86594 ( .A(n66459), .Z(n66460) );
  NOR U86595 ( .A(n66460), .B(n73468), .Z(n66461) );
  IV U86596 ( .A(n66461), .Z(n73466) );
  NOR U86597 ( .A(n66466), .B(n73466), .Z(n66465) );
  IV U86598 ( .A(n66462), .Z(n66463) );
  NOR U86599 ( .A(n66463), .B(n73468), .Z(n66464) );
  NOR U86600 ( .A(n66465), .B(n66464), .Z(n68520) );
  IV U86601 ( .A(n66466), .Z(n66470) );
  NOR U86602 ( .A(n66467), .B(n73468), .Z(n66468) );
  IV U86603 ( .A(n66468), .Z(n66469) );
  NOR U86604 ( .A(n66470), .B(n66469), .Z(n66471) );
  IV U86605 ( .A(n66471), .Z(n76787) );
  IV U86606 ( .A(n66472), .Z(n66473) );
  NOR U86607 ( .A(n71413), .B(n66473), .Z(n73457) );
  IV U86608 ( .A(n66474), .Z(n66475) );
  NOR U86609 ( .A(n66476), .B(n66475), .Z(n71410) );
  NOR U86610 ( .A(n73457), .B(n71410), .Z(n68519) );
  NOR U86611 ( .A(n66477), .B(n71413), .Z(n68518) );
  IV U86612 ( .A(n66478), .Z(n66480) );
  NOR U86613 ( .A(n66480), .B(n66479), .Z(n71422) );
  IV U86614 ( .A(n66481), .Z(n66483) );
  NOR U86615 ( .A(n66483), .B(n66482), .Z(n71419) );
  NOR U86616 ( .A(n71422), .B(n71419), .Z(n68517) );
  NOR U86617 ( .A(n66484), .B(n68507), .Z(n68504) );
  IV U86618 ( .A(n66485), .Z(n66486) );
  NOR U86619 ( .A(n66487), .B(n66486), .Z(n71430) );
  IV U86620 ( .A(n66488), .Z(n66489) );
  NOR U86621 ( .A(n66489), .B(n68485), .Z(n73448) );
  IV U86622 ( .A(n66490), .Z(n66494) );
  NOR U86623 ( .A(n66491), .B(n68485), .Z(n66492) );
  IV U86624 ( .A(n66492), .Z(n66493) );
  NOR U86625 ( .A(n66494), .B(n66493), .Z(n73441) );
  IV U86626 ( .A(n66495), .Z(n66496) );
  NOR U86627 ( .A(n68482), .B(n66496), .Z(n73438) );
  IV U86628 ( .A(n66497), .Z(n66498) );
  NOR U86629 ( .A(n66498), .B(n68474), .Z(n71451) );
  IV U86630 ( .A(n66499), .Z(n66500) );
  NOR U86631 ( .A(n66500), .B(n68474), .Z(n73430) );
  IV U86632 ( .A(n66501), .Z(n66502) );
  NOR U86633 ( .A(n66503), .B(n66502), .Z(n73420) );
  IV U86634 ( .A(n66504), .Z(n66505) );
  NOR U86635 ( .A(n68465), .B(n66505), .Z(n73423) );
  NOR U86636 ( .A(n73420), .B(n73423), .Z(n68461) );
  IV U86637 ( .A(n66506), .Z(n66513) );
  IV U86638 ( .A(n66507), .Z(n66508) );
  NOR U86639 ( .A(n66513), .B(n66508), .Z(n66509) );
  IV U86640 ( .A(n66509), .Z(n73412) );
  NOR U86641 ( .A(n66511), .B(n66510), .Z(n73405) );
  IV U86642 ( .A(n66512), .Z(n66514) );
  NOR U86643 ( .A(n66514), .B(n66513), .Z(n73408) );
  NOR U86644 ( .A(n73405), .B(n73408), .Z(n68453) );
  IV U86645 ( .A(n66515), .Z(n66517) );
  IV U86646 ( .A(n66516), .Z(n66519) );
  NOR U86647 ( .A(n66517), .B(n66519), .Z(n73402) );
  IV U86648 ( .A(n66518), .Z(n66520) );
  NOR U86649 ( .A(n66520), .B(n66519), .Z(n73398) );
  IV U86650 ( .A(n66521), .Z(n66524) );
  NOR U86651 ( .A(n66530), .B(n66522), .Z(n66523) );
  IV U86652 ( .A(n66523), .Z(n66526) );
  NOR U86653 ( .A(n66524), .B(n66526), .Z(n73395) );
  IV U86654 ( .A(n66525), .Z(n66527) );
  NOR U86655 ( .A(n66527), .B(n66526), .Z(n73391) );
  IV U86656 ( .A(n66528), .Z(n66529) );
  NOR U86657 ( .A(n66530), .B(n66529), .Z(n73388) );
  IV U86658 ( .A(n66531), .Z(n66535) );
  NOR U86659 ( .A(n66533), .B(n66532), .Z(n66534) );
  IV U86660 ( .A(n66534), .Z(n66537) );
  NOR U86661 ( .A(n66535), .B(n66537), .Z(n73384) );
  IV U86662 ( .A(n66536), .Z(n66538) );
  NOR U86663 ( .A(n66538), .B(n66537), .Z(n73381) );
  NOR U86664 ( .A(n68442), .B(n66539), .Z(n66540) );
  IV U86665 ( .A(n66540), .Z(n71474) );
  IV U86666 ( .A(n66541), .Z(n66542) );
  NOR U86667 ( .A(n66543), .B(n66542), .Z(n71482) );
  IV U86668 ( .A(n66544), .Z(n66546) );
  NOR U86669 ( .A(n66546), .B(n66545), .Z(n71480) );
  NOR U86670 ( .A(n71482), .B(n71480), .Z(n68440) );
  IV U86671 ( .A(n66547), .Z(n66548) );
  NOR U86672 ( .A(n66549), .B(n66548), .Z(n73375) );
  IV U86673 ( .A(n66550), .Z(n66552) );
  IV U86674 ( .A(n66551), .Z(n66557) );
  NOR U86675 ( .A(n66552), .B(n66557), .Z(n66553) );
  IV U86676 ( .A(n66553), .Z(n73373) );
  NOR U86677 ( .A(n66555), .B(n66554), .Z(n71485) );
  IV U86678 ( .A(n66556), .Z(n66558) );
  NOR U86679 ( .A(n66558), .B(n66557), .Z(n73369) );
  NOR U86680 ( .A(n71485), .B(n73369), .Z(n68438) );
  IV U86681 ( .A(n66559), .Z(n66561) );
  NOR U86682 ( .A(n66561), .B(n66560), .Z(n66562) );
  IV U86683 ( .A(n66562), .Z(n68432) );
  IV U86684 ( .A(n66563), .Z(n66565) );
  IV U86685 ( .A(n66564), .Z(n68430) );
  NOR U86686 ( .A(n66565), .B(n68430), .Z(n71500) );
  IV U86687 ( .A(n66566), .Z(n66567) );
  NOR U86688 ( .A(n66567), .B(n66569), .Z(n71503) );
  IV U86689 ( .A(n66568), .Z(n66570) );
  NOR U86690 ( .A(n66570), .B(n66569), .Z(n73355) );
  NOR U86691 ( .A(n71503), .B(n73355), .Z(n68416) );
  IV U86692 ( .A(n66571), .Z(n66572) );
  NOR U86693 ( .A(n66572), .B(n66576), .Z(n71513) );
  IV U86694 ( .A(n66573), .Z(n66574) );
  NOR U86695 ( .A(n66574), .B(n66576), .Z(n73342) );
  IV U86696 ( .A(n66575), .Z(n66577) );
  NOR U86697 ( .A(n66577), .B(n66576), .Z(n71516) );
  IV U86698 ( .A(n66578), .Z(n66581) );
  NOR U86699 ( .A(n68398), .B(n66579), .Z(n66580) );
  IV U86700 ( .A(n66580), .Z(n66583) );
  NOR U86701 ( .A(n66581), .B(n66583), .Z(n73336) );
  IV U86702 ( .A(n66582), .Z(n66584) );
  NOR U86703 ( .A(n66584), .B(n66583), .Z(n73333) );
  IV U86704 ( .A(n66585), .Z(n66587) );
  IV U86705 ( .A(n66586), .Z(n66591) );
  NOR U86706 ( .A(n66587), .B(n66591), .Z(n66588) );
  IV U86707 ( .A(n66588), .Z(n73319) );
  IV U86708 ( .A(n66589), .Z(n66590) );
  NOR U86709 ( .A(n66591), .B(n66590), .Z(n73325) );
  NOR U86710 ( .A(n73313), .B(n73325), .Z(n68395) );
  IV U86711 ( .A(n66592), .Z(n66594) );
  NOR U86712 ( .A(n66594), .B(n66593), .Z(n66595) );
  IV U86713 ( .A(n66595), .Z(n73312) );
  IV U86714 ( .A(n66596), .Z(n66598) );
  NOR U86715 ( .A(n66598), .B(n66597), .Z(n68393) );
  IV U86716 ( .A(n68393), .Z(n68386) );
  IV U86717 ( .A(n66599), .Z(n66601) );
  NOR U86718 ( .A(n66601), .B(n66600), .Z(n76932) );
  IV U86719 ( .A(n66602), .Z(n66603) );
  NOR U86720 ( .A(n66603), .B(n68383), .Z(n76927) );
  NOR U86721 ( .A(n76932), .B(n76927), .Z(n71521) );
  IV U86722 ( .A(n71521), .Z(n68378) );
  IV U86723 ( .A(n66604), .Z(n66609) );
  IV U86724 ( .A(n66605), .Z(n66606) );
  NOR U86725 ( .A(n66609), .B(n66606), .Z(n71529) );
  IV U86726 ( .A(n66607), .Z(n66608) );
  NOR U86727 ( .A(n66609), .B(n66608), .Z(n71526) );
  IV U86728 ( .A(n66610), .Z(n66611) );
  NOR U86729 ( .A(n66611), .B(n66613), .Z(n71535) );
  IV U86730 ( .A(n66612), .Z(n66614) );
  NOR U86731 ( .A(n66614), .B(n66613), .Z(n71532) );
  IV U86732 ( .A(n66615), .Z(n66620) );
  IV U86733 ( .A(n66616), .Z(n66617) );
  NOR U86734 ( .A(n66620), .B(n66617), .Z(n71541) );
  IV U86735 ( .A(n66618), .Z(n66622) );
  NOR U86736 ( .A(n66620), .B(n66619), .Z(n66621) );
  IV U86737 ( .A(n66621), .Z(n66624) );
  NOR U86738 ( .A(n66622), .B(n66624), .Z(n71538) );
  IV U86739 ( .A(n66623), .Z(n66625) );
  NOR U86740 ( .A(n66625), .B(n66624), .Z(n73304) );
  IV U86741 ( .A(n66626), .Z(n66628) );
  NOR U86742 ( .A(n66628), .B(n66627), .Z(n73301) );
  NOR U86743 ( .A(n66630), .B(n66629), .Z(n66631) );
  XOR U86744 ( .A(n66632), .B(n66631), .Z(n66633) );
  NOR U86745 ( .A(n66633), .B(n66638), .Z(n66634) );
  IV U86746 ( .A(n66634), .Z(n66635) );
  NOR U86747 ( .A(n66636), .B(n66635), .Z(n73290) );
  IV U86748 ( .A(n66637), .Z(n66639) );
  NOR U86749 ( .A(n66639), .B(n66638), .Z(n71544) );
  IV U86750 ( .A(n66640), .Z(n66644) );
  IV U86751 ( .A(n66641), .Z(n68374) );
  NOR U86752 ( .A(n68374), .B(n66642), .Z(n66643) );
  IV U86753 ( .A(n66643), .Z(n68376) );
  NOR U86754 ( .A(n66644), .B(n68376), .Z(n66645) );
  IV U86755 ( .A(n66645), .Z(n73280) );
  IV U86756 ( .A(n66646), .Z(n66647) );
  NOR U86757 ( .A(n66648), .B(n66647), .Z(n78675) );
  IV U86758 ( .A(n66649), .Z(n66650) );
  NOR U86759 ( .A(n66650), .B(n68370), .Z(n76943) );
  NOR U86760 ( .A(n78675), .B(n76943), .Z(n73275) );
  IV U86761 ( .A(n73275), .Z(n68368) );
  IV U86762 ( .A(n66651), .Z(n66652) );
  NOR U86763 ( .A(n66652), .B(n66658), .Z(n66653) );
  IV U86764 ( .A(n66653), .Z(n73274) );
  IV U86765 ( .A(n66654), .Z(n66655) );
  NOR U86766 ( .A(n66656), .B(n66655), .Z(n73265) );
  IV U86767 ( .A(n66657), .Z(n66659) );
  NOR U86768 ( .A(n66659), .B(n66658), .Z(n71548) );
  NOR U86769 ( .A(n73265), .B(n71548), .Z(n68367) );
  IV U86770 ( .A(n66660), .Z(n66661) );
  IV U86771 ( .A(n68349), .Z(n66663) );
  NOR U86772 ( .A(n66661), .B(n66663), .Z(n73268) );
  IV U86773 ( .A(n66662), .Z(n68350) );
  NOR U86774 ( .A(n68350), .B(n66663), .Z(n68359) );
  IV U86775 ( .A(n68359), .Z(n68347) );
  IV U86776 ( .A(n66664), .Z(n66665) );
  NOR U86777 ( .A(n68355), .B(n66665), .Z(n71553) );
  IV U86778 ( .A(n66666), .Z(n66668) );
  IV U86779 ( .A(n66667), .Z(n68345) );
  NOR U86780 ( .A(n66668), .B(n68345), .Z(n71559) );
  IV U86781 ( .A(n66669), .Z(n66670) );
  NOR U86782 ( .A(n66673), .B(n66670), .Z(n71556) );
  IV U86783 ( .A(n66671), .Z(n66672) );
  NOR U86784 ( .A(n66673), .B(n66672), .Z(n71565) );
  IV U86785 ( .A(n66674), .Z(n66675) );
  NOR U86786 ( .A(n66675), .B(n68329), .Z(n66676) );
  IV U86787 ( .A(n66676), .Z(n71576) );
  IV U86788 ( .A(n66677), .Z(n66678) );
  NOR U86789 ( .A(n66679), .B(n66678), .Z(n66680) );
  IV U86790 ( .A(n66680), .Z(n68333) );
  IV U86791 ( .A(n66681), .Z(n68332) );
  IV U86792 ( .A(n66682), .Z(n66683) );
  NOR U86793 ( .A(n68332), .B(n66683), .Z(n71577) );
  IV U86794 ( .A(n66684), .Z(n66685) );
  NOR U86795 ( .A(n66685), .B(n66689), .Z(n66686) );
  IV U86796 ( .A(n66686), .Z(n71585) );
  IV U86797 ( .A(n66687), .Z(n66688) );
  NOR U86798 ( .A(n66689), .B(n66688), .Z(n71591) );
  IV U86799 ( .A(n66690), .Z(n66691) );
  NOR U86800 ( .A(n66692), .B(n66691), .Z(n71589) );
  NOR U86801 ( .A(n71591), .B(n71589), .Z(n68316) );
  IV U86802 ( .A(n66693), .Z(n66694) );
  NOR U86803 ( .A(n66694), .B(n66700), .Z(n66695) );
  IV U86804 ( .A(n66695), .Z(n71601) );
  IV U86805 ( .A(n66696), .Z(n66698) );
  NOR U86806 ( .A(n66698), .B(n66697), .Z(n73237) );
  IV U86807 ( .A(n66699), .Z(n66701) );
  NOR U86808 ( .A(n66701), .B(n66700), .Z(n73241) );
  NOR U86809 ( .A(n73237), .B(n73241), .Z(n68302) );
  NOR U86810 ( .A(n66702), .B(n73226), .Z(n73232) );
  IV U86811 ( .A(n66703), .Z(n66709) );
  IV U86812 ( .A(n66704), .Z(n66705) );
  NOR U86813 ( .A(n66709), .B(n66705), .Z(n73222) );
  XOR U86814 ( .A(n66707), .B(n66706), .Z(n66712) );
  NOR U86815 ( .A(n66709), .B(n66708), .Z(n66710) );
  IV U86816 ( .A(n66710), .Z(n66711) );
  NOR U86817 ( .A(n66712), .B(n66711), .Z(n71608) );
  IV U86818 ( .A(n66713), .Z(n66714) );
  NOR U86819 ( .A(n66714), .B(n66716), .Z(n71605) );
  IV U86820 ( .A(n66715), .Z(n66717) );
  NOR U86821 ( .A(n66717), .B(n66716), .Z(n73218) );
  IV U86822 ( .A(n66718), .Z(n66721) );
  IV U86823 ( .A(n66719), .Z(n66720) );
  NOR U86824 ( .A(n66721), .B(n66720), .Z(n73215) );
  IV U86825 ( .A(n66722), .Z(n66723) );
  NOR U86826 ( .A(n66723), .B(n68294), .Z(n73211) );
  IV U86827 ( .A(n66724), .Z(n66725) );
  NOR U86828 ( .A(n66725), .B(n68294), .Z(n73208) );
  IV U86829 ( .A(n66726), .Z(n66727) );
  NOR U86830 ( .A(n66728), .B(n66727), .Z(n66729) );
  IV U86831 ( .A(n66729), .Z(n71618) );
  IV U86832 ( .A(n66730), .Z(n66731) );
  NOR U86833 ( .A(n66731), .B(n66736), .Z(n73192) );
  IV U86834 ( .A(n66732), .Z(n66733) );
  NOR U86835 ( .A(n66734), .B(n66733), .Z(n71624) );
  IV U86836 ( .A(n66735), .Z(n66737) );
  NOR U86837 ( .A(n66737), .B(n66736), .Z(n73189) );
  NOR U86838 ( .A(n71624), .B(n73189), .Z(n66738) );
  IV U86839 ( .A(n66738), .Z(n68274) );
  IV U86840 ( .A(n66739), .Z(n66743) );
  IV U86841 ( .A(n66740), .Z(n68268) );
  NOR U86842 ( .A(n66741), .B(n68268), .Z(n66742) );
  IV U86843 ( .A(n66742), .Z(n68272) );
  NOR U86844 ( .A(n66743), .B(n68272), .Z(n71622) );
  IV U86845 ( .A(n66744), .Z(n66745) );
  NOR U86846 ( .A(n68266), .B(n66745), .Z(n73163) );
  IV U86847 ( .A(n66746), .Z(n66748) );
  IV U86848 ( .A(n66747), .Z(n68260) );
  NOR U86849 ( .A(n66748), .B(n68260), .Z(n71627) );
  NOR U86850 ( .A(n73163), .B(n71627), .Z(n68263) );
  IV U86851 ( .A(n66749), .Z(n66750) );
  NOR U86852 ( .A(n66751), .B(n66750), .Z(n71637) );
  NOR U86853 ( .A(n71637), .B(n71632), .Z(n68255) );
  IV U86854 ( .A(n66752), .Z(n66757) );
  IV U86855 ( .A(n66753), .Z(n66754) );
  NOR U86856 ( .A(n66757), .B(n66754), .Z(n73157) );
  IV U86857 ( .A(n66755), .Z(n66759) );
  NOR U86858 ( .A(n66757), .B(n66756), .Z(n66758) );
  IV U86859 ( .A(n66758), .Z(n68249) );
  NOR U86860 ( .A(n66759), .B(n68249), .Z(n73154) );
  IV U86861 ( .A(n66760), .Z(n66761) );
  NOR U86862 ( .A(n66762), .B(n66761), .Z(n66763) );
  IV U86863 ( .A(n66763), .Z(n68243) );
  IV U86864 ( .A(n66764), .Z(n66766) );
  NOR U86865 ( .A(n66766), .B(n66765), .Z(n73130) );
  IV U86866 ( .A(n66767), .Z(n66768) );
  NOR U86867 ( .A(n66769), .B(n66768), .Z(n71647) );
  IV U86868 ( .A(n66770), .Z(n66771) );
  NOR U86869 ( .A(n66771), .B(n68229), .Z(n71645) );
  NOR U86870 ( .A(n71647), .B(n71645), .Z(n68226) );
  IV U86871 ( .A(n66772), .Z(n66776) );
  IV U86872 ( .A(n66773), .Z(n68218) );
  NOR U86873 ( .A(n66774), .B(n68218), .Z(n66775) );
  IV U86874 ( .A(n66775), .Z(n66779) );
  NOR U86875 ( .A(n66776), .B(n66779), .Z(n66777) );
  IV U86876 ( .A(n66777), .Z(n71652) );
  IV U86877 ( .A(n66778), .Z(n66780) );
  NOR U86878 ( .A(n66780), .B(n66779), .Z(n68222) );
  IV U86879 ( .A(n66781), .Z(n66782) );
  NOR U86880 ( .A(n68215), .B(n66782), .Z(n73111) );
  IV U86881 ( .A(n66783), .Z(n66784) );
  NOR U86882 ( .A(n66787), .B(n66784), .Z(n73108) );
  IV U86883 ( .A(n66785), .Z(n66786) );
  NOR U86884 ( .A(n66787), .B(n66786), .Z(n71654) );
  IV U86885 ( .A(n66788), .Z(n66790) );
  IV U86886 ( .A(n66789), .Z(n66794) );
  NOR U86887 ( .A(n66790), .B(n66794), .Z(n71656) );
  NOR U86888 ( .A(n71654), .B(n71656), .Z(n68213) );
  NOR U86889 ( .A(n66791), .B(n71660), .Z(n66795) );
  IV U86890 ( .A(n66792), .Z(n66793) );
  NOR U86891 ( .A(n66794), .B(n66793), .Z(n73105) );
  NOR U86892 ( .A(n66795), .B(n73105), .Z(n68212) );
  IV U86893 ( .A(n66796), .Z(n66797) );
  NOR U86894 ( .A(n66798), .B(n66797), .Z(n77134) );
  IV U86895 ( .A(n66799), .Z(n66801) );
  NOR U86896 ( .A(n66801), .B(n66800), .Z(n78595) );
  NOR U86897 ( .A(n77134), .B(n78595), .Z(n71664) );
  IV U86898 ( .A(n66802), .Z(n66804) );
  NOR U86899 ( .A(n66804), .B(n66803), .Z(n73093) );
  NOR U86900 ( .A(n71667), .B(n71665), .Z(n66805) );
  NOR U86901 ( .A(n73093), .B(n66805), .Z(n68211) );
  IV U86902 ( .A(n66806), .Z(n66807) );
  NOR U86903 ( .A(n68205), .B(n66807), .Z(n73077) );
  IV U86904 ( .A(n66808), .Z(n66809) );
  NOR U86905 ( .A(n66810), .B(n66809), .Z(n78575) );
  IV U86906 ( .A(n66811), .Z(n66814) );
  NOR U86907 ( .A(n66812), .B(n68205), .Z(n66813) );
  IV U86908 ( .A(n66813), .Z(n68208) );
  NOR U86909 ( .A(n66814), .B(n68208), .Z(n78585) );
  NOR U86910 ( .A(n78575), .B(n78585), .Z(n71669) );
  IV U86911 ( .A(n66815), .Z(n68202) );
  IV U86912 ( .A(n66816), .Z(n66817) );
  NOR U86913 ( .A(n68202), .B(n66817), .Z(n71673) );
  NOR U86914 ( .A(n66819), .B(n66818), .Z(n71680) );
  IV U86915 ( .A(n66820), .Z(n66821) );
  NOR U86916 ( .A(n66822), .B(n66821), .Z(n71685) );
  NOR U86917 ( .A(n71680), .B(n71685), .Z(n68199) );
  IV U86918 ( .A(n66823), .Z(n66826) );
  NOR U86919 ( .A(n66824), .B(n78562), .Z(n66825) );
  IV U86920 ( .A(n66825), .Z(n66828) );
  NOR U86921 ( .A(n66826), .B(n66828), .Z(n71682) );
  IV U86922 ( .A(n66827), .Z(n66829) );
  NOR U86923 ( .A(n66829), .B(n66828), .Z(n71688) );
  IV U86924 ( .A(n66830), .Z(n66831) );
  NOR U86925 ( .A(n66831), .B(n66839), .Z(n78563) );
  IV U86926 ( .A(n66832), .Z(n66833) );
  NOR U86927 ( .A(n78562), .B(n66833), .Z(n66834) );
  NOR U86928 ( .A(n78563), .B(n66834), .Z(n73069) );
  IV U86929 ( .A(n66835), .Z(n66836) );
  NOR U86930 ( .A(n66837), .B(n66836), .Z(n73062) );
  IV U86931 ( .A(n66838), .Z(n66840) );
  NOR U86932 ( .A(n66840), .B(n66839), .Z(n78564) );
  NOR U86933 ( .A(n73062), .B(n78564), .Z(n68198) );
  IV U86934 ( .A(n66841), .Z(n68195) );
  IV U86935 ( .A(n66842), .Z(n66843) );
  NOR U86936 ( .A(n68195), .B(n66843), .Z(n73059) );
  IV U86937 ( .A(n66844), .Z(n66846) );
  NOR U86938 ( .A(n66846), .B(n66845), .Z(n71694) );
  IV U86939 ( .A(n66847), .Z(n66850) );
  NOR U86940 ( .A(n66848), .B(n66852), .Z(n66849) );
  IV U86941 ( .A(n66849), .Z(n68191) );
  NOR U86942 ( .A(n66850), .B(n68191), .Z(n73043) );
  IV U86943 ( .A(n66851), .Z(n66853) );
  NOR U86944 ( .A(n66853), .B(n66852), .Z(n73039) );
  IV U86945 ( .A(n66854), .Z(n66859) );
  IV U86946 ( .A(n66855), .Z(n66856) );
  NOR U86947 ( .A(n66859), .B(n66856), .Z(n73036) );
  IV U86948 ( .A(n66857), .Z(n66858) );
  NOR U86949 ( .A(n66859), .B(n66858), .Z(n71697) );
  IV U86950 ( .A(n66860), .Z(n66861) );
  NOR U86951 ( .A(n66862), .B(n66861), .Z(n77177) );
  IV U86952 ( .A(n66863), .Z(n66864) );
  NOR U86953 ( .A(n66864), .B(n68187), .Z(n77171) );
  NOR U86954 ( .A(n77177), .B(n77171), .Z(n71700) );
  IV U86955 ( .A(n66865), .Z(n66869) );
  NOR U86956 ( .A(n66867), .B(n66866), .Z(n66868) );
  IV U86957 ( .A(n66868), .Z(n66873) );
  NOR U86958 ( .A(n66869), .B(n66873), .Z(n73026) );
  IV U86959 ( .A(n66870), .Z(n66871) );
  NOR U86960 ( .A(n66871), .B(n66873), .Z(n71708) );
  NOR U86961 ( .A(n73026), .B(n71708), .Z(n68178) );
  IV U86962 ( .A(n66872), .Z(n66874) );
  NOR U86963 ( .A(n66874), .B(n66873), .Z(n73011) );
  IV U86964 ( .A(n66875), .Z(n66880) );
  IV U86965 ( .A(n66876), .Z(n66877) );
  NOR U86966 ( .A(n66880), .B(n66877), .Z(n73014) );
  IV U86967 ( .A(n66878), .Z(n66879) );
  NOR U86968 ( .A(n66880), .B(n66879), .Z(n71710) );
  IV U86969 ( .A(n66881), .Z(n66887) );
  IV U86970 ( .A(n66882), .Z(n66883) );
  NOR U86971 ( .A(n66887), .B(n66883), .Z(n66884) );
  IV U86972 ( .A(n66884), .Z(n71717) );
  IV U86973 ( .A(n66885), .Z(n66886) );
  NOR U86974 ( .A(n66887), .B(n66886), .Z(n73006) );
  IV U86975 ( .A(n66888), .Z(n66889) );
  NOR U86976 ( .A(n66889), .B(n68159), .Z(n73003) );
  NOR U86977 ( .A(n73006), .B(n73003), .Z(n68167) );
  IV U86978 ( .A(n66890), .Z(n66891) );
  NOR U86979 ( .A(n66892), .B(n66891), .Z(n66893) );
  IV U86980 ( .A(n66893), .Z(n68150) );
  IV U86981 ( .A(n66894), .Z(n66897) );
  IV U86982 ( .A(n66895), .Z(n66896) );
  NOR U86983 ( .A(n66897), .B(n66896), .Z(n71725) );
  IV U86984 ( .A(n66898), .Z(n66900) );
  NOR U86985 ( .A(n66900), .B(n66899), .Z(n72978) );
  IV U86986 ( .A(n66901), .Z(n66904) );
  IV U86987 ( .A(n66902), .Z(n66903) );
  NOR U86988 ( .A(n66904), .B(n66903), .Z(n72975) );
  IV U86989 ( .A(n68136), .Z(n66905) );
  NOR U86990 ( .A(n66908), .B(n66905), .Z(n71737) );
  IV U86991 ( .A(n66906), .Z(n66907) );
  NOR U86992 ( .A(n66908), .B(n66907), .Z(n71735) );
  NOR U86993 ( .A(n71737), .B(n71735), .Z(n68135) );
  IV U86994 ( .A(n66909), .Z(n66912) );
  IV U86995 ( .A(n66910), .Z(n66911) );
  NOR U86996 ( .A(n66912), .B(n66911), .Z(n66913) );
  IV U86997 ( .A(n66913), .Z(n72967) );
  IV U86998 ( .A(n66914), .Z(n66915) );
  NOR U86999 ( .A(n66916), .B(n66915), .Z(n72969) );
  NOR U87000 ( .A(n71740), .B(n72969), .Z(n68134) );
  IV U87001 ( .A(n66917), .Z(n66918) );
  NOR U87002 ( .A(n66919), .B(n66918), .Z(n68127) );
  NOR U87003 ( .A(n66920), .B(n72944), .Z(n68099) );
  IV U87004 ( .A(n66921), .Z(n66924) );
  NOR U87005 ( .A(n66922), .B(n66929), .Z(n66923) );
  IV U87006 ( .A(n66923), .Z(n68084) );
  NOR U87007 ( .A(n66924), .B(n68084), .Z(n72935) );
  IV U87008 ( .A(n66925), .Z(n66927) );
  NOR U87009 ( .A(n66927), .B(n66926), .Z(n71761) );
  IV U87010 ( .A(n66928), .Z(n66930) );
  NOR U87011 ( .A(n66930), .B(n66929), .Z(n72938) );
  NOR U87012 ( .A(n71761), .B(n72938), .Z(n68081) );
  IV U87013 ( .A(n66931), .Z(n66932) );
  NOR U87014 ( .A(n68080), .B(n66932), .Z(n71767) );
  IV U87015 ( .A(n66933), .Z(n66935) );
  IV U87016 ( .A(n66934), .Z(n68068) );
  NOR U87017 ( .A(n66935), .B(n68068), .Z(n68071) );
  IV U87018 ( .A(n66936), .Z(n66937) );
  NOR U87019 ( .A(n66937), .B(n68063), .Z(n66938) );
  IV U87020 ( .A(n66938), .Z(n72928) );
  IV U87021 ( .A(n66939), .Z(n66940) );
  NOR U87022 ( .A(n66941), .B(n66940), .Z(n71770) );
  IV U87023 ( .A(n66942), .Z(n66943) );
  NOR U87024 ( .A(n66944), .B(n66943), .Z(n72924) );
  NOR U87025 ( .A(n71770), .B(n72924), .Z(n68061) );
  IV U87026 ( .A(n66945), .Z(n66948) );
  IV U87027 ( .A(n66946), .Z(n66947) );
  NOR U87028 ( .A(n66948), .B(n66947), .Z(n72920) );
  IV U87029 ( .A(n66949), .Z(n66951) );
  XOR U87030 ( .A(n68045), .B(n68058), .Z(n66950) );
  NOR U87031 ( .A(n66951), .B(n66950), .Z(n72917) );
  NOR U87032 ( .A(n66953), .B(n66952), .Z(n66954) );
  IV U87033 ( .A(n66954), .Z(n71777) );
  NOR U87034 ( .A(n66955), .B(n71777), .Z(n66956) );
  NOR U87035 ( .A(n72910), .B(n66956), .Z(n68041) );
  IV U87036 ( .A(n66957), .Z(n66958) );
  NOR U87037 ( .A(n68023), .B(n66958), .Z(n66959) );
  IV U87038 ( .A(n66959), .Z(n71786) );
  IV U87039 ( .A(n66960), .Z(n68028) );
  IV U87040 ( .A(n66961), .Z(n66963) );
  NOR U87041 ( .A(n66963), .B(n66962), .Z(n71807) );
  IV U87042 ( .A(n66964), .Z(n66974) );
  NOR U87043 ( .A(n66966), .B(n66965), .Z(n66967) );
  IV U87044 ( .A(n66967), .Z(n66972) );
  NOR U87045 ( .A(n66969), .B(n66968), .Z(n66970) );
  IV U87046 ( .A(n66970), .Z(n66971) );
  NOR U87047 ( .A(n66972), .B(n66971), .Z(n66973) );
  IV U87048 ( .A(n66973), .Z(n68015) );
  NOR U87049 ( .A(n66974), .B(n68015), .Z(n71802) );
  NOR U87050 ( .A(n71807), .B(n71802), .Z(n68010) );
  IV U87051 ( .A(n66975), .Z(n66978) );
  NOR U87052 ( .A(n66976), .B(n68000), .Z(n66977) );
  IV U87053 ( .A(n66977), .Z(n68007) );
  NOR U87054 ( .A(n66978), .B(n68007), .Z(n72899) );
  NOR U87055 ( .A(n66980), .B(n66979), .Z(n72860) );
  IV U87056 ( .A(n66981), .Z(n66983) );
  NOR U87057 ( .A(n66983), .B(n66982), .Z(n77296) );
  NOR U87058 ( .A(n77296), .B(n77291), .Z(n72857) );
  IV U87059 ( .A(n66984), .Z(n66985) );
  NOR U87060 ( .A(n66986), .B(n66985), .Z(n71828) );
  IV U87061 ( .A(n66987), .Z(n66991) );
  IV U87062 ( .A(n66988), .Z(n66993) );
  NOR U87063 ( .A(n66989), .B(n66993), .Z(n66990) );
  IV U87064 ( .A(n66990), .Z(n66996) );
  NOR U87065 ( .A(n66991), .B(n66996), .Z(n72850) );
  NOR U87066 ( .A(n71828), .B(n72850), .Z(n67951) );
  IV U87067 ( .A(n66992), .Z(n66994) );
  NOR U87068 ( .A(n66994), .B(n66993), .Z(n71833) );
  IV U87069 ( .A(n66995), .Z(n66997) );
  NOR U87070 ( .A(n66997), .B(n66996), .Z(n71830) );
  NOR U87071 ( .A(n71833), .B(n71830), .Z(n67950) );
  IV U87072 ( .A(n66998), .Z(n66999) );
  NOR U87073 ( .A(n67933), .B(n66999), .Z(n72833) );
  IV U87074 ( .A(n67000), .Z(n67001) );
  NOR U87075 ( .A(n67929), .B(n67001), .Z(n72824) );
  NOR U87076 ( .A(n72833), .B(n72824), .Z(n67930) );
  IV U87077 ( .A(n67002), .Z(n67003) );
  NOR U87078 ( .A(n67003), .B(n67015), .Z(n78271) );
  IV U87079 ( .A(n67004), .Z(n67005) );
  NOR U87080 ( .A(n67006), .B(n67005), .Z(n78279) );
  NOR U87081 ( .A(n78271), .B(n78279), .Z(n84108) );
  IV U87082 ( .A(n67007), .Z(n67010) );
  XOR U87083 ( .A(n67008), .B(n67015), .Z(n67009) );
  NOR U87084 ( .A(n67010), .B(n67009), .Z(n72799) );
  NOR U87085 ( .A(n67012), .B(n67011), .Z(n67013) );
  IV U87086 ( .A(n67013), .Z(n67018) );
  NOR U87087 ( .A(n67015), .B(n67014), .Z(n67016) );
  IV U87088 ( .A(n67016), .Z(n67017) );
  NOR U87089 ( .A(n67018), .B(n67017), .Z(n67019) );
  IV U87090 ( .A(n67019), .Z(n72797) );
  IV U87091 ( .A(n67020), .Z(n67022) );
  NOR U87092 ( .A(n67022), .B(n67021), .Z(n71842) );
  IV U87093 ( .A(n67023), .Z(n67024) );
  NOR U87094 ( .A(n67025), .B(n67024), .Z(n71839) );
  NOR U87095 ( .A(n71842), .B(n71839), .Z(n67916) );
  IV U87096 ( .A(n67026), .Z(n67027) );
  NOR U87097 ( .A(n67027), .B(n67029), .Z(n71845) );
  IV U87098 ( .A(n67028), .Z(n67030) );
  NOR U87099 ( .A(n67030), .B(n67029), .Z(n71847) );
  NOR U87100 ( .A(n71845), .B(n71847), .Z(n67915) );
  IV U87101 ( .A(n67031), .Z(n67910) );
  IV U87102 ( .A(n67032), .Z(n67034) );
  NOR U87103 ( .A(n67034), .B(n67033), .Z(n78244) );
  IV U87104 ( .A(n67035), .Z(n67037) );
  NOR U87105 ( .A(n67037), .B(n67036), .Z(n78253) );
  NOR U87106 ( .A(n78244), .B(n78253), .Z(n72787) );
  NOR U87107 ( .A(n67038), .B(n71854), .Z(n67902) );
  IV U87108 ( .A(n67039), .Z(n67041) );
  NOR U87109 ( .A(n67041), .B(n67040), .Z(n72772) );
  IV U87110 ( .A(n67042), .Z(n67044) );
  NOR U87111 ( .A(n67044), .B(n67043), .Z(n72766) );
  NOR U87112 ( .A(n72772), .B(n72766), .Z(n67045) );
  IV U87113 ( .A(n67045), .Z(n67901) );
  IV U87114 ( .A(n67046), .Z(n67047) );
  NOR U87115 ( .A(n67048), .B(n67047), .Z(n72770) );
  IV U87116 ( .A(n67049), .Z(n67050) );
  NOR U87117 ( .A(n67050), .B(n67897), .Z(n67051) );
  IV U87118 ( .A(n67051), .Z(n71861) );
  IV U87119 ( .A(n67052), .Z(n67053) );
  NOR U87120 ( .A(n67054), .B(n67053), .Z(n72755) );
  IV U87121 ( .A(n67055), .Z(n67056) );
  NOR U87122 ( .A(n67057), .B(n67056), .Z(n71858) );
  NOR U87123 ( .A(n72755), .B(n71858), .Z(n67893) );
  IV U87124 ( .A(n67058), .Z(n67059) );
  NOR U87125 ( .A(n67881), .B(n67059), .Z(n72734) );
  NOR U87126 ( .A(n78221), .B(n67060), .Z(n71873) );
  IV U87127 ( .A(n67061), .Z(n67062) );
  NOR U87128 ( .A(n67867), .B(n67062), .Z(n72720) );
  IV U87129 ( .A(n67063), .Z(n67069) );
  IV U87130 ( .A(n67064), .Z(n67065) );
  NOR U87131 ( .A(n67069), .B(n67065), .Z(n67066) );
  IV U87132 ( .A(n67066), .Z(n71894) );
  IV U87133 ( .A(n67068), .Z(n67067) );
  NOR U87134 ( .A(n67069), .B(n67067), .Z(n72704) );
  XOR U87135 ( .A(n67069), .B(n67068), .Z(n67072) );
  IV U87136 ( .A(n67070), .Z(n67071) );
  NOR U87137 ( .A(n67072), .B(n67071), .Z(n71896) );
  NOR U87138 ( .A(n72704), .B(n71896), .Z(n67838) );
  IV U87139 ( .A(n67073), .Z(n67075) );
  NOR U87140 ( .A(n67075), .B(n67074), .Z(n72695) );
  IV U87141 ( .A(n67076), .Z(n67077) );
  NOR U87142 ( .A(n67828), .B(n67077), .Z(n71898) );
  IV U87143 ( .A(n67078), .Z(n67083) );
  IV U87144 ( .A(n67079), .Z(n67080) );
  NOR U87145 ( .A(n67828), .B(n67080), .Z(n67081) );
  IV U87146 ( .A(n67081), .Z(n67082) );
  NOR U87147 ( .A(n67083), .B(n67082), .Z(n72692) );
  IV U87148 ( .A(n67084), .Z(n67085) );
  NOR U87149 ( .A(n67085), .B(n67813), .Z(n67086) );
  IV U87150 ( .A(n67086), .Z(n71908) );
  IV U87151 ( .A(n67087), .Z(n67089) );
  NOR U87152 ( .A(n67089), .B(n67088), .Z(n72671) );
  IV U87153 ( .A(n67090), .Z(n67092) );
  NOR U87154 ( .A(n67092), .B(n67091), .Z(n72679) );
  NOR U87155 ( .A(n72671), .B(n72679), .Z(n67807) );
  IV U87156 ( .A(n67093), .Z(n67094) );
  NOR U87157 ( .A(n67094), .B(n67097), .Z(n71916) );
  IV U87158 ( .A(n67095), .Z(n67096) );
  NOR U87159 ( .A(n67097), .B(n67096), .Z(n71921) );
  IV U87160 ( .A(n67098), .Z(n67099) );
  NOR U87161 ( .A(n67100), .B(n67099), .Z(n71919) );
  NOR U87162 ( .A(n72663), .B(n71919), .Z(n67799) );
  IV U87163 ( .A(n67101), .Z(n67102) );
  NOR U87164 ( .A(n67102), .B(n67104), .Z(n72660) );
  IV U87165 ( .A(n67103), .Z(n67105) );
  NOR U87166 ( .A(n67105), .B(n67104), .Z(n67106) );
  IV U87167 ( .A(n67106), .Z(n71925) );
  IV U87168 ( .A(n67107), .Z(n67109) );
  NOR U87169 ( .A(n67109), .B(n67108), .Z(n72653) );
  IV U87170 ( .A(n67110), .Z(n67111) );
  NOR U87171 ( .A(n67112), .B(n67111), .Z(n67113) );
  IV U87172 ( .A(n67113), .Z(n67789) );
  IV U87173 ( .A(n67114), .Z(n67115) );
  NOR U87174 ( .A(n67115), .B(n67120), .Z(n72643) );
  IV U87175 ( .A(n67116), .Z(n67117) );
  NOR U87176 ( .A(n67118), .B(n67117), .Z(n83212) );
  IV U87177 ( .A(n67119), .Z(n67121) );
  NOR U87178 ( .A(n67121), .B(n67120), .Z(n83207) );
  NOR U87179 ( .A(n83212), .B(n83207), .Z(n78129) );
  IV U87180 ( .A(n67122), .Z(n67123) );
  NOR U87181 ( .A(n67126), .B(n67123), .Z(n71942) );
  IV U87182 ( .A(n67124), .Z(n67125) );
  NOR U87183 ( .A(n67126), .B(n67125), .Z(n71947) );
  IV U87184 ( .A(n67127), .Z(n67131) );
  NOR U87185 ( .A(n67129), .B(n67128), .Z(n67130) );
  IV U87186 ( .A(n67130), .Z(n67133) );
  NOR U87187 ( .A(n67131), .B(n67133), .Z(n72630) );
  IV U87188 ( .A(n67132), .Z(n67134) );
  NOR U87189 ( .A(n67134), .B(n67133), .Z(n71950) );
  XOR U87190 ( .A(n72630), .B(n71950), .Z(n67135) );
  NOR U87191 ( .A(n71947), .B(n67135), .Z(n67752) );
  IV U87192 ( .A(n67136), .Z(n67139) );
  NOR U87193 ( .A(n67137), .B(n67144), .Z(n67138) );
  IV U87194 ( .A(n67138), .Z(n67141) );
  NOR U87195 ( .A(n67139), .B(n67141), .Z(n71953) );
  IV U87196 ( .A(n67140), .Z(n67142) );
  NOR U87197 ( .A(n67142), .B(n67141), .Z(n72623) );
  IV U87198 ( .A(n67143), .Z(n67145) );
  NOR U87199 ( .A(n67145), .B(n67144), .Z(n72620) );
  IV U87200 ( .A(n67146), .Z(n67147) );
  NOR U87201 ( .A(n67147), .B(n67750), .Z(n71956) );
  IV U87202 ( .A(n67148), .Z(n67150) );
  NOR U87203 ( .A(n67150), .B(n67149), .Z(n67151) );
  IV U87204 ( .A(n67151), .Z(n71963) );
  IV U87205 ( .A(n67152), .Z(n67153) );
  NOR U87206 ( .A(n67153), .B(n67739), .Z(n72612) );
  IV U87207 ( .A(n67154), .Z(n67155) );
  NOR U87208 ( .A(n67155), .B(n67729), .Z(n71967) );
  IV U87209 ( .A(n67156), .Z(n67157) );
  NOR U87210 ( .A(n67158), .B(n67157), .Z(n72588) );
  NOR U87211 ( .A(n71970), .B(n72588), .Z(n72576) );
  IV U87212 ( .A(n72576), .Z(n67727) );
  IV U87213 ( .A(n67159), .Z(n67160) );
  NOR U87214 ( .A(n67160), .B(n67723), .Z(n72577) );
  IV U87215 ( .A(n67161), .Z(n67162) );
  NOR U87216 ( .A(n67163), .B(n67162), .Z(n78068) );
  IV U87217 ( .A(n67164), .Z(n67166) );
  IV U87218 ( .A(n67165), .Z(n67710) );
  NOR U87219 ( .A(n67166), .B(n67710), .Z(n78059) );
  NOR U87220 ( .A(n78068), .B(n78059), .Z(n71979) );
  IV U87221 ( .A(n67167), .Z(n67169) );
  NOR U87222 ( .A(n67169), .B(n67168), .Z(n72003) );
  IV U87223 ( .A(n67170), .Z(n67171) );
  NOR U87224 ( .A(n67171), .B(n67173), .Z(n72018) );
  IV U87225 ( .A(n67172), .Z(n67174) );
  NOR U87226 ( .A(n67174), .B(n67173), .Z(n72015) );
  IV U87227 ( .A(n67175), .Z(n67176) );
  NOR U87228 ( .A(n67177), .B(n67176), .Z(n72536) );
  IV U87229 ( .A(n67178), .Z(n67179) );
  NOR U87230 ( .A(n67180), .B(n67179), .Z(n72021) );
  NOR U87231 ( .A(n72536), .B(n72021), .Z(n67181) );
  IV U87232 ( .A(n67181), .Z(n67670) );
  IV U87233 ( .A(n67182), .Z(n67183) );
  NOR U87234 ( .A(n67183), .B(n67185), .Z(n72533) );
  IV U87235 ( .A(n67184), .Z(n67186) );
  NOR U87236 ( .A(n67186), .B(n67185), .Z(n72026) );
  IV U87237 ( .A(n67187), .Z(n67192) );
  IV U87238 ( .A(n67188), .Z(n67190) );
  NOR U87239 ( .A(n67190), .B(n67189), .Z(n67191) );
  IV U87240 ( .A(n67191), .Z(n67668) );
  NOR U87241 ( .A(n67192), .B(n67668), .Z(n67193) );
  IV U87242 ( .A(n67193), .Z(n72024) );
  NOR U87243 ( .A(n67194), .B(n67644), .Z(n67642) );
  IV U87244 ( .A(n67195), .Z(n67197) );
  NOR U87245 ( .A(n67197), .B(n67196), .Z(n72520) );
  IV U87246 ( .A(n67198), .Z(n67200) );
  NOR U87247 ( .A(n67200), .B(n67199), .Z(n72510) );
  IV U87248 ( .A(n67201), .Z(n67203) );
  NOR U87249 ( .A(n67203), .B(n67202), .Z(n72041) );
  NOR U87250 ( .A(n72510), .B(n72041), .Z(n67637) );
  IV U87251 ( .A(n67204), .Z(n67205) );
  NOR U87252 ( .A(n67206), .B(n67205), .Z(n72513) );
  IV U87253 ( .A(n67207), .Z(n67209) );
  IV U87254 ( .A(n67208), .Z(n67214) );
  NOR U87255 ( .A(n67209), .B(n67214), .Z(n72043) );
  NOR U87256 ( .A(n72513), .B(n72043), .Z(n67210) );
  IV U87257 ( .A(n67210), .Z(n67636) );
  IV U87258 ( .A(n67211), .Z(n67212) );
  NOR U87259 ( .A(n67212), .B(n67631), .Z(n72501) );
  IV U87260 ( .A(n67213), .Z(n67215) );
  NOR U87261 ( .A(n67215), .B(n67214), .Z(n72506) );
  NOR U87262 ( .A(n72501), .B(n72506), .Z(n67635) );
  IV U87263 ( .A(n67216), .Z(n67217) );
  NOR U87264 ( .A(n67217), .B(n67634), .Z(n72045) );
  IV U87265 ( .A(n67218), .Z(n67219) );
  NOR U87266 ( .A(n67225), .B(n67219), .Z(n67220) );
  IV U87267 ( .A(n67220), .Z(n72485) );
  IV U87268 ( .A(n67221), .Z(n67222) );
  NOR U87269 ( .A(n67223), .B(n67222), .Z(n77930) );
  IV U87270 ( .A(n67224), .Z(n67226) );
  NOR U87271 ( .A(n67226), .B(n67225), .Z(n77953) );
  NOR U87272 ( .A(n77930), .B(n77953), .Z(n72056) );
  IV U87273 ( .A(n67227), .Z(n67229) );
  NOR U87274 ( .A(n67229), .B(n67228), .Z(n72060) );
  IV U87275 ( .A(n67230), .Z(n67231) );
  NOR U87276 ( .A(n67231), .B(n67614), .Z(n72057) );
  IV U87277 ( .A(n67232), .Z(n67234) );
  IV U87278 ( .A(n67233), .Z(n67237) );
  NOR U87279 ( .A(n67234), .B(n67237), .Z(n72475) );
  NOR U87280 ( .A(n67235), .B(n72463), .Z(n67239) );
  IV U87281 ( .A(n67236), .Z(n67238) );
  NOR U87282 ( .A(n67238), .B(n67237), .Z(n72468) );
  NOR U87283 ( .A(n67239), .B(n72468), .Z(n67609) );
  IV U87284 ( .A(n67240), .Z(n67241) );
  NOR U87285 ( .A(n67243), .B(n67241), .Z(n72069) );
  IV U87286 ( .A(n67242), .Z(n67244) );
  NOR U87287 ( .A(n67244), .B(n67243), .Z(n72435) );
  IV U87288 ( .A(n67245), .Z(n67246) );
  NOR U87289 ( .A(n67246), .B(n67257), .Z(n72432) );
  IV U87290 ( .A(n67247), .Z(n67249) );
  NOR U87291 ( .A(n67249), .B(n67248), .Z(n72438) );
  NOR U87292 ( .A(n72432), .B(n72438), .Z(n67577) );
  IV U87293 ( .A(n67250), .Z(n67251) );
  NOR U87294 ( .A(n67251), .B(n67257), .Z(n72428) );
  NOR U87295 ( .A(n67253), .B(n67252), .Z(n67254) );
  IV U87296 ( .A(n67254), .Z(n67255) );
  NOR U87297 ( .A(n67255), .B(n67257), .Z(n72425) );
  IV U87298 ( .A(n67256), .Z(n67261) );
  NOR U87299 ( .A(n67258), .B(n67257), .Z(n67259) );
  IV U87300 ( .A(n67259), .Z(n67260) );
  NOR U87301 ( .A(n67261), .B(n67260), .Z(n72420) );
  IV U87302 ( .A(n67262), .Z(n67267) );
  IV U87303 ( .A(n67263), .Z(n67264) );
  NOR U87304 ( .A(n67267), .B(n67264), .Z(n77563) );
  IV U87305 ( .A(n67265), .Z(n67269) );
  NOR U87306 ( .A(n67267), .B(n67266), .Z(n67268) );
  IV U87307 ( .A(n67268), .Z(n67271) );
  NOR U87308 ( .A(n67269), .B(n67271), .Z(n77568) );
  NOR U87309 ( .A(n77563), .B(n77568), .Z(n72419) );
  IV U87310 ( .A(n67270), .Z(n67272) );
  NOR U87311 ( .A(n67272), .B(n67271), .Z(n72408) );
  IV U87312 ( .A(n67273), .Z(n67274) );
  NOR U87313 ( .A(n67275), .B(n67274), .Z(n72078) );
  IV U87314 ( .A(n67276), .Z(n67277) );
  NOR U87315 ( .A(n67277), .B(n67574), .Z(n72411) );
  NOR U87316 ( .A(n72078), .B(n72411), .Z(n67278) );
  IV U87317 ( .A(n67278), .Z(n67572) );
  IV U87318 ( .A(n67279), .Z(n67280) );
  NOR U87319 ( .A(n67280), .B(n67569), .Z(n67281) );
  IV U87320 ( .A(n67281), .Z(n72403) );
  NOR U87321 ( .A(n67282), .B(n72391), .Z(n67564) );
  IV U87322 ( .A(n67283), .Z(n67284) );
  NOR U87323 ( .A(n67285), .B(n67284), .Z(n72387) );
  NOR U87324 ( .A(n72384), .B(n72387), .Z(n67562) );
  IV U87325 ( .A(n67286), .Z(n67290) );
  NOR U87326 ( .A(n67288), .B(n67287), .Z(n67289) );
  IV U87327 ( .A(n67289), .Z(n67292) );
  NOR U87328 ( .A(n67290), .B(n67292), .Z(n72381) );
  IV U87329 ( .A(n67291), .Z(n67293) );
  NOR U87330 ( .A(n67293), .B(n67292), .Z(n72377) );
  IV U87331 ( .A(n67294), .Z(n67299) );
  IV U87332 ( .A(n67295), .Z(n67296) );
  NOR U87333 ( .A(n67299), .B(n67296), .Z(n72374) );
  IV U87334 ( .A(n67297), .Z(n67298) );
  NOR U87335 ( .A(n67299), .B(n67298), .Z(n72361) );
  IV U87336 ( .A(n67300), .Z(n67302) );
  NOR U87337 ( .A(n67302), .B(n67301), .Z(n72358) );
  IV U87338 ( .A(n67303), .Z(n67305) );
  NOR U87339 ( .A(n67305), .B(n67304), .Z(n72080) );
  NOR U87340 ( .A(n67307), .B(n67306), .Z(n67308) );
  IV U87341 ( .A(n67308), .Z(n67315) );
  XOR U87342 ( .A(n67310), .B(n67309), .Z(n67311) );
  NOR U87343 ( .A(n67312), .B(n67311), .Z(n67313) );
  IV U87344 ( .A(n67313), .Z(n67314) );
  NOR U87345 ( .A(n67315), .B(n67314), .Z(n72086) );
  IV U87346 ( .A(n67316), .Z(n67317) );
  NOR U87347 ( .A(n67320), .B(n67317), .Z(n72349) );
  IV U87348 ( .A(n67318), .Z(n67322) );
  NOR U87349 ( .A(n67320), .B(n67319), .Z(n67321) );
  IV U87350 ( .A(n67321), .Z(n67324) );
  NOR U87351 ( .A(n67322), .B(n67324), .Z(n72346) );
  IV U87352 ( .A(n67323), .Z(n67325) );
  NOR U87353 ( .A(n67325), .B(n67324), .Z(n72341) );
  IV U87354 ( .A(n67326), .Z(n67330) );
  IV U87355 ( .A(n67327), .Z(n67328) );
  NOR U87356 ( .A(n67330), .B(n67328), .Z(n72094) );
  IV U87357 ( .A(n67329), .Z(n67331) );
  NOR U87358 ( .A(n67331), .B(n67330), .Z(n72100) );
  NOR U87359 ( .A(n72103), .B(n72100), .Z(n67551) );
  IV U87360 ( .A(n67332), .Z(n67334) );
  NOR U87361 ( .A(n67334), .B(n67333), .Z(n72320) );
  IV U87362 ( .A(n67335), .Z(n67338) );
  IV U87363 ( .A(n67336), .Z(n67337) );
  NOR U87364 ( .A(n67338), .B(n67337), .Z(n72317) );
  IV U87365 ( .A(n67339), .Z(n67341) );
  NOR U87366 ( .A(n67341), .B(n67340), .Z(n72106) );
  NOR U87367 ( .A(n72108), .B(n72106), .Z(n67545) );
  NOR U87368 ( .A(n67343), .B(n67342), .Z(n67344) );
  IV U87369 ( .A(n67344), .Z(n67345) );
  NOR U87370 ( .A(n67346), .B(n67345), .Z(n72310) );
  IV U87371 ( .A(n67347), .Z(n67348) );
  NOR U87372 ( .A(n67349), .B(n67348), .Z(n72111) );
  IV U87373 ( .A(n67350), .Z(n67351) );
  NOR U87374 ( .A(n67354), .B(n67351), .Z(n72293) );
  NOR U87375 ( .A(n72111), .B(n72293), .Z(n67537) );
  IV U87376 ( .A(n67352), .Z(n67356) );
  NOR U87377 ( .A(n67354), .B(n67353), .Z(n67355) );
  IV U87378 ( .A(n67355), .Z(n67358) );
  NOR U87379 ( .A(n67356), .B(n67358), .Z(n72290) );
  IV U87380 ( .A(n67357), .Z(n67359) );
  NOR U87381 ( .A(n67359), .B(n67358), .Z(n72286) );
  IV U87382 ( .A(n67360), .Z(n67361) );
  NOR U87383 ( .A(n67361), .B(n72115), .Z(n72283) );
  NOR U87384 ( .A(n67362), .B(n72115), .Z(n67536) );
  IV U87385 ( .A(n67363), .Z(n67364) );
  NOR U87386 ( .A(n67366), .B(n67364), .Z(n77812) );
  IV U87387 ( .A(n67365), .Z(n67367) );
  NOR U87388 ( .A(n67367), .B(n67366), .Z(n77655) );
  NOR U87389 ( .A(n77812), .B(n77655), .Z(n72276) );
  IV U87390 ( .A(n67368), .Z(n67373) );
  IV U87391 ( .A(n67369), .Z(n67370) );
  NOR U87392 ( .A(n67373), .B(n67370), .Z(n72118) );
  IV U87393 ( .A(n67371), .Z(n67372) );
  NOR U87394 ( .A(n67373), .B(n67372), .Z(n72120) );
  NOR U87395 ( .A(n72118), .B(n72120), .Z(n67535) );
  NOR U87396 ( .A(n67375), .B(n67374), .Z(n77772) );
  IV U87397 ( .A(n67376), .Z(n67524) );
  IV U87398 ( .A(n67377), .Z(n67378) );
  NOR U87399 ( .A(n67524), .B(n67378), .Z(n77786) );
  NOR U87400 ( .A(n77772), .B(n77786), .Z(n72135) );
  IV U87401 ( .A(n67379), .Z(n67517) );
  IV U87402 ( .A(n67380), .Z(n67381) );
  NOR U87403 ( .A(n67517), .B(n67381), .Z(n72138) );
  IV U87404 ( .A(n67382), .Z(n67383) );
  NOR U87405 ( .A(n67384), .B(n67383), .Z(n72268) );
  IV U87406 ( .A(n67385), .Z(n67512) );
  IV U87407 ( .A(n67511), .Z(n67387) );
  NOR U87408 ( .A(n67512), .B(n67387), .Z(n72146) );
  IV U87409 ( .A(n67386), .Z(n67388) );
  NOR U87410 ( .A(n67388), .B(n67387), .Z(n72144) );
  NOR U87411 ( .A(n72146), .B(n72144), .Z(n67509) );
  IV U87412 ( .A(n67389), .Z(n67390) );
  NOR U87413 ( .A(n67390), .B(n67393), .Z(n67391) );
  IV U87414 ( .A(n67391), .Z(n72152) );
  IV U87415 ( .A(n67392), .Z(n67394) );
  NOR U87416 ( .A(n67394), .B(n67393), .Z(n72148) );
  IV U87417 ( .A(n67395), .Z(n67400) );
  IV U87418 ( .A(n67396), .Z(n67397) );
  NOR U87419 ( .A(n67400), .B(n67397), .Z(n72153) );
  IV U87420 ( .A(n67398), .Z(n67399) );
  NOR U87421 ( .A(n67400), .B(n67399), .Z(n72259) );
  NOR U87422 ( .A(n72153), .B(n72259), .Z(n67401) );
  IV U87423 ( .A(n67401), .Z(n67405) );
  IV U87424 ( .A(n67402), .Z(n67404) );
  NOR U87425 ( .A(n67404), .B(n67403), .Z(n72155) );
  NOR U87426 ( .A(n67405), .B(n72155), .Z(n67506) );
  IV U87427 ( .A(n67406), .Z(n67408) );
  IV U87428 ( .A(n67407), .Z(n67413) );
  NOR U87429 ( .A(n67408), .B(n67413), .Z(n72248) );
  IV U87430 ( .A(n67409), .Z(n67411) );
  NOR U87431 ( .A(n67411), .B(n67410), .Z(n72157) );
  NOR U87432 ( .A(n72248), .B(n72157), .Z(n67496) );
  IV U87433 ( .A(n67412), .Z(n67414) );
  NOR U87434 ( .A(n67414), .B(n67413), .Z(n72245) );
  IV U87435 ( .A(n67415), .Z(n67419) );
  IV U87436 ( .A(n67416), .Z(n67423) );
  XOR U87437 ( .A(n67417), .B(n67423), .Z(n67418) );
  NOR U87438 ( .A(n67419), .B(n67418), .Z(n72164) );
  IV U87439 ( .A(n67420), .Z(n67421) );
  NOR U87440 ( .A(n67421), .B(n67423), .Z(n72240) );
  IV U87441 ( .A(n67422), .Z(n67426) );
  NOR U87442 ( .A(n67424), .B(n67423), .Z(n67425) );
  IV U87443 ( .A(n67425), .Z(n67429) );
  NOR U87444 ( .A(n67426), .B(n67429), .Z(n72237) );
  NOR U87445 ( .A(n67427), .B(n72228), .Z(n67431) );
  IV U87446 ( .A(n67428), .Z(n67430) );
  NOR U87447 ( .A(n67430), .B(n67429), .Z(n72234) );
  NOR U87448 ( .A(n67431), .B(n72234), .Z(n67486) );
  IV U87449 ( .A(n67432), .Z(n67434) );
  IV U87450 ( .A(n67433), .Z(n72207) );
  NOR U87451 ( .A(n67434), .B(n72207), .Z(n67435) );
  IV U87452 ( .A(n67435), .Z(n67436) );
  NOR U87453 ( .A(n67437), .B(n67436), .Z(n72172) );
  IV U87454 ( .A(n67438), .Z(n67439) );
  NOR U87455 ( .A(n67440), .B(n67439), .Z(n67441) );
  IV U87456 ( .A(n67441), .Z(n72206) );
  NOR U87457 ( .A(n67442), .B(n72206), .Z(n72211) );
  NOR U87458 ( .A(n67443), .B(n67442), .Z(n67444) );
  IV U87459 ( .A(n67444), .Z(n72214) );
  IV U87460 ( .A(n67445), .Z(n67447) );
  NOR U87461 ( .A(n67447), .B(n67446), .Z(n72217) );
  IV U87462 ( .A(n67448), .Z(n67450) );
  NOR U87463 ( .A(n67450), .B(n67449), .Z(n72219) );
  NOR U87464 ( .A(n72217), .B(n72219), .Z(n67479) );
  IV U87465 ( .A(n67451), .Z(n67452) );
  NOR U87466 ( .A(n67453), .B(n67452), .Z(n72191) );
  IV U87467 ( .A(n67454), .Z(n67457) );
  IV U87468 ( .A(n67455), .Z(n67456) );
  NOR U87469 ( .A(n67457), .B(n67456), .Z(n72178) );
  IV U87470 ( .A(n67458), .Z(n67459) );
  NOR U87471 ( .A(n67459), .B(n67468), .Z(n72179) );
  XOR U87472 ( .A(n72178), .B(n72179), .Z(n67465) );
  NOR U87473 ( .A(n67461), .B(n67460), .Z(n67462) );
  IV U87474 ( .A(n67462), .Z(n67463) );
  NOR U87475 ( .A(n72179), .B(n67463), .Z(n67464) );
  NOR U87476 ( .A(n67465), .B(n67464), .Z(n72184) );
  IV U87477 ( .A(n67466), .Z(n67467) );
  NOR U87478 ( .A(n67468), .B(n67467), .Z(n72182) );
  XOR U87479 ( .A(n72184), .B(n72182), .Z(n72189) );
  XOR U87480 ( .A(n72191), .B(n72189), .Z(n72201) );
  IV U87481 ( .A(n72201), .Z(n67475) );
  IV U87482 ( .A(n67469), .Z(n67470) );
  NOR U87483 ( .A(n67471), .B(n67470), .Z(n72188) );
  IV U87484 ( .A(n67472), .Z(n67473) );
  NOR U87485 ( .A(n67473), .B(n67478), .Z(n72199) );
  NOR U87486 ( .A(n72188), .B(n72199), .Z(n67474) );
  XOR U87487 ( .A(n67475), .B(n67474), .Z(n72198) );
  IV U87488 ( .A(n67476), .Z(n67477) );
  NOR U87489 ( .A(n67478), .B(n67477), .Z(n72196) );
  XOR U87490 ( .A(n72198), .B(n72196), .Z(n72220) );
  XOR U87491 ( .A(n67479), .B(n72220), .Z(n72204) );
  XOR U87492 ( .A(n72214), .B(n72204), .Z(n72212) );
  XOR U87493 ( .A(n72211), .B(n72212), .Z(n72173) );
  XOR U87494 ( .A(n72172), .B(n72173), .Z(n72177) );
  IV U87495 ( .A(n67480), .Z(n67481) );
  NOR U87496 ( .A(n67482), .B(n67481), .Z(n72170) );
  IV U87497 ( .A(n67483), .Z(n67484) );
  NOR U87498 ( .A(n72207), .B(n67484), .Z(n72175) );
  NOR U87499 ( .A(n72170), .B(n72175), .Z(n67485) );
  XOR U87500 ( .A(n72177), .B(n67485), .Z(n72227) );
  XOR U87501 ( .A(n67486), .B(n72227), .Z(n72239) );
  XOR U87502 ( .A(n72237), .B(n72239), .Z(n72241) );
  XOR U87503 ( .A(n72240), .B(n72241), .Z(n72165) );
  XOR U87504 ( .A(n72164), .B(n72165), .Z(n72169) );
  IV U87505 ( .A(n72169), .Z(n67495) );
  IV U87506 ( .A(n67487), .Z(n67490) );
  IV U87507 ( .A(n67488), .Z(n67489) );
  NOR U87508 ( .A(n67490), .B(n67489), .Z(n72162) );
  IV U87509 ( .A(n67491), .Z(n67493) );
  NOR U87510 ( .A(n67493), .B(n67492), .Z(n72167) );
  NOR U87511 ( .A(n72162), .B(n72167), .Z(n67494) );
  XOR U87512 ( .A(n67495), .B(n67494), .Z(n72247) );
  XOR U87513 ( .A(n72245), .B(n72247), .Z(n72249) );
  XOR U87514 ( .A(n67496), .B(n72249), .Z(n72160) );
  IV U87515 ( .A(n67497), .Z(n67498) );
  NOR U87516 ( .A(n67498), .B(n67500), .Z(n72159) );
  IV U87517 ( .A(n67499), .Z(n67501) );
  NOR U87518 ( .A(n67501), .B(n67500), .Z(n72255) );
  NOR U87519 ( .A(n72159), .B(n72255), .Z(n67502) );
  XOR U87520 ( .A(n72160), .B(n67502), .Z(n83558) );
  IV U87521 ( .A(n67503), .Z(n67505) );
  NOR U87522 ( .A(n67505), .B(n67504), .Z(n72253) );
  XOR U87523 ( .A(n83558), .B(n72253), .Z(n72260) );
  XOR U87524 ( .A(n67506), .B(n72260), .Z(n67507) );
  IV U87525 ( .A(n67507), .Z(n72150) );
  XOR U87526 ( .A(n72148), .B(n72150), .Z(n72151) );
  XOR U87527 ( .A(n72152), .B(n72151), .Z(n67508) );
  XOR U87528 ( .A(n67509), .B(n67508), .Z(n72267) );
  IV U87529 ( .A(n67510), .Z(n67514) );
  XOR U87530 ( .A(n67512), .B(n67511), .Z(n67513) );
  NOR U87531 ( .A(n67514), .B(n67513), .Z(n72265) );
  XOR U87532 ( .A(n72267), .B(n72265), .Z(n72269) );
  XOR U87533 ( .A(n72268), .B(n72269), .Z(n72139) );
  XOR U87534 ( .A(n72138), .B(n72139), .Z(n72142) );
  IV U87535 ( .A(n67515), .Z(n67516) );
  NOR U87536 ( .A(n67517), .B(n67516), .Z(n72141) );
  IV U87537 ( .A(n67518), .Z(n67519) );
  NOR U87538 ( .A(n67520), .B(n67519), .Z(n72136) );
  NOR U87539 ( .A(n72141), .B(n72136), .Z(n67521) );
  XOR U87540 ( .A(n72142), .B(n67521), .Z(n72134) );
  XOR U87541 ( .A(n72135), .B(n72134), .Z(n72130) );
  IV U87542 ( .A(n67522), .Z(n67523) );
  NOR U87543 ( .A(n67524), .B(n67523), .Z(n72128) );
  XOR U87544 ( .A(n72130), .B(n72128), .Z(n72132) );
  IV U87545 ( .A(n67525), .Z(n67526) );
  NOR U87546 ( .A(n67527), .B(n67526), .Z(n72131) );
  IV U87547 ( .A(n67528), .Z(n67529) );
  NOR U87548 ( .A(n67534), .B(n67529), .Z(n72126) );
  NOR U87549 ( .A(n72131), .B(n72126), .Z(n67530) );
  XOR U87550 ( .A(n72132), .B(n67530), .Z(n67531) );
  IV U87551 ( .A(n67531), .Z(n72125) );
  IV U87552 ( .A(n67532), .Z(n67533) );
  NOR U87553 ( .A(n67534), .B(n67533), .Z(n72123) );
  XOR U87554 ( .A(n72125), .B(n72123), .Z(n72121) );
  XOR U87555 ( .A(n67535), .B(n72121), .Z(n72275) );
  XOR U87556 ( .A(n72276), .B(n72275), .Z(n72114) );
  XOR U87557 ( .A(n67536), .B(n72114), .Z(n72285) );
  XOR U87558 ( .A(n72283), .B(n72285), .Z(n72287) );
  XOR U87559 ( .A(n72286), .B(n72287), .Z(n72291) );
  XOR U87560 ( .A(n72290), .B(n72291), .Z(n72295) );
  XOR U87561 ( .A(n67537), .B(n72295), .Z(n72298) );
  IV U87562 ( .A(n67538), .Z(n67540) );
  NOR U87563 ( .A(n67540), .B(n67539), .Z(n72297) );
  IV U87564 ( .A(n67541), .Z(n67543) );
  NOR U87565 ( .A(n67543), .B(n67542), .Z(n72300) );
  NOR U87566 ( .A(n72297), .B(n72300), .Z(n67544) );
  XOR U87567 ( .A(n72298), .B(n67544), .Z(n72305) );
  XOR U87568 ( .A(n72303), .B(n72305), .Z(n72307) );
  XOR U87569 ( .A(n72306), .B(n72307), .Z(n72312) );
  XOR U87570 ( .A(n72310), .B(n72312), .Z(n72314) );
  XOR U87571 ( .A(n72313), .B(n72314), .Z(n72109) );
  XOR U87572 ( .A(n67545), .B(n72109), .Z(n67546) );
  IV U87573 ( .A(n67546), .Z(n72318) );
  XOR U87574 ( .A(n72317), .B(n72318), .Z(n72321) );
  XOR U87575 ( .A(n72320), .B(n72321), .Z(n72328) );
  IV U87576 ( .A(n67547), .Z(n67548) );
  NOR U87577 ( .A(n67549), .B(n67548), .Z(n72327) );
  NOR U87578 ( .A(n72325), .B(n72327), .Z(n67550) );
  XOR U87579 ( .A(n72328), .B(n67550), .Z(n72101) );
  XOR U87580 ( .A(n67551), .B(n72101), .Z(n72096) );
  XOR U87581 ( .A(n72094), .B(n72096), .Z(n72098) );
  IV U87582 ( .A(n67552), .Z(n67553) );
  NOR U87583 ( .A(n67554), .B(n67553), .Z(n72097) );
  IV U87584 ( .A(n67555), .Z(n67556) );
  NOR U87585 ( .A(n67560), .B(n67556), .Z(n72092) );
  NOR U87586 ( .A(n72097), .B(n72092), .Z(n67557) );
  XOR U87587 ( .A(n72098), .B(n67557), .Z(n67558) );
  IV U87588 ( .A(n67558), .Z(n72340) );
  IV U87589 ( .A(n67559), .Z(n67561) );
  NOR U87590 ( .A(n67561), .B(n67560), .Z(n72338) );
  XOR U87591 ( .A(n72340), .B(n72338), .Z(n72343) );
  XOR U87592 ( .A(n72341), .B(n72343), .Z(n72348) );
  XOR U87593 ( .A(n72346), .B(n72348), .Z(n72350) );
  XOR U87594 ( .A(n72349), .B(n72350), .Z(n72090) );
  XOR U87595 ( .A(n72089), .B(n72090), .Z(n72084) );
  XOR U87596 ( .A(n72083), .B(n72084), .Z(n72087) );
  XOR U87597 ( .A(n72086), .B(n72087), .Z(n72082) );
  XOR U87598 ( .A(n72080), .B(n72082), .Z(n72360) );
  XOR U87599 ( .A(n72358), .B(n72360), .Z(n72363) );
  XOR U87600 ( .A(n72361), .B(n72363), .Z(n72375) );
  XOR U87601 ( .A(n72374), .B(n72375), .Z(n72378) );
  XOR U87602 ( .A(n72377), .B(n72378), .Z(n72382) );
  XOR U87603 ( .A(n72381), .B(n72382), .Z(n72388) );
  XOR U87604 ( .A(n67562), .B(n72388), .Z(n67563) );
  IV U87605 ( .A(n67563), .Z(n72399) );
  XOR U87606 ( .A(n67564), .B(n72399), .Z(n72406) );
  IV U87607 ( .A(n67565), .Z(n67566) );
  NOR U87608 ( .A(n67567), .B(n67566), .Z(n72398) );
  IV U87609 ( .A(n67568), .Z(n67570) );
  NOR U87610 ( .A(n67570), .B(n67569), .Z(n72405) );
  NOR U87611 ( .A(n72398), .B(n72405), .Z(n67571) );
  XOR U87612 ( .A(n72406), .B(n67571), .Z(n72402) );
  XOR U87613 ( .A(n72403), .B(n72402), .Z(n72413) );
  XOR U87614 ( .A(n67572), .B(n72413), .Z(n72076) );
  IV U87615 ( .A(n67573), .Z(n67575) );
  NOR U87616 ( .A(n67575), .B(n67574), .Z(n72074) );
  XOR U87617 ( .A(n72076), .B(n72074), .Z(n72409) );
  XOR U87618 ( .A(n72408), .B(n72409), .Z(n77565) );
  XOR U87619 ( .A(n72419), .B(n77565), .Z(n67576) );
  IV U87620 ( .A(n67576), .Z(n72422) );
  XOR U87621 ( .A(n72420), .B(n72422), .Z(n72427) );
  XOR U87622 ( .A(n72425), .B(n72427), .Z(n72429) );
  XOR U87623 ( .A(n72428), .B(n72429), .Z(n72439) );
  XOR U87624 ( .A(n67577), .B(n72439), .Z(n67578) );
  IV U87625 ( .A(n67578), .Z(n72437) );
  XOR U87626 ( .A(n72435), .B(n72437), .Z(n72070) );
  XOR U87627 ( .A(n72069), .B(n72070), .Z(n72443) );
  IV U87628 ( .A(n67579), .Z(n67580) );
  NOR U87629 ( .A(n67581), .B(n67580), .Z(n72072) );
  IV U87630 ( .A(n67582), .Z(n67583) );
  NOR U87631 ( .A(n67583), .B(n67589), .Z(n72441) );
  NOR U87632 ( .A(n72072), .B(n72441), .Z(n67584) );
  XOR U87633 ( .A(n72443), .B(n67584), .Z(n72444) );
  IV U87634 ( .A(n67585), .Z(n67587) );
  NOR U87635 ( .A(n67587), .B(n67586), .Z(n77895) );
  IV U87636 ( .A(n67588), .Z(n67590) );
  NOR U87637 ( .A(n67590), .B(n67589), .Z(n77886) );
  NOR U87638 ( .A(n77895), .B(n77886), .Z(n72445) );
  XOR U87639 ( .A(n72444), .B(n72445), .Z(n72454) );
  IV U87640 ( .A(n67591), .Z(n67592) );
  NOR U87641 ( .A(n67592), .B(n67594), .Z(n72446) );
  IV U87642 ( .A(n67593), .Z(n67595) );
  NOR U87643 ( .A(n67595), .B(n67594), .Z(n72453) );
  NOR U87644 ( .A(n72446), .B(n72453), .Z(n67596) );
  XOR U87645 ( .A(n72454), .B(n67596), .Z(n72450) );
  IV U87646 ( .A(n67597), .Z(n67599) );
  NOR U87647 ( .A(n67599), .B(n67598), .Z(n72457) );
  NOR U87648 ( .A(n72451), .B(n72457), .Z(n67600) );
  XOR U87649 ( .A(n72450), .B(n67600), .Z(n72068) );
  IV U87650 ( .A(n67601), .Z(n67602) );
  NOR U87651 ( .A(n67602), .B(n67608), .Z(n72066) );
  XOR U87652 ( .A(n72068), .B(n72066), .Z(n77907) );
  IV U87653 ( .A(n67603), .Z(n67605) );
  NOR U87654 ( .A(n67605), .B(n67604), .Z(n77911) );
  IV U87655 ( .A(n67606), .Z(n67607) );
  NOR U87656 ( .A(n67608), .B(n67607), .Z(n77905) );
  NOR U87657 ( .A(n77911), .B(n77905), .Z(n72460) );
  XOR U87658 ( .A(n77907), .B(n72460), .Z(n72462) );
  XOR U87659 ( .A(n67609), .B(n72462), .Z(n72477) );
  XOR U87660 ( .A(n72475), .B(n72477), .Z(n72479) );
  IV U87661 ( .A(n72479), .Z(n67617) );
  IV U87662 ( .A(n67610), .Z(n67611) );
  NOR U87663 ( .A(n67612), .B(n67611), .Z(n72478) );
  IV U87664 ( .A(n67613), .Z(n67615) );
  NOR U87665 ( .A(n67615), .B(n67614), .Z(n72063) );
  NOR U87666 ( .A(n72478), .B(n72063), .Z(n67616) );
  XOR U87667 ( .A(n67617), .B(n67616), .Z(n72058) );
  XOR U87668 ( .A(n72057), .B(n72058), .Z(n72061) );
  XOR U87669 ( .A(n72060), .B(n72061), .Z(n77932) );
  XOR U87670 ( .A(n72056), .B(n77932), .Z(n72483) );
  XOR U87671 ( .A(n72485), .B(n72483), .Z(n72487) );
  IV U87672 ( .A(n67618), .Z(n67619) );
  NOR U87673 ( .A(n67620), .B(n67619), .Z(n72486) );
  IV U87674 ( .A(n67621), .Z(n67622) );
  NOR U87675 ( .A(n67623), .B(n67622), .Z(n72054) );
  NOR U87676 ( .A(n72486), .B(n72054), .Z(n67624) );
  XOR U87677 ( .A(n72487), .B(n67624), .Z(n72048) );
  IV U87678 ( .A(n67625), .Z(n67627) );
  NOR U87679 ( .A(n67627), .B(n67626), .Z(n72051) );
  NOR U87680 ( .A(n72051), .B(n72049), .Z(n67628) );
  XOR U87681 ( .A(n72048), .B(n67628), .Z(n72046) );
  XOR U87682 ( .A(n72045), .B(n72046), .Z(n77973) );
  IV U87683 ( .A(n67629), .Z(n67630) );
  NOR U87684 ( .A(n67631), .B(n67630), .Z(n77977) );
  IV U87685 ( .A(n67632), .Z(n67633) );
  NOR U87686 ( .A(n67634), .B(n67633), .Z(n77971) );
  NOR U87687 ( .A(n77977), .B(n77971), .Z(n72500) );
  XOR U87688 ( .A(n77973), .B(n72500), .Z(n72502) );
  XOR U87689 ( .A(n67635), .B(n72502), .Z(n72515) );
  XOR U87690 ( .A(n67636), .B(n72515), .Z(n72511) );
  XOR U87691 ( .A(n67637), .B(n72511), .Z(n72518) );
  IV U87692 ( .A(n67638), .Z(n67640) );
  NOR U87693 ( .A(n67640), .B(n67639), .Z(n77998) );
  NOR U87694 ( .A(n77998), .B(n77523), .Z(n72519) );
  XOR U87695 ( .A(n72518), .B(n72519), .Z(n72521) );
  XOR U87696 ( .A(n72520), .B(n72521), .Z(n77519) );
  IV U87697 ( .A(n77519), .Z(n67641) );
  NOR U87698 ( .A(n67642), .B(n67641), .Z(n67652) );
  IV U87699 ( .A(n67643), .Z(n67646) );
  NOR U87700 ( .A(n67644), .B(n72521), .Z(n67645) );
  IV U87701 ( .A(n67645), .Z(n67648) );
  NOR U87702 ( .A(n67646), .B(n67648), .Z(n78006) );
  IV U87703 ( .A(n67647), .Z(n67649) );
  NOR U87704 ( .A(n67649), .B(n67648), .Z(n72040) );
  NOR U87705 ( .A(n78006), .B(n72040), .Z(n67650) );
  IV U87706 ( .A(n67650), .Z(n67651) );
  NOR U87707 ( .A(n67652), .B(n67651), .Z(n67653) );
  IV U87708 ( .A(n67653), .Z(n72037) );
  XOR U87709 ( .A(n72034), .B(n72037), .Z(n72031) );
  IV U87710 ( .A(n67654), .Z(n67656) );
  NOR U87711 ( .A(n67656), .B(n67655), .Z(n72036) );
  IV U87712 ( .A(n67657), .Z(n67658) );
  NOR U87713 ( .A(n67658), .B(n78031), .Z(n72030) );
  NOR U87714 ( .A(n72036), .B(n72030), .Z(n67659) );
  XOR U87715 ( .A(n72031), .B(n67659), .Z(n78030) );
  IV U87716 ( .A(n67660), .Z(n78026) );
  NOR U87717 ( .A(n78026), .B(n67665), .Z(n72526) );
  IV U87718 ( .A(n67661), .Z(n67662) );
  NOR U87719 ( .A(n67662), .B(n78031), .Z(n72029) );
  NOR U87720 ( .A(n72526), .B(n72029), .Z(n67663) );
  XOR U87721 ( .A(n78030), .B(n67663), .Z(n77509) );
  IV U87722 ( .A(n67664), .Z(n67666) );
  NOR U87723 ( .A(n67666), .B(n67665), .Z(n77512) );
  IV U87724 ( .A(n67667), .Z(n67669) );
  NOR U87725 ( .A(n67669), .B(n67668), .Z(n77507) );
  NOR U87726 ( .A(n77512), .B(n77507), .Z(n72529) );
  XOR U87727 ( .A(n77509), .B(n72529), .Z(n72023) );
  XOR U87728 ( .A(n72024), .B(n72023), .Z(n72028) );
  XOR U87729 ( .A(n72026), .B(n72028), .Z(n72535) );
  XOR U87730 ( .A(n72533), .B(n72535), .Z(n72537) );
  XOR U87731 ( .A(n67670), .B(n72537), .Z(n72017) );
  XOR U87732 ( .A(n72015), .B(n72017), .Z(n72019) );
  XOR U87733 ( .A(n72018), .B(n72019), .Z(n72544) );
  IV U87734 ( .A(n67671), .Z(n67674) );
  IV U87735 ( .A(n67673), .Z(n67679) );
  NOR U87736 ( .A(n67674), .B(n67679), .Z(n72013) );
  IV U87737 ( .A(n67672), .Z(n67676) );
  XOR U87738 ( .A(n67674), .B(n67673), .Z(n67675) );
  NOR U87739 ( .A(n67676), .B(n67675), .Z(n72543) );
  NOR U87740 ( .A(n72013), .B(n72543), .Z(n67677) );
  XOR U87741 ( .A(n72544), .B(n67677), .Z(n72007) );
  IV U87742 ( .A(n67678), .Z(n67680) );
  NOR U87743 ( .A(n67680), .B(n67679), .Z(n72010) );
  IV U87744 ( .A(n67681), .Z(n67682) );
  NOR U87745 ( .A(n67682), .B(n67685), .Z(n72008) );
  NOR U87746 ( .A(n72010), .B(n72008), .Z(n67683) );
  XOR U87747 ( .A(n72007), .B(n67683), .Z(n72548) );
  IV U87748 ( .A(n67684), .Z(n67686) );
  NOR U87749 ( .A(n67686), .B(n67685), .Z(n72546) );
  XOR U87750 ( .A(n72548), .B(n72546), .Z(n72004) );
  XOR U87751 ( .A(n72003), .B(n72004), .Z(n72565) );
  IV U87752 ( .A(n67687), .Z(n67689) );
  NOR U87753 ( .A(n67689), .B(n67688), .Z(n72553) );
  IV U87754 ( .A(n67690), .Z(n67692) );
  NOR U87755 ( .A(n67692), .B(n67691), .Z(n72564) );
  NOR U87756 ( .A(n72553), .B(n72564), .Z(n67693) );
  XOR U87757 ( .A(n72565), .B(n67693), .Z(n72000) );
  IV U87758 ( .A(n67694), .Z(n67696) );
  NOR U87759 ( .A(n67696), .B(n67695), .Z(n72561) );
  IV U87760 ( .A(n67697), .Z(n67698) );
  NOR U87761 ( .A(n67698), .B(n67701), .Z(n72001) );
  NOR U87762 ( .A(n72561), .B(n72001), .Z(n67699) );
  XOR U87763 ( .A(n72000), .B(n67699), .Z(n71999) );
  IV U87764 ( .A(n67700), .Z(n67702) );
  NOR U87765 ( .A(n67702), .B(n67701), .Z(n71997) );
  XOR U87766 ( .A(n71999), .B(n71997), .Z(n71994) );
  NOR U87767 ( .A(n67704), .B(n67703), .Z(n71993) );
  IV U87768 ( .A(n67705), .Z(n67706) );
  NOR U87769 ( .A(n67714), .B(n67706), .Z(n71991) );
  NOR U87770 ( .A(n71993), .B(n71991), .Z(n67707) );
  XOR U87771 ( .A(n71994), .B(n67707), .Z(n67708) );
  IV U87772 ( .A(n67708), .Z(n71987) );
  IV U87773 ( .A(n67709), .Z(n67711) );
  NOR U87774 ( .A(n67711), .B(n67710), .Z(n67712) );
  IV U87775 ( .A(n67712), .Z(n67716) );
  NOR U87776 ( .A(n71987), .B(n67716), .Z(n78057) );
  IV U87777 ( .A(n67713), .Z(n67715) );
  NOR U87778 ( .A(n67715), .B(n67714), .Z(n71988) );
  XOR U87779 ( .A(n71985), .B(n71987), .Z(n71989) );
  IV U87780 ( .A(n71989), .Z(n67717) );
  XOR U87781 ( .A(n71988), .B(n67717), .Z(n67719) );
  NOR U87782 ( .A(n67717), .B(n67716), .Z(n67718) );
  NOR U87783 ( .A(n67719), .B(n67718), .Z(n67720) );
  NOR U87784 ( .A(n78057), .B(n67720), .Z(n67721) );
  IV U87785 ( .A(n67721), .Z(n78061) );
  XOR U87786 ( .A(n71979), .B(n78061), .Z(n71972) );
  NOR U87787 ( .A(n67722), .B(n71976), .Z(n67725) );
  NOR U87788 ( .A(n67724), .B(n67723), .Z(n71971) );
  NOR U87789 ( .A(n67725), .B(n71971), .Z(n67726) );
  XOR U87790 ( .A(n71972), .B(n67726), .Z(n72579) );
  XOR U87791 ( .A(n72577), .B(n72579), .Z(n72575) );
  XOR U87792 ( .A(n67727), .B(n72575), .Z(n71968) );
  XOR U87793 ( .A(n71967), .B(n71968), .Z(n72608) );
  IV U87794 ( .A(n67728), .Z(n67730) );
  NOR U87795 ( .A(n67730), .B(n67729), .Z(n72599) );
  IV U87796 ( .A(n67731), .Z(n67732) );
  NOR U87797 ( .A(n67733), .B(n67732), .Z(n72607) );
  NOR U87798 ( .A(n72599), .B(n72607), .Z(n67734) );
  XOR U87799 ( .A(n72608), .B(n67734), .Z(n72601) );
  IV U87800 ( .A(n67735), .Z(n67736) );
  NOR U87801 ( .A(n67737), .B(n67736), .Z(n72604) );
  IV U87802 ( .A(n67738), .Z(n67740) );
  NOR U87803 ( .A(n67740), .B(n67739), .Z(n72602) );
  NOR U87804 ( .A(n72604), .B(n72602), .Z(n67741) );
  XOR U87805 ( .A(n72601), .B(n67741), .Z(n72613) );
  XOR U87806 ( .A(n72612), .B(n72613), .Z(n72617) );
  IV U87807 ( .A(n67742), .Z(n67744) );
  NOR U87808 ( .A(n67744), .B(n67743), .Z(n72615) );
  XOR U87809 ( .A(n72617), .B(n72615), .Z(n71962) );
  XOR U87810 ( .A(n71963), .B(n71962), .Z(n71960) );
  IV U87811 ( .A(n67745), .Z(n67747) );
  NOR U87812 ( .A(n67747), .B(n67746), .Z(n71964) );
  IV U87813 ( .A(n67748), .Z(n67749) );
  NOR U87814 ( .A(n67750), .B(n67749), .Z(n71959) );
  NOR U87815 ( .A(n71964), .B(n71959), .Z(n67751) );
  XOR U87816 ( .A(n71960), .B(n67751), .Z(n71957) );
  XOR U87817 ( .A(n71956), .B(n71957), .Z(n72621) );
  XOR U87818 ( .A(n72620), .B(n72621), .Z(n72624) );
  XOR U87819 ( .A(n72623), .B(n72624), .Z(n71955) );
  XOR U87820 ( .A(n71953), .B(n71955), .Z(n72632) );
  XOR U87821 ( .A(n67752), .B(n72632), .Z(n67753) );
  IV U87822 ( .A(n67753), .Z(n71943) );
  XOR U87823 ( .A(n71942), .B(n71943), .Z(n72638) );
  IV U87824 ( .A(n67754), .Z(n67764) );
  IV U87825 ( .A(n67755), .Z(n67756) );
  NOR U87826 ( .A(n67764), .B(n67756), .Z(n71945) );
  NOR U87827 ( .A(n72637), .B(n71945), .Z(n67757) );
  XOR U87828 ( .A(n72638), .B(n67757), .Z(n71933) );
  IV U87829 ( .A(n67758), .Z(n67762) );
  NOR U87830 ( .A(n67760), .B(n67759), .Z(n67761) );
  IV U87831 ( .A(n67761), .Z(n67768) );
  NOR U87832 ( .A(n67762), .B(n67768), .Z(n71934) );
  IV U87833 ( .A(n67763), .Z(n67765) );
  NOR U87834 ( .A(n67765), .B(n67764), .Z(n71939) );
  NOR U87835 ( .A(n71934), .B(n71939), .Z(n67766) );
  XOR U87836 ( .A(n71933), .B(n67766), .Z(n71938) );
  IV U87837 ( .A(n67767), .Z(n67769) );
  NOR U87838 ( .A(n67769), .B(n67768), .Z(n71936) );
  XOR U87839 ( .A(n71938), .B(n71936), .Z(n78127) );
  XOR U87840 ( .A(n78129), .B(n78127), .Z(n67779) );
  XOR U87841 ( .A(n72643), .B(n67779), .Z(n67776) );
  IV U87842 ( .A(n67776), .Z(n67770) );
  NOR U87843 ( .A(n67789), .B(n67770), .Z(n77432) );
  IV U87844 ( .A(n67771), .Z(n67772) );
  NOR U87845 ( .A(n67773), .B(n67772), .Z(n72649) );
  IV U87846 ( .A(n67774), .Z(n67780) );
  NOR U87847 ( .A(n67775), .B(n67780), .Z(n67777) );
  NOR U87848 ( .A(n67777), .B(n67776), .Z(n67788) );
  IV U87849 ( .A(n67778), .Z(n67782) );
  IV U87850 ( .A(n67779), .Z(n72644) );
  NOR U87851 ( .A(n67780), .B(n72644), .Z(n67781) );
  IV U87852 ( .A(n67781), .Z(n67784) );
  NOR U87853 ( .A(n67782), .B(n67784), .Z(n77437) );
  IV U87854 ( .A(n67783), .Z(n67785) );
  NOR U87855 ( .A(n67785), .B(n67784), .Z(n77434) );
  NOR U87856 ( .A(n77437), .B(n77434), .Z(n67786) );
  IV U87857 ( .A(n67786), .Z(n67787) );
  NOR U87858 ( .A(n67788), .B(n67787), .Z(n72650) );
  XOR U87859 ( .A(n72649), .B(n72650), .Z(n67791) );
  NOR U87860 ( .A(n72650), .B(n67789), .Z(n67790) );
  NOR U87861 ( .A(n67791), .B(n67790), .Z(n67792) );
  NOR U87862 ( .A(n77432), .B(n67792), .Z(n67793) );
  IV U87863 ( .A(n67793), .Z(n72657) );
  XOR U87864 ( .A(n72653), .B(n72657), .Z(n71930) );
  IV U87865 ( .A(n67794), .Z(n67795) );
  NOR U87866 ( .A(n67796), .B(n67795), .Z(n72656) );
  NOR U87867 ( .A(n72656), .B(n67797), .Z(n67798) );
  XOR U87868 ( .A(n71930), .B(n67798), .Z(n71924) );
  XOR U87869 ( .A(n71925), .B(n71924), .Z(n72661) );
  XOR U87870 ( .A(n72660), .B(n72661), .Z(n72664) );
  XOR U87871 ( .A(n67799), .B(n72664), .Z(n67800) );
  IV U87872 ( .A(n67800), .Z(n71922) );
  XOR U87873 ( .A(n71921), .B(n71922), .Z(n71917) );
  XOR U87874 ( .A(n71916), .B(n71917), .Z(n77417) );
  IV U87875 ( .A(n67801), .Z(n78168) );
  NOR U87876 ( .A(n67802), .B(n78168), .Z(n72672) );
  IV U87877 ( .A(n67803), .Z(n67804) );
  NOR U87878 ( .A(n67805), .B(n67804), .Z(n72669) );
  NOR U87879 ( .A(n72672), .B(n72669), .Z(n67806) );
  XOR U87880 ( .A(n77417), .B(n67806), .Z(n72680) );
  XOR U87881 ( .A(n67807), .B(n72680), .Z(n71915) );
  IV U87882 ( .A(n67808), .Z(n67810) );
  NOR U87883 ( .A(n67810), .B(n67809), .Z(n71913) );
  IV U87884 ( .A(n67811), .Z(n67812) );
  NOR U87885 ( .A(n67813), .B(n67812), .Z(n71911) );
  NOR U87886 ( .A(n71913), .B(n71911), .Z(n67814) );
  XOR U87887 ( .A(n71915), .B(n67814), .Z(n71906) );
  XOR U87888 ( .A(n71908), .B(n71906), .Z(n72687) );
  IV U87889 ( .A(n67815), .Z(n67817) );
  NOR U87890 ( .A(n67817), .B(n67816), .Z(n71909) );
  IV U87891 ( .A(n67818), .Z(n67819) );
  NOR U87892 ( .A(n67820), .B(n67819), .Z(n72686) );
  NOR U87893 ( .A(n71909), .B(n72686), .Z(n67821) );
  XOR U87894 ( .A(n72687), .B(n67821), .Z(n72684) );
  IV U87895 ( .A(n67822), .Z(n67823) );
  NOR U87896 ( .A(n67824), .B(n67823), .Z(n78188) );
  IV U87897 ( .A(n67825), .Z(n67826) );
  NOR U87898 ( .A(n67826), .B(n67834), .Z(n78193) );
  NOR U87899 ( .A(n78188), .B(n78193), .Z(n72685) );
  XOR U87900 ( .A(n72684), .B(n72685), .Z(n71905) );
  IV U87901 ( .A(n71905), .Z(n67837) );
  IV U87902 ( .A(n67827), .Z(n67832) );
  NOR U87903 ( .A(n67829), .B(n67828), .Z(n67830) );
  IV U87904 ( .A(n67830), .Z(n67831) );
  NOR U87905 ( .A(n67832), .B(n67831), .Z(n71901) );
  IV U87906 ( .A(n67833), .Z(n67835) );
  NOR U87907 ( .A(n67835), .B(n67834), .Z(n71903) );
  NOR U87908 ( .A(n71901), .B(n71903), .Z(n67836) );
  XOR U87909 ( .A(n67837), .B(n67836), .Z(n72694) );
  XOR U87910 ( .A(n72692), .B(n72694), .Z(n71900) );
  XOR U87911 ( .A(n71898), .B(n71900), .Z(n72697) );
  XOR U87912 ( .A(n72695), .B(n72697), .Z(n72705) );
  XOR U87913 ( .A(n67838), .B(n72705), .Z(n71891) );
  XOR U87914 ( .A(n71894), .B(n71891), .Z(n72717) );
  IV U87915 ( .A(n67839), .Z(n67841) );
  NOR U87916 ( .A(n67841), .B(n67840), .Z(n71892) );
  IV U87917 ( .A(n67842), .Z(n67843) );
  NOR U87918 ( .A(n67843), .B(n67847), .Z(n72716) );
  NOR U87919 ( .A(n71892), .B(n72716), .Z(n67844) );
  XOR U87920 ( .A(n72717), .B(n67844), .Z(n71882) );
  IV U87921 ( .A(n67845), .Z(n67846) );
  NOR U87922 ( .A(n67847), .B(n67846), .Z(n71888) );
  IV U87923 ( .A(n67848), .Z(n67852) );
  IV U87924 ( .A(n67849), .Z(n67861) );
  NOR U87925 ( .A(n67850), .B(n67861), .Z(n67851) );
  IV U87926 ( .A(n67851), .Z(n67857) );
  NOR U87927 ( .A(n67852), .B(n67857), .Z(n71883) );
  NOR U87928 ( .A(n71888), .B(n71883), .Z(n67853) );
  XOR U87929 ( .A(n71882), .B(n67853), .Z(n71886) );
  IV U87930 ( .A(n67854), .Z(n67855) );
  NOR U87931 ( .A(n67855), .B(n67861), .Z(n71880) );
  IV U87932 ( .A(n67856), .Z(n67858) );
  NOR U87933 ( .A(n67858), .B(n67857), .Z(n71885) );
  NOR U87934 ( .A(n71880), .B(n71885), .Z(n67859) );
  XOR U87935 ( .A(n71886), .B(n67859), .Z(n72723) );
  IV U87936 ( .A(n67860), .Z(n67862) );
  NOR U87937 ( .A(n67862), .B(n67861), .Z(n77376) );
  IV U87938 ( .A(n67863), .Z(n67864) );
  NOR U87939 ( .A(n67867), .B(n67864), .Z(n77369) );
  NOR U87940 ( .A(n77376), .B(n77369), .Z(n72724) );
  XOR U87941 ( .A(n72723), .B(n72724), .Z(n71878) );
  IV U87942 ( .A(n67865), .Z(n67866) );
  NOR U87943 ( .A(n67867), .B(n67866), .Z(n71876) );
  XOR U87944 ( .A(n71878), .B(n71876), .Z(n72721) );
  XOR U87945 ( .A(n72720), .B(n72721), .Z(n71872) );
  IV U87946 ( .A(n67868), .Z(n67871) );
  IV U87947 ( .A(n67869), .Z(n67870) );
  NOR U87948 ( .A(n67871), .B(n67870), .Z(n71870) );
  XOR U87949 ( .A(n71872), .B(n71870), .Z(n78209) );
  XOR U87950 ( .A(n71873), .B(n78209), .Z(n71869) );
  IV U87951 ( .A(n67872), .Z(n67875) );
  NOR U87952 ( .A(n78221), .B(n67873), .Z(n67874) );
  IV U87953 ( .A(n67874), .Z(n67877) );
  NOR U87954 ( .A(n67875), .B(n67877), .Z(n71867) );
  XOR U87955 ( .A(n71869), .B(n71867), .Z(n72733) );
  IV U87956 ( .A(n67876), .Z(n67878) );
  NOR U87957 ( .A(n67878), .B(n67877), .Z(n72731) );
  XOR U87958 ( .A(n72733), .B(n72731), .Z(n72735) );
  XOR U87959 ( .A(n72734), .B(n72735), .Z(n72741) );
  IV U87960 ( .A(n67879), .Z(n67883) );
  NOR U87961 ( .A(n67881), .B(n67880), .Z(n67882) );
  IV U87962 ( .A(n67882), .Z(n67885) );
  NOR U87963 ( .A(n67883), .B(n67885), .Z(n72739) );
  XOR U87964 ( .A(n72741), .B(n72739), .Z(n72744) );
  IV U87965 ( .A(n67884), .Z(n67886) );
  NOR U87966 ( .A(n67886), .B(n67885), .Z(n72742) );
  XOR U87967 ( .A(n72744), .B(n72742), .Z(n71865) );
  NOR U87968 ( .A(n67888), .B(n67887), .Z(n71864) );
  NOR U87969 ( .A(n67890), .B(n67889), .Z(n71862) );
  NOR U87970 ( .A(n71864), .B(n71862), .Z(n67891) );
  XOR U87971 ( .A(n71865), .B(n67891), .Z(n67892) );
  IV U87972 ( .A(n67892), .Z(n72753) );
  XOR U87973 ( .A(n72752), .B(n72753), .Z(n72756) );
  XOR U87974 ( .A(n67893), .B(n72756), .Z(n71860) );
  XOR U87975 ( .A(n71861), .B(n71860), .Z(n72765) );
  IV U87976 ( .A(n72765), .Z(n67900) );
  IV U87977 ( .A(n67894), .Z(n67895) );
  NOR U87978 ( .A(n67897), .B(n67895), .Z(n72763) );
  IV U87979 ( .A(n67896), .Z(n67898) );
  NOR U87980 ( .A(n67898), .B(n67897), .Z(n72760) );
  NOR U87981 ( .A(n72763), .B(n72760), .Z(n67899) );
  XOR U87982 ( .A(n67900), .B(n67899), .Z(n72774) );
  XOR U87983 ( .A(n72770), .B(n72774), .Z(n72767) );
  XOR U87984 ( .A(n67901), .B(n72767), .Z(n71855) );
  XOR U87985 ( .A(n67902), .B(n71855), .Z(n78246) );
  XOR U87986 ( .A(n72787), .B(n78246), .Z(n67909) );
  IV U87987 ( .A(n67909), .Z(n72788) );
  NOR U87988 ( .A(n67910), .B(n72788), .Z(n77325) );
  IV U87989 ( .A(n67903), .Z(n67905) );
  NOR U87990 ( .A(n67905), .B(n67904), .Z(n71850) );
  NOR U87991 ( .A(n67907), .B(n67906), .Z(n67908) );
  IV U87992 ( .A(n67908), .Z(n72789) );
  XOR U87993 ( .A(n72789), .B(n67909), .Z(n71851) );
  IV U87994 ( .A(n71851), .Z(n67911) );
  XOR U87995 ( .A(n71850), .B(n67911), .Z(n67913) );
  NOR U87996 ( .A(n67911), .B(n67910), .Z(n67912) );
  NOR U87997 ( .A(n67913), .B(n67912), .Z(n67914) );
  NOR U87998 ( .A(n77325), .B(n67914), .Z(n71843) );
  XOR U87999 ( .A(n67915), .B(n71843), .Z(n71841) );
  XOR U88000 ( .A(n67916), .B(n71841), .Z(n72796) );
  XOR U88001 ( .A(n72797), .B(n72796), .Z(n72800) );
  XOR U88002 ( .A(n72799), .B(n72800), .Z(n78273) );
  XOR U88003 ( .A(n84108), .B(n78273), .Z(n67917) );
  IV U88004 ( .A(n67917), .Z(n72815) );
  IV U88005 ( .A(n67918), .Z(n67919) );
  NOR U88006 ( .A(n67919), .B(n67923), .Z(n72813) );
  XOR U88007 ( .A(n72815), .B(n72813), .Z(n72819) );
  IV U88008 ( .A(n67920), .Z(n67921) );
  NOR U88009 ( .A(n67929), .B(n67921), .Z(n72818) );
  IV U88010 ( .A(n67922), .Z(n67924) );
  NOR U88011 ( .A(n67924), .B(n67923), .Z(n71837) );
  NOR U88012 ( .A(n72818), .B(n71837), .Z(n67925) );
  XOR U88013 ( .A(n72819), .B(n67925), .Z(n67926) );
  IV U88014 ( .A(n67926), .Z(n72823) );
  IV U88015 ( .A(n67927), .Z(n67928) );
  NOR U88016 ( .A(n67929), .B(n67928), .Z(n72821) );
  XOR U88017 ( .A(n72823), .B(n72821), .Z(n72834) );
  XOR U88018 ( .A(n67930), .B(n72834), .Z(n67931) );
  IV U88019 ( .A(n67931), .Z(n72832) );
  IV U88020 ( .A(n67932), .Z(n67936) );
  NOR U88021 ( .A(n67934), .B(n67933), .Z(n67935) );
  IV U88022 ( .A(n67935), .Z(n67938) );
  NOR U88023 ( .A(n67936), .B(n67938), .Z(n72830) );
  XOR U88024 ( .A(n72832), .B(n72830), .Z(n72829) );
  IV U88025 ( .A(n67937), .Z(n67939) );
  NOR U88026 ( .A(n67939), .B(n67938), .Z(n72827) );
  XOR U88027 ( .A(n72829), .B(n72827), .Z(n72846) );
  IV U88028 ( .A(n72846), .Z(n67949) );
  IV U88029 ( .A(n67940), .Z(n67941) );
  NOR U88030 ( .A(n67941), .B(n67943), .Z(n71835) );
  IV U88031 ( .A(n67942), .Z(n67944) );
  NOR U88032 ( .A(n67944), .B(n67943), .Z(n72845) );
  NOR U88033 ( .A(n71835), .B(n72845), .Z(n67945) );
  IV U88034 ( .A(n67945), .Z(n67946) );
  NOR U88035 ( .A(n67947), .B(n67946), .Z(n67948) );
  XOR U88036 ( .A(n67949), .B(n67948), .Z(n72844) );
  XOR U88037 ( .A(n72842), .B(n72844), .Z(n71832) );
  XOR U88038 ( .A(n67950), .B(n71832), .Z(n71827) );
  XOR U88039 ( .A(n67951), .B(n71827), .Z(n72855) );
  XOR U88040 ( .A(n72857), .B(n72855), .Z(n67952) );
  IV U88041 ( .A(n67952), .Z(n72861) );
  XOR U88042 ( .A(n72860), .B(n72861), .Z(n72865) );
  IV U88043 ( .A(n67953), .Z(n67955) );
  IV U88044 ( .A(n67954), .Z(n67957) );
  NOR U88045 ( .A(n67955), .B(n67957), .Z(n72863) );
  XOR U88046 ( .A(n72865), .B(n72863), .Z(n72869) );
  IV U88047 ( .A(n67956), .Z(n67958) );
  NOR U88048 ( .A(n67958), .B(n67957), .Z(n72867) );
  XOR U88049 ( .A(n72869), .B(n72867), .Z(n72872) );
  IV U88050 ( .A(n67959), .Z(n67960) );
  NOR U88051 ( .A(n67963), .B(n67960), .Z(n72870) );
  XOR U88052 ( .A(n72872), .B(n72870), .Z(n71825) );
  IV U88053 ( .A(n67961), .Z(n67962) );
  NOR U88054 ( .A(n67963), .B(n67962), .Z(n71823) );
  XOR U88055 ( .A(n71825), .B(n71823), .Z(n67975) );
  IV U88056 ( .A(n67975), .Z(n67971) );
  IV U88057 ( .A(n67964), .Z(n67966) );
  NOR U88058 ( .A(n67966), .B(n67965), .Z(n67972) );
  IV U88059 ( .A(n67967), .Z(n67968) );
  NOR U88060 ( .A(n67968), .B(n67983), .Z(n67974) );
  NOR U88061 ( .A(n67972), .B(n67974), .Z(n67969) );
  IV U88062 ( .A(n67969), .Z(n67970) );
  NOR U88063 ( .A(n67971), .B(n67970), .Z(n67978) );
  IV U88064 ( .A(n67972), .Z(n67973) );
  NOR U88065 ( .A(n67973), .B(n71825), .Z(n83025) );
  IV U88066 ( .A(n67974), .Z(n67976) );
  NOR U88067 ( .A(n67976), .B(n67975), .Z(n83020) );
  NOR U88068 ( .A(n83025), .B(n83020), .Z(n67977) );
  IV U88069 ( .A(n67977), .Z(n71826) );
  NOR U88070 ( .A(n67978), .B(n71826), .Z(n72875) );
  IV U88071 ( .A(n67979), .Z(n67988) );
  IV U88072 ( .A(n67980), .Z(n67981) );
  NOR U88073 ( .A(n67988), .B(n67981), .Z(n72874) );
  IV U88074 ( .A(n67982), .Z(n67984) );
  NOR U88075 ( .A(n67984), .B(n67983), .Z(n72877) );
  NOR U88076 ( .A(n72874), .B(n72877), .Z(n67985) );
  XOR U88077 ( .A(n72875), .B(n67985), .Z(n72889) );
  IV U88078 ( .A(n72889), .Z(n67993) );
  IV U88079 ( .A(n67986), .Z(n67987) );
  NOR U88080 ( .A(n67988), .B(n67987), .Z(n71821) );
  IV U88081 ( .A(n67989), .Z(n67990) );
  NOR U88082 ( .A(n67991), .B(n67990), .Z(n72887) );
  NOR U88083 ( .A(n71821), .B(n72887), .Z(n67992) );
  XOR U88084 ( .A(n67993), .B(n67992), .Z(n71819) );
  XOR U88085 ( .A(n71818), .B(n71819), .Z(n71814) );
  IV U88086 ( .A(n67994), .Z(n67998) );
  NOR U88087 ( .A(n67996), .B(n67995), .Z(n67997) );
  IV U88088 ( .A(n67997), .Z(n68003) );
  NOR U88089 ( .A(n67998), .B(n68003), .Z(n71812) );
  XOR U88090 ( .A(n71814), .B(n71812), .Z(n71817) );
  IV U88091 ( .A(n67999), .Z(n68001) );
  NOR U88092 ( .A(n68001), .B(n68000), .Z(n71810) );
  IV U88093 ( .A(n68002), .Z(n68004) );
  NOR U88094 ( .A(n68004), .B(n68003), .Z(n71815) );
  NOR U88095 ( .A(n71810), .B(n71815), .Z(n68005) );
  XOR U88096 ( .A(n71817), .B(n68005), .Z(n72896) );
  IV U88097 ( .A(n68006), .Z(n68008) );
  NOR U88098 ( .A(n68008), .B(n68007), .Z(n68009) );
  IV U88099 ( .A(n68009), .Z(n72897) );
  XOR U88100 ( .A(n72896), .B(n72897), .Z(n72901) );
  XOR U88101 ( .A(n72899), .B(n72901), .Z(n71808) );
  XOR U88102 ( .A(n68010), .B(n71808), .Z(n71800) );
  IV U88103 ( .A(n68011), .Z(n68012) );
  NOR U88104 ( .A(n68013), .B(n68012), .Z(n71799) );
  IV U88105 ( .A(n68014), .Z(n68016) );
  NOR U88106 ( .A(n68016), .B(n68015), .Z(n71804) );
  NOR U88107 ( .A(n71799), .B(n71804), .Z(n68017) );
  XOR U88108 ( .A(n71800), .B(n68017), .Z(n71798) );
  IV U88109 ( .A(n68018), .Z(n68020) );
  NOR U88110 ( .A(n68020), .B(n68019), .Z(n71796) );
  XOR U88111 ( .A(n71798), .B(n71796), .Z(n71794) );
  NOR U88112 ( .A(n68028), .B(n71794), .Z(n77259) );
  IV U88113 ( .A(n68021), .Z(n68022) );
  NOR U88114 ( .A(n68023), .B(n68022), .Z(n71790) );
  IV U88115 ( .A(n68024), .Z(n68027) );
  IV U88116 ( .A(n68025), .Z(n68026) );
  NOR U88117 ( .A(n68027), .B(n68026), .Z(n71793) );
  XOR U88118 ( .A(n71793), .B(n71794), .Z(n71791) );
  IV U88119 ( .A(n71791), .Z(n68029) );
  XOR U88120 ( .A(n71790), .B(n68029), .Z(n68031) );
  NOR U88121 ( .A(n68029), .B(n68028), .Z(n68030) );
  NOR U88122 ( .A(n68031), .B(n68030), .Z(n68032) );
  NOR U88123 ( .A(n77259), .B(n68032), .Z(n71784) );
  XOR U88124 ( .A(n71786), .B(n71784), .Z(n71788) );
  IV U88125 ( .A(n68033), .Z(n68035) );
  IV U88126 ( .A(n68034), .Z(n68038) );
  NOR U88127 ( .A(n68035), .B(n68038), .Z(n71782) );
  NOR U88128 ( .A(n71787), .B(n71782), .Z(n68036) );
  XOR U88129 ( .A(n71788), .B(n68036), .Z(n71776) );
  IV U88130 ( .A(n68037), .Z(n68039) );
  NOR U88131 ( .A(n68039), .B(n68038), .Z(n71780) );
  XOR U88132 ( .A(n71776), .B(n71780), .Z(n68040) );
  XOR U88133 ( .A(n68041), .B(n68040), .Z(n71774) );
  XOR U88134 ( .A(n71772), .B(n71774), .Z(n68051) );
  IV U88135 ( .A(n68051), .Z(n68049) );
  IV U88136 ( .A(n68042), .Z(n68043) );
  NOR U88137 ( .A(n68044), .B(n68043), .Z(n68050) );
  IV U88138 ( .A(n68045), .Z(n68046) );
  NOR U88139 ( .A(n68046), .B(n68058), .Z(n68053) );
  NOR U88140 ( .A(n68050), .B(n68053), .Z(n68047) );
  IV U88141 ( .A(n68047), .Z(n68048) );
  NOR U88142 ( .A(n68049), .B(n68048), .Z(n68056) );
  IV U88143 ( .A(n68050), .Z(n68052) );
  NOR U88144 ( .A(n68052), .B(n68051), .Z(n78394) );
  IV U88145 ( .A(n68053), .Z(n68054) );
  NOR U88146 ( .A(n71774), .B(n68054), .Z(n78410) );
  NOR U88147 ( .A(n78394), .B(n78410), .Z(n68055) );
  IV U88148 ( .A(n68055), .Z(n77252) );
  NOR U88149 ( .A(n68056), .B(n77252), .Z(n72913) );
  IV U88150 ( .A(n68057), .Z(n68059) );
  NOR U88151 ( .A(n68059), .B(n68058), .Z(n68060) );
  IV U88152 ( .A(n68060), .Z(n72915) );
  XOR U88153 ( .A(n72913), .B(n72915), .Z(n72919) );
  XOR U88154 ( .A(n72917), .B(n72919), .Z(n72922) );
  XOR U88155 ( .A(n72920), .B(n72922), .Z(n72925) );
  XOR U88156 ( .A(n68061), .B(n72925), .Z(n72927) );
  XOR U88157 ( .A(n72928), .B(n72927), .Z(n72930) );
  IV U88158 ( .A(n68062), .Z(n68064) );
  NOR U88159 ( .A(n68064), .B(n68063), .Z(n68065) );
  IV U88160 ( .A(n68065), .Z(n72931) );
  XOR U88161 ( .A(n72930), .B(n72931), .Z(n68066) );
  NOR U88162 ( .A(n68071), .B(n68066), .Z(n68073) );
  IV U88163 ( .A(n68067), .Z(n68069) );
  NOR U88164 ( .A(n68069), .B(n68068), .Z(n68075) );
  IV U88165 ( .A(n68075), .Z(n68070) );
  NOR U88166 ( .A(n68073), .B(n68070), .Z(n78435) );
  IV U88167 ( .A(n68071), .Z(n68072) );
  NOR U88168 ( .A(n72930), .B(n68072), .Z(n78442) );
  NOR U88169 ( .A(n78442), .B(n68073), .Z(n68074) );
  NOR U88170 ( .A(n68075), .B(n68074), .Z(n68076) );
  NOR U88171 ( .A(n78435), .B(n68076), .Z(n68077) );
  IV U88172 ( .A(n68077), .Z(n71765) );
  IV U88173 ( .A(n68078), .Z(n68079) );
  NOR U88174 ( .A(n68080), .B(n68079), .Z(n71764) );
  XOR U88175 ( .A(n71765), .B(n71764), .Z(n71768) );
  XOR U88176 ( .A(n71767), .B(n71768), .Z(n72940) );
  XOR U88177 ( .A(n68081), .B(n72940), .Z(n68082) );
  IV U88178 ( .A(n68082), .Z(n72937) );
  XOR U88179 ( .A(n72935), .B(n72937), .Z(n71757) );
  IV U88180 ( .A(n68083), .Z(n68085) );
  NOR U88181 ( .A(n68085), .B(n68084), .Z(n71755) );
  XOR U88182 ( .A(n71757), .B(n71755), .Z(n71760) );
  IV U88183 ( .A(n68086), .Z(n68090) );
  IV U88184 ( .A(n68087), .Z(n68088) );
  NOR U88185 ( .A(n68090), .B(n68088), .Z(n71758) );
  XOR U88186 ( .A(n71760), .B(n71758), .Z(n72953) );
  NOR U88187 ( .A(n68090), .B(n68089), .Z(n68091) );
  IV U88188 ( .A(n68091), .Z(n68098) );
  XOR U88189 ( .A(n68093), .B(n68092), .Z(n68094) );
  NOR U88190 ( .A(n68095), .B(n68094), .Z(n68096) );
  IV U88191 ( .A(n68096), .Z(n68097) );
  NOR U88192 ( .A(n68098), .B(n68097), .Z(n72951) );
  XOR U88193 ( .A(n72953), .B(n72951), .Z(n72943) );
  XOR U88194 ( .A(n68099), .B(n72943), .Z(n68111) );
  IV U88195 ( .A(n68111), .Z(n68107) );
  NOR U88196 ( .A(n68101), .B(n68100), .Z(n68108) );
  IV U88197 ( .A(n68102), .Z(n68104) );
  NOR U88198 ( .A(n68104), .B(n68103), .Z(n68110) );
  NOR U88199 ( .A(n68108), .B(n68110), .Z(n68105) );
  IV U88200 ( .A(n68105), .Z(n68106) );
  NOR U88201 ( .A(n68107), .B(n68106), .Z(n68114) );
  IV U88202 ( .A(n68108), .Z(n68109) );
  NOR U88203 ( .A(n68109), .B(n72943), .Z(n77233) );
  IV U88204 ( .A(n68110), .Z(n68112) );
  NOR U88205 ( .A(n68112), .B(n68111), .Z(n77230) );
  NOR U88206 ( .A(n77233), .B(n77230), .Z(n68113) );
  IV U88207 ( .A(n68113), .Z(n71754) );
  NOR U88208 ( .A(n68114), .B(n71754), .Z(n71749) );
  IV U88209 ( .A(n68115), .Z(n68117) );
  NOR U88210 ( .A(n68117), .B(n68116), .Z(n71748) );
  NOR U88211 ( .A(n71751), .B(n71748), .Z(n68118) );
  XOR U88212 ( .A(n71749), .B(n68118), .Z(n71747) );
  IV U88213 ( .A(n68119), .Z(n68121) );
  NOR U88214 ( .A(n68121), .B(n68120), .Z(n71745) );
  IV U88215 ( .A(n68122), .Z(n68124) );
  NOR U88216 ( .A(n68124), .B(n68123), .Z(n71742) );
  NOR U88217 ( .A(n71745), .B(n71742), .Z(n68125) );
  XOR U88218 ( .A(n71747), .B(n68125), .Z(n68126) );
  NOR U88219 ( .A(n68127), .B(n68126), .Z(n68130) );
  IV U88220 ( .A(n68127), .Z(n68129) );
  XOR U88221 ( .A(n71745), .B(n71747), .Z(n68128) );
  NOR U88222 ( .A(n68129), .B(n68128), .Z(n77222) );
  NOR U88223 ( .A(n68130), .B(n77222), .Z(n68131) );
  IV U88224 ( .A(n68131), .Z(n72959) );
  NOR U88225 ( .A(n68133), .B(n68132), .Z(n72958) );
  XOR U88226 ( .A(n72959), .B(n72958), .Z(n72962) );
  XOR U88227 ( .A(n72961), .B(n72962), .Z(n72971) );
  XOR U88228 ( .A(n68134), .B(n72971), .Z(n72966) );
  XOR U88229 ( .A(n72967), .B(n72966), .Z(n71738) );
  XOR U88230 ( .A(n68135), .B(n71738), .Z(n71732) );
  NOR U88231 ( .A(n68137), .B(n68136), .Z(n68143) );
  IV U88232 ( .A(n68138), .Z(n68140) );
  NOR U88233 ( .A(n68140), .B(n68139), .Z(n68141) );
  IV U88234 ( .A(n68141), .Z(n68142) );
  NOR U88235 ( .A(n68143), .B(n68142), .Z(n68144) );
  IV U88236 ( .A(n68144), .Z(n71733) );
  XOR U88237 ( .A(n71732), .B(n71733), .Z(n72977) );
  XOR U88238 ( .A(n72975), .B(n72977), .Z(n72980) );
  XOR U88239 ( .A(n72978), .B(n72980), .Z(n71727) );
  XOR U88240 ( .A(n71725), .B(n71727), .Z(n71729) );
  NOR U88241 ( .A(n68150), .B(n71729), .Z(n78494) );
  IV U88242 ( .A(n68145), .Z(n68146) );
  NOR U88243 ( .A(n68146), .B(n68156), .Z(n72983) );
  IV U88244 ( .A(n68147), .Z(n68148) );
  NOR U88245 ( .A(n68149), .B(n68148), .Z(n71728) );
  XOR U88246 ( .A(n71728), .B(n71729), .Z(n72984) );
  IV U88247 ( .A(n72984), .Z(n68151) );
  XOR U88248 ( .A(n72983), .B(n68151), .Z(n68153) );
  NOR U88249 ( .A(n68151), .B(n68150), .Z(n68152) );
  NOR U88250 ( .A(n68153), .B(n68152), .Z(n68154) );
  NOR U88251 ( .A(n78494), .B(n68154), .Z(n71722) );
  IV U88252 ( .A(n68155), .Z(n68157) );
  NOR U88253 ( .A(n68157), .B(n68156), .Z(n72986) );
  IV U88254 ( .A(n68158), .Z(n68162) );
  NOR U88255 ( .A(n68160), .B(n68159), .Z(n68161) );
  IV U88256 ( .A(n68161), .Z(n68165) );
  NOR U88257 ( .A(n68162), .B(n68165), .Z(n71723) );
  NOR U88258 ( .A(n72986), .B(n71723), .Z(n68163) );
  XOR U88259 ( .A(n71722), .B(n68163), .Z(n73002) );
  IV U88260 ( .A(n68164), .Z(n68166) );
  NOR U88261 ( .A(n68166), .B(n68165), .Z(n73000) );
  XOR U88262 ( .A(n73002), .B(n73000), .Z(n73007) );
  XOR U88263 ( .A(n68167), .B(n73007), .Z(n71716) );
  XOR U88264 ( .A(n71717), .B(n71716), .Z(n71720) );
  IV U88265 ( .A(n68168), .Z(n68169) );
  NOR U88266 ( .A(n68170), .B(n68169), .Z(n71719) );
  IV U88267 ( .A(n68171), .Z(n68172) );
  NOR U88268 ( .A(n68172), .B(n68176), .Z(n71713) );
  NOR U88269 ( .A(n71719), .B(n71713), .Z(n68173) );
  XOR U88270 ( .A(n71720), .B(n68173), .Z(n68174) );
  IV U88271 ( .A(n68174), .Z(n73020) );
  IV U88272 ( .A(n68175), .Z(n68177) );
  NOR U88273 ( .A(n68177), .B(n68176), .Z(n73018) );
  XOR U88274 ( .A(n73020), .B(n73018), .Z(n71712) );
  XOR U88275 ( .A(n71710), .B(n71712), .Z(n73015) );
  XOR U88276 ( .A(n73014), .B(n73015), .Z(n73012) );
  XOR U88277 ( .A(n73011), .B(n73012), .Z(n73028) );
  XOR U88278 ( .A(n68178), .B(n73028), .Z(n71706) );
  IV U88279 ( .A(n68179), .Z(n68180) );
  NOR U88280 ( .A(n68181), .B(n68180), .Z(n73029) );
  IV U88281 ( .A(n68182), .Z(n68183) );
  NOR U88282 ( .A(n68184), .B(n68183), .Z(n71705) );
  NOR U88283 ( .A(n73029), .B(n71705), .Z(n68185) );
  XOR U88284 ( .A(n71706), .B(n68185), .Z(n77173) );
  XOR U88285 ( .A(n71700), .B(n77173), .Z(n71701) );
  IV U88286 ( .A(n68186), .Z(n68188) );
  NOR U88287 ( .A(n68188), .B(n68187), .Z(n68189) );
  IV U88288 ( .A(n68189), .Z(n71702) );
  XOR U88289 ( .A(n71701), .B(n71702), .Z(n71698) );
  XOR U88290 ( .A(n71697), .B(n71698), .Z(n73037) );
  XOR U88291 ( .A(n73036), .B(n73037), .Z(n73040) );
  XOR U88292 ( .A(n73039), .B(n73040), .Z(n73044) );
  XOR U88293 ( .A(n73043), .B(n73044), .Z(n73048) );
  IV U88294 ( .A(n68190), .Z(n68192) );
  NOR U88295 ( .A(n68192), .B(n68191), .Z(n73046) );
  XOR U88296 ( .A(n73048), .B(n73046), .Z(n71695) );
  XOR U88297 ( .A(n71694), .B(n71695), .Z(n73056) );
  IV U88298 ( .A(n73056), .Z(n68197) );
  IV U88299 ( .A(n68193), .Z(n68194) );
  NOR U88300 ( .A(n68195), .B(n68194), .Z(n71692) );
  NOR U88301 ( .A(n73055), .B(n71692), .Z(n68196) );
  XOR U88302 ( .A(n68197), .B(n68196), .Z(n73061) );
  XOR U88303 ( .A(n73059), .B(n73061), .Z(n78566) );
  XOR U88304 ( .A(n68198), .B(n78566), .Z(n73067) );
  XOR U88305 ( .A(n73069), .B(n73067), .Z(n71690) );
  XOR U88306 ( .A(n71688), .B(n71690), .Z(n71684) );
  XOR U88307 ( .A(n71682), .B(n71684), .Z(n71687) );
  XOR U88308 ( .A(n68199), .B(n71687), .Z(n71670) );
  IV U88309 ( .A(n68200), .Z(n68201) );
  NOR U88310 ( .A(n68202), .B(n68201), .Z(n71671) );
  NOR U88311 ( .A(n71676), .B(n71671), .Z(n68203) );
  XOR U88312 ( .A(n71670), .B(n68203), .Z(n71675) );
  XOR U88313 ( .A(n71673), .B(n71675), .Z(n78576) );
  XOR U88314 ( .A(n71669), .B(n78576), .Z(n73083) );
  IV U88315 ( .A(n68204), .Z(n68206) );
  NOR U88316 ( .A(n68206), .B(n68205), .Z(n73082) );
  IV U88317 ( .A(n68207), .Z(n68209) );
  NOR U88318 ( .A(n68209), .B(n68208), .Z(n73085) );
  NOR U88319 ( .A(n73082), .B(n73085), .Z(n68210) );
  XOR U88320 ( .A(n73083), .B(n68210), .Z(n73078) );
  XOR U88321 ( .A(n73077), .B(n73078), .Z(n73094) );
  XOR U88322 ( .A(n68211), .B(n73094), .Z(n71663) );
  XOR U88323 ( .A(n71664), .B(n71663), .Z(n73107) );
  XOR U88324 ( .A(n68212), .B(n73107), .Z(n71653) );
  XOR U88325 ( .A(n68213), .B(n71653), .Z(n73109) );
  XOR U88326 ( .A(n73108), .B(n73109), .Z(n73112) );
  XOR U88327 ( .A(n73111), .B(n73112), .Z(n73118) );
  IV U88328 ( .A(n68214), .Z(n68216) );
  NOR U88329 ( .A(n68216), .B(n68215), .Z(n73115) );
  IV U88330 ( .A(n68217), .Z(n68219) );
  NOR U88331 ( .A(n68219), .B(n68218), .Z(n73117) );
  NOR U88332 ( .A(n73115), .B(n73117), .Z(n68220) );
  XOR U88333 ( .A(n73118), .B(n68220), .Z(n68221) );
  NOR U88334 ( .A(n68222), .B(n68221), .Z(n68225) );
  IV U88335 ( .A(n68222), .Z(n68224) );
  XOR U88336 ( .A(n73115), .B(n73118), .Z(n68223) );
  NOR U88337 ( .A(n68224), .B(n68223), .Z(n77108) );
  NOR U88338 ( .A(n68225), .B(n77108), .Z(n71650) );
  XOR U88339 ( .A(n71652), .B(n71650), .Z(n71648) );
  XOR U88340 ( .A(n68226), .B(n71648), .Z(n68227) );
  IV U88341 ( .A(n68227), .Z(n73125) );
  IV U88342 ( .A(n68228), .Z(n68230) );
  NOR U88343 ( .A(n68230), .B(n68229), .Z(n73123) );
  XOR U88344 ( .A(n73125), .B(n73123), .Z(n73127) );
  IV U88345 ( .A(n73127), .Z(n68237) );
  IV U88346 ( .A(n68231), .Z(n68235) );
  NOR U88347 ( .A(n68235), .B(n68232), .Z(n73126) );
  IV U88348 ( .A(n68233), .Z(n68234) );
  NOR U88349 ( .A(n68235), .B(n68234), .Z(n71642) );
  NOR U88350 ( .A(n73126), .B(n71642), .Z(n68236) );
  XOR U88351 ( .A(n68237), .B(n68236), .Z(n73132) );
  XOR U88352 ( .A(n73130), .B(n73132), .Z(n73134) );
  NOR U88353 ( .A(n68243), .B(n73134), .Z(n77084) );
  IV U88354 ( .A(n68238), .Z(n68240) );
  NOR U88355 ( .A(n68240), .B(n68239), .Z(n73133) );
  XOR U88356 ( .A(n73133), .B(n73134), .Z(n71641) );
  IV U88357 ( .A(n68241), .Z(n68242) );
  NOR U88358 ( .A(n68242), .B(n68252), .Z(n68244) );
  IV U88359 ( .A(n68244), .Z(n71640) );
  XOR U88360 ( .A(n71641), .B(n71640), .Z(n68246) );
  NOR U88361 ( .A(n68244), .B(n68243), .Z(n68245) );
  NOR U88362 ( .A(n68246), .B(n68245), .Z(n68247) );
  NOR U88363 ( .A(n77084), .B(n68247), .Z(n73138) );
  IV U88364 ( .A(n68248), .Z(n68250) );
  NOR U88365 ( .A(n68250), .B(n68249), .Z(n73137) );
  IV U88366 ( .A(n68251), .Z(n68253) );
  NOR U88367 ( .A(n68253), .B(n68252), .Z(n73142) );
  NOR U88368 ( .A(n73137), .B(n73142), .Z(n68254) );
  XOR U88369 ( .A(n73138), .B(n68254), .Z(n73156) );
  XOR U88370 ( .A(n73154), .B(n73156), .Z(n73159) );
  XOR U88371 ( .A(n73157), .B(n73159), .Z(n71638) );
  XOR U88372 ( .A(n68255), .B(n71638), .Z(n71629) );
  IV U88373 ( .A(n68256), .Z(n68258) );
  NOR U88374 ( .A(n68258), .B(n68257), .Z(n71634) );
  IV U88375 ( .A(n68259), .Z(n68261) );
  NOR U88376 ( .A(n68261), .B(n68260), .Z(n71630) );
  NOR U88377 ( .A(n71634), .B(n71630), .Z(n68262) );
  XOR U88378 ( .A(n71629), .B(n68262), .Z(n73164) );
  XOR U88379 ( .A(n68263), .B(n73164), .Z(n73167) );
  IV U88380 ( .A(n68264), .Z(n68265) );
  NOR U88381 ( .A(n68266), .B(n68265), .Z(n73166) );
  IV U88382 ( .A(n68267), .Z(n68269) );
  NOR U88383 ( .A(n68269), .B(n68268), .Z(n73183) );
  NOR U88384 ( .A(n73166), .B(n73183), .Z(n68270) );
  XOR U88385 ( .A(n73167), .B(n68270), .Z(n73182) );
  IV U88386 ( .A(n68271), .Z(n68273) );
  NOR U88387 ( .A(n68273), .B(n68272), .Z(n73180) );
  XOR U88388 ( .A(n73182), .B(n73180), .Z(n71625) );
  XOR U88389 ( .A(n71622), .B(n71625), .Z(n73191) );
  XOR U88390 ( .A(n68274), .B(n73191), .Z(n73194) );
  XOR U88391 ( .A(n73192), .B(n73194), .Z(n73197) );
  XOR U88392 ( .A(n68276), .B(n68275), .Z(n68280) );
  IV U88393 ( .A(n68277), .Z(n68289) );
  NOR U88394 ( .A(n68289), .B(n68278), .Z(n68279) );
  IV U88395 ( .A(n68279), .Z(n68285) );
  NOR U88396 ( .A(n68280), .B(n68285), .Z(n68281) );
  IV U88397 ( .A(n68281), .Z(n68282) );
  NOR U88398 ( .A(n68283), .B(n68282), .Z(n73195) );
  XOR U88399 ( .A(n73197), .B(n73195), .Z(n71621) );
  IV U88400 ( .A(n68284), .Z(n68286) );
  NOR U88401 ( .A(n68286), .B(n68285), .Z(n71619) );
  XOR U88402 ( .A(n71621), .B(n71619), .Z(n71616) );
  IV U88403 ( .A(n68287), .Z(n68288) );
  NOR U88404 ( .A(n68289), .B(n68288), .Z(n71614) );
  XOR U88405 ( .A(n71616), .B(n71614), .Z(n71617) );
  XOR U88406 ( .A(n71618), .B(n71617), .Z(n71612) );
  IV U88407 ( .A(n68290), .Z(n68291) );
  NOR U88408 ( .A(n68292), .B(n68291), .Z(n71611) );
  IV U88409 ( .A(n68293), .Z(n68297) );
  NOR U88410 ( .A(n68295), .B(n68294), .Z(n68296) );
  IV U88411 ( .A(n68296), .Z(n68300) );
  NOR U88412 ( .A(n68297), .B(n68300), .Z(n73204) );
  NOR U88413 ( .A(n71611), .B(n73204), .Z(n68298) );
  XOR U88414 ( .A(n71612), .B(n68298), .Z(n73203) );
  IV U88415 ( .A(n68299), .Z(n68301) );
  NOR U88416 ( .A(n68301), .B(n68300), .Z(n73201) );
  XOR U88417 ( .A(n73203), .B(n73201), .Z(n73209) );
  XOR U88418 ( .A(n73208), .B(n73209), .Z(n73212) );
  XOR U88419 ( .A(n73211), .B(n73212), .Z(n73217) );
  XOR U88420 ( .A(n73215), .B(n73217), .Z(n73220) );
  XOR U88421 ( .A(n73218), .B(n73220), .Z(n71607) );
  XOR U88422 ( .A(n71605), .B(n71607), .Z(n71610) );
  XOR U88423 ( .A(n71608), .B(n71610), .Z(n73223) );
  XOR U88424 ( .A(n73222), .B(n73223), .Z(n73238) );
  XOR U88425 ( .A(n73232), .B(n73238), .Z(n73243) );
  XOR U88426 ( .A(n68302), .B(n73243), .Z(n71600) );
  XOR U88427 ( .A(n71601), .B(n71600), .Z(n71599) );
  IV U88428 ( .A(n71599), .Z(n68312) );
  IV U88429 ( .A(n68303), .Z(n68308) );
  IV U88430 ( .A(n68304), .Z(n68305) );
  NOR U88431 ( .A(n68308), .B(n68305), .Z(n71602) );
  IV U88432 ( .A(n68306), .Z(n68310) );
  NOR U88433 ( .A(n68308), .B(n68307), .Z(n68309) );
  IV U88434 ( .A(n68309), .Z(n68314) );
  NOR U88435 ( .A(n68310), .B(n68314), .Z(n71597) );
  NOR U88436 ( .A(n71602), .B(n71597), .Z(n68311) );
  XOR U88437 ( .A(n68312), .B(n68311), .Z(n71596) );
  IV U88438 ( .A(n68313), .Z(n68315) );
  NOR U88439 ( .A(n68315), .B(n68314), .Z(n71594) );
  XOR U88440 ( .A(n71596), .B(n71594), .Z(n71592) );
  XOR U88441 ( .A(n68316), .B(n71592), .Z(n71584) );
  XOR U88442 ( .A(n71585), .B(n71584), .Z(n73252) );
  IV U88443 ( .A(n68317), .Z(n68325) );
  NOR U88444 ( .A(n68325), .B(n68318), .Z(n71587) );
  IV U88445 ( .A(n68319), .Z(n68321) );
  NOR U88446 ( .A(n68321), .B(n68320), .Z(n73250) );
  NOR U88447 ( .A(n71587), .B(n73250), .Z(n68322) );
  XOR U88448 ( .A(n73252), .B(n68322), .Z(n73247) );
  IV U88449 ( .A(n68323), .Z(n68324) );
  NOR U88450 ( .A(n68325), .B(n68324), .Z(n68326) );
  IV U88451 ( .A(n68326), .Z(n73248) );
  XOR U88452 ( .A(n73247), .B(n73248), .Z(n71579) );
  XOR U88453 ( .A(n71577), .B(n71579), .Z(n71581) );
  NOR U88454 ( .A(n68333), .B(n71581), .Z(n76984) );
  IV U88455 ( .A(n68327), .Z(n68328) );
  NOR U88456 ( .A(n68329), .B(n68328), .Z(n71571) );
  IV U88457 ( .A(n68330), .Z(n68331) );
  NOR U88458 ( .A(n68332), .B(n68331), .Z(n71580) );
  XOR U88459 ( .A(n71580), .B(n71581), .Z(n71572) );
  IV U88460 ( .A(n71572), .Z(n68334) );
  XOR U88461 ( .A(n71571), .B(n68334), .Z(n68336) );
  NOR U88462 ( .A(n68334), .B(n68333), .Z(n68335) );
  NOR U88463 ( .A(n68336), .B(n68335), .Z(n68337) );
  NOR U88464 ( .A(n76984), .B(n68337), .Z(n71574) );
  XOR U88465 ( .A(n71576), .B(n71574), .Z(n71570) );
  IV U88466 ( .A(n68338), .Z(n68340) );
  IV U88467 ( .A(n68339), .Z(n68342) );
  NOR U88468 ( .A(n68340), .B(n68342), .Z(n71568) );
  XOR U88469 ( .A(n71570), .B(n71568), .Z(n71564) );
  IV U88470 ( .A(n68341), .Z(n68343) );
  NOR U88471 ( .A(n68343), .B(n68342), .Z(n71562) );
  XOR U88472 ( .A(n71564), .B(n71562), .Z(n71566) );
  XOR U88473 ( .A(n71565), .B(n71566), .Z(n71557) );
  XOR U88474 ( .A(n71556), .B(n71557), .Z(n71560) );
  XOR U88475 ( .A(n71559), .B(n71560), .Z(n71552) );
  IV U88476 ( .A(n68344), .Z(n68346) );
  NOR U88477 ( .A(n68346), .B(n68345), .Z(n71550) );
  XOR U88478 ( .A(n71552), .B(n71550), .Z(n71554) );
  XOR U88479 ( .A(n71553), .B(n71554), .Z(n73260) );
  NOR U88480 ( .A(n68347), .B(n73260), .Z(n76956) );
  IV U88481 ( .A(n68348), .Z(n68352) );
  XOR U88482 ( .A(n68350), .B(n68349), .Z(n68351) );
  NOR U88483 ( .A(n68352), .B(n68351), .Z(n68362) );
  IV U88484 ( .A(n68362), .Z(n68356) );
  IV U88485 ( .A(n68353), .Z(n68354) );
  NOR U88486 ( .A(n68355), .B(n68354), .Z(n73259) );
  XOR U88487 ( .A(n73259), .B(n73260), .Z(n73269) );
  NOR U88488 ( .A(n68356), .B(n73269), .Z(n78668) );
  NOR U88489 ( .A(n76956), .B(n78668), .Z(n73263) );
  IV U88490 ( .A(n73263), .Z(n68357) );
  NOR U88491 ( .A(n73268), .B(n68357), .Z(n68358) );
  IV U88492 ( .A(n68358), .Z(n68361) );
  IV U88493 ( .A(n73269), .Z(n68364) );
  NOR U88494 ( .A(n68359), .B(n68364), .Z(n68360) );
  NOR U88495 ( .A(n68361), .B(n68360), .Z(n68366) );
  NOR U88496 ( .A(n73268), .B(n68362), .Z(n68363) );
  NOR U88497 ( .A(n68364), .B(n68363), .Z(n68365) );
  NOR U88498 ( .A(n68366), .B(n68365), .Z(n73267) );
  XOR U88499 ( .A(n68367), .B(n73267), .Z(n73272) );
  XOR U88500 ( .A(n73274), .B(n73272), .Z(n76945) );
  XOR U88501 ( .A(n68368), .B(n76945), .Z(n73284) );
  IV U88502 ( .A(n68369), .Z(n68371) );
  NOR U88503 ( .A(n68371), .B(n68370), .Z(n73282) );
  XOR U88504 ( .A(n73284), .B(n73282), .Z(n73279) );
  XOR U88505 ( .A(n73280), .B(n73279), .Z(n73294) );
  IV U88506 ( .A(n68372), .Z(n68373) );
  NOR U88507 ( .A(n68374), .B(n68373), .Z(n84467) );
  IV U88508 ( .A(n68375), .Z(n68377) );
  NOR U88509 ( .A(n68377), .B(n68376), .Z(n82643) );
  NOR U88510 ( .A(n84467), .B(n82643), .Z(n73295) );
  XOR U88511 ( .A(n73294), .B(n73295), .Z(n71545) );
  XOR U88512 ( .A(n71544), .B(n71545), .Z(n73292) );
  XOR U88513 ( .A(n73290), .B(n73292), .Z(n73303) );
  XOR U88514 ( .A(n73301), .B(n73303), .Z(n73305) );
  XOR U88515 ( .A(n73304), .B(n73305), .Z(n71540) );
  XOR U88516 ( .A(n71538), .B(n71540), .Z(n71543) );
  XOR U88517 ( .A(n71541), .B(n71543), .Z(n71534) );
  XOR U88518 ( .A(n71532), .B(n71534), .Z(n71537) );
  XOR U88519 ( .A(n71535), .B(n71537), .Z(n71527) );
  XOR U88520 ( .A(n71526), .B(n71527), .Z(n71530) );
  XOR U88521 ( .A(n71529), .B(n71530), .Z(n76929) );
  XOR U88522 ( .A(n68378), .B(n76929), .Z(n76921) );
  IV U88523 ( .A(n68379), .Z(n68389) );
  IV U88524 ( .A(n68380), .Z(n68381) );
  NOR U88525 ( .A(n68389), .B(n68381), .Z(n76920) );
  IV U88526 ( .A(n68382), .Z(n68384) );
  NOR U88527 ( .A(n68384), .B(n68383), .Z(n76924) );
  NOR U88528 ( .A(n76920), .B(n76924), .Z(n71522) );
  IV U88529 ( .A(n71522), .Z(n68390) );
  XOR U88530 ( .A(n76921), .B(n68390), .Z(n68385) );
  NOR U88531 ( .A(n68386), .B(n68385), .Z(n76915) );
  IV U88532 ( .A(n68387), .Z(n68388) );
  NOR U88533 ( .A(n68389), .B(n68388), .Z(n71519) );
  NOR U88534 ( .A(n71519), .B(n68390), .Z(n68391) );
  XOR U88535 ( .A(n76921), .B(n68391), .Z(n68392) );
  NOR U88536 ( .A(n68393), .B(n68392), .Z(n68394) );
  NOR U88537 ( .A(n76915), .B(n68394), .Z(n73311) );
  XOR U88538 ( .A(n73312), .B(n73311), .Z(n73314) );
  XOR U88539 ( .A(n68395), .B(n73314), .Z(n73318) );
  XOR U88540 ( .A(n73319), .B(n73318), .Z(n73324) );
  IV U88541 ( .A(n68396), .Z(n68397) );
  NOR U88542 ( .A(n68398), .B(n68397), .Z(n73322) );
  XOR U88543 ( .A(n73324), .B(n73322), .Z(n73334) );
  XOR U88544 ( .A(n73333), .B(n73334), .Z(n73337) );
  XOR U88545 ( .A(n73336), .B(n73337), .Z(n71517) );
  XOR U88546 ( .A(n71516), .B(n71517), .Z(n73343) );
  XOR U88547 ( .A(n73342), .B(n73343), .Z(n71514) );
  XOR U88548 ( .A(n71513), .B(n71514), .Z(n71509) );
  IV U88549 ( .A(n68399), .Z(n68402) );
  IV U88550 ( .A(n68400), .Z(n68401) );
  NOR U88551 ( .A(n68402), .B(n68401), .Z(n71507) );
  XOR U88552 ( .A(n71509), .B(n71507), .Z(n71511) );
  IV U88553 ( .A(n68403), .Z(n68404) );
  NOR U88554 ( .A(n68405), .B(n68404), .Z(n71510) );
  IV U88555 ( .A(n68406), .Z(n68407) );
  NOR U88556 ( .A(n68410), .B(n68407), .Z(n71505) );
  NOR U88557 ( .A(n71510), .B(n71505), .Z(n68408) );
  XOR U88558 ( .A(n71511), .B(n68408), .Z(n73349) );
  IV U88559 ( .A(n68409), .Z(n68411) );
  NOR U88560 ( .A(n68411), .B(n68410), .Z(n73350) );
  IV U88561 ( .A(n68412), .Z(n68414) );
  NOR U88562 ( .A(n68414), .B(n68413), .Z(n73352) );
  NOR U88563 ( .A(n73350), .B(n73352), .Z(n68415) );
  XOR U88564 ( .A(n73349), .B(n68415), .Z(n73357) );
  XOR U88565 ( .A(n68416), .B(n73357), .Z(n73358) );
  IV U88566 ( .A(n68417), .Z(n68418) );
  NOR U88567 ( .A(n68425), .B(n68418), .Z(n73363) );
  IV U88568 ( .A(n68419), .Z(n68420) );
  NOR U88569 ( .A(n68421), .B(n68420), .Z(n73359) );
  NOR U88570 ( .A(n73363), .B(n73359), .Z(n68422) );
  XOR U88571 ( .A(n73358), .B(n68422), .Z(n71499) );
  IV U88572 ( .A(n68423), .Z(n68424) );
  NOR U88573 ( .A(n68425), .B(n68424), .Z(n71497) );
  XOR U88574 ( .A(n71499), .B(n71497), .Z(n71501) );
  XOR U88575 ( .A(n71500), .B(n71501), .Z(n71495) );
  NOR U88576 ( .A(n68432), .B(n71495), .Z(n78769) );
  IV U88577 ( .A(n68426), .Z(n68427) );
  NOR U88578 ( .A(n68428), .B(n68427), .Z(n71487) );
  IV U88579 ( .A(n68429), .Z(n68431) );
  NOR U88580 ( .A(n68431), .B(n68430), .Z(n71494) );
  XOR U88581 ( .A(n71494), .B(n71495), .Z(n71488) );
  IV U88582 ( .A(n71488), .Z(n68433) );
  XOR U88583 ( .A(n71487), .B(n68433), .Z(n68435) );
  NOR U88584 ( .A(n68433), .B(n68432), .Z(n68434) );
  NOR U88585 ( .A(n68435), .B(n68434), .Z(n68436) );
  NOR U88586 ( .A(n78769), .B(n68436), .Z(n68437) );
  IV U88587 ( .A(n68437), .Z(n71491) );
  XOR U88588 ( .A(n71491), .B(n71490), .Z(n73371) );
  XOR U88589 ( .A(n68438), .B(n73371), .Z(n73372) );
  XOR U88590 ( .A(n73373), .B(n73372), .Z(n73376) );
  XOR U88591 ( .A(n73375), .B(n73376), .Z(n68439) );
  XOR U88592 ( .A(n68440), .B(n68439), .Z(n71478) );
  IV U88593 ( .A(n68441), .Z(n68443) );
  NOR U88594 ( .A(n68443), .B(n68442), .Z(n78783) );
  NOR U88595 ( .A(n68445), .B(n68444), .Z(n76860) );
  NOR U88596 ( .A(n78783), .B(n76860), .Z(n71479) );
  XOR U88597 ( .A(n71478), .B(n71479), .Z(n71473) );
  XOR U88598 ( .A(n71474), .B(n71473), .Z(n71471) );
  IV U88599 ( .A(n68446), .Z(n68448) );
  NOR U88600 ( .A(n68448), .B(n68447), .Z(n71475) );
  IV U88601 ( .A(n68449), .Z(n68451) );
  NOR U88602 ( .A(n68451), .B(n68450), .Z(n71470) );
  NOR U88603 ( .A(n71475), .B(n71470), .Z(n68452) );
  XOR U88604 ( .A(n71471), .B(n68452), .Z(n71469) );
  XOR U88605 ( .A(n71467), .B(n71469), .Z(n73382) );
  XOR U88606 ( .A(n73381), .B(n73382), .Z(n73386) );
  XOR U88607 ( .A(n73384), .B(n73386), .Z(n73390) );
  XOR U88608 ( .A(n73388), .B(n73390), .Z(n73392) );
  XOR U88609 ( .A(n73391), .B(n73392), .Z(n73396) );
  XOR U88610 ( .A(n73395), .B(n73396), .Z(n73400) );
  XOR U88611 ( .A(n73398), .B(n73400), .Z(n73404) );
  XOR U88612 ( .A(n73402), .B(n73404), .Z(n73409) );
  XOR U88613 ( .A(n68453), .B(n73409), .Z(n73411) );
  XOR U88614 ( .A(n73412), .B(n73411), .Z(n73418) );
  IV U88615 ( .A(n68454), .Z(n68455) );
  NOR U88616 ( .A(n68456), .B(n68455), .Z(n73414) );
  IV U88617 ( .A(n68457), .Z(n68459) );
  NOR U88618 ( .A(n68459), .B(n68458), .Z(n73417) );
  NOR U88619 ( .A(n73414), .B(n73417), .Z(n68460) );
  XOR U88620 ( .A(n73418), .B(n68460), .Z(n73421) );
  XOR U88621 ( .A(n68461), .B(n73421), .Z(n73427) );
  IV U88622 ( .A(n68462), .Z(n71461) );
  NOR U88623 ( .A(n71461), .B(n68463), .Z(n68467) );
  IV U88624 ( .A(n68464), .Z(n68466) );
  NOR U88625 ( .A(n68466), .B(n68465), .Z(n73426) );
  NOR U88626 ( .A(n68467), .B(n73426), .Z(n68468) );
  XOR U88627 ( .A(n73427), .B(n68468), .Z(n71457) );
  IV U88628 ( .A(n68469), .Z(n68470) );
  NOR U88629 ( .A(n68471), .B(n68470), .Z(n71458) );
  IV U88630 ( .A(n68472), .Z(n68473) );
  NOR U88631 ( .A(n68474), .B(n68473), .Z(n73433) );
  NOR U88632 ( .A(n71458), .B(n73433), .Z(n68475) );
  XOR U88633 ( .A(n71457), .B(n68475), .Z(n73431) );
  XOR U88634 ( .A(n73430), .B(n73431), .Z(n71452) );
  XOR U88635 ( .A(n71451), .B(n71452), .Z(n71456) );
  IV U88636 ( .A(n68476), .Z(n68479) );
  IV U88637 ( .A(n68477), .Z(n68478) );
  NOR U88638 ( .A(n68479), .B(n68478), .Z(n71454) );
  XOR U88639 ( .A(n71456), .B(n71454), .Z(n71449) );
  IV U88640 ( .A(n68480), .Z(n68481) );
  NOR U88641 ( .A(n68482), .B(n68481), .Z(n71447) );
  XOR U88642 ( .A(n71449), .B(n71447), .Z(n73439) );
  XOR U88643 ( .A(n73438), .B(n73439), .Z(n73442) );
  XOR U88644 ( .A(n73441), .B(n73442), .Z(n73447) );
  IV U88645 ( .A(n68483), .Z(n68489) );
  IV U88646 ( .A(n68484), .Z(n68486) );
  NOR U88647 ( .A(n68486), .B(n68485), .Z(n68487) );
  IV U88648 ( .A(n68487), .Z(n68488) );
  NOR U88649 ( .A(n68489), .B(n68488), .Z(n73445) );
  XOR U88650 ( .A(n73447), .B(n73445), .Z(n73449) );
  XOR U88651 ( .A(n73448), .B(n73449), .Z(n71442) );
  XOR U88652 ( .A(n71441), .B(n71442), .Z(n71445) );
  XOR U88653 ( .A(n71444), .B(n71445), .Z(n71437) );
  IV U88654 ( .A(n68490), .Z(n68495) );
  IV U88655 ( .A(n68491), .Z(n68492) );
  NOR U88656 ( .A(n68493), .B(n68492), .Z(n68494) );
  IV U88657 ( .A(n68494), .Z(n68497) );
  NOR U88658 ( .A(n68495), .B(n68497), .Z(n71435) );
  XOR U88659 ( .A(n71437), .B(n71435), .Z(n71440) );
  IV U88660 ( .A(n68496), .Z(n68498) );
  NOR U88661 ( .A(n68498), .B(n68497), .Z(n71438) );
  XOR U88662 ( .A(n71440), .B(n71438), .Z(n71429) );
  IV U88663 ( .A(n68499), .Z(n68502) );
  IV U88664 ( .A(n68500), .Z(n68501) );
  NOR U88665 ( .A(n68502), .B(n68501), .Z(n71427) );
  XOR U88666 ( .A(n71429), .B(n71427), .Z(n71431) );
  IV U88667 ( .A(n71431), .Z(n68506) );
  XOR U88668 ( .A(n71430), .B(n68506), .Z(n68503) );
  NOR U88669 ( .A(n68504), .B(n68503), .Z(n68516) );
  IV U88670 ( .A(n68505), .Z(n68510) );
  NOR U88671 ( .A(n71430), .B(n68506), .Z(n68508) );
  NOR U88672 ( .A(n68508), .B(n68507), .Z(n68509) );
  IV U88673 ( .A(n68509), .Z(n68512) );
  NOR U88674 ( .A(n68510), .B(n68512), .Z(n78849) );
  IV U88675 ( .A(n68511), .Z(n68513) );
  NOR U88676 ( .A(n68513), .B(n68512), .Z(n71426) );
  NOR U88677 ( .A(n78849), .B(n71426), .Z(n68514) );
  IV U88678 ( .A(n68514), .Z(n68515) );
  NOR U88679 ( .A(n68516), .B(n68515), .Z(n71420) );
  XOR U88680 ( .A(n68517), .B(n71420), .Z(n71414) );
  XOR U88681 ( .A(n68518), .B(n71414), .Z(n73459) );
  XOR U88682 ( .A(n68519), .B(n73459), .Z(n73465) );
  XOR U88683 ( .A(n76787), .B(n73465), .Z(n73467) );
  XOR U88684 ( .A(n68520), .B(n73467), .Z(n68521) );
  IV U88685 ( .A(n68521), .Z(n71406) );
  XOR U88686 ( .A(n71404), .B(n71406), .Z(n71409) );
  IV U88687 ( .A(n68522), .Z(n68524) );
  NOR U88688 ( .A(n68524), .B(n68523), .Z(n71407) );
  XOR U88689 ( .A(n71409), .B(n71407), .Z(n71399) );
  XOR U88690 ( .A(n71398), .B(n71399), .Z(n71402) );
  IV U88691 ( .A(n68525), .Z(n68527) );
  NOR U88692 ( .A(n68527), .B(n68526), .Z(n71401) );
  IV U88693 ( .A(n68528), .Z(n68530) );
  NOR U88694 ( .A(n68530), .B(n68529), .Z(n71396) );
  NOR U88695 ( .A(n71401), .B(n71396), .Z(n68531) );
  XOR U88696 ( .A(n71402), .B(n68531), .Z(n68532) );
  IV U88697 ( .A(n68532), .Z(n71395) );
  XOR U88698 ( .A(n71393), .B(n71395), .Z(n68538) );
  NOR U88699 ( .A(n68540), .B(n68538), .Z(n78907) );
  IV U88700 ( .A(n68533), .Z(n68534) );
  NOR U88701 ( .A(n68535), .B(n68534), .Z(n73477) );
  IV U88702 ( .A(n68536), .Z(n71387) );
  NOR U88703 ( .A(n68537), .B(n71387), .Z(n68539) );
  XOR U88704 ( .A(n68539), .B(n68538), .Z(n73478) );
  IV U88705 ( .A(n73478), .Z(n68541) );
  XOR U88706 ( .A(n73477), .B(n68541), .Z(n68543) );
  NOR U88707 ( .A(n68541), .B(n68540), .Z(n68542) );
  NOR U88708 ( .A(n68543), .B(n68542), .Z(n68544) );
  NOR U88709 ( .A(n78907), .B(n68544), .Z(n71382) );
  XOR U88710 ( .A(n71384), .B(n71382), .Z(n71377) );
  XOR U88711 ( .A(n68545), .B(n71377), .Z(n68546) );
  XOR U88712 ( .A(n68547), .B(n68546), .Z(n71365) );
  XOR U88713 ( .A(n71364), .B(n71365), .Z(n71362) );
  XOR U88714 ( .A(n71361), .B(n71362), .Z(n73489) );
  NOR U88715 ( .A(n68552), .B(n73489), .Z(n76752) );
  IV U88716 ( .A(n68548), .Z(n68551) );
  IV U88717 ( .A(n68549), .Z(n68550) );
  NOR U88718 ( .A(n68551), .B(n68550), .Z(n73491) );
  XOR U88719 ( .A(n73488), .B(n73489), .Z(n73492) );
  IV U88720 ( .A(n73492), .Z(n68553) );
  XOR U88721 ( .A(n73491), .B(n68553), .Z(n68555) );
  NOR U88722 ( .A(n68553), .B(n68552), .Z(n68554) );
  NOR U88723 ( .A(n68555), .B(n68554), .Z(n68556) );
  NOR U88724 ( .A(n76752), .B(n68556), .Z(n71346) );
  IV U88725 ( .A(n68557), .Z(n68559) );
  NOR U88726 ( .A(n68559), .B(n68558), .Z(n68562) );
  IV U88727 ( .A(n68560), .Z(n68561) );
  NOR U88728 ( .A(n68561), .B(n68565), .Z(n71345) );
  NOR U88729 ( .A(n68562), .B(n71345), .Z(n68563) );
  XOR U88730 ( .A(n71346), .B(n68563), .Z(n73499) );
  IV U88731 ( .A(n68564), .Z(n68566) );
  NOR U88732 ( .A(n68566), .B(n68565), .Z(n71343) );
  IV U88733 ( .A(n68567), .Z(n68569) );
  NOR U88734 ( .A(n68569), .B(n68568), .Z(n73497) );
  NOR U88735 ( .A(n71343), .B(n73497), .Z(n68570) );
  XOR U88736 ( .A(n73499), .B(n68570), .Z(n71341) );
  XOR U88737 ( .A(n68571), .B(n71341), .Z(n73505) );
  XOR U88738 ( .A(n68572), .B(n73505), .Z(n68573) );
  IV U88739 ( .A(n68573), .Z(n73519) );
  XOR U88740 ( .A(n73506), .B(n73519), .Z(n73510) );
  XOR U88741 ( .A(n73508), .B(n73510), .Z(n73514) );
  XOR U88742 ( .A(n68574), .B(n73514), .Z(n68575) );
  IV U88743 ( .A(n68575), .Z(n71334) );
  XOR U88744 ( .A(n71332), .B(n71334), .Z(n71336) );
  XOR U88745 ( .A(n71335), .B(n71336), .Z(n71330) );
  XOR U88746 ( .A(n71327), .B(n71330), .Z(n71325) );
  IV U88747 ( .A(n68576), .Z(n68578) );
  NOR U88748 ( .A(n68578), .B(n68577), .Z(n71329) );
  IV U88749 ( .A(n68579), .Z(n68580) );
  NOR U88750 ( .A(n68580), .B(n68583), .Z(n71323) );
  NOR U88751 ( .A(n71329), .B(n71323), .Z(n68581) );
  XOR U88752 ( .A(n71325), .B(n68581), .Z(n71317) );
  IV U88753 ( .A(n68582), .Z(n68584) );
  NOR U88754 ( .A(n68584), .B(n68583), .Z(n68585) );
  IV U88755 ( .A(n68585), .Z(n71318) );
  XOR U88756 ( .A(n71317), .B(n71318), .Z(n71322) );
  XOR U88757 ( .A(n71320), .B(n71322), .Z(n71315) );
  XOR U88758 ( .A(n71313), .B(n71315), .Z(n73530) );
  XOR U88759 ( .A(n73529), .B(n73530), .Z(n73542) );
  XOR U88760 ( .A(n68586), .B(n73542), .Z(n73536) );
  NOR U88761 ( .A(n73545), .B(n68587), .Z(n68591) );
  IV U88762 ( .A(n68588), .Z(n68590) );
  NOR U88763 ( .A(n68590), .B(n68589), .Z(n73537) );
  NOR U88764 ( .A(n68591), .B(n73537), .Z(n68592) );
  XOR U88765 ( .A(n73536), .B(n68592), .Z(n73550) );
  XOR U88766 ( .A(n73548), .B(n73550), .Z(n71311) );
  XOR U88767 ( .A(n71310), .B(n71311), .Z(n71306) );
  XOR U88768 ( .A(n71304), .B(n71306), .Z(n71309) );
  XOR U88769 ( .A(n71307), .B(n71309), .Z(n76696) );
  XOR U88770 ( .A(n71299), .B(n76696), .Z(n71296) );
  IV U88771 ( .A(n68593), .Z(n68595) );
  NOR U88772 ( .A(n68595), .B(n68594), .Z(n71300) );
  IV U88773 ( .A(n68596), .Z(n68598) );
  NOR U88774 ( .A(n68598), .B(n68597), .Z(n71297) );
  NOR U88775 ( .A(n71300), .B(n71297), .Z(n68599) );
  XOR U88776 ( .A(n71296), .B(n68599), .Z(n73562) );
  IV U88777 ( .A(n68600), .Z(n68602) );
  NOR U88778 ( .A(n68602), .B(n68601), .Z(n73560) );
  XOR U88779 ( .A(n73562), .B(n73560), .Z(n73568) );
  XOR U88780 ( .A(n71294), .B(n73568), .Z(n68603) );
  NOR U88781 ( .A(n68604), .B(n68603), .Z(n79000) );
  IV U88782 ( .A(n68605), .Z(n68606) );
  NOR U88783 ( .A(n68607), .B(n68606), .Z(n73567) );
  NOR U88784 ( .A(n73567), .B(n71294), .Z(n68608) );
  XOR U88785 ( .A(n68608), .B(n73568), .Z(n68616) );
  NOR U88786 ( .A(n68609), .B(n68616), .Z(n68610) );
  NOR U88787 ( .A(n79000), .B(n68610), .Z(n68623) );
  IV U88788 ( .A(n68623), .Z(n68611) );
  NOR U88789 ( .A(n68612), .B(n68611), .Z(n82317) );
  IV U88790 ( .A(n68613), .Z(n68615) );
  NOR U88791 ( .A(n68615), .B(n68614), .Z(n68620) );
  IV U88792 ( .A(n68620), .Z(n68618) );
  IV U88793 ( .A(n68616), .Z(n68617) );
  NOR U88794 ( .A(n68618), .B(n68617), .Z(n79003) );
  NOR U88795 ( .A(n68620), .B(n68619), .Z(n68621) );
  IV U88796 ( .A(n68621), .Z(n68622) );
  NOR U88797 ( .A(n68623), .B(n68622), .Z(n68624) );
  NOR U88798 ( .A(n79003), .B(n68624), .Z(n68625) );
  IV U88799 ( .A(n68625), .Z(n71291) );
  NOR U88800 ( .A(n82317), .B(n71291), .Z(n73573) );
  IV U88801 ( .A(n68626), .Z(n68628) );
  NOR U88802 ( .A(n68628), .B(n68627), .Z(n71290) );
  IV U88803 ( .A(n68629), .Z(n68630) );
  NOR U88804 ( .A(n68631), .B(n68630), .Z(n73572) );
  NOR U88805 ( .A(n71290), .B(n73572), .Z(n68632) );
  XOR U88806 ( .A(n73573), .B(n68632), .Z(n73577) );
  XOR U88807 ( .A(n73575), .B(n73577), .Z(n73579) );
  XOR U88808 ( .A(n73578), .B(n73579), .Z(n71288) );
  XOR U88809 ( .A(n71285), .B(n71288), .Z(n68633) );
  NOR U88810 ( .A(n68634), .B(n68633), .Z(n71284) );
  IV U88811 ( .A(n68635), .Z(n68637) );
  NOR U88812 ( .A(n68637), .B(n68636), .Z(n71287) );
  NOR U88813 ( .A(n71285), .B(n71287), .Z(n68638) );
  XOR U88814 ( .A(n71288), .B(n68638), .Z(n68639) );
  NOR U88815 ( .A(n68640), .B(n68639), .Z(n68641) );
  NOR U88816 ( .A(n71284), .B(n68641), .Z(n71278) );
  IV U88817 ( .A(n68642), .Z(n68644) );
  NOR U88818 ( .A(n68644), .B(n68643), .Z(n73587) );
  IV U88819 ( .A(n68645), .Z(n68647) );
  NOR U88820 ( .A(n68647), .B(n68646), .Z(n71280) );
  NOR U88821 ( .A(n73587), .B(n71280), .Z(n68648) );
  XOR U88822 ( .A(n71278), .B(n68648), .Z(n71275) );
  XOR U88823 ( .A(n71273), .B(n71275), .Z(n73598) );
  XOR U88824 ( .A(n68649), .B(n73598), .Z(n71270) );
  XOR U88825 ( .A(n68650), .B(n71270), .Z(n71266) );
  XOR U88826 ( .A(n71264), .B(n71266), .Z(n71268) );
  XOR U88827 ( .A(n71267), .B(n71268), .Z(n73603) );
  XOR U88828 ( .A(n73602), .B(n73603), .Z(n73608) );
  XOR U88829 ( .A(n68651), .B(n73608), .Z(n73612) );
  IV U88830 ( .A(n68652), .Z(n68653) );
  NOR U88831 ( .A(n68653), .B(n68656), .Z(n68654) );
  IV U88832 ( .A(n68654), .Z(n73613) );
  XOR U88833 ( .A(n73612), .B(n73613), .Z(n76638) );
  IV U88834 ( .A(n68655), .Z(n68657) );
  NOR U88835 ( .A(n68657), .B(n68656), .Z(n73615) );
  XOR U88836 ( .A(n76638), .B(n73615), .Z(n73624) );
  NOR U88837 ( .A(n76636), .B(n68658), .Z(n73619) );
  IV U88838 ( .A(n68659), .Z(n68661) );
  NOR U88839 ( .A(n68661), .B(n68660), .Z(n73623) );
  NOR U88840 ( .A(n73619), .B(n73623), .Z(n68662) );
  XOR U88841 ( .A(n73624), .B(n68662), .Z(n68663) );
  IV U88842 ( .A(n68663), .Z(n79022) );
  XOR U88843 ( .A(n73621), .B(n79022), .Z(n73628) );
  XOR U88844 ( .A(n73629), .B(n73628), .Z(n68664) );
  IV U88845 ( .A(n68664), .Z(n73631) );
  XOR U88846 ( .A(n73630), .B(n73631), .Z(n71262) );
  IV U88847 ( .A(n68665), .Z(n68667) );
  NOR U88848 ( .A(n68667), .B(n68666), .Z(n71261) );
  NOR U88849 ( .A(n68669), .B(n68668), .Z(n71256) );
  NOR U88850 ( .A(n71261), .B(n71256), .Z(n68670) );
  XOR U88851 ( .A(n71262), .B(n68670), .Z(n68671) );
  IV U88852 ( .A(n68671), .Z(n71259) );
  IV U88853 ( .A(n68677), .Z(n68672) );
  NOR U88854 ( .A(n68676), .B(n68672), .Z(n71254) );
  NOR U88855 ( .A(n71258), .B(n71254), .Z(n68673) );
  XOR U88856 ( .A(n71259), .B(n68673), .Z(n68674) );
  NOR U88857 ( .A(n68675), .B(n68674), .Z(n68683) );
  XOR U88858 ( .A(n68677), .B(n68676), .Z(n68679) );
  XOR U88859 ( .A(n71258), .B(n71259), .Z(n68678) );
  NOR U88860 ( .A(n68679), .B(n68678), .Z(n68680) );
  IV U88861 ( .A(n68680), .Z(n68681) );
  NOR U88862 ( .A(n68682), .B(n68681), .Z(n79036) );
  NOR U88863 ( .A(n68683), .B(n79036), .Z(n68684) );
  IV U88864 ( .A(n68684), .Z(n73641) );
  IV U88865 ( .A(n68685), .Z(n68686) );
  NOR U88866 ( .A(n68686), .B(n68689), .Z(n73639) );
  XOR U88867 ( .A(n73641), .B(n73639), .Z(n73644) );
  IV U88868 ( .A(n68696), .Z(n71248) );
  IV U88869 ( .A(n68687), .Z(n68697) );
  NOR U88870 ( .A(n71248), .B(n68697), .Z(n68691) );
  IV U88871 ( .A(n68688), .Z(n68690) );
  NOR U88872 ( .A(n68690), .B(n68689), .Z(n73643) );
  XOR U88873 ( .A(n68691), .B(n73643), .Z(n68692) );
  XOR U88874 ( .A(n73644), .B(n68692), .Z(n76611) );
  IV U88875 ( .A(n68693), .Z(n68694) );
  NOR U88876 ( .A(n71248), .B(n68694), .Z(n79050) );
  IV U88877 ( .A(n68695), .Z(n68699) );
  XOR U88878 ( .A(n68697), .B(n68696), .Z(n68698) );
  NOR U88879 ( .A(n68699), .B(n68698), .Z(n76609) );
  NOR U88880 ( .A(n79050), .B(n76609), .Z(n73650) );
  XOR U88881 ( .A(n76611), .B(n73650), .Z(n73651) );
  XOR U88882 ( .A(n73652), .B(n73651), .Z(n73658) );
  XOR U88883 ( .A(n73656), .B(n73658), .Z(n73661) );
  XOR U88884 ( .A(n68700), .B(n73661), .Z(n71239) );
  XOR U88885 ( .A(n68701), .B(n71239), .Z(n73664) );
  XOR U88886 ( .A(n73662), .B(n73664), .Z(n73666) );
  XOR U88887 ( .A(n73665), .B(n73666), .Z(n71237) );
  XOR U88888 ( .A(n68702), .B(n71237), .Z(n71227) );
  XOR U88889 ( .A(n71228), .B(n71227), .Z(n71232) );
  IV U88890 ( .A(n68703), .Z(n68704) );
  NOR U88891 ( .A(n68714), .B(n68704), .Z(n68705) );
  IV U88892 ( .A(n68705), .Z(n68706) );
  NOR U88893 ( .A(n68707), .B(n68706), .Z(n71225) );
  IV U88894 ( .A(n68708), .Z(n68710) );
  NOR U88895 ( .A(n68710), .B(n68709), .Z(n71230) );
  NOR U88896 ( .A(n71225), .B(n71230), .Z(n68711) );
  XOR U88897 ( .A(n71232), .B(n68711), .Z(n71222) );
  IV U88898 ( .A(n68712), .Z(n68713) );
  NOR U88899 ( .A(n68714), .B(n68713), .Z(n71223) );
  NOR U88900 ( .A(n73671), .B(n71223), .Z(n68715) );
  XOR U88901 ( .A(n71222), .B(n68715), .Z(n73675) );
  XOR U88902 ( .A(n73674), .B(n73675), .Z(n73680) );
  IV U88903 ( .A(n68716), .Z(n68718) );
  NOR U88904 ( .A(n68718), .B(n68717), .Z(n71220) );
  NOR U88905 ( .A(n73679), .B(n71220), .Z(n68719) );
  XOR U88906 ( .A(n73680), .B(n68719), .Z(n71209) );
  NOR U88907 ( .A(n68720), .B(n71213), .Z(n68723) );
  NOR U88908 ( .A(n68722), .B(n68721), .Z(n71210) );
  NOR U88909 ( .A(n68723), .B(n71210), .Z(n68724) );
  XOR U88910 ( .A(n71209), .B(n68724), .Z(n71207) );
  XOR U88911 ( .A(n71206), .B(n71207), .Z(n71204) );
  IV U88912 ( .A(n71204), .Z(n68729) );
  IV U88913 ( .A(n68725), .Z(n68727) );
  NOR U88914 ( .A(n68727), .B(n68726), .Z(n71201) );
  NOR U88915 ( .A(n71203), .B(n71201), .Z(n68728) );
  XOR U88916 ( .A(n68729), .B(n68728), .Z(n71199) );
  XOR U88917 ( .A(n71198), .B(n71199), .Z(n84893) );
  XOR U88918 ( .A(n73686), .B(n84893), .Z(n71195) );
  IV U88919 ( .A(n68730), .Z(n68731) );
  NOR U88920 ( .A(n68732), .B(n68731), .Z(n68733) );
  IV U88921 ( .A(n68733), .Z(n68734) );
  NOR U88922 ( .A(n68735), .B(n68734), .Z(n68736) );
  IV U88923 ( .A(n68736), .Z(n71196) );
  XOR U88924 ( .A(n71195), .B(n71196), .Z(n73701) );
  XOR U88925 ( .A(n73700), .B(n73701), .Z(n71193) );
  IV U88926 ( .A(n68737), .Z(n68738) );
  NOR U88927 ( .A(n68739), .B(n68738), .Z(n71191) );
  XOR U88928 ( .A(n71193), .B(n71191), .Z(n73699) );
  IV U88929 ( .A(n68740), .Z(n68742) );
  NOR U88930 ( .A(n68742), .B(n68741), .Z(n73697) );
  XOR U88931 ( .A(n73699), .B(n73697), .Z(n71188) );
  XOR U88932 ( .A(n71187), .B(n71188), .Z(n71179) );
  IV U88933 ( .A(n68743), .Z(n68746) );
  NOR U88934 ( .A(n68746), .B(n71170), .Z(n71178) );
  IV U88935 ( .A(n68744), .Z(n68748) );
  XOR U88936 ( .A(n68746), .B(n68745), .Z(n68747) );
  NOR U88937 ( .A(n68748), .B(n68747), .Z(n71176) );
  NOR U88938 ( .A(n71178), .B(n71176), .Z(n68749) );
  XOR U88939 ( .A(n71179), .B(n68749), .Z(n71169) );
  XOR U88940 ( .A(n68750), .B(n71169), .Z(n73719) );
  XOR U88941 ( .A(n73717), .B(n73719), .Z(n73722) );
  IV U88942 ( .A(n68751), .Z(n68755) );
  NOR U88943 ( .A(n68753), .B(n68752), .Z(n68754) );
  IV U88944 ( .A(n68754), .Z(n68757) );
  NOR U88945 ( .A(n68755), .B(n68757), .Z(n73720) );
  XOR U88946 ( .A(n73722), .B(n73720), .Z(n71164) );
  IV U88947 ( .A(n68756), .Z(n68758) );
  NOR U88948 ( .A(n68758), .B(n68757), .Z(n71162) );
  XOR U88949 ( .A(n71164), .B(n71162), .Z(n71167) );
  IV U88950 ( .A(n68759), .Z(n68762) );
  NOR U88951 ( .A(n68773), .B(n68760), .Z(n68761) );
  IV U88952 ( .A(n68761), .Z(n68764) );
  NOR U88953 ( .A(n68762), .B(n68764), .Z(n71165) );
  XOR U88954 ( .A(n71167), .B(n71165), .Z(n73727) );
  IV U88955 ( .A(n68763), .Z(n68765) );
  NOR U88956 ( .A(n68765), .B(n68764), .Z(n73725) );
  XOR U88957 ( .A(n73727), .B(n73725), .Z(n73730) );
  IV U88958 ( .A(n68766), .Z(n68770) );
  NOR U88959 ( .A(n68768), .B(n68767), .Z(n68769) );
  IV U88960 ( .A(n68769), .Z(n68776) );
  NOR U88961 ( .A(n68770), .B(n68776), .Z(n73723) );
  IV U88962 ( .A(n68771), .Z(n68772) );
  NOR U88963 ( .A(n68773), .B(n68772), .Z(n73728) );
  NOR U88964 ( .A(n73723), .B(n73728), .Z(n68774) );
  XOR U88965 ( .A(n73730), .B(n68774), .Z(n71155) );
  IV U88966 ( .A(n68775), .Z(n68777) );
  NOR U88967 ( .A(n68777), .B(n68776), .Z(n68778) );
  IV U88968 ( .A(n68778), .Z(n71156) );
  XOR U88969 ( .A(n71155), .B(n71156), .Z(n71160) );
  XOR U88970 ( .A(n71158), .B(n71160), .Z(n79140) );
  XOR U88971 ( .A(n71154), .B(n79140), .Z(n71148) );
  IV U88972 ( .A(n68779), .Z(n68780) );
  NOR U88973 ( .A(n68781), .B(n68780), .Z(n76559) );
  IV U88974 ( .A(n68782), .Z(n68783) );
  NOR U88975 ( .A(n68784), .B(n68783), .Z(n76555) );
  NOR U88976 ( .A(n76559), .B(n76555), .Z(n71149) );
  XOR U88977 ( .A(n71148), .B(n71149), .Z(n71152) );
  XOR U88978 ( .A(n71150), .B(n71152), .Z(n71143) );
  XOR U88979 ( .A(n71142), .B(n71143), .Z(n71146) );
  NOR U88980 ( .A(n68791), .B(n71146), .Z(n76543) );
  IV U88981 ( .A(n68785), .Z(n68786) );
  NOR U88982 ( .A(n68787), .B(n68786), .Z(n71145) );
  XOR U88983 ( .A(n71145), .B(n71146), .Z(n71141) );
  IV U88984 ( .A(n68788), .Z(n68790) );
  NOR U88985 ( .A(n68790), .B(n68789), .Z(n68792) );
  IV U88986 ( .A(n68792), .Z(n71140) );
  XOR U88987 ( .A(n71141), .B(n71140), .Z(n68794) );
  NOR U88988 ( .A(n68792), .B(n68791), .Z(n68793) );
  NOR U88989 ( .A(n68794), .B(n68793), .Z(n68795) );
  NOR U88990 ( .A(n76543), .B(n68795), .Z(n73737) );
  XOR U88991 ( .A(n73739), .B(n73737), .Z(n73741) );
  XOR U88992 ( .A(n73740), .B(n73741), .Z(n73747) );
  IV U88993 ( .A(n68796), .Z(n68798) );
  NOR U88994 ( .A(n68798), .B(n68797), .Z(n73745) );
  XOR U88995 ( .A(n73747), .B(n73745), .Z(n76535) );
  IV U88996 ( .A(n68799), .Z(n68801) );
  NOR U88997 ( .A(n68801), .B(n68800), .Z(n79167) );
  IV U88998 ( .A(n68802), .Z(n68803) );
  NOR U88999 ( .A(n68804), .B(n68803), .Z(n76534) );
  NOR U89000 ( .A(n79167), .B(n76534), .Z(n73748) );
  XOR U89001 ( .A(n76535), .B(n73748), .Z(n68805) );
  IV U89002 ( .A(n68805), .Z(n73753) );
  XOR U89003 ( .A(n73751), .B(n73753), .Z(n73755) );
  XOR U89004 ( .A(n73754), .B(n73755), .Z(n71139) );
  XOR U89005 ( .A(n68806), .B(n71139), .Z(n71134) );
  XOR U89006 ( .A(n71132), .B(n71134), .Z(n73759) );
  XOR U89007 ( .A(n73758), .B(n73759), .Z(n73766) );
  IV U89008 ( .A(n68807), .Z(n68808) );
  NOR U89009 ( .A(n68809), .B(n68808), .Z(n73761) );
  IV U89010 ( .A(n68810), .Z(n68811) );
  NOR U89011 ( .A(n68812), .B(n68811), .Z(n73764) );
  NOR U89012 ( .A(n73761), .B(n73764), .Z(n68813) );
  XOR U89013 ( .A(n73766), .B(n68813), .Z(n73769) );
  IV U89014 ( .A(n68814), .Z(n68816) );
  NOR U89015 ( .A(n68816), .B(n68815), .Z(n68817) );
  IV U89016 ( .A(n68817), .Z(n73770) );
  XOR U89017 ( .A(n73769), .B(n73770), .Z(n71131) );
  XOR U89018 ( .A(n71129), .B(n71131), .Z(n73779) );
  XOR U89019 ( .A(n68818), .B(n73779), .Z(n73781) );
  IV U89020 ( .A(n68819), .Z(n68821) );
  NOR U89021 ( .A(n68821), .B(n68820), .Z(n73780) );
  IV U89022 ( .A(n68822), .Z(n68823) );
  NOR U89023 ( .A(n68827), .B(n68823), .Z(n73787) );
  NOR U89024 ( .A(n73780), .B(n73787), .Z(n68824) );
  XOR U89025 ( .A(n73781), .B(n68824), .Z(n73786) );
  IV U89026 ( .A(n68825), .Z(n68826) );
  NOR U89027 ( .A(n68827), .B(n68826), .Z(n73784) );
  XOR U89028 ( .A(n73786), .B(n73784), .Z(n73792) );
  XOR U89029 ( .A(n68828), .B(n73792), .Z(n68829) );
  IV U89030 ( .A(n68829), .Z(n73795) );
  IV U89031 ( .A(n68830), .Z(n68831) );
  NOR U89032 ( .A(n68831), .B(n68834), .Z(n71123) );
  NOR U89033 ( .A(n73794), .B(n71123), .Z(n68832) );
  XOR U89034 ( .A(n73795), .B(n68832), .Z(n71120) );
  IV U89035 ( .A(n68833), .Z(n68835) );
  NOR U89036 ( .A(n68835), .B(n68834), .Z(n71121) );
  IV U89037 ( .A(n68836), .Z(n68838) );
  NOR U89038 ( .A(n68838), .B(n68837), .Z(n73799) );
  NOR U89039 ( .A(n71121), .B(n73799), .Z(n68839) );
  XOR U89040 ( .A(n71120), .B(n68839), .Z(n73803) );
  XOR U89041 ( .A(n73802), .B(n73803), .Z(n73806) );
  XOR U89042 ( .A(n73805), .B(n73806), .Z(n71119) );
  IV U89043 ( .A(n68840), .Z(n68843) );
  IV U89044 ( .A(n68841), .Z(n68842) );
  NOR U89045 ( .A(n68843), .B(n68842), .Z(n71117) );
  XOR U89046 ( .A(n71119), .B(n71117), .Z(n71112) );
  XOR U89047 ( .A(n71111), .B(n71112), .Z(n71115) );
  IV U89048 ( .A(n68844), .Z(n68845) );
  NOR U89049 ( .A(n68846), .B(n68845), .Z(n71114) );
  IV U89050 ( .A(n68847), .Z(n68849) );
  NOR U89051 ( .A(n68849), .B(n68848), .Z(n71109) );
  NOR U89052 ( .A(n71114), .B(n71109), .Z(n68850) );
  XOR U89053 ( .A(n71115), .B(n68850), .Z(n71106) );
  IV U89054 ( .A(n68851), .Z(n68852) );
  NOR U89055 ( .A(n68852), .B(n68856), .Z(n73811) );
  IV U89056 ( .A(n68857), .Z(n68853) );
  NOR U89057 ( .A(n68853), .B(n68856), .Z(n71107) );
  NOR U89058 ( .A(n73811), .B(n71107), .Z(n68854) );
  XOR U89059 ( .A(n71106), .B(n68854), .Z(n73816) );
  IV U89060 ( .A(n68855), .Z(n68859) );
  XOR U89061 ( .A(n68857), .B(n68856), .Z(n68858) );
  NOR U89062 ( .A(n68859), .B(n68858), .Z(n73814) );
  XOR U89063 ( .A(n73816), .B(n73814), .Z(n73833) );
  IV U89064 ( .A(n68860), .Z(n68863) );
  IV U89065 ( .A(n68861), .Z(n68862) );
  NOR U89066 ( .A(n68863), .B(n68862), .Z(n73822) );
  XOR U89067 ( .A(n73833), .B(n73822), .Z(n71101) );
  XOR U89068 ( .A(n71102), .B(n71101), .Z(n68864) );
  IV U89069 ( .A(n68864), .Z(n71099) );
  XOR U89070 ( .A(n71098), .B(n71099), .Z(n73841) );
  NOR U89071 ( .A(n68868), .B(n73841), .Z(n82113) );
  IV U89072 ( .A(n68865), .Z(n68866) );
  NOR U89073 ( .A(n68867), .B(n68866), .Z(n71095) );
  XOR U89074 ( .A(n73840), .B(n73841), .Z(n71096) );
  IV U89075 ( .A(n71096), .Z(n68869) );
  XOR U89076 ( .A(n71095), .B(n68869), .Z(n68871) );
  NOR U89077 ( .A(n68869), .B(n68868), .Z(n68870) );
  NOR U89078 ( .A(n68871), .B(n68870), .Z(n68872) );
  NOR U89079 ( .A(n82113), .B(n68872), .Z(n68873) );
  IV U89080 ( .A(n68873), .Z(n71091) );
  XOR U89081 ( .A(n71090), .B(n71091), .Z(n73846) );
  IV U89082 ( .A(n68874), .Z(n68875) );
  NOR U89083 ( .A(n68875), .B(n68877), .Z(n71093) );
  IV U89084 ( .A(n68876), .Z(n68878) );
  NOR U89085 ( .A(n68878), .B(n68877), .Z(n73844) );
  NOR U89086 ( .A(n71093), .B(n73844), .Z(n68879) );
  XOR U89087 ( .A(n73846), .B(n68879), .Z(n73847) );
  XOR U89088 ( .A(n73848), .B(n73847), .Z(n73863) );
  XOR U89089 ( .A(n73861), .B(n73863), .Z(n73856) );
  XOR U89090 ( .A(n68880), .B(n73856), .Z(n73875) );
  XOR U89091 ( .A(n73876), .B(n73875), .Z(n73882) );
  XOR U89092 ( .A(n73877), .B(n73882), .Z(n68881) );
  NOR U89093 ( .A(n68882), .B(n68881), .Z(n76463) );
  IV U89094 ( .A(n68883), .Z(n68885) );
  NOR U89095 ( .A(n68885), .B(n68884), .Z(n73881) );
  NOR U89096 ( .A(n73877), .B(n73881), .Z(n68886) );
  XOR U89097 ( .A(n73882), .B(n68886), .Z(n68887) );
  NOR U89098 ( .A(n68888), .B(n68887), .Z(n68889) );
  NOR U89099 ( .A(n76463), .B(n68889), .Z(n71085) );
  IV U89100 ( .A(n68890), .Z(n68892) );
  NOR U89101 ( .A(n68892), .B(n68891), .Z(n71087) );
  IV U89102 ( .A(n68893), .Z(n68897) );
  NOR U89103 ( .A(n68895), .B(n68894), .Z(n68896) );
  IV U89104 ( .A(n68896), .Z(n68900) );
  NOR U89105 ( .A(n68897), .B(n68900), .Z(n71084) );
  NOR U89106 ( .A(n71087), .B(n71084), .Z(n68898) );
  XOR U89107 ( .A(n71085), .B(n68898), .Z(n71083) );
  IV U89108 ( .A(n68899), .Z(n68901) );
  NOR U89109 ( .A(n68901), .B(n68900), .Z(n71081) );
  XOR U89110 ( .A(n71083), .B(n71081), .Z(n73889) );
  XOR U89111 ( .A(n73887), .B(n73889), .Z(n76454) );
  XOR U89112 ( .A(n73890), .B(n76454), .Z(n68902) );
  IV U89113 ( .A(n68902), .Z(n73894) );
  XOR U89114 ( .A(n73893), .B(n73894), .Z(n73898) );
  IV U89115 ( .A(n68903), .Z(n68905) );
  NOR U89116 ( .A(n68905), .B(n68904), .Z(n73896) );
  XOR U89117 ( .A(n73898), .B(n73896), .Z(n82042) );
  NOR U89118 ( .A(n82040), .B(n68906), .Z(n71077) );
  IV U89119 ( .A(n68907), .Z(n68910) );
  IV U89120 ( .A(n68908), .Z(n68909) );
  NOR U89121 ( .A(n68910), .B(n68909), .Z(n71079) );
  NOR U89122 ( .A(n71077), .B(n71079), .Z(n68911) );
  XOR U89123 ( .A(n82042), .B(n68911), .Z(n73899) );
  XOR U89124 ( .A(n73900), .B(n73899), .Z(n73902) );
  XOR U89125 ( .A(n73901), .B(n73902), .Z(n82020) );
  IV U89126 ( .A(n68912), .Z(n68914) );
  IV U89127 ( .A(n68913), .Z(n73906) );
  NOR U89128 ( .A(n68914), .B(n73906), .Z(n82016) );
  NOR U89129 ( .A(n82026), .B(n82016), .Z(n68915) );
  IV U89130 ( .A(n68915), .Z(n85132) );
  XOR U89131 ( .A(n82020), .B(n85132), .Z(n71073) );
  NOR U89132 ( .A(n68917), .B(n68916), .Z(n68918) );
  IV U89133 ( .A(n68918), .Z(n68919) );
  NOR U89134 ( .A(n68919), .B(n73906), .Z(n71071) );
  XOR U89135 ( .A(n71073), .B(n71071), .Z(n71067) );
  XOR U89136 ( .A(n71065), .B(n71067), .Z(n71069) );
  XOR U89137 ( .A(n71068), .B(n71069), .Z(n73913) );
  XOR U89138 ( .A(n73912), .B(n73913), .Z(n73917) );
  XOR U89139 ( .A(n73915), .B(n73917), .Z(n79298) );
  XOR U89140 ( .A(n79297), .B(n79298), .Z(n79305) );
  XOR U89141 ( .A(n68920), .B(n79305), .Z(n71063) );
  XOR U89142 ( .A(n71061), .B(n71063), .Z(n71056) );
  XOR U89143 ( .A(n71055), .B(n71056), .Z(n71060) );
  XOR U89144 ( .A(n68922), .B(n68921), .Z(n68924) );
  IV U89145 ( .A(n68923), .Z(n68929) );
  NOR U89146 ( .A(n68924), .B(n68929), .Z(n68925) );
  IV U89147 ( .A(n68925), .Z(n68926) );
  NOR U89148 ( .A(n68927), .B(n68926), .Z(n71058) );
  XOR U89149 ( .A(n71060), .B(n71058), .Z(n71052) );
  IV U89150 ( .A(n68928), .Z(n68930) );
  NOR U89151 ( .A(n68930), .B(n68929), .Z(n71050) );
  XOR U89152 ( .A(n71052), .B(n71050), .Z(n76401) );
  IV U89153 ( .A(n68931), .Z(n68932) );
  NOR U89154 ( .A(n68933), .B(n68932), .Z(n76400) );
  IV U89155 ( .A(n68934), .Z(n68936) );
  NOR U89156 ( .A(n68936), .B(n68935), .Z(n79312) );
  NOR U89157 ( .A(n76400), .B(n79312), .Z(n71053) );
  XOR U89158 ( .A(n76401), .B(n71053), .Z(n71046) );
  XOR U89159 ( .A(n71048), .B(n71046), .Z(n73934) );
  XOR U89160 ( .A(n73933), .B(n73934), .Z(n73937) );
  XOR U89161 ( .A(n73936), .B(n73937), .Z(n71042) );
  XOR U89162 ( .A(n71040), .B(n71042), .Z(n71045) );
  XOR U89163 ( .A(n71043), .B(n71045), .Z(n73944) );
  XOR U89164 ( .A(n73943), .B(n73944), .Z(n71039) );
  XOR U89165 ( .A(n71037), .B(n71039), .Z(n71036) );
  XOR U89166 ( .A(n71034), .B(n71036), .Z(n73956) );
  XOR U89167 ( .A(n73955), .B(n73956), .Z(n73960) );
  XOR U89168 ( .A(n73958), .B(n73960), .Z(n71030) );
  XOR U89169 ( .A(n71028), .B(n71030), .Z(n71032) );
  XOR U89170 ( .A(n71031), .B(n71032), .Z(n73962) );
  XOR U89171 ( .A(n73961), .B(n73962), .Z(n73965) );
  XOR U89172 ( .A(n73964), .B(n73965), .Z(n71023) );
  XOR U89173 ( .A(n71022), .B(n71023), .Z(n71026) );
  XOR U89174 ( .A(n71025), .B(n71026), .Z(n73969) );
  XOR U89175 ( .A(n73968), .B(n73969), .Z(n81946) );
  XOR U89176 ( .A(n73971), .B(n81946), .Z(n71015) );
  IV U89177 ( .A(n68937), .Z(n68939) );
  NOR U89178 ( .A(n68939), .B(n68938), .Z(n71019) );
  IV U89179 ( .A(n68940), .Z(n68942) );
  NOR U89180 ( .A(n68942), .B(n68941), .Z(n71016) );
  NOR U89181 ( .A(n71019), .B(n71016), .Z(n68943) );
  XOR U89182 ( .A(n71015), .B(n68943), .Z(n73978) );
  XOR U89183 ( .A(n73976), .B(n73978), .Z(n73989) );
  XOR U89184 ( .A(n71013), .B(n73989), .Z(n73997) );
  XOR U89185 ( .A(n68944), .B(n73997), .Z(n68945) );
  IV U89186 ( .A(n68945), .Z(n90895) );
  XOR U89187 ( .A(n71008), .B(n90895), .Z(n73994) );
  IV U89188 ( .A(n68946), .Z(n68950) );
  NOR U89189 ( .A(n68956), .B(n68947), .Z(n68948) );
  IV U89190 ( .A(n68948), .Z(n68949) );
  NOR U89191 ( .A(n68950), .B(n68949), .Z(n73992) );
  XOR U89192 ( .A(n73994), .B(n73992), .Z(n68966) );
  IV U89193 ( .A(n68966), .Z(n68962) );
  IV U89194 ( .A(n68951), .Z(n68952) );
  NOR U89195 ( .A(n68956), .B(n68952), .Z(n68963) );
  IV U89196 ( .A(n68953), .Z(n68959) );
  IV U89197 ( .A(n68954), .Z(n68955) );
  NOR U89198 ( .A(n68956), .B(n68955), .Z(n68957) );
  IV U89199 ( .A(n68957), .Z(n68958) );
  NOR U89200 ( .A(n68959), .B(n68958), .Z(n68965) );
  NOR U89201 ( .A(n68963), .B(n68965), .Z(n68960) );
  IV U89202 ( .A(n68960), .Z(n68961) );
  NOR U89203 ( .A(n68962), .B(n68961), .Z(n68968) );
  IV U89204 ( .A(n68963), .Z(n68964) );
  NOR U89205 ( .A(n68964), .B(n73994), .Z(n76368) );
  IV U89206 ( .A(n68965), .Z(n68967) );
  NOR U89207 ( .A(n68967), .B(n68966), .Z(n76370) );
  NOR U89208 ( .A(n76368), .B(n76370), .Z(n74003) );
  IV U89209 ( .A(n74003), .Z(n74013) );
  NOR U89210 ( .A(n68968), .B(n74013), .Z(n68969) );
  IV U89211 ( .A(n68969), .Z(n74011) );
  XOR U89212 ( .A(n74010), .B(n74011), .Z(n74005) );
  XOR U89213 ( .A(n74004), .B(n74005), .Z(n74023) );
  XOR U89214 ( .A(n74022), .B(n74023), .Z(n71005) );
  XOR U89215 ( .A(n71004), .B(n71005), .Z(n74020) );
  XOR U89216 ( .A(n74019), .B(n74020), .Z(n70999) );
  XOR U89217 ( .A(n70998), .B(n70999), .Z(n71002) );
  XOR U89218 ( .A(n68970), .B(n71002), .Z(n70992) );
  XOR U89219 ( .A(n70993), .B(n70992), .Z(n70989) );
  IV U89220 ( .A(n68971), .Z(n68973) );
  NOR U89221 ( .A(n68973), .B(n68972), .Z(n70987) );
  XOR U89222 ( .A(n70989), .B(n70987), .Z(n74034) );
  IV U89223 ( .A(n68974), .Z(n68982) );
  NOR U89224 ( .A(n68982), .B(n68975), .Z(n70990) );
  IV U89225 ( .A(n68976), .Z(n68978) );
  NOR U89226 ( .A(n68978), .B(n68977), .Z(n74033) );
  NOR U89227 ( .A(n70990), .B(n74033), .Z(n68979) );
  XOR U89228 ( .A(n74034), .B(n68979), .Z(n70983) );
  IV U89229 ( .A(n68980), .Z(n68981) );
  NOR U89230 ( .A(n68982), .B(n68981), .Z(n68983) );
  IV U89231 ( .A(n68983), .Z(n70984) );
  XOR U89232 ( .A(n70983), .B(n70984), .Z(n70982) );
  XOR U89233 ( .A(n68984), .B(n70982), .Z(n70974) );
  IV U89234 ( .A(n68985), .Z(n68986) );
  NOR U89235 ( .A(n68986), .B(n68988), .Z(n70972) );
  XOR U89236 ( .A(n70974), .B(n70972), .Z(n70977) );
  IV U89237 ( .A(n68987), .Z(n68989) );
  NOR U89238 ( .A(n68989), .B(n68988), .Z(n70975) );
  IV U89239 ( .A(n68990), .Z(n68996) );
  IV U89240 ( .A(n68991), .Z(n68992) );
  NOR U89241 ( .A(n68996), .B(n68992), .Z(n70970) );
  NOR U89242 ( .A(n70975), .B(n70970), .Z(n68993) );
  XOR U89243 ( .A(n70977), .B(n68993), .Z(n70961) );
  IV U89244 ( .A(n68994), .Z(n68995) );
  NOR U89245 ( .A(n68996), .B(n68995), .Z(n68997) );
  IV U89246 ( .A(n68997), .Z(n70968) );
  XOR U89247 ( .A(n70961), .B(n70968), .Z(n69002) );
  NOR U89248 ( .A(n69004), .B(n69002), .Z(n79386) );
  IV U89249 ( .A(n68998), .Z(n69000) );
  NOR U89250 ( .A(n69000), .B(n68999), .Z(n70954) );
  NOR U89251 ( .A(n69001), .B(n70962), .Z(n69003) );
  XOR U89252 ( .A(n69003), .B(n69002), .Z(n70955) );
  IV U89253 ( .A(n70955), .Z(n69005) );
  XOR U89254 ( .A(n70954), .B(n69005), .Z(n69007) );
  NOR U89255 ( .A(n69005), .B(n69004), .Z(n69006) );
  NOR U89256 ( .A(n69007), .B(n69006), .Z(n69008) );
  NOR U89257 ( .A(n79386), .B(n69008), .Z(n69009) );
  IV U89258 ( .A(n69009), .Z(n70958) );
  XOR U89259 ( .A(n70957), .B(n70958), .Z(n70949) );
  XOR U89260 ( .A(n70948), .B(n70949), .Z(n70952) );
  XOR U89261 ( .A(n70951), .B(n70952), .Z(n70946) );
  XOR U89262 ( .A(n70945), .B(n70946), .Z(n74049) );
  XOR U89263 ( .A(n74048), .B(n74049), .Z(n74052) );
  XOR U89264 ( .A(n74051), .B(n74052), .Z(n70940) );
  XOR U89265 ( .A(n70939), .B(n70940), .Z(n70944) );
  IV U89266 ( .A(n69010), .Z(n69012) );
  NOR U89267 ( .A(n69012), .B(n69011), .Z(n70942) );
  XOR U89268 ( .A(n70944), .B(n70942), .Z(n70934) );
  XOR U89269 ( .A(n70933), .B(n70934), .Z(n76324) );
  XOR U89270 ( .A(n70936), .B(n76324), .Z(n79422) );
  XOR U89271 ( .A(n69013), .B(n79422), .Z(n74069) );
  XOR U89272 ( .A(n74062), .B(n74069), .Z(n69014) );
  XOR U89273 ( .A(n69015), .B(n69014), .Z(n70924) );
  XOR U89274 ( .A(n69016), .B(n70924), .Z(n70928) );
  XOR U89275 ( .A(n69017), .B(n70928), .Z(n69018) );
  IV U89276 ( .A(n69018), .Z(n70921) );
  XOR U89277 ( .A(n70919), .B(n70921), .Z(n74075) );
  IV U89278 ( .A(n69019), .Z(n69021) );
  NOR U89279 ( .A(n69021), .B(n69020), .Z(n74073) );
  XOR U89280 ( .A(n74075), .B(n74073), .Z(n74076) );
  XOR U89281 ( .A(n74077), .B(n74076), .Z(n70913) );
  IV U89282 ( .A(n69022), .Z(n69023) );
  NOR U89283 ( .A(n69024), .B(n69023), .Z(n70915) );
  IV U89284 ( .A(n69025), .Z(n69027) );
  NOR U89285 ( .A(n69027), .B(n69026), .Z(n70912) );
  NOR U89286 ( .A(n70915), .B(n70912), .Z(n69028) );
  XOR U89287 ( .A(n70913), .B(n69028), .Z(n70907) );
  XOR U89288 ( .A(n70906), .B(n70907), .Z(n70911) );
  XOR U89289 ( .A(n70909), .B(n70911), .Z(n70902) );
  XOR U89290 ( .A(n70900), .B(n70902), .Z(n70904) );
  XOR U89291 ( .A(n70903), .B(n70904), .Z(n70898) );
  XOR U89292 ( .A(n69029), .B(n70898), .Z(n70890) );
  IV U89293 ( .A(n69030), .Z(n69031) );
  NOR U89294 ( .A(n69031), .B(n69033), .Z(n70894) );
  IV U89295 ( .A(n69032), .Z(n69034) );
  NOR U89296 ( .A(n69034), .B(n69033), .Z(n70889) );
  NOR U89297 ( .A(n70894), .B(n70889), .Z(n69035) );
  XOR U89298 ( .A(n70890), .B(n69035), .Z(n74085) );
  IV U89299 ( .A(n69036), .Z(n69038) );
  NOR U89300 ( .A(n69038), .B(n69037), .Z(n74083) );
  XOR U89301 ( .A(n74085), .B(n74083), .Z(n74087) );
  XOR U89302 ( .A(n74086), .B(n74087), .Z(n70885) );
  XOR U89303 ( .A(n70884), .B(n70885), .Z(n76304) );
  XOR U89304 ( .A(n70887), .B(n76304), .Z(n70876) );
  IV U89305 ( .A(n69039), .Z(n69040) );
  NOR U89306 ( .A(n69041), .B(n69040), .Z(n70881) );
  IV U89307 ( .A(n69042), .Z(n69045) );
  IV U89308 ( .A(n69043), .Z(n69044) );
  NOR U89309 ( .A(n69045), .B(n69044), .Z(n70875) );
  NOR U89310 ( .A(n70881), .B(n70875), .Z(n69046) );
  XOR U89311 ( .A(n70876), .B(n69046), .Z(n70880) );
  XOR U89312 ( .A(n70878), .B(n70880), .Z(n70871) );
  XOR U89313 ( .A(n70870), .B(n70871), .Z(n76296) );
  XOR U89314 ( .A(n70873), .B(n76296), .Z(n70868) );
  IV U89315 ( .A(n69047), .Z(n69049) );
  NOR U89316 ( .A(n69049), .B(n69048), .Z(n79516) );
  IV U89317 ( .A(n69050), .Z(n69051) );
  NOR U89318 ( .A(n69052), .B(n69051), .Z(n79524) );
  NOR U89319 ( .A(n79516), .B(n79524), .Z(n70869) );
  XOR U89320 ( .A(n70868), .B(n70869), .Z(n70864) );
  XOR U89321 ( .A(n70862), .B(n70864), .Z(n70866) );
  XOR U89322 ( .A(n70865), .B(n70866), .Z(n70858) );
  XOR U89323 ( .A(n70856), .B(n70858), .Z(n70860) );
  XOR U89324 ( .A(n69053), .B(n70860), .Z(n70845) );
  XOR U89325 ( .A(n70846), .B(n70845), .Z(n79549) );
  XOR U89326 ( .A(n69054), .B(n79549), .Z(n70838) );
  IV U89327 ( .A(n69055), .Z(n69057) );
  NOR U89328 ( .A(n69057), .B(n69056), .Z(n70842) );
  IV U89329 ( .A(n69058), .Z(n69060) );
  NOR U89330 ( .A(n69060), .B(n69059), .Z(n70837) );
  NOR U89331 ( .A(n70842), .B(n70837), .Z(n69061) );
  XOR U89332 ( .A(n70838), .B(n69061), .Z(n70835) );
  XOR U89333 ( .A(n70833), .B(n70835), .Z(n70829) );
  XOR U89334 ( .A(n69062), .B(n70829), .Z(n74105) );
  NOR U89335 ( .A(n69063), .B(n76271), .Z(n69065) );
  NOR U89336 ( .A(n69065), .B(n69064), .Z(n69066) );
  XOR U89337 ( .A(n74105), .B(n69066), .Z(n76262) );
  XOR U89338 ( .A(n70824), .B(n76262), .Z(n70825) );
  XOR U89339 ( .A(n70826), .B(n70825), .Z(n70823) );
  XOR U89340 ( .A(n69067), .B(n70823), .Z(n70809) );
  XOR U89341 ( .A(n70810), .B(n70809), .Z(n74111) );
  IV U89342 ( .A(n69068), .Z(n69069) );
  NOR U89343 ( .A(n69070), .B(n69069), .Z(n74109) );
  XOR U89344 ( .A(n74111), .B(n74109), .Z(n74113) );
  IV U89345 ( .A(n69071), .Z(n69073) );
  NOR U89346 ( .A(n69073), .B(n69072), .Z(n74112) );
  IV U89347 ( .A(n69074), .Z(n69076) );
  NOR U89348 ( .A(n69076), .B(n69075), .Z(n70806) );
  NOR U89349 ( .A(n74112), .B(n70806), .Z(n69077) );
  XOR U89350 ( .A(n74113), .B(n69077), .Z(n69078) );
  IV U89351 ( .A(n69078), .Z(n70804) );
  XOR U89352 ( .A(n70802), .B(n70804), .Z(n74119) );
  XOR U89353 ( .A(n69079), .B(n74119), .Z(n69080) );
  IV U89354 ( .A(n69080), .Z(n70794) );
  XOR U89355 ( .A(n70793), .B(n70794), .Z(n74128) );
  IV U89356 ( .A(n69081), .Z(n69082) );
  NOR U89357 ( .A(n69083), .B(n69082), .Z(n70790) );
  IV U89358 ( .A(n69084), .Z(n69085) );
  NOR U89359 ( .A(n69085), .B(n74122), .Z(n74126) );
  NOR U89360 ( .A(n70790), .B(n74126), .Z(n69086) );
  XOR U89361 ( .A(n74128), .B(n69086), .Z(n70787) );
  IV U89362 ( .A(n69087), .Z(n69088) );
  NOR U89363 ( .A(n69089), .B(n69088), .Z(n70788) );
  IV U89364 ( .A(n69090), .Z(n69091) );
  NOR U89365 ( .A(n69091), .B(n69095), .Z(n74130) );
  NOR U89366 ( .A(n70788), .B(n74130), .Z(n69092) );
  XOR U89367 ( .A(n70787), .B(n69092), .Z(n81741) );
  IV U89368 ( .A(n69093), .Z(n69094) );
  NOR U89369 ( .A(n69095), .B(n69094), .Z(n81740) );
  IV U89370 ( .A(n69096), .Z(n69097) );
  NOR U89371 ( .A(n81733), .B(n69097), .Z(n69098) );
  NOR U89372 ( .A(n81740), .B(n69098), .Z(n74129) );
  XOR U89373 ( .A(n81741), .B(n74129), .Z(n70780) );
  XOR U89374 ( .A(n70786), .B(n70780), .Z(n70775) );
  XOR U89375 ( .A(n69099), .B(n70775), .Z(n70764) );
  XOR U89376 ( .A(n69100), .B(n70764), .Z(n79605) );
  XOR U89377 ( .A(n70763), .B(n79605), .Z(n70753) );
  IV U89378 ( .A(n69101), .Z(n69102) );
  NOR U89379 ( .A(n69103), .B(n69102), .Z(n70760) );
  NOR U89380 ( .A(n69104), .B(n70754), .Z(n69105) );
  NOR U89381 ( .A(n70760), .B(n69105), .Z(n69106) );
  XOR U89382 ( .A(n70753), .B(n69106), .Z(n76196) );
  XOR U89383 ( .A(n69107), .B(n76196), .Z(n74144) );
  IV U89384 ( .A(n69108), .Z(n69110) );
  NOR U89385 ( .A(n69110), .B(n69109), .Z(n70749) );
  IV U89386 ( .A(n69111), .Z(n69113) );
  NOR U89387 ( .A(n69113), .B(n69112), .Z(n74143) );
  NOR U89388 ( .A(n70749), .B(n74143), .Z(n69114) );
  XOR U89389 ( .A(n74144), .B(n69114), .Z(n70744) );
  IV U89390 ( .A(n69115), .Z(n69117) );
  NOR U89391 ( .A(n69117), .B(n69116), .Z(n74138) );
  NOR U89392 ( .A(n69118), .B(n70745), .Z(n69119) );
  NOR U89393 ( .A(n74138), .B(n69119), .Z(n69120) );
  XOR U89394 ( .A(n70744), .B(n69120), .Z(n74164) );
  IV U89395 ( .A(n69121), .Z(n69122) );
  NOR U89396 ( .A(n69122), .B(n70745), .Z(n74162) );
  XOR U89397 ( .A(n74164), .B(n74162), .Z(n74165) );
  XOR U89398 ( .A(n74166), .B(n74165), .Z(n70738) );
  IV U89399 ( .A(n69123), .Z(n69124) );
  NOR U89400 ( .A(n69125), .B(n69124), .Z(n70740) );
  IV U89401 ( .A(n69126), .Z(n69128) );
  NOR U89402 ( .A(n69128), .B(n69127), .Z(n70737) );
  NOR U89403 ( .A(n70740), .B(n70737), .Z(n69129) );
  XOR U89404 ( .A(n70738), .B(n69129), .Z(n74171) );
  XOR U89405 ( .A(n74169), .B(n74171), .Z(n74174) );
  XOR U89406 ( .A(n74172), .B(n74174), .Z(n74183) );
  XOR U89407 ( .A(n69130), .B(n74183), .Z(n70734) );
  XOR U89408 ( .A(n70732), .B(n70734), .Z(n74189) );
  IV U89409 ( .A(n69131), .Z(n69133) );
  NOR U89410 ( .A(n69133), .B(n69132), .Z(n74187) );
  XOR U89411 ( .A(n74189), .B(n74187), .Z(n70731) );
  IV U89412 ( .A(n69134), .Z(n69136) );
  NOR U89413 ( .A(n69136), .B(n69135), .Z(n70729) );
  XOR U89414 ( .A(n70731), .B(n70729), .Z(n74205) );
  IV U89415 ( .A(n69137), .Z(n70726) );
  NOR U89416 ( .A(n70726), .B(n69138), .Z(n69142) );
  IV U89417 ( .A(n69139), .Z(n69141) );
  NOR U89418 ( .A(n69141), .B(n69140), .Z(n74204) );
  NOR U89419 ( .A(n69142), .B(n74204), .Z(n69143) );
  XOR U89420 ( .A(n74205), .B(n69143), .Z(n70721) );
  NOR U89421 ( .A(n69145), .B(n69144), .Z(n69146) );
  IV U89422 ( .A(n69146), .Z(n69147) );
  NOR U89423 ( .A(n69148), .B(n69147), .Z(n69149) );
  IV U89424 ( .A(n69149), .Z(n70722) );
  XOR U89425 ( .A(n70721), .B(n70722), .Z(n74218) );
  XOR U89426 ( .A(n74216), .B(n74218), .Z(n74226) );
  XOR U89427 ( .A(n74219), .B(n74226), .Z(n74224) );
  XOR U89428 ( .A(n74222), .B(n74224), .Z(n74242) );
  XOR U89429 ( .A(n69150), .B(n74242), .Z(n70718) );
  XOR U89430 ( .A(n70719), .B(n70718), .Z(n76167) );
  IV U89431 ( .A(n76167), .Z(n69157) );
  IV U89432 ( .A(n69151), .Z(n69152) );
  NOR U89433 ( .A(n69153), .B(n69152), .Z(n76170) );
  IV U89434 ( .A(n69154), .Z(n69156) );
  NOR U89435 ( .A(n69156), .B(n69155), .Z(n76164) );
  NOR U89436 ( .A(n76170), .B(n76164), .Z(n70713) );
  XOR U89437 ( .A(n69157), .B(n70713), .Z(n70715) );
  XOR U89438 ( .A(n70714), .B(n70715), .Z(n85470) );
  XOR U89439 ( .A(n70709), .B(n85470), .Z(n70704) );
  IV U89440 ( .A(n69158), .Z(n69160) );
  NOR U89441 ( .A(n69160), .B(n69159), .Z(n70710) );
  IV U89442 ( .A(n69161), .Z(n69163) );
  NOR U89443 ( .A(n69163), .B(n69162), .Z(n70703) );
  NOR U89444 ( .A(n70710), .B(n70703), .Z(n69164) );
  XOR U89445 ( .A(n70704), .B(n69164), .Z(n70707) );
  XOR U89446 ( .A(n70706), .B(n70707), .Z(n76148) );
  XOR U89447 ( .A(n69165), .B(n76148), .Z(n74255) );
  IV U89448 ( .A(n69166), .Z(n69168) );
  NOR U89449 ( .A(n69168), .B(n69167), .Z(n74253) );
  XOR U89450 ( .A(n74255), .B(n74253), .Z(n74259) );
  XOR U89451 ( .A(n74258), .B(n74259), .Z(n76144) );
  IV U89452 ( .A(n76144), .Z(n69175) );
  IV U89453 ( .A(n69169), .Z(n69170) );
  NOR U89454 ( .A(n69171), .B(n69170), .Z(n76142) );
  IV U89455 ( .A(n69172), .Z(n69173) );
  NOR U89456 ( .A(n69174), .B(n69173), .Z(n79696) );
  NOR U89457 ( .A(n76142), .B(n79696), .Z(n74261) );
  XOR U89458 ( .A(n69175), .B(n74261), .Z(n74265) );
  XOR U89459 ( .A(n74264), .B(n74265), .Z(n74275) );
  XOR U89460 ( .A(n69176), .B(n74275), .Z(n74270) );
  XOR U89461 ( .A(n74271), .B(n74270), .Z(n70701) );
  IV U89462 ( .A(n70701), .Z(n69184) );
  IV U89463 ( .A(n69177), .Z(n69179) );
  NOR U89464 ( .A(n69179), .B(n69178), .Z(n70700) );
  IV U89465 ( .A(n69180), .Z(n69182) );
  NOR U89466 ( .A(n69182), .B(n69181), .Z(n70698) );
  NOR U89467 ( .A(n70700), .B(n70698), .Z(n69183) );
  XOR U89468 ( .A(n69184), .B(n69183), .Z(n74277) );
  XOR U89469 ( .A(n74276), .B(n74277), .Z(n74280) );
  NOR U89470 ( .A(n69187), .B(n74280), .Z(n76119) );
  XOR U89471 ( .A(n74279), .B(n74280), .Z(n74288) );
  IV U89472 ( .A(n69185), .Z(n69186) );
  NOR U89473 ( .A(n69186), .B(n69196), .Z(n69188) );
  IV U89474 ( .A(n69188), .Z(n74287) );
  XOR U89475 ( .A(n74288), .B(n74287), .Z(n69190) );
  NOR U89476 ( .A(n69188), .B(n69187), .Z(n69189) );
  NOR U89477 ( .A(n69190), .B(n69189), .Z(n69191) );
  NOR U89478 ( .A(n76119), .B(n69191), .Z(n74283) );
  IV U89479 ( .A(n69192), .Z(n69193) );
  NOR U89480 ( .A(n69194), .B(n69193), .Z(n74294) );
  IV U89481 ( .A(n69195), .Z(n69197) );
  NOR U89482 ( .A(n69197), .B(n69196), .Z(n74284) );
  NOR U89483 ( .A(n74294), .B(n74284), .Z(n69198) );
  XOR U89484 ( .A(n74283), .B(n69198), .Z(n74302) );
  XOR U89485 ( .A(n74298), .B(n74302), .Z(n74312) );
  XOR U89486 ( .A(n69199), .B(n74312), .Z(n69200) );
  IV U89487 ( .A(n69200), .Z(n74310) );
  XOR U89488 ( .A(n74308), .B(n74310), .Z(n79727) );
  XOR U89489 ( .A(n74304), .B(n79727), .Z(n76103) );
  XOR U89490 ( .A(n74322), .B(n76103), .Z(n74323) );
  XOR U89491 ( .A(n74325), .B(n74323), .Z(n74329) );
  XOR U89492 ( .A(n74328), .B(n74329), .Z(n74333) );
  XOR U89493 ( .A(n74331), .B(n74333), .Z(n74336) );
  NOR U89494 ( .A(n69206), .B(n74336), .Z(n76090) );
  NOR U89495 ( .A(n69202), .B(n69201), .Z(n70695) );
  IV U89496 ( .A(n69203), .Z(n69204) );
  NOR U89497 ( .A(n69205), .B(n69204), .Z(n74335) );
  XOR U89498 ( .A(n74335), .B(n74336), .Z(n70696) );
  IV U89499 ( .A(n70696), .Z(n69207) );
  XOR U89500 ( .A(n70695), .B(n69207), .Z(n69209) );
  NOR U89501 ( .A(n69207), .B(n69206), .Z(n69208) );
  NOR U89502 ( .A(n69209), .B(n69208), .Z(n69210) );
  NOR U89503 ( .A(n76090), .B(n69210), .Z(n69211) );
  IV U89504 ( .A(n69211), .Z(n70693) );
  XOR U89505 ( .A(n70692), .B(n70693), .Z(n74343) );
  NOR U89506 ( .A(n69213), .B(n69212), .Z(n74341) );
  XOR U89507 ( .A(n74343), .B(n74341), .Z(n70690) );
  XOR U89508 ( .A(n69214), .B(n70690), .Z(n74350) );
  IV U89509 ( .A(n74350), .Z(n69219) );
  IV U89510 ( .A(n69215), .Z(n69217) );
  NOR U89511 ( .A(n69217), .B(n69216), .Z(n74349) );
  NOR U89512 ( .A(n70688), .B(n74349), .Z(n69218) );
  XOR U89513 ( .A(n69219), .B(n69218), .Z(n70684) );
  XOR U89514 ( .A(n70682), .B(n70684), .Z(n70686) );
  XOR U89515 ( .A(n69220), .B(n70686), .Z(n70680) );
  IV U89516 ( .A(n69221), .Z(n69223) );
  NOR U89517 ( .A(n69223), .B(n69222), .Z(n70679) );
  IV U89518 ( .A(n69224), .Z(n69225) );
  NOR U89519 ( .A(n69225), .B(n74353), .Z(n79743) );
  NOR U89520 ( .A(n70679), .B(n79743), .Z(n69226) );
  XOR U89521 ( .A(n70680), .B(n69226), .Z(n76068) );
  IV U89522 ( .A(n69227), .Z(n69228) );
  NOR U89523 ( .A(n69228), .B(n74353), .Z(n76066) );
  XOR U89524 ( .A(n76068), .B(n76066), .Z(n70673) );
  XOR U89525 ( .A(n70672), .B(n70673), .Z(n74372) );
  XOR U89526 ( .A(n69229), .B(n74372), .Z(n74367) );
  XOR U89527 ( .A(n74368), .B(n74367), .Z(n76056) );
  IV U89528 ( .A(n76056), .Z(n69236) );
  IV U89529 ( .A(n69230), .Z(n69231) );
  NOR U89530 ( .A(n69232), .B(n69231), .Z(n76062) );
  IV U89531 ( .A(n69233), .Z(n69235) );
  NOR U89532 ( .A(n69235), .B(n69234), .Z(n76054) );
  NOR U89533 ( .A(n76062), .B(n76054), .Z(n74375) );
  XOR U89534 ( .A(n69236), .B(n74375), .Z(n70670) );
  XOR U89535 ( .A(n70669), .B(n70670), .Z(n76049) );
  XOR U89536 ( .A(n70668), .B(n76049), .Z(n74385) );
  IV U89537 ( .A(n69237), .Z(n69239) );
  NOR U89538 ( .A(n69239), .B(n69238), .Z(n74386) );
  IV U89539 ( .A(n69240), .Z(n69241) );
  NOR U89540 ( .A(n69245), .B(n69241), .Z(n74390) );
  NOR U89541 ( .A(n74386), .B(n74390), .Z(n69242) );
  XOR U89542 ( .A(n74385), .B(n69242), .Z(n70666) );
  IV U89543 ( .A(n69243), .Z(n69244) );
  NOR U89544 ( .A(n69245), .B(n69244), .Z(n70664) );
  XOR U89545 ( .A(n70666), .B(n70664), .Z(n74400) );
  XOR U89546 ( .A(n74388), .B(n74400), .Z(n74404) );
  XOR U89547 ( .A(n69246), .B(n74404), .Z(n69247) );
  IV U89548 ( .A(n69247), .Z(n74407) );
  XOR U89549 ( .A(n74405), .B(n74407), .Z(n74409) );
  XOR U89550 ( .A(n74408), .B(n74409), .Z(n79794) );
  XOR U89551 ( .A(n74412), .B(n79794), .Z(n74416) );
  IV U89552 ( .A(n69248), .Z(n69249) );
  NOR U89553 ( .A(n79800), .B(n69249), .Z(n74414) );
  XOR U89554 ( .A(n74416), .B(n74414), .Z(n70660) );
  IV U89555 ( .A(n69250), .Z(n69252) );
  NOR U89556 ( .A(n69252), .B(n69251), .Z(n70658) );
  XOR U89557 ( .A(n70660), .B(n70658), .Z(n70662) );
  XOR U89558 ( .A(n70661), .B(n70662), .Z(n85544) );
  XOR U89559 ( .A(n85543), .B(n85544), .Z(n70655) );
  IV U89560 ( .A(n70655), .Z(n69260) );
  IV U89561 ( .A(n69253), .Z(n69255) );
  NOR U89562 ( .A(n69255), .B(n69254), .Z(n85552) );
  IV U89563 ( .A(n69256), .Z(n69258) );
  IV U89564 ( .A(n69257), .Z(n69262) );
  NOR U89565 ( .A(n69258), .B(n69262), .Z(n70653) );
  NOR U89566 ( .A(n85552), .B(n70653), .Z(n69259) );
  XOR U89567 ( .A(n69260), .B(n69259), .Z(n74422) );
  NOR U89568 ( .A(n69262), .B(n69261), .Z(n69263) );
  IV U89569 ( .A(n69263), .Z(n69268) );
  NOR U89570 ( .A(n69265), .B(n69264), .Z(n69266) );
  IV U89571 ( .A(n69266), .Z(n69267) );
  NOR U89572 ( .A(n69268), .B(n69267), .Z(n69269) );
  IV U89573 ( .A(n69269), .Z(n69270) );
  NOR U89574 ( .A(n69271), .B(n69270), .Z(n74420) );
  XOR U89575 ( .A(n74422), .B(n74420), .Z(n74432) );
  XOR U89576 ( .A(n69272), .B(n74432), .Z(n69273) );
  IV U89577 ( .A(n69273), .Z(n74429) );
  XOR U89578 ( .A(n74427), .B(n74429), .Z(n74435) );
  XOR U89579 ( .A(n74434), .B(n74435), .Z(n74438) );
  XOR U89580 ( .A(n74437), .B(n74438), .Z(n74442) );
  XOR U89581 ( .A(n74441), .B(n74442), .Z(n74446) );
  IV U89582 ( .A(n69274), .Z(n69277) );
  IV U89583 ( .A(n69275), .Z(n69276) );
  NOR U89584 ( .A(n69277), .B(n69276), .Z(n74444) );
  XOR U89585 ( .A(n74446), .B(n74444), .Z(n85590) );
  XOR U89586 ( .A(n69278), .B(n85590), .Z(n70646) );
  XOR U89587 ( .A(n70645), .B(n70646), .Z(n74449) );
  XOR U89588 ( .A(n74448), .B(n74449), .Z(n74452) );
  XOR U89589 ( .A(n74451), .B(n74452), .Z(n74458) );
  NOR U89590 ( .A(n69285), .B(n74458), .Z(n79822) );
  NOR U89591 ( .A(n69279), .B(n75998), .Z(n69282) );
  IV U89592 ( .A(n69280), .Z(n69281) );
  NOR U89593 ( .A(n69282), .B(n69281), .Z(n74459) );
  IV U89594 ( .A(n69283), .Z(n69284) );
  NOR U89595 ( .A(n69284), .B(n76001), .Z(n74456) );
  XOR U89596 ( .A(n74458), .B(n74456), .Z(n75999) );
  IV U89597 ( .A(n75999), .Z(n69286) );
  XOR U89598 ( .A(n74459), .B(n69286), .Z(n69288) );
  NOR U89599 ( .A(n69286), .B(n69285), .Z(n69287) );
  NOR U89600 ( .A(n69288), .B(n69287), .Z(n69289) );
  NOR U89601 ( .A(n79822), .B(n69289), .Z(n70642) );
  IV U89602 ( .A(n69290), .Z(n69291) );
  NOR U89603 ( .A(n69291), .B(n69293), .Z(n70641) );
  IV U89604 ( .A(n69292), .Z(n69294) );
  NOR U89605 ( .A(n69294), .B(n69293), .Z(n74463) );
  NOR U89606 ( .A(n70641), .B(n74463), .Z(n69295) );
  XOR U89607 ( .A(n70642), .B(n69295), .Z(n70636) );
  XOR U89608 ( .A(n70635), .B(n70636), .Z(n70640) );
  XOR U89609 ( .A(n70638), .B(n70640), .Z(n70633) );
  XOR U89610 ( .A(n70630), .B(n70633), .Z(n70628) );
  XOR U89611 ( .A(n69296), .B(n70628), .Z(n70618) );
  XOR U89612 ( .A(n69297), .B(n70618), .Z(n79846) );
  XOR U89613 ( .A(n69298), .B(n79846), .Z(n74476) );
  XOR U89614 ( .A(n74478), .B(n74476), .Z(n74472) );
  IV U89615 ( .A(n69299), .Z(n69301) );
  NOR U89616 ( .A(n69301), .B(n69300), .Z(n70609) );
  IV U89617 ( .A(n69302), .Z(n69304) );
  NOR U89618 ( .A(n69304), .B(n69303), .Z(n74470) );
  NOR U89619 ( .A(n70609), .B(n74470), .Z(n69305) );
  XOR U89620 ( .A(n74472), .B(n69305), .Z(n70607) );
  XOR U89621 ( .A(n69306), .B(n70607), .Z(n70603) );
  XOR U89622 ( .A(n70601), .B(n70603), .Z(n74482) );
  IV U89623 ( .A(n69307), .Z(n69321) );
  IV U89624 ( .A(n69308), .Z(n69309) );
  NOR U89625 ( .A(n69321), .B(n69309), .Z(n74480) );
  IV U89626 ( .A(n69310), .Z(n69312) );
  NOR U89627 ( .A(n69312), .B(n69311), .Z(n70604) );
  NOR U89628 ( .A(n74480), .B(n70604), .Z(n69313) );
  XOR U89629 ( .A(n74482), .B(n69313), .Z(n69323) );
  IV U89630 ( .A(n69323), .Z(n74484) );
  IV U89631 ( .A(n69314), .Z(n69315) );
  NOR U89632 ( .A(n69315), .B(n69317), .Z(n69316) );
  IV U89633 ( .A(n69316), .Z(n69324) );
  NOR U89634 ( .A(n74484), .B(n69324), .Z(n75951) );
  NOR U89635 ( .A(n69318), .B(n69317), .Z(n70598) );
  IV U89636 ( .A(n69319), .Z(n69320) );
  NOR U89637 ( .A(n69321), .B(n69320), .Z(n69322) );
  IV U89638 ( .A(n69322), .Z(n74483) );
  XOR U89639 ( .A(n69323), .B(n74483), .Z(n70599) );
  IV U89640 ( .A(n70599), .Z(n69325) );
  XOR U89641 ( .A(n70598), .B(n69325), .Z(n69327) );
  NOR U89642 ( .A(n69325), .B(n69324), .Z(n69326) );
  NOR U89643 ( .A(n69327), .B(n69326), .Z(n69328) );
  NOR U89644 ( .A(n75951), .B(n69328), .Z(n70592) );
  IV U89645 ( .A(n69329), .Z(n69332) );
  IV U89646 ( .A(n69330), .Z(n69331) );
  NOR U89647 ( .A(n69332), .B(n69331), .Z(n69333) );
  IV U89648 ( .A(n69333), .Z(n70593) );
  XOR U89649 ( .A(n70592), .B(n70593), .Z(n70596) );
  XOR U89650 ( .A(n70595), .B(n70596), .Z(n70585) );
  XOR U89651 ( .A(n70584), .B(n70585), .Z(n70588) );
  XOR U89652 ( .A(n70587), .B(n70588), .Z(n70582) );
  XOR U89653 ( .A(n70581), .B(n70582), .Z(n70576) );
  XOR U89654 ( .A(n70575), .B(n70576), .Z(n70579) );
  XOR U89655 ( .A(n70578), .B(n70579), .Z(n74491) );
  XOR U89656 ( .A(n74488), .B(n74491), .Z(n70574) );
  XOR U89657 ( .A(n69334), .B(n70574), .Z(n69335) );
  IV U89658 ( .A(n69335), .Z(n70568) );
  XOR U89659 ( .A(n70566), .B(n70568), .Z(n70570) );
  IV U89660 ( .A(n69336), .Z(n69337) );
  NOR U89661 ( .A(n69338), .B(n69337), .Z(n70569) );
  IV U89662 ( .A(n69339), .Z(n69341) );
  NOR U89663 ( .A(n69341), .B(n69340), .Z(n70563) );
  NOR U89664 ( .A(n70569), .B(n70563), .Z(n69342) );
  XOR U89665 ( .A(n70570), .B(n69342), .Z(n74499) );
  XOR U89666 ( .A(n69343), .B(n74499), .Z(n79893) );
  XOR U89667 ( .A(n70557), .B(n79893), .Z(n74506) );
  XOR U89668 ( .A(n74508), .B(n74506), .Z(n74504) );
  XOR U89669 ( .A(n69344), .B(n74504), .Z(n70546) );
  XOR U89670 ( .A(n70547), .B(n70546), .Z(n70549) );
  XOR U89671 ( .A(n70548), .B(n70549), .Z(n70542) );
  XOR U89672 ( .A(n70540), .B(n70542), .Z(n70545) );
  XOR U89673 ( .A(n70543), .B(n70545), .Z(n70535) );
  XOR U89674 ( .A(n70534), .B(n70535), .Z(n70538) );
  XOR U89675 ( .A(n69345), .B(n70538), .Z(n74518) );
  XOR U89676 ( .A(n74520), .B(n74518), .Z(n74522) );
  XOR U89677 ( .A(n74521), .B(n74522), .Z(n79950) );
  XOR U89678 ( .A(n79949), .B(n79950), .Z(n70516) );
  XOR U89679 ( .A(n69346), .B(n70516), .Z(n70524) );
  XOR U89680 ( .A(n70523), .B(n70524), .Z(n70522) );
  IV U89681 ( .A(n69347), .Z(n69349) );
  NOR U89682 ( .A(n69349), .B(n69348), .Z(n70520) );
  XOR U89683 ( .A(n70522), .B(n70520), .Z(n70510) );
  XOR U89684 ( .A(n70509), .B(n70510), .Z(n70513) );
  XOR U89685 ( .A(n70512), .B(n70513), .Z(n70508) );
  IV U89686 ( .A(n69350), .Z(n69351) );
  NOR U89687 ( .A(n69351), .B(n69353), .Z(n70506) );
  XOR U89688 ( .A(n70508), .B(n70506), .Z(n70502) );
  IV U89689 ( .A(n69352), .Z(n69354) );
  NOR U89690 ( .A(n69354), .B(n69353), .Z(n70500) );
  XOR U89691 ( .A(n70502), .B(n70500), .Z(n70504) );
  IV U89692 ( .A(n69355), .Z(n69356) );
  NOR U89693 ( .A(n69359), .B(n69356), .Z(n70503) );
  IV U89694 ( .A(n69357), .Z(n69358) );
  NOR U89695 ( .A(n69359), .B(n69358), .Z(n70497) );
  NOR U89696 ( .A(n70503), .B(n70497), .Z(n69360) );
  XOR U89697 ( .A(n70504), .B(n69360), .Z(n74529) );
  IV U89698 ( .A(n69361), .Z(n69363) );
  NOR U89699 ( .A(n69363), .B(n69362), .Z(n74528) );
  IV U89700 ( .A(n74528), .Z(n74530) );
  XOR U89701 ( .A(n74529), .B(n74530), .Z(n74537) );
  XOR U89702 ( .A(n69364), .B(n74537), .Z(n74538) );
  XOR U89703 ( .A(n74539), .B(n74538), .Z(n74548) );
  IV U89704 ( .A(n69365), .Z(n69366) );
  NOR U89705 ( .A(n69367), .B(n69366), .Z(n74541) );
  IV U89706 ( .A(n69368), .Z(n69370) );
  NOR U89707 ( .A(n69370), .B(n69369), .Z(n74547) );
  NOR U89708 ( .A(n74541), .B(n74547), .Z(n69371) );
  XOR U89709 ( .A(n74548), .B(n69371), .Z(n74544) );
  IV U89710 ( .A(n69372), .Z(n69374) );
  NOR U89711 ( .A(n69374), .B(n69373), .Z(n69375) );
  IV U89712 ( .A(n69375), .Z(n74545) );
  XOR U89713 ( .A(n74544), .B(n74545), .Z(n74553) );
  XOR U89714 ( .A(n74551), .B(n74553), .Z(n74556) );
  XOR U89715 ( .A(n74554), .B(n74556), .Z(n74561) );
  XOR U89716 ( .A(n74559), .B(n74561), .Z(n74564) );
  XOR U89717 ( .A(n74562), .B(n74564), .Z(n74567) );
  XOR U89718 ( .A(n74566), .B(n74567), .Z(n74572) );
  XOR U89719 ( .A(n69376), .B(n74572), .Z(n70495) );
  XOR U89720 ( .A(n70496), .B(n70495), .Z(n74579) );
  XOR U89721 ( .A(n74578), .B(n74579), .Z(n74586) );
  XOR U89722 ( .A(n69377), .B(n74586), .Z(n70492) );
  XOR U89723 ( .A(n70490), .B(n70492), .Z(n74593) );
  IV U89724 ( .A(n69378), .Z(n69380) );
  NOR U89725 ( .A(n69380), .B(n69379), .Z(n74591) );
  XOR U89726 ( .A(n74593), .B(n74591), .Z(n74603) );
  IV U89727 ( .A(n74603), .Z(n69389) );
  IV U89728 ( .A(n69383), .Z(n69382) );
  NOR U89729 ( .A(n69382), .B(n69381), .Z(n74594) );
  NOR U89730 ( .A(n69384), .B(n69383), .Z(n69387) );
  IV U89731 ( .A(n69385), .Z(n69386) );
  NOR U89732 ( .A(n69387), .B(n69386), .Z(n74601) );
  NOR U89733 ( .A(n74594), .B(n74601), .Z(n69388) );
  XOR U89734 ( .A(n69389), .B(n69388), .Z(n74600) );
  IV U89735 ( .A(n69390), .Z(n69392) );
  NOR U89736 ( .A(n69392), .B(n69391), .Z(n74598) );
  XOR U89737 ( .A(n74600), .B(n74598), .Z(n70488) );
  XOR U89738 ( .A(n69393), .B(n70488), .Z(n69394) );
  IV U89739 ( .A(n69394), .Z(n75819) );
  XOR U89740 ( .A(n70484), .B(n75819), .Z(n70480) );
  XOR U89741 ( .A(n70477), .B(n70480), .Z(n70476) );
  IV U89742 ( .A(n69395), .Z(n69397) );
  NOR U89743 ( .A(n69397), .B(n69396), .Z(n70479) );
  IV U89744 ( .A(n69398), .Z(n69399) );
  NOR U89745 ( .A(n69399), .B(n69403), .Z(n70474) );
  NOR U89746 ( .A(n70479), .B(n70474), .Z(n69400) );
  XOR U89747 ( .A(n70476), .B(n69400), .Z(n70465) );
  IV U89748 ( .A(n69410), .Z(n69408) );
  IV U89749 ( .A(n69401), .Z(n69411) );
  NOR U89750 ( .A(n69408), .B(n69411), .Z(n70466) );
  IV U89751 ( .A(n69402), .Z(n69404) );
  NOR U89752 ( .A(n69404), .B(n69403), .Z(n70471) );
  NOR U89753 ( .A(n70466), .B(n70471), .Z(n69405) );
  XOR U89754 ( .A(n70465), .B(n69405), .Z(n70469) );
  IV U89755 ( .A(n70469), .Z(n69415) );
  IV U89756 ( .A(n69406), .Z(n69407) );
  NOR U89757 ( .A(n69408), .B(n69407), .Z(n70468) );
  IV U89758 ( .A(n69409), .Z(n69413) );
  XOR U89759 ( .A(n69411), .B(n69410), .Z(n69412) );
  NOR U89760 ( .A(n69413), .B(n69412), .Z(n70460) );
  NOR U89761 ( .A(n70468), .B(n70460), .Z(n69414) );
  XOR U89762 ( .A(n69415), .B(n69414), .Z(n70464) );
  XOR U89763 ( .A(n70462), .B(n70464), .Z(n70457) );
  XOR U89764 ( .A(n70456), .B(n70457), .Z(n74612) );
  XOR U89765 ( .A(n74610), .B(n74612), .Z(n74634) );
  XOR U89766 ( .A(n69416), .B(n74634), .Z(n70450) );
  XOR U89767 ( .A(n69417), .B(n70450), .Z(n70455) );
  XOR U89768 ( .A(n70453), .B(n70455), .Z(n70448) );
  XOR U89769 ( .A(n70445), .B(n70448), .Z(n69418) );
  NOR U89770 ( .A(n69419), .B(n69418), .Z(n75795) );
  IV U89771 ( .A(n69420), .Z(n69421) );
  NOR U89772 ( .A(n69422), .B(n69421), .Z(n70447) );
  NOR U89773 ( .A(n70445), .B(n70447), .Z(n69423) );
  XOR U89774 ( .A(n70448), .B(n69423), .Z(n69424) );
  NOR U89775 ( .A(n69425), .B(n69424), .Z(n69426) );
  NOR U89776 ( .A(n75795), .B(n69426), .Z(n70442) );
  IV U89777 ( .A(n69427), .Z(n69428) );
  NOR U89778 ( .A(n69429), .B(n69428), .Z(n75790) );
  IV U89779 ( .A(n69430), .Z(n69432) );
  NOR U89780 ( .A(n69432), .B(n69431), .Z(n80060) );
  NOR U89781 ( .A(n75790), .B(n80060), .Z(n70443) );
  XOR U89782 ( .A(n70442), .B(n70443), .Z(n70441) );
  XOR U89783 ( .A(n70439), .B(n70441), .Z(n74642) );
  XOR U89784 ( .A(n69433), .B(n74642), .Z(n74654) );
  XOR U89785 ( .A(n74653), .B(n74654), .Z(n74658) );
  NOR U89786 ( .A(n69435), .B(n69434), .Z(n69436) );
  IV U89787 ( .A(n69436), .Z(n69441) );
  NOR U89788 ( .A(n69438), .B(n69437), .Z(n69439) );
  IV U89789 ( .A(n69439), .Z(n69440) );
  NOR U89790 ( .A(n69441), .B(n69440), .Z(n74656) );
  XOR U89791 ( .A(n74658), .B(n74656), .Z(n70437) );
  XOR U89792 ( .A(n70438), .B(n70437), .Z(n74667) );
  IV U89793 ( .A(n69442), .Z(n69443) );
  NOR U89794 ( .A(n69444), .B(n69443), .Z(n74666) );
  IV U89795 ( .A(n69445), .Z(n69446) );
  NOR U89796 ( .A(n69446), .B(n69449), .Z(n74669) );
  NOR U89797 ( .A(n74666), .B(n74669), .Z(n69447) );
  XOR U89798 ( .A(n74667), .B(n69447), .Z(n74676) );
  IV U89799 ( .A(n69448), .Z(n69450) );
  NOR U89800 ( .A(n69450), .B(n69449), .Z(n74672) );
  IV U89801 ( .A(n69451), .Z(n69453) );
  NOR U89802 ( .A(n69453), .B(n69452), .Z(n74674) );
  NOR U89803 ( .A(n74672), .B(n74674), .Z(n69454) );
  XOR U89804 ( .A(n74676), .B(n69454), .Z(n69455) );
  NOR U89805 ( .A(n69456), .B(n69455), .Z(n69459) );
  IV U89806 ( .A(n69456), .Z(n69458) );
  XOR U89807 ( .A(n74672), .B(n74676), .Z(n69457) );
  NOR U89808 ( .A(n69458), .B(n69457), .Z(n75784) );
  NOR U89809 ( .A(n69459), .B(n75784), .Z(n69460) );
  IV U89810 ( .A(n69460), .Z(n70433) );
  IV U89811 ( .A(n69461), .Z(n69463) );
  NOR U89812 ( .A(n69463), .B(n69462), .Z(n70431) );
  XOR U89813 ( .A(n70433), .B(n70431), .Z(n70436) );
  XOR U89814 ( .A(n70434), .B(n70436), .Z(n74686) );
  XOR U89815 ( .A(n69464), .B(n74686), .Z(n74682) );
  XOR U89816 ( .A(n74683), .B(n74682), .Z(n70429) );
  IV U89817 ( .A(n69465), .Z(n69467) );
  NOR U89818 ( .A(n69467), .B(n69466), .Z(n70428) );
  NOR U89819 ( .A(n69469), .B(n69468), .Z(n70421) );
  NOR U89820 ( .A(n70428), .B(n70421), .Z(n69470) );
  XOR U89821 ( .A(n70429), .B(n69470), .Z(n69471) );
  IV U89822 ( .A(n69471), .Z(n70424) );
  XOR U89823 ( .A(n69472), .B(n70424), .Z(n70414) );
  IV U89824 ( .A(n69473), .Z(n69474) );
  NOR U89825 ( .A(n69474), .B(n69476), .Z(n70416) );
  IV U89826 ( .A(n69475), .Z(n69477) );
  NOR U89827 ( .A(n69477), .B(n69476), .Z(n70413) );
  NOR U89828 ( .A(n70416), .B(n70413), .Z(n69478) );
  XOR U89829 ( .A(n70414), .B(n69478), .Z(n70411) );
  XOR U89830 ( .A(n70409), .B(n70411), .Z(n70407) );
  XOR U89831 ( .A(n70404), .B(n70407), .Z(n74694) );
  XOR U89832 ( .A(n69479), .B(n74694), .Z(n70401) );
  XOR U89833 ( .A(n69480), .B(n70401), .Z(n74700) );
  XOR U89834 ( .A(n69481), .B(n74700), .Z(n70398) );
  XOR U89835 ( .A(n70400), .B(n70398), .Z(n74705) );
  XOR U89836 ( .A(n69483), .B(n69482), .Z(n69484) );
  NOR U89837 ( .A(n69485), .B(n69484), .Z(n69486) );
  IV U89838 ( .A(n69486), .Z(n69487) );
  NOR U89839 ( .A(n69488), .B(n69487), .Z(n74704) );
  IV U89840 ( .A(n69489), .Z(n69491) );
  NOR U89841 ( .A(n69491), .B(n69490), .Z(n70394) );
  NOR U89842 ( .A(n74704), .B(n70394), .Z(n69492) );
  XOR U89843 ( .A(n74705), .B(n69492), .Z(n69493) );
  IV U89844 ( .A(n69493), .Z(n74709) );
  XOR U89845 ( .A(n74707), .B(n74709), .Z(n70392) );
  XOR U89846 ( .A(n70391), .B(n70392), .Z(n74714) );
  XOR U89847 ( .A(n74713), .B(n74714), .Z(n70389) );
  XOR U89848 ( .A(n70388), .B(n70389), .Z(n74727) );
  XOR U89849 ( .A(n74725), .B(n74727), .Z(n74729) );
  XOR U89850 ( .A(n74728), .B(n74729), .Z(n74733) );
  XOR U89851 ( .A(n74732), .B(n74733), .Z(n74739) );
  XOR U89852 ( .A(n69494), .B(n74739), .Z(n74742) );
  XOR U89853 ( .A(n74743), .B(n74742), .Z(n74746) );
  IV U89854 ( .A(n69495), .Z(n69497) );
  NOR U89855 ( .A(n69497), .B(n69496), .Z(n69498) );
  IV U89856 ( .A(n69498), .Z(n74745) );
  XOR U89857 ( .A(n74746), .B(n74745), .Z(n70386) );
  IV U89858 ( .A(n69499), .Z(n69501) );
  NOR U89859 ( .A(n69501), .B(n69500), .Z(n74750) );
  IV U89860 ( .A(n69502), .Z(n69504) );
  NOR U89861 ( .A(n69504), .B(n69503), .Z(n70385) );
  NOR U89862 ( .A(n74750), .B(n70385), .Z(n69505) );
  XOR U89863 ( .A(n70386), .B(n69505), .Z(n74762) );
  XOR U89864 ( .A(n74761), .B(n74762), .Z(n75741) );
  XOR U89865 ( .A(n74764), .B(n75741), .Z(n69506) );
  IV U89866 ( .A(n69506), .Z(n70382) );
  XOR U89867 ( .A(n70381), .B(n70382), .Z(n70376) );
  XOR U89868 ( .A(n70375), .B(n70376), .Z(n70379) );
  IV U89869 ( .A(n69507), .Z(n69509) );
  NOR U89870 ( .A(n69509), .B(n69508), .Z(n70372) );
  NOR U89871 ( .A(n70378), .B(n70372), .Z(n69510) );
  XOR U89872 ( .A(n70379), .B(n69510), .Z(n69520) );
  IV U89873 ( .A(n69520), .Z(n69511) );
  NOR U89874 ( .A(n69512), .B(n69511), .Z(n75724) );
  IV U89875 ( .A(n69513), .Z(n69514) );
  NOR U89876 ( .A(n69515), .B(n69514), .Z(n74768) );
  IV U89877 ( .A(n69516), .Z(n69517) );
  NOR U89878 ( .A(n69518), .B(n69517), .Z(n69521) );
  IV U89879 ( .A(n69521), .Z(n69519) );
  NOR U89880 ( .A(n69519), .B(n70379), .Z(n75727) );
  NOR U89881 ( .A(n69521), .B(n69520), .Z(n69522) );
  NOR U89882 ( .A(n75727), .B(n69522), .Z(n74769) );
  XOR U89883 ( .A(n74768), .B(n74769), .Z(n69523) );
  NOR U89884 ( .A(n69524), .B(n69523), .Z(n69525) );
  NOR U89885 ( .A(n75724), .B(n69525), .Z(n69526) );
  IV U89886 ( .A(n69526), .Z(n74775) );
  XOR U89887 ( .A(n70370), .B(n74775), .Z(n74779) );
  IV U89888 ( .A(n69527), .Z(n69529) );
  NOR U89889 ( .A(n69529), .B(n69528), .Z(n74774) );
  IV U89890 ( .A(n69530), .Z(n69532) );
  IV U89891 ( .A(n69531), .Z(n69535) );
  NOR U89892 ( .A(n69532), .B(n69535), .Z(n74777) );
  NOR U89893 ( .A(n74774), .B(n74777), .Z(n69533) );
  XOR U89894 ( .A(n74779), .B(n69533), .Z(n70366) );
  IV U89895 ( .A(n69534), .Z(n69536) );
  NOR U89896 ( .A(n69536), .B(n69535), .Z(n69537) );
  IV U89897 ( .A(n69537), .Z(n70367) );
  XOR U89898 ( .A(n70366), .B(n70367), .Z(n74781) );
  XOR U89899 ( .A(n74780), .B(n74781), .Z(n74784) );
  XOR U89900 ( .A(n69538), .B(n74784), .Z(n70357) );
  XOR U89901 ( .A(n69539), .B(n70357), .Z(n70351) );
  IV U89902 ( .A(n69540), .Z(n69541) );
  NOR U89903 ( .A(n69541), .B(n70358), .Z(n70349) );
  XOR U89904 ( .A(n70351), .B(n70349), .Z(n70352) );
  XOR U89905 ( .A(n70353), .B(n70352), .Z(n74788) );
  IV U89906 ( .A(n69542), .Z(n69543) );
  NOR U89907 ( .A(n69544), .B(n69543), .Z(n75700) );
  IV U89908 ( .A(n69545), .Z(n69547) );
  NOR U89909 ( .A(n69547), .B(n69546), .Z(n80201) );
  NOR U89910 ( .A(n75700), .B(n80201), .Z(n74789) );
  XOR U89911 ( .A(n74788), .B(n74789), .Z(n74792) );
  XOR U89912 ( .A(n74791), .B(n74792), .Z(n74796) );
  XOR U89913 ( .A(n74794), .B(n74796), .Z(n70346) );
  XOR U89914 ( .A(n70345), .B(n70346), .Z(n74803) );
  XOR U89915 ( .A(n74801), .B(n74803), .Z(n70344) );
  XOR U89916 ( .A(n70342), .B(n70344), .Z(n75686) );
  XOR U89917 ( .A(n69548), .B(n75686), .Z(n74816) );
  IV U89918 ( .A(n69549), .Z(n69551) );
  NOR U89919 ( .A(n69551), .B(n69550), .Z(n74814) );
  XOR U89920 ( .A(n74816), .B(n74814), .Z(n74826) );
  IV U89921 ( .A(n74826), .Z(n69559) );
  IV U89922 ( .A(n69552), .Z(n69553) );
  NOR U89923 ( .A(n69554), .B(n69553), .Z(n70340) );
  IV U89924 ( .A(n69555), .Z(n69557) );
  NOR U89925 ( .A(n69557), .B(n69556), .Z(n74825) );
  NOR U89926 ( .A(n70340), .B(n74825), .Z(n69558) );
  XOR U89927 ( .A(n69559), .B(n69558), .Z(n74822) );
  XOR U89928 ( .A(n74821), .B(n74822), .Z(n70338) );
  IV U89929 ( .A(n69560), .Z(n69566) );
  IV U89930 ( .A(n69561), .Z(n69562) );
  NOR U89931 ( .A(n69563), .B(n69562), .Z(n69564) );
  IV U89932 ( .A(n69564), .Z(n69565) );
  NOR U89933 ( .A(n69566), .B(n69565), .Z(n70337) );
  NOR U89934 ( .A(n70334), .B(n70336), .Z(n69567) );
  NOR U89935 ( .A(n70337), .B(n69567), .Z(n69568) );
  XOR U89936 ( .A(n70338), .B(n69568), .Z(n69569) );
  IV U89937 ( .A(n69569), .Z(n74837) );
  IV U89938 ( .A(n69570), .Z(n69572) );
  NOR U89939 ( .A(n69572), .B(n69571), .Z(n74835) );
  XOR U89940 ( .A(n74837), .B(n74835), .Z(n70333) );
  XOR U89941 ( .A(n69573), .B(n70333), .Z(n74850) );
  XOR U89942 ( .A(n74848), .B(n74850), .Z(n70327) );
  NOR U89943 ( .A(n69575), .B(n69574), .Z(n74852) );
  NOR U89944 ( .A(n69577), .B(n69576), .Z(n70326) );
  NOR U89945 ( .A(n74852), .B(n70326), .Z(n69578) );
  XOR U89946 ( .A(n70327), .B(n69578), .Z(n70320) );
  IV U89947 ( .A(n69579), .Z(n69580) );
  NOR U89948 ( .A(n69581), .B(n69580), .Z(n70321) );
  NOR U89949 ( .A(n70323), .B(n70321), .Z(n69582) );
  XOR U89950 ( .A(n70320), .B(n69582), .Z(n75670) );
  XOR U89951 ( .A(n74868), .B(n75670), .Z(n74870) );
  XOR U89952 ( .A(n69583), .B(n74870), .Z(n70319) );
  XOR U89953 ( .A(n69584), .B(n70319), .Z(n74879) );
  XOR U89954 ( .A(n70313), .B(n74879), .Z(n69585) );
  NOR U89955 ( .A(n69586), .B(n69585), .Z(n75655) );
  NOR U89956 ( .A(n69588), .B(n69587), .Z(n74878) );
  NOR U89957 ( .A(n70313), .B(n74878), .Z(n69589) );
  XOR U89958 ( .A(n74879), .B(n69589), .Z(n69590) );
  NOR U89959 ( .A(n69591), .B(n69590), .Z(n69592) );
  NOR U89960 ( .A(n75655), .B(n69592), .Z(n70311) );
  XOR U89961 ( .A(n69593), .B(n70311), .Z(n70306) );
  XOR U89962 ( .A(n70304), .B(n70306), .Z(n70309) );
  IV U89963 ( .A(n69594), .Z(n69595) );
  NOR U89964 ( .A(n69595), .B(n69600), .Z(n69596) );
  IV U89965 ( .A(n69596), .Z(n69597) );
  NOR U89966 ( .A(n69598), .B(n69597), .Z(n70307) );
  XOR U89967 ( .A(n70309), .B(n70307), .Z(n70300) );
  IV U89968 ( .A(n69599), .Z(n69603) );
  NOR U89969 ( .A(n69601), .B(n69600), .Z(n69602) );
  IV U89970 ( .A(n69602), .Z(n69605) );
  NOR U89971 ( .A(n69603), .B(n69605), .Z(n70298) );
  XOR U89972 ( .A(n70300), .B(n70298), .Z(n70303) );
  IV U89973 ( .A(n69604), .Z(n69606) );
  NOR U89974 ( .A(n69606), .B(n69605), .Z(n70301) );
  XOR U89975 ( .A(n70303), .B(n70301), .Z(n70297) );
  IV U89976 ( .A(n69607), .Z(n69612) );
  IV U89977 ( .A(n69608), .Z(n69609) );
  NOR U89978 ( .A(n69612), .B(n69609), .Z(n70295) );
  XOR U89979 ( .A(n70297), .B(n70295), .Z(n70291) );
  IV U89980 ( .A(n69610), .Z(n69611) );
  NOR U89981 ( .A(n69612), .B(n69611), .Z(n70289) );
  XOR U89982 ( .A(n70291), .B(n70289), .Z(n70293) );
  XOR U89983 ( .A(n70292), .B(n70293), .Z(n74895) );
  IV U89984 ( .A(n69613), .Z(n69615) );
  NOR U89985 ( .A(n69615), .B(n69614), .Z(n70287) );
  IV U89986 ( .A(n69616), .Z(n69617) );
  NOR U89987 ( .A(n69617), .B(n69621), .Z(n74893) );
  NOR U89988 ( .A(n70287), .B(n74893), .Z(n69618) );
  XOR U89989 ( .A(n74895), .B(n69618), .Z(n69619) );
  IV U89990 ( .A(n69619), .Z(n74898) );
  IV U89991 ( .A(n69620), .Z(n69622) );
  NOR U89992 ( .A(n69622), .B(n69621), .Z(n74896) );
  XOR U89993 ( .A(n74898), .B(n74896), .Z(n75621) );
  XOR U89994 ( .A(n74899), .B(n75621), .Z(n70285) );
  IV U89995 ( .A(n69623), .Z(n69625) );
  NOR U89996 ( .A(n69625), .B(n69624), .Z(n75613) );
  NOR U89997 ( .A(n75624), .B(n75613), .Z(n70286) );
  XOR U89998 ( .A(n70285), .B(n70286), .Z(n70281) );
  XOR U89999 ( .A(n70279), .B(n70281), .Z(n70283) );
  XOR U90000 ( .A(n70282), .B(n70283), .Z(n70277) );
  XOR U90001 ( .A(n69626), .B(n70277), .Z(n70269) );
  IV U90002 ( .A(n69627), .Z(n69628) );
  NOR U90003 ( .A(n69630), .B(n69628), .Z(n70268) );
  IV U90004 ( .A(n69629), .Z(n69631) );
  NOR U90005 ( .A(n69631), .B(n69630), .Z(n70271) );
  NOR U90006 ( .A(n70268), .B(n70271), .Z(n69632) );
  XOR U90007 ( .A(n70269), .B(n69632), .Z(n70267) );
  IV U90008 ( .A(n69633), .Z(n69634) );
  NOR U90009 ( .A(n69644), .B(n69634), .Z(n69648) );
  IV U90010 ( .A(n69648), .Z(n69635) );
  NOR U90011 ( .A(n70267), .B(n69635), .Z(n75605) );
  IV U90012 ( .A(n70267), .Z(n69642) );
  IV U90013 ( .A(n69636), .Z(n69638) );
  NOR U90014 ( .A(n69638), .B(n69637), .Z(n70265) );
  IV U90015 ( .A(n69639), .Z(n69640) );
  NOR U90016 ( .A(n69640), .B(n69644), .Z(n70261) );
  NOR U90017 ( .A(n70265), .B(n70261), .Z(n69641) );
  XOR U90018 ( .A(n69642), .B(n69641), .Z(n70264) );
  IV U90019 ( .A(n69643), .Z(n69645) );
  NOR U90020 ( .A(n69645), .B(n69644), .Z(n69646) );
  IV U90021 ( .A(n69646), .Z(n70263) );
  XOR U90022 ( .A(n70264), .B(n70263), .Z(n69647) );
  NOR U90023 ( .A(n69648), .B(n69647), .Z(n69649) );
  NOR U90024 ( .A(n75605), .B(n69649), .Z(n70258) );
  XOR U90025 ( .A(n70260), .B(n70258), .Z(n70254) );
  IV U90026 ( .A(n69650), .Z(n69652) );
  NOR U90027 ( .A(n69652), .B(n69651), .Z(n70252) );
  XOR U90028 ( .A(n70254), .B(n70252), .Z(n70256) );
  IV U90029 ( .A(n69653), .Z(n69654) );
  NOR U90030 ( .A(n69655), .B(n69654), .Z(n70255) );
  IV U90031 ( .A(n69656), .Z(n69658) );
  NOR U90032 ( .A(n69658), .B(n69657), .Z(n70250) );
  NOR U90033 ( .A(n70255), .B(n70250), .Z(n69659) );
  XOR U90034 ( .A(n70256), .B(n69659), .Z(n69660) );
  IV U90035 ( .A(n69660), .Z(n74909) );
  XOR U90036 ( .A(n74907), .B(n74909), .Z(n75585) );
  XOR U90037 ( .A(n74910), .B(n75585), .Z(n74919) );
  IV U90038 ( .A(n69661), .Z(n69663) );
  NOR U90039 ( .A(n69663), .B(n69662), .Z(n74921) );
  IV U90040 ( .A(n69664), .Z(n69666) );
  NOR U90041 ( .A(n69666), .B(n69665), .Z(n74918) );
  NOR U90042 ( .A(n74921), .B(n74918), .Z(n69667) );
  XOR U90043 ( .A(n74919), .B(n69667), .Z(n74915) );
  XOR U90044 ( .A(n74914), .B(n74915), .Z(n74932) );
  XOR U90045 ( .A(n69668), .B(n74932), .Z(n70243) );
  XOR U90046 ( .A(n70244), .B(n70243), .Z(n70242) );
  IV U90047 ( .A(n69669), .Z(n69670) );
  NOR U90048 ( .A(n69671), .B(n69670), .Z(n70245) );
  IV U90049 ( .A(n69672), .Z(n69673) );
  NOR U90050 ( .A(n69673), .B(n69678), .Z(n70240) );
  NOR U90051 ( .A(n70245), .B(n70240), .Z(n69674) );
  XOR U90052 ( .A(n70242), .B(n69674), .Z(n69675) );
  IV U90053 ( .A(n69675), .Z(n70239) );
  IV U90054 ( .A(n69676), .Z(n69677) );
  NOR U90055 ( .A(n69678), .B(n69677), .Z(n70237) );
  XOR U90056 ( .A(n70239), .B(n70237), .Z(n69679) );
  NOR U90057 ( .A(n69680), .B(n69679), .Z(n75577) );
  IV U90058 ( .A(n69681), .Z(n69683) );
  NOR U90059 ( .A(n69683), .B(n69682), .Z(n70235) );
  NOR U90060 ( .A(n70235), .B(n70237), .Z(n69684) );
  XOR U90061 ( .A(n70239), .B(n69684), .Z(n69685) );
  NOR U90062 ( .A(n69686), .B(n69685), .Z(n69687) );
  NOR U90063 ( .A(n75577), .B(n69687), .Z(n69688) );
  IV U90064 ( .A(n69688), .Z(n74936) );
  XOR U90065 ( .A(n74935), .B(n74936), .Z(n70231) );
  XOR U90066 ( .A(n70230), .B(n70231), .Z(n75565) );
  XOR U90067 ( .A(n69689), .B(n75565), .Z(n70225) );
  XOR U90068 ( .A(n70224), .B(n70225), .Z(n70228) );
  IV U90069 ( .A(n69690), .Z(n69691) );
  NOR U90070 ( .A(n69692), .B(n69691), .Z(n70227) );
  IV U90071 ( .A(n69693), .Z(n69695) );
  NOR U90072 ( .A(n69695), .B(n69694), .Z(n70221) );
  NOR U90073 ( .A(n70227), .B(n70221), .Z(n69696) );
  XOR U90074 ( .A(n70228), .B(n69696), .Z(n69697) );
  NOR U90075 ( .A(n69698), .B(n69697), .Z(n69701) );
  IV U90076 ( .A(n69698), .Z(n69700) );
  XOR U90077 ( .A(n70227), .B(n70228), .Z(n69699) );
  NOR U90078 ( .A(n69700), .B(n69699), .Z(n80349) );
  NOR U90079 ( .A(n69701), .B(n80349), .Z(n69702) );
  IV U90080 ( .A(n69702), .Z(n74943) );
  IV U90081 ( .A(n69703), .Z(n69705) );
  NOR U90082 ( .A(n69705), .B(n69704), .Z(n74941) );
  XOR U90083 ( .A(n74943), .B(n74941), .Z(n75556) );
  XOR U90084 ( .A(n74946), .B(n75556), .Z(n74948) );
  IV U90085 ( .A(n69706), .Z(n69708) );
  NOR U90086 ( .A(n69708), .B(n69707), .Z(n74947) );
  IV U90087 ( .A(n69709), .Z(n69710) );
  NOR U90088 ( .A(n69711), .B(n69710), .Z(n74952) );
  NOR U90089 ( .A(n74947), .B(n74952), .Z(n69712) );
  XOR U90090 ( .A(n74948), .B(n69712), .Z(n74959) );
  XOR U90091 ( .A(n69713), .B(n74959), .Z(n70215) );
  XOR U90092 ( .A(n69714), .B(n70215), .Z(n70214) );
  XOR U90093 ( .A(n70212), .B(n70214), .Z(n75528) );
  XOR U90094 ( .A(n70207), .B(n75528), .Z(n70208) );
  IV U90095 ( .A(n69715), .Z(n69719) );
  NOR U90096 ( .A(n69717), .B(n69716), .Z(n69718) );
  IV U90097 ( .A(n69718), .Z(n69722) );
  NOR U90098 ( .A(n69719), .B(n69722), .Z(n69720) );
  IV U90099 ( .A(n69720), .Z(n70209) );
  XOR U90100 ( .A(n70208), .B(n70209), .Z(n70203) );
  IV U90101 ( .A(n69721), .Z(n69723) );
  NOR U90102 ( .A(n69723), .B(n69722), .Z(n70201) );
  XOR U90103 ( .A(n70203), .B(n70201), .Z(n70205) );
  XOR U90104 ( .A(n70204), .B(n70205), .Z(n74966) );
  XOR U90105 ( .A(n74965), .B(n74966), .Z(n74972) );
  IV U90106 ( .A(n69724), .Z(n69725) );
  NOR U90107 ( .A(n69726), .B(n69725), .Z(n74968) );
  IV U90108 ( .A(n69727), .Z(n69729) );
  NOR U90109 ( .A(n69729), .B(n69728), .Z(n74971) );
  NOR U90110 ( .A(n74968), .B(n74971), .Z(n69730) );
  XOR U90111 ( .A(n74972), .B(n69730), .Z(n70198) );
  IV U90112 ( .A(n69731), .Z(n69733) );
  NOR U90113 ( .A(n69733), .B(n69732), .Z(n74975) );
  IV U90114 ( .A(n69734), .Z(n69735) );
  NOR U90115 ( .A(n69737), .B(n69735), .Z(n70199) );
  IV U90116 ( .A(n69736), .Z(n69738) );
  NOR U90117 ( .A(n69738), .B(n69737), .Z(n74979) );
  NOR U90118 ( .A(n70199), .B(n74979), .Z(n69739) );
  IV U90119 ( .A(n69739), .Z(n69740) );
  NOR U90120 ( .A(n74975), .B(n69740), .Z(n69741) );
  XOR U90121 ( .A(n70198), .B(n69741), .Z(n70193) );
  XOR U90122 ( .A(n70192), .B(n70193), .Z(n70197) );
  IV U90123 ( .A(n69742), .Z(n69743) );
  NOR U90124 ( .A(n69743), .B(n69745), .Z(n70195) );
  XOR U90125 ( .A(n70197), .B(n70195), .Z(n70191) );
  IV U90126 ( .A(n69744), .Z(n69746) );
  NOR U90127 ( .A(n69746), .B(n69745), .Z(n70189) );
  XOR U90128 ( .A(n70191), .B(n70189), .Z(n74989) );
  IV U90129 ( .A(n74989), .Z(n69751) );
  NOR U90130 ( .A(n69747), .B(n69751), .Z(n69760) );
  IV U90131 ( .A(n69752), .Z(n69748) );
  NOR U90132 ( .A(n69748), .B(n70197), .Z(n69749) );
  IV U90133 ( .A(n69749), .Z(n69750) );
  NOR U90134 ( .A(n69755), .B(n69750), .Z(n80382) );
  NOR U90135 ( .A(n69752), .B(n69751), .Z(n69758) );
  IV U90136 ( .A(n69753), .Z(n69754) );
  NOR U90137 ( .A(n69755), .B(n69754), .Z(n69756) );
  IV U90138 ( .A(n69756), .Z(n69757) );
  NOR U90139 ( .A(n69758), .B(n69757), .Z(n75499) );
  NOR U90140 ( .A(n80382), .B(n75499), .Z(n69759) );
  IV U90141 ( .A(n69759), .Z(n74990) );
  NOR U90142 ( .A(n69760), .B(n74990), .Z(n74995) );
  NOR U90143 ( .A(n69761), .B(n75496), .Z(n74987) );
  IV U90144 ( .A(n69762), .Z(n69763) );
  NOR U90145 ( .A(n69764), .B(n69763), .Z(n74994) );
  NOR U90146 ( .A(n74987), .B(n74994), .Z(n69765) );
  XOR U90147 ( .A(n74995), .B(n69765), .Z(n75002) );
  IV U90148 ( .A(n69766), .Z(n69767) );
  NOR U90149 ( .A(n69768), .B(n69767), .Z(n75000) );
  XOR U90150 ( .A(n75002), .B(n75000), .Z(n70187) );
  XOR U90151 ( .A(n70185), .B(n70187), .Z(n74998) );
  XOR U90152 ( .A(n69769), .B(n74998), .Z(n69770) );
  IV U90153 ( .A(n69770), .Z(n75009) );
  XOR U90154 ( .A(n75008), .B(n75009), .Z(n75014) );
  IV U90155 ( .A(n75014), .Z(n75017) );
  IV U90156 ( .A(n69771), .Z(n69773) );
  NOR U90157 ( .A(n69773), .B(n69772), .Z(n75015) );
  IV U90158 ( .A(n69774), .Z(n69776) );
  NOR U90159 ( .A(n69776), .B(n69775), .Z(n75013) );
  NOR U90160 ( .A(n75015), .B(n75013), .Z(n69777) );
  XOR U90161 ( .A(n75017), .B(n69777), .Z(n75030) );
  XOR U90162 ( .A(n69785), .B(n75030), .Z(n69778) );
  NOR U90163 ( .A(n69779), .B(n69778), .Z(n75476) );
  IV U90164 ( .A(n69780), .Z(n69782) );
  IV U90165 ( .A(n69781), .Z(n70172) );
  NOR U90166 ( .A(n69782), .B(n70172), .Z(n69787) );
  IV U90167 ( .A(n69783), .Z(n69784) );
  NOR U90168 ( .A(n70172), .B(n69784), .Z(n75029) );
  NOR U90169 ( .A(n69785), .B(n75029), .Z(n69786) );
  XOR U90170 ( .A(n69786), .B(n75030), .Z(n70165) );
  XOR U90171 ( .A(n69787), .B(n70165), .Z(n69788) );
  NOR U90172 ( .A(n69789), .B(n69788), .Z(n69790) );
  NOR U90173 ( .A(n75476), .B(n69790), .Z(n70162) );
  IV U90174 ( .A(n69791), .Z(n69793) );
  NOR U90175 ( .A(n69793), .B(n69792), .Z(n69794) );
  IV U90176 ( .A(n69794), .Z(n70164) );
  XOR U90177 ( .A(n70162), .B(n70164), .Z(n70160) );
  XOR U90178 ( .A(n70159), .B(n70160), .Z(n75046) );
  XOR U90179 ( .A(n75045), .B(n75046), .Z(n75049) );
  XOR U90180 ( .A(n69795), .B(n75049), .Z(n69796) );
  IV U90181 ( .A(n69796), .Z(n70153) );
  XOR U90182 ( .A(n70151), .B(n70153), .Z(n70155) );
  XOR U90183 ( .A(n70154), .B(n70155), .Z(n70144) );
  IV U90184 ( .A(n69797), .Z(n70148) );
  NOR U90185 ( .A(n69798), .B(n70148), .Z(n69802) );
  IV U90186 ( .A(n69799), .Z(n69801) );
  NOR U90187 ( .A(n69801), .B(n69800), .Z(n70143) );
  NOR U90188 ( .A(n69802), .B(n70143), .Z(n69803) );
  XOR U90189 ( .A(n70144), .B(n69803), .Z(n75056) );
  IV U90190 ( .A(n69804), .Z(n69816) );
  IV U90191 ( .A(n69805), .Z(n69806) );
  NOR U90192 ( .A(n69816), .B(n69806), .Z(n75064) );
  IV U90193 ( .A(n69807), .Z(n69808) );
  NOR U90194 ( .A(n69810), .B(n69808), .Z(n75058) );
  IV U90195 ( .A(n69809), .Z(n69811) );
  NOR U90196 ( .A(n69811), .B(n69810), .Z(n75059) );
  XOR U90197 ( .A(n75058), .B(n75059), .Z(n69812) );
  NOR U90198 ( .A(n75064), .B(n69812), .Z(n69813) );
  XOR U90199 ( .A(n75056), .B(n69813), .Z(n75068) );
  IV U90200 ( .A(n69814), .Z(n69815) );
  NOR U90201 ( .A(n69816), .B(n69815), .Z(n75067) );
  IV U90202 ( .A(n69817), .Z(n69822) );
  NOR U90203 ( .A(n69819), .B(n69818), .Z(n69820) );
  IV U90204 ( .A(n69820), .Z(n69821) );
  NOR U90205 ( .A(n69822), .B(n69821), .Z(n75062) );
  NOR U90206 ( .A(n75067), .B(n75062), .Z(n69823) );
  XOR U90207 ( .A(n75068), .B(n69823), .Z(n70141) );
  XOR U90208 ( .A(n70142), .B(n70141), .Z(n70136) );
  XOR U90209 ( .A(n70135), .B(n70136), .Z(n70140) );
  IV U90210 ( .A(n69824), .Z(n69828) );
  NOR U90211 ( .A(n69826), .B(n69825), .Z(n69827) );
  IV U90212 ( .A(n69827), .Z(n69830) );
  NOR U90213 ( .A(n69828), .B(n69830), .Z(n70138) );
  XOR U90214 ( .A(n70140), .B(n70138), .Z(n75090) );
  IV U90215 ( .A(n69829), .Z(n69831) );
  NOR U90216 ( .A(n69831), .B(n69830), .Z(n75088) );
  XOR U90217 ( .A(n75090), .B(n75088), .Z(n75091) );
  XOR U90218 ( .A(n75092), .B(n75091), .Z(n70127) );
  IV U90219 ( .A(n69832), .Z(n69834) );
  NOR U90220 ( .A(n69834), .B(n69833), .Z(n70126) );
  IV U90221 ( .A(n69835), .Z(n69836) );
  NOR U90222 ( .A(n69837), .B(n69836), .Z(n70132) );
  NOR U90223 ( .A(n70126), .B(n70132), .Z(n69838) );
  XOR U90224 ( .A(n70127), .B(n69838), .Z(n70130) );
  XOR U90225 ( .A(n70129), .B(n70130), .Z(n75097) );
  XOR U90226 ( .A(n75096), .B(n75097), .Z(n75100) );
  XOR U90227 ( .A(n75099), .B(n75100), .Z(n70120) );
  NOR U90228 ( .A(n69845), .B(n70120), .Z(n75443) );
  IV U90229 ( .A(n69839), .Z(n69841) );
  NOR U90230 ( .A(n69841), .B(n69840), .Z(n70122) );
  IV U90231 ( .A(n69842), .Z(n69844) );
  NOR U90232 ( .A(n69844), .B(n69843), .Z(n70119) );
  XOR U90233 ( .A(n70119), .B(n70120), .Z(n70123) );
  IV U90234 ( .A(n70123), .Z(n69846) );
  XOR U90235 ( .A(n70122), .B(n69846), .Z(n69848) );
  NOR U90236 ( .A(n69846), .B(n69845), .Z(n69847) );
  NOR U90237 ( .A(n69848), .B(n69847), .Z(n69849) );
  NOR U90238 ( .A(n75443), .B(n69849), .Z(n70116) );
  NOR U90239 ( .A(n69851), .B(n69850), .Z(n70115) );
  IV U90240 ( .A(n69852), .Z(n69854) );
  NOR U90241 ( .A(n69854), .B(n69853), .Z(n75105) );
  NOR U90242 ( .A(n70115), .B(n75105), .Z(n69855) );
  XOR U90243 ( .A(n70116), .B(n69855), .Z(n75110) );
  XOR U90244 ( .A(n75108), .B(n75110), .Z(n75427) );
  XOR U90245 ( .A(n70114), .B(n75427), .Z(n75116) );
  IV U90246 ( .A(n69856), .Z(n69857) );
  NOR U90247 ( .A(n69858), .B(n69857), .Z(n69859) );
  IV U90248 ( .A(n69859), .Z(n75117) );
  XOR U90249 ( .A(n75116), .B(n75117), .Z(n75128) );
  IV U90250 ( .A(n69860), .Z(n69861) );
  NOR U90251 ( .A(n69861), .B(n69866), .Z(n75124) );
  IV U90252 ( .A(n69862), .Z(n69863) );
  NOR U90253 ( .A(n69864), .B(n69863), .Z(n75112) );
  IV U90254 ( .A(n69865), .Z(n69867) );
  NOR U90255 ( .A(n69867), .B(n69866), .Z(n75127) );
  NOR U90256 ( .A(n75112), .B(n75127), .Z(n69868) );
  IV U90257 ( .A(n69868), .Z(n69869) );
  NOR U90258 ( .A(n75124), .B(n69869), .Z(n69870) );
  XOR U90259 ( .A(n75128), .B(n69870), .Z(n69873) );
  IV U90260 ( .A(n69873), .Z(n69872) );
  IV U90261 ( .A(n69874), .Z(n69871) );
  NOR U90262 ( .A(n69872), .B(n69871), .Z(n75132) );
  NOR U90263 ( .A(n69874), .B(n69873), .Z(n70112) );
  XOR U90264 ( .A(n70112), .B(n70110), .Z(n69875) );
  NOR U90265 ( .A(n75132), .B(n69875), .Z(n69876) );
  IV U90266 ( .A(n69876), .Z(n75141) );
  NOR U90267 ( .A(n69880), .B(n75141), .Z(n75414) );
  IV U90268 ( .A(n69877), .Z(n69879) );
  NOR U90269 ( .A(n69879), .B(n69878), .Z(n75144) );
  XOR U90270 ( .A(n75140), .B(n75141), .Z(n75145) );
  IV U90271 ( .A(n75145), .Z(n69881) );
  XOR U90272 ( .A(n75144), .B(n69881), .Z(n69883) );
  NOR U90273 ( .A(n69881), .B(n69880), .Z(n69882) );
  NOR U90274 ( .A(n69883), .B(n69882), .Z(n69884) );
  NOR U90275 ( .A(n75414), .B(n69884), .Z(n69885) );
  IV U90276 ( .A(n69885), .Z(n75152) );
  XOR U90277 ( .A(n75151), .B(n75152), .Z(n75156) );
  XOR U90278 ( .A(n75155), .B(n75156), .Z(n75160) );
  IV U90279 ( .A(n69886), .Z(n69888) );
  NOR U90280 ( .A(n69888), .B(n69887), .Z(n75158) );
  XOR U90281 ( .A(n75160), .B(n75158), .Z(n75164) );
  IV U90282 ( .A(n69889), .Z(n69893) );
  NOR U90283 ( .A(n69896), .B(n69890), .Z(n69891) );
  IV U90284 ( .A(n69891), .Z(n69892) );
  NOR U90285 ( .A(n69893), .B(n69892), .Z(n75162) );
  XOR U90286 ( .A(n75164), .B(n75162), .Z(n75167) );
  IV U90287 ( .A(n69894), .Z(n69899) );
  NOR U90288 ( .A(n69896), .B(n69895), .Z(n69897) );
  IV U90289 ( .A(n69897), .Z(n69898) );
  NOR U90290 ( .A(n69899), .B(n69898), .Z(n75165) );
  XOR U90291 ( .A(n75167), .B(n75165), .Z(n75171) );
  XOR U90292 ( .A(n75170), .B(n75171), .Z(n80472) );
  IV U90293 ( .A(n80472), .Z(n69906) );
  IV U90294 ( .A(n69900), .Z(n69902) );
  NOR U90295 ( .A(n69902), .B(n69901), .Z(n80475) );
  IV U90296 ( .A(n69903), .Z(n69905) );
  NOR U90297 ( .A(n69905), .B(n69904), .Z(n80470) );
  NOR U90298 ( .A(n80475), .B(n80470), .Z(n75173) );
  XOR U90299 ( .A(n69906), .B(n75173), .Z(n75179) );
  XOR U90300 ( .A(n75176), .B(n75179), .Z(n75188) );
  XOR U90301 ( .A(n69907), .B(n75188), .Z(n70108) );
  XOR U90302 ( .A(n69908), .B(n70108), .Z(n75199) );
  XOR U90303 ( .A(n75193), .B(n75199), .Z(n70106) );
  XOR U90304 ( .A(n69909), .B(n70106), .Z(n70099) );
  XOR U90305 ( .A(n69910), .B(n70099), .Z(n70095) );
  XOR U90306 ( .A(n69911), .B(n70095), .Z(n70088) );
  XOR U90307 ( .A(n70089), .B(n70088), .Z(n75206) );
  IV U90308 ( .A(n69912), .Z(n69913) );
  NOR U90309 ( .A(n69914), .B(n69913), .Z(n75202) );
  IV U90310 ( .A(n69915), .Z(n69917) );
  NOR U90311 ( .A(n69917), .B(n69916), .Z(n75204) );
  NOR U90312 ( .A(n75202), .B(n75204), .Z(n69918) );
  XOR U90313 ( .A(n75206), .B(n69918), .Z(n69919) );
  NOR U90314 ( .A(n69920), .B(n69919), .Z(n69923) );
  IV U90315 ( .A(n69920), .Z(n69922) );
  XOR U90316 ( .A(n75204), .B(n75206), .Z(n69921) );
  NOR U90317 ( .A(n69922), .B(n69921), .Z(n75382) );
  NOR U90318 ( .A(n69923), .B(n75382), .Z(n75208) );
  IV U90319 ( .A(n69924), .Z(n69938) );
  XOR U90320 ( .A(n69926), .B(n69925), .Z(n69927) );
  NOR U90321 ( .A(n69928), .B(n69927), .Z(n69929) );
  IV U90322 ( .A(n69929), .Z(n69935) );
  IV U90323 ( .A(n69930), .Z(n69932) );
  NOR U90324 ( .A(n69932), .B(n69931), .Z(n69933) );
  IV U90325 ( .A(n69933), .Z(n69934) );
  NOR U90326 ( .A(n69935), .B(n69934), .Z(n69936) );
  IV U90327 ( .A(n69936), .Z(n69937) );
  NOR U90328 ( .A(n69938), .B(n69937), .Z(n69939) );
  IV U90329 ( .A(n69939), .Z(n69940) );
  NOR U90330 ( .A(n69941), .B(n69940), .Z(n69942) );
  IV U90331 ( .A(n69942), .Z(n75209) );
  XOR U90332 ( .A(n75208), .B(n75209), .Z(n75213) );
  XOR U90333 ( .A(n75212), .B(n75213), .Z(n75216) );
  XOR U90334 ( .A(n75215), .B(n75216), .Z(n70083) );
  XOR U90335 ( .A(n70082), .B(n70083), .Z(n70086) );
  XOR U90336 ( .A(n70085), .B(n70086), .Z(n70078) );
  IV U90337 ( .A(n69943), .Z(n69945) );
  IV U90338 ( .A(n69944), .Z(n69951) );
  NOR U90339 ( .A(n69945), .B(n69951), .Z(n69946) );
  IV U90340 ( .A(n69946), .Z(n70077) );
  XOR U90341 ( .A(n70078), .B(n70077), .Z(n70079) );
  IV U90342 ( .A(n69947), .Z(n69948) );
  NOR U90343 ( .A(n69949), .B(n69948), .Z(n75224) );
  IV U90344 ( .A(n69950), .Z(n69952) );
  NOR U90345 ( .A(n69952), .B(n69951), .Z(n70080) );
  NOR U90346 ( .A(n75224), .B(n70080), .Z(n69953) );
  XOR U90347 ( .A(n70079), .B(n69953), .Z(n70075) );
  XOR U90348 ( .A(n70074), .B(n70075), .Z(n70072) );
  XOR U90349 ( .A(n69954), .B(n70072), .Z(n70069) );
  XOR U90350 ( .A(n70068), .B(n70069), .Z(n75237) );
  XOR U90351 ( .A(n75236), .B(n75237), .Z(n75241) );
  IV U90352 ( .A(n69955), .Z(n69956) );
  NOR U90353 ( .A(n69957), .B(n69956), .Z(n75239) );
  XOR U90354 ( .A(n75241), .B(n75239), .Z(n80756) );
  IV U90355 ( .A(n69958), .Z(n69959) );
  NOR U90356 ( .A(n69960), .B(n69959), .Z(n80759) );
  IV U90357 ( .A(n69961), .Z(n69963) );
  NOR U90358 ( .A(n69963), .B(n69962), .Z(n80751) );
  NOR U90359 ( .A(n80759), .B(n80751), .Z(n86472) );
  XOR U90360 ( .A(n80756), .B(n86472), .Z(n70063) );
  XOR U90361 ( .A(n69964), .B(n70063), .Z(n75350) );
  XOR U90362 ( .A(n69965), .B(n75350), .Z(n70058) );
  XOR U90363 ( .A(n70056), .B(n70058), .Z(n70061) );
  XOR U90364 ( .A(n70059), .B(n70061), .Z(n75251) );
  XOR U90365 ( .A(n75249), .B(n75251), .Z(n75253) );
  XOR U90366 ( .A(n75252), .B(n75253), .Z(n75259) );
  XOR U90367 ( .A(n75257), .B(n75259), .Z(n75262) );
  XOR U90368 ( .A(n75260), .B(n75262), .Z(n75273) );
  XOR U90369 ( .A(n69966), .B(n75273), .Z(n75269) );
  XOR U90370 ( .A(n69967), .B(n75269), .Z(n70052) );
  XOR U90371 ( .A(n70051), .B(n70052), .Z(n75281) );
  XOR U90372 ( .A(n75280), .B(n75281), .Z(n80704) );
  XOR U90373 ( .A(n70050), .B(n80704), .Z(n70049) );
  IV U90374 ( .A(n69968), .Z(n69969) );
  NOR U90375 ( .A(n69970), .B(n69969), .Z(n80584) );
  IV U90376 ( .A(n69971), .Z(n69973) );
  NOR U90377 ( .A(n69973), .B(n69972), .Z(n80580) );
  NOR U90378 ( .A(n80584), .B(n80580), .Z(n75297) );
  XOR U90379 ( .A(n70049), .B(n75297), .Z(n75300) );
  XOR U90380 ( .A(n75299), .B(n75300), .Z(n75303) );
  XOR U90381 ( .A(n75302), .B(n75303), .Z(n69974) );
  NOR U90382 ( .A(n69981), .B(n69974), .Z(n75344) );
  IV U90383 ( .A(n69975), .Z(n69976) );
  NOR U90384 ( .A(n69976), .B(n69986), .Z(n70041) );
  IV U90385 ( .A(n69977), .Z(n69979) );
  NOR U90386 ( .A(n69979), .B(n69978), .Z(n70047) );
  NOR U90387 ( .A(n75302), .B(n70047), .Z(n69980) );
  XOR U90388 ( .A(n69980), .B(n75303), .Z(n70042) );
  XOR U90389 ( .A(n70041), .B(n70042), .Z(n69983) );
  NOR U90390 ( .A(n70042), .B(n69981), .Z(n69982) );
  NOR U90391 ( .A(n69983), .B(n69982), .Z(n69984) );
  NOR U90392 ( .A(n75344), .B(n69984), .Z(n70045) );
  IV U90393 ( .A(n69985), .Z(n69987) );
  NOR U90394 ( .A(n69987), .B(n69986), .Z(n80598) );
  NOR U90395 ( .A(n69989), .B(n69988), .Z(n69990) );
  IV U90396 ( .A(n69990), .Z(n69996) );
  IV U90397 ( .A(n69991), .Z(n69992) );
  NOR U90398 ( .A(n69993), .B(n69992), .Z(n69994) );
  IV U90399 ( .A(n69994), .Z(n69995) );
  NOR U90400 ( .A(n69996), .B(n69995), .Z(n69997) );
  IV U90401 ( .A(n69997), .Z(n69998) );
  NOR U90402 ( .A(n69999), .B(n69998), .Z(n80616) );
  NOR U90403 ( .A(n80598), .B(n80616), .Z(n86337) );
  XOR U90404 ( .A(n70045), .B(n86337), .Z(n75312) );
  XOR U90405 ( .A(n70000), .B(n75312), .Z(n70038) );
  XOR U90406 ( .A(n70040), .B(n70038), .Z(n70033) );
  XOR U90407 ( .A(n70032), .B(n70033), .Z(n70037) );
  IV U90408 ( .A(n70001), .Z(n70002) );
  NOR U90409 ( .A(n70003), .B(n70002), .Z(n70035) );
  XOR U90410 ( .A(n70037), .B(n70035), .Z(n70027) );
  XOR U90411 ( .A(n70026), .B(n70027), .Z(n75335) );
  XOR U90412 ( .A(n70029), .B(n75335), .Z(n80642) );
  IV U90413 ( .A(n80642), .Z(n75332) );
  XOR U90414 ( .A(n70005), .B(n70004), .Z(n75318) );
  IV U90415 ( .A(n80645), .Z(n70008) );
  NOR U90416 ( .A(n70007), .B(n70006), .Z(n80646) );
  XOR U90417 ( .A(n70008), .B(n80646), .Z(n86386) );
  NOR U90418 ( .A(n70010), .B(n70009), .Z(n70011) );
  XOR U90419 ( .A(n70012), .B(n70011), .Z(n70013) );
  IV U90420 ( .A(n70013), .Z(n80647) );
  NOR U90421 ( .A(n86386), .B(n80647), .Z(n70014) );
  IV U90422 ( .A(n70014), .Z(n80651) );
  XOR U90423 ( .A(n70016), .B(n70015), .Z(n80652) );
  NOR U90424 ( .A(n80651), .B(n80652), .Z(n70017) );
  IV U90425 ( .A(n70017), .Z(n75324) );
  IV U90426 ( .A(n70018), .Z(n70020) );
  NOR U90427 ( .A(n70020), .B(n70019), .Z(n80650) );
  IV U90428 ( .A(n80650), .Z(n70021) );
  NOR U90429 ( .A(n75324), .B(n70021), .Z(n75325) );
  IV U90430 ( .A(n75325), .Z(n70022) );
  NOR U90431 ( .A(n70023), .B(n70022), .Z(n75319) );
  IV U90432 ( .A(n75319), .Z(n70024) );
  NOR U90433 ( .A(n75318), .B(n70024), .Z(n80640) );
  IV U90434 ( .A(n80640), .Z(n70025) );
  NOR U90435 ( .A(n75332), .B(n70025), .Z(n80664) );
  IV U90436 ( .A(n70026), .Z(n70028) );
  NOR U90437 ( .A(n70028), .B(n70027), .Z(n80635) );
  NOR U90438 ( .A(n70029), .B(n75335), .Z(n70030) );
  NOR U90439 ( .A(n80635), .B(n70030), .Z(n70031) );
  IV U90440 ( .A(n70031), .Z(n75317) );
  IV U90441 ( .A(n70032), .Z(n70034) );
  NOR U90442 ( .A(n70034), .B(n70033), .Z(n80628) );
  IV U90443 ( .A(n70035), .Z(n70036) );
  NOR U90444 ( .A(n70037), .B(n70036), .Z(n75339) );
  NOR U90445 ( .A(n80628), .B(n75339), .Z(n75316) );
  IV U90446 ( .A(n70038), .Z(n70039) );
  NOR U90447 ( .A(n70040), .B(n70039), .Z(n75314) );
  IV U90448 ( .A(n75314), .Z(n75307) );
  IV U90449 ( .A(n70041), .Z(n70044) );
  IV U90450 ( .A(n70042), .Z(n70043) );
  NOR U90451 ( .A(n70044), .B(n70043), .Z(n80604) );
  IV U90452 ( .A(n70045), .Z(n80600) );
  NOR U90453 ( .A(n86337), .B(n80600), .Z(n70046) );
  NOR U90454 ( .A(n80604), .B(n70046), .Z(n75306) );
  IV U90455 ( .A(n70047), .Z(n70048) );
  NOR U90456 ( .A(n70048), .B(n75303), .Z(n80593) );
  NOR U90457 ( .A(n80593), .B(n75344), .Z(n75305) );
  IV U90458 ( .A(n70049), .Z(n75295) );
  NOR U90459 ( .A(n75297), .B(n75295), .Z(n75292) );
  NOR U90460 ( .A(n70050), .B(n80704), .Z(n75289) );
  IV U90461 ( .A(n75289), .Z(n75286) );
  IV U90462 ( .A(n70051), .Z(n70053) );
  NOR U90463 ( .A(n70053), .B(n70052), .Z(n75346) );
  IV U90464 ( .A(n70054), .Z(n70055) );
  NOR U90465 ( .A(n75273), .B(n70055), .Z(n75265) );
  IV U90466 ( .A(n70056), .Z(n70057) );
  NOR U90467 ( .A(n70058), .B(n70057), .Z(n80733) );
  IV U90468 ( .A(n70059), .Z(n70060) );
  NOR U90469 ( .A(n70061), .B(n70060), .Z(n86287) );
  NOR U90470 ( .A(n80733), .B(n86287), .Z(n80546) );
  IV U90471 ( .A(n70062), .Z(n70064) );
  IV U90472 ( .A(n70063), .Z(n75245) );
  NOR U90473 ( .A(n70064), .B(n75245), .Z(n80533) );
  NOR U90474 ( .A(n75350), .B(n70065), .Z(n75247) );
  IV U90475 ( .A(n70066), .Z(n70067) );
  NOR U90476 ( .A(n70067), .B(n70072), .Z(n75368) );
  IV U90477 ( .A(n70068), .Z(n70070) );
  NOR U90478 ( .A(n70070), .B(n70069), .Z(n75364) );
  NOR U90479 ( .A(n75368), .B(n75364), .Z(n80769) );
  IV U90480 ( .A(n80769), .Z(n75235) );
  IV U90481 ( .A(n70071), .Z(n70073) );
  NOR U90482 ( .A(n70073), .B(n70072), .Z(n80770) );
  IV U90483 ( .A(n70074), .Z(n70076) );
  NOR U90484 ( .A(n70076), .B(n70075), .Z(n75232) );
  IV U90485 ( .A(n75232), .Z(n75223) );
  NOR U90486 ( .A(n70078), .B(n70077), .Z(n80519) );
  IV U90487 ( .A(n70079), .Z(n75225) );
  IV U90488 ( .A(n70080), .Z(n70081) );
  NOR U90489 ( .A(n75225), .B(n70081), .Z(n75370) );
  NOR U90490 ( .A(n80519), .B(n75370), .Z(n75221) );
  IV U90491 ( .A(n70082), .Z(n70084) );
  NOR U90492 ( .A(n70084), .B(n70083), .Z(n75372) );
  IV U90493 ( .A(n70085), .Z(n70087) );
  NOR U90494 ( .A(n70087), .B(n70086), .Z(n80522) );
  NOR U90495 ( .A(n75372), .B(n80522), .Z(n75219) );
  IV U90496 ( .A(n70088), .Z(n70090) );
  NOR U90497 ( .A(n70090), .B(n70089), .Z(n80506) );
  IV U90498 ( .A(n70091), .Z(n70092) );
  NOR U90499 ( .A(n70095), .B(n70092), .Z(n75391) );
  IV U90500 ( .A(n70093), .Z(n70094) );
  NOR U90501 ( .A(n70095), .B(n70094), .Z(n75385) );
  XOR U90502 ( .A(n75391), .B(n75385), .Z(n70096) );
  NOR U90503 ( .A(n80506), .B(n70096), .Z(n75201) );
  IV U90504 ( .A(n70097), .Z(n70101) );
  NOR U90505 ( .A(n70099), .B(n70098), .Z(n70100) );
  IV U90506 ( .A(n70100), .Z(n70103) );
  NOR U90507 ( .A(n70101), .B(n70103), .Z(n75388) );
  IV U90508 ( .A(n70102), .Z(n70104) );
  NOR U90509 ( .A(n70104), .B(n70103), .Z(n75396) );
  IV U90510 ( .A(n70105), .Z(n70107) );
  NOR U90511 ( .A(n70107), .B(n70106), .Z(n75393) );
  IV U90512 ( .A(n70108), .Z(n80496) );
  NOR U90513 ( .A(n70109), .B(n80496), .Z(n75192) );
  IV U90514 ( .A(n70110), .Z(n70111) );
  NOR U90515 ( .A(n70112), .B(n70111), .Z(n75134) );
  NOR U90516 ( .A(n75132), .B(n75134), .Z(n70113) );
  IV U90517 ( .A(n70113), .Z(n75131) );
  NOR U90518 ( .A(n70114), .B(n75427), .Z(n75119) );
  IV U90519 ( .A(n70115), .Z(n70117) );
  IV U90520 ( .A(n70116), .Z(n75106) );
  NOR U90521 ( .A(n70117), .B(n75106), .Z(n70118) );
  IV U90522 ( .A(n70118), .Z(n75440) );
  IV U90523 ( .A(n70119), .Z(n70121) );
  NOR U90524 ( .A(n70121), .B(n70120), .Z(n75445) );
  NOR U90525 ( .A(n75445), .B(n75443), .Z(n75104) );
  IV U90526 ( .A(n70122), .Z(n70124) );
  NOR U90527 ( .A(n70124), .B(n70123), .Z(n70125) );
  IV U90528 ( .A(n70125), .Z(n75442) );
  IV U90529 ( .A(n70126), .Z(n70128) );
  IV U90530 ( .A(n70127), .Z(n70134) );
  NOR U90531 ( .A(n70128), .B(n70134), .Z(n75450) );
  IV U90532 ( .A(n70129), .Z(n70131) );
  NOR U90533 ( .A(n70131), .B(n70130), .Z(n75453) );
  NOR U90534 ( .A(n75450), .B(n75453), .Z(n75095) );
  IV U90535 ( .A(n70132), .Z(n70133) );
  NOR U90536 ( .A(n70134), .B(n70133), .Z(n80429) );
  IV U90537 ( .A(n70135), .Z(n70137) );
  NOR U90538 ( .A(n70137), .B(n70136), .Z(n80890) );
  IV U90539 ( .A(n70138), .Z(n70139) );
  NOR U90540 ( .A(n70140), .B(n70139), .Z(n80883) );
  NOR U90541 ( .A(n80890), .B(n80883), .Z(n80424) );
  IV U90542 ( .A(n70141), .Z(n75081) );
  NOR U90543 ( .A(n70142), .B(n75081), .Z(n75071) );
  IV U90544 ( .A(n70143), .Z(n70145) );
  NOR U90545 ( .A(n70145), .B(n70144), .Z(n70146) );
  IV U90546 ( .A(n70146), .Z(n75464) );
  IV U90547 ( .A(n70147), .Z(n70150) );
  NOR U90548 ( .A(n70153), .B(n70148), .Z(n70149) );
  IV U90549 ( .A(n70149), .Z(n75054) );
  NOR U90550 ( .A(n70150), .B(n75054), .Z(n80414) );
  IV U90551 ( .A(n70151), .Z(n70152) );
  NOR U90552 ( .A(n70153), .B(n70152), .Z(n80406) );
  IV U90553 ( .A(n70154), .Z(n70156) );
  NOR U90554 ( .A(n70156), .B(n70155), .Z(n75468) );
  NOR U90555 ( .A(n80406), .B(n75468), .Z(n86116) );
  IV U90556 ( .A(n70157), .Z(n70158) );
  NOR U90557 ( .A(n75049), .B(n70158), .Z(n80404) );
  IV U90558 ( .A(n70159), .Z(n70161) );
  NOR U90559 ( .A(n70161), .B(n70160), .Z(n75473) );
  IV U90560 ( .A(n70162), .Z(n70163) );
  NOR U90561 ( .A(n70164), .B(n70163), .Z(n75470) );
  NOR U90562 ( .A(n75476), .B(n75470), .Z(n75044) );
  IV U90563 ( .A(n70165), .Z(n70167) );
  NOR U90564 ( .A(n70167), .B(n70166), .Z(n70168) );
  IV U90565 ( .A(n70168), .Z(n70175) );
  XOR U90566 ( .A(n70170), .B(n70169), .Z(n70171) );
  NOR U90567 ( .A(n70172), .B(n70171), .Z(n70173) );
  IV U90568 ( .A(n70173), .Z(n70174) );
  NOR U90569 ( .A(n70175), .B(n70174), .Z(n70176) );
  IV U90570 ( .A(n70176), .Z(n70177) );
  NOR U90571 ( .A(n70178), .B(n70177), .Z(n75040) );
  IV U90572 ( .A(n70179), .Z(n70180) );
  NOR U90573 ( .A(n70180), .B(n75014), .Z(n70181) );
  IV U90574 ( .A(n70181), .Z(n70182) );
  NOR U90575 ( .A(n75022), .B(n70182), .Z(n75033) );
  IV U90576 ( .A(n70183), .Z(n70184) );
  NOR U90577 ( .A(n70184), .B(n74998), .Z(n75488) );
  IV U90578 ( .A(n70185), .Z(n70186) );
  NOR U90579 ( .A(n70187), .B(n70186), .Z(n70188) );
  IV U90580 ( .A(n70188), .Z(n75003) );
  IV U90581 ( .A(n70189), .Z(n70190) );
  NOR U90582 ( .A(n70191), .B(n70190), .Z(n80376) );
  IV U90583 ( .A(n70192), .Z(n70194) );
  NOR U90584 ( .A(n70194), .B(n70193), .Z(n80372) );
  IV U90585 ( .A(n70195), .Z(n70196) );
  NOR U90586 ( .A(n70197), .B(n70196), .Z(n80378) );
  NOR U90587 ( .A(n80372), .B(n80378), .Z(n74986) );
  IV U90588 ( .A(n70198), .Z(n74981) );
  IV U90589 ( .A(n70199), .Z(n70200) );
  NOR U90590 ( .A(n74981), .B(n70200), .Z(n75505) );
  IV U90591 ( .A(n70201), .Z(n70202) );
  NOR U90592 ( .A(n70203), .B(n70202), .Z(n75522) );
  IV U90593 ( .A(n70204), .Z(n70206) );
  NOR U90594 ( .A(n70206), .B(n70205), .Z(n75512) );
  NOR U90595 ( .A(n75522), .B(n75512), .Z(n74964) );
  NOR U90596 ( .A(n70207), .B(n75528), .Z(n70211) );
  IV U90597 ( .A(n70208), .Z(n70210) );
  NOR U90598 ( .A(n70210), .B(n70209), .Z(n75525) );
  NOR U90599 ( .A(n70211), .B(n75525), .Z(n74963) );
  IV U90600 ( .A(n70212), .Z(n70213) );
  NOR U90601 ( .A(n70214), .B(n70213), .Z(n75537) );
  IV U90602 ( .A(n70215), .Z(n70220) );
  IV U90603 ( .A(n70216), .Z(n70217) );
  NOR U90604 ( .A(n70220), .B(n70217), .Z(n75535) );
  NOR U90605 ( .A(n75537), .B(n75535), .Z(n74961) );
  IV U90606 ( .A(n70218), .Z(n70219) );
  NOR U90607 ( .A(n70220), .B(n70219), .Z(n75544) );
  IV U90608 ( .A(n70221), .Z(n70222) );
  NOR U90609 ( .A(n70222), .B(n70228), .Z(n70223) );
  IV U90610 ( .A(n70223), .Z(n80348) );
  IV U90611 ( .A(n70224), .Z(n70226) );
  NOR U90612 ( .A(n70226), .B(n70225), .Z(n80342) );
  IV U90613 ( .A(n70227), .Z(n70229) );
  NOR U90614 ( .A(n70229), .B(n70228), .Z(n80344) );
  NOR U90615 ( .A(n80342), .B(n80344), .Z(n74940) );
  IV U90616 ( .A(n70230), .Z(n70232) );
  NOR U90617 ( .A(n70232), .B(n70231), .Z(n75568) );
  NOR U90618 ( .A(n70233), .B(n75565), .Z(n70234) );
  NOR U90619 ( .A(n75568), .B(n70234), .Z(n74939) );
  IV U90620 ( .A(n70235), .Z(n70236) );
  NOR U90621 ( .A(n70239), .B(n70236), .Z(n75581) );
  IV U90622 ( .A(n70237), .Z(n70238) );
  NOR U90623 ( .A(n70239), .B(n70238), .Z(n80332) );
  IV U90624 ( .A(n70240), .Z(n70241) );
  NOR U90625 ( .A(n70242), .B(n70241), .Z(n80329) );
  IV U90626 ( .A(n70243), .Z(n70247) );
  NOR U90627 ( .A(n70247), .B(n70244), .Z(n80322) );
  IV U90628 ( .A(n70245), .Z(n70246) );
  NOR U90629 ( .A(n70247), .B(n70246), .Z(n80326) );
  NOR U90630 ( .A(n80322), .B(n80326), .Z(n74933) );
  IV U90631 ( .A(n70248), .Z(n70249) );
  NOR U90632 ( .A(n70249), .B(n74932), .Z(n80320) );
  IV U90633 ( .A(n70250), .Z(n70251) );
  NOR U90634 ( .A(n70256), .B(n70251), .Z(n80296) );
  IV U90635 ( .A(n70252), .Z(n70253) );
  NOR U90636 ( .A(n70254), .B(n70253), .Z(n75595) );
  IV U90637 ( .A(n70255), .Z(n70257) );
  NOR U90638 ( .A(n70257), .B(n70256), .Z(n75592) );
  NOR U90639 ( .A(n75595), .B(n75592), .Z(n74905) );
  IV U90640 ( .A(n70258), .Z(n70259) );
  NOR U90641 ( .A(n70260), .B(n70259), .Z(n75599) );
  NOR U90642 ( .A(n75605), .B(n75599), .Z(n74904) );
  IV U90643 ( .A(n70261), .Z(n70262) );
  NOR U90644 ( .A(n70267), .B(n70262), .Z(n80287) );
  NOR U90645 ( .A(n70264), .B(n70263), .Z(n75602) );
  NOR U90646 ( .A(n80287), .B(n75602), .Z(n74903) );
  IV U90647 ( .A(n70265), .Z(n70266) );
  NOR U90648 ( .A(n70267), .B(n70266), .Z(n75611) );
  IV U90649 ( .A(n70268), .Z(n70270) );
  IV U90650 ( .A(n70269), .Z(n70272) );
  NOR U90651 ( .A(n70270), .B(n70272), .Z(n75608) );
  IV U90652 ( .A(n70271), .Z(n70273) );
  NOR U90653 ( .A(n70273), .B(n70272), .Z(n80275) );
  IV U90654 ( .A(n70274), .Z(n70275) );
  NOR U90655 ( .A(n70277), .B(n70275), .Z(n85983) );
  IV U90656 ( .A(n70276), .Z(n70278) );
  NOR U90657 ( .A(n70278), .B(n70277), .Z(n85963) );
  NOR U90658 ( .A(n85983), .B(n85963), .Z(n80280) );
  IV U90659 ( .A(n70279), .Z(n70280) );
  NOR U90660 ( .A(n70281), .B(n70280), .Z(n85975) );
  IV U90661 ( .A(n70282), .Z(n70284) );
  NOR U90662 ( .A(n70284), .B(n70283), .Z(n85969) );
  NOR U90663 ( .A(n85975), .B(n85969), .Z(n80274) );
  IV U90664 ( .A(n70285), .Z(n75625) );
  NOR U90665 ( .A(n70286), .B(n75625), .Z(n75614) );
  IV U90666 ( .A(n70287), .Z(n70288) );
  NOR U90667 ( .A(n70288), .B(n70293), .Z(n80261) );
  IV U90668 ( .A(n70289), .Z(n70290) );
  NOR U90669 ( .A(n70291), .B(n70290), .Z(n80257) );
  IV U90670 ( .A(n70292), .Z(n70294) );
  NOR U90671 ( .A(n70294), .B(n70293), .Z(n75636) );
  NOR U90672 ( .A(n80257), .B(n75636), .Z(n74892) );
  IV U90673 ( .A(n70295), .Z(n70296) );
  NOR U90674 ( .A(n70297), .B(n70296), .Z(n74891) );
  IV U90675 ( .A(n74891), .Z(n74889) );
  IV U90676 ( .A(n70298), .Z(n70299) );
  NOR U90677 ( .A(n70300), .B(n70299), .Z(n75643) );
  IV U90678 ( .A(n70301), .Z(n70302) );
  NOR U90679 ( .A(n70303), .B(n70302), .Z(n75641) );
  NOR U90680 ( .A(n75643), .B(n75641), .Z(n74887) );
  IV U90681 ( .A(n70304), .Z(n70305) );
  NOR U90682 ( .A(n70306), .B(n70305), .Z(n75646) );
  IV U90683 ( .A(n70307), .Z(n70308) );
  NOR U90684 ( .A(n70309), .B(n70308), .Z(n80254) );
  NOR U90685 ( .A(n75646), .B(n80254), .Z(n74885) );
  IV U90686 ( .A(n70310), .Z(n70312) );
  IV U90687 ( .A(n70311), .Z(n74883) );
  NOR U90688 ( .A(n70312), .B(n74883), .Z(n75652) );
  IV U90689 ( .A(n70313), .Z(n70314) );
  NOR U90690 ( .A(n70314), .B(n74879), .Z(n81092) );
  IV U90691 ( .A(n70315), .Z(n70316) );
  NOR U90692 ( .A(n70319), .B(n70316), .Z(n85937) );
  NOR U90693 ( .A(n81092), .B(n85937), .Z(n75658) );
  IV U90694 ( .A(n70317), .Z(n70318) );
  NOR U90695 ( .A(n70319), .B(n70318), .Z(n75666) );
  IV U90696 ( .A(n70320), .Z(n70325) );
  IV U90697 ( .A(n70321), .Z(n70322) );
  NOR U90698 ( .A(n70325), .B(n70322), .Z(n75676) );
  IV U90699 ( .A(n70323), .Z(n70324) );
  NOR U90700 ( .A(n70325), .B(n70324), .Z(n75673) );
  IV U90701 ( .A(n70326), .Z(n70328) );
  NOR U90702 ( .A(n70328), .B(n70327), .Z(n80234) );
  IV U90703 ( .A(n70329), .Z(n70330) );
  NOR U90704 ( .A(n70333), .B(n70330), .Z(n74844) );
  IV U90705 ( .A(n70331), .Z(n70332) );
  NOR U90706 ( .A(n70333), .B(n70332), .Z(n74842) );
  IV U90707 ( .A(n74842), .Z(n74834) );
  NOR U90708 ( .A(n70334), .B(n70338), .Z(n70335) );
  IV U90709 ( .A(n70335), .Z(n80224) );
  NOR U90710 ( .A(n70336), .B(n80224), .Z(n74838) );
  IV U90711 ( .A(n70337), .Z(n70339) );
  NOR U90712 ( .A(n70339), .B(n70338), .Z(n74831) );
  IV U90713 ( .A(n74831), .Z(n74820) );
  IV U90714 ( .A(n70340), .Z(n70341) );
  NOR U90715 ( .A(n70341), .B(n74826), .Z(n80213) );
  IV U90716 ( .A(n70342), .Z(n70343) );
  NOR U90717 ( .A(n70344), .B(n70343), .Z(n74805) );
  IV U90718 ( .A(n74805), .Z(n74800) );
  IV U90719 ( .A(n70345), .Z(n70347) );
  NOR U90720 ( .A(n70347), .B(n70346), .Z(n70348) );
  IV U90721 ( .A(n70348), .Z(n75695) );
  IV U90722 ( .A(n70349), .Z(n70350) );
  NOR U90723 ( .A(n70351), .B(n70350), .Z(n70355) );
  NOR U90724 ( .A(n70353), .B(n70352), .Z(n70354) );
  NOR U90725 ( .A(n70355), .B(n70354), .Z(n75705) );
  IV U90726 ( .A(n70356), .Z(n70360) );
  NOR U90727 ( .A(n70358), .B(n70357), .Z(n70359) );
  IV U90728 ( .A(n70359), .Z(n70362) );
  NOR U90729 ( .A(n70360), .B(n70362), .Z(n80184) );
  IV U90730 ( .A(n70361), .Z(n70363) );
  NOR U90731 ( .A(n70363), .B(n70362), .Z(n75709) );
  IV U90732 ( .A(n70364), .Z(n70365) );
  NOR U90733 ( .A(n70365), .B(n74784), .Z(n75706) );
  IV U90734 ( .A(n70366), .Z(n70368) );
  NOR U90735 ( .A(n70368), .B(n70367), .Z(n70369) );
  IV U90736 ( .A(n70369), .Z(n80175) );
  IV U90737 ( .A(n70370), .Z(n70371) );
  NOR U90738 ( .A(n70371), .B(n74775), .Z(n75719) );
  NOR U90739 ( .A(n75724), .B(n75719), .Z(n74773) );
  IV U90740 ( .A(n70372), .Z(n70373) );
  NOR U90741 ( .A(n70373), .B(n70379), .Z(n70374) );
  IV U90742 ( .A(n70374), .Z(n80163) );
  IV U90743 ( .A(n70375), .Z(n70377) );
  NOR U90744 ( .A(n70377), .B(n70376), .Z(n75730) );
  IV U90745 ( .A(n70378), .Z(n70380) );
  NOR U90746 ( .A(n70380), .B(n70379), .Z(n80165) );
  NOR U90747 ( .A(n75730), .B(n80165), .Z(n74767) );
  IV U90748 ( .A(n70381), .Z(n70383) );
  NOR U90749 ( .A(n70383), .B(n70382), .Z(n70384) );
  IV U90750 ( .A(n70384), .Z(n75732) );
  IV U90751 ( .A(n70385), .Z(n70387) );
  IV U90752 ( .A(n70386), .Z(n74751) );
  NOR U90753 ( .A(n70387), .B(n74751), .Z(n74754) );
  IV U90754 ( .A(n74754), .Z(n74749) );
  IV U90755 ( .A(n70388), .Z(n70390) );
  NOR U90756 ( .A(n70390), .B(n70389), .Z(n74718) );
  IV U90757 ( .A(n74718), .Z(n74712) );
  IV U90758 ( .A(n70391), .Z(n70393) );
  NOR U90759 ( .A(n70393), .B(n70392), .Z(n80133) );
  IV U90760 ( .A(n70394), .Z(n70395) );
  NOR U90761 ( .A(n74705), .B(n70395), .Z(n75764) );
  IV U90762 ( .A(n70396), .Z(n70397) );
  NOR U90763 ( .A(n70397), .B(n74700), .Z(n75769) );
  IV U90764 ( .A(n70398), .Z(n70399) );
  NOR U90765 ( .A(n70400), .B(n70399), .Z(n75761) );
  NOR U90766 ( .A(n75769), .B(n75761), .Z(n74703) );
  IV U90767 ( .A(n70401), .Z(n74698) );
  IV U90768 ( .A(n70402), .Z(n70403) );
  NOR U90769 ( .A(n74698), .B(n70403), .Z(n75772) );
  IV U90770 ( .A(n70404), .Z(n70405) );
  NOR U90771 ( .A(n70405), .B(n70407), .Z(n75778) );
  IV U90772 ( .A(n70406), .Z(n70408) );
  NOR U90773 ( .A(n70408), .B(n70407), .Z(n75776) );
  NOR U90774 ( .A(n75778), .B(n75776), .Z(n74692) );
  IV U90775 ( .A(n70409), .Z(n70410) );
  NOR U90776 ( .A(n70411), .B(n70410), .Z(n70412) );
  IV U90777 ( .A(n70412), .Z(n80113) );
  IV U90778 ( .A(n70413), .Z(n70415) );
  IV U90779 ( .A(n70414), .Z(n70417) );
  NOR U90780 ( .A(n70415), .B(n70417), .Z(n80109) );
  IV U90781 ( .A(n70416), .Z(n70418) );
  NOR U90782 ( .A(n70418), .B(n70417), .Z(n80101) );
  IV U90783 ( .A(n70419), .Z(n70420) );
  NOR U90784 ( .A(n70420), .B(n70424), .Z(n85802) );
  IV U90785 ( .A(n70421), .Z(n70422) );
  NOR U90786 ( .A(n70422), .B(n70429), .Z(n85798) );
  IV U90787 ( .A(n70423), .Z(n70425) );
  NOR U90788 ( .A(n70425), .B(n70424), .Z(n85803) );
  NOR U90789 ( .A(n85798), .B(n85803), .Z(n70426) );
  IV U90790 ( .A(n70426), .Z(n70427) );
  NOR U90791 ( .A(n85802), .B(n70427), .Z(n74689) );
  IV U90792 ( .A(n70428), .Z(n70430) );
  NOR U90793 ( .A(n70430), .B(n70429), .Z(n80092) );
  IV U90794 ( .A(n70431), .Z(n70432) );
  NOR U90795 ( .A(n70433), .B(n70432), .Z(n81241) );
  IV U90796 ( .A(n70434), .Z(n70435) );
  NOR U90797 ( .A(n70436), .B(n70435), .Z(n81233) );
  NOR U90798 ( .A(n81241), .B(n81233), .Z(n75786) );
  IV U90799 ( .A(n75786), .Z(n74679) );
  NOR U90800 ( .A(n70438), .B(n70437), .Z(n74661) );
  IV U90801 ( .A(n70439), .Z(n70440) );
  NOR U90802 ( .A(n70441), .B(n70440), .Z(n80056) );
  IV U90803 ( .A(n70442), .Z(n75792) );
  NOR U90804 ( .A(n70443), .B(n75792), .Z(n70444) );
  NOR U90805 ( .A(n75795), .B(n70444), .Z(n74637) );
  IV U90806 ( .A(n70445), .Z(n70446) );
  NOR U90807 ( .A(n70446), .B(n70448), .Z(n85761) );
  IV U90808 ( .A(n70447), .Z(n70449) );
  NOR U90809 ( .A(n70449), .B(n70448), .Z(n85768) );
  NOR U90810 ( .A(n85761), .B(n85768), .Z(n80045) );
  IV U90811 ( .A(n70450), .Z(n74631) );
  IV U90812 ( .A(n70451), .Z(n70452) );
  NOR U90813 ( .A(n74631), .B(n70452), .Z(n75801) );
  IV U90814 ( .A(n70453), .Z(n70454) );
  NOR U90815 ( .A(n70455), .B(n70454), .Z(n75798) );
  NOR U90816 ( .A(n75801), .B(n75798), .Z(n74636) );
  IV U90817 ( .A(n70456), .Z(n70458) );
  NOR U90818 ( .A(n70458), .B(n70457), .Z(n70459) );
  IV U90819 ( .A(n70459), .Z(n75809) );
  IV U90820 ( .A(n70460), .Z(n70461) );
  NOR U90821 ( .A(n70469), .B(n70461), .Z(n75812) );
  IV U90822 ( .A(n70462), .Z(n70463) );
  NOR U90823 ( .A(n70464), .B(n70463), .Z(n75806) );
  NOR U90824 ( .A(n75812), .B(n75806), .Z(n74609) );
  IV U90825 ( .A(n70465), .Z(n70473) );
  IV U90826 ( .A(n70466), .Z(n70467) );
  NOR U90827 ( .A(n70473), .B(n70467), .Z(n81281) );
  IV U90828 ( .A(n70468), .Z(n70470) );
  NOR U90829 ( .A(n70470), .B(n70469), .Z(n85733) );
  NOR U90830 ( .A(n81281), .B(n85733), .Z(n75811) );
  IV U90831 ( .A(n70471), .Z(n70472) );
  NOR U90832 ( .A(n70473), .B(n70472), .Z(n75816) );
  IV U90833 ( .A(n70474), .Z(n70475) );
  NOR U90834 ( .A(n70476), .B(n70475), .Z(n80011) );
  NOR U90835 ( .A(n75816), .B(n80011), .Z(n74608) );
  IV U90836 ( .A(n70477), .Z(n70478) );
  NOR U90837 ( .A(n70478), .B(n70480), .Z(n80018) );
  IV U90838 ( .A(n70479), .Z(n70481) );
  NOR U90839 ( .A(n70481), .B(n70480), .Z(n80016) );
  NOR U90840 ( .A(n80018), .B(n80016), .Z(n74607) );
  IV U90841 ( .A(n70482), .Z(n70483) );
  NOR U90842 ( .A(n70488), .B(n70483), .Z(n75829) );
  IV U90843 ( .A(n70484), .Z(n70485) );
  NOR U90844 ( .A(n70485), .B(n75819), .Z(n70486) );
  NOR U90845 ( .A(n75829), .B(n70486), .Z(n74606) );
  IV U90846 ( .A(n70487), .Z(n70489) );
  NOR U90847 ( .A(n70489), .B(n70488), .Z(n80003) );
  IV U90848 ( .A(n70490), .Z(n70491) );
  NOR U90849 ( .A(n70492), .B(n70491), .Z(n80000) );
  IV U90850 ( .A(n70493), .Z(n70494) );
  NOR U90851 ( .A(n70494), .B(n74586), .Z(n75836) );
  NOR U90852 ( .A(n80000), .B(n75836), .Z(n74590) );
  IV U90853 ( .A(n70495), .Z(n75846) );
  NOR U90854 ( .A(n70496), .B(n75846), .Z(n74577) );
  IV U90855 ( .A(n70497), .Z(n70498) );
  NOR U90856 ( .A(n70508), .B(n70498), .Z(n70499) );
  IV U90857 ( .A(n70499), .Z(n79978) );
  IV U90858 ( .A(n70500), .Z(n70501) );
  NOR U90859 ( .A(n70502), .B(n70501), .Z(n79963) );
  IV U90860 ( .A(n70503), .Z(n70505) );
  NOR U90861 ( .A(n70505), .B(n70504), .Z(n79979) );
  NOR U90862 ( .A(n79963), .B(n79979), .Z(n74527) );
  IV U90863 ( .A(n70506), .Z(n70507) );
  NOR U90864 ( .A(n70508), .B(n70507), .Z(n79968) );
  IV U90865 ( .A(n70509), .Z(n70511) );
  NOR U90866 ( .A(n70511), .B(n70510), .Z(n81357) );
  IV U90867 ( .A(n70512), .Z(n70514) );
  NOR U90868 ( .A(n70514), .B(n70513), .Z(n81353) );
  NOR U90869 ( .A(n81357), .B(n81353), .Z(n79967) );
  IV U90870 ( .A(n70515), .Z(n70519) );
  NOR U90871 ( .A(n70529), .B(n70516), .Z(n70517) );
  IV U90872 ( .A(n70517), .Z(n70518) );
  NOR U90873 ( .A(n70519), .B(n70518), .Z(n79959) );
  IV U90874 ( .A(n70520), .Z(n70521) );
  NOR U90875 ( .A(n70522), .B(n70521), .Z(n79957) );
  IV U90876 ( .A(n70523), .Z(n70525) );
  NOR U90877 ( .A(n70525), .B(n70524), .Z(n79955) );
  NOR U90878 ( .A(n79957), .B(n79955), .Z(n70526) );
  IV U90879 ( .A(n70526), .Z(n70527) );
  NOR U90880 ( .A(n79959), .B(n70527), .Z(n74526) );
  IV U90881 ( .A(n70528), .Z(n75896) );
  NOR U90882 ( .A(n70529), .B(n75896), .Z(n70530) );
  NOR U90883 ( .A(n79949), .B(n70530), .Z(n70531) );
  NOR U90884 ( .A(n70531), .B(n79950), .Z(n74525) );
  IV U90885 ( .A(n70532), .Z(n70533) );
  NOR U90886 ( .A(n70538), .B(n70533), .Z(n79937) );
  IV U90887 ( .A(n70534), .Z(n70536) );
  NOR U90888 ( .A(n70536), .B(n70535), .Z(n79928) );
  IV U90889 ( .A(n70537), .Z(n70539) );
  NOR U90890 ( .A(n70539), .B(n70538), .Z(n79923) );
  NOR U90891 ( .A(n79928), .B(n79923), .Z(n74517) );
  IV U90892 ( .A(n70540), .Z(n70541) );
  NOR U90893 ( .A(n70542), .B(n70541), .Z(n79916) );
  IV U90894 ( .A(n70543), .Z(n70544) );
  NOR U90895 ( .A(n70545), .B(n70544), .Z(n75907) );
  NOR U90896 ( .A(n79916), .B(n75907), .Z(n74516) );
  IV U90897 ( .A(n70546), .Z(n75910) );
  NOR U90898 ( .A(n75910), .B(n70547), .Z(n70551) );
  IV U90899 ( .A(n70548), .Z(n70550) );
  NOR U90900 ( .A(n70550), .B(n70549), .Z(n79919) );
  NOR U90901 ( .A(n70551), .B(n79919), .Z(n74515) );
  IV U90902 ( .A(n70552), .Z(n70555) );
  NOR U90903 ( .A(n70553), .B(n74504), .Z(n70554) );
  IV U90904 ( .A(n70554), .Z(n74510) );
  NOR U90905 ( .A(n70555), .B(n74510), .Z(n70556) );
  IV U90906 ( .A(n70556), .Z(n75914) );
  NOR U90907 ( .A(n70557), .B(n79893), .Z(n74502) );
  IV U90908 ( .A(n70558), .Z(n70562) );
  XOR U90909 ( .A(n70569), .B(n70570), .Z(n70559) );
  NOR U90910 ( .A(n70560), .B(n70559), .Z(n70561) );
  IV U90911 ( .A(n70561), .Z(n74496) );
  NOR U90912 ( .A(n70562), .B(n74496), .Z(n79880) );
  IV U90913 ( .A(n70563), .Z(n70564) );
  NOR U90914 ( .A(n70564), .B(n70570), .Z(n70565) );
  IV U90915 ( .A(n70565), .Z(n79878) );
  IV U90916 ( .A(n70566), .Z(n70567) );
  NOR U90917 ( .A(n70568), .B(n70567), .Z(n75927) );
  IV U90918 ( .A(n70569), .Z(n70571) );
  NOR U90919 ( .A(n70571), .B(n70570), .Z(n79874) );
  NOR U90920 ( .A(n75927), .B(n79874), .Z(n74494) );
  IV U90921 ( .A(n70572), .Z(n70573) );
  NOR U90922 ( .A(n70574), .B(n70573), .Z(n75930) );
  IV U90923 ( .A(n70575), .Z(n70577) );
  NOR U90924 ( .A(n70577), .B(n70576), .Z(n75939) );
  IV U90925 ( .A(n70578), .Z(n70580) );
  NOR U90926 ( .A(n70580), .B(n70579), .Z(n75936) );
  NOR U90927 ( .A(n75939), .B(n75936), .Z(n74487) );
  IV U90928 ( .A(n70581), .Z(n70583) );
  NOR U90929 ( .A(n70583), .B(n70582), .Z(n75941) );
  IV U90930 ( .A(n70584), .Z(n70586) );
  NOR U90931 ( .A(n70586), .B(n70585), .Z(n70591) );
  IV U90932 ( .A(n70587), .Z(n70589) );
  NOR U90933 ( .A(n70589), .B(n70588), .Z(n70590) );
  NOR U90934 ( .A(n70591), .B(n70590), .Z(n79863) );
  IV U90935 ( .A(n70592), .Z(n70594) );
  NOR U90936 ( .A(n70594), .B(n70593), .Z(n75945) );
  IV U90937 ( .A(n70595), .Z(n70597) );
  NOR U90938 ( .A(n70597), .B(n70596), .Z(n79865) );
  NOR U90939 ( .A(n75945), .B(n79865), .Z(n74486) );
  IV U90940 ( .A(n70598), .Z(n70600) );
  NOR U90941 ( .A(n70600), .B(n70599), .Z(n75948) );
  IV U90942 ( .A(n70601), .Z(n70602) );
  NOR U90943 ( .A(n70603), .B(n70602), .Z(n75965) );
  IV U90944 ( .A(n70604), .Z(n70605) );
  NOR U90945 ( .A(n74482), .B(n70605), .Z(n75957) );
  NOR U90946 ( .A(n75965), .B(n75957), .Z(n74479) );
  IV U90947 ( .A(n70606), .Z(n70608) );
  IV U90948 ( .A(n70607), .Z(n74474) );
  NOR U90949 ( .A(n70608), .B(n74474), .Z(n75962) );
  IV U90950 ( .A(n70609), .Z(n70610) );
  NOR U90951 ( .A(n70610), .B(n74472), .Z(n70611) );
  IV U90952 ( .A(n70611), .Z(n74469) );
  IV U90953 ( .A(n70612), .Z(n70613) );
  NOR U90954 ( .A(n79846), .B(n70613), .Z(n79842) );
  IV U90955 ( .A(n70614), .Z(n70615) );
  NOR U90956 ( .A(n79846), .B(n70615), .Z(n75976) );
  IV U90957 ( .A(n70616), .Z(n70623) );
  NOR U90958 ( .A(n70618), .B(n70617), .Z(n70619) );
  IV U90959 ( .A(n70619), .Z(n70620) );
  NOR U90960 ( .A(n70621), .B(n70620), .Z(n70622) );
  IV U90961 ( .A(n70622), .Z(n70625) );
  NOR U90962 ( .A(n70623), .B(n70625), .Z(n75973) );
  IV U90963 ( .A(n70624), .Z(n70626) );
  NOR U90964 ( .A(n70626), .B(n70625), .Z(n79837) );
  IV U90965 ( .A(n70627), .Z(n70629) );
  NOR U90966 ( .A(n70629), .B(n70628), .Z(n79834) );
  IV U90967 ( .A(n70630), .Z(n70631) );
  NOR U90968 ( .A(n70631), .B(n70633), .Z(n75984) );
  IV U90969 ( .A(n70632), .Z(n70634) );
  NOR U90970 ( .A(n70634), .B(n70633), .Z(n75982) );
  NOR U90971 ( .A(n75984), .B(n75982), .Z(n74468) );
  IV U90972 ( .A(n70635), .Z(n70637) );
  NOR U90973 ( .A(n70637), .B(n70636), .Z(n75989) );
  IV U90974 ( .A(n70638), .Z(n70639) );
  NOR U90975 ( .A(n70640), .B(n70639), .Z(n75987) );
  NOR U90976 ( .A(n75989), .B(n75987), .Z(n74467) );
  IV U90977 ( .A(n70641), .Z(n70643) );
  IV U90978 ( .A(n70642), .Z(n74464) );
  NOR U90979 ( .A(n70643), .B(n74464), .Z(n75992) );
  NOR U90980 ( .A(n70644), .B(n85590), .Z(n76020) );
  IV U90981 ( .A(n70645), .Z(n70647) );
  NOR U90982 ( .A(n70647), .B(n70646), .Z(n76011) );
  NOR U90983 ( .A(n76020), .B(n76011), .Z(n74447) );
  IV U90984 ( .A(n70648), .Z(n70651) );
  NOR U90985 ( .A(n70649), .B(n74432), .Z(n70650) );
  IV U90986 ( .A(n70650), .Z(n74424) );
  NOR U90987 ( .A(n70651), .B(n74424), .Z(n70652) );
  IV U90988 ( .A(n70652), .Z(n79813) );
  IV U90989 ( .A(n70653), .Z(n70654) );
  NOR U90990 ( .A(n70655), .B(n70654), .Z(n76033) );
  NOR U90991 ( .A(n85543), .B(n85552), .Z(n70656) );
  NOR U90992 ( .A(n70656), .B(n85544), .Z(n70657) );
  IV U90993 ( .A(n70657), .Z(n76039) );
  IV U90994 ( .A(n70658), .Z(n70659) );
  NOR U90995 ( .A(n70660), .B(n70659), .Z(n76042) );
  IV U90996 ( .A(n70661), .Z(n70663) );
  NOR U90997 ( .A(n70663), .B(n70662), .Z(n76040) );
  NOR U90998 ( .A(n76042), .B(n76040), .Z(n74419) );
  IV U90999 ( .A(n70664), .Z(n70665) );
  NOR U91000 ( .A(n70666), .B(n70665), .Z(n70667) );
  IV U91001 ( .A(n70667), .Z(n74393) );
  NOR U91002 ( .A(n70668), .B(n76049), .Z(n74380) );
  IV U91003 ( .A(n70669), .Z(n70671) );
  NOR U91004 ( .A(n70671), .B(n70670), .Z(n74377) );
  IV U91005 ( .A(n74377), .Z(n74373) );
  IV U91006 ( .A(n70672), .Z(n70674) );
  NOR U91007 ( .A(n70674), .B(n70673), .Z(n74361) );
  IV U91008 ( .A(n70675), .Z(n70676) );
  NOR U91009 ( .A(n70676), .B(n74372), .Z(n74363) );
  IV U91010 ( .A(n70677), .Z(n70678) );
  NOR U91011 ( .A(n70678), .B(n70686), .Z(n79738) );
  IV U91012 ( .A(n70679), .Z(n70681) );
  IV U91013 ( .A(n70680), .Z(n79744) );
  NOR U91014 ( .A(n70681), .B(n79744), .Z(n79736) );
  NOR U91015 ( .A(n79738), .B(n79736), .Z(n74352) );
  IV U91016 ( .A(n70682), .Z(n70683) );
  NOR U91017 ( .A(n70684), .B(n70683), .Z(n85534) );
  IV U91018 ( .A(n70685), .Z(n70687) );
  NOR U91019 ( .A(n70687), .B(n70686), .Z(n81565) );
  NOR U91020 ( .A(n85534), .B(n81565), .Z(n76076) );
  IV U91021 ( .A(n70688), .Z(n70689) );
  NOR U91022 ( .A(n70689), .B(n70690), .Z(n76078) );
  NOR U91023 ( .A(n70691), .B(n70690), .Z(n74346) );
  IV U91024 ( .A(n74346), .Z(n74340) );
  IV U91025 ( .A(n70692), .Z(n70694) );
  NOR U91026 ( .A(n70694), .B(n70693), .Z(n76083) );
  IV U91027 ( .A(n70695), .Z(n70697) );
  NOR U91028 ( .A(n70697), .B(n70696), .Z(n76086) );
  IV U91029 ( .A(n70698), .Z(n70699) );
  NOR U91030 ( .A(n70699), .B(n70701), .Z(n76125) );
  IV U91031 ( .A(n70700), .Z(n70702) );
  NOR U91032 ( .A(n70702), .B(n70701), .Z(n76133) );
  IV U91033 ( .A(n70703), .Z(n70705) );
  IV U91034 ( .A(n70704), .Z(n70711) );
  NOR U91035 ( .A(n70705), .B(n70711), .Z(n76157) );
  IV U91036 ( .A(n70706), .Z(n70708) );
  NOR U91037 ( .A(n70708), .B(n70707), .Z(n76154) );
  NOR U91038 ( .A(n76157), .B(n76154), .Z(n74251) );
  NOR U91039 ( .A(n70709), .B(n85470), .Z(n76162) );
  IV U91040 ( .A(n70710), .Z(n70712) );
  NOR U91041 ( .A(n70712), .B(n70711), .Z(n76160) );
  NOR U91042 ( .A(n76162), .B(n76160), .Z(n74250) );
  NOR U91043 ( .A(n70713), .B(n76167), .Z(n70717) );
  IV U91044 ( .A(n70714), .Z(n70716) );
  NOR U91045 ( .A(n70716), .B(n70715), .Z(n79680) );
  NOR U91046 ( .A(n70717), .B(n79680), .Z(n74249) );
  IV U91047 ( .A(n70718), .Z(n70720) );
  NOR U91048 ( .A(n70720), .B(n70719), .Z(n74247) );
  IV U91049 ( .A(n74247), .Z(n74239) );
  IV U91050 ( .A(n70721), .Z(n70723) );
  NOR U91051 ( .A(n70723), .B(n70722), .Z(n70724) );
  IV U91052 ( .A(n70724), .Z(n74212) );
  IV U91053 ( .A(n70725), .Z(n70728) );
  NOR U91054 ( .A(n70726), .B(n74205), .Z(n70727) );
  IV U91055 ( .A(n70727), .Z(n74200) );
  NOR U91056 ( .A(n70728), .B(n74200), .Z(n74194) );
  IV U91057 ( .A(n70729), .Z(n70730) );
  NOR U91058 ( .A(n70731), .B(n70730), .Z(n74191) );
  IV U91059 ( .A(n74191), .Z(n74186) );
  IV U91060 ( .A(n70732), .Z(n70733) );
  NOR U91061 ( .A(n70734), .B(n70733), .Z(n79647) );
  IV U91062 ( .A(n70735), .Z(n70736) );
  NOR U91063 ( .A(n70736), .B(n74183), .Z(n74177) );
  IV U91064 ( .A(n70737), .Z(n70739) );
  IV U91065 ( .A(n70738), .Z(n70741) );
  NOR U91066 ( .A(n70739), .B(n70741), .Z(n76187) );
  IV U91067 ( .A(n70740), .Z(n70742) );
  NOR U91068 ( .A(n70742), .B(n70741), .Z(n76184) );
  IV U91069 ( .A(n70743), .Z(n70747) );
  IV U91070 ( .A(n70744), .Z(n74140) );
  NOR U91071 ( .A(n74140), .B(n70745), .Z(n70746) );
  IV U91072 ( .A(n70746), .Z(n74159) );
  NOR U91073 ( .A(n70747), .B(n74159), .Z(n74153) );
  NOR U91074 ( .A(n70748), .B(n76196), .Z(n70751) );
  IV U91075 ( .A(n70749), .Z(n70750) );
  NOR U91076 ( .A(n70750), .B(n74144), .Z(n76192) );
  NOR U91077 ( .A(n70751), .B(n76192), .Z(n74137) );
  IV U91078 ( .A(n70752), .Z(n70756) );
  IV U91079 ( .A(n70753), .Z(n70761) );
  NOR U91080 ( .A(n70754), .B(n70761), .Z(n70755) );
  IV U91081 ( .A(n70755), .Z(n70758) );
  NOR U91082 ( .A(n70756), .B(n70758), .Z(n79620) );
  IV U91083 ( .A(n70757), .Z(n70759) );
  NOR U91084 ( .A(n70759), .B(n70758), .Z(n79623) );
  IV U91085 ( .A(n70760), .Z(n70762) );
  NOR U91086 ( .A(n70762), .B(n70761), .Z(n79614) );
  NOR U91087 ( .A(n79623), .B(n79614), .Z(n74136) );
  NOR U91088 ( .A(n70763), .B(n79605), .Z(n70771) );
  IV U91089 ( .A(n70764), .Z(n70769) );
  IV U91090 ( .A(n70765), .Z(n70766) );
  NOR U91091 ( .A(n70769), .B(n70766), .Z(n79601) );
  IV U91092 ( .A(n70767), .Z(n70768) );
  NOR U91093 ( .A(n70769), .B(n70768), .Z(n79600) );
  XOR U91094 ( .A(n79601), .B(n79600), .Z(n70770) );
  NOR U91095 ( .A(n70771), .B(n70770), .Z(n74135) );
  IV U91096 ( .A(n70772), .Z(n70773) );
  NOR U91097 ( .A(n70773), .B(n70775), .Z(n79592) );
  IV U91098 ( .A(n70774), .Z(n70778) );
  NOR U91099 ( .A(n70781), .B(n70775), .Z(n70776) );
  IV U91100 ( .A(n70776), .Z(n70777) );
  NOR U91101 ( .A(n70778), .B(n70777), .Z(n76203) );
  IV U91102 ( .A(n70779), .Z(n70784) );
  IV U91103 ( .A(n70780), .Z(n70785) );
  NOR U91104 ( .A(n70781), .B(n70785), .Z(n70782) );
  IV U91105 ( .A(n70782), .Z(n70783) );
  NOR U91106 ( .A(n70784), .B(n70783), .Z(n76200) );
  NOR U91107 ( .A(n70786), .B(n70785), .Z(n76208) );
  IV U91108 ( .A(n70787), .Z(n74132) );
  IV U91109 ( .A(n70788), .Z(n70789) );
  NOR U91110 ( .A(n74132), .B(n70789), .Z(n76218) );
  IV U91111 ( .A(n70790), .Z(n70791) );
  NOR U91112 ( .A(n70791), .B(n74128), .Z(n76215) );
  IV U91113 ( .A(n70792), .Z(n70798) );
  IV U91114 ( .A(n70793), .Z(n70795) );
  NOR U91115 ( .A(n70795), .B(n70794), .Z(n70796) );
  IV U91116 ( .A(n70796), .Z(n70797) );
  NOR U91117 ( .A(n70798), .B(n70797), .Z(n76220) );
  IV U91118 ( .A(n70799), .Z(n70800) );
  NOR U91119 ( .A(n70800), .B(n74119), .Z(n70801) );
  IV U91120 ( .A(n70801), .Z(n79583) );
  IV U91121 ( .A(n70802), .Z(n70803) );
  NOR U91122 ( .A(n70804), .B(n70803), .Z(n76230) );
  IV U91123 ( .A(n74120), .Z(n70805) );
  NOR U91124 ( .A(n70805), .B(n74119), .Z(n79578) );
  NOR U91125 ( .A(n76230), .B(n79578), .Z(n74117) );
  IV U91126 ( .A(n70806), .Z(n70807) );
  NOR U91127 ( .A(n70807), .B(n74113), .Z(n76232) );
  IV U91128 ( .A(n70808), .Z(n70814) );
  IV U91129 ( .A(n70809), .Z(n70811) );
  NOR U91130 ( .A(n70811), .B(n70810), .Z(n70812) );
  IV U91131 ( .A(n70812), .Z(n70813) );
  NOR U91132 ( .A(n70814), .B(n70813), .Z(n76240) );
  IV U91133 ( .A(n70815), .Z(n70818) );
  NOR U91134 ( .A(n70823), .B(n70816), .Z(n70817) );
  IV U91135 ( .A(n70817), .Z(n70819) );
  NOR U91136 ( .A(n70818), .B(n70819), .Z(n76237) );
  NOR U91137 ( .A(n70820), .B(n70819), .Z(n76248) );
  IV U91138 ( .A(n70821), .Z(n70822) );
  NOR U91139 ( .A(n70823), .B(n70822), .Z(n76245) );
  NOR U91140 ( .A(n70824), .B(n76262), .Z(n70828) );
  IV U91141 ( .A(n70825), .Z(n76254) );
  NOR U91142 ( .A(n70826), .B(n76254), .Z(n70827) );
  NOR U91143 ( .A(n70828), .B(n70827), .Z(n74107) );
  NOR U91144 ( .A(n70830), .B(n70829), .Z(n70831) );
  IV U91145 ( .A(n70831), .Z(n76277) );
  NOR U91146 ( .A(n70832), .B(n76277), .Z(n74100) );
  IV U91147 ( .A(n70833), .Z(n70834) );
  NOR U91148 ( .A(n70835), .B(n70834), .Z(n70836) );
  IV U91149 ( .A(n70836), .Z(n76276) );
  IV U91150 ( .A(n70837), .Z(n70839) );
  IV U91151 ( .A(n70838), .Z(n70843) );
  NOR U91152 ( .A(n70839), .B(n70843), .Z(n76282) );
  IV U91153 ( .A(n70840), .Z(n70841) );
  NOR U91154 ( .A(n70841), .B(n79549), .Z(n76285) );
  IV U91155 ( .A(n70842), .Z(n70844) );
  NOR U91156 ( .A(n70844), .B(n70843), .Z(n79556) );
  NOR U91157 ( .A(n76285), .B(n79556), .Z(n74098) );
  IV U91158 ( .A(n70845), .Z(n85333) );
  NOR U91159 ( .A(n70846), .B(n85333), .Z(n76288) );
  IV U91160 ( .A(n70847), .Z(n70850) );
  NOR U91161 ( .A(n70848), .B(n70860), .Z(n70849) );
  IV U91162 ( .A(n70849), .Z(n70854) );
  NOR U91163 ( .A(n70850), .B(n70854), .Z(n79543) );
  NOR U91164 ( .A(n76288), .B(n79543), .Z(n74097) );
  IV U91165 ( .A(n70851), .Z(n70852) );
  NOR U91166 ( .A(n79549), .B(n70852), .Z(n74095) );
  IV U91167 ( .A(n70853), .Z(n70855) );
  NOR U91168 ( .A(n70855), .B(n70854), .Z(n79536) );
  IV U91169 ( .A(n70856), .Z(n70857) );
  NOR U91170 ( .A(n70858), .B(n70857), .Z(n76290) );
  IV U91171 ( .A(n70859), .Z(n70861) );
  NOR U91172 ( .A(n70861), .B(n70860), .Z(n79533) );
  NOR U91173 ( .A(n76290), .B(n79533), .Z(n74094) );
  IV U91174 ( .A(n70862), .Z(n70863) );
  NOR U91175 ( .A(n70864), .B(n70863), .Z(n79527) );
  IV U91176 ( .A(n70865), .Z(n70867) );
  NOR U91177 ( .A(n70867), .B(n70866), .Z(n79530) );
  NOR U91178 ( .A(n79527), .B(n79530), .Z(n74093) );
  IV U91179 ( .A(n70868), .Z(n79520) );
  NOR U91180 ( .A(n70869), .B(n79520), .Z(n74092) );
  IV U91181 ( .A(n70870), .Z(n70872) );
  NOR U91182 ( .A(n70872), .B(n70871), .Z(n76293) );
  NOR U91183 ( .A(n70873), .B(n76296), .Z(n70874) );
  NOR U91184 ( .A(n76293), .B(n70874), .Z(n74091) );
  IV U91185 ( .A(n70875), .Z(n70877) );
  IV U91186 ( .A(n70876), .Z(n70882) );
  NOR U91187 ( .A(n70877), .B(n70882), .Z(n85295) );
  IV U91188 ( .A(n70878), .Z(n70879) );
  NOR U91189 ( .A(n70880), .B(n70879), .Z(n76299) );
  NOR U91190 ( .A(n85295), .B(n76299), .Z(n74090) );
  IV U91191 ( .A(n70881), .Z(n70883) );
  NOR U91192 ( .A(n70883), .B(n70882), .Z(n85281) );
  IV U91193 ( .A(n70884), .Z(n70886) );
  NOR U91194 ( .A(n70886), .B(n70885), .Z(n79501) );
  NOR U91195 ( .A(n70887), .B(n76304), .Z(n70888) );
  NOR U91196 ( .A(n79501), .B(n70888), .Z(n74089) );
  IV U91197 ( .A(n70889), .Z(n70891) );
  IV U91198 ( .A(n70890), .Z(n70895) );
  NOR U91199 ( .A(n70891), .B(n70895), .Z(n79490) );
  IV U91200 ( .A(n70892), .Z(n70893) );
  NOR U91201 ( .A(n70893), .B(n70898), .Z(n79486) );
  IV U91202 ( .A(n70894), .Z(n70896) );
  NOR U91203 ( .A(n70896), .B(n70895), .Z(n79481) );
  NOR U91204 ( .A(n79486), .B(n79481), .Z(n74081) );
  IV U91205 ( .A(n70897), .Z(n70899) );
  NOR U91206 ( .A(n70899), .B(n70898), .Z(n79483) );
  IV U91207 ( .A(n70900), .Z(n70901) );
  NOR U91208 ( .A(n70902), .B(n70901), .Z(n79477) );
  IV U91209 ( .A(n70903), .Z(n70905) );
  NOR U91210 ( .A(n70905), .B(n70904), .Z(n76308) );
  NOR U91211 ( .A(n79477), .B(n76308), .Z(n74080) );
  IV U91212 ( .A(n70906), .Z(n70908) );
  NOR U91213 ( .A(n70908), .B(n70907), .Z(n76313) );
  IV U91214 ( .A(n70909), .Z(n70910) );
  NOR U91215 ( .A(n70911), .B(n70910), .Z(n76310) );
  NOR U91216 ( .A(n76313), .B(n76310), .Z(n74079) );
  IV U91217 ( .A(n70912), .Z(n70914) );
  IV U91218 ( .A(n70913), .Z(n70916) );
  NOR U91219 ( .A(n70914), .B(n70916), .Z(n79461) );
  IV U91220 ( .A(n70915), .Z(n70917) );
  NOR U91221 ( .A(n70917), .B(n70916), .Z(n70918) );
  IV U91222 ( .A(n70918), .Z(n79454) );
  IV U91223 ( .A(n70919), .Z(n70920) );
  NOR U91224 ( .A(n70921), .B(n70920), .Z(n79448) );
  IV U91225 ( .A(n70922), .Z(n70923) );
  NOR U91226 ( .A(n70923), .B(n70928), .Z(n79440) );
  IV U91227 ( .A(n70924), .Z(n70932) );
  IV U91228 ( .A(n70925), .Z(n70926) );
  NOR U91229 ( .A(n70932), .B(n70926), .Z(n79437) );
  IV U91230 ( .A(n70927), .Z(n70929) );
  NOR U91231 ( .A(n70929), .B(n70928), .Z(n79443) );
  NOR U91232 ( .A(n79437), .B(n79443), .Z(n74071) );
  IV U91233 ( .A(n70930), .Z(n70931) );
  NOR U91234 ( .A(n70932), .B(n70931), .Z(n76317) );
  IV U91235 ( .A(n70933), .Z(n70935) );
  NOR U91236 ( .A(n70935), .B(n70934), .Z(n79412) );
  NOR U91237 ( .A(n70936), .B(n76324), .Z(n70937) );
  NOR U91238 ( .A(n79412), .B(n70937), .Z(n70938) );
  IV U91239 ( .A(n70938), .Z(n74056) );
  IV U91240 ( .A(n70939), .Z(n70941) );
  NOR U91241 ( .A(n70941), .B(n70940), .Z(n79400) );
  IV U91242 ( .A(n70942), .Z(n70943) );
  NOR U91243 ( .A(n70944), .B(n70943), .Z(n79405) );
  NOR U91244 ( .A(n79400), .B(n79405), .Z(n74055) );
  IV U91245 ( .A(n70945), .Z(n70947) );
  NOR U91246 ( .A(n70947), .B(n70946), .Z(n76330) );
  IV U91247 ( .A(n70948), .Z(n70950) );
  NOR U91248 ( .A(n70950), .B(n70949), .Z(n79394) );
  IV U91249 ( .A(n70951), .Z(n70953) );
  NOR U91250 ( .A(n70953), .B(n70952), .Z(n76335) );
  NOR U91251 ( .A(n79394), .B(n76335), .Z(n74046) );
  IV U91252 ( .A(n70954), .Z(n70956) );
  NOR U91253 ( .A(n70956), .B(n70955), .Z(n81892) );
  IV U91254 ( .A(n70957), .Z(n70959) );
  NOR U91255 ( .A(n70959), .B(n70958), .Z(n81887) );
  NOR U91256 ( .A(n81892), .B(n81887), .Z(n79392) );
  IV U91257 ( .A(n70960), .Z(n70964) );
  IV U91258 ( .A(n70961), .Z(n70969) );
  NOR U91259 ( .A(n70969), .B(n70962), .Z(n70963) );
  IV U91260 ( .A(n70963), .Z(n70966) );
  NOR U91261 ( .A(n70964), .B(n70966), .Z(n76341) );
  NOR U91262 ( .A(n79386), .B(n76341), .Z(n74045) );
  IV U91263 ( .A(n70965), .Z(n70967) );
  NOR U91264 ( .A(n70967), .B(n70966), .Z(n76338) );
  NOR U91265 ( .A(n70969), .B(n70968), .Z(n81903) );
  IV U91266 ( .A(n70970), .Z(n70971) );
  NOR U91267 ( .A(n70974), .B(n70971), .Z(n81908) );
  NOR U91268 ( .A(n81903), .B(n81908), .Z(n76345) );
  IV U91269 ( .A(n70972), .Z(n70973) );
  NOR U91270 ( .A(n70974), .B(n70973), .Z(n76349) );
  IV U91271 ( .A(n70975), .Z(n70976) );
  NOR U91272 ( .A(n70977), .B(n70976), .Z(n76346) );
  NOR U91273 ( .A(n76349), .B(n76346), .Z(n74044) );
  IV U91274 ( .A(n70978), .Z(n70979) );
  NOR U91275 ( .A(n70979), .B(n70982), .Z(n79376) );
  IV U91276 ( .A(n70980), .Z(n70981) );
  NOR U91277 ( .A(n70982), .B(n70981), .Z(n79373) );
  IV U91278 ( .A(n70983), .Z(n70985) );
  NOR U91279 ( .A(n70985), .B(n70984), .Z(n70986) );
  IV U91280 ( .A(n70986), .Z(n74040) );
  IV U91281 ( .A(n70987), .Z(n70988) );
  NOR U91282 ( .A(n70989), .B(n70988), .Z(n85219) );
  IV U91283 ( .A(n70990), .Z(n70991) );
  NOR U91284 ( .A(n70991), .B(n74034), .Z(n81922) );
  NOR U91285 ( .A(n85219), .B(n81922), .Z(n76352) );
  IV U91286 ( .A(n70992), .Z(n70994) );
  NOR U91287 ( .A(n70994), .B(n70993), .Z(n76353) );
  IV U91288 ( .A(n70995), .Z(n70996) );
  NOR U91289 ( .A(n70996), .B(n71002), .Z(n79367) );
  NOR U91290 ( .A(n76353), .B(n79367), .Z(n70997) );
  IV U91291 ( .A(n70997), .Z(n74031) );
  IV U91292 ( .A(n70998), .Z(n71000) );
  NOR U91293 ( .A(n71000), .B(n70999), .Z(n76358) );
  IV U91294 ( .A(n71001), .Z(n71003) );
  NOR U91295 ( .A(n71003), .B(n71002), .Z(n79364) );
  NOR U91296 ( .A(n76358), .B(n79364), .Z(n74030) );
  IV U91297 ( .A(n71004), .Z(n71006) );
  NOR U91298 ( .A(n71006), .B(n71005), .Z(n71007) );
  IV U91299 ( .A(n71007), .Z(n74025) );
  IV U91300 ( .A(n71008), .Z(n71009) );
  NOR U91301 ( .A(n90895), .B(n71009), .Z(n71010) );
  IV U91302 ( .A(n71010), .Z(n73998) );
  IV U91303 ( .A(n71011), .Z(n71012) );
  NOR U91304 ( .A(n71012), .B(n73997), .Z(n76379) );
  IV U91305 ( .A(n71013), .Z(n71014) );
  NOR U91306 ( .A(n71014), .B(n73989), .Z(n73983) );
  IV U91307 ( .A(n73983), .Z(n73975) );
  IV U91308 ( .A(n71015), .Z(n71020) );
  IV U91309 ( .A(n71016), .Z(n71017) );
  NOR U91310 ( .A(n71020), .B(n71017), .Z(n71018) );
  IV U91311 ( .A(n71018), .Z(n79349) );
  IV U91312 ( .A(n71019), .Z(n71021) );
  NOR U91313 ( .A(n71021), .B(n71020), .Z(n79342) );
  IV U91314 ( .A(n71022), .Z(n71024) );
  NOR U91315 ( .A(n71024), .B(n71023), .Z(n76388) );
  IV U91316 ( .A(n71025), .Z(n71027) );
  NOR U91317 ( .A(n71027), .B(n71026), .Z(n76384) );
  NOR U91318 ( .A(n76388), .B(n76384), .Z(n73967) );
  IV U91319 ( .A(n71028), .Z(n71029) );
  NOR U91320 ( .A(n71030), .B(n71029), .Z(n81974) );
  IV U91321 ( .A(n71031), .Z(n71033) );
  NOR U91322 ( .A(n71033), .B(n71032), .Z(n81969) );
  NOR U91323 ( .A(n81974), .B(n81969), .Z(n79334) );
  IV U91324 ( .A(n71034), .Z(n71035) );
  NOR U91325 ( .A(n71036), .B(n71035), .Z(n79326) );
  IV U91326 ( .A(n71037), .Z(n71038) );
  NOR U91327 ( .A(n71039), .B(n71038), .Z(n73952) );
  IV U91328 ( .A(n73952), .Z(n73942) );
  IV U91329 ( .A(n71040), .Z(n71041) );
  NOR U91330 ( .A(n71042), .B(n71041), .Z(n76395) );
  IV U91331 ( .A(n71043), .Z(n71044) );
  NOR U91332 ( .A(n71045), .B(n71044), .Z(n76393) );
  NOR U91333 ( .A(n76395), .B(n76393), .Z(n73940) );
  IV U91334 ( .A(n71046), .Z(n71047) );
  NOR U91335 ( .A(n71048), .B(n71047), .Z(n71049) );
  IV U91336 ( .A(n71049), .Z(n79311) );
  IV U91337 ( .A(n71050), .Z(n71051) );
  NOR U91338 ( .A(n71052), .B(n71051), .Z(n76404) );
  NOR U91339 ( .A(n71053), .B(n76401), .Z(n71054) );
  NOR U91340 ( .A(n76404), .B(n71054), .Z(n73931) );
  IV U91341 ( .A(n71055), .Z(n71057) );
  NOR U91342 ( .A(n71057), .B(n71056), .Z(n76411) );
  IV U91343 ( .A(n71058), .Z(n71059) );
  NOR U91344 ( .A(n71060), .B(n71059), .Z(n76407) );
  NOR U91345 ( .A(n76411), .B(n76407), .Z(n73930) );
  IV U91346 ( .A(n71061), .Z(n71062) );
  NOR U91347 ( .A(n71063), .B(n71062), .Z(n73928) );
  IV U91348 ( .A(n73928), .Z(n73920) );
  NOR U91349 ( .A(n79297), .B(n79303), .Z(n71064) );
  NOR U91350 ( .A(n79298), .B(n71064), .Z(n73919) );
  IV U91351 ( .A(n71065), .Z(n71066) );
  NOR U91352 ( .A(n71067), .B(n71066), .Z(n76423) );
  IV U91353 ( .A(n71068), .Z(n71070) );
  NOR U91354 ( .A(n71070), .B(n71069), .Z(n76418) );
  NOR U91355 ( .A(n76423), .B(n76418), .Z(n73911) );
  IV U91356 ( .A(n71071), .Z(n71072) );
  NOR U91357 ( .A(n71073), .B(n71072), .Z(n71074) );
  IV U91358 ( .A(n71074), .Z(n71075) );
  NOR U91359 ( .A(n71076), .B(n71075), .Z(n76420) );
  IV U91360 ( .A(n71077), .Z(n71078) );
  NOR U91361 ( .A(n71078), .B(n82042), .Z(n76442) );
  IV U91362 ( .A(n71079), .Z(n71080) );
  NOR U91363 ( .A(n82042), .B(n71080), .Z(n76439) );
  IV U91364 ( .A(n71081), .Z(n71082) );
  NOR U91365 ( .A(n71083), .B(n71082), .Z(n76458) );
  IV U91366 ( .A(n71084), .Z(n71086) );
  IV U91367 ( .A(n71085), .Z(n71088) );
  NOR U91368 ( .A(n71086), .B(n71088), .Z(n76460) );
  NOR U91369 ( .A(n76458), .B(n76460), .Z(n73885) );
  IV U91370 ( .A(n71087), .Z(n71089) );
  NOR U91371 ( .A(n71089), .B(n71088), .Z(n79265) );
  IV U91372 ( .A(n71090), .Z(n71092) );
  NOR U91373 ( .A(n71092), .B(n71091), .Z(n76482) );
  IV U91374 ( .A(n71093), .Z(n71094) );
  NOR U91375 ( .A(n71094), .B(n73846), .Z(n76477) );
  NOR U91376 ( .A(n76482), .B(n76477), .Z(n73843) );
  IV U91377 ( .A(n71095), .Z(n71097) );
  NOR U91378 ( .A(n71097), .B(n71096), .Z(n76479) );
  IV U91379 ( .A(n71098), .Z(n71100) );
  NOR U91380 ( .A(n71100), .B(n71099), .Z(n76485) );
  NOR U91381 ( .A(n71102), .B(n71101), .Z(n71103) );
  IV U91382 ( .A(n71103), .Z(n71104) );
  NOR U91383 ( .A(n71105), .B(n71104), .Z(n76487) );
  NOR U91384 ( .A(n76485), .B(n76487), .Z(n73839) );
  IV U91385 ( .A(n71106), .Z(n73813) );
  IV U91386 ( .A(n71107), .Z(n71108) );
  NOR U91387 ( .A(n73813), .B(n71108), .Z(n79225) );
  IV U91388 ( .A(n71109), .Z(n71110) );
  NOR U91389 ( .A(n71110), .B(n71115), .Z(n79222) );
  IV U91390 ( .A(n71111), .Z(n71113) );
  NOR U91391 ( .A(n71113), .B(n71112), .Z(n79216) );
  IV U91392 ( .A(n71114), .Z(n71116) );
  NOR U91393 ( .A(n71116), .B(n71115), .Z(n79219) );
  NOR U91394 ( .A(n79216), .B(n79219), .Z(n73809) );
  IV U91395 ( .A(n71117), .Z(n71118) );
  NOR U91396 ( .A(n71119), .B(n71118), .Z(n76503) );
  IV U91397 ( .A(n71120), .Z(n73801) );
  IV U91398 ( .A(n71121), .Z(n71122) );
  NOR U91399 ( .A(n73801), .B(n71122), .Z(n76511) );
  IV U91400 ( .A(n71123), .Z(n71124) );
  NOR U91401 ( .A(n71124), .B(n73795), .Z(n76515) );
  NOR U91402 ( .A(n76511), .B(n76515), .Z(n73798) );
  IV U91403 ( .A(n71125), .Z(n71126) );
  NOR U91404 ( .A(n73792), .B(n71126), .Z(n79207) );
  IV U91405 ( .A(n71127), .Z(n71128) );
  NOR U91406 ( .A(n71128), .B(n73779), .Z(n76526) );
  IV U91407 ( .A(n71129), .Z(n71130) );
  NOR U91408 ( .A(n71131), .B(n71130), .Z(n73774) );
  IV U91409 ( .A(n73774), .Z(n73768) );
  IV U91410 ( .A(n71132), .Z(n71133) );
  NOR U91411 ( .A(n71134), .B(n71133), .Z(n82157) );
  IV U91412 ( .A(n71135), .Z(n71136) );
  NOR U91413 ( .A(n71139), .B(n71136), .Z(n85005) );
  NOR U91414 ( .A(n82157), .B(n85005), .Z(n76533) );
  IV U91415 ( .A(n71137), .Z(n71138) );
  NOR U91416 ( .A(n71139), .B(n71138), .Z(n79174) );
  NOR U91417 ( .A(n71141), .B(n71140), .Z(n79157) );
  IV U91418 ( .A(n71142), .Z(n71144) );
  NOR U91419 ( .A(n71144), .B(n71143), .Z(n76549) );
  IV U91420 ( .A(n71145), .Z(n71147) );
  NOR U91421 ( .A(n71147), .B(n71146), .Z(n76546) );
  NOR U91422 ( .A(n76549), .B(n76546), .Z(n73736) );
  IV U91423 ( .A(n71148), .Z(n76556) );
  NOR U91424 ( .A(n71149), .B(n76556), .Z(n71153) );
  IV U91425 ( .A(n71150), .Z(n71151) );
  NOR U91426 ( .A(n71152), .B(n71151), .Z(n76552) );
  NOR U91427 ( .A(n71153), .B(n76552), .Z(n73735) );
  NOR U91428 ( .A(n71154), .B(n79140), .Z(n73734) );
  IV U91429 ( .A(n71155), .Z(n71157) );
  NOR U91430 ( .A(n71157), .B(n71156), .Z(n79137) );
  IV U91431 ( .A(n71158), .Z(n71159) );
  NOR U91432 ( .A(n71160), .B(n71159), .Z(n79144) );
  NOR U91433 ( .A(n79137), .B(n79144), .Z(n71161) );
  IV U91434 ( .A(n71161), .Z(n73733) );
  IV U91435 ( .A(n71162), .Z(n71163) );
  NOR U91436 ( .A(n71164), .B(n71163), .Z(n84917) );
  IV U91437 ( .A(n71165), .Z(n71166) );
  NOR U91438 ( .A(n71167), .B(n71166), .Z(n82189) );
  NOR U91439 ( .A(n84917), .B(n82189), .Z(n79132) );
  IV U91440 ( .A(n71168), .Z(n71175) );
  IV U91441 ( .A(n71169), .Z(n73710) );
  NOR U91442 ( .A(n71170), .B(n73710), .Z(n71171) );
  IV U91443 ( .A(n71171), .Z(n71172) );
  NOR U91444 ( .A(n71173), .B(n71172), .Z(n71174) );
  IV U91445 ( .A(n71174), .Z(n71183) );
  NOR U91446 ( .A(n71175), .B(n71183), .Z(n76566) );
  IV U91447 ( .A(n71176), .Z(n71177) );
  NOR U91448 ( .A(n71177), .B(n71179), .Z(n79120) );
  IV U91449 ( .A(n71178), .Z(n71180) );
  NOR U91450 ( .A(n71180), .B(n71179), .Z(n79116) );
  NOR U91451 ( .A(n79120), .B(n79116), .Z(n71181) );
  IV U91452 ( .A(n71181), .Z(n71185) );
  IV U91453 ( .A(n71182), .Z(n71184) );
  NOR U91454 ( .A(n71184), .B(n71183), .Z(n76572) );
  NOR U91455 ( .A(n71185), .B(n76572), .Z(n71186) );
  IV U91456 ( .A(n71186), .Z(n73708) );
  IV U91457 ( .A(n71187), .Z(n71189) );
  NOR U91458 ( .A(n71189), .B(n71188), .Z(n71190) );
  IV U91459 ( .A(n71190), .Z(n79115) );
  IV U91460 ( .A(n71191), .Z(n71192) );
  NOR U91461 ( .A(n71193), .B(n71192), .Z(n71194) );
  IV U91462 ( .A(n71194), .Z(n73703) );
  IV U91463 ( .A(n71195), .Z(n71197) );
  NOR U91464 ( .A(n71197), .B(n71196), .Z(n73688) );
  IV U91465 ( .A(n71198), .Z(n71200) );
  NOR U91466 ( .A(n71200), .B(n71199), .Z(n79104) );
  IV U91467 ( .A(n71201), .Z(n71202) );
  NOR U91468 ( .A(n71202), .B(n71204), .Z(n79101) );
  IV U91469 ( .A(n71203), .Z(n71205) );
  NOR U91470 ( .A(n71205), .B(n71204), .Z(n79096) );
  IV U91471 ( .A(n71206), .Z(n71208) );
  NOR U91472 ( .A(n71208), .B(n71207), .Z(n79093) );
  IV U91473 ( .A(n71209), .Z(n71214) );
  IV U91474 ( .A(n71210), .Z(n71211) );
  NOR U91475 ( .A(n71214), .B(n71211), .Z(n79090) );
  NOR U91476 ( .A(n79093), .B(n79090), .Z(n73682) );
  IV U91477 ( .A(n71212), .Z(n71216) );
  NOR U91478 ( .A(n71214), .B(n71213), .Z(n71215) );
  IV U91479 ( .A(n71215), .Z(n71218) );
  NOR U91480 ( .A(n71216), .B(n71218), .Z(n79087) );
  IV U91481 ( .A(n71217), .Z(n71219) );
  NOR U91482 ( .A(n71219), .B(n71218), .Z(n76578) );
  IV U91483 ( .A(n71220), .Z(n71221) );
  NOR U91484 ( .A(n71221), .B(n73680), .Z(n79079) );
  IV U91485 ( .A(n71222), .Z(n73673) );
  IV U91486 ( .A(n71223), .Z(n71224) );
  NOR U91487 ( .A(n73673), .B(n71224), .Z(n79069) );
  IV U91488 ( .A(n71225), .Z(n71226) );
  NOR U91489 ( .A(n71232), .B(n71226), .Z(n79066) );
  IV U91490 ( .A(n71227), .Z(n71229) );
  NOR U91491 ( .A(n71229), .B(n71228), .Z(n79063) );
  IV U91492 ( .A(n71230), .Z(n71231) );
  NOR U91493 ( .A(n71232), .B(n71231), .Z(n76584) );
  NOR U91494 ( .A(n79063), .B(n76584), .Z(n71233) );
  IV U91495 ( .A(n71233), .Z(n73670) );
  IV U91496 ( .A(n71234), .Z(n71235) );
  NOR U91497 ( .A(n73666), .B(n71235), .Z(n79062) );
  IV U91498 ( .A(n71236), .Z(n71238) );
  NOR U91499 ( .A(n71238), .B(n71237), .Z(n76589) );
  IV U91500 ( .A(n71239), .Z(n71244) );
  IV U91501 ( .A(n71240), .Z(n71241) );
  NOR U91502 ( .A(n71244), .B(n71241), .Z(n76593) );
  IV U91503 ( .A(n71242), .Z(n71243) );
  NOR U91504 ( .A(n71244), .B(n71243), .Z(n76602) );
  IV U91505 ( .A(n71245), .Z(n71246) );
  NOR U91506 ( .A(n71246), .B(n73661), .Z(n76599) );
  IV U91507 ( .A(n71247), .Z(n71253) );
  NOR U91508 ( .A(n71248), .B(n73641), .Z(n71249) );
  IV U91509 ( .A(n71249), .Z(n71250) );
  NOR U91510 ( .A(n71251), .B(n71250), .Z(n71252) );
  IV U91511 ( .A(n71252), .Z(n73647) );
  NOR U91512 ( .A(n71253), .B(n73647), .Z(n79045) );
  IV U91513 ( .A(n71254), .Z(n71255) );
  NOR U91514 ( .A(n71255), .B(n71259), .Z(n79033) );
  IV U91515 ( .A(n71256), .Z(n71257) );
  NOR U91516 ( .A(n71257), .B(n71262), .Z(n79026) );
  IV U91517 ( .A(n71258), .Z(n71260) );
  NOR U91518 ( .A(n71260), .B(n71259), .Z(n79029) );
  NOR U91519 ( .A(n79026), .B(n79029), .Z(n73638) );
  IV U91520 ( .A(n71261), .Z(n71263) );
  NOR U91521 ( .A(n71263), .B(n71262), .Z(n73635) );
  IV U91522 ( .A(n71264), .Z(n71265) );
  NOR U91523 ( .A(n71266), .B(n71265), .Z(n76667) );
  IV U91524 ( .A(n71267), .Z(n71269) );
  NOR U91525 ( .A(n71269), .B(n71268), .Z(n76658) );
  NOR U91526 ( .A(n76667), .B(n76658), .Z(n73601) );
  IV U91527 ( .A(n71270), .Z(n73596) );
  IV U91528 ( .A(n71271), .Z(n71272) );
  NOR U91529 ( .A(n73596), .B(n71272), .Z(n76664) );
  IV U91530 ( .A(n71273), .Z(n71274) );
  NOR U91531 ( .A(n71275), .B(n71274), .Z(n76671) );
  IV U91532 ( .A(n71276), .Z(n71277) );
  NOR U91533 ( .A(n71277), .B(n73598), .Z(n79013) );
  NOR U91534 ( .A(n76671), .B(n79013), .Z(n73593) );
  IV U91535 ( .A(n73587), .Z(n71279) );
  IV U91536 ( .A(n71278), .Z(n71281) );
  NOR U91537 ( .A(n71279), .B(n71281), .Z(n73584) );
  IV U91538 ( .A(n71280), .Z(n71282) );
  NOR U91539 ( .A(n71282), .B(n71281), .Z(n73588) );
  NOR U91540 ( .A(n73584), .B(n73588), .Z(n71283) );
  IV U91541 ( .A(n71283), .Z(n73583) );
  IV U91542 ( .A(n71284), .Z(n76675) );
  IV U91543 ( .A(n71285), .Z(n71286) );
  NOR U91544 ( .A(n71286), .B(n71288), .Z(n76679) );
  IV U91545 ( .A(n71287), .Z(n71289) );
  NOR U91546 ( .A(n71289), .B(n71288), .Z(n76676) );
  NOR U91547 ( .A(n76679), .B(n76676), .Z(n73582) );
  IV U91548 ( .A(n71290), .Z(n71292) );
  NOR U91549 ( .A(n71292), .B(n71291), .Z(n71293) );
  NOR U91550 ( .A(n82317), .B(n71293), .Z(n76691) );
  IV U91551 ( .A(n71294), .Z(n71295) );
  NOR U91552 ( .A(n73568), .B(n71295), .Z(n73565) );
  IV U91553 ( .A(n73565), .Z(n73559) );
  IV U91554 ( .A(n71296), .Z(n71301) );
  IV U91555 ( .A(n71297), .Z(n71298) );
  NOR U91556 ( .A(n71301), .B(n71298), .Z(n78988) );
  NOR U91557 ( .A(n71299), .B(n76696), .Z(n71303) );
  IV U91558 ( .A(n71300), .Z(n71302) );
  NOR U91559 ( .A(n71302), .B(n71301), .Z(n76693) );
  NOR U91560 ( .A(n71303), .B(n76693), .Z(n73557) );
  IV U91561 ( .A(n71304), .Z(n71305) );
  NOR U91562 ( .A(n71306), .B(n71305), .Z(n76700) );
  IV U91563 ( .A(n71307), .Z(n71308) );
  NOR U91564 ( .A(n71309), .B(n71308), .Z(n78979) );
  NOR U91565 ( .A(n76700), .B(n78979), .Z(n73556) );
  IV U91566 ( .A(n71310), .Z(n71312) );
  NOR U91567 ( .A(n71312), .B(n71311), .Z(n76702) );
  IV U91568 ( .A(n71313), .Z(n71314) );
  NOR U91569 ( .A(n71315), .B(n71314), .Z(n71316) );
  IV U91570 ( .A(n71316), .Z(n76719) );
  IV U91571 ( .A(n71317), .Z(n71319) );
  NOR U91572 ( .A(n71319), .B(n71318), .Z(n76725) );
  IV U91573 ( .A(n71320), .Z(n71321) );
  NOR U91574 ( .A(n71322), .B(n71321), .Z(n76720) );
  NOR U91575 ( .A(n76725), .B(n76720), .Z(n73528) );
  IV U91576 ( .A(n71323), .Z(n71324) );
  NOR U91577 ( .A(n71325), .B(n71324), .Z(n71326) );
  IV U91578 ( .A(n71326), .Z(n76723) );
  IV U91579 ( .A(n71327), .Z(n71328) );
  NOR U91580 ( .A(n71328), .B(n71330), .Z(n76730) );
  IV U91581 ( .A(n71329), .Z(n71331) );
  NOR U91582 ( .A(n71331), .B(n71330), .Z(n76728) );
  NOR U91583 ( .A(n76730), .B(n76728), .Z(n73527) );
  IV U91584 ( .A(n71332), .Z(n71333) );
  NOR U91585 ( .A(n71334), .B(n71333), .Z(n78957) );
  IV U91586 ( .A(n71335), .Z(n71337) );
  NOR U91587 ( .A(n71337), .B(n71336), .Z(n78962) );
  NOR U91588 ( .A(n78957), .B(n78962), .Z(n73526) );
  IV U91589 ( .A(n71338), .Z(n71339) );
  NOR U91590 ( .A(n73505), .B(n71339), .Z(n76735) );
  IV U91591 ( .A(n71340), .Z(n71342) );
  IV U91592 ( .A(n71341), .Z(n73501) );
  NOR U91593 ( .A(n71342), .B(n73501), .Z(n78948) );
  IV U91594 ( .A(n71343), .Z(n71344) );
  NOR U91595 ( .A(n73499), .B(n71344), .Z(n84654) );
  IV U91596 ( .A(n71345), .Z(n71347) );
  IV U91597 ( .A(n71346), .Z(n71351) );
  NOR U91598 ( .A(n71347), .B(n71351), .Z(n84660) );
  NOR U91599 ( .A(n84654), .B(n84660), .Z(n76745) );
  IV U91600 ( .A(n76745), .Z(n73496) );
  IV U91601 ( .A(n71348), .Z(n71357) );
  NOR U91602 ( .A(n71350), .B(n71349), .Z(n71352) );
  NOR U91603 ( .A(n71352), .B(n71351), .Z(n71353) );
  IV U91604 ( .A(n71353), .Z(n71354) );
  NOR U91605 ( .A(n71355), .B(n71354), .Z(n71356) );
  IV U91606 ( .A(n71356), .Z(n71359) );
  NOR U91607 ( .A(n71357), .B(n71359), .Z(n76749) );
  IV U91608 ( .A(n71358), .Z(n71360) );
  NOR U91609 ( .A(n71360), .B(n71359), .Z(n78941) );
  IV U91610 ( .A(n71361), .Z(n71363) );
  NOR U91611 ( .A(n71363), .B(n71362), .Z(n78928) );
  IV U91612 ( .A(n71364), .Z(n71366) );
  NOR U91613 ( .A(n71366), .B(n71365), .Z(n78931) );
  IV U91614 ( .A(n71367), .Z(n71368) );
  XOR U91615 ( .A(n71376), .B(n71377), .Z(n71370) );
  NOR U91616 ( .A(n71368), .B(n71370), .Z(n76758) );
  NOR U91617 ( .A(n78931), .B(n76758), .Z(n73487) );
  IV U91618 ( .A(n71369), .Z(n71371) );
  NOR U91619 ( .A(n71371), .B(n71370), .Z(n76760) );
  IV U91620 ( .A(n71372), .Z(n71375) );
  NOR U91621 ( .A(n71373), .B(n71377), .Z(n71374) );
  IV U91622 ( .A(n71374), .Z(n71380) );
  NOR U91623 ( .A(n71375), .B(n71380), .Z(n76762) );
  NOR U91624 ( .A(n76760), .B(n76762), .Z(n73486) );
  IV U91625 ( .A(n71376), .Z(n71378) );
  NOR U91626 ( .A(n71378), .B(n71377), .Z(n78911) );
  IV U91627 ( .A(n71379), .Z(n71381) );
  NOR U91628 ( .A(n71381), .B(n71380), .Z(n78923) );
  NOR U91629 ( .A(n78911), .B(n78923), .Z(n73485) );
  IV U91630 ( .A(n71382), .Z(n71383) );
  NOR U91631 ( .A(n71384), .B(n71383), .Z(n71385) );
  IV U91632 ( .A(n71385), .Z(n73480) );
  IV U91633 ( .A(n71386), .Z(n71389) );
  NOR U91634 ( .A(n71395), .B(n71387), .Z(n71388) );
  IV U91635 ( .A(n71388), .Z(n71391) );
  NOR U91636 ( .A(n71389), .B(n71391), .Z(n78904) );
  IV U91637 ( .A(n71390), .Z(n71392) );
  NOR U91638 ( .A(n71392), .B(n71391), .Z(n78899) );
  IV U91639 ( .A(n71393), .Z(n71394) );
  NOR U91640 ( .A(n71395), .B(n71394), .Z(n82421) );
  IV U91641 ( .A(n71396), .Z(n71397) );
  NOR U91642 ( .A(n71397), .B(n71402), .Z(n82426) );
  NOR U91643 ( .A(n82421), .B(n82426), .Z(n78898) );
  IV U91644 ( .A(n71398), .Z(n71400) );
  NOR U91645 ( .A(n71400), .B(n71399), .Z(n76767) );
  IV U91646 ( .A(n71401), .Z(n71403) );
  NOR U91647 ( .A(n71403), .B(n71402), .Z(n76765) );
  NOR U91648 ( .A(n76767), .B(n76765), .Z(n73476) );
  IV U91649 ( .A(n71404), .Z(n71405) );
  NOR U91650 ( .A(n71406), .B(n71405), .Z(n82437) );
  IV U91651 ( .A(n71407), .Z(n71408) );
  NOR U91652 ( .A(n71409), .B(n71408), .Z(n82431) );
  NOR U91653 ( .A(n82437), .B(n82431), .Z(n78888) );
  IV U91654 ( .A(n71410), .Z(n71411) );
  NOR U91655 ( .A(n73459), .B(n71411), .Z(n76788) );
  IV U91656 ( .A(n71412), .Z(n71418) );
  NOR U91657 ( .A(n71414), .B(n71413), .Z(n71415) );
  IV U91658 ( .A(n71415), .Z(n73461) );
  NOR U91659 ( .A(n71416), .B(n73461), .Z(n71417) );
  IV U91660 ( .A(n71417), .Z(n73455) );
  NOR U91661 ( .A(n71418), .B(n73455), .Z(n76792) );
  IV U91662 ( .A(n71419), .Z(n71421) );
  IV U91663 ( .A(n71420), .Z(n71423) );
  NOR U91664 ( .A(n71421), .B(n71423), .Z(n78857) );
  IV U91665 ( .A(n71422), .Z(n71424) );
  NOR U91666 ( .A(n71424), .B(n71423), .Z(n78852) );
  NOR U91667 ( .A(n78849), .B(n78852), .Z(n71425) );
  IV U91668 ( .A(n71425), .Z(n73453) );
  IV U91669 ( .A(n71426), .Z(n78848) );
  IV U91670 ( .A(n71427), .Z(n71428) );
  NOR U91671 ( .A(n71429), .B(n71428), .Z(n71434) );
  IV U91672 ( .A(n71430), .Z(n71432) );
  NOR U91673 ( .A(n71432), .B(n71431), .Z(n71433) );
  NOR U91674 ( .A(n71434), .B(n71433), .Z(n78840) );
  IV U91675 ( .A(n71435), .Z(n71436) );
  NOR U91676 ( .A(n71437), .B(n71436), .Z(n78835) );
  IV U91677 ( .A(n71438), .Z(n71439) );
  NOR U91678 ( .A(n71440), .B(n71439), .Z(n78842) );
  NOR U91679 ( .A(n78835), .B(n78842), .Z(n73452) );
  IV U91680 ( .A(n71441), .Z(n71443) );
  NOR U91681 ( .A(n71443), .B(n71442), .Z(n82463) );
  IV U91682 ( .A(n71444), .Z(n71446) );
  NOR U91683 ( .A(n71446), .B(n71445), .Z(n82458) );
  NOR U91684 ( .A(n82463), .B(n82458), .Z(n78834) );
  IV U91685 ( .A(n71447), .Z(n71448) );
  NOR U91686 ( .A(n71449), .B(n71448), .Z(n71450) );
  IV U91687 ( .A(n71450), .Z(n76808) );
  IV U91688 ( .A(n71451), .Z(n71453) );
  NOR U91689 ( .A(n71453), .B(n71452), .Z(n78828) );
  IV U91690 ( .A(n71454), .Z(n71455) );
  NOR U91691 ( .A(n71456), .B(n71455), .Z(n76812) );
  NOR U91692 ( .A(n78828), .B(n76812), .Z(n73437) );
  IV U91693 ( .A(n71457), .Z(n73435) );
  IV U91694 ( .A(n71458), .Z(n71459) );
  NOR U91695 ( .A(n73435), .B(n71459), .Z(n78819) );
  IV U91696 ( .A(n71460), .Z(n71463) );
  NOR U91697 ( .A(n71461), .B(n73427), .Z(n71462) );
  IV U91698 ( .A(n71462), .Z(n71465) );
  NOR U91699 ( .A(n71463), .B(n71465), .Z(n76821) );
  NOR U91700 ( .A(n78819), .B(n76821), .Z(n90424) );
  IV U91701 ( .A(n71464), .Z(n71466) );
  NOR U91702 ( .A(n71466), .B(n71465), .Z(n76820) );
  IV U91703 ( .A(n71467), .Z(n71468) );
  NOR U91704 ( .A(n71469), .B(n71468), .Z(n76847) );
  IV U91705 ( .A(n71470), .Z(n71472) );
  IV U91706 ( .A(n71471), .Z(n71476) );
  NOR U91707 ( .A(n71472), .B(n71476), .Z(n76850) );
  NOR U91708 ( .A(n71474), .B(n71473), .Z(n76858) );
  IV U91709 ( .A(n71475), .Z(n71477) );
  NOR U91710 ( .A(n71477), .B(n71476), .Z(n76855) );
  NOR U91711 ( .A(n76858), .B(n76855), .Z(n73379) );
  IV U91712 ( .A(n71478), .Z(n78785) );
  NOR U91713 ( .A(n78785), .B(n71479), .Z(n76861) );
  IV U91714 ( .A(n71480), .Z(n71481) );
  NOR U91715 ( .A(n71481), .B(n73376), .Z(n78778) );
  IV U91716 ( .A(n71482), .Z(n71483) );
  NOR U91717 ( .A(n71483), .B(n73376), .Z(n71484) );
  IV U91718 ( .A(n71484), .Z(n78776) );
  IV U91719 ( .A(n71485), .Z(n71486) );
  NOR U91720 ( .A(n71486), .B(n73371), .Z(n76876) );
  IV U91721 ( .A(n71487), .Z(n71489) );
  NOR U91722 ( .A(n71489), .B(n71488), .Z(n78766) );
  IV U91723 ( .A(n71490), .Z(n71492) );
  NOR U91724 ( .A(n71492), .B(n71491), .Z(n76871) );
  NOR U91725 ( .A(n78766), .B(n76871), .Z(n71493) );
  IV U91726 ( .A(n71493), .Z(n73368) );
  IV U91727 ( .A(n71494), .Z(n71496) );
  NOR U91728 ( .A(n71496), .B(n71495), .Z(n76880) );
  NOR U91729 ( .A(n76880), .B(n78769), .Z(n73367) );
  IV U91730 ( .A(n71497), .Z(n71498) );
  NOR U91731 ( .A(n71499), .B(n71498), .Z(n76884) );
  IV U91732 ( .A(n71500), .Z(n71502) );
  NOR U91733 ( .A(n71502), .B(n71501), .Z(n76882) );
  NOR U91734 ( .A(n76884), .B(n76882), .Z(n73366) );
  IV U91735 ( .A(n71503), .Z(n71504) );
  NOR U91736 ( .A(n71504), .B(n73357), .Z(n78738) );
  IV U91737 ( .A(n71505), .Z(n71506) );
  NOR U91738 ( .A(n71506), .B(n71511), .Z(n76890) );
  IV U91739 ( .A(n71507), .Z(n71508) );
  NOR U91740 ( .A(n71509), .B(n71508), .Z(n76897) );
  IV U91741 ( .A(n71510), .Z(n71512) );
  NOR U91742 ( .A(n71512), .B(n71511), .Z(n76894) );
  NOR U91743 ( .A(n76897), .B(n76894), .Z(n73348) );
  IV U91744 ( .A(n71513), .Z(n71515) );
  NOR U91745 ( .A(n71515), .B(n71514), .Z(n73346) );
  IV U91746 ( .A(n73346), .Z(n73341) );
  IV U91747 ( .A(n71516), .Z(n71518) );
  NOR U91748 ( .A(n71518), .B(n71517), .Z(n78716) );
  IV U91749 ( .A(n71519), .Z(n71520) );
  NOR U91750 ( .A(n71520), .B(n76921), .Z(n76917) );
  NOR U91751 ( .A(n71521), .B(n76929), .Z(n71524) );
  NOR U91752 ( .A(n71522), .B(n76921), .Z(n71523) );
  NOR U91753 ( .A(n71524), .B(n71523), .Z(n71525) );
  IV U91754 ( .A(n71525), .Z(n73310) );
  IV U91755 ( .A(n71526), .Z(n71528) );
  NOR U91756 ( .A(n71528), .B(n71527), .Z(n82619) );
  IV U91757 ( .A(n71529), .Z(n71531) );
  NOR U91758 ( .A(n71531), .B(n71530), .Z(n82612) );
  NOR U91759 ( .A(n82619), .B(n82612), .Z(n78703) );
  IV U91760 ( .A(n71532), .Z(n71533) );
  NOR U91761 ( .A(n71534), .B(n71533), .Z(n76940) );
  IV U91762 ( .A(n71535), .Z(n71536) );
  NOR U91763 ( .A(n71537), .B(n71536), .Z(n76935) );
  NOR U91764 ( .A(n76940), .B(n76935), .Z(n73309) );
  IV U91765 ( .A(n71538), .Z(n71539) );
  NOR U91766 ( .A(n71540), .B(n71539), .Z(n78690) );
  IV U91767 ( .A(n71541), .Z(n71542) );
  NOR U91768 ( .A(n71543), .B(n71542), .Z(n76938) );
  NOR U91769 ( .A(n78690), .B(n76938), .Z(n73308) );
  IV U91770 ( .A(n71544), .Z(n71546) );
  NOR U91771 ( .A(n71546), .B(n71545), .Z(n71547) );
  IV U91772 ( .A(n71547), .Z(n73293) );
  IV U91773 ( .A(n71548), .Z(n71549) );
  NOR U91774 ( .A(n73267), .B(n71549), .Z(n76949) );
  IV U91775 ( .A(n71550), .Z(n71551) );
  NOR U91776 ( .A(n71552), .B(n71551), .Z(n76962) );
  IV U91777 ( .A(n71553), .Z(n71555) );
  NOR U91778 ( .A(n71555), .B(n71554), .Z(n76959) );
  NOR U91779 ( .A(n76962), .B(n76959), .Z(n73258) );
  IV U91780 ( .A(n71556), .Z(n71558) );
  NOR U91781 ( .A(n71558), .B(n71557), .Z(n76968) );
  IV U91782 ( .A(n71559), .Z(n71561) );
  NOR U91783 ( .A(n71561), .B(n71560), .Z(n76966) );
  NOR U91784 ( .A(n76968), .B(n76966), .Z(n73257) );
  IV U91785 ( .A(n71562), .Z(n71563) );
  NOR U91786 ( .A(n71564), .B(n71563), .Z(n76974) );
  IV U91787 ( .A(n71565), .Z(n71567) );
  NOR U91788 ( .A(n71567), .B(n71566), .Z(n76971) );
  NOR U91789 ( .A(n76974), .B(n76971), .Z(n73256) );
  IV U91790 ( .A(n71568), .Z(n71569) );
  NOR U91791 ( .A(n71570), .B(n71569), .Z(n76975) );
  IV U91792 ( .A(n71571), .Z(n71573) );
  NOR U91793 ( .A(n71573), .B(n71572), .Z(n76981) );
  IV U91794 ( .A(n71574), .Z(n71575) );
  NOR U91795 ( .A(n71576), .B(n71575), .Z(n76979) );
  NOR U91796 ( .A(n76981), .B(n76979), .Z(n73255) );
  IV U91797 ( .A(n71577), .Z(n71578) );
  NOR U91798 ( .A(n71579), .B(n71578), .Z(n82686) );
  IV U91799 ( .A(n71580), .Z(n71582) );
  NOR U91800 ( .A(n71582), .B(n71581), .Z(n84420) );
  NOR U91801 ( .A(n82686), .B(n84420), .Z(n76986) );
  IV U91802 ( .A(n76986), .Z(n71583) );
  NOR U91803 ( .A(n71583), .B(n76984), .Z(n73254) );
  IV U91804 ( .A(n71584), .Z(n71586) );
  NOR U91805 ( .A(n71586), .B(n71585), .Z(n76996) );
  IV U91806 ( .A(n71587), .Z(n71588) );
  NOR U91807 ( .A(n71588), .B(n73252), .Z(n76994) );
  NOR U91808 ( .A(n76996), .B(n76994), .Z(n73246) );
  IV U91809 ( .A(n71589), .Z(n71590) );
  NOR U91810 ( .A(n71592), .B(n71590), .Z(n77002) );
  IV U91811 ( .A(n71591), .Z(n71593) );
  NOR U91812 ( .A(n71593), .B(n71592), .Z(n76999) );
  IV U91813 ( .A(n71594), .Z(n71595) );
  NOR U91814 ( .A(n71596), .B(n71595), .Z(n77007) );
  IV U91815 ( .A(n71597), .Z(n71598) );
  NOR U91816 ( .A(n71599), .B(n71598), .Z(n77012) );
  NOR U91817 ( .A(n77007), .B(n77012), .Z(n73245) );
  IV U91818 ( .A(n71600), .Z(n71604) );
  NOR U91819 ( .A(n71604), .B(n71601), .Z(n77020) );
  IV U91820 ( .A(n71602), .Z(n71603) );
  NOR U91821 ( .A(n71604), .B(n71603), .Z(n77009) );
  NOR U91822 ( .A(n77020), .B(n77009), .Z(n73244) );
  IV U91823 ( .A(n71605), .Z(n71606) );
  NOR U91824 ( .A(n71607), .B(n71606), .Z(n77040) );
  IV U91825 ( .A(n71608), .Z(n71609) );
  NOR U91826 ( .A(n71610), .B(n71609), .Z(n77036) );
  NOR U91827 ( .A(n77040), .B(n77036), .Z(n73221) );
  IV U91828 ( .A(n71611), .Z(n71613) );
  IV U91829 ( .A(n71612), .Z(n73206) );
  NOR U91830 ( .A(n71613), .B(n73206), .Z(n77055) );
  IV U91831 ( .A(n77055), .Z(n77057) );
  IV U91832 ( .A(n71614), .Z(n71615) );
  NOR U91833 ( .A(n71616), .B(n71615), .Z(n77066) );
  NOR U91834 ( .A(n71618), .B(n71617), .Z(n77063) );
  NOR U91835 ( .A(n77066), .B(n77063), .Z(n73200) );
  IV U91836 ( .A(n71619), .Z(n71620) );
  NOR U91837 ( .A(n71621), .B(n71620), .Z(n77068) );
  IV U91838 ( .A(n71622), .Z(n71623) );
  NOR U91839 ( .A(n71625), .B(n71623), .Z(n78653) );
  IV U91840 ( .A(n71624), .Z(n71626) );
  NOR U91841 ( .A(n71626), .B(n71625), .Z(n77079) );
  NOR U91842 ( .A(n78653), .B(n77079), .Z(n73187) );
  IV U91843 ( .A(n71627), .Z(n71628) );
  NOR U91844 ( .A(n73164), .B(n71628), .Z(n78641) );
  IV U91845 ( .A(n71629), .Z(n71635) );
  IV U91846 ( .A(n71630), .Z(n71631) );
  NOR U91847 ( .A(n71635), .B(n71631), .Z(n78638) );
  IV U91848 ( .A(n71632), .Z(n71633) );
  NOR U91849 ( .A(n71633), .B(n71638), .Z(n84348) );
  IV U91850 ( .A(n71634), .Z(n71636) );
  NOR U91851 ( .A(n71636), .B(n71635), .Z(n77081) );
  NOR U91852 ( .A(n84348), .B(n77081), .Z(n73161) );
  IV U91853 ( .A(n71637), .Z(n71639) );
  NOR U91854 ( .A(n71639), .B(n71638), .Z(n84343) );
  NOR U91855 ( .A(n71641), .B(n71640), .Z(n78609) );
  IV U91856 ( .A(n71642), .Z(n71643) );
  NOR U91857 ( .A(n71643), .B(n73127), .Z(n71644) );
  IV U91858 ( .A(n71644), .Z(n77091) );
  IV U91859 ( .A(n71645), .Z(n71646) );
  NOR U91860 ( .A(n71648), .B(n71646), .Z(n77103) );
  IV U91861 ( .A(n71647), .Z(n71649) );
  NOR U91862 ( .A(n71649), .B(n71648), .Z(n77097) );
  NOR U91863 ( .A(n77103), .B(n77097), .Z(n73122) );
  IV U91864 ( .A(n71650), .Z(n71651) );
  NOR U91865 ( .A(n71652), .B(n71651), .Z(n77106) );
  NOR U91866 ( .A(n77108), .B(n77106), .Z(n73121) );
  IV U91867 ( .A(n71653), .Z(n71658) );
  IV U91868 ( .A(n71654), .Z(n71655) );
  NOR U91869 ( .A(n71658), .B(n71655), .Z(n77122) );
  IV U91870 ( .A(n71656), .Z(n71657) );
  NOR U91871 ( .A(n71658), .B(n71657), .Z(n77131) );
  IV U91872 ( .A(n71659), .Z(n71662) );
  NOR U91873 ( .A(n71660), .B(n73107), .Z(n71661) );
  IV U91874 ( .A(n71661), .Z(n73103) );
  NOR U91875 ( .A(n71662), .B(n73103), .Z(n78598) );
  IV U91876 ( .A(n71663), .Z(n77136) );
  NOR U91877 ( .A(n71664), .B(n77136), .Z(n71668) );
  NOR U91878 ( .A(n71665), .B(n73094), .Z(n71666) );
  IV U91879 ( .A(n71666), .Z(n78591) );
  NOR U91880 ( .A(n71667), .B(n78591), .Z(n77139) );
  NOR U91881 ( .A(n71668), .B(n77139), .Z(n73101) );
  NOR U91882 ( .A(n71669), .B(n78576), .Z(n73088) );
  IV U91883 ( .A(n71670), .Z(n71677) );
  IV U91884 ( .A(n71671), .Z(n71672) );
  NOR U91885 ( .A(n71677), .B(n71672), .Z(n78573) );
  IV U91886 ( .A(n71673), .Z(n71674) );
  NOR U91887 ( .A(n71675), .B(n71674), .Z(n78580) );
  NOR U91888 ( .A(n78573), .B(n78580), .Z(n73076) );
  IV U91889 ( .A(n71676), .Z(n71678) );
  NOR U91890 ( .A(n71678), .B(n71677), .Z(n71679) );
  IV U91891 ( .A(n71679), .Z(n77154) );
  IV U91892 ( .A(n71680), .Z(n71681) );
  NOR U91893 ( .A(n71681), .B(n71687), .Z(n77151) );
  IV U91894 ( .A(n71682), .Z(n71683) );
  NOR U91895 ( .A(n71684), .B(n71683), .Z(n77161) );
  IV U91896 ( .A(n71685), .Z(n71686) );
  NOR U91897 ( .A(n71687), .B(n71686), .Z(n77157) );
  NOR U91898 ( .A(n77161), .B(n77157), .Z(n73074) );
  IV U91899 ( .A(n71688), .Z(n71689) );
  NOR U91900 ( .A(n71690), .B(n71689), .Z(n73072) );
  IV U91901 ( .A(n73072), .Z(n73066) );
  IV U91902 ( .A(n78564), .Z(n71691) );
  NOR U91903 ( .A(n71691), .B(n78566), .Z(n73070) );
  IV U91904 ( .A(n71692), .Z(n71693) );
  NOR U91905 ( .A(n71693), .B(n73056), .Z(n77168) );
  IV U91906 ( .A(n71694), .Z(n71696) );
  NOR U91907 ( .A(n71696), .B(n71695), .Z(n73051) );
  IV U91908 ( .A(n71697), .Z(n71699) );
  NOR U91909 ( .A(n71699), .B(n71698), .Z(n78533) );
  NOR U91910 ( .A(n71700), .B(n77173), .Z(n71704) );
  IV U91911 ( .A(n71701), .Z(n71703) );
  NOR U91912 ( .A(n71703), .B(n71702), .Z(n78530) );
  NOR U91913 ( .A(n71704), .B(n78530), .Z(n73034) );
  IV U91914 ( .A(n71705), .Z(n71707) );
  IV U91915 ( .A(n71706), .Z(n73030) );
  NOR U91916 ( .A(n71707), .B(n73030), .Z(n77183) );
  IV U91917 ( .A(n71708), .Z(n71709) );
  NOR U91918 ( .A(n73028), .B(n71709), .Z(n78525) );
  IV U91919 ( .A(n71710), .Z(n71711) );
  NOR U91920 ( .A(n71712), .B(n71711), .Z(n73023) );
  IV U91921 ( .A(n73023), .Z(n73010) );
  IV U91922 ( .A(n71713), .Z(n71714) );
  NOR U91923 ( .A(n71720), .B(n71714), .Z(n71715) );
  IV U91924 ( .A(n71715), .Z(n78515) );
  IV U91925 ( .A(n71716), .Z(n71718) );
  NOR U91926 ( .A(n71718), .B(n71717), .Z(n78511) );
  IV U91927 ( .A(n71719), .Z(n71721) );
  NOR U91928 ( .A(n71721), .B(n71720), .Z(n78517) );
  NOR U91929 ( .A(n78511), .B(n78517), .Z(n73009) );
  IV U91930 ( .A(n71722), .Z(n72987) );
  IV U91931 ( .A(n71723), .Z(n71724) );
  NOR U91932 ( .A(n72987), .B(n71724), .Z(n78499) );
  IV U91933 ( .A(n71725), .Z(n71726) );
  NOR U91934 ( .A(n71727), .B(n71726), .Z(n77199) );
  IV U91935 ( .A(n71728), .Z(n71730) );
  NOR U91936 ( .A(n71730), .B(n71729), .Z(n78491) );
  NOR U91937 ( .A(n77199), .B(n78491), .Z(n71731) );
  IV U91938 ( .A(n71731), .Z(n72982) );
  IV U91939 ( .A(n71732), .Z(n71734) );
  NOR U91940 ( .A(n71734), .B(n71733), .Z(n78483) );
  IV U91941 ( .A(n71735), .Z(n71736) );
  NOR U91942 ( .A(n71736), .B(n71738), .Z(n77203) );
  NOR U91943 ( .A(n78483), .B(n77203), .Z(n72974) );
  IV U91944 ( .A(n71737), .Z(n71739) );
  NOR U91945 ( .A(n71739), .B(n71738), .Z(n77207) );
  IV U91946 ( .A(n71740), .Z(n71741) );
  NOR U91947 ( .A(n71741), .B(n72971), .Z(n78472) );
  IV U91948 ( .A(n71742), .Z(n71743) );
  NOR U91949 ( .A(n71747), .B(n71743), .Z(n71744) );
  IV U91950 ( .A(n71744), .Z(n77221) );
  IV U91951 ( .A(n71745), .Z(n71746) );
  NOR U91952 ( .A(n71747), .B(n71746), .Z(n82934) );
  IV U91953 ( .A(n71748), .Z(n71750) );
  IV U91954 ( .A(n71749), .Z(n71752) );
  NOR U91955 ( .A(n71750), .B(n71752), .Z(n84225) );
  NOR U91956 ( .A(n82934), .B(n84225), .Z(n77225) );
  IV U91957 ( .A(n71751), .Z(n71753) );
  NOR U91958 ( .A(n71753), .B(n71752), .Z(n77227) );
  NOR U91959 ( .A(n71754), .B(n77227), .Z(n72957) );
  IV U91960 ( .A(n71755), .Z(n71756) );
  NOR U91961 ( .A(n71757), .B(n71756), .Z(n84202) );
  IV U91962 ( .A(n71758), .Z(n71759) );
  NOR U91963 ( .A(n71760), .B(n71759), .Z(n84196) );
  NOR U91964 ( .A(n84202), .B(n84196), .Z(n78462) );
  IV U91965 ( .A(n71761), .Z(n71762) );
  NOR U91966 ( .A(n71762), .B(n72940), .Z(n71763) );
  IV U91967 ( .A(n71763), .Z(n78456) );
  IV U91968 ( .A(n71764), .Z(n71766) );
  NOR U91969 ( .A(n71766), .B(n71765), .Z(n78449) );
  IV U91970 ( .A(n71767), .Z(n71769) );
  NOR U91971 ( .A(n71769), .B(n71768), .Z(n78452) );
  NOR U91972 ( .A(n78449), .B(n78452), .Z(n72934) );
  NOR U91973 ( .A(n78442), .B(n78435), .Z(n72933) );
  IV U91974 ( .A(n71770), .Z(n71771) );
  NOR U91975 ( .A(n71771), .B(n72925), .Z(n78428) );
  IV U91976 ( .A(n71772), .Z(n71773) );
  NOR U91977 ( .A(n71774), .B(n71773), .Z(n78396) );
  IV U91978 ( .A(n71775), .Z(n71779) );
  IV U91979 ( .A(n71776), .Z(n72911) );
  NOR U91980 ( .A(n71777), .B(n72911), .Z(n71778) );
  IV U91981 ( .A(n71778), .Z(n72908) );
  NOR U91982 ( .A(n71779), .B(n72908), .Z(n77256) );
  IV U91983 ( .A(n71780), .Z(n71781) );
  NOR U91984 ( .A(n72911), .B(n71781), .Z(n78382) );
  IV U91985 ( .A(n71782), .Z(n71783) );
  NOR U91986 ( .A(n71788), .B(n71783), .Z(n78379) );
  IV U91987 ( .A(n71784), .Z(n71785) );
  NOR U91988 ( .A(n71786), .B(n71785), .Z(n82976) );
  IV U91989 ( .A(n71787), .Z(n71789) );
  NOR U91990 ( .A(n71789), .B(n71788), .Z(n84173) );
  NOR U91991 ( .A(n82976), .B(n84173), .Z(n78376) );
  IV U91992 ( .A(n71790), .Z(n71792) );
  NOR U91993 ( .A(n71792), .B(n71791), .Z(n78373) );
  IV U91994 ( .A(n71793), .Z(n71795) );
  NOR U91995 ( .A(n71795), .B(n71794), .Z(n78363) );
  IV U91996 ( .A(n71796), .Z(n71797) );
  NOR U91997 ( .A(n71798), .B(n71797), .Z(n78355) );
  IV U91998 ( .A(n71799), .Z(n71801) );
  IV U91999 ( .A(n71800), .Z(n71806) );
  NOR U92000 ( .A(n71801), .B(n71806), .Z(n78357) );
  NOR U92001 ( .A(n78355), .B(n78357), .Z(n72905) );
  IV U92002 ( .A(n71802), .Z(n71803) );
  NOR U92003 ( .A(n71808), .B(n71803), .Z(n77265) );
  IV U92004 ( .A(n71804), .Z(n71805) );
  NOR U92005 ( .A(n71806), .B(n71805), .Z(n78350) );
  NOR U92006 ( .A(n77265), .B(n78350), .Z(n72904) );
  IV U92007 ( .A(n71807), .Z(n71809) );
  NOR U92008 ( .A(n71809), .B(n71808), .Z(n77262) );
  IV U92009 ( .A(n71810), .Z(n71811) );
  NOR U92010 ( .A(n71817), .B(n71811), .Z(n78341) );
  IV U92011 ( .A(n71812), .Z(n71813) );
  NOR U92012 ( .A(n71814), .B(n71813), .Z(n77269) );
  IV U92013 ( .A(n71815), .Z(n71816) );
  NOR U92014 ( .A(n71817), .B(n71816), .Z(n78337) );
  NOR U92015 ( .A(n77269), .B(n78337), .Z(n72895) );
  IV U92016 ( .A(n71818), .Z(n71820) );
  NOR U92017 ( .A(n71820), .B(n71819), .Z(n72893) );
  IV U92018 ( .A(n72893), .Z(n72886) );
  IV U92019 ( .A(n71821), .Z(n71822) );
  NOR U92020 ( .A(n72889), .B(n71822), .Z(n72882) );
  IV U92021 ( .A(n71823), .Z(n71824) );
  NOR U92022 ( .A(n71825), .B(n71824), .Z(n83029) );
  NOR U92023 ( .A(n83029), .B(n71826), .Z(n77277) );
  NOR U92024 ( .A(n72857), .B(n72855), .Z(n72854) );
  IV U92025 ( .A(n71827), .Z(n72852) );
  IV U92026 ( .A(n71828), .Z(n71829) );
  NOR U92027 ( .A(n72852), .B(n71829), .Z(n77293) );
  IV U92028 ( .A(n71830), .Z(n71831) );
  NOR U92029 ( .A(n71832), .B(n71831), .Z(n77300) );
  IV U92030 ( .A(n71833), .Z(n71834) );
  NOR U92031 ( .A(n72844), .B(n71834), .Z(n78318) );
  IV U92032 ( .A(n71835), .Z(n71836) );
  NOR U92033 ( .A(n71836), .B(n72846), .Z(n78310) );
  IV U92034 ( .A(n71837), .Z(n71838) );
  NOR U92035 ( .A(n71838), .B(n72815), .Z(n78283) );
  IV U92036 ( .A(n71839), .Z(n71840) );
  NOR U92037 ( .A(n71841), .B(n71840), .Z(n77314) );
  IV U92038 ( .A(n71842), .Z(n71844) );
  IV U92039 ( .A(n71843), .Z(n71848) );
  NOR U92040 ( .A(n71844), .B(n71848), .Z(n78261) );
  NOR U92041 ( .A(n77314), .B(n78261), .Z(n72795) );
  IV U92042 ( .A(n71845), .Z(n71846) );
  NOR U92043 ( .A(n71846), .B(n71848), .Z(n77319) );
  IV U92044 ( .A(n71847), .Z(n71849) );
  NOR U92045 ( .A(n71849), .B(n71848), .Z(n77316) );
  IV U92046 ( .A(n71850), .Z(n71852) );
  NOR U92047 ( .A(n71852), .B(n71851), .Z(n77322) );
  IV U92048 ( .A(n71853), .Z(n71857) );
  NOR U92049 ( .A(n71855), .B(n71854), .Z(n71856) );
  IV U92050 ( .A(n71856), .Z(n72784) );
  NOR U92051 ( .A(n71857), .B(n72784), .Z(n72779) );
  IV U92052 ( .A(n71858), .Z(n71859) );
  NOR U92053 ( .A(n71859), .B(n72756), .Z(n78231) );
  IV U92054 ( .A(n71860), .Z(n72762) );
  NOR U92055 ( .A(n71861), .B(n72762), .Z(n77343) );
  NOR U92056 ( .A(n78231), .B(n77343), .Z(n72759) );
  IV U92057 ( .A(n71862), .Z(n71863) );
  NOR U92058 ( .A(n71863), .B(n71865), .Z(n77351) );
  IV U92059 ( .A(n71864), .Z(n71866) );
  NOR U92060 ( .A(n71866), .B(n71865), .Z(n72747) );
  IV U92061 ( .A(n71867), .Z(n71868) );
  NOR U92062 ( .A(n71869), .B(n71868), .Z(n78216) );
  IV U92063 ( .A(n71870), .Z(n71871) );
  NOR U92064 ( .A(n71872), .B(n71871), .Z(n78212) );
  IV U92065 ( .A(n71873), .Z(n71874) );
  NOR U92066 ( .A(n71874), .B(n78209), .Z(n71875) );
  NOR U92067 ( .A(n78212), .B(n71875), .Z(n72730) );
  IV U92068 ( .A(n71876), .Z(n71877) );
  NOR U92069 ( .A(n71878), .B(n71877), .Z(n71879) );
  IV U92070 ( .A(n71879), .Z(n72725) );
  IV U92071 ( .A(n71880), .Z(n71881) );
  NOR U92072 ( .A(n71881), .B(n71886), .Z(n77382) );
  IV U92073 ( .A(n71882), .Z(n71890) );
  IV U92074 ( .A(n71883), .Z(n71884) );
  NOR U92075 ( .A(n71890), .B(n71884), .Z(n83996) );
  IV U92076 ( .A(n71885), .Z(n71887) );
  NOR U92077 ( .A(n71887), .B(n71886), .Z(n84010) );
  NOR U92078 ( .A(n83996), .B(n84010), .Z(n77381) );
  IV U92079 ( .A(n71888), .Z(n71889) );
  NOR U92080 ( .A(n71890), .B(n71889), .Z(n77389) );
  IV U92081 ( .A(n71891), .Z(n71895) );
  IV U92082 ( .A(n71892), .Z(n71893) );
  NOR U92083 ( .A(n71895), .B(n71893), .Z(n77394) );
  NOR U92084 ( .A(n71895), .B(n71894), .Z(n77398) );
  IV U92085 ( .A(n71896), .Z(n71897) );
  NOR U92086 ( .A(n71897), .B(n72705), .Z(n77401) );
  IV U92087 ( .A(n71898), .Z(n71899) );
  NOR U92088 ( .A(n71900), .B(n71899), .Z(n72698) );
  IV U92089 ( .A(n72698), .Z(n72691) );
  IV U92090 ( .A(n71901), .Z(n71902) );
  NOR U92091 ( .A(n71905), .B(n71902), .Z(n78199) );
  IV U92092 ( .A(n71903), .Z(n71904) );
  NOR U92093 ( .A(n71905), .B(n71904), .Z(n78196) );
  IV U92094 ( .A(n71906), .Z(n71907) );
  NOR U92095 ( .A(n71908), .B(n71907), .Z(n77415) );
  IV U92096 ( .A(n71909), .Z(n71910) );
  NOR U92097 ( .A(n71910), .B(n72687), .Z(n78181) );
  NOR U92098 ( .A(n77415), .B(n78181), .Z(n72683) );
  IV U92099 ( .A(n71911), .Z(n71912) );
  NOR U92100 ( .A(n71915), .B(n71912), .Z(n77412) );
  IV U92101 ( .A(n71913), .Z(n71914) );
  NOR U92102 ( .A(n71915), .B(n71914), .Z(n77409) );
  IV U92103 ( .A(n71916), .Z(n71918) );
  NOR U92104 ( .A(n71918), .B(n71917), .Z(n78159) );
  IV U92105 ( .A(n71919), .Z(n71920) );
  NOR U92106 ( .A(n71920), .B(n72664), .Z(n78155) );
  IV U92107 ( .A(n71921), .Z(n71923) );
  NOR U92108 ( .A(n71923), .B(n71922), .Z(n78162) );
  NOR U92109 ( .A(n78155), .B(n78162), .Z(n72667) );
  IV U92110 ( .A(n71924), .Z(n71926) );
  NOR U92111 ( .A(n71926), .B(n71925), .Z(n78147) );
  IV U92112 ( .A(n71927), .Z(n71928) );
  NOR U92113 ( .A(n71928), .B(n72657), .Z(n78142) );
  IV U92114 ( .A(n71929), .Z(n71931) );
  NOR U92115 ( .A(n71931), .B(n71930), .Z(n77426) );
  XOR U92116 ( .A(n78142), .B(n77426), .Z(n71932) );
  NOR U92117 ( .A(n78147), .B(n71932), .Z(n72659) );
  NOR U92118 ( .A(n77437), .B(n77432), .Z(n72648) );
  IV U92119 ( .A(n71933), .Z(n71941) );
  IV U92120 ( .A(n71934), .Z(n71935) );
  NOR U92121 ( .A(n71941), .B(n71935), .Z(n83219) );
  IV U92122 ( .A(n71936), .Z(n71937) );
  NOR U92123 ( .A(n71938), .B(n71937), .Z(n83215) );
  NOR U92124 ( .A(n83219), .B(n83215), .Z(n78122) );
  IV U92125 ( .A(n71939), .Z(n71940) );
  NOR U92126 ( .A(n71941), .B(n71940), .Z(n78119) );
  IV U92127 ( .A(n71942), .Z(n71944) );
  NOR U92128 ( .A(n71944), .B(n71943), .Z(n78113) );
  IV U92129 ( .A(n71945), .Z(n71946) );
  NOR U92130 ( .A(n72638), .B(n71946), .Z(n78116) );
  NOR U92131 ( .A(n78113), .B(n78116), .Z(n72642) );
  IV U92132 ( .A(n71947), .Z(n71948) );
  NOR U92133 ( .A(n71948), .B(n72632), .Z(n71949) );
  IV U92134 ( .A(n71949), .Z(n78106) );
  XOR U92135 ( .A(n72630), .B(n72632), .Z(n71952) );
  IV U92136 ( .A(n71950), .Z(n71951) );
  NOR U92137 ( .A(n71952), .B(n71951), .Z(n72635) );
  IV U92138 ( .A(n72635), .Z(n72629) );
  IV U92139 ( .A(n71953), .Z(n71954) );
  NOR U92140 ( .A(n71955), .B(n71954), .Z(n77441) );
  IV U92141 ( .A(n71956), .Z(n71958) );
  NOR U92142 ( .A(n71958), .B(n71957), .Z(n77446) );
  IV U92143 ( .A(n71959), .Z(n71961) );
  IV U92144 ( .A(n71960), .Z(n71965) );
  NOR U92145 ( .A(n71961), .B(n71965), .Z(n77449) );
  NOR U92146 ( .A(n71963), .B(n71962), .Z(n83239) );
  IV U92147 ( .A(n71964), .Z(n71966) );
  NOR U92148 ( .A(n71966), .B(n71965), .Z(n83234) );
  NOR U92149 ( .A(n83239), .B(n83234), .Z(n77448) );
  IV U92150 ( .A(n77448), .Z(n72619) );
  IV U92151 ( .A(n71967), .Z(n71969) );
  NOR U92152 ( .A(n71969), .B(n71968), .Z(n72591) );
  IV U92153 ( .A(n71970), .Z(n72574) );
  IV U92154 ( .A(n71971), .Z(n71973) );
  IV U92155 ( .A(n71972), .Z(n71975) );
  NOR U92156 ( .A(n71973), .B(n71975), .Z(n77457) );
  IV U92157 ( .A(n71974), .Z(n71978) );
  NOR U92158 ( .A(n71976), .B(n71975), .Z(n71977) );
  IV U92159 ( .A(n71977), .Z(n71981) );
  NOR U92160 ( .A(n71978), .B(n71981), .Z(n77459) );
  NOR U92161 ( .A(n77457), .B(n77459), .Z(n72571) );
  NOR U92162 ( .A(n71979), .B(n78061), .Z(n71983) );
  IV U92163 ( .A(n71980), .Z(n71982) );
  NOR U92164 ( .A(n71982), .B(n71981), .Z(n78065) );
  NOR U92165 ( .A(n71983), .B(n78065), .Z(n71984) );
  IV U92166 ( .A(n71984), .Z(n72570) );
  IV U92167 ( .A(n71985), .Z(n71986) );
  NOR U92168 ( .A(n71987), .B(n71986), .Z(n83869) );
  IV U92169 ( .A(n71988), .Z(n71990) );
  NOR U92170 ( .A(n71990), .B(n71989), .Z(n83266) );
  NOR U92171 ( .A(n83869), .B(n83266), .Z(n77465) );
  IV U92172 ( .A(n71991), .Z(n71992) );
  NOR U92173 ( .A(n71992), .B(n71994), .Z(n77470) );
  IV U92174 ( .A(n71993), .Z(n71995) );
  NOR U92175 ( .A(n71995), .B(n71994), .Z(n71996) );
  IV U92176 ( .A(n71996), .Z(n77468) );
  IV U92177 ( .A(n71997), .Z(n71998) );
  NOR U92178 ( .A(n71999), .B(n71998), .Z(n77473) );
  IV U92179 ( .A(n72000), .Z(n72563) );
  IV U92180 ( .A(n72001), .Z(n72002) );
  NOR U92181 ( .A(n72563), .B(n72002), .Z(n77478) );
  NOR U92182 ( .A(n77473), .B(n77478), .Z(n72568) );
  IV U92183 ( .A(n72003), .Z(n72005) );
  NOR U92184 ( .A(n72005), .B(n72004), .Z(n72006) );
  IV U92185 ( .A(n72006), .Z(n72557) );
  IV U92186 ( .A(n72007), .Z(n72012) );
  IV U92187 ( .A(n72008), .Z(n72009) );
  NOR U92188 ( .A(n72012), .B(n72009), .Z(n78047) );
  IV U92189 ( .A(n72010), .Z(n72011) );
  NOR U92190 ( .A(n72012), .B(n72011), .Z(n78042) );
  IV U92191 ( .A(n72013), .Z(n72014) );
  NOR U92192 ( .A(n72014), .B(n72544), .Z(n77488) );
  IV U92193 ( .A(n72015), .Z(n72016) );
  NOR U92194 ( .A(n72017), .B(n72016), .Z(n77493) );
  IV U92195 ( .A(n72018), .Z(n72020) );
  NOR U92196 ( .A(n72020), .B(n72019), .Z(n77491) );
  NOR U92197 ( .A(n77493), .B(n77491), .Z(n72541) );
  IV U92198 ( .A(n72021), .Z(n72022) );
  NOR U92199 ( .A(n72022), .B(n72537), .Z(n77498) );
  IV U92200 ( .A(n72023), .Z(n72025) );
  NOR U92201 ( .A(n72025), .B(n72024), .Z(n83310) );
  IV U92202 ( .A(n72026), .Z(n72027) );
  NOR U92203 ( .A(n72028), .B(n72027), .Z(n83839) );
  NOR U92204 ( .A(n83310), .B(n83839), .Z(n77502) );
  IV U92205 ( .A(n78030), .Z(n72528) );
  IV U92206 ( .A(n72029), .Z(n78029) );
  NOR U92207 ( .A(n72528), .B(n78029), .Z(n78022) );
  IV U92208 ( .A(n72030), .Z(n72032) );
  NOR U92209 ( .A(n72032), .B(n72031), .Z(n72033) );
  IV U92210 ( .A(n72033), .Z(n78020) );
  IV U92211 ( .A(n72034), .Z(n72035) );
  NOR U92212 ( .A(n72035), .B(n72037), .Z(n72039) );
  IV U92213 ( .A(n72036), .Z(n72038) );
  NOR U92214 ( .A(n72038), .B(n72037), .Z(n78016) );
  NOR U92215 ( .A(n72039), .B(n78016), .Z(n72525) );
  IV U92216 ( .A(n72040), .Z(n78004) );
  IV U92217 ( .A(n72041), .Z(n72042) );
  NOR U92218 ( .A(n72042), .B(n72511), .Z(n77995) );
  IV U92219 ( .A(n72043), .Z(n72044) );
  NOR U92220 ( .A(n72515), .B(n72044), .Z(n77532) );
  IV U92221 ( .A(n72045), .Z(n72047) );
  NOR U92222 ( .A(n72047), .B(n72046), .Z(n77969) );
  IV U92223 ( .A(n72048), .Z(n72053) );
  IV U92224 ( .A(n72049), .Z(n72050) );
  NOR U92225 ( .A(n72053), .B(n72050), .Z(n77962) );
  IV U92226 ( .A(n72051), .Z(n72052) );
  NOR U92227 ( .A(n72053), .B(n72052), .Z(n77965) );
  IV U92228 ( .A(n72054), .Z(n72055) );
  NOR U92229 ( .A(n72055), .B(n72487), .Z(n77957) );
  NOR U92230 ( .A(n77965), .B(n77957), .Z(n72499) );
  NOR U92231 ( .A(n72056), .B(n77932), .Z(n72482) );
  IV U92232 ( .A(n72057), .Z(n72059) );
  NOR U92233 ( .A(n72059), .B(n72058), .Z(n77937) );
  IV U92234 ( .A(n72060), .Z(n72062) );
  NOR U92235 ( .A(n72062), .B(n72061), .Z(n77942) );
  NOR U92236 ( .A(n77937), .B(n77942), .Z(n77935) );
  IV U92237 ( .A(n72063), .Z(n72064) );
  NOR U92238 ( .A(n72064), .B(n72479), .Z(n72065) );
  IV U92239 ( .A(n72065), .Z(n77540) );
  IV U92240 ( .A(n72066), .Z(n72067) );
  NOR U92241 ( .A(n72068), .B(n72067), .Z(n77547) );
  IV U92242 ( .A(n72069), .Z(n72071) );
  NOR U92243 ( .A(n72071), .B(n72070), .Z(n83390) );
  IV U92244 ( .A(n72072), .Z(n72073) );
  NOR U92245 ( .A(n72073), .B(n72443), .Z(n83385) );
  NOR U92246 ( .A(n83390), .B(n83385), .Z(n77880) );
  IV U92247 ( .A(n72074), .Z(n72075) );
  NOR U92248 ( .A(n72076), .B(n72075), .Z(n72077) );
  IV U92249 ( .A(n72077), .Z(n72414) );
  IV U92250 ( .A(n72078), .Z(n72079) );
  NOR U92251 ( .A(n72079), .B(n72413), .Z(n77574) );
  IV U92252 ( .A(n72080), .Z(n72081) );
  NOR U92253 ( .A(n72082), .B(n72081), .Z(n77592) );
  IV U92254 ( .A(n72083), .Z(n72085) );
  NOR U92255 ( .A(n72085), .B(n72084), .Z(n83461) );
  IV U92256 ( .A(n72086), .Z(n72088) );
  NOR U92257 ( .A(n72088), .B(n72087), .Z(n83457) );
  NOR U92258 ( .A(n83461), .B(n83457), .Z(n77853) );
  IV U92259 ( .A(n72089), .Z(n72091) );
  NOR U92260 ( .A(n72091), .B(n72090), .Z(n72354) );
  IV U92261 ( .A(n72092), .Z(n72093) );
  NOR U92262 ( .A(n72098), .B(n72093), .Z(n77602) );
  IV U92263 ( .A(n72094), .Z(n72095) );
  NOR U92264 ( .A(n72096), .B(n72095), .Z(n77613) );
  IV U92265 ( .A(n72097), .Z(n72099) );
  NOR U92266 ( .A(n72099), .B(n72098), .Z(n77608) );
  NOR U92267 ( .A(n77613), .B(n77608), .Z(n72337) );
  IV U92268 ( .A(n72100), .Z(n72102) );
  IV U92269 ( .A(n72101), .Z(n72104) );
  NOR U92270 ( .A(n72102), .B(n72104), .Z(n72333) );
  IV U92271 ( .A(n72103), .Z(n72105) );
  NOR U92272 ( .A(n72105), .B(n72104), .Z(n72331) );
  IV U92273 ( .A(n72331), .Z(n72324) );
  IV U92274 ( .A(n72106), .Z(n72107) );
  NOR U92275 ( .A(n72107), .B(n72109), .Z(n77628) );
  IV U92276 ( .A(n72108), .Z(n72110) );
  NOR U92277 ( .A(n72110), .B(n72109), .Z(n77635) );
  IV U92278 ( .A(n72111), .Z(n72112) );
  NOR U92279 ( .A(n72112), .B(n72295), .Z(n77828) );
  IV U92280 ( .A(n72113), .Z(n72117) );
  NOR U92281 ( .A(n72115), .B(n72114), .Z(n72116) );
  IV U92282 ( .A(n72116), .Z(n72278) );
  NOR U92283 ( .A(n72117), .B(n72278), .Z(n77819) );
  IV U92284 ( .A(n72118), .Z(n72119) );
  NOR U92285 ( .A(n72119), .B(n72121), .Z(n77808) );
  IV U92286 ( .A(n72120), .Z(n72122) );
  NOR U92287 ( .A(n72122), .B(n72121), .Z(n77805) );
  IV U92288 ( .A(n72123), .Z(n72124) );
  NOR U92289 ( .A(n72125), .B(n72124), .Z(n77660) );
  IV U92290 ( .A(n72126), .Z(n72127) );
  NOR U92291 ( .A(n72132), .B(n72127), .Z(n77798) );
  NOR U92292 ( .A(n77660), .B(n77798), .Z(n72274) );
  IV U92293 ( .A(n72128), .Z(n72129) );
  NOR U92294 ( .A(n72130), .B(n72129), .Z(n77783) );
  IV U92295 ( .A(n72131), .Z(n72133) );
  NOR U92296 ( .A(n72133), .B(n72132), .Z(n77801) );
  NOR U92297 ( .A(n77783), .B(n77801), .Z(n72273) );
  IV U92298 ( .A(n72134), .Z(n77774) );
  NOR U92299 ( .A(n72135), .B(n77774), .Z(n77787) );
  IV U92300 ( .A(n72136), .Z(n72137) );
  NOR U92301 ( .A(n72137), .B(n72142), .Z(n77662) );
  IV U92302 ( .A(n72138), .Z(n72140) );
  NOR U92303 ( .A(n72140), .B(n72139), .Z(n77767) );
  IV U92304 ( .A(n72141), .Z(n72143) );
  NOR U92305 ( .A(n72143), .B(n72142), .Z(n77769) );
  NOR U92306 ( .A(n77767), .B(n77769), .Z(n72272) );
  IV U92307 ( .A(n72144), .Z(n72145) );
  NOR U92308 ( .A(n72145), .B(n72151), .Z(n77758) );
  IV U92309 ( .A(n72146), .Z(n72147) );
  NOR U92310 ( .A(n72147), .B(n72151), .Z(n77668) );
  IV U92311 ( .A(n72148), .Z(n72149) );
  NOR U92312 ( .A(n72150), .B(n72149), .Z(n77671) );
  NOR U92313 ( .A(n72152), .B(n72151), .Z(n77666) );
  NOR U92314 ( .A(n77671), .B(n77666), .Z(n72264) );
  IV U92315 ( .A(n72153), .Z(n72154) );
  NOR U92316 ( .A(n72154), .B(n72260), .Z(n77748) );
  IV U92317 ( .A(n72155), .Z(n72156) );
  NOR U92318 ( .A(n72156), .B(n72260), .Z(n77674) );
  NOR U92319 ( .A(n77748), .B(n77674), .Z(n72263) );
  IV U92320 ( .A(n72157), .Z(n72158) );
  NOR U92321 ( .A(n72158), .B(n72249), .Z(n83623) );
  IV U92322 ( .A(n72159), .Z(n72161) );
  IV U92323 ( .A(n72160), .Z(n72257) );
  NOR U92324 ( .A(n72161), .B(n72257), .Z(n83559) );
  NOR U92325 ( .A(n83623), .B(n83559), .Z(n77676) );
  IV U92326 ( .A(n72162), .Z(n72163) );
  NOR U92327 ( .A(n72163), .B(n72169), .Z(n77680) );
  IV U92328 ( .A(n72164), .Z(n72166) );
  NOR U92329 ( .A(n72166), .B(n72165), .Z(n77690) );
  IV U92330 ( .A(n72167), .Z(n72168) );
  NOR U92331 ( .A(n72169), .B(n72168), .Z(n77687) );
  NOR U92332 ( .A(n77690), .B(n77687), .Z(n72244) );
  IV U92333 ( .A(n72170), .Z(n72171) );
  NOR U92334 ( .A(n72171), .B(n72177), .Z(n77723) );
  IV U92335 ( .A(n72172), .Z(n72174) );
  NOR U92336 ( .A(n72174), .B(n72173), .Z(n77696) );
  IV U92337 ( .A(n72175), .Z(n72176) );
  NOR U92338 ( .A(n72177), .B(n72176), .Z(n77693) );
  NOR U92339 ( .A(n77696), .B(n77693), .Z(n72225) );
  IV U92340 ( .A(n72178), .Z(n72181) );
  IV U92341 ( .A(n72179), .Z(n72180) );
  NOR U92342 ( .A(n72181), .B(n72180), .Z(n72186) );
  IV U92343 ( .A(n72182), .Z(n72183) );
  NOR U92344 ( .A(n72184), .B(n72183), .Z(n72185) );
  NOR U92345 ( .A(n72186), .B(n72185), .Z(n77702) );
  IV U92346 ( .A(n77702), .Z(n77700) );
  IV U92347 ( .A(n72191), .Z(n72187) );
  NOR U92348 ( .A(n72187), .B(n72189), .Z(n72195) );
  IV U92349 ( .A(n72188), .Z(n72193) );
  IV U92350 ( .A(n72189), .Z(n72190) );
  NOR U92351 ( .A(n72191), .B(n72190), .Z(n72192) );
  NOR U92352 ( .A(n72193), .B(n72192), .Z(n72194) );
  NOR U92353 ( .A(n72195), .B(n72194), .Z(n77701) );
  XOR U92354 ( .A(n77700), .B(n77701), .Z(n77712) );
  IV U92355 ( .A(n72196), .Z(n72197) );
  NOR U92356 ( .A(n72198), .B(n72197), .Z(n77710) );
  IV U92357 ( .A(n72199), .Z(n72200) );
  NOR U92358 ( .A(n72201), .B(n72200), .Z(n77703) );
  NOR U92359 ( .A(n77710), .B(n77703), .Z(n72202) );
  XOR U92360 ( .A(n77712), .B(n72202), .Z(n72203) );
  IV U92361 ( .A(n72203), .Z(n77709) );
  IV U92362 ( .A(n72204), .Z(n72215) );
  NOR U92363 ( .A(n77709), .B(n72215), .Z(n72205) );
  IV U92364 ( .A(n72205), .Z(n72210) );
  NOR U92365 ( .A(n72207), .B(n72206), .Z(n72208) );
  IV U92366 ( .A(n72208), .Z(n72209) );
  NOR U92367 ( .A(n72210), .B(n72209), .Z(n83581) );
  IV U92368 ( .A(n72211), .Z(n72213) );
  NOR U92369 ( .A(n72213), .B(n72212), .Z(n72223) );
  NOR U92370 ( .A(n72215), .B(n72214), .Z(n72216) );
  IV U92371 ( .A(n72216), .Z(n77719) );
  IV U92372 ( .A(n72217), .Z(n72218) );
  NOR U92373 ( .A(n72218), .B(n72220), .Z(n77707) );
  XOR U92374 ( .A(n77707), .B(n77709), .Z(n77717) );
  IV U92375 ( .A(n72219), .Z(n72221) );
  NOR U92376 ( .A(n72221), .B(n72220), .Z(n77715) );
  XOR U92377 ( .A(n77717), .B(n77715), .Z(n77718) );
  XOR U92378 ( .A(n77719), .B(n77718), .Z(n72222) );
  NOR U92379 ( .A(n72223), .B(n72222), .Z(n72224) );
  NOR U92380 ( .A(n83581), .B(n72224), .Z(n77694) );
  XOR U92381 ( .A(n72225), .B(n77694), .Z(n77724) );
  XOR U92382 ( .A(n77723), .B(n77724), .Z(n77728) );
  IV U92383 ( .A(n72226), .Z(n72230) );
  IV U92384 ( .A(n72227), .Z(n72235) );
  NOR U92385 ( .A(n72228), .B(n72235), .Z(n72229) );
  IV U92386 ( .A(n72229), .Z(n72232) );
  NOR U92387 ( .A(n72230), .B(n72232), .Z(n77726) );
  XOR U92388 ( .A(n77728), .B(n77726), .Z(n77733) );
  IV U92389 ( .A(n72231), .Z(n72233) );
  NOR U92390 ( .A(n72233), .B(n72232), .Z(n77731) );
  XOR U92391 ( .A(n77733), .B(n77731), .Z(n77736) );
  IV U92392 ( .A(n72234), .Z(n72236) );
  NOR U92393 ( .A(n72236), .B(n72235), .Z(n77734) );
  XOR U92394 ( .A(n77736), .B(n77734), .Z(n77742) );
  IV U92395 ( .A(n72237), .Z(n72238) );
  NOR U92396 ( .A(n72239), .B(n72238), .Z(n77739) );
  IV U92397 ( .A(n72240), .Z(n72242) );
  NOR U92398 ( .A(n72242), .B(n72241), .Z(n77741) );
  NOR U92399 ( .A(n77739), .B(n77741), .Z(n72243) );
  XOR U92400 ( .A(n77742), .B(n72243), .Z(n77686) );
  XOR U92401 ( .A(n72244), .B(n77686), .Z(n77682) );
  XOR U92402 ( .A(n77680), .B(n77682), .Z(n77684) );
  IV U92403 ( .A(n72245), .Z(n72246) );
  NOR U92404 ( .A(n72247), .B(n72246), .Z(n77683) );
  IV U92405 ( .A(n72248), .Z(n72250) );
  NOR U92406 ( .A(n72250), .B(n72249), .Z(n77677) );
  NOR U92407 ( .A(n77683), .B(n77677), .Z(n72251) );
  XOR U92408 ( .A(n77684), .B(n72251), .Z(n72252) );
  IV U92409 ( .A(n72252), .Z(n83561) );
  XOR U92410 ( .A(n77676), .B(n83561), .Z(n77751) );
  IV U92411 ( .A(n72253), .Z(n72254) );
  NOR U92412 ( .A(n83558), .B(n72254), .Z(n72258) );
  IV U92413 ( .A(n72255), .Z(n72256) );
  NOR U92414 ( .A(n72257), .B(n72256), .Z(n83638) );
  NOR U92415 ( .A(n72258), .B(n83638), .Z(n77752) );
  XOR U92416 ( .A(n77751), .B(n77752), .Z(n77749) );
  IV U92417 ( .A(n72259), .Z(n72261) );
  NOR U92418 ( .A(n72261), .B(n72260), .Z(n77746) );
  XOR U92419 ( .A(n77749), .B(n77746), .Z(n72262) );
  XOR U92420 ( .A(n72263), .B(n72262), .Z(n77665) );
  XOR U92421 ( .A(n72264), .B(n77665), .Z(n77670) );
  XOR U92422 ( .A(n77668), .B(n77670), .Z(n77760) );
  XOR U92423 ( .A(n77758), .B(n77760), .Z(n77762) );
  IV U92424 ( .A(n72265), .Z(n72266) );
  NOR U92425 ( .A(n72267), .B(n72266), .Z(n77755) );
  IV U92426 ( .A(n72268), .Z(n72270) );
  NOR U92427 ( .A(n72270), .B(n72269), .Z(n77761) );
  NOR U92428 ( .A(n77755), .B(n77761), .Z(n72271) );
  XOR U92429 ( .A(n77762), .B(n72271), .Z(n77766) );
  XOR U92430 ( .A(n72272), .B(n77766), .Z(n77773) );
  XOR U92431 ( .A(n77662), .B(n77773), .Z(n77788) );
  XOR U92432 ( .A(n77787), .B(n77788), .Z(n77802) );
  XOR U92433 ( .A(n72273), .B(n77802), .Z(n77659) );
  XOR U92434 ( .A(n72274), .B(n77659), .Z(n77807) );
  XOR U92435 ( .A(n77805), .B(n77807), .Z(n77810) );
  XOR U92436 ( .A(n77808), .B(n77810), .Z(n77818) );
  IV U92437 ( .A(n77818), .Z(n72282) );
  IV U92438 ( .A(n72275), .Z(n77656) );
  NOR U92439 ( .A(n77656), .B(n72276), .Z(n72280) );
  IV U92440 ( .A(n72277), .Z(n72279) );
  NOR U92441 ( .A(n72279), .B(n72278), .Z(n77816) );
  NOR U92442 ( .A(n72280), .B(n77816), .Z(n72281) );
  XOR U92443 ( .A(n72282), .B(n72281), .Z(n77821) );
  XOR U92444 ( .A(n77819), .B(n77821), .Z(n77823) );
  IV U92445 ( .A(n72283), .Z(n72284) );
  NOR U92446 ( .A(n72285), .B(n72284), .Z(n77822) );
  IV U92447 ( .A(n72286), .Z(n72288) );
  NOR U92448 ( .A(n72288), .B(n72287), .Z(n77653) );
  NOR U92449 ( .A(n77822), .B(n77653), .Z(n72289) );
  XOR U92450 ( .A(n77823), .B(n72289), .Z(n77647) );
  IV U92451 ( .A(n72290), .Z(n72292) );
  NOR U92452 ( .A(n72292), .B(n72291), .Z(n77650) );
  IV U92453 ( .A(n72293), .Z(n72294) );
  NOR U92454 ( .A(n72295), .B(n72294), .Z(n77648) );
  NOR U92455 ( .A(n77650), .B(n77648), .Z(n72296) );
  XOR U92456 ( .A(n77647), .B(n72296), .Z(n77829) );
  XOR U92457 ( .A(n77828), .B(n77829), .Z(n77833) );
  IV U92458 ( .A(n72297), .Z(n72299) );
  IV U92459 ( .A(n72298), .Z(n72301) );
  NOR U92460 ( .A(n72299), .B(n72301), .Z(n77831) );
  XOR U92461 ( .A(n77833), .B(n77831), .Z(n77643) );
  IV U92462 ( .A(n72300), .Z(n72302) );
  NOR U92463 ( .A(n72302), .B(n72301), .Z(n77641) );
  XOR U92464 ( .A(n77643), .B(n77641), .Z(n77645) );
  IV U92465 ( .A(n72303), .Z(n72304) );
  NOR U92466 ( .A(n72305), .B(n72304), .Z(n77644) );
  IV U92467 ( .A(n72306), .Z(n72308) );
  NOR U92468 ( .A(n72308), .B(n72307), .Z(n77638) );
  NOR U92469 ( .A(n77644), .B(n77638), .Z(n72309) );
  XOR U92470 ( .A(n77645), .B(n72309), .Z(n77838) );
  IV U92471 ( .A(n72310), .Z(n72311) );
  NOR U92472 ( .A(n72312), .B(n72311), .Z(n77839) );
  IV U92473 ( .A(n72313), .Z(n72315) );
  NOR U92474 ( .A(n72315), .B(n72314), .Z(n77841) );
  NOR U92475 ( .A(n77839), .B(n77841), .Z(n72316) );
  XOR U92476 ( .A(n77838), .B(n72316), .Z(n77636) );
  XOR U92477 ( .A(n77635), .B(n77636), .Z(n77626) );
  XOR U92478 ( .A(n77628), .B(n77626), .Z(n83691) );
  IV U92479 ( .A(n72317), .Z(n72319) );
  NOR U92480 ( .A(n72319), .B(n72318), .Z(n77629) );
  IV U92481 ( .A(n72320), .Z(n72322) );
  NOR U92482 ( .A(n72322), .B(n72321), .Z(n77630) );
  NOR U92483 ( .A(n77629), .B(n77630), .Z(n83692) );
  XOR U92484 ( .A(n83691), .B(n83692), .Z(n72323) );
  IV U92485 ( .A(n72323), .Z(n77618) );
  NOR U92486 ( .A(n72324), .B(n77618), .Z(n83697) );
  IV U92487 ( .A(n72325), .Z(n72326) );
  NOR U92488 ( .A(n72326), .B(n72328), .Z(n77620) );
  IV U92489 ( .A(n72327), .Z(n72329) );
  NOR U92490 ( .A(n72329), .B(n72328), .Z(n77617) );
  XOR U92491 ( .A(n77617), .B(n77618), .Z(n77621) );
  XOR U92492 ( .A(n77620), .B(n77621), .Z(n72334) );
  IV U92493 ( .A(n72334), .Z(n72330) );
  NOR U92494 ( .A(n72331), .B(n72330), .Z(n72332) );
  NOR U92495 ( .A(n83697), .B(n72332), .Z(n77614) );
  NOR U92496 ( .A(n72333), .B(n77614), .Z(n72336) );
  IV U92497 ( .A(n72333), .Z(n72335) );
  NOR U92498 ( .A(n72335), .B(n72334), .Z(n83700) );
  NOR U92499 ( .A(n72336), .B(n83700), .Z(n77609) );
  XOR U92500 ( .A(n72337), .B(n77609), .Z(n77604) );
  XOR U92501 ( .A(n77602), .B(n77604), .Z(n77606) );
  IV U92502 ( .A(n72338), .Z(n72339) );
  NOR U92503 ( .A(n72340), .B(n72339), .Z(n77600) );
  IV U92504 ( .A(n72341), .Z(n72342) );
  NOR U92505 ( .A(n72343), .B(n72342), .Z(n77605) );
  NOR U92506 ( .A(n77600), .B(n77605), .Z(n72344) );
  XOR U92507 ( .A(n77606), .B(n72344), .Z(n72345) );
  IV U92508 ( .A(n72345), .Z(n77599) );
  IV U92509 ( .A(n72346), .Z(n72347) );
  NOR U92510 ( .A(n72348), .B(n72347), .Z(n77597) );
  IV U92511 ( .A(n72349), .Z(n72351) );
  NOR U92512 ( .A(n72351), .B(n72350), .Z(n77595) );
  NOR U92513 ( .A(n77597), .B(n77595), .Z(n72352) );
  XOR U92514 ( .A(n77599), .B(n72352), .Z(n72353) );
  NOR U92515 ( .A(n72354), .B(n72353), .Z(n72357) );
  IV U92516 ( .A(n72354), .Z(n72356) );
  XOR U92517 ( .A(n77597), .B(n77599), .Z(n72355) );
  NOR U92518 ( .A(n72356), .B(n72355), .Z(n83711) );
  NOR U92519 ( .A(n72357), .B(n83711), .Z(n77852) );
  XOR U92520 ( .A(n77853), .B(n77852), .Z(n77593) );
  XOR U92521 ( .A(n77592), .B(n77593), .Z(n72368) );
  IV U92522 ( .A(n72368), .Z(n72366) );
  IV U92523 ( .A(n72358), .Z(n72359) );
  NOR U92524 ( .A(n72360), .B(n72359), .Z(n72370) );
  IV U92525 ( .A(n72361), .Z(n72362) );
  NOR U92526 ( .A(n72363), .B(n72362), .Z(n72367) );
  NOR U92527 ( .A(n72370), .B(n72367), .Z(n72364) );
  IV U92528 ( .A(n72364), .Z(n72365) );
  NOR U92529 ( .A(n72366), .B(n72365), .Z(n72373) );
  IV U92530 ( .A(n72367), .Z(n72369) );
  NOR U92531 ( .A(n72369), .B(n72368), .Z(n83446) );
  IV U92532 ( .A(n72370), .Z(n72371) );
  NOR U92533 ( .A(n72371), .B(n77593), .Z(n83452) );
  NOR U92534 ( .A(n83446), .B(n83452), .Z(n72372) );
  IV U92535 ( .A(n72372), .Z(n77591) );
  NOR U92536 ( .A(n72373), .B(n77591), .Z(n77585) );
  IV U92537 ( .A(n72374), .Z(n72376) );
  NOR U92538 ( .A(n72376), .B(n72375), .Z(n77588) );
  IV U92539 ( .A(n72377), .Z(n72379) );
  NOR U92540 ( .A(n72379), .B(n72378), .Z(n77584) );
  NOR U92541 ( .A(n77588), .B(n77584), .Z(n72380) );
  XOR U92542 ( .A(n77585), .B(n72380), .Z(n77859) );
  IV U92543 ( .A(n72381), .Z(n72383) );
  NOR U92544 ( .A(n72383), .B(n72382), .Z(n77582) );
  IV U92545 ( .A(n72384), .Z(n72385) );
  NOR U92546 ( .A(n72385), .B(n72388), .Z(n77857) );
  NOR U92547 ( .A(n77582), .B(n77857), .Z(n72386) );
  XOR U92548 ( .A(n77859), .B(n72386), .Z(n77861) );
  IV U92549 ( .A(n72387), .Z(n72389) );
  NOR U92550 ( .A(n72389), .B(n72388), .Z(n77860) );
  IV U92551 ( .A(n72390), .Z(n72393) );
  NOR U92552 ( .A(n72391), .B(n72399), .Z(n72392) );
  IV U92553 ( .A(n72392), .Z(n72396) );
  NOR U92554 ( .A(n72393), .B(n72396), .Z(n77864) );
  NOR U92555 ( .A(n77860), .B(n77864), .Z(n72394) );
  XOR U92556 ( .A(n77861), .B(n72394), .Z(n77872) );
  IV U92557 ( .A(n72395), .Z(n72397) );
  NOR U92558 ( .A(n72397), .B(n72396), .Z(n77580) );
  IV U92559 ( .A(n72398), .Z(n72400) );
  NOR U92560 ( .A(n72400), .B(n72399), .Z(n77870) );
  NOR U92561 ( .A(n77580), .B(n77870), .Z(n72401) );
  XOR U92562 ( .A(n77872), .B(n72401), .Z(n77868) );
  IV U92563 ( .A(n72402), .Z(n72404) );
  NOR U92564 ( .A(n72404), .B(n72403), .Z(n83427) );
  IV U92565 ( .A(n72405), .Z(n72407) );
  NOR U92566 ( .A(n72407), .B(n72406), .Z(n83431) );
  NOR U92567 ( .A(n83427), .B(n83431), .Z(n77869) );
  XOR U92568 ( .A(n77868), .B(n77869), .Z(n77575) );
  XOR U92569 ( .A(n77574), .B(n77575), .Z(n77578) );
  NOR U92570 ( .A(n72414), .B(n77578), .Z(n83413) );
  IV U92571 ( .A(n72408), .Z(n72410) );
  NOR U92572 ( .A(n72410), .B(n72409), .Z(n77571) );
  IV U92573 ( .A(n72411), .Z(n72412) );
  NOR U92574 ( .A(n72413), .B(n72412), .Z(n77577) );
  XOR U92575 ( .A(n77577), .B(n77578), .Z(n77572) );
  IV U92576 ( .A(n77572), .Z(n72415) );
  XOR U92577 ( .A(n77571), .B(n72415), .Z(n72417) );
  NOR U92578 ( .A(n72415), .B(n72414), .Z(n72416) );
  NOR U92579 ( .A(n72417), .B(n72416), .Z(n72418) );
  NOR U92580 ( .A(n83413), .B(n72418), .Z(n77561) );
  NOR U92581 ( .A(n72419), .B(n77565), .Z(n72423) );
  IV U92582 ( .A(n72420), .Z(n72421) );
  NOR U92583 ( .A(n72422), .B(n72421), .Z(n77560) );
  NOR U92584 ( .A(n72423), .B(n77560), .Z(n72424) );
  XOR U92585 ( .A(n77561), .B(n72424), .Z(n77559) );
  IV U92586 ( .A(n72425), .Z(n72426) );
  NOR U92587 ( .A(n72427), .B(n72426), .Z(n77557) );
  IV U92588 ( .A(n72428), .Z(n72430) );
  NOR U92589 ( .A(n72430), .B(n72429), .Z(n77555) );
  NOR U92590 ( .A(n77557), .B(n77555), .Z(n72431) );
  XOR U92591 ( .A(n77559), .B(n72431), .Z(n77552) );
  IV U92592 ( .A(n72432), .Z(n72433) );
  NOR U92593 ( .A(n72433), .B(n72439), .Z(n72434) );
  IV U92594 ( .A(n72434), .Z(n77553) );
  XOR U92595 ( .A(n77552), .B(n77553), .Z(n83395) );
  IV U92596 ( .A(n72435), .Z(n72436) );
  NOR U92597 ( .A(n72437), .B(n72436), .Z(n83394) );
  IV U92598 ( .A(n72438), .Z(n72440) );
  NOR U92599 ( .A(n72440), .B(n72439), .Z(n83401) );
  NOR U92600 ( .A(n83394), .B(n83401), .Z(n77878) );
  XOR U92601 ( .A(n83395), .B(n77878), .Z(n77879) );
  XOR U92602 ( .A(n77880), .B(n77879), .Z(n77887) );
  IV U92603 ( .A(n72441), .Z(n72442) );
  NOR U92604 ( .A(n72443), .B(n72442), .Z(n77884) );
  XOR U92605 ( .A(n77887), .B(n77884), .Z(n77894) );
  IV U92606 ( .A(n72444), .Z(n77888) );
  NOR U92607 ( .A(n77888), .B(n72445), .Z(n72448) );
  IV U92608 ( .A(n72446), .Z(n72447) );
  NOR U92609 ( .A(n72447), .B(n72454), .Z(n77892) );
  NOR U92610 ( .A(n72448), .B(n77892), .Z(n72449) );
  XOR U92611 ( .A(n77894), .B(n72449), .Z(n77549) );
  IV U92612 ( .A(n72450), .Z(n72459) );
  IV U92613 ( .A(n72451), .Z(n72452) );
  NOR U92614 ( .A(n72459), .B(n72452), .Z(n77550) );
  IV U92615 ( .A(n72453), .Z(n72455) );
  NOR U92616 ( .A(n72455), .B(n72454), .Z(n77900) );
  NOR U92617 ( .A(n77550), .B(n77900), .Z(n72456) );
  XOR U92618 ( .A(n77549), .B(n72456), .Z(n77546) );
  IV U92619 ( .A(n72457), .Z(n72458) );
  NOR U92620 ( .A(n72459), .B(n72458), .Z(n77544) );
  XOR U92621 ( .A(n77546), .B(n77544), .Z(n77906) );
  XOR U92622 ( .A(n77547), .B(n77906), .Z(n77920) );
  NOR U92623 ( .A(n72460), .B(n77907), .Z(n72466) );
  IV U92624 ( .A(n72461), .Z(n72465) );
  IV U92625 ( .A(n72462), .Z(n72470) );
  NOR U92626 ( .A(n72463), .B(n72470), .Z(n72464) );
  IV U92627 ( .A(n72464), .Z(n72472) );
  NOR U92628 ( .A(n72465), .B(n72472), .Z(n77919) );
  NOR U92629 ( .A(n72466), .B(n77919), .Z(n72467) );
  XOR U92630 ( .A(n77920), .B(n72467), .Z(n77541) );
  IV U92631 ( .A(n72468), .Z(n72469) );
  NOR U92632 ( .A(n72470), .B(n72469), .Z(n77542) );
  IV U92633 ( .A(n72471), .Z(n72473) );
  NOR U92634 ( .A(n72473), .B(n72472), .Z(n77916) );
  NOR U92635 ( .A(n77542), .B(n77916), .Z(n72474) );
  XOR U92636 ( .A(n77541), .B(n72474), .Z(n89106) );
  IV U92637 ( .A(n72475), .Z(n72476) );
  NOR U92638 ( .A(n72477), .B(n72476), .Z(n89111) );
  IV U92639 ( .A(n72478), .Z(n72480) );
  NOR U92640 ( .A(n72480), .B(n72479), .Z(n89101) );
  NOR U92641 ( .A(n89111), .B(n89101), .Z(n77924) );
  XOR U92642 ( .A(n89106), .B(n77924), .Z(n77538) );
  XOR U92643 ( .A(n77540), .B(n77538), .Z(n77939) );
  XOR U92644 ( .A(n77935), .B(n77939), .Z(n72481) );
  IV U92645 ( .A(n72481), .Z(n77931) );
  XOR U92646 ( .A(n72482), .B(n77931), .Z(n72493) );
  IV U92647 ( .A(n72493), .Z(n72491) );
  IV U92648 ( .A(n72483), .Z(n72484) );
  NOR U92649 ( .A(n72485), .B(n72484), .Z(n72495) );
  IV U92650 ( .A(n72486), .Z(n72488) );
  NOR U92651 ( .A(n72488), .B(n72487), .Z(n72492) );
  NOR U92652 ( .A(n72495), .B(n72492), .Z(n72489) );
  IV U92653 ( .A(n72489), .Z(n72490) );
  NOR U92654 ( .A(n72491), .B(n72490), .Z(n72498) );
  IV U92655 ( .A(n72492), .Z(n72494) );
  NOR U92656 ( .A(n72494), .B(n72493), .Z(n83349) );
  IV U92657 ( .A(n72495), .Z(n72496) );
  NOR U92658 ( .A(n72496), .B(n77931), .Z(n83352) );
  NOR U92659 ( .A(n83349), .B(n83352), .Z(n72497) );
  IV U92660 ( .A(n72497), .Z(n77959) );
  NOR U92661 ( .A(n72498), .B(n77959), .Z(n77956) );
  XOR U92662 ( .A(n72499), .B(n77956), .Z(n77964) );
  XOR U92663 ( .A(n77962), .B(n77964), .Z(n77972) );
  XOR U92664 ( .A(n77969), .B(n77972), .Z(n77537) );
  NOR U92665 ( .A(n72500), .B(n77973), .Z(n72504) );
  IV U92666 ( .A(n72501), .Z(n72503) );
  IV U92667 ( .A(n72502), .Z(n72508) );
  NOR U92668 ( .A(n72503), .B(n72508), .Z(n77535) );
  NOR U92669 ( .A(n72504), .B(n77535), .Z(n72505) );
  XOR U92670 ( .A(n77537), .B(n72505), .Z(n77980) );
  IV U92671 ( .A(n72506), .Z(n72507) );
  NOR U92672 ( .A(n72508), .B(n72507), .Z(n72509) );
  IV U92673 ( .A(n72509), .Z(n77981) );
  XOR U92674 ( .A(n77980), .B(n77981), .Z(n77992) );
  XOR U92675 ( .A(n77532), .B(n77992), .Z(n77985) );
  IV U92676 ( .A(n72510), .Z(n72512) );
  NOR U92677 ( .A(n72512), .B(n72511), .Z(n77991) );
  IV U92678 ( .A(n72513), .Z(n72514) );
  NOR U92679 ( .A(n72515), .B(n72514), .Z(n77983) );
  NOR U92680 ( .A(n77991), .B(n77983), .Z(n72516) );
  XOR U92681 ( .A(n77985), .B(n72516), .Z(n72517) );
  IV U92682 ( .A(n72517), .Z(n77997) );
  XOR U92683 ( .A(n77995), .B(n77997), .Z(n77529) );
  IV U92684 ( .A(n72518), .Z(n77524) );
  NOR U92685 ( .A(n72519), .B(n77524), .Z(n72523) );
  IV U92686 ( .A(n72520), .Z(n72522) );
  NOR U92687 ( .A(n72522), .B(n72521), .Z(n77528) );
  NOR U92688 ( .A(n72523), .B(n77528), .Z(n72524) );
  XOR U92689 ( .A(n77529), .B(n72524), .Z(n78003) );
  XOR U92690 ( .A(n78004), .B(n78003), .Z(n78007) );
  XOR U92691 ( .A(n78006), .B(n78007), .Z(n78018) );
  XOR U92692 ( .A(n72525), .B(n78018), .Z(n78019) );
  XOR U92693 ( .A(n78020), .B(n78019), .Z(n78027) );
  XOR U92694 ( .A(n78022), .B(n78027), .Z(n77508) );
  IV U92695 ( .A(n72526), .Z(n72527) );
  NOR U92696 ( .A(n72528), .B(n72527), .Z(n72531) );
  NOR U92697 ( .A(n72529), .B(n77509), .Z(n72530) );
  NOR U92698 ( .A(n72531), .B(n72530), .Z(n72532) );
  XOR U92699 ( .A(n77508), .B(n72532), .Z(n77501) );
  XOR U92700 ( .A(n77502), .B(n77501), .Z(n77504) );
  IV U92701 ( .A(n77504), .Z(n72540) );
  IV U92702 ( .A(n72533), .Z(n72534) );
  NOR U92703 ( .A(n72535), .B(n72534), .Z(n77503) );
  IV U92704 ( .A(n72536), .Z(n72538) );
  NOR U92705 ( .A(n72538), .B(n72537), .Z(n77496) );
  NOR U92706 ( .A(n77503), .B(n77496), .Z(n72539) );
  XOR U92707 ( .A(n72540), .B(n72539), .Z(n77500) );
  XOR U92708 ( .A(n77498), .B(n77500), .Z(n77494) );
  XOR U92709 ( .A(n72541), .B(n77494), .Z(n72542) );
  IV U92710 ( .A(n72542), .Z(n77490) );
  XOR U92711 ( .A(n77488), .B(n77490), .Z(n78041) );
  IV U92712 ( .A(n72543), .Z(n72545) );
  NOR U92713 ( .A(n72545), .B(n72544), .Z(n78039) );
  XOR U92714 ( .A(n78041), .B(n78039), .Z(n78043) );
  XOR U92715 ( .A(n78042), .B(n78043), .Z(n78048) );
  IV U92716 ( .A(n78048), .Z(n72550) );
  XOR U92717 ( .A(n78047), .B(n72550), .Z(n72552) );
  IV U92718 ( .A(n72546), .Z(n72547) );
  NOR U92719 ( .A(n72548), .B(n72547), .Z(n72549) );
  IV U92720 ( .A(n72549), .Z(n72555) );
  NOR U92721 ( .A(n72550), .B(n72555), .Z(n72551) );
  NOR U92722 ( .A(n72552), .B(n72551), .Z(n72556) );
  NOR U92723 ( .A(n72557), .B(n72556), .Z(n78046) );
  IV U92724 ( .A(n72553), .Z(n72554) );
  NOR U92725 ( .A(n72554), .B(n72565), .Z(n77481) );
  NOR U92726 ( .A(n72555), .B(n78048), .Z(n83287) );
  NOR U92727 ( .A(n83287), .B(n72556), .Z(n77482) );
  XOR U92728 ( .A(n77481), .B(n77482), .Z(n72559) );
  NOR U92729 ( .A(n77482), .B(n72557), .Z(n72558) );
  NOR U92730 ( .A(n72559), .B(n72558), .Z(n72560) );
  NOR U92731 ( .A(n78046), .B(n72560), .Z(n77476) );
  IV U92732 ( .A(n72561), .Z(n72562) );
  NOR U92733 ( .A(n72563), .B(n72562), .Z(n77475) );
  IV U92734 ( .A(n72564), .Z(n72566) );
  NOR U92735 ( .A(n72566), .B(n72565), .Z(n77485) );
  NOR U92736 ( .A(n77475), .B(n77485), .Z(n72567) );
  XOR U92737 ( .A(n77476), .B(n72567), .Z(n77480) );
  XOR U92738 ( .A(n72568), .B(n77480), .Z(n77467) );
  XOR U92739 ( .A(n77468), .B(n77467), .Z(n77471) );
  XOR U92740 ( .A(n77470), .B(n77471), .Z(n83870) );
  XOR U92741 ( .A(n77465), .B(n83870), .Z(n72569) );
  IV U92742 ( .A(n72569), .Z(n78060) );
  XOR U92743 ( .A(n78057), .B(n78060), .Z(n78067) );
  XOR U92744 ( .A(n72570), .B(n78067), .Z(n77461) );
  XOR U92745 ( .A(n72571), .B(n77461), .Z(n72582) );
  IV U92746 ( .A(n72582), .Z(n72572) );
  NOR U92747 ( .A(n72575), .B(n72572), .Z(n72573) );
  IV U92748 ( .A(n72573), .Z(n72589) );
  NOR U92749 ( .A(n72574), .B(n72589), .Z(n83894) );
  NOR U92750 ( .A(n72576), .B(n72575), .Z(n72585) );
  IV U92751 ( .A(n72577), .Z(n72578) );
  NOR U92752 ( .A(n72579), .B(n72578), .Z(n72583) );
  IV U92753 ( .A(n72583), .Z(n72581) );
  XOR U92754 ( .A(n77461), .B(n77459), .Z(n72580) );
  NOR U92755 ( .A(n72581), .B(n72580), .Z(n83257) );
  NOR U92756 ( .A(n72583), .B(n72582), .Z(n72584) );
  NOR U92757 ( .A(n83257), .B(n72584), .Z(n72592) );
  NOR U92758 ( .A(n72585), .B(n72592), .Z(n72586) );
  NOR U92759 ( .A(n83894), .B(n72586), .Z(n72587) );
  NOR U92760 ( .A(n72591), .B(n72587), .Z(n72597) );
  IV U92761 ( .A(n72588), .Z(n72590) );
  NOR U92762 ( .A(n72590), .B(n72589), .Z(n83897) );
  IV U92763 ( .A(n72591), .Z(n72594) );
  IV U92764 ( .A(n72592), .Z(n72593) );
  NOR U92765 ( .A(n72594), .B(n72593), .Z(n83901) );
  NOR U92766 ( .A(n83897), .B(n83901), .Z(n72595) );
  IV U92767 ( .A(n72595), .Z(n72596) );
  NOR U92768 ( .A(n72597), .B(n72596), .Z(n72598) );
  IV U92769 ( .A(n72598), .Z(n78076) );
  IV U92770 ( .A(n72599), .Z(n72600) );
  NOR U92771 ( .A(n72600), .B(n72608), .Z(n78074) );
  XOR U92772 ( .A(n78076), .B(n78074), .Z(n83248) );
  IV U92773 ( .A(n72601), .Z(n72606) );
  IV U92774 ( .A(n72602), .Z(n72603) );
  NOR U92775 ( .A(n72606), .B(n72603), .Z(n78084) );
  IV U92776 ( .A(n72604), .Z(n72605) );
  NOR U92777 ( .A(n72606), .B(n72605), .Z(n83247) );
  IV U92778 ( .A(n72607), .Z(n72609) );
  NOR U92779 ( .A(n72609), .B(n72608), .Z(n83252) );
  NOR U92780 ( .A(n83247), .B(n83252), .Z(n77456) );
  IV U92781 ( .A(n77456), .Z(n72610) );
  NOR U92782 ( .A(n78084), .B(n72610), .Z(n72611) );
  XOR U92783 ( .A(n83248), .B(n72611), .Z(n77454) );
  IV U92784 ( .A(n72612), .Z(n72614) );
  NOR U92785 ( .A(n72614), .B(n72613), .Z(n78080) );
  IV U92786 ( .A(n72615), .Z(n72616) );
  NOR U92787 ( .A(n72617), .B(n72616), .Z(n77453) );
  NOR U92788 ( .A(n78080), .B(n77453), .Z(n72618) );
  XOR U92789 ( .A(n77454), .B(n72618), .Z(n83236) );
  XOR U92790 ( .A(n72619), .B(n83236), .Z(n77450) );
  XOR U92791 ( .A(n77449), .B(n77450), .Z(n78095) );
  XOR U92792 ( .A(n77446), .B(n78095), .Z(n77444) );
  IV U92793 ( .A(n72620), .Z(n72622) );
  NOR U92794 ( .A(n72622), .B(n72621), .Z(n78094) );
  IV U92795 ( .A(n72623), .Z(n72625) );
  NOR U92796 ( .A(n72625), .B(n72624), .Z(n77443) );
  NOR U92797 ( .A(n78094), .B(n77443), .Z(n72626) );
  XOR U92798 ( .A(n77444), .B(n72626), .Z(n72627) );
  IV U92799 ( .A(n72627), .Z(n78109) );
  XOR U92800 ( .A(n77441), .B(n78109), .Z(n72628) );
  NOR U92801 ( .A(n72629), .B(n72628), .Z(n83228) );
  IV U92802 ( .A(n72630), .Z(n72631) );
  NOR U92803 ( .A(n72632), .B(n72631), .Z(n78107) );
  NOR U92804 ( .A(n77441), .B(n78107), .Z(n72633) );
  XOR U92805 ( .A(n78109), .B(n72633), .Z(n72634) );
  NOR U92806 ( .A(n72635), .B(n72634), .Z(n72636) );
  NOR U92807 ( .A(n83228), .B(n72636), .Z(n78105) );
  XOR U92808 ( .A(n78106), .B(n78105), .Z(n78117) );
  IV U92809 ( .A(n72637), .Z(n72639) );
  NOR U92810 ( .A(n72639), .B(n72638), .Z(n72640) );
  IV U92811 ( .A(n72640), .Z(n77440) );
  XOR U92812 ( .A(n78117), .B(n77440), .Z(n72641) );
  XOR U92813 ( .A(n72642), .B(n72641), .Z(n78121) );
  XOR U92814 ( .A(n78119), .B(n78121), .Z(n83216) );
  XOR U92815 ( .A(n78122), .B(n83216), .Z(n78126) );
  NOR U92816 ( .A(n78129), .B(n78127), .Z(n72646) );
  IV U92817 ( .A(n72643), .Z(n72645) );
  NOR U92818 ( .A(n72645), .B(n72644), .Z(n78131) );
  NOR U92819 ( .A(n72646), .B(n78131), .Z(n72647) );
  XOR U92820 ( .A(n78126), .B(n72647), .Z(n77436) );
  XOR U92821 ( .A(n77434), .B(n77436), .Z(n77438) );
  XOR U92822 ( .A(n72648), .B(n77438), .Z(n77430) );
  IV U92823 ( .A(n72649), .Z(n72652) );
  IV U92824 ( .A(n72650), .Z(n72651) );
  NOR U92825 ( .A(n72652), .B(n72651), .Z(n78136) );
  IV U92826 ( .A(n72653), .Z(n72654) );
  NOR U92827 ( .A(n72654), .B(n72657), .Z(n77429) );
  NOR U92828 ( .A(n78136), .B(n77429), .Z(n72655) );
  XOR U92829 ( .A(n77430), .B(n72655), .Z(n78141) );
  IV U92830 ( .A(n72656), .Z(n72658) );
  NOR U92831 ( .A(n72658), .B(n72657), .Z(n78139) );
  XOR U92832 ( .A(n78141), .B(n78139), .Z(n78148) );
  XOR U92833 ( .A(n72659), .B(n78148), .Z(n77424) );
  IV U92834 ( .A(n72660), .Z(n72662) );
  NOR U92835 ( .A(n72662), .B(n72661), .Z(n77423) );
  IV U92836 ( .A(n72663), .Z(n72665) );
  NOR U92837 ( .A(n72665), .B(n72664), .Z(n78152) );
  NOR U92838 ( .A(n77423), .B(n78152), .Z(n72666) );
  XOR U92839 ( .A(n77424), .B(n72666), .Z(n78163) );
  XOR U92840 ( .A(n72667), .B(n78163), .Z(n72668) );
  IV U92841 ( .A(n72668), .Z(n78161) );
  XOR U92842 ( .A(n78159), .B(n78161), .Z(n83966) );
  IV U92843 ( .A(n72672), .Z(n77419) );
  NOR U92844 ( .A(n77419), .B(n77417), .Z(n72676) );
  IV U92845 ( .A(n72669), .Z(n72670) );
  NOR U92846 ( .A(n72670), .B(n77417), .Z(n83964) );
  IV U92847 ( .A(n72671), .Z(n72674) );
  XOR U92848 ( .A(n72672), .B(n77417), .Z(n72673) );
  NOR U92849 ( .A(n72674), .B(n72673), .Z(n83970) );
  NOR U92850 ( .A(n83964), .B(n83970), .Z(n78176) );
  IV U92851 ( .A(n78176), .Z(n72675) );
  NOR U92852 ( .A(n72676), .B(n72675), .Z(n72677) );
  XOR U92853 ( .A(n83966), .B(n72677), .Z(n72678) );
  IV U92854 ( .A(n72678), .Z(n78175) );
  IV U92855 ( .A(n72679), .Z(n72682) );
  IV U92856 ( .A(n72680), .Z(n72681) );
  NOR U92857 ( .A(n72682), .B(n72681), .Z(n78173) );
  XOR U92858 ( .A(n78175), .B(n78173), .Z(n77410) );
  XOR U92859 ( .A(n77409), .B(n77410), .Z(n77414) );
  XOR U92860 ( .A(n77412), .B(n77414), .Z(n78182) );
  XOR U92861 ( .A(n72683), .B(n78182), .Z(n78185) );
  IV U92862 ( .A(n72684), .Z(n78190) );
  NOR U92863 ( .A(n78190), .B(n72685), .Z(n72689) );
  IV U92864 ( .A(n72686), .Z(n72688) );
  NOR U92865 ( .A(n72688), .B(n72687), .Z(n78184) );
  NOR U92866 ( .A(n72689), .B(n78184), .Z(n72690) );
  XOR U92867 ( .A(n78185), .B(n72690), .Z(n78198) );
  XOR U92868 ( .A(n78196), .B(n78198), .Z(n78200) );
  XOR U92869 ( .A(n78199), .B(n78200), .Z(n77407) );
  NOR U92870 ( .A(n72691), .B(n77407), .Z(n83148) );
  IV U92871 ( .A(n72692), .Z(n72693) );
  NOR U92872 ( .A(n72694), .B(n72693), .Z(n77406) );
  XOR U92873 ( .A(n77406), .B(n77407), .Z(n72709) );
  IV U92874 ( .A(n72709), .Z(n72701) );
  IV U92875 ( .A(n72695), .Z(n72696) );
  NOR U92876 ( .A(n72697), .B(n72696), .Z(n72708) );
  NOR U92877 ( .A(n72698), .B(n72708), .Z(n72699) );
  IV U92878 ( .A(n72699), .Z(n72700) );
  NOR U92879 ( .A(n72701), .B(n72700), .Z(n72702) );
  NOR U92880 ( .A(n83148), .B(n72702), .Z(n72703) );
  IV U92881 ( .A(n72703), .Z(n72711) );
  IV U92882 ( .A(n72704), .Z(n72706) );
  NOR U92883 ( .A(n72706), .B(n72705), .Z(n72713) );
  IV U92884 ( .A(n72713), .Z(n72707) );
  NOR U92885 ( .A(n72711), .B(n72707), .Z(n83975) );
  IV U92886 ( .A(n72708), .Z(n72710) );
  NOR U92887 ( .A(n72710), .B(n72709), .Z(n83977) );
  NOR U92888 ( .A(n83977), .B(n72711), .Z(n72712) );
  NOR U92889 ( .A(n72713), .B(n72712), .Z(n72714) );
  NOR U92890 ( .A(n83975), .B(n72714), .Z(n72715) );
  IV U92891 ( .A(n72715), .Z(n77402) );
  XOR U92892 ( .A(n77401), .B(n77402), .Z(n77399) );
  XOR U92893 ( .A(n77398), .B(n77399), .Z(n77395) );
  XOR U92894 ( .A(n77394), .B(n77395), .Z(n77388) );
  IV U92895 ( .A(n72716), .Z(n72718) );
  NOR U92896 ( .A(n72718), .B(n72717), .Z(n77386) );
  XOR U92897 ( .A(n77388), .B(n77386), .Z(n77390) );
  XOR U92898 ( .A(n77389), .B(n77390), .Z(n83998) );
  XOR U92899 ( .A(n77381), .B(n83998), .Z(n72719) );
  IV U92900 ( .A(n72719), .Z(n77384) );
  XOR U92901 ( .A(n77382), .B(n77384), .Z(n77371) );
  NOR U92902 ( .A(n72725), .B(n77371), .Z(n84017) );
  IV U92903 ( .A(n72720), .Z(n72722) );
  NOR U92904 ( .A(n72722), .B(n72721), .Z(n77365) );
  IV U92905 ( .A(n72723), .Z(n77380) );
  NOR U92906 ( .A(n77380), .B(n72724), .Z(n77370) );
  XOR U92907 ( .A(n77370), .B(n77371), .Z(n77366) );
  IV U92908 ( .A(n77366), .Z(n72726) );
  XOR U92909 ( .A(n77365), .B(n72726), .Z(n72728) );
  NOR U92910 ( .A(n72726), .B(n72725), .Z(n72727) );
  NOR U92911 ( .A(n72728), .B(n72727), .Z(n72729) );
  NOR U92912 ( .A(n84017), .B(n72729), .Z(n78208) );
  XOR U92913 ( .A(n72730), .B(n78208), .Z(n78218) );
  XOR U92914 ( .A(n78216), .B(n78218), .Z(n77361) );
  IV U92915 ( .A(n72731), .Z(n72732) );
  NOR U92916 ( .A(n72733), .B(n72732), .Z(n77363) );
  IV U92917 ( .A(n72734), .Z(n72736) );
  NOR U92918 ( .A(n72736), .B(n72735), .Z(n77360) );
  NOR U92919 ( .A(n77363), .B(n77360), .Z(n72737) );
  XOR U92920 ( .A(n77361), .B(n72737), .Z(n72738) );
  IV U92921 ( .A(n72738), .Z(n77358) );
  IV U92922 ( .A(n72739), .Z(n72740) );
  NOR U92923 ( .A(n72741), .B(n72740), .Z(n77356) );
  IV U92924 ( .A(n72742), .Z(n72743) );
  NOR U92925 ( .A(n72744), .B(n72743), .Z(n77354) );
  NOR U92926 ( .A(n77356), .B(n77354), .Z(n72745) );
  XOR U92927 ( .A(n77358), .B(n72745), .Z(n72746) );
  NOR U92928 ( .A(n72747), .B(n72746), .Z(n72750) );
  IV U92929 ( .A(n72747), .Z(n72749) );
  XOR U92930 ( .A(n77356), .B(n77358), .Z(n72748) );
  NOR U92931 ( .A(n72749), .B(n72748), .Z(n84051) );
  NOR U92932 ( .A(n72750), .B(n84051), .Z(n72751) );
  IV U92933 ( .A(n72751), .Z(n77352) );
  XOR U92934 ( .A(n77351), .B(n77352), .Z(n77349) );
  IV U92935 ( .A(n72752), .Z(n72754) );
  NOR U92936 ( .A(n72754), .B(n72753), .Z(n77348) );
  IV U92937 ( .A(n72755), .Z(n72757) );
  NOR U92938 ( .A(n72757), .B(n72756), .Z(n77346) );
  NOR U92939 ( .A(n77348), .B(n77346), .Z(n72758) );
  XOR U92940 ( .A(n77349), .B(n72758), .Z(n77344) );
  XOR U92941 ( .A(n72759), .B(n77344), .Z(n77339) );
  IV U92942 ( .A(n72760), .Z(n72761) );
  NOR U92943 ( .A(n72762), .B(n72761), .Z(n77337) );
  XOR U92944 ( .A(n77339), .B(n77337), .Z(n77342) );
  IV U92945 ( .A(n72763), .Z(n72764) );
  NOR U92946 ( .A(n72765), .B(n72764), .Z(n77340) );
  XOR U92947 ( .A(n77342), .B(n77340), .Z(n77332) );
  IV U92948 ( .A(n72766), .Z(n72768) );
  NOR U92949 ( .A(n72768), .B(n72767), .Z(n72776) );
  IV U92950 ( .A(n72776), .Z(n72769) );
  NOR U92951 ( .A(n77332), .B(n72769), .Z(n84075) );
  IV U92952 ( .A(n72770), .Z(n72771) );
  NOR U92953 ( .A(n72774), .B(n72771), .Z(n77331) );
  XOR U92954 ( .A(n77331), .B(n77332), .Z(n77336) );
  IV U92955 ( .A(n72772), .Z(n72773) );
  NOR U92956 ( .A(n72774), .B(n72773), .Z(n77334) );
  XOR U92957 ( .A(n77336), .B(n77334), .Z(n72780) );
  IV U92958 ( .A(n72780), .Z(n72775) );
  NOR U92959 ( .A(n72776), .B(n72775), .Z(n72777) );
  NOR U92960 ( .A(n84075), .B(n72777), .Z(n72778) );
  NOR U92961 ( .A(n72779), .B(n72778), .Z(n72782) );
  IV U92962 ( .A(n72779), .Z(n72781) );
  NOR U92963 ( .A(n72781), .B(n72780), .Z(n77330) );
  NOR U92964 ( .A(n72782), .B(n77330), .Z(n77327) );
  IV U92965 ( .A(n72783), .Z(n72785) );
  NOR U92966 ( .A(n72785), .B(n72784), .Z(n72786) );
  IV U92967 ( .A(n72786), .Z(n77328) );
  XOR U92968 ( .A(n77327), .B(n77328), .Z(n78251) );
  NOR U92969 ( .A(n78246), .B(n72787), .Z(n72790) );
  NOR U92970 ( .A(n72789), .B(n72788), .Z(n78250) );
  NOR U92971 ( .A(n72790), .B(n78250), .Z(n72791) );
  IV U92972 ( .A(n72791), .Z(n72792) );
  NOR U92973 ( .A(n77325), .B(n72792), .Z(n72793) );
  XOR U92974 ( .A(n78251), .B(n72793), .Z(n72794) );
  IV U92975 ( .A(n72794), .Z(n77324) );
  XOR U92976 ( .A(n77322), .B(n77324), .Z(n77318) );
  XOR U92977 ( .A(n77316), .B(n77318), .Z(n77321) );
  XOR U92978 ( .A(n77319), .B(n77321), .Z(n78263) );
  XOR U92979 ( .A(n72795), .B(n78263), .Z(n72805) );
  IV U92980 ( .A(n72796), .Z(n72798) );
  NOR U92981 ( .A(n72798), .B(n72797), .Z(n72808) );
  IV U92982 ( .A(n72799), .Z(n72801) );
  NOR U92983 ( .A(n72801), .B(n72800), .Z(n72804) );
  NOR U92984 ( .A(n72808), .B(n72804), .Z(n72802) );
  IV U92985 ( .A(n72802), .Z(n72803) );
  NOR U92986 ( .A(n72805), .B(n72803), .Z(n72812) );
  IV U92987 ( .A(n72804), .Z(n72807) );
  IV U92988 ( .A(n72805), .Z(n72806) );
  NOR U92989 ( .A(n72807), .B(n72806), .Z(n83102) );
  IV U92990 ( .A(n72808), .Z(n72810) );
  XOR U92991 ( .A(n78261), .B(n78263), .Z(n72809) );
  NOR U92992 ( .A(n72810), .B(n72809), .Z(n84100) );
  NOR U92993 ( .A(n83102), .B(n84100), .Z(n72811) );
  IV U92994 ( .A(n72811), .Z(n78276) );
  NOR U92995 ( .A(n72812), .B(n78276), .Z(n78272) );
  NOR U92996 ( .A(n84108), .B(n78273), .Z(n72816) );
  IV U92997 ( .A(n72813), .Z(n72814) );
  NOR U92998 ( .A(n72815), .B(n72814), .Z(n78286) );
  NOR U92999 ( .A(n72816), .B(n78286), .Z(n72817) );
  XOR U93000 ( .A(n78272), .B(n72817), .Z(n78285) );
  XOR U93001 ( .A(n78283), .B(n78285), .Z(n78292) );
  IV U93002 ( .A(n72818), .Z(n72820) );
  NOR U93003 ( .A(n72820), .B(n72819), .Z(n78290) );
  XOR U93004 ( .A(n78292), .B(n78290), .Z(n78297) );
  IV U93005 ( .A(n72821), .Z(n72822) );
  NOR U93006 ( .A(n72823), .B(n72822), .Z(n78293) );
  IV U93007 ( .A(n72824), .Z(n72825) );
  NOR U93008 ( .A(n72834), .B(n72825), .Z(n78296) );
  NOR U93009 ( .A(n78293), .B(n78296), .Z(n72826) );
  XOR U93010 ( .A(n78297), .B(n72826), .Z(n77308) );
  IV U93011 ( .A(n72827), .Z(n72828) );
  NOR U93012 ( .A(n72829), .B(n72828), .Z(n78300) );
  IV U93013 ( .A(n72830), .Z(n72831) );
  NOR U93014 ( .A(n72832), .B(n72831), .Z(n77310) );
  IV U93015 ( .A(n72833), .Z(n72835) );
  NOR U93016 ( .A(n72835), .B(n72834), .Z(n77311) );
  XOR U93017 ( .A(n77310), .B(n77311), .Z(n72836) );
  NOR U93018 ( .A(n78300), .B(n72836), .Z(n72837) );
  XOR U93019 ( .A(n77308), .B(n72837), .Z(n78305) );
  IV U93020 ( .A(n72838), .Z(n72839) );
  NOR U93021 ( .A(n72839), .B(n72846), .Z(n78303) );
  XOR U93022 ( .A(n78305), .B(n78303), .Z(n78309) );
  IV U93023 ( .A(n72840), .Z(n72841) );
  NOR U93024 ( .A(n72841), .B(n72846), .Z(n78307) );
  XOR U93025 ( .A(n78309), .B(n78307), .Z(n78311) );
  XOR U93026 ( .A(n78310), .B(n78311), .Z(n78316) );
  IV U93027 ( .A(n72842), .Z(n72843) );
  NOR U93028 ( .A(n72844), .B(n72843), .Z(n78315) );
  IV U93029 ( .A(n72845), .Z(n72847) );
  NOR U93030 ( .A(n72847), .B(n72846), .Z(n77306) );
  NOR U93031 ( .A(n78315), .B(n77306), .Z(n72848) );
  XOR U93032 ( .A(n78316), .B(n72848), .Z(n72849) );
  IV U93033 ( .A(n72849), .Z(n78319) );
  XOR U93034 ( .A(n78318), .B(n78319), .Z(n77302) );
  XOR U93035 ( .A(n77300), .B(n77302), .Z(n77305) );
  IV U93036 ( .A(n72850), .Z(n72851) );
  NOR U93037 ( .A(n72852), .B(n72851), .Z(n77303) );
  XOR U93038 ( .A(n77305), .B(n77303), .Z(n77294) );
  XOR U93039 ( .A(n77293), .B(n77294), .Z(n77289) );
  IV U93040 ( .A(n77289), .Z(n72853) );
  NOR U93041 ( .A(n72854), .B(n72853), .Z(n72859) );
  NOR U93042 ( .A(n72855), .B(n77305), .Z(n72856) );
  IV U93043 ( .A(n72856), .Z(n77297) );
  NOR U93044 ( .A(n77297), .B(n72857), .Z(n72858) );
  NOR U93045 ( .A(n72859), .B(n72858), .Z(n77285) );
  IV U93046 ( .A(n72860), .Z(n72862) );
  NOR U93047 ( .A(n72862), .B(n72861), .Z(n77288) );
  IV U93048 ( .A(n72863), .Z(n72864) );
  NOR U93049 ( .A(n72865), .B(n72864), .Z(n77284) );
  NOR U93050 ( .A(n77288), .B(n77284), .Z(n72866) );
  XOR U93051 ( .A(n77285), .B(n72866), .Z(n77282) );
  IV U93052 ( .A(n72867), .Z(n72868) );
  NOR U93053 ( .A(n72869), .B(n72868), .Z(n77278) );
  IV U93054 ( .A(n72870), .Z(n72871) );
  NOR U93055 ( .A(n72872), .B(n72871), .Z(n77280) );
  NOR U93056 ( .A(n77278), .B(n77280), .Z(n72873) );
  XOR U93057 ( .A(n77282), .B(n72873), .Z(n77276) );
  XOR U93058 ( .A(n77277), .B(n77276), .Z(n78330) );
  IV U93059 ( .A(n72874), .Z(n72876) );
  IV U93060 ( .A(n72875), .Z(n72879) );
  NOR U93061 ( .A(n72876), .B(n72879), .Z(n78328) );
  IV U93062 ( .A(n72877), .Z(n72878) );
  NOR U93063 ( .A(n72879), .B(n72878), .Z(n77274) );
  NOR U93064 ( .A(n78328), .B(n77274), .Z(n72880) );
  XOR U93065 ( .A(n78330), .B(n72880), .Z(n72881) );
  NOR U93066 ( .A(n72882), .B(n72881), .Z(n72885) );
  IV U93067 ( .A(n72882), .Z(n72884) );
  XOR U93068 ( .A(n77274), .B(n78330), .Z(n72883) );
  NOR U93069 ( .A(n72884), .B(n72883), .Z(n78327) );
  NOR U93070 ( .A(n72885), .B(n78327), .Z(n72891) );
  IV U93071 ( .A(n72891), .Z(n77273) );
  NOR U93072 ( .A(n72886), .B(n77273), .Z(n83010) );
  IV U93073 ( .A(n72887), .Z(n72888) );
  NOR U93074 ( .A(n72889), .B(n72888), .Z(n72890) );
  IV U93075 ( .A(n72890), .Z(n77272) );
  XOR U93076 ( .A(n72891), .B(n77272), .Z(n77270) );
  IV U93077 ( .A(n77270), .Z(n72892) );
  NOR U93078 ( .A(n72893), .B(n72892), .Z(n72894) );
  NOR U93079 ( .A(n83010), .B(n72894), .Z(n78338) );
  XOR U93080 ( .A(n72895), .B(n78338), .Z(n78343) );
  XOR U93081 ( .A(n78341), .B(n78343), .Z(n78345) );
  IV U93082 ( .A(n78345), .Z(n72903) );
  IV U93083 ( .A(n72896), .Z(n72898) );
  NOR U93084 ( .A(n72898), .B(n72897), .Z(n78344) );
  IV U93085 ( .A(n72899), .Z(n72900) );
  NOR U93086 ( .A(n72901), .B(n72900), .Z(n77267) );
  NOR U93087 ( .A(n78344), .B(n77267), .Z(n72902) );
  XOR U93088 ( .A(n72903), .B(n72902), .Z(n77263) );
  XOR U93089 ( .A(n77262), .B(n77263), .Z(n78352) );
  XOR U93090 ( .A(n72904), .B(n78352), .Z(n78354) );
  XOR U93091 ( .A(n72905), .B(n78354), .Z(n78364) );
  XOR U93092 ( .A(n78363), .B(n78364), .Z(n77260) );
  XOR U93093 ( .A(n77259), .B(n77260), .Z(n78374) );
  XOR U93094 ( .A(n78373), .B(n78374), .Z(n82979) );
  XOR U93095 ( .A(n78376), .B(n82979), .Z(n72906) );
  IV U93096 ( .A(n72906), .Z(n78380) );
  XOR U93097 ( .A(n78379), .B(n78380), .Z(n78383) );
  XOR U93098 ( .A(n78382), .B(n78383), .Z(n77257) );
  XOR U93099 ( .A(n77256), .B(n77257), .Z(n78389) );
  IV U93100 ( .A(n72907), .Z(n72909) );
  NOR U93101 ( .A(n72909), .B(n72908), .Z(n78387) );
  XOR U93102 ( .A(n78389), .B(n78387), .Z(n78392) );
  IV U93103 ( .A(n72910), .Z(n72912) );
  NOR U93104 ( .A(n72912), .B(n72911), .Z(n78390) );
  XOR U93105 ( .A(n78392), .B(n78390), .Z(n78397) );
  XOR U93106 ( .A(n78396), .B(n78397), .Z(n78414) );
  IV U93107 ( .A(n72913), .Z(n72914) );
  NOR U93108 ( .A(n72915), .B(n72914), .Z(n78413) );
  NOR U93109 ( .A(n78413), .B(n77252), .Z(n72916) );
  XOR U93110 ( .A(n78414), .B(n72916), .Z(n77249) );
  IV U93111 ( .A(n72917), .Z(n72918) );
  NOR U93112 ( .A(n72919), .B(n72918), .Z(n77253) );
  IV U93113 ( .A(n72920), .Z(n72921) );
  NOR U93114 ( .A(n72922), .B(n72921), .Z(n77248) );
  NOR U93115 ( .A(n77253), .B(n77248), .Z(n72923) );
  XOR U93116 ( .A(n77249), .B(n72923), .Z(n78430) );
  XOR U93117 ( .A(n78428), .B(n78430), .Z(n78433) );
  IV U93118 ( .A(n72924), .Z(n72926) );
  NOR U93119 ( .A(n72926), .B(n72925), .Z(n78431) );
  XOR U93120 ( .A(n78433), .B(n78431), .Z(n77246) );
  IV U93121 ( .A(n72927), .Z(n72929) );
  NOR U93122 ( .A(n72929), .B(n72928), .Z(n77245) );
  NOR U93123 ( .A(n72931), .B(n72930), .Z(n77243) );
  NOR U93124 ( .A(n77245), .B(n77243), .Z(n72932) );
  XOR U93125 ( .A(n77246), .B(n72932), .Z(n78436) );
  XOR U93126 ( .A(n72933), .B(n78436), .Z(n78454) );
  XOR U93127 ( .A(n72934), .B(n78454), .Z(n78455) );
  XOR U93128 ( .A(n78456), .B(n78455), .Z(n78464) );
  IV U93129 ( .A(n72935), .Z(n72936) );
  NOR U93130 ( .A(n72937), .B(n72936), .Z(n78463) );
  IV U93131 ( .A(n72938), .Z(n72939) );
  NOR U93132 ( .A(n72940), .B(n72939), .Z(n78458) );
  NOR U93133 ( .A(n78463), .B(n78458), .Z(n72941) );
  XOR U93134 ( .A(n78464), .B(n72941), .Z(n78461) );
  XOR U93135 ( .A(n78462), .B(n78461), .Z(n77237) );
  IV U93136 ( .A(n72942), .Z(n72946) );
  NOR U93137 ( .A(n72944), .B(n72943), .Z(n72945) );
  IV U93138 ( .A(n72945), .Z(n72949) );
  NOR U93139 ( .A(n72946), .B(n72949), .Z(n72955) );
  IV U93140 ( .A(n72955), .Z(n72947) );
  NOR U93141 ( .A(n77237), .B(n72947), .Z(n84215) );
  IV U93142 ( .A(n72948), .Z(n72950) );
  NOR U93143 ( .A(n72950), .B(n72949), .Z(n77239) );
  IV U93144 ( .A(n72951), .Z(n72952) );
  NOR U93145 ( .A(n72953), .B(n72952), .Z(n77236) );
  XOR U93146 ( .A(n77236), .B(n77237), .Z(n77240) );
  XOR U93147 ( .A(n77239), .B(n77240), .Z(n77234) );
  IV U93148 ( .A(n77234), .Z(n72954) );
  NOR U93149 ( .A(n72955), .B(n72954), .Z(n72956) );
  NOR U93150 ( .A(n84215), .B(n72956), .Z(n77226) );
  XOR U93151 ( .A(n72957), .B(n77226), .Z(n82935) );
  XOR U93152 ( .A(n77225), .B(n82935), .Z(n77219) );
  XOR U93153 ( .A(n77221), .B(n77219), .Z(n77223) );
  XOR U93154 ( .A(n77222), .B(n77223), .Z(n77214) );
  IV U93155 ( .A(n72958), .Z(n72960) );
  NOR U93156 ( .A(n72960), .B(n72959), .Z(n77217) );
  IV U93157 ( .A(n72961), .Z(n72963) );
  NOR U93158 ( .A(n72963), .B(n72962), .Z(n77213) );
  NOR U93159 ( .A(n77217), .B(n77213), .Z(n72964) );
  XOR U93160 ( .A(n77214), .B(n72964), .Z(n72965) );
  IV U93161 ( .A(n72965), .Z(n78474) );
  XOR U93162 ( .A(n78472), .B(n78474), .Z(n77211) );
  IV U93163 ( .A(n77211), .Z(n72973) );
  IV U93164 ( .A(n72966), .Z(n72968) );
  NOR U93165 ( .A(n72968), .B(n72967), .Z(n77205) );
  IV U93166 ( .A(n72969), .Z(n72970) );
  NOR U93167 ( .A(n72971), .B(n72970), .Z(n77210) );
  NOR U93168 ( .A(n77205), .B(n77210), .Z(n72972) );
  XOR U93169 ( .A(n72973), .B(n72972), .Z(n77209) );
  XOR U93170 ( .A(n77207), .B(n77209), .Z(n78484) );
  XOR U93171 ( .A(n72974), .B(n78484), .Z(n77197) );
  IV U93172 ( .A(n72975), .Z(n72976) );
  NOR U93173 ( .A(n72977), .B(n72976), .Z(n78486) );
  IV U93174 ( .A(n72978), .Z(n72979) );
  NOR U93175 ( .A(n72980), .B(n72979), .Z(n77196) );
  NOR U93176 ( .A(n78486), .B(n77196), .Z(n72981) );
  XOR U93177 ( .A(n77197), .B(n72981), .Z(n78492) );
  XOR U93178 ( .A(n72982), .B(n78492), .Z(n78496) );
  XOR U93179 ( .A(n78494), .B(n78496), .Z(n72995) );
  IV U93180 ( .A(n72995), .Z(n72991) );
  IV U93181 ( .A(n72983), .Z(n72985) );
  NOR U93182 ( .A(n72985), .B(n72984), .Z(n72994) );
  IV U93183 ( .A(n72986), .Z(n72988) );
  NOR U93184 ( .A(n72988), .B(n72987), .Z(n72992) );
  NOR U93185 ( .A(n72994), .B(n72992), .Z(n72989) );
  IV U93186 ( .A(n72989), .Z(n72990) );
  NOR U93187 ( .A(n72991), .B(n72990), .Z(n72998) );
  IV U93188 ( .A(n72992), .Z(n72993) );
  NOR U93189 ( .A(n78496), .B(n72993), .Z(n78501) );
  IV U93190 ( .A(n72994), .Z(n72996) );
  NOR U93191 ( .A(n72996), .B(n72995), .Z(n78497) );
  NOR U93192 ( .A(n78501), .B(n78497), .Z(n84257) );
  IV U93193 ( .A(n84257), .Z(n72997) );
  NOR U93194 ( .A(n72998), .B(n72997), .Z(n72999) );
  IV U93195 ( .A(n72999), .Z(n78504) );
  XOR U93196 ( .A(n78499), .B(n78504), .Z(n77195) );
  IV U93197 ( .A(n73000), .Z(n73001) );
  NOR U93198 ( .A(n73002), .B(n73001), .Z(n78503) );
  IV U93199 ( .A(n73003), .Z(n73004) );
  NOR U93200 ( .A(n73007), .B(n73004), .Z(n77193) );
  NOR U93201 ( .A(n78503), .B(n77193), .Z(n73005) );
  XOR U93202 ( .A(n77195), .B(n73005), .Z(n78507) );
  IV U93203 ( .A(n73006), .Z(n73008) );
  NOR U93204 ( .A(n73008), .B(n73007), .Z(n78506) );
  IV U93205 ( .A(n78506), .Z(n78508) );
  XOR U93206 ( .A(n78507), .B(n78508), .Z(n78519) );
  XOR U93207 ( .A(n73009), .B(n78519), .Z(n78514) );
  XOR U93208 ( .A(n78515), .B(n78514), .Z(n78521) );
  NOR U93209 ( .A(n73010), .B(n78521), .Z(n78523) );
  IV U93210 ( .A(n78523), .Z(n82898) );
  IV U93211 ( .A(n73011), .Z(n73013) );
  NOR U93212 ( .A(n73013), .B(n73012), .Z(n73024) );
  IV U93213 ( .A(n73014), .Z(n73016) );
  NOR U93214 ( .A(n73016), .B(n73015), .Z(n73017) );
  IV U93215 ( .A(n73017), .Z(n77191) );
  IV U93216 ( .A(n73018), .Z(n73019) );
  NOR U93217 ( .A(n73020), .B(n73019), .Z(n73021) );
  IV U93218 ( .A(n73021), .Z(n78522) );
  XOR U93219 ( .A(n78522), .B(n78521), .Z(n73022) );
  NOR U93220 ( .A(n73023), .B(n73022), .Z(n77192) );
  IV U93221 ( .A(n73024), .Z(n73025) );
  NOR U93222 ( .A(n73025), .B(n78521), .Z(n82892) );
  XOR U93223 ( .A(n78525), .B(n78526), .Z(n77189) );
  IV U93224 ( .A(n73026), .Z(n73027) );
  NOR U93225 ( .A(n73028), .B(n73027), .Z(n77188) );
  IV U93226 ( .A(n73029), .Z(n73031) );
  NOR U93227 ( .A(n73031), .B(n73030), .Z(n77181) );
  NOR U93228 ( .A(n77188), .B(n77181), .Z(n73032) );
  XOR U93229 ( .A(n77189), .B(n73032), .Z(n73033) );
  IV U93230 ( .A(n73033), .Z(n77184) );
  XOR U93231 ( .A(n77183), .B(n77184), .Z(n78531) );
  XOR U93232 ( .A(n73034), .B(n78531), .Z(n73035) );
  IV U93233 ( .A(n73035), .Z(n78535) );
  XOR U93234 ( .A(n78533), .B(n78535), .Z(n84282) );
  IV U93235 ( .A(n73036), .Z(n73038) );
  NOR U93236 ( .A(n73038), .B(n73037), .Z(n84281) );
  IV U93237 ( .A(n73039), .Z(n73041) );
  NOR U93238 ( .A(n73041), .B(n73040), .Z(n84296) );
  NOR U93239 ( .A(n84281), .B(n84296), .Z(n78536) );
  XOR U93240 ( .A(n84282), .B(n78536), .Z(n73042) );
  IV U93241 ( .A(n73042), .Z(n78544) );
  IV U93242 ( .A(n73043), .Z(n73045) );
  NOR U93243 ( .A(n73045), .B(n73044), .Z(n78543) );
  IV U93244 ( .A(n73046), .Z(n73047) );
  NOR U93245 ( .A(n73048), .B(n73047), .Z(n78541) );
  NOR U93246 ( .A(n78543), .B(n78541), .Z(n73049) );
  XOR U93247 ( .A(n78544), .B(n73049), .Z(n73050) );
  NOR U93248 ( .A(n73051), .B(n73050), .Z(n73054) );
  IV U93249 ( .A(n73051), .Z(n73053) );
  XOR U93250 ( .A(n78543), .B(n78544), .Z(n73052) );
  NOR U93251 ( .A(n73053), .B(n73052), .Z(n78553) );
  NOR U93252 ( .A(n73054), .B(n78553), .Z(n77165) );
  IV U93253 ( .A(n73055), .Z(n73057) );
  NOR U93254 ( .A(n73057), .B(n73056), .Z(n73058) );
  IV U93255 ( .A(n73058), .Z(n77166) );
  XOR U93256 ( .A(n77165), .B(n77166), .Z(n77169) );
  XOR U93257 ( .A(n77168), .B(n77169), .Z(n82855) );
  IV U93258 ( .A(n73059), .Z(n73060) );
  NOR U93259 ( .A(n73061), .B(n73060), .Z(n82863) );
  IV U93260 ( .A(n73062), .Z(n73063) );
  NOR U93261 ( .A(n73063), .B(n78566), .Z(n82854) );
  NOR U93262 ( .A(n82863), .B(n82854), .Z(n78556) );
  XOR U93263 ( .A(n82855), .B(n78556), .Z(n73064) );
  IV U93264 ( .A(n73064), .Z(n78565) );
  XOR U93265 ( .A(n73070), .B(n78565), .Z(n73065) );
  NOR U93266 ( .A(n73066), .B(n73065), .Z(n82851) );
  IV U93267 ( .A(n73067), .Z(n73068) );
  NOR U93268 ( .A(n73069), .B(n73068), .Z(n78558) );
  NOR U93269 ( .A(n73070), .B(n78558), .Z(n73071) );
  XOR U93270 ( .A(n73071), .B(n78565), .Z(n77162) );
  NOR U93271 ( .A(n73072), .B(n77162), .Z(n73073) );
  NOR U93272 ( .A(n82851), .B(n73073), .Z(n77158) );
  XOR U93273 ( .A(n73074), .B(n77158), .Z(n77153) );
  XOR U93274 ( .A(n77151), .B(n77153), .Z(n78581) );
  XOR U93275 ( .A(n77154), .B(n78581), .Z(n73075) );
  XOR U93276 ( .A(n73076), .B(n73075), .Z(n78577) );
  XOR U93277 ( .A(n73088), .B(n78577), .Z(n73081) );
  IV U93278 ( .A(n73077), .Z(n73079) );
  NOR U93279 ( .A(n73079), .B(n73078), .Z(n73080) );
  IV U93280 ( .A(n73080), .Z(n73096) );
  NOR U93281 ( .A(n73081), .B(n73096), .Z(n82839) );
  IV U93282 ( .A(n78577), .Z(n73092) );
  IV U93283 ( .A(n73082), .Z(n73084) );
  IV U93284 ( .A(n73083), .Z(n73086) );
  NOR U93285 ( .A(n73084), .B(n73086), .Z(n77146) );
  IV U93286 ( .A(n73085), .Z(n73087) );
  NOR U93287 ( .A(n73087), .B(n73086), .Z(n77149) );
  NOR U93288 ( .A(n73088), .B(n77149), .Z(n73089) );
  IV U93289 ( .A(n73089), .Z(n73090) );
  NOR U93290 ( .A(n77146), .B(n73090), .Z(n73091) );
  XOR U93291 ( .A(n73092), .B(n73091), .Z(n77145) );
  IV U93292 ( .A(n73093), .Z(n73095) );
  NOR U93293 ( .A(n73095), .B(n73094), .Z(n73097) );
  IV U93294 ( .A(n73097), .Z(n77144) );
  XOR U93295 ( .A(n77145), .B(n77144), .Z(n73099) );
  NOR U93296 ( .A(n73097), .B(n73096), .Z(n73098) );
  NOR U93297 ( .A(n73099), .B(n73098), .Z(n73100) );
  NOR U93298 ( .A(n82839), .B(n73100), .Z(n77135) );
  XOR U93299 ( .A(n73101), .B(n77135), .Z(n78600) );
  XOR U93300 ( .A(n78598), .B(n78600), .Z(n78603) );
  IV U93301 ( .A(n73102), .Z(n73104) );
  NOR U93302 ( .A(n73104), .B(n73103), .Z(n78601) );
  XOR U93303 ( .A(n78603), .B(n78601), .Z(n77130) );
  IV U93304 ( .A(n73105), .Z(n73106) );
  NOR U93305 ( .A(n73107), .B(n73106), .Z(n77128) );
  XOR U93306 ( .A(n77130), .B(n77128), .Z(n77132) );
  XOR U93307 ( .A(n77131), .B(n77132), .Z(n77123) );
  XOR U93308 ( .A(n77122), .B(n77123), .Z(n77126) );
  IV U93309 ( .A(n73108), .Z(n73110) );
  NOR U93310 ( .A(n73110), .B(n73109), .Z(n77125) );
  IV U93311 ( .A(n73111), .Z(n73113) );
  NOR U93312 ( .A(n73113), .B(n73112), .Z(n77119) );
  NOR U93313 ( .A(n77125), .B(n77119), .Z(n73114) );
  XOR U93314 ( .A(n77126), .B(n73114), .Z(n77113) );
  IV U93315 ( .A(n73115), .Z(n73116) );
  NOR U93316 ( .A(n73116), .B(n73118), .Z(n77116) );
  IV U93317 ( .A(n73117), .Z(n73119) );
  NOR U93318 ( .A(n73119), .B(n73118), .Z(n77112) );
  NOR U93319 ( .A(n77116), .B(n77112), .Z(n73120) );
  XOR U93320 ( .A(n77113), .B(n73120), .Z(n77110) );
  XOR U93321 ( .A(n73121), .B(n77110), .Z(n77099) );
  IV U93322 ( .A(n77099), .Z(n77104) );
  XOR U93323 ( .A(n73122), .B(n77104), .Z(n77094) );
  IV U93324 ( .A(n73123), .Z(n73124) );
  NOR U93325 ( .A(n73125), .B(n73124), .Z(n77098) );
  IV U93326 ( .A(n73126), .Z(n73128) );
  NOR U93327 ( .A(n73128), .B(n73127), .Z(n77093) );
  NOR U93328 ( .A(n77098), .B(n77093), .Z(n73129) );
  XOR U93329 ( .A(n77094), .B(n73129), .Z(n77092) );
  XOR U93330 ( .A(n77091), .B(n77092), .Z(n77089) );
  IV U93331 ( .A(n73130), .Z(n73131) );
  NOR U93332 ( .A(n73132), .B(n73131), .Z(n77088) );
  IV U93333 ( .A(n73133), .Z(n73135) );
  NOR U93334 ( .A(n73135), .B(n73134), .Z(n78612) );
  NOR U93335 ( .A(n77088), .B(n78612), .Z(n73136) );
  XOR U93336 ( .A(n77089), .B(n73136), .Z(n77086) );
  XOR U93337 ( .A(n77084), .B(n77086), .Z(n78610) );
  XOR U93338 ( .A(n78609), .B(n78610), .Z(n73145) );
  IV U93339 ( .A(n73145), .Z(n73151) );
  NOR U93340 ( .A(n73142), .B(n73151), .Z(n73141) );
  IV U93341 ( .A(n73137), .Z(n73139) );
  IV U93342 ( .A(n73138), .Z(n73144) );
  NOR U93343 ( .A(n73139), .B(n73144), .Z(n73148) );
  IV U93344 ( .A(n73148), .Z(n73140) );
  NOR U93345 ( .A(n73141), .B(n73140), .Z(n78624) );
  IV U93346 ( .A(n73142), .Z(n73143) );
  NOR U93347 ( .A(n73144), .B(n73143), .Z(n73147) );
  IV U93348 ( .A(n73147), .Z(n73146) );
  NOR U93349 ( .A(n73146), .B(n73145), .Z(n82765) );
  NOR U93350 ( .A(n73148), .B(n73147), .Z(n73149) );
  IV U93351 ( .A(n73149), .Z(n73150) );
  NOR U93352 ( .A(n73151), .B(n73150), .Z(n73152) );
  NOR U93353 ( .A(n82765), .B(n73152), .Z(n73153) );
  IV U93354 ( .A(n73153), .Z(n78621) );
  NOR U93355 ( .A(n78624), .B(n78621), .Z(n78628) );
  IV U93356 ( .A(n73154), .Z(n73155) );
  NOR U93357 ( .A(n73156), .B(n73155), .Z(n78620) );
  IV U93358 ( .A(n73157), .Z(n73158) );
  NOR U93359 ( .A(n73159), .B(n73158), .Z(n78627) );
  NOR U93360 ( .A(n78620), .B(n78627), .Z(n73160) );
  XOR U93361 ( .A(n78628), .B(n73160), .Z(n84350) );
  XOR U93362 ( .A(n84343), .B(n84350), .Z(n77082) );
  XOR U93363 ( .A(n73161), .B(n77082), .Z(n73162) );
  IV U93364 ( .A(n73162), .Z(n78640) );
  XOR U93365 ( .A(n78638), .B(n78640), .Z(n78642) );
  XOR U93366 ( .A(n78641), .B(n78642), .Z(n73173) );
  IV U93367 ( .A(n73173), .Z(n73171) );
  IV U93368 ( .A(n73163), .Z(n73165) );
  NOR U93369 ( .A(n73165), .B(n73164), .Z(n73175) );
  IV U93370 ( .A(n73166), .Z(n73168) );
  IV U93371 ( .A(n73167), .Z(n73184) );
  NOR U93372 ( .A(n73168), .B(n73184), .Z(n73172) );
  NOR U93373 ( .A(n73175), .B(n73172), .Z(n73169) );
  IV U93374 ( .A(n73169), .Z(n73170) );
  NOR U93375 ( .A(n73171), .B(n73170), .Z(n73179) );
  IV U93376 ( .A(n73172), .Z(n73174) );
  NOR U93377 ( .A(n73174), .B(n73173), .Z(n73178) );
  IV U93378 ( .A(n73175), .Z(n73176) );
  NOR U93379 ( .A(n78642), .B(n73176), .Z(n73177) );
  NOR U93380 ( .A(n73178), .B(n73177), .Z(n82754) );
  IV U93381 ( .A(n82754), .Z(n78648) );
  NOR U93382 ( .A(n73179), .B(n78648), .Z(n78646) );
  IV U93383 ( .A(n73180), .Z(n73181) );
  NOR U93384 ( .A(n73182), .B(n73181), .Z(n78650) );
  IV U93385 ( .A(n73183), .Z(n73185) );
  NOR U93386 ( .A(n73185), .B(n73184), .Z(n78645) );
  NOR U93387 ( .A(n78650), .B(n78645), .Z(n73186) );
  XOR U93388 ( .A(n78646), .B(n73186), .Z(n78654) );
  XOR U93389 ( .A(n73187), .B(n78654), .Z(n73188) );
  IV U93390 ( .A(n73188), .Z(n77075) );
  IV U93391 ( .A(n73189), .Z(n73190) );
  NOR U93392 ( .A(n73191), .B(n73190), .Z(n77073) );
  XOR U93393 ( .A(n77075), .B(n77073), .Z(n77077) );
  IV U93394 ( .A(n77077), .Z(n73199) );
  IV U93395 ( .A(n73192), .Z(n73193) );
  NOR U93396 ( .A(n73194), .B(n73193), .Z(n77076) );
  IV U93397 ( .A(n73195), .Z(n73196) );
  NOR U93398 ( .A(n73197), .B(n73196), .Z(n77071) );
  NOR U93399 ( .A(n77076), .B(n77071), .Z(n73198) );
  XOR U93400 ( .A(n73199), .B(n73198), .Z(n77070) );
  XOR U93401 ( .A(n77068), .B(n77070), .Z(n77064) );
  XOR U93402 ( .A(n73200), .B(n77064), .Z(n77056) );
  XOR U93403 ( .A(n77057), .B(n77056), .Z(n77053) );
  IV U93404 ( .A(n73201), .Z(n73202) );
  NOR U93405 ( .A(n73203), .B(n73202), .Z(n77052) );
  IV U93406 ( .A(n73204), .Z(n73205) );
  NOR U93407 ( .A(n73206), .B(n73205), .Z(n77059) );
  NOR U93408 ( .A(n77052), .B(n77059), .Z(n73207) );
  XOR U93409 ( .A(n77053), .B(n73207), .Z(n77046) );
  IV U93410 ( .A(n73208), .Z(n73210) );
  NOR U93411 ( .A(n73210), .B(n73209), .Z(n77049) );
  IV U93412 ( .A(n73211), .Z(n73213) );
  NOR U93413 ( .A(n73213), .B(n73212), .Z(n77047) );
  NOR U93414 ( .A(n77049), .B(n77047), .Z(n73214) );
  XOR U93415 ( .A(n77046), .B(n73214), .Z(n82725) );
  IV U93416 ( .A(n73215), .Z(n73216) );
  NOR U93417 ( .A(n73217), .B(n73216), .Z(n82728) );
  IV U93418 ( .A(n73218), .Z(n73219) );
  NOR U93419 ( .A(n73220), .B(n73219), .Z(n82724) );
  NOR U93420 ( .A(n82728), .B(n82724), .Z(n77039) );
  XOR U93421 ( .A(n82725), .B(n77039), .Z(n77037) );
  XOR U93422 ( .A(n73221), .B(n77037), .Z(n77035) );
  IV U93423 ( .A(n73222), .Z(n73224) );
  NOR U93424 ( .A(n73224), .B(n73223), .Z(n77033) );
  IV U93425 ( .A(n73225), .Z(n73229) );
  NOR U93426 ( .A(n73226), .B(n73238), .Z(n73227) );
  IV U93427 ( .A(n73227), .Z(n73228) );
  NOR U93428 ( .A(n73229), .B(n73228), .Z(n77028) );
  NOR U93429 ( .A(n77033), .B(n77028), .Z(n73230) );
  XOR U93430 ( .A(n77035), .B(n73230), .Z(n77025) );
  IV U93431 ( .A(n73231), .Z(n73236) );
  IV U93432 ( .A(n73232), .Z(n73233) );
  NOR U93433 ( .A(n73233), .B(n73238), .Z(n73234) );
  IV U93434 ( .A(n73234), .Z(n73235) );
  NOR U93435 ( .A(n73236), .B(n73235), .Z(n77030) );
  IV U93436 ( .A(n73237), .Z(n73239) );
  NOR U93437 ( .A(n73239), .B(n73238), .Z(n77026) );
  NOR U93438 ( .A(n77030), .B(n77026), .Z(n73240) );
  XOR U93439 ( .A(n77025), .B(n73240), .Z(n77017) );
  IV U93440 ( .A(n73241), .Z(n73242) );
  NOR U93441 ( .A(n73243), .B(n73242), .Z(n77019) );
  XOR U93442 ( .A(n77017), .B(n77019), .Z(n77011) );
  XOR U93443 ( .A(n73244), .B(n77011), .Z(n77006) );
  XOR U93444 ( .A(n73245), .B(n77006), .Z(n77001) );
  XOR U93445 ( .A(n76999), .B(n77001), .Z(n77003) );
  XOR U93446 ( .A(n77002), .B(n77003), .Z(n76997) );
  XOR U93447 ( .A(n73246), .B(n76997), .Z(n76988) );
  IV U93448 ( .A(n73247), .Z(n73249) );
  NOR U93449 ( .A(n73249), .B(n73248), .Z(n76987) );
  IV U93450 ( .A(n73250), .Z(n73251) );
  NOR U93451 ( .A(n73252), .B(n73251), .Z(n76990) );
  NOR U93452 ( .A(n76987), .B(n76990), .Z(n73253) );
  XOR U93453 ( .A(n76988), .B(n73253), .Z(n82688) );
  XOR U93454 ( .A(n73254), .B(n82688), .Z(n76978) );
  XOR U93455 ( .A(n73255), .B(n76978), .Z(n76976) );
  XOR U93456 ( .A(n76975), .B(n76976), .Z(n76972) );
  XOR U93457 ( .A(n73256), .B(n76972), .Z(n76965) );
  XOR U93458 ( .A(n73257), .B(n76965), .Z(n76963) );
  XOR U93459 ( .A(n73258), .B(n76963), .Z(n76957) );
  IV U93460 ( .A(n73259), .Z(n73261) );
  NOR U93461 ( .A(n73261), .B(n73260), .Z(n73262) );
  IV U93462 ( .A(n73262), .Z(n76961) );
  XOR U93463 ( .A(n76961), .B(n73263), .Z(n73264) );
  XOR U93464 ( .A(n76957), .B(n73264), .Z(n76953) );
  IV U93465 ( .A(n73265), .Z(n73266) );
  NOR U93466 ( .A(n73267), .B(n73266), .Z(n76954) );
  IV U93467 ( .A(n73268), .Z(n73270) );
  NOR U93468 ( .A(n73270), .B(n73269), .Z(n78665) );
  NOR U93469 ( .A(n76954), .B(n78665), .Z(n73271) );
  XOR U93470 ( .A(n76953), .B(n73271), .Z(n76950) );
  XOR U93471 ( .A(n76949), .B(n76950), .Z(n76944) );
  IV U93472 ( .A(n73272), .Z(n73273) );
  NOR U93473 ( .A(n73274), .B(n73273), .Z(n76948) );
  NOR U93474 ( .A(n73275), .B(n76945), .Z(n73276) );
  NOR U93475 ( .A(n76948), .B(n73276), .Z(n73277) );
  XOR U93476 ( .A(n76944), .B(n73277), .Z(n73278) );
  IV U93477 ( .A(n73278), .Z(n78674) );
  NOR U93478 ( .A(n73280), .B(n73279), .Z(n73281) );
  IV U93479 ( .A(n73281), .Z(n73285) );
  NOR U93480 ( .A(n78674), .B(n73285), .Z(n78680) );
  IV U93481 ( .A(n73282), .Z(n73283) );
  NOR U93482 ( .A(n73284), .B(n73283), .Z(n73286) );
  IV U93483 ( .A(n73286), .Z(n78673) );
  XOR U93484 ( .A(n78674), .B(n78673), .Z(n73288) );
  NOR U93485 ( .A(n73286), .B(n73285), .Z(n73287) );
  NOR U93486 ( .A(n73288), .B(n73287), .Z(n82644) );
  NOR U93487 ( .A(n78680), .B(n82644), .Z(n73297) );
  IV U93488 ( .A(n73297), .Z(n73289) );
  NOR U93489 ( .A(n73293), .B(n73289), .Z(n82629) );
  IV U93490 ( .A(n73290), .Z(n73291) );
  NOR U93491 ( .A(n73292), .B(n73291), .Z(n78681) );
  IV U93492 ( .A(n73294), .Z(n82647) );
  NOR U93493 ( .A(n73295), .B(n82647), .Z(n73298) );
  IV U93494 ( .A(n73298), .Z(n73296) );
  NOR U93495 ( .A(n73296), .B(n82644), .Z(n78684) );
  NOR U93496 ( .A(n73298), .B(n73297), .Z(n73299) );
  NOR U93497 ( .A(n78684), .B(n73299), .Z(n73300) );
  IV U93498 ( .A(n73300), .Z(n78682) );
  IV U93499 ( .A(n73301), .Z(n73302) );
  NOR U93500 ( .A(n73303), .B(n73302), .Z(n78688) );
  IV U93501 ( .A(n73304), .Z(n73306) );
  NOR U93502 ( .A(n73306), .B(n73305), .Z(n78693) );
  NOR U93503 ( .A(n78688), .B(n78693), .Z(n73307) );
  XOR U93504 ( .A(n78694), .B(n73307), .Z(n76937) );
  XOR U93505 ( .A(n73308), .B(n76937), .Z(n76941) );
  XOR U93506 ( .A(n73309), .B(n76941), .Z(n78702) );
  XOR U93507 ( .A(n78703), .B(n78702), .Z(n76928) );
  XOR U93508 ( .A(n73310), .B(n76928), .Z(n76919) );
  XOR U93509 ( .A(n76917), .B(n76919), .Z(n78708) );
  XOR U93510 ( .A(n76915), .B(n78708), .Z(n76913) );
  IV U93511 ( .A(n73311), .Z(n73327) );
  NOR U93512 ( .A(n73312), .B(n73327), .Z(n78707) );
  IV U93513 ( .A(n73313), .Z(n73315) );
  NOR U93514 ( .A(n73315), .B(n73314), .Z(n76911) );
  NOR U93515 ( .A(n78707), .B(n76911), .Z(n73316) );
  XOR U93516 ( .A(n76913), .B(n73316), .Z(n73317) );
  IV U93517 ( .A(n73317), .Z(n78712) );
  IV U93518 ( .A(n73318), .Z(n73320) );
  NOR U93519 ( .A(n73320), .B(n73319), .Z(n73321) );
  IV U93520 ( .A(n73321), .Z(n73328) );
  NOR U93521 ( .A(n78712), .B(n73328), .Z(n82593) );
  IV U93522 ( .A(n73322), .Z(n73323) );
  NOR U93523 ( .A(n73324), .B(n73323), .Z(n76908) );
  IV U93524 ( .A(n73325), .Z(n73326) );
  NOR U93525 ( .A(n73327), .B(n73326), .Z(n78710) );
  XOR U93526 ( .A(n78710), .B(n78712), .Z(n76909) );
  IV U93527 ( .A(n76909), .Z(n73329) );
  XOR U93528 ( .A(n76908), .B(n73329), .Z(n73331) );
  NOR U93529 ( .A(n73329), .B(n73328), .Z(n73330) );
  NOR U93530 ( .A(n73331), .B(n73330), .Z(n73332) );
  NOR U93531 ( .A(n82593), .B(n73332), .Z(n76903) );
  IV U93532 ( .A(n73333), .Z(n73335) );
  NOR U93533 ( .A(n73335), .B(n73334), .Z(n76905) );
  IV U93534 ( .A(n73336), .Z(n73338) );
  NOR U93535 ( .A(n73338), .B(n73337), .Z(n76902) );
  NOR U93536 ( .A(n76905), .B(n76902), .Z(n73339) );
  XOR U93537 ( .A(n76903), .B(n73339), .Z(n78718) );
  XOR U93538 ( .A(n78716), .B(n78718), .Z(n73340) );
  NOR U93539 ( .A(n73341), .B(n73340), .Z(n76901) );
  IV U93540 ( .A(n73342), .Z(n73344) );
  NOR U93541 ( .A(n73344), .B(n73343), .Z(n78714) );
  NOR U93542 ( .A(n78716), .B(n78714), .Z(n73345) );
  XOR U93543 ( .A(n78718), .B(n73345), .Z(n76898) );
  NOR U93544 ( .A(n73346), .B(n76898), .Z(n73347) );
  NOR U93545 ( .A(n76901), .B(n73347), .Z(n76893) );
  XOR U93546 ( .A(n73348), .B(n76893), .Z(n76892) );
  XOR U93547 ( .A(n76890), .B(n76892), .Z(n78729) );
  IV U93548 ( .A(n73349), .Z(n73354) );
  IV U93549 ( .A(n73350), .Z(n73351) );
  NOR U93550 ( .A(n73354), .B(n73351), .Z(n78727) );
  XOR U93551 ( .A(n78729), .B(n78727), .Z(n76889) );
  IV U93552 ( .A(n73352), .Z(n73353) );
  NOR U93553 ( .A(n73354), .B(n73353), .Z(n76887) );
  XOR U93554 ( .A(n76889), .B(n76887), .Z(n78755) );
  XOR U93555 ( .A(n78738), .B(n78755), .Z(n78734) );
  IV U93556 ( .A(n73355), .Z(n73356) );
  NOR U93557 ( .A(n73357), .B(n73356), .Z(n78733) );
  IV U93558 ( .A(n73358), .Z(n73365) );
  IV U93559 ( .A(n73359), .Z(n73360) );
  NOR U93560 ( .A(n73365), .B(n73360), .Z(n78753) );
  NOR U93561 ( .A(n78733), .B(n78753), .Z(n73361) );
  XOR U93562 ( .A(n78734), .B(n73361), .Z(n73362) );
  IV U93563 ( .A(n73362), .Z(n78752) );
  IV U93564 ( .A(n73363), .Z(n73364) );
  NOR U93565 ( .A(n73365), .B(n73364), .Z(n78750) );
  XOR U93566 ( .A(n78752), .B(n78750), .Z(n76885) );
  XOR U93567 ( .A(n73366), .B(n76885), .Z(n76879) );
  XOR U93568 ( .A(n73367), .B(n76879), .Z(n78767) );
  XOR U93569 ( .A(n73368), .B(n78767), .Z(n76877) );
  XOR U93570 ( .A(n76876), .B(n76877), .Z(n76875) );
  IV U93571 ( .A(n73369), .Z(n73370) );
  NOR U93572 ( .A(n73371), .B(n73370), .Z(n76873) );
  XOR U93573 ( .A(n76875), .B(n76873), .Z(n76869) );
  IV U93574 ( .A(n73372), .Z(n73374) );
  NOR U93575 ( .A(n73374), .B(n73373), .Z(n76868) );
  IV U93576 ( .A(n73375), .Z(n73377) );
  NOR U93577 ( .A(n73377), .B(n73376), .Z(n76866) );
  NOR U93578 ( .A(n76868), .B(n76866), .Z(n73378) );
  XOR U93579 ( .A(n76869), .B(n73378), .Z(n78775) );
  XOR U93580 ( .A(n78776), .B(n78775), .Z(n78780) );
  XOR U93581 ( .A(n78778), .B(n78780), .Z(n78784) );
  XOR U93582 ( .A(n76861), .B(n78784), .Z(n76856) );
  XOR U93583 ( .A(n73379), .B(n76856), .Z(n73380) );
  IV U93584 ( .A(n73380), .Z(n76852) );
  XOR U93585 ( .A(n76850), .B(n76852), .Z(n76848) );
  XOR U93586 ( .A(n76847), .B(n76848), .Z(n76842) );
  IV U93587 ( .A(n73381), .Z(n73383) );
  NOR U93588 ( .A(n73383), .B(n73382), .Z(n76845) );
  IV U93589 ( .A(n73384), .Z(n73385) );
  NOR U93590 ( .A(n73386), .B(n73385), .Z(n76841) );
  NOR U93591 ( .A(n76845), .B(n76841), .Z(n73387) );
  XOR U93592 ( .A(n76842), .B(n73387), .Z(n78790) );
  IV U93593 ( .A(n73388), .Z(n73389) );
  NOR U93594 ( .A(n73390), .B(n73389), .Z(n78791) );
  IV U93595 ( .A(n73391), .Z(n73393) );
  NOR U93596 ( .A(n73393), .B(n73392), .Z(n78795) );
  NOR U93597 ( .A(n78791), .B(n78795), .Z(n73394) );
  XOR U93598 ( .A(n78790), .B(n73394), .Z(n78800) );
  IV U93599 ( .A(n73395), .Z(n73397) );
  NOR U93600 ( .A(n73397), .B(n73396), .Z(n78793) );
  IV U93601 ( .A(n73398), .Z(n73399) );
  NOR U93602 ( .A(n73400), .B(n73399), .Z(n78799) );
  NOR U93603 ( .A(n78793), .B(n78799), .Z(n73401) );
  XOR U93604 ( .A(n78800), .B(n73401), .Z(n76838) );
  IV U93605 ( .A(n73402), .Z(n73403) );
  NOR U93606 ( .A(n73404), .B(n73403), .Z(n76839) );
  IV U93607 ( .A(n73405), .Z(n73406) );
  NOR U93608 ( .A(n73406), .B(n73409), .Z(n78806) );
  NOR U93609 ( .A(n76839), .B(n78806), .Z(n73407) );
  XOR U93610 ( .A(n76838), .B(n73407), .Z(n78805) );
  IV U93611 ( .A(n73408), .Z(n73410) );
  NOR U93612 ( .A(n73410), .B(n73409), .Z(n78803) );
  XOR U93613 ( .A(n78805), .B(n78803), .Z(n76836) );
  IV U93614 ( .A(n73411), .Z(n73413) );
  NOR U93615 ( .A(n73413), .B(n73412), .Z(n76835) );
  IV U93616 ( .A(n73414), .Z(n73415) );
  NOR U93617 ( .A(n73415), .B(n73418), .Z(n76832) );
  NOR U93618 ( .A(n76835), .B(n76832), .Z(n73416) );
  XOR U93619 ( .A(n76836), .B(n73416), .Z(n76830) );
  IV U93620 ( .A(n73417), .Z(n73419) );
  NOR U93621 ( .A(n73419), .B(n73418), .Z(n84562) );
  IV U93622 ( .A(n73420), .Z(n73422) );
  IV U93623 ( .A(n73421), .Z(n73424) );
  NOR U93624 ( .A(n73422), .B(n73424), .Z(n82496) );
  NOR U93625 ( .A(n84562), .B(n82496), .Z(n76831) );
  XOR U93626 ( .A(n76830), .B(n76831), .Z(n76828) );
  IV U93627 ( .A(n73423), .Z(n73425) );
  NOR U93628 ( .A(n73425), .B(n73424), .Z(n76827) );
  IV U93629 ( .A(n73426), .Z(n73428) );
  NOR U93630 ( .A(n73428), .B(n73427), .Z(n76825) );
  NOR U93631 ( .A(n76827), .B(n76825), .Z(n73429) );
  XOR U93632 ( .A(n76828), .B(n73429), .Z(n76819) );
  IV U93633 ( .A(n76819), .Z(n76817) );
  XOR U93634 ( .A(n76820), .B(n76817), .Z(n90423) );
  XOR U93635 ( .A(n90424), .B(n90423), .Z(n78829) );
  IV U93636 ( .A(n73430), .Z(n73432) );
  NOR U93637 ( .A(n73432), .B(n73431), .Z(n78816) );
  IV U93638 ( .A(n73433), .Z(n73434) );
  NOR U93639 ( .A(n73435), .B(n73434), .Z(n76815) );
  NOR U93640 ( .A(n78816), .B(n76815), .Z(n73436) );
  XOR U93641 ( .A(n78829), .B(n73436), .Z(n76813) );
  XOR U93642 ( .A(n73437), .B(n76813), .Z(n76802) );
  XOR U93643 ( .A(n76808), .B(n76802), .Z(n76806) );
  IV U93644 ( .A(n73438), .Z(n73440) );
  NOR U93645 ( .A(n73440), .B(n73439), .Z(n76803) );
  IV U93646 ( .A(n73441), .Z(n73443) );
  NOR U93647 ( .A(n73443), .B(n73442), .Z(n76805) );
  NOR U93648 ( .A(n76803), .B(n76805), .Z(n73444) );
  XOR U93649 ( .A(n76806), .B(n73444), .Z(n76795) );
  IV U93650 ( .A(n73445), .Z(n73446) );
  NOR U93651 ( .A(n73447), .B(n73446), .Z(n76798) );
  IV U93652 ( .A(n73448), .Z(n73450) );
  NOR U93653 ( .A(n73450), .B(n73449), .Z(n76796) );
  NOR U93654 ( .A(n76798), .B(n76796), .Z(n73451) );
  XOR U93655 ( .A(n76795), .B(n73451), .Z(n82460) );
  XOR U93656 ( .A(n78834), .B(n82460), .Z(n78836) );
  XOR U93657 ( .A(n73452), .B(n78836), .Z(n78841) );
  XOR U93658 ( .A(n78840), .B(n78841), .Z(n78846) );
  XOR U93659 ( .A(n78848), .B(n78846), .Z(n78854) );
  XOR U93660 ( .A(n73453), .B(n78854), .Z(n78859) );
  XOR U93661 ( .A(n78857), .B(n78859), .Z(n76793) );
  XOR U93662 ( .A(n76792), .B(n76793), .Z(n78871) );
  IV U93663 ( .A(n73454), .Z(n73456) );
  NOR U93664 ( .A(n73456), .B(n73455), .Z(n78869) );
  XOR U93665 ( .A(n78871), .B(n78869), .Z(n78882) );
  IV U93666 ( .A(n78882), .Z(n73464) );
  IV U93667 ( .A(n73457), .Z(n73458) );
  NOR U93668 ( .A(n73459), .B(n73458), .Z(n78880) );
  IV U93669 ( .A(n73460), .Z(n73462) );
  NOR U93670 ( .A(n73462), .B(n73461), .Z(n78865) );
  NOR U93671 ( .A(n78880), .B(n78865), .Z(n73463) );
  XOR U93672 ( .A(n73464), .B(n73463), .Z(n76791) );
  XOR U93673 ( .A(n76788), .B(n76791), .Z(n76782) );
  IV U93674 ( .A(n73465), .Z(n76786) );
  NOR U93675 ( .A(n73466), .B(n76786), .Z(n76780) );
  NOR U93676 ( .A(n73468), .B(n73467), .Z(n73469) );
  IV U93677 ( .A(n73469), .Z(n73470) );
  NOR U93678 ( .A(n73471), .B(n73470), .Z(n73472) );
  IV U93679 ( .A(n73472), .Z(n76775) );
  NOR U93680 ( .A(n73473), .B(n76775), .Z(n73474) );
  NOR U93681 ( .A(n76780), .B(n73474), .Z(n73475) );
  XOR U93682 ( .A(n76782), .B(n73475), .Z(n78887) );
  XOR U93683 ( .A(n78888), .B(n78887), .Z(n76768) );
  XOR U93684 ( .A(n73476), .B(n76768), .Z(n78897) );
  XOR U93685 ( .A(n78898), .B(n78897), .Z(n78901) );
  XOR U93686 ( .A(n78899), .B(n78901), .Z(n78906) );
  XOR U93687 ( .A(n78904), .B(n78906), .Z(n78908) );
  NOR U93688 ( .A(n73480), .B(n78908), .Z(n84615) );
  IV U93689 ( .A(n73477), .Z(n73479) );
  NOR U93690 ( .A(n73479), .B(n73478), .Z(n78915) );
  XOR U93691 ( .A(n78907), .B(n78908), .Z(n78916) );
  IV U93692 ( .A(n78916), .Z(n73481) );
  XOR U93693 ( .A(n78915), .B(n73481), .Z(n73483) );
  NOR U93694 ( .A(n73481), .B(n73480), .Z(n73482) );
  NOR U93695 ( .A(n73483), .B(n73482), .Z(n73484) );
  NOR U93696 ( .A(n84615), .B(n73484), .Z(n78912) );
  XOR U93697 ( .A(n73485), .B(n78912), .Z(n76764) );
  XOR U93698 ( .A(n73486), .B(n76764), .Z(n76757) );
  XOR U93699 ( .A(n73487), .B(n76757), .Z(n78930) );
  XOR U93700 ( .A(n78928), .B(n78930), .Z(n78937) );
  IV U93701 ( .A(n78937), .Z(n73495) );
  IV U93702 ( .A(n73488), .Z(n73490) );
  NOR U93703 ( .A(n73490), .B(n73489), .Z(n76755) );
  IV U93704 ( .A(n73491), .Z(n73493) );
  NOR U93705 ( .A(n73493), .B(n73492), .Z(n78936) );
  NOR U93706 ( .A(n76755), .B(n78936), .Z(n73494) );
  XOR U93707 ( .A(n73495), .B(n73494), .Z(n76754) );
  XOR U93708 ( .A(n76752), .B(n76754), .Z(n78943) );
  XOR U93709 ( .A(n78941), .B(n78943), .Z(n76751) );
  XOR U93710 ( .A(n76749), .B(n76751), .Z(n84657) );
  XOR U93711 ( .A(n73496), .B(n84657), .Z(n76748) );
  IV U93712 ( .A(n73497), .Z(n73498) );
  NOR U93713 ( .A(n73499), .B(n73498), .Z(n76746) );
  XOR U93714 ( .A(n76748), .B(n76746), .Z(n78949) );
  XOR U93715 ( .A(n78948), .B(n78949), .Z(n78953) );
  IV U93716 ( .A(n73500), .Z(n73502) );
  NOR U93717 ( .A(n73502), .B(n73501), .Z(n78951) );
  XOR U93718 ( .A(n78953), .B(n78951), .Z(n76743) );
  IV U93719 ( .A(n73503), .Z(n73504) );
  NOR U93720 ( .A(n73505), .B(n73504), .Z(n76741) );
  XOR U93721 ( .A(n76743), .B(n76741), .Z(n76736) );
  XOR U93722 ( .A(n76735), .B(n76736), .Z(n76739) );
  IV U93723 ( .A(n73506), .Z(n73507) );
  NOR U93724 ( .A(n73519), .B(n73507), .Z(n76738) );
  IV U93725 ( .A(n73508), .Z(n73509) );
  NOR U93726 ( .A(n73510), .B(n73509), .Z(n76733) );
  NOR U93727 ( .A(n76738), .B(n76733), .Z(n73511) );
  XOR U93728 ( .A(n76739), .B(n73511), .Z(n73520) );
  IV U93729 ( .A(n73520), .Z(n73516) );
  IV U93730 ( .A(n73512), .Z(n73513) );
  NOR U93731 ( .A(n73514), .B(n73513), .Z(n73524) );
  IV U93732 ( .A(n73524), .Z(n73515) );
  NOR U93733 ( .A(n73516), .B(n73515), .Z(n82373) );
  IV U93734 ( .A(n73517), .Z(n73518) );
  NOR U93735 ( .A(n73519), .B(n73518), .Z(n73521) );
  NOR U93736 ( .A(n73520), .B(n73521), .Z(n73523) );
  IV U93737 ( .A(n73521), .Z(n73522) );
  NOR U93738 ( .A(n76739), .B(n73522), .Z(n82375) );
  NOR U93739 ( .A(n73523), .B(n82375), .Z(n78958) );
  NOR U93740 ( .A(n73524), .B(n78958), .Z(n73525) );
  NOR U93741 ( .A(n82373), .B(n73525), .Z(n78963) );
  XOR U93742 ( .A(n73526), .B(n78963), .Z(n76732) );
  XOR U93743 ( .A(n73527), .B(n76732), .Z(n76722) );
  XOR U93744 ( .A(n76723), .B(n76722), .Z(n76726) );
  XOR U93745 ( .A(n73528), .B(n76726), .Z(n76716) );
  XOR U93746 ( .A(n76719), .B(n76716), .Z(n76713) );
  IV U93747 ( .A(n73529), .Z(n73531) );
  NOR U93748 ( .A(n73531), .B(n73530), .Z(n76715) );
  IV U93749 ( .A(n73543), .Z(n73532) );
  NOR U93750 ( .A(n73532), .B(n73542), .Z(n76712) );
  NOR U93751 ( .A(n76715), .B(n76712), .Z(n73533) );
  XOR U93752 ( .A(n76713), .B(n73533), .Z(n76706) );
  IV U93753 ( .A(n73534), .Z(n73535) );
  NOR U93754 ( .A(n73535), .B(n73542), .Z(n76709) );
  IV U93755 ( .A(n73536), .Z(n73539) );
  IV U93756 ( .A(n73537), .Z(n73538) );
  NOR U93757 ( .A(n73539), .B(n73538), .Z(n76707) );
  NOR U93758 ( .A(n76709), .B(n76707), .Z(n73540) );
  XOR U93759 ( .A(n76706), .B(n73540), .Z(n78971) );
  IV U93760 ( .A(n73541), .Z(n73547) );
  XOR U93761 ( .A(n73543), .B(n73542), .Z(n73544) );
  NOR U93762 ( .A(n73545), .B(n73544), .Z(n73546) );
  IV U93763 ( .A(n73546), .Z(n73552) );
  NOR U93764 ( .A(n73547), .B(n73552), .Z(n78969) );
  XOR U93765 ( .A(n78971), .B(n78969), .Z(n78976) );
  IV U93766 ( .A(n73548), .Z(n73549) );
  NOR U93767 ( .A(n73550), .B(n73549), .Z(n78975) );
  IV U93768 ( .A(n73551), .Z(n73553) );
  NOR U93769 ( .A(n73553), .B(n73552), .Z(n78972) );
  NOR U93770 ( .A(n78975), .B(n78972), .Z(n73554) );
  XOR U93771 ( .A(n78976), .B(n73554), .Z(n73555) );
  IV U93772 ( .A(n73555), .Z(n76704) );
  XOR U93773 ( .A(n76702), .B(n76704), .Z(n78980) );
  XOR U93774 ( .A(n73556), .B(n78980), .Z(n76692) );
  XOR U93775 ( .A(n73557), .B(n76692), .Z(n78991) );
  XOR U93776 ( .A(n78988), .B(n78991), .Z(n73558) );
  NOR U93777 ( .A(n73559), .B(n73558), .Z(n82323) );
  IV U93778 ( .A(n73560), .Z(n73561) );
  NOR U93779 ( .A(n73562), .B(n73561), .Z(n78990) );
  NOR U93780 ( .A(n78990), .B(n78988), .Z(n73563) );
  XOR U93781 ( .A(n78991), .B(n73563), .Z(n73564) );
  NOR U93782 ( .A(n73565), .B(n73564), .Z(n73566) );
  NOR U93783 ( .A(n82323), .B(n73566), .Z(n78996) );
  IV U93784 ( .A(n73567), .Z(n73569) );
  NOR U93785 ( .A(n73569), .B(n73568), .Z(n73570) );
  IV U93786 ( .A(n73570), .Z(n78998) );
  XOR U93787 ( .A(n78996), .B(n78998), .Z(n79001) );
  XOR U93788 ( .A(n79000), .B(n79001), .Z(n79004) );
  XOR U93789 ( .A(n79003), .B(n79004), .Z(n82319) );
  XOR U93790 ( .A(n76691), .B(n82319), .Z(n73571) );
  IV U93791 ( .A(n73571), .Z(n76687) );
  IV U93792 ( .A(n73572), .Z(n73574) );
  IV U93793 ( .A(n73573), .Z(n82313) );
  NOR U93794 ( .A(n73574), .B(n82313), .Z(n76685) );
  XOR U93795 ( .A(n76687), .B(n76685), .Z(n76689) );
  IV U93796 ( .A(n73575), .Z(n73576) );
  NOR U93797 ( .A(n73577), .B(n73576), .Z(n76688) );
  IV U93798 ( .A(n73578), .Z(n73580) );
  NOR U93799 ( .A(n73580), .B(n73579), .Z(n76682) );
  NOR U93800 ( .A(n76688), .B(n76682), .Z(n73581) );
  XOR U93801 ( .A(n76689), .B(n73581), .Z(n76677) );
  XOR U93802 ( .A(n73582), .B(n76677), .Z(n76674) );
  XOR U93803 ( .A(n76675), .B(n76674), .Z(n73586) );
  NOR U93804 ( .A(n73583), .B(n73586), .Z(n73592) );
  IV U93805 ( .A(n73584), .Z(n73585) );
  NOR U93806 ( .A(n73585), .B(n76674), .Z(n84740) );
  NOR U93807 ( .A(n73587), .B(n73586), .Z(n73590) );
  IV U93808 ( .A(n73588), .Z(n73589) );
  NOR U93809 ( .A(n73590), .B(n73589), .Z(n84743) );
  NOR U93810 ( .A(n84740), .B(n84743), .Z(n73591) );
  IV U93811 ( .A(n73591), .Z(n79008) );
  NOR U93812 ( .A(n73592), .B(n79008), .Z(n76672) );
  XOR U93813 ( .A(n73593), .B(n76672), .Z(n82303) );
  IV U93814 ( .A(n82303), .Z(n73600) );
  IV U93815 ( .A(n73594), .Z(n73595) );
  NOR U93816 ( .A(n73596), .B(n73595), .Z(n82302) );
  IV U93817 ( .A(n73597), .Z(n73599) );
  NOR U93818 ( .A(n73599), .B(n73598), .Z(n84752) );
  NOR U93819 ( .A(n82302), .B(n84752), .Z(n76670) );
  XOR U93820 ( .A(n73600), .B(n76670), .Z(n76666) );
  XOR U93821 ( .A(n76664), .B(n76666), .Z(n76668) );
  XOR U93822 ( .A(n73601), .B(n76668), .Z(n76651) );
  IV U93823 ( .A(n73602), .Z(n73604) );
  NOR U93824 ( .A(n73604), .B(n73603), .Z(n76660) );
  IV U93825 ( .A(n73605), .Z(n73606) );
  NOR U93826 ( .A(n73606), .B(n73608), .Z(n84771) );
  IV U93827 ( .A(n73607), .Z(n73609) );
  NOR U93828 ( .A(n73609), .B(n73608), .Z(n84776) );
  NOR U93829 ( .A(n84771), .B(n84776), .Z(n76652) );
  IV U93830 ( .A(n76652), .Z(n73610) );
  NOR U93831 ( .A(n76660), .B(n73610), .Z(n73611) );
  XOR U93832 ( .A(n76651), .B(n73611), .Z(n76655) );
  IV U93833 ( .A(n73612), .Z(n73614) );
  NOR U93834 ( .A(n73614), .B(n73613), .Z(n76653) );
  IV U93835 ( .A(n73615), .Z(n73616) );
  NOR U93836 ( .A(n76638), .B(n73616), .Z(n76649) );
  NOR U93837 ( .A(n76653), .B(n76649), .Z(n73617) );
  XOR U93838 ( .A(n76655), .B(n73617), .Z(n73618) );
  IV U93839 ( .A(n73618), .Z(n76645) );
  IV U93840 ( .A(n73619), .Z(n73620) );
  NOR U93841 ( .A(n73620), .B(n73624), .Z(n76643) );
  XOR U93842 ( .A(n76645), .B(n76643), .Z(n76633) );
  IV U93843 ( .A(n73621), .Z(n73622) );
  NOR U93844 ( .A(n79022), .B(n73622), .Z(n76629) );
  IV U93845 ( .A(n73623), .Z(n73625) );
  NOR U93846 ( .A(n73625), .B(n73624), .Z(n76631) );
  NOR U93847 ( .A(n76629), .B(n76631), .Z(n73626) );
  XOR U93848 ( .A(n76633), .B(n73626), .Z(n73627) );
  IV U93849 ( .A(n73627), .Z(n79021) );
  NOR U93850 ( .A(n73629), .B(n73628), .Z(n76624) );
  IV U93851 ( .A(n73630), .Z(n73632) );
  NOR U93852 ( .A(n73632), .B(n73631), .Z(n76621) );
  NOR U93853 ( .A(n76624), .B(n76621), .Z(n73633) );
  XOR U93854 ( .A(n79021), .B(n73633), .Z(n73634) );
  NOR U93855 ( .A(n73635), .B(n73634), .Z(n73637) );
  IV U93856 ( .A(n73635), .Z(n73636) );
  XOR U93857 ( .A(n76624), .B(n79021), .Z(n79027) );
  NOR U93858 ( .A(n73636), .B(n79027), .Z(n82280) );
  NOR U93859 ( .A(n73637), .B(n82280), .Z(n79030) );
  XOR U93860 ( .A(n73638), .B(n79030), .Z(n79035) );
  XOR U93861 ( .A(n79033), .B(n79035), .Z(n79041) );
  IV U93862 ( .A(n73639), .Z(n73640) );
  NOR U93863 ( .A(n73641), .B(n73640), .Z(n79040) );
  NOR U93864 ( .A(n79036), .B(n79040), .Z(n73642) );
  XOR U93865 ( .A(n79041), .B(n73642), .Z(n76614) );
  IV U93866 ( .A(n73643), .Z(n73645) );
  NOR U93867 ( .A(n73645), .B(n73644), .Z(n76617) );
  IV U93868 ( .A(n73646), .Z(n73648) );
  NOR U93869 ( .A(n73648), .B(n73647), .Z(n76615) );
  NOR U93870 ( .A(n76617), .B(n76615), .Z(n73649) );
  XOR U93871 ( .A(n76614), .B(n73649), .Z(n79046) );
  XOR U93872 ( .A(n79045), .B(n79046), .Z(n76610) );
  NOR U93873 ( .A(n73650), .B(n76611), .Z(n73654) );
  IV U93874 ( .A(n73651), .Z(n73653) );
  NOR U93875 ( .A(n73653), .B(n73652), .Z(n76607) );
  NOR U93876 ( .A(n73654), .B(n76607), .Z(n73655) );
  XOR U93877 ( .A(n76610), .B(n73655), .Z(n76605) );
  IV U93878 ( .A(n73656), .Z(n73657) );
  NOR U93879 ( .A(n73658), .B(n73657), .Z(n84822) );
  IV U93880 ( .A(n73659), .Z(n73660) );
  NOR U93881 ( .A(n73661), .B(n73660), .Z(n84832) );
  NOR U93882 ( .A(n84822), .B(n84832), .Z(n76606) );
  XOR U93883 ( .A(n76605), .B(n76606), .Z(n76600) );
  XOR U93884 ( .A(n76599), .B(n76600), .Z(n76603) );
  XOR U93885 ( .A(n76602), .B(n76603), .Z(n76594) );
  XOR U93886 ( .A(n76593), .B(n76594), .Z(n76597) );
  IV U93887 ( .A(n73662), .Z(n73663) );
  NOR U93888 ( .A(n73664), .B(n73663), .Z(n76596) );
  IV U93889 ( .A(n73665), .Z(n73667) );
  NOR U93890 ( .A(n73667), .B(n73666), .Z(n76587) );
  NOR U93891 ( .A(n76596), .B(n76587), .Z(n73668) );
  XOR U93892 ( .A(n76597), .B(n73668), .Z(n73669) );
  IV U93893 ( .A(n73669), .Z(n76591) );
  XOR U93894 ( .A(n76589), .B(n76591), .Z(n79064) );
  XOR U93895 ( .A(n79062), .B(n79064), .Z(n76585) );
  XOR U93896 ( .A(n73670), .B(n76585), .Z(n79068) );
  XOR U93897 ( .A(n79066), .B(n79068), .Z(n79073) );
  XOR U93898 ( .A(n79069), .B(n79073), .Z(n76582) );
  IV U93899 ( .A(n73671), .Z(n73672) );
  NOR U93900 ( .A(n73673), .B(n73672), .Z(n79072) );
  IV U93901 ( .A(n73674), .Z(n73676) );
  NOR U93902 ( .A(n73676), .B(n73675), .Z(n76581) );
  NOR U93903 ( .A(n79072), .B(n76581), .Z(n73677) );
  XOR U93904 ( .A(n76582), .B(n73677), .Z(n73678) );
  IV U93905 ( .A(n73678), .Z(n79078) );
  IV U93906 ( .A(n73679), .Z(n73681) );
  NOR U93907 ( .A(n73681), .B(n73680), .Z(n79076) );
  XOR U93908 ( .A(n79078), .B(n79076), .Z(n79081) );
  XOR U93909 ( .A(n79079), .B(n79081), .Z(n76579) );
  XOR U93910 ( .A(n76578), .B(n76579), .Z(n79089) );
  XOR U93911 ( .A(n79087), .B(n79089), .Z(n79094) );
  XOR U93912 ( .A(n73682), .B(n79094), .Z(n73683) );
  IV U93913 ( .A(n73683), .Z(n79097) );
  XOR U93914 ( .A(n79096), .B(n79097), .Z(n79102) );
  XOR U93915 ( .A(n79101), .B(n79102), .Z(n84889) );
  XOR U93916 ( .A(n79104), .B(n84889), .Z(n73689) );
  IV U93917 ( .A(n73689), .Z(n73684) );
  NOR U93918 ( .A(n73688), .B(n73684), .Z(n73685) );
  IV U93919 ( .A(n73685), .Z(n73687) );
  NOR U93920 ( .A(n73686), .B(n84893), .Z(n73691) );
  NOR U93921 ( .A(n73687), .B(n73691), .Z(n73695) );
  IV U93922 ( .A(n73688), .Z(n73690) );
  NOR U93923 ( .A(n73690), .B(n73689), .Z(n82219) );
  IV U93924 ( .A(n73691), .Z(n73692) );
  NOR U93925 ( .A(n73692), .B(n84889), .Z(n73693) );
  NOR U93926 ( .A(n82219), .B(n73693), .Z(n73694) );
  IV U93927 ( .A(n73694), .Z(n79112) );
  NOR U93928 ( .A(n73695), .B(n79112), .Z(n73696) );
  IV U93929 ( .A(n73696), .Z(n79108) );
  NOR U93930 ( .A(n73703), .B(n79108), .Z(n82215) );
  IV U93931 ( .A(n73697), .Z(n73698) );
  NOR U93932 ( .A(n73699), .B(n73698), .Z(n76575) );
  IV U93933 ( .A(n73700), .Z(n73702) );
  NOR U93934 ( .A(n73702), .B(n73701), .Z(n79107) );
  XOR U93935 ( .A(n79107), .B(n79108), .Z(n76576) );
  IV U93936 ( .A(n76576), .Z(n73704) );
  XOR U93937 ( .A(n76575), .B(n73704), .Z(n73706) );
  NOR U93938 ( .A(n73704), .B(n73703), .Z(n73705) );
  NOR U93939 ( .A(n73706), .B(n73705), .Z(n73707) );
  NOR U93940 ( .A(n82215), .B(n73707), .Z(n79114) );
  XOR U93941 ( .A(n79115), .B(n79114), .Z(n76574) );
  XOR U93942 ( .A(n73708), .B(n76574), .Z(n76568) );
  XOR U93943 ( .A(n76566), .B(n76568), .Z(n76571) );
  IV U93944 ( .A(n73709), .Z(n73713) );
  NOR U93945 ( .A(n73711), .B(n73710), .Z(n73712) );
  IV U93946 ( .A(n73712), .Z(n73715) );
  NOR U93947 ( .A(n73713), .B(n73715), .Z(n76569) );
  XOR U93948 ( .A(n76571), .B(n76569), .Z(n79127) );
  IV U93949 ( .A(n73714), .Z(n73716) );
  NOR U93950 ( .A(n73716), .B(n73715), .Z(n79125) );
  XOR U93951 ( .A(n79127), .B(n79125), .Z(n82195) );
  IV U93952 ( .A(n73717), .Z(n73718) );
  NOR U93953 ( .A(n73719), .B(n73718), .Z(n82198) );
  IV U93954 ( .A(n73720), .Z(n73721) );
  NOR U93955 ( .A(n73722), .B(n73721), .Z(n82194) );
  NOR U93956 ( .A(n82198), .B(n82194), .Z(n79128) );
  XOR U93957 ( .A(n82195), .B(n79128), .Z(n79131) );
  XOR U93958 ( .A(n79132), .B(n79131), .Z(n82186) );
  IV U93959 ( .A(n82186), .Z(n73732) );
  IV U93960 ( .A(n73723), .Z(n73724) );
  NOR U93961 ( .A(n73730), .B(n73724), .Z(n76563) );
  IV U93962 ( .A(n73725), .Z(n73726) );
  NOR U93963 ( .A(n73727), .B(n73726), .Z(n84930) );
  IV U93964 ( .A(n73728), .Z(n73729) );
  NOR U93965 ( .A(n73730), .B(n73729), .Z(n82184) );
  NOR U93966 ( .A(n84930), .B(n82184), .Z(n79133) );
  IV U93967 ( .A(n79133), .Z(n76562) );
  NOR U93968 ( .A(n76563), .B(n76562), .Z(n73731) );
  XOR U93969 ( .A(n73732), .B(n73731), .Z(n79145) );
  XOR U93970 ( .A(n73733), .B(n79145), .Z(n79141) );
  XOR U93971 ( .A(n73734), .B(n79141), .Z(n76554) );
  XOR U93972 ( .A(n73735), .B(n76554), .Z(n76547) );
  XOR U93973 ( .A(n73736), .B(n76547), .Z(n76544) );
  XOR U93974 ( .A(n76543), .B(n76544), .Z(n79158) );
  XOR U93975 ( .A(n79157), .B(n79158), .Z(n79153) );
  IV U93976 ( .A(n73737), .Z(n73738) );
  NOR U93977 ( .A(n73739), .B(n73738), .Z(n79152) );
  IV U93978 ( .A(n73740), .Z(n73742) );
  NOR U93979 ( .A(n73742), .B(n73741), .Z(n76538) );
  NOR U93980 ( .A(n79152), .B(n76538), .Z(n73743) );
  XOR U93981 ( .A(n79153), .B(n73743), .Z(n73744) );
  IV U93982 ( .A(n73744), .Z(n76542) );
  IV U93983 ( .A(n73745), .Z(n73746) );
  NOR U93984 ( .A(n73747), .B(n73746), .Z(n76540) );
  NOR U93985 ( .A(n73748), .B(n76535), .Z(n73749) );
  NOR U93986 ( .A(n76540), .B(n73749), .Z(n73750) );
  XOR U93987 ( .A(n76542), .B(n73750), .Z(n79165) );
  IV U93988 ( .A(n73751), .Z(n73752) );
  NOR U93989 ( .A(n73753), .B(n73752), .Z(n79164) );
  IV U93990 ( .A(n73754), .Z(n73756) );
  NOR U93991 ( .A(n73756), .B(n73755), .Z(n79171) );
  NOR U93992 ( .A(n79164), .B(n79171), .Z(n73757) );
  XOR U93993 ( .A(n79165), .B(n73757), .Z(n79176) );
  XOR U93994 ( .A(n79174), .B(n79176), .Z(n82159) );
  XOR U93995 ( .A(n76533), .B(n82159), .Z(n79182) );
  IV U93996 ( .A(n73758), .Z(n73760) );
  NOR U93997 ( .A(n73760), .B(n73759), .Z(n79181) );
  IV U93998 ( .A(n73761), .Z(n73762) );
  NOR U93999 ( .A(n73762), .B(n73766), .Z(n79187) );
  NOR U94000 ( .A(n79181), .B(n79187), .Z(n73763) );
  XOR U94001 ( .A(n79182), .B(n73763), .Z(n79196) );
  IV U94002 ( .A(n73764), .Z(n73765) );
  NOR U94003 ( .A(n73766), .B(n73765), .Z(n76531) );
  XOR U94004 ( .A(n79196), .B(n76531), .Z(n73767) );
  NOR U94005 ( .A(n73768), .B(n73767), .Z(n85024) );
  IV U94006 ( .A(n73769), .Z(n73771) );
  NOR U94007 ( .A(n73771), .B(n73770), .Z(n79194) );
  NOR U94008 ( .A(n79194), .B(n76531), .Z(n73772) );
  XOR U94009 ( .A(n79196), .B(n73772), .Z(n73773) );
  NOR U94010 ( .A(n73774), .B(n73773), .Z(n73775) );
  NOR U94011 ( .A(n85024), .B(n73775), .Z(n73776) );
  IV U94012 ( .A(n73776), .Z(n76527) );
  XOR U94013 ( .A(n76526), .B(n76527), .Z(n79200) );
  IV U94014 ( .A(n73777), .Z(n73778) );
  NOR U94015 ( .A(n73779), .B(n73778), .Z(n76529) );
  IV U94016 ( .A(n73780), .Z(n73782) );
  IV U94017 ( .A(n73781), .Z(n73788) );
  NOR U94018 ( .A(n73782), .B(n73788), .Z(n79198) );
  NOR U94019 ( .A(n76529), .B(n79198), .Z(n73783) );
  XOR U94020 ( .A(n79200), .B(n73783), .Z(n76522) );
  IV U94021 ( .A(n73784), .Z(n73785) );
  NOR U94022 ( .A(n73786), .B(n73785), .Z(n76523) );
  IV U94023 ( .A(n73787), .Z(n73789) );
  NOR U94024 ( .A(n73789), .B(n73788), .Z(n79204) );
  NOR U94025 ( .A(n76523), .B(n79204), .Z(n73790) );
  XOR U94026 ( .A(n76522), .B(n73790), .Z(n79208) );
  XOR U94027 ( .A(n79207), .B(n79208), .Z(n76519) );
  IV U94028 ( .A(n73791), .Z(n73793) );
  NOR U94029 ( .A(n73793), .B(n73792), .Z(n76518) );
  IV U94030 ( .A(n73794), .Z(n73796) );
  NOR U94031 ( .A(n73796), .B(n73795), .Z(n76513) );
  NOR U94032 ( .A(n76518), .B(n76513), .Z(n73797) );
  XOR U94033 ( .A(n76519), .B(n73797), .Z(n76510) );
  XOR U94034 ( .A(n73798), .B(n76510), .Z(n76507) );
  IV U94035 ( .A(n73799), .Z(n73800) );
  NOR U94036 ( .A(n73801), .B(n73800), .Z(n76505) );
  XOR U94037 ( .A(n76507), .B(n76505), .Z(n82137) );
  IV U94038 ( .A(n73802), .Z(n73804) );
  NOR U94039 ( .A(n73804), .B(n73803), .Z(n82136) );
  IV U94040 ( .A(n73805), .Z(n73807) );
  NOR U94041 ( .A(n73807), .B(n73806), .Z(n85062) );
  NOR U94042 ( .A(n82136), .B(n85062), .Z(n76508) );
  XOR U94043 ( .A(n82137), .B(n76508), .Z(n73808) );
  IV U94044 ( .A(n73808), .Z(n79217) );
  XOR U94045 ( .A(n76503), .B(n79217), .Z(n79221) );
  XOR U94046 ( .A(n73809), .B(n79221), .Z(n73810) );
  IV U94047 ( .A(n73810), .Z(n79224) );
  XOR U94048 ( .A(n79222), .B(n79224), .Z(n79226) );
  XOR U94049 ( .A(n79225), .B(n79226), .Z(n76501) );
  IV U94050 ( .A(n73811), .Z(n73812) );
  NOR U94051 ( .A(n73813), .B(n73812), .Z(n76500) );
  IV U94052 ( .A(n73814), .Z(n73815) );
  NOR U94053 ( .A(n73816), .B(n73815), .Z(n76498) );
  NOR U94054 ( .A(n76500), .B(n76498), .Z(n73817) );
  XOR U94055 ( .A(n76501), .B(n73817), .Z(n73826) );
  IV U94056 ( .A(n73826), .Z(n73821) );
  IV U94057 ( .A(n73818), .Z(n73819) );
  NOR U94058 ( .A(n73819), .B(n73833), .Z(n73830) );
  IV U94059 ( .A(n73830), .Z(n73820) );
  NOR U94060 ( .A(n73821), .B(n73820), .Z(n79234) );
  IV U94061 ( .A(n73822), .Z(n73823) );
  NOR U94062 ( .A(n73833), .B(n73823), .Z(n73827) );
  IV U94063 ( .A(n73827), .Z(n73825) );
  XOR U94064 ( .A(n76500), .B(n76501), .Z(n73824) );
  NOR U94065 ( .A(n73825), .B(n73824), .Z(n76497) );
  NOR U94066 ( .A(n73827), .B(n73826), .Z(n73828) );
  NOR U94067 ( .A(n76497), .B(n73828), .Z(n73829) );
  NOR U94068 ( .A(n73830), .B(n73829), .Z(n73831) );
  NOR U94069 ( .A(n79234), .B(n73831), .Z(n76494) );
  IV U94070 ( .A(n73832), .Z(n73834) );
  NOR U94071 ( .A(n73834), .B(n73833), .Z(n73835) );
  IV U94072 ( .A(n73835), .Z(n73836) );
  NOR U94073 ( .A(n73837), .B(n73836), .Z(n73838) );
  IV U94074 ( .A(n73838), .Z(n76495) );
  XOR U94075 ( .A(n76494), .B(n76495), .Z(n76488) );
  XOR U94076 ( .A(n73839), .B(n76488), .Z(n76490) );
  IV U94077 ( .A(n73840), .Z(n73842) );
  NOR U94078 ( .A(n73842), .B(n73841), .Z(n82118) );
  NOR U94079 ( .A(n82118), .B(n82113), .Z(n76491) );
  XOR U94080 ( .A(n76490), .B(n76491), .Z(n76480) );
  XOR U94081 ( .A(n76479), .B(n76480), .Z(n76483) );
  XOR U94082 ( .A(n73843), .B(n76483), .Z(n76474) );
  IV U94083 ( .A(n73844), .Z(n73845) );
  NOR U94084 ( .A(n73846), .B(n73845), .Z(n76475) );
  IV U94085 ( .A(n73847), .Z(n73849) );
  NOR U94086 ( .A(n73849), .B(n73848), .Z(n79241) );
  NOR U94087 ( .A(n76475), .B(n79241), .Z(n73850) );
  XOR U94088 ( .A(n76474), .B(n73850), .Z(n76472) );
  IV U94089 ( .A(n73851), .Z(n73854) );
  NOR U94090 ( .A(n73852), .B(n73856), .Z(n73853) );
  IV U94091 ( .A(n73853), .Z(n73865) );
  NOR U94092 ( .A(n73854), .B(n73865), .Z(n73868) );
  IV U94093 ( .A(n73868), .Z(n73855) );
  NOR U94094 ( .A(n76472), .B(n73855), .Z(n82089) );
  NOR U94095 ( .A(n73857), .B(n73856), .Z(n73858) );
  IV U94096 ( .A(n73858), .Z(n79246) );
  NOR U94097 ( .A(n73859), .B(n79246), .Z(n73871) );
  NOR U94098 ( .A(n82089), .B(n73871), .Z(n73860) );
  IV U94099 ( .A(n73860), .Z(n73870) );
  IV U94100 ( .A(n73861), .Z(n73862) );
  NOR U94101 ( .A(n73863), .B(n73862), .Z(n76471) );
  IV U94102 ( .A(n73864), .Z(n73866) );
  NOR U94103 ( .A(n73866), .B(n73865), .Z(n76469) );
  NOR U94104 ( .A(n76471), .B(n76469), .Z(n73867) );
  XOR U94105 ( .A(n73867), .B(n76472), .Z(n79245) );
  NOR U94106 ( .A(n73868), .B(n79245), .Z(n73869) );
  NOR U94107 ( .A(n73870), .B(n73869), .Z(n73874) );
  IV U94108 ( .A(n73871), .Z(n73872) );
  NOR U94109 ( .A(n79245), .B(n73872), .Z(n73873) );
  NOR U94110 ( .A(n73874), .B(n73873), .Z(n79264) );
  IV U94111 ( .A(n73875), .Z(n79255) );
  NOR U94112 ( .A(n73876), .B(n79255), .Z(n73879) );
  IV U94113 ( .A(n73877), .Z(n73878) );
  NOR U94114 ( .A(n73878), .B(n73882), .Z(n79262) );
  NOR U94115 ( .A(n73879), .B(n79262), .Z(n73880) );
  XOR U94116 ( .A(n79264), .B(n73880), .Z(n76464) );
  IV U94117 ( .A(n73881), .Z(n73883) );
  NOR U94118 ( .A(n73883), .B(n73882), .Z(n76466) );
  NOR U94119 ( .A(n76463), .B(n76466), .Z(n73884) );
  XOR U94120 ( .A(n76464), .B(n73884), .Z(n79267) );
  XOR U94121 ( .A(n79265), .B(n79267), .Z(n76461) );
  XOR U94122 ( .A(n73885), .B(n76461), .Z(n73886) );
  IV U94123 ( .A(n73886), .Z(n79283) );
  IV U94124 ( .A(n73887), .Z(n73888) );
  NOR U94125 ( .A(n73889), .B(n73888), .Z(n79282) );
  NOR U94126 ( .A(n73890), .B(n76454), .Z(n73891) );
  NOR U94127 ( .A(n79282), .B(n73891), .Z(n73892) );
  XOR U94128 ( .A(n79283), .B(n73892), .Z(n76448) );
  IV U94129 ( .A(n73893), .Z(n73895) );
  NOR U94130 ( .A(n73895), .B(n73894), .Z(n85109) );
  IV U94131 ( .A(n73896), .Z(n73897) );
  NOR U94132 ( .A(n73898), .B(n73897), .Z(n82055) );
  NOR U94133 ( .A(n85109), .B(n82055), .Z(n76446) );
  XOR U94134 ( .A(n76448), .B(n76446), .Z(n76440) );
  XOR U94135 ( .A(n76439), .B(n76440), .Z(n82043) );
  XOR U94136 ( .A(n76442), .B(n82043), .Z(n76430) );
  IV U94137 ( .A(n73899), .Z(n76433) );
  NOR U94138 ( .A(n73900), .B(n76433), .Z(n73904) );
  IV U94139 ( .A(n73901), .Z(n73903) );
  NOR U94140 ( .A(n73903), .B(n73902), .Z(n76429) );
  NOR U94141 ( .A(n73904), .B(n76429), .Z(n73905) );
  XOR U94142 ( .A(n76430), .B(n73905), .Z(n76427) );
  NOR U94143 ( .A(n73907), .B(n73906), .Z(n73908) );
  NOR U94144 ( .A(n82026), .B(n73908), .Z(n73909) );
  NOR U94145 ( .A(n73909), .B(n82020), .Z(n73910) );
  IV U94146 ( .A(n73910), .Z(n76428) );
  XOR U94147 ( .A(n76427), .B(n76428), .Z(n76422) );
  XOR U94148 ( .A(n76420), .B(n76422), .Z(n76424) );
  XOR U94149 ( .A(n73911), .B(n76424), .Z(n76416) );
  IV U94150 ( .A(n73912), .Z(n73914) );
  NOR U94151 ( .A(n73914), .B(n73913), .Z(n76415) );
  IV U94152 ( .A(n73915), .Z(n73916) );
  NOR U94153 ( .A(n73917), .B(n73916), .Z(n79294) );
  NOR U94154 ( .A(n76415), .B(n79294), .Z(n73918) );
  XOR U94155 ( .A(n76416), .B(n73918), .Z(n79304) );
  XOR U94156 ( .A(n73919), .B(n79304), .Z(n73924) );
  NOR U94157 ( .A(n73920), .B(n73924), .Z(n85152) );
  IV U94158 ( .A(n73921), .Z(n73922) );
  NOR U94159 ( .A(n73922), .B(n79305), .Z(n73925) );
  IV U94160 ( .A(n73925), .Z(n73923) );
  NOR U94161 ( .A(n79304), .B(n73923), .Z(n85148) );
  IV U94162 ( .A(n73924), .Z(n73926) );
  NOR U94163 ( .A(n73926), .B(n73925), .Z(n73927) );
  NOR U94164 ( .A(n85148), .B(n73927), .Z(n76412) );
  NOR U94165 ( .A(n73928), .B(n76412), .Z(n73929) );
  NOR U94166 ( .A(n85152), .B(n73929), .Z(n76408) );
  XOR U94167 ( .A(n73930), .B(n76408), .Z(n76406) );
  XOR U94168 ( .A(n73931), .B(n76406), .Z(n73932) );
  IV U94169 ( .A(n73932), .Z(n79310) );
  XOR U94170 ( .A(n79311), .B(n79310), .Z(n79322) );
  IV U94171 ( .A(n73933), .Z(n73935) );
  NOR U94172 ( .A(n73935), .B(n73934), .Z(n76398) );
  IV U94173 ( .A(n73936), .Z(n73938) );
  NOR U94174 ( .A(n73938), .B(n73937), .Z(n79321) );
  NOR U94175 ( .A(n76398), .B(n79321), .Z(n73939) );
  XOR U94176 ( .A(n79322), .B(n73939), .Z(n76397) );
  XOR U94177 ( .A(n73940), .B(n76397), .Z(n73948) );
  IV U94178 ( .A(n73948), .Z(n73941) );
  NOR U94179 ( .A(n73942), .B(n73941), .Z(n81986) );
  IV U94180 ( .A(n73943), .Z(n73945) );
  NOR U94181 ( .A(n73945), .B(n73944), .Z(n73949) );
  IV U94182 ( .A(n73949), .Z(n73947) );
  XOR U94183 ( .A(n76395), .B(n76397), .Z(n73946) );
  NOR U94184 ( .A(n73947), .B(n73946), .Z(n76392) );
  NOR U94185 ( .A(n73949), .B(n73948), .Z(n73950) );
  NOR U94186 ( .A(n76392), .B(n73950), .Z(n73951) );
  NOR U94187 ( .A(n73952), .B(n73951), .Z(n73953) );
  NOR U94188 ( .A(n81986), .B(n73953), .Z(n73954) );
  IV U94189 ( .A(n73954), .Z(n79331) );
  XOR U94190 ( .A(n79326), .B(n79331), .Z(n81977) );
  IV U94191 ( .A(n73955), .Z(n73957) );
  NOR U94192 ( .A(n73957), .B(n73956), .Z(n79329) );
  IV U94193 ( .A(n73958), .Z(n73959) );
  NOR U94194 ( .A(n73960), .B(n73959), .Z(n79335) );
  NOR U94195 ( .A(n79329), .B(n79335), .Z(n81978) );
  XOR U94196 ( .A(n81977), .B(n81978), .Z(n79333) );
  XOR U94197 ( .A(n79334), .B(n79333), .Z(n81963) );
  IV U94198 ( .A(n73961), .Z(n73963) );
  NOR U94199 ( .A(n73963), .B(n73962), .Z(n81966) );
  IV U94200 ( .A(n73964), .Z(n73966) );
  NOR U94201 ( .A(n73966), .B(n73965), .Z(n81961) );
  NOR U94202 ( .A(n81966), .B(n81961), .Z(n76387) );
  XOR U94203 ( .A(n81963), .B(n76387), .Z(n76385) );
  XOR U94204 ( .A(n73967), .B(n76385), .Z(n81944) );
  IV U94205 ( .A(n73968), .Z(n73970) );
  NOR U94206 ( .A(n73970), .B(n73969), .Z(n81953) );
  NOR U94207 ( .A(n73971), .B(n81946), .Z(n73972) );
  NOR U94208 ( .A(n81953), .B(n73972), .Z(n79341) );
  XOR U94209 ( .A(n81944), .B(n79341), .Z(n73973) );
  IV U94210 ( .A(n73973), .Z(n79343) );
  XOR U94211 ( .A(n79342), .B(n79343), .Z(n79348) );
  XOR U94212 ( .A(n79349), .B(n79348), .Z(n73986) );
  IV U94213 ( .A(n73986), .Z(n73974) );
  NOR U94214 ( .A(n73975), .B(n73974), .Z(n73981) );
  IV U94215 ( .A(n73976), .Z(n73977) );
  NOR U94216 ( .A(n73978), .B(n73977), .Z(n73982) );
  IV U94217 ( .A(n73982), .Z(n73979) );
  NOR U94218 ( .A(n73979), .B(n79348), .Z(n73980) );
  NOR U94219 ( .A(n73981), .B(n73980), .Z(n79347) );
  IV U94220 ( .A(n79347), .Z(n79356) );
  NOR U94221 ( .A(n73983), .B(n73982), .Z(n73984) );
  IV U94222 ( .A(n73984), .Z(n73985) );
  NOR U94223 ( .A(n73986), .B(n73985), .Z(n73987) );
  NOR U94224 ( .A(n79356), .B(n73987), .Z(n76376) );
  IV U94225 ( .A(n73988), .Z(n73990) );
  NOR U94226 ( .A(n73990), .B(n73989), .Z(n73991) );
  IV U94227 ( .A(n73991), .Z(n76377) );
  XOR U94228 ( .A(n76376), .B(n76377), .Z(n76380) );
  XOR U94229 ( .A(n76379), .B(n76380), .Z(n90894) );
  NOR U94230 ( .A(n73998), .B(n90894), .Z(n81938) );
  IV U94231 ( .A(n73992), .Z(n73993) );
  NOR U94232 ( .A(n73994), .B(n73993), .Z(n76373) );
  IV U94233 ( .A(n73995), .Z(n73996) );
  NOR U94234 ( .A(n73997), .B(n73996), .Z(n79359) );
  XOR U94235 ( .A(n90894), .B(n79359), .Z(n76374) );
  IV U94236 ( .A(n76374), .Z(n73999) );
  XOR U94237 ( .A(n76373), .B(n73999), .Z(n74001) );
  NOR U94238 ( .A(n73999), .B(n73998), .Z(n74000) );
  NOR U94239 ( .A(n74001), .B(n74000), .Z(n74002) );
  NOR U94240 ( .A(n81938), .B(n74002), .Z(n74009) );
  XOR U94241 ( .A(n74003), .B(n74009), .Z(n74008) );
  IV U94242 ( .A(n74004), .Z(n74006) );
  NOR U94243 ( .A(n74006), .B(n74005), .Z(n74016) );
  IV U94244 ( .A(n74016), .Z(n74007) );
  NOR U94245 ( .A(n74008), .B(n74007), .Z(n85209) );
  IV U94246 ( .A(n74009), .Z(n76371) );
  IV U94247 ( .A(n74010), .Z(n74012) );
  NOR U94248 ( .A(n74012), .B(n74011), .Z(n76366) );
  NOR U94249 ( .A(n76366), .B(n74013), .Z(n74014) );
  XOR U94250 ( .A(n76371), .B(n74014), .Z(n74015) );
  NOR U94251 ( .A(n74016), .B(n74015), .Z(n74017) );
  NOR U94252 ( .A(n85209), .B(n74017), .Z(n74018) );
  IV U94253 ( .A(n74018), .Z(n76362) );
  NOR U94254 ( .A(n74025), .B(n76362), .Z(n76364) );
  IV U94255 ( .A(n74019), .Z(n74021) );
  NOR U94256 ( .A(n74021), .B(n74020), .Z(n76355) );
  IV U94257 ( .A(n74022), .Z(n74024) );
  NOR U94258 ( .A(n74024), .B(n74023), .Z(n76361) );
  XOR U94259 ( .A(n76361), .B(n76362), .Z(n76356) );
  IV U94260 ( .A(n76356), .Z(n74026) );
  XOR U94261 ( .A(n76355), .B(n74026), .Z(n74028) );
  NOR U94262 ( .A(n74026), .B(n74025), .Z(n74027) );
  NOR U94263 ( .A(n74028), .B(n74027), .Z(n74029) );
  NOR U94264 ( .A(n76364), .B(n74029), .Z(n76359) );
  XOR U94265 ( .A(n74030), .B(n76359), .Z(n79369) );
  XOR U94266 ( .A(n74031), .B(n79369), .Z(n81923) );
  XOR U94267 ( .A(n76352), .B(n81923), .Z(n74041) );
  IV U94268 ( .A(n74041), .Z(n74032) );
  NOR U94269 ( .A(n74040), .B(n74032), .Z(n81915) );
  IV U94270 ( .A(n74033), .Z(n74035) );
  NOR U94271 ( .A(n74035), .B(n74034), .Z(n74038) );
  IV U94272 ( .A(n74038), .Z(n74036) );
  NOR U94273 ( .A(n81923), .B(n74036), .Z(n81919) );
  NOR U94274 ( .A(n81915), .B(n81919), .Z(n74037) );
  IV U94275 ( .A(n74037), .Z(n79372) );
  NOR U94276 ( .A(n74038), .B(n74041), .Z(n74039) );
  NOR U94277 ( .A(n79372), .B(n74039), .Z(n74043) );
  NOR U94278 ( .A(n74041), .B(n74040), .Z(n74042) );
  NOR U94279 ( .A(n74043), .B(n74042), .Z(n79375) );
  XOR U94280 ( .A(n79373), .B(n79375), .Z(n79377) );
  XOR U94281 ( .A(n79376), .B(n79377), .Z(n76350) );
  XOR U94282 ( .A(n74044), .B(n76350), .Z(n76344) );
  XOR U94283 ( .A(n76345), .B(n76344), .Z(n76340) );
  XOR U94284 ( .A(n76338), .B(n76340), .Z(n79387) );
  XOR U94285 ( .A(n74045), .B(n79387), .Z(n79391) );
  XOR U94286 ( .A(n79392), .B(n79391), .Z(n76336) );
  XOR U94287 ( .A(n74046), .B(n76336), .Z(n74047) );
  IV U94288 ( .A(n74047), .Z(n76332) );
  XOR U94289 ( .A(n76330), .B(n76332), .Z(n79398) );
  IV U94290 ( .A(n74048), .Z(n74050) );
  NOR U94291 ( .A(n74050), .B(n74049), .Z(n76333) );
  IV U94292 ( .A(n74051), .Z(n74053) );
  NOR U94293 ( .A(n74053), .B(n74052), .Z(n79397) );
  NOR U94294 ( .A(n76333), .B(n79397), .Z(n74054) );
  XOR U94295 ( .A(n79398), .B(n74054), .Z(n79401) );
  XOR U94296 ( .A(n74055), .B(n79401), .Z(n79411) );
  XOR U94297 ( .A(n74056), .B(n79411), .Z(n79417) );
  IV U94298 ( .A(n74057), .Z(n74058) );
  IV U94299 ( .A(n79422), .Z(n74060) );
  NOR U94300 ( .A(n74058), .B(n74060), .Z(n79415) );
  IV U94301 ( .A(n74059), .Z(n79423) );
  NOR U94302 ( .A(n79423), .B(n74060), .Z(n79410) );
  NOR U94303 ( .A(n79415), .B(n79410), .Z(n74061) );
  XOR U94304 ( .A(n79417), .B(n74061), .Z(n76321) );
  IV U94305 ( .A(n74062), .Z(n74063) );
  NOR U94306 ( .A(n74063), .B(n74069), .Z(n74066) );
  IV U94307 ( .A(n74064), .Z(n74065) );
  NOR U94308 ( .A(n74065), .B(n74069), .Z(n76320) );
  NOR U94309 ( .A(n74066), .B(n76320), .Z(n74067) );
  XOR U94310 ( .A(n76321), .B(n74067), .Z(n79439) );
  IV U94311 ( .A(n74068), .Z(n74070) );
  NOR U94312 ( .A(n74070), .B(n74069), .Z(n76315) );
  XOR U94313 ( .A(n79439), .B(n76315), .Z(n76319) );
  XOR U94314 ( .A(n76317), .B(n76319), .Z(n79444) );
  XOR U94315 ( .A(n74071), .B(n79444), .Z(n74072) );
  IV U94316 ( .A(n74072), .Z(n79442) );
  XOR U94317 ( .A(n79440), .B(n79442), .Z(n79451) );
  XOR U94318 ( .A(n79448), .B(n79451), .Z(n79457) );
  IV U94319 ( .A(n74073), .Z(n74074) );
  NOR U94320 ( .A(n74075), .B(n74074), .Z(n79450) );
  NOR U94321 ( .A(n74077), .B(n74076), .Z(n79456) );
  NOR U94322 ( .A(n79450), .B(n79456), .Z(n74078) );
  XOR U94323 ( .A(n79457), .B(n74078), .Z(n79453) );
  XOR U94324 ( .A(n79454), .B(n79453), .Z(n79462) );
  XOR U94325 ( .A(n79461), .B(n79462), .Z(n76311) );
  XOR U94326 ( .A(n74079), .B(n76311), .Z(n76307) );
  XOR U94327 ( .A(n74080), .B(n76307), .Z(n79484) );
  XOR U94328 ( .A(n79483), .B(n79484), .Z(n79487) );
  XOR U94329 ( .A(n74081), .B(n79487), .Z(n74082) );
  IV U94330 ( .A(n74082), .Z(n79492) );
  XOR U94331 ( .A(n79490), .B(n79492), .Z(n79496) );
  IV U94332 ( .A(n74083), .Z(n74084) );
  NOR U94333 ( .A(n74085), .B(n74084), .Z(n79493) );
  IV U94334 ( .A(n74086), .Z(n79500) );
  NOR U94335 ( .A(n79500), .B(n74087), .Z(n74088) );
  NOR U94336 ( .A(n79493), .B(n74088), .Z(n79497) );
  XOR U94337 ( .A(n79496), .B(n79497), .Z(n76303) );
  XOR U94338 ( .A(n74089), .B(n76303), .Z(n85283) );
  XOR U94339 ( .A(n85281), .B(n85283), .Z(n76301) );
  XOR U94340 ( .A(n74090), .B(n76301), .Z(n79517) );
  XOR U94341 ( .A(n74091), .B(n79517), .Z(n79529) );
  XOR U94342 ( .A(n74092), .B(n79529), .Z(n79532) );
  XOR U94343 ( .A(n74093), .B(n79532), .Z(n76291) );
  XOR U94344 ( .A(n74094), .B(n76291), .Z(n79538) );
  XOR U94345 ( .A(n79536), .B(n79538), .Z(n85329) );
  XOR U94346 ( .A(n74095), .B(n85329), .Z(n74096) );
  XOR U94347 ( .A(n74097), .B(n74096), .Z(n76286) );
  XOR U94348 ( .A(n74098), .B(n76286), .Z(n76284) );
  XOR U94349 ( .A(n76282), .B(n76284), .Z(n76280) );
  XOR U94350 ( .A(n76276), .B(n76280), .Z(n74099) );
  XOR U94351 ( .A(n74100), .B(n74099), .Z(n74101) );
  IV U94352 ( .A(n74101), .Z(n76270) );
  NOR U94353 ( .A(n74103), .B(n74102), .Z(n74104) );
  IV U94354 ( .A(n74104), .Z(n74106) );
  NOR U94355 ( .A(n74106), .B(n74105), .Z(n76268) );
  XOR U94356 ( .A(n76270), .B(n76268), .Z(n76261) );
  XOR U94357 ( .A(n74107), .B(n76261), .Z(n74108) );
  IV U94358 ( .A(n74108), .Z(n76247) );
  XOR U94359 ( .A(n76245), .B(n76247), .Z(n76249) );
  XOR U94360 ( .A(n76248), .B(n76249), .Z(n76238) );
  XOR U94361 ( .A(n76237), .B(n76238), .Z(n76241) );
  XOR U94362 ( .A(n76240), .B(n76241), .Z(n79567) );
  IV U94363 ( .A(n79567), .Z(n74116) );
  IV U94364 ( .A(n74109), .Z(n74110) );
  NOR U94365 ( .A(n74111), .B(n74110), .Z(n76235) );
  IV U94366 ( .A(n74112), .Z(n74114) );
  NOR U94367 ( .A(n74114), .B(n74113), .Z(n79566) );
  NOR U94368 ( .A(n76235), .B(n79566), .Z(n74115) );
  XOR U94369 ( .A(n74116), .B(n74115), .Z(n76233) );
  XOR U94370 ( .A(n76232), .B(n76233), .Z(n79579) );
  XOR U94371 ( .A(n74117), .B(n79579), .Z(n79581) );
  XOR U94372 ( .A(n79583), .B(n79581), .Z(n76228) );
  IV U94373 ( .A(n74118), .Z(n74125) );
  XOR U94374 ( .A(n74120), .B(n74119), .Z(n74121) );
  NOR U94375 ( .A(n74122), .B(n74121), .Z(n74123) );
  IV U94376 ( .A(n74123), .Z(n74124) );
  NOR U94377 ( .A(n74125), .B(n74124), .Z(n76226) );
  XOR U94378 ( .A(n76228), .B(n76226), .Z(n76221) );
  XOR U94379 ( .A(n76220), .B(n76221), .Z(n76225) );
  IV U94380 ( .A(n74126), .Z(n74127) );
  NOR U94381 ( .A(n74128), .B(n74127), .Z(n76223) );
  XOR U94382 ( .A(n76225), .B(n76223), .Z(n76216) );
  XOR U94383 ( .A(n76215), .B(n76216), .Z(n81738) );
  XOR U94384 ( .A(n76218), .B(n81738), .Z(n76213) );
  NOR U94385 ( .A(n74129), .B(n81741), .Z(n79589) );
  IV U94386 ( .A(n74130), .Z(n74131) );
  NOR U94387 ( .A(n74132), .B(n74131), .Z(n76211) );
  NOR U94388 ( .A(n79589), .B(n76211), .Z(n74133) );
  XOR U94389 ( .A(n76213), .B(n74133), .Z(n74134) );
  IV U94390 ( .A(n74134), .Z(n76210) );
  XOR U94391 ( .A(n76208), .B(n76210), .Z(n76202) );
  XOR U94392 ( .A(n76200), .B(n76202), .Z(n76204) );
  XOR U94393 ( .A(n76203), .B(n76204), .Z(n79594) );
  XOR U94394 ( .A(n79592), .B(n79594), .Z(n79604) );
  XOR U94395 ( .A(n74135), .B(n79604), .Z(n79613) );
  XOR U94396 ( .A(n74136), .B(n79613), .Z(n79622) );
  XOR U94397 ( .A(n79620), .B(n79622), .Z(n76194) );
  XOR U94398 ( .A(n74137), .B(n76194), .Z(n74147) );
  IV U94399 ( .A(n74147), .Z(n74142) );
  IV U94400 ( .A(n74138), .Z(n74139) );
  NOR U94401 ( .A(n74140), .B(n74139), .Z(n74150) );
  IV U94402 ( .A(n74150), .Z(n74141) );
  NOR U94403 ( .A(n74142), .B(n74141), .Z(n81696) );
  IV U94404 ( .A(n74143), .Z(n74145) );
  NOR U94405 ( .A(n74145), .B(n74144), .Z(n74148) );
  IV U94406 ( .A(n74148), .Z(n74146) );
  NOR U94407 ( .A(n76194), .B(n74146), .Z(n85402) );
  NOR U94408 ( .A(n74148), .B(n74147), .Z(n74149) );
  NOR U94409 ( .A(n85402), .B(n74149), .Z(n74154) );
  NOR U94410 ( .A(n74150), .B(n74154), .Z(n74151) );
  NOR U94411 ( .A(n81696), .B(n74151), .Z(n74152) );
  NOR U94412 ( .A(n74153), .B(n74152), .Z(n74157) );
  IV U94413 ( .A(n74153), .Z(n74156) );
  IV U94414 ( .A(n74154), .Z(n74155) );
  NOR U94415 ( .A(n74156), .B(n74155), .Z(n79633) );
  NOR U94416 ( .A(n74157), .B(n79633), .Z(n79635) );
  IV U94417 ( .A(n74158), .Z(n74160) );
  NOR U94418 ( .A(n74160), .B(n74159), .Z(n74161) );
  IV U94419 ( .A(n74161), .Z(n79636) );
  XOR U94420 ( .A(n79635), .B(n79636), .Z(n79639) );
  IV U94421 ( .A(n74162), .Z(n74163) );
  NOR U94422 ( .A(n74164), .B(n74163), .Z(n79638) );
  NOR U94423 ( .A(n74166), .B(n74165), .Z(n76190) );
  NOR U94424 ( .A(n79638), .B(n76190), .Z(n74167) );
  XOR U94425 ( .A(n79639), .B(n74167), .Z(n74168) );
  IV U94426 ( .A(n74168), .Z(n76185) );
  XOR U94427 ( .A(n76184), .B(n76185), .Z(n76188) );
  XOR U94428 ( .A(n76187), .B(n76188), .Z(n76182) );
  IV U94429 ( .A(n74169), .Z(n74170) );
  NOR U94430 ( .A(n74171), .B(n74170), .Z(n76181) );
  IV U94431 ( .A(n74172), .Z(n74173) );
  NOR U94432 ( .A(n74174), .B(n74173), .Z(n76179) );
  NOR U94433 ( .A(n76181), .B(n76179), .Z(n74175) );
  XOR U94434 ( .A(n76182), .B(n74175), .Z(n74176) );
  NOR U94435 ( .A(n74177), .B(n74176), .Z(n74180) );
  IV U94436 ( .A(n74177), .Z(n74179) );
  XOR U94437 ( .A(n76181), .B(n76182), .Z(n74178) );
  NOR U94438 ( .A(n74179), .B(n74178), .Z(n81679) );
  NOR U94439 ( .A(n74180), .B(n81679), .Z(n74181) );
  IV U94440 ( .A(n74181), .Z(n79646) );
  IV U94441 ( .A(n74182), .Z(n74184) );
  NOR U94442 ( .A(n74184), .B(n74183), .Z(n79644) );
  XOR U94443 ( .A(n79646), .B(n79644), .Z(n79648) );
  XOR U94444 ( .A(n79647), .B(n79648), .Z(n74185) );
  NOR U94445 ( .A(n74186), .B(n74185), .Z(n81674) );
  IV U94446 ( .A(n74187), .Z(n74188) );
  NOR U94447 ( .A(n74189), .B(n74188), .Z(n76177) );
  NOR U94448 ( .A(n79647), .B(n76177), .Z(n74190) );
  XOR U94449 ( .A(n74190), .B(n79648), .Z(n74195) );
  NOR U94450 ( .A(n74191), .B(n74195), .Z(n74192) );
  NOR U94451 ( .A(n81674), .B(n74192), .Z(n74193) );
  NOR U94452 ( .A(n74194), .B(n74193), .Z(n74198) );
  IV U94453 ( .A(n74194), .Z(n74197) );
  IV U94454 ( .A(n74195), .Z(n74196) );
  NOR U94455 ( .A(n74197), .B(n74196), .Z(n81668) );
  NOR U94456 ( .A(n74198), .B(n81668), .Z(n74203) );
  IV U94457 ( .A(n74199), .Z(n74201) );
  NOR U94458 ( .A(n74201), .B(n74200), .Z(n74202) );
  IV U94459 ( .A(n74202), .Z(n76175) );
  XOR U94460 ( .A(n74203), .B(n76175), .Z(n74209) );
  NOR U94461 ( .A(n74212), .B(n74209), .Z(n85440) );
  IV U94462 ( .A(n74203), .Z(n76176) );
  IV U94463 ( .A(n74204), .Z(n74206) );
  NOR U94464 ( .A(n74206), .B(n74205), .Z(n74210) );
  IV U94465 ( .A(n74210), .Z(n74207) );
  NOR U94466 ( .A(n76176), .B(n74207), .Z(n85446) );
  NOR U94467 ( .A(n85440), .B(n85446), .Z(n74208) );
  IV U94468 ( .A(n74208), .Z(n79661) );
  IV U94469 ( .A(n74209), .Z(n74213) );
  NOR U94470 ( .A(n74210), .B(n74213), .Z(n74211) );
  NOR U94471 ( .A(n79661), .B(n74211), .Z(n74215) );
  NOR U94472 ( .A(n74213), .B(n74212), .Z(n74214) );
  NOR U94473 ( .A(n74215), .B(n74214), .Z(n79664) );
  IV U94474 ( .A(n74216), .Z(n74217) );
  NOR U94475 ( .A(n74218), .B(n74217), .Z(n79662) );
  IV U94476 ( .A(n74219), .Z(n74220) );
  NOR U94477 ( .A(n74226), .B(n74220), .Z(n76173) );
  NOR U94478 ( .A(n79662), .B(n76173), .Z(n74221) );
  XOR U94479 ( .A(n79664), .B(n74221), .Z(n79671) );
  IV U94480 ( .A(n74222), .Z(n74223) );
  NOR U94481 ( .A(n74224), .B(n74223), .Z(n79670) );
  IV U94482 ( .A(n74225), .Z(n74232) );
  NOR U94483 ( .A(n74227), .B(n74226), .Z(n74228) );
  IV U94484 ( .A(n74228), .Z(n74229) );
  NOR U94485 ( .A(n74230), .B(n74229), .Z(n74231) );
  IV U94486 ( .A(n74231), .Z(n74235) );
  NOR U94487 ( .A(n74232), .B(n74235), .Z(n79676) );
  NOR U94488 ( .A(n79670), .B(n79676), .Z(n74233) );
  XOR U94489 ( .A(n79671), .B(n74233), .Z(n79675) );
  IV U94490 ( .A(n74234), .Z(n74236) );
  NOR U94491 ( .A(n74236), .B(n74235), .Z(n74237) );
  IV U94492 ( .A(n74237), .Z(n79674) );
  XOR U94493 ( .A(n79675), .B(n79674), .Z(n74244) );
  IV U94494 ( .A(n74244), .Z(n74238) );
  NOR U94495 ( .A(n74239), .B(n74238), .Z(n81660) );
  IV U94496 ( .A(n74240), .Z(n74241) );
  NOR U94497 ( .A(n74242), .B(n74241), .Z(n74245) );
  IV U94498 ( .A(n74245), .Z(n74243) );
  NOR U94499 ( .A(n79675), .B(n74243), .Z(n81657) );
  NOR U94500 ( .A(n74245), .B(n74244), .Z(n74246) );
  NOR U94501 ( .A(n81657), .B(n74246), .Z(n76165) );
  NOR U94502 ( .A(n74247), .B(n76165), .Z(n74248) );
  NOR U94503 ( .A(n81660), .B(n74248), .Z(n79681) );
  XOR U94504 ( .A(n74249), .B(n79681), .Z(n85467) );
  XOR U94505 ( .A(n74250), .B(n85467), .Z(n76155) );
  XOR U94506 ( .A(n74251), .B(n76155), .Z(n79689) );
  NOR U94507 ( .A(n74252), .B(n76148), .Z(n74256) );
  IV U94508 ( .A(n74253), .Z(n74254) );
  NOR U94509 ( .A(n74255), .B(n74254), .Z(n79688) );
  NOR U94510 ( .A(n74256), .B(n79688), .Z(n74257) );
  XOR U94511 ( .A(n79689), .B(n74257), .Z(n76143) );
  IV U94512 ( .A(n74258), .Z(n74260) );
  NOR U94513 ( .A(n74260), .B(n74259), .Z(n79691) );
  NOR U94514 ( .A(n74261), .B(n76144), .Z(n74262) );
  NOR U94515 ( .A(n79691), .B(n74262), .Z(n74263) );
  XOR U94516 ( .A(n76143), .B(n74263), .Z(n76140) );
  IV U94517 ( .A(n74264), .Z(n74266) );
  NOR U94518 ( .A(n74266), .B(n74265), .Z(n76139) );
  IV U94519 ( .A(n74267), .Z(n74268) );
  NOR U94520 ( .A(n74268), .B(n74275), .Z(n76137) );
  NOR U94521 ( .A(n76139), .B(n76137), .Z(n74269) );
  XOR U94522 ( .A(n76140), .B(n74269), .Z(n76131) );
  IV U94523 ( .A(n74270), .Z(n74272) );
  NOR U94524 ( .A(n74272), .B(n74271), .Z(n81609) );
  IV U94525 ( .A(n74273), .Z(n74274) );
  NOR U94526 ( .A(n74275), .B(n74274), .Z(n81616) );
  NOR U94527 ( .A(n81609), .B(n81616), .Z(n76132) );
  XOR U94528 ( .A(n76131), .B(n76132), .Z(n76134) );
  XOR U94529 ( .A(n76133), .B(n76134), .Z(n76126) );
  XOR U94530 ( .A(n76125), .B(n76126), .Z(n85504) );
  IV U94531 ( .A(n74276), .Z(n74278) );
  NOR U94532 ( .A(n74278), .B(n74277), .Z(n76128) );
  IV U94533 ( .A(n74279), .Z(n74281) );
  NOR U94534 ( .A(n74281), .B(n74280), .Z(n76122) );
  NOR U94535 ( .A(n76128), .B(n76122), .Z(n85505) );
  XOR U94536 ( .A(n85504), .B(n85505), .Z(n74282) );
  IV U94537 ( .A(n74282), .Z(n76120) );
  IV U94538 ( .A(n74283), .Z(n74295) );
  IV U94539 ( .A(n74284), .Z(n74285) );
  NOR U94540 ( .A(n74295), .B(n74285), .Z(n74286) );
  IV U94541 ( .A(n74286), .Z(n74289) );
  NOR U94542 ( .A(n76120), .B(n74289), .Z(n76115) );
  NOR U94543 ( .A(n74288), .B(n74287), .Z(n76116) );
  XOR U94544 ( .A(n76119), .B(n76120), .Z(n76117) );
  IV U94545 ( .A(n76117), .Z(n74290) );
  XOR U94546 ( .A(n76116), .B(n74290), .Z(n74292) );
  NOR U94547 ( .A(n74290), .B(n74289), .Z(n74291) );
  NOR U94548 ( .A(n74292), .B(n74291), .Z(n74293) );
  NOR U94549 ( .A(n76115), .B(n74293), .Z(n79703) );
  IV U94550 ( .A(n74294), .Z(n74296) );
  NOR U94551 ( .A(n74296), .B(n74295), .Z(n74297) );
  IV U94552 ( .A(n74297), .Z(n79704) );
  XOR U94553 ( .A(n79703), .B(n79704), .Z(n79711) );
  IV U94554 ( .A(n74298), .Z(n74299) );
  NOR U94555 ( .A(n74302), .B(n74299), .Z(n79706) );
  IV U94556 ( .A(n74300), .Z(n74301) );
  NOR U94557 ( .A(n74302), .B(n74301), .Z(n79709) );
  NOR U94558 ( .A(n79706), .B(n79709), .Z(n74303) );
  XOR U94559 ( .A(n79711), .B(n74303), .Z(n74315) );
  IV U94560 ( .A(n74315), .Z(n74307) );
  IV U94561 ( .A(n74304), .Z(n74305) );
  NOR U94562 ( .A(n74305), .B(n79727), .Z(n74320) );
  IV U94563 ( .A(n74320), .Z(n74306) );
  NOR U94564 ( .A(n74307), .B(n74306), .Z(n81594) );
  IV U94565 ( .A(n74308), .Z(n74309) );
  NOR U94566 ( .A(n74310), .B(n74309), .Z(n76112) );
  IV U94567 ( .A(n74311), .Z(n74313) );
  NOR U94568 ( .A(n74313), .B(n74312), .Z(n74316) );
  IV U94569 ( .A(n74316), .Z(n74314) );
  NOR U94570 ( .A(n79711), .B(n74314), .Z(n79717) );
  NOR U94571 ( .A(n74316), .B(n74315), .Z(n74317) );
  NOR U94572 ( .A(n79717), .B(n74317), .Z(n74318) );
  IV U94573 ( .A(n74318), .Z(n76113) );
  XOR U94574 ( .A(n76112), .B(n76113), .Z(n76102) );
  IV U94575 ( .A(n76102), .Z(n74319) );
  NOR U94576 ( .A(n74320), .B(n74319), .Z(n74321) );
  NOR U94577 ( .A(n81594), .B(n74321), .Z(n76109) );
  NOR U94578 ( .A(n74322), .B(n76103), .Z(n74326) );
  IV U94579 ( .A(n74323), .Z(n74324) );
  NOR U94580 ( .A(n74325), .B(n74324), .Z(n76108) );
  NOR U94581 ( .A(n74326), .B(n76108), .Z(n74327) );
  XOR U94582 ( .A(n76109), .B(n74327), .Z(n76100) );
  IV U94583 ( .A(n74328), .Z(n74330) );
  NOR U94584 ( .A(n74330), .B(n74329), .Z(n76098) );
  IV U94585 ( .A(n74331), .Z(n74332) );
  NOR U94586 ( .A(n74333), .B(n74332), .Z(n76096) );
  NOR U94587 ( .A(n76098), .B(n76096), .Z(n74334) );
  XOR U94588 ( .A(n76100), .B(n74334), .Z(n76091) );
  IV U94589 ( .A(n74335), .Z(n74337) );
  NOR U94590 ( .A(n74337), .B(n74336), .Z(n76093) );
  NOR U94591 ( .A(n76093), .B(n76090), .Z(n74338) );
  XOR U94592 ( .A(n76091), .B(n74338), .Z(n76088) );
  XOR U94593 ( .A(n76086), .B(n76088), .Z(n76085) );
  XOR U94594 ( .A(n76083), .B(n76085), .Z(n74339) );
  NOR U94595 ( .A(n74340), .B(n74339), .Z(n76082) );
  IV U94596 ( .A(n74341), .Z(n74342) );
  NOR U94597 ( .A(n74343), .B(n74342), .Z(n76084) );
  NOR U94598 ( .A(n76083), .B(n76084), .Z(n74344) );
  XOR U94599 ( .A(n76085), .B(n74344), .Z(n74345) );
  NOR U94600 ( .A(n74346), .B(n74345), .Z(n74347) );
  NOR U94601 ( .A(n76082), .B(n74347), .Z(n74348) );
  IV U94602 ( .A(n74348), .Z(n76079) );
  XOR U94603 ( .A(n76078), .B(n76079), .Z(n76075) );
  IV U94604 ( .A(n74349), .Z(n74351) );
  NOR U94605 ( .A(n74351), .B(n74350), .Z(n76073) );
  XOR U94606 ( .A(n76075), .B(n76073), .Z(n81566) );
  XOR U94607 ( .A(n76076), .B(n81566), .Z(n79740) );
  XOR U94608 ( .A(n74352), .B(n79740), .Z(n76070) );
  NOR U94609 ( .A(n74354), .B(n74353), .Z(n74355) );
  IV U94610 ( .A(n74355), .Z(n74356) );
  NOR U94611 ( .A(n79744), .B(n74356), .Z(n74357) );
  XOR U94612 ( .A(n76070), .B(n74357), .Z(n74364) );
  IV U94613 ( .A(n74364), .Z(n74358) );
  NOR U94614 ( .A(n74363), .B(n74358), .Z(n74359) );
  IV U94615 ( .A(n74359), .Z(n74360) );
  NOR U94616 ( .A(n74361), .B(n74360), .Z(n81541) );
  IV U94617 ( .A(n74361), .Z(n74362) );
  NOR U94618 ( .A(n74362), .B(n74364), .Z(n81555) );
  IV U94619 ( .A(n74363), .Z(n74365) );
  NOR U94620 ( .A(n74365), .B(n74364), .Z(n81548) );
  NOR U94621 ( .A(n81555), .B(n81548), .Z(n74366) );
  IV U94622 ( .A(n74366), .Z(n81538) );
  NOR U94623 ( .A(n81541), .B(n81538), .Z(n76059) );
  IV U94624 ( .A(n74367), .Z(n74369) );
  NOR U94625 ( .A(n74369), .B(n74368), .Z(n81537) );
  IV U94626 ( .A(n74370), .Z(n74371) );
  NOR U94627 ( .A(n74372), .B(n74371), .Z(n81545) );
  NOR U94628 ( .A(n81537), .B(n81545), .Z(n76061) );
  XOR U94629 ( .A(n76059), .B(n76061), .Z(n76055) );
  NOR U94630 ( .A(n74373), .B(n76055), .Z(n76053) );
  NOR U94631 ( .A(n74380), .B(n76053), .Z(n74374) );
  IV U94632 ( .A(n74374), .Z(n74379) );
  NOR U94633 ( .A(n74375), .B(n76056), .Z(n74376) );
  XOR U94634 ( .A(n74376), .B(n76055), .Z(n76048) );
  IV U94635 ( .A(n76048), .Z(n74382) );
  NOR U94636 ( .A(n74377), .B(n74382), .Z(n74378) );
  NOR U94637 ( .A(n74379), .B(n74378), .Z(n74384) );
  IV U94638 ( .A(n74380), .Z(n74381) );
  NOR U94639 ( .A(n74382), .B(n74381), .Z(n74383) );
  NOR U94640 ( .A(n74384), .B(n74383), .Z(n79759) );
  IV U94641 ( .A(n74385), .Z(n74392) );
  IV U94642 ( .A(n74386), .Z(n74387) );
  NOR U94643 ( .A(n74392), .B(n74387), .Z(n79757) );
  XOR U94644 ( .A(n79759), .B(n79757), .Z(n79761) );
  NOR U94645 ( .A(n74393), .B(n79761), .Z(n81517) );
  IV U94646 ( .A(n74388), .Z(n74389) );
  NOR U94647 ( .A(n74389), .B(n74400), .Z(n79774) );
  IV U94648 ( .A(n74390), .Z(n74391) );
  NOR U94649 ( .A(n74392), .B(n74391), .Z(n79760) );
  XOR U94650 ( .A(n79760), .B(n79761), .Z(n79775) );
  IV U94651 ( .A(n79775), .Z(n74394) );
  XOR U94652 ( .A(n79774), .B(n74394), .Z(n74396) );
  NOR U94653 ( .A(n74394), .B(n74393), .Z(n74395) );
  NOR U94654 ( .A(n74396), .B(n74395), .Z(n74397) );
  NOR U94655 ( .A(n81517), .B(n74397), .Z(n74398) );
  IV U94656 ( .A(n74398), .Z(n79768) );
  IV U94657 ( .A(n74399), .Z(n74401) );
  NOR U94658 ( .A(n74401), .B(n74400), .Z(n79766) );
  XOR U94659 ( .A(n79768), .B(n79766), .Z(n79773) );
  IV U94660 ( .A(n74402), .Z(n74403) );
  NOR U94661 ( .A(n74404), .B(n74403), .Z(n79771) );
  XOR U94662 ( .A(n79773), .B(n79771), .Z(n79787) );
  IV U94663 ( .A(n74405), .Z(n74406) );
  NOR U94664 ( .A(n74407), .B(n74406), .Z(n76045) );
  IV U94665 ( .A(n74408), .Z(n74410) );
  NOR U94666 ( .A(n74410), .B(n74409), .Z(n79786) );
  NOR U94667 ( .A(n76045), .B(n79786), .Z(n74411) );
  XOR U94668 ( .A(n79787), .B(n74411), .Z(n79789) );
  IV U94669 ( .A(n74412), .Z(n74413) );
  NOR U94670 ( .A(n74413), .B(n79794), .Z(n74417) );
  IV U94671 ( .A(n74414), .Z(n74415) );
  NOR U94672 ( .A(n74416), .B(n74415), .Z(n79803) );
  NOR U94673 ( .A(n74417), .B(n79803), .Z(n74418) );
  XOR U94674 ( .A(n79789), .B(n74418), .Z(n76044) );
  XOR U94675 ( .A(n74419), .B(n76044), .Z(n76038) );
  XOR U94676 ( .A(n76039), .B(n76038), .Z(n76035) );
  XOR U94677 ( .A(n76033), .B(n76035), .Z(n79816) );
  IV U94678 ( .A(n74420), .Z(n74421) );
  NOR U94679 ( .A(n74422), .B(n74421), .Z(n76036) );
  IV U94680 ( .A(n74423), .Z(n74425) );
  NOR U94681 ( .A(n74425), .B(n74424), .Z(n79815) );
  NOR U94682 ( .A(n76036), .B(n79815), .Z(n74426) );
  XOR U94683 ( .A(n79816), .B(n74426), .Z(n79812) );
  XOR U94684 ( .A(n79813), .B(n79812), .Z(n79809) );
  IV U94685 ( .A(n74427), .Z(n74428) );
  NOR U94686 ( .A(n74429), .B(n74428), .Z(n76031) );
  IV U94687 ( .A(n74430), .Z(n74431) );
  NOR U94688 ( .A(n74432), .B(n74431), .Z(n79808) );
  NOR U94689 ( .A(n76031), .B(n79808), .Z(n74433) );
  XOR U94690 ( .A(n79809), .B(n74433), .Z(n76024) );
  IV U94691 ( .A(n74434), .Z(n74436) );
  NOR U94692 ( .A(n74436), .B(n74435), .Z(n76027) );
  IV U94693 ( .A(n74437), .Z(n74439) );
  NOR U94694 ( .A(n74439), .B(n74438), .Z(n76025) );
  NOR U94695 ( .A(n76027), .B(n76025), .Z(n74440) );
  XOR U94696 ( .A(n76024), .B(n74440), .Z(n85579) );
  IV U94697 ( .A(n74441), .Z(n74443) );
  NOR U94698 ( .A(n74443), .B(n74442), .Z(n85577) );
  IV U94699 ( .A(n74444), .Z(n74445) );
  NOR U94700 ( .A(n74446), .B(n74445), .Z(n81490) );
  NOR U94701 ( .A(n85577), .B(n81490), .Z(n76019) );
  XOR U94702 ( .A(n85579), .B(n76019), .Z(n76012) );
  XOR U94703 ( .A(n74447), .B(n76012), .Z(n76009) );
  IV U94704 ( .A(n74448), .Z(n74450) );
  NOR U94705 ( .A(n74450), .B(n74449), .Z(n76014) );
  IV U94706 ( .A(n74451), .Z(n74453) );
  NOR U94707 ( .A(n74453), .B(n74452), .Z(n76008) );
  NOR U94708 ( .A(n76014), .B(n76008), .Z(n74454) );
  XOR U94709 ( .A(n76009), .B(n74454), .Z(n74455) );
  IV U94710 ( .A(n74455), .Z(n76007) );
  IV U94711 ( .A(n74456), .Z(n74457) );
  NOR U94712 ( .A(n74458), .B(n74457), .Z(n76005) );
  IV U94713 ( .A(n74459), .Z(n74460) );
  NOR U94714 ( .A(n74460), .B(n75999), .Z(n74461) );
  NOR U94715 ( .A(n76005), .B(n74461), .Z(n74462) );
  XOR U94716 ( .A(n76007), .B(n74462), .Z(n75996) );
  IV U94717 ( .A(n74463), .Z(n74465) );
  NOR U94718 ( .A(n74465), .B(n74464), .Z(n75995) );
  NOR U94719 ( .A(n79822), .B(n75995), .Z(n74466) );
  XOR U94720 ( .A(n75996), .B(n74466), .Z(n75994) );
  XOR U94721 ( .A(n75992), .B(n75994), .Z(n75990) );
  XOR U94722 ( .A(n74467), .B(n75990), .Z(n75981) );
  XOR U94723 ( .A(n74468), .B(n75981), .Z(n79836) );
  XOR U94724 ( .A(n79834), .B(n79836), .Z(n79838) );
  XOR U94725 ( .A(n79837), .B(n79838), .Z(n75975) );
  XOR U94726 ( .A(n75973), .B(n75975), .Z(n75977) );
  XOR U94727 ( .A(n75976), .B(n75977), .Z(n79843) );
  XOR U94728 ( .A(n79842), .B(n79843), .Z(n79854) );
  NOR U94729 ( .A(n74469), .B(n79854), .Z(n85620) );
  IV U94730 ( .A(n74470), .Z(n74471) );
  NOR U94731 ( .A(n74472), .B(n74471), .Z(n75971) );
  IV U94732 ( .A(n74473), .Z(n74475) );
  NOR U94733 ( .A(n74475), .B(n74474), .Z(n75968) );
  IV U94734 ( .A(n74476), .Z(n74477) );
  NOR U94735 ( .A(n74478), .B(n74477), .Z(n79853) );
  XOR U94736 ( .A(n79853), .B(n79854), .Z(n75970) );
  XOR U94737 ( .A(n75962), .B(n75964), .Z(n75966) );
  XOR U94738 ( .A(n74479), .B(n75966), .Z(n75955) );
  IV U94739 ( .A(n74480), .Z(n74481) );
  NOR U94740 ( .A(n74482), .B(n74481), .Z(n75959) );
  NOR U94741 ( .A(n74484), .B(n74483), .Z(n75954) );
  NOR U94742 ( .A(n75959), .B(n75954), .Z(n74485) );
  XOR U94743 ( .A(n75955), .B(n74485), .Z(n75949) );
  XOR U94744 ( .A(n75948), .B(n75949), .Z(n75952) );
  XOR U94745 ( .A(n75951), .B(n75952), .Z(n79866) );
  XOR U94746 ( .A(n74486), .B(n79866), .Z(n79862) );
  XOR U94747 ( .A(n79863), .B(n79862), .Z(n75942) );
  XOR U94748 ( .A(n75941), .B(n75942), .Z(n75937) );
  XOR U94749 ( .A(n74487), .B(n75937), .Z(n75933) );
  IV U94750 ( .A(n74488), .Z(n74489) );
  NOR U94751 ( .A(n74489), .B(n74491), .Z(n79869) );
  IV U94752 ( .A(n74490), .Z(n74492) );
  NOR U94753 ( .A(n74492), .B(n74491), .Z(n75934) );
  NOR U94754 ( .A(n79869), .B(n75934), .Z(n74493) );
  XOR U94755 ( .A(n75933), .B(n74493), .Z(n75932) );
  XOR U94756 ( .A(n75930), .B(n75932), .Z(n79875) );
  XOR U94757 ( .A(n74494), .B(n79875), .Z(n79877) );
  XOR U94758 ( .A(n79878), .B(n79877), .Z(n79881) );
  XOR U94759 ( .A(n79880), .B(n79881), .Z(n75924) );
  IV U94760 ( .A(n74495), .Z(n74497) );
  NOR U94761 ( .A(n74497), .B(n74496), .Z(n75922) );
  XOR U94762 ( .A(n75924), .B(n75922), .Z(n79892) );
  IV U94763 ( .A(n74498), .Z(n74501) );
  IV U94764 ( .A(n74499), .Z(n74500) );
  NOR U94765 ( .A(n74501), .B(n74500), .Z(n75925) );
  XOR U94766 ( .A(n79892), .B(n75925), .Z(n79907) );
  XOR U94767 ( .A(n74502), .B(n79907), .Z(n79902) );
  IV U94768 ( .A(n74503), .Z(n74505) );
  NOR U94769 ( .A(n74505), .B(n74504), .Z(n75919) );
  IV U94770 ( .A(n74506), .Z(n74507) );
  NOR U94771 ( .A(n74508), .B(n74507), .Z(n79906) );
  IV U94772 ( .A(n74509), .Z(n74511) );
  NOR U94773 ( .A(n74511), .B(n74510), .Z(n79901) );
  NOR U94774 ( .A(n79906), .B(n79901), .Z(n74512) );
  IV U94775 ( .A(n74512), .Z(n74513) );
  NOR U94776 ( .A(n75919), .B(n74513), .Z(n74514) );
  XOR U94777 ( .A(n79902), .B(n74514), .Z(n75913) );
  XOR U94778 ( .A(n75914), .B(n75913), .Z(n79920) );
  XOR U94779 ( .A(n74515), .B(n79920), .Z(n75906) );
  XOR U94780 ( .A(n74516), .B(n75906), .Z(n79929) );
  XOR U94781 ( .A(n74517), .B(n79929), .Z(n79938) );
  XOR U94782 ( .A(n79937), .B(n79938), .Z(n79942) );
  IV U94783 ( .A(n74518), .Z(n74519) );
  NOR U94784 ( .A(n74520), .B(n74519), .Z(n79941) );
  IV U94785 ( .A(n74521), .Z(n74523) );
  NOR U94786 ( .A(n74523), .B(n74522), .Z(n79946) );
  NOR U94787 ( .A(n79941), .B(n79946), .Z(n74524) );
  XOR U94788 ( .A(n79942), .B(n74524), .Z(n79953) );
  XOR U94789 ( .A(n74525), .B(n79953), .Z(n79960) );
  XOR U94790 ( .A(n74526), .B(n79960), .Z(n79966) );
  XOR U94791 ( .A(n79967), .B(n79966), .Z(n79969) );
  XOR U94792 ( .A(n79968), .B(n79969), .Z(n79981) );
  XOR U94793 ( .A(n74527), .B(n79981), .Z(n79977) );
  XOR U94794 ( .A(n79978), .B(n79977), .Z(n75882) );
  NOR U94795 ( .A(n74528), .B(n74529), .Z(n74533) );
  IV U94796 ( .A(n74529), .Z(n75883) );
  NOR U94797 ( .A(n75883), .B(n74530), .Z(n79983) );
  NOR U94798 ( .A(n74531), .B(n79983), .Z(n74532) );
  NOR U94799 ( .A(n74533), .B(n74532), .Z(n74534) );
  XOR U94800 ( .A(n75882), .B(n74534), .Z(n75876) );
  IV U94801 ( .A(n75876), .Z(n75874) );
  IV U94802 ( .A(n74535), .Z(n74536) );
  NOR U94803 ( .A(n74537), .B(n74536), .Z(n75873) );
  IV U94804 ( .A(n75873), .Z(n75875) );
  XOR U94805 ( .A(n75874), .B(n75875), .Z(n75872) );
  IV U94806 ( .A(n74538), .Z(n74540) );
  NOR U94807 ( .A(n74540), .B(n74539), .Z(n75878) );
  IV U94808 ( .A(n74541), .Z(n74542) );
  NOR U94809 ( .A(n74542), .B(n74548), .Z(n75870) );
  NOR U94810 ( .A(n75878), .B(n75870), .Z(n74543) );
  XOR U94811 ( .A(n75872), .B(n74543), .Z(n75861) );
  IV U94812 ( .A(n74544), .Z(n74546) );
  NOR U94813 ( .A(n74546), .B(n74545), .Z(n75862) );
  IV U94814 ( .A(n74547), .Z(n74549) );
  NOR U94815 ( .A(n74549), .B(n74548), .Z(n75867) );
  NOR U94816 ( .A(n75862), .B(n75867), .Z(n74550) );
  XOR U94817 ( .A(n75861), .B(n74550), .Z(n75865) );
  IV U94818 ( .A(n75865), .Z(n74558) );
  IV U94819 ( .A(n74551), .Z(n74552) );
  NOR U94820 ( .A(n74553), .B(n74552), .Z(n75864) );
  IV U94821 ( .A(n74554), .Z(n74555) );
  NOR U94822 ( .A(n74556), .B(n74555), .Z(n75859) );
  NOR U94823 ( .A(n75864), .B(n75859), .Z(n74557) );
  XOR U94824 ( .A(n74558), .B(n74557), .Z(n79994) );
  IV U94825 ( .A(n74559), .Z(n74560) );
  NOR U94826 ( .A(n74561), .B(n74560), .Z(n79992) );
  IV U94827 ( .A(n74562), .Z(n74563) );
  NOR U94828 ( .A(n74564), .B(n74563), .Z(n79990) );
  NOR U94829 ( .A(n79992), .B(n79990), .Z(n74565) );
  XOR U94830 ( .A(n79994), .B(n74565), .Z(n75854) );
  IV U94831 ( .A(n74566), .Z(n74568) );
  NOR U94832 ( .A(n74568), .B(n74567), .Z(n79987) );
  IV U94833 ( .A(n74569), .Z(n74570) );
  NOR U94834 ( .A(n74570), .B(n74572), .Z(n75853) );
  IV U94835 ( .A(n74571), .Z(n74573) );
  NOR U94836 ( .A(n74573), .B(n74572), .Z(n75856) );
  NOR U94837 ( .A(n75853), .B(n75856), .Z(n74574) );
  IV U94838 ( .A(n74574), .Z(n74575) );
  NOR U94839 ( .A(n79987), .B(n74575), .Z(n74576) );
  XOR U94840 ( .A(n75854), .B(n74576), .Z(n75847) );
  XOR U94841 ( .A(n74577), .B(n75847), .Z(n75844) );
  IV U94842 ( .A(n74578), .Z(n74580) );
  NOR U94843 ( .A(n74580), .B(n74579), .Z(n75842) );
  IV U94844 ( .A(n74581), .Z(n74582) );
  NOR U94845 ( .A(n74582), .B(n74586), .Z(n75840) );
  NOR U94846 ( .A(n75842), .B(n75840), .Z(n74583) );
  XOR U94847 ( .A(n75844), .B(n74583), .Z(n74584) );
  IV U94848 ( .A(n74584), .Z(n80001) );
  IV U94849 ( .A(n74585), .Z(n74587) );
  NOR U94850 ( .A(n74587), .B(n74586), .Z(n74588) );
  IV U94851 ( .A(n74588), .Z(n75839) );
  XOR U94852 ( .A(n80001), .B(n75839), .Z(n74589) );
  XOR U94853 ( .A(n74590), .B(n74589), .Z(n75835) );
  IV U94854 ( .A(n74591), .Z(n74592) );
  NOR U94855 ( .A(n74593), .B(n74592), .Z(n74597) );
  IV U94856 ( .A(n74594), .Z(n74595) );
  NOR U94857 ( .A(n74595), .B(n74603), .Z(n74596) );
  NOR U94858 ( .A(n74597), .B(n74596), .Z(n75834) );
  XOR U94859 ( .A(n75835), .B(n75834), .Z(n75831) );
  IV U94860 ( .A(n74598), .Z(n74599) );
  NOR U94861 ( .A(n74600), .B(n74599), .Z(n80006) );
  IV U94862 ( .A(n74601), .Z(n74602) );
  NOR U94863 ( .A(n74603), .B(n74602), .Z(n75832) );
  NOR U94864 ( .A(n80006), .B(n75832), .Z(n74604) );
  XOR U94865 ( .A(n75831), .B(n74604), .Z(n80005) );
  XOR U94866 ( .A(n80003), .B(n80005), .Z(n74605) );
  XOR U94867 ( .A(n74606), .B(n74605), .Z(n80015) );
  XOR U94868 ( .A(n74607), .B(n80015), .Z(n80012) );
  XOR U94869 ( .A(n74608), .B(n80012), .Z(n75810) );
  XOR U94870 ( .A(n75811), .B(n75810), .Z(n75813) );
  XOR U94871 ( .A(n74609), .B(n75813), .Z(n74622) );
  XOR U94872 ( .A(n75809), .B(n74622), .Z(n74619) );
  IV U94873 ( .A(n74619), .Z(n74617) );
  IV U94874 ( .A(n74610), .Z(n74611) );
  NOR U94875 ( .A(n74612), .B(n74611), .Z(n74621) );
  IV U94876 ( .A(n74613), .Z(n74614) );
  NOR U94877 ( .A(n74614), .B(n74634), .Z(n74618) );
  NOR U94878 ( .A(n74621), .B(n74618), .Z(n74615) );
  IV U94879 ( .A(n74615), .Z(n74616) );
  NOR U94880 ( .A(n74617), .B(n74616), .Z(n74625) );
  IV U94881 ( .A(n74618), .Z(n74620) );
  NOR U94882 ( .A(n74620), .B(n74619), .Z(n81272) );
  IV U94883 ( .A(n74621), .Z(n74623) );
  IV U94884 ( .A(n74622), .Z(n75808) );
  NOR U94885 ( .A(n74623), .B(n75808), .Z(n81270) );
  NOR U94886 ( .A(n81272), .B(n81270), .Z(n74624) );
  IV U94887 ( .A(n74624), .Z(n80033) );
  NOR U94888 ( .A(n74625), .B(n80033), .Z(n74626) );
  IV U94889 ( .A(n74626), .Z(n80030) );
  IV U94890 ( .A(n74627), .Z(n74628) );
  NOR U94891 ( .A(n74628), .B(n74634), .Z(n80028) );
  XOR U94892 ( .A(n80030), .B(n80028), .Z(n80040) );
  IV U94893 ( .A(n74629), .Z(n74630) );
  NOR U94894 ( .A(n74631), .B(n74630), .Z(n80039) );
  IV U94895 ( .A(n74632), .Z(n74633) );
  NOR U94896 ( .A(n74634), .B(n74633), .Z(n75804) );
  NOR U94897 ( .A(n80039), .B(n75804), .Z(n74635) );
  XOR U94898 ( .A(n80040), .B(n74635), .Z(n75799) );
  XOR U94899 ( .A(n74636), .B(n75799), .Z(n85763) );
  XOR U94900 ( .A(n80045), .B(n85763), .Z(n75791) );
  XOR U94901 ( .A(n74637), .B(n75791), .Z(n80058) );
  XOR U94902 ( .A(n80056), .B(n80058), .Z(n74649) );
  IV U94903 ( .A(n74649), .Z(n74645) );
  IV U94904 ( .A(n74638), .Z(n74639) );
  NOR U94905 ( .A(n74642), .B(n74639), .Z(n74648) );
  IV U94906 ( .A(n74640), .Z(n74641) );
  NOR U94907 ( .A(n74642), .B(n74641), .Z(n74646) );
  NOR U94908 ( .A(n74648), .B(n74646), .Z(n74643) );
  IV U94909 ( .A(n74643), .Z(n74644) );
  NOR U94910 ( .A(n74645), .B(n74644), .Z(n74651) );
  IV U94911 ( .A(n74646), .Z(n74647) );
  NOR U94912 ( .A(n80058), .B(n74647), .Z(n85773) );
  IV U94913 ( .A(n74648), .Z(n74650) );
  NOR U94914 ( .A(n74650), .B(n74649), .Z(n85782) );
  NOR U94915 ( .A(n85773), .B(n85782), .Z(n87015) );
  IV U94916 ( .A(n87015), .Z(n80074) );
  NOR U94917 ( .A(n74651), .B(n80074), .Z(n74652) );
  IV U94918 ( .A(n74652), .Z(n80072) );
  IV U94919 ( .A(n74653), .Z(n74655) );
  NOR U94920 ( .A(n74655), .B(n74654), .Z(n80071) );
  IV U94921 ( .A(n74656), .Z(n74657) );
  NOR U94922 ( .A(n74658), .B(n74657), .Z(n80069) );
  NOR U94923 ( .A(n80071), .B(n80069), .Z(n74659) );
  XOR U94924 ( .A(n80072), .B(n74659), .Z(n74660) );
  NOR U94925 ( .A(n74661), .B(n74660), .Z(n74664) );
  IV U94926 ( .A(n74661), .Z(n74663) );
  XOR U94927 ( .A(n80071), .B(n80072), .Z(n74662) );
  NOR U94928 ( .A(n74663), .B(n74662), .Z(n80077) );
  NOR U94929 ( .A(n74664), .B(n80077), .Z(n74665) );
  IV U94930 ( .A(n74665), .Z(n80081) );
  IV U94931 ( .A(n74666), .Z(n74668) );
  IV U94932 ( .A(n74667), .Z(n74670) );
  NOR U94933 ( .A(n74668), .B(n74670), .Z(n80079) );
  XOR U94934 ( .A(n80081), .B(n80079), .Z(n80084) );
  IV U94935 ( .A(n74669), .Z(n74671) );
  NOR U94936 ( .A(n74671), .B(n74670), .Z(n80082) );
  XOR U94937 ( .A(n80084), .B(n80082), .Z(n80087) );
  IV U94938 ( .A(n80087), .Z(n74678) );
  IV U94939 ( .A(n74672), .Z(n74673) );
  NOR U94940 ( .A(n74676), .B(n74673), .Z(n80086) );
  IV U94941 ( .A(n74674), .Z(n74675) );
  NOR U94942 ( .A(n74676), .B(n74675), .Z(n75788) );
  NOR U94943 ( .A(n80086), .B(n75788), .Z(n74677) );
  XOR U94944 ( .A(n74678), .B(n74677), .Z(n81242) );
  XOR U94945 ( .A(n75784), .B(n81242), .Z(n81235) );
  XOR U94946 ( .A(n74679), .B(n81235), .Z(n75782) );
  IV U94947 ( .A(n74680), .Z(n74681) );
  NOR U94948 ( .A(n74681), .B(n74686), .Z(n75780) );
  XOR U94949 ( .A(n75782), .B(n75780), .Z(n81228) );
  IV U94950 ( .A(n74682), .Z(n74684) );
  NOR U94951 ( .A(n74684), .B(n74683), .Z(n85792) );
  IV U94952 ( .A(n74685), .Z(n74687) );
  NOR U94953 ( .A(n74687), .B(n74686), .Z(n81226) );
  NOR U94954 ( .A(n85792), .B(n81226), .Z(n80091) );
  XOR U94955 ( .A(n81228), .B(n80091), .Z(n74688) );
  IV U94956 ( .A(n74688), .Z(n80093) );
  XOR U94957 ( .A(n80092), .B(n80093), .Z(n85799) );
  XOR U94958 ( .A(n74689), .B(n85799), .Z(n74690) );
  IV U94959 ( .A(n74690), .Z(n80102) );
  XOR U94960 ( .A(n80101), .B(n80102), .Z(n80110) );
  XOR U94961 ( .A(n80109), .B(n80110), .Z(n80112) );
  XOR U94962 ( .A(n80113), .B(n80112), .Z(n74691) );
  XOR U94963 ( .A(n74692), .B(n74691), .Z(n80119) );
  IV U94964 ( .A(n74693), .Z(n74695) );
  NOR U94965 ( .A(n74695), .B(n74694), .Z(n80117) );
  XOR U94966 ( .A(n80119), .B(n80117), .Z(n75773) );
  XOR U94967 ( .A(n75772), .B(n75773), .Z(n80126) );
  IV U94968 ( .A(n74696), .Z(n74697) );
  NOR U94969 ( .A(n74698), .B(n74697), .Z(n80115) );
  IV U94970 ( .A(n74699), .Z(n74701) );
  NOR U94971 ( .A(n74701), .B(n74700), .Z(n80125) );
  NOR U94972 ( .A(n80115), .B(n80125), .Z(n74702) );
  XOR U94973 ( .A(n80126), .B(n74702), .Z(n75762) );
  XOR U94974 ( .A(n74703), .B(n75762), .Z(n75765) );
  XOR U94975 ( .A(n75764), .B(n75765), .Z(n80131) );
  IV U94976 ( .A(n74704), .Z(n74706) );
  NOR U94977 ( .A(n74706), .B(n74705), .Z(n75759) );
  IV U94978 ( .A(n74707), .Z(n74708) );
  NOR U94979 ( .A(n74709), .B(n74708), .Z(n80130) );
  NOR U94980 ( .A(n75759), .B(n80130), .Z(n74710) );
  XOR U94981 ( .A(n80131), .B(n74710), .Z(n74716) );
  XOR U94982 ( .A(n80133), .B(n74716), .Z(n74722) );
  IV U94983 ( .A(n74722), .Z(n74711) );
  NOR U94984 ( .A(n74712), .B(n74711), .Z(n80144) );
  IV U94985 ( .A(n74713), .Z(n74715) );
  NOR U94986 ( .A(n74715), .B(n74714), .Z(n74719) );
  IV U94987 ( .A(n74719), .Z(n74717) );
  IV U94988 ( .A(n74716), .Z(n80134) );
  NOR U94989 ( .A(n74717), .B(n80134), .Z(n81188) );
  NOR U94990 ( .A(n74719), .B(n74718), .Z(n74720) );
  IV U94991 ( .A(n74720), .Z(n74721) );
  NOR U94992 ( .A(n74722), .B(n74721), .Z(n74723) );
  NOR U94993 ( .A(n81188), .B(n74723), .Z(n74724) );
  IV U94994 ( .A(n74724), .Z(n80141) );
  NOR U94995 ( .A(n80144), .B(n80141), .Z(n80149) );
  IV U94996 ( .A(n74725), .Z(n74726) );
  NOR U94997 ( .A(n74727), .B(n74726), .Z(n80140) );
  IV U94998 ( .A(n74728), .Z(n74730) );
  NOR U94999 ( .A(n74730), .B(n74729), .Z(n80148) );
  NOR U95000 ( .A(n80140), .B(n80148), .Z(n74731) );
  XOR U95001 ( .A(n80149), .B(n74731), .Z(n80147) );
  IV U95002 ( .A(n74732), .Z(n74734) );
  NOR U95003 ( .A(n74734), .B(n74733), .Z(n80145) );
  IV U95004 ( .A(n74735), .Z(n74736) );
  NOR U95005 ( .A(n74736), .B(n74739), .Z(n75757) );
  NOR U95006 ( .A(n80145), .B(n75757), .Z(n74737) );
  XOR U95007 ( .A(n80147), .B(n74737), .Z(n75748) );
  IV U95008 ( .A(n74738), .Z(n74740) );
  NOR U95009 ( .A(n74740), .B(n74739), .Z(n74741) );
  IV U95010 ( .A(n74741), .Z(n75749) );
  XOR U95011 ( .A(n75748), .B(n75749), .Z(n75755) );
  IV U95012 ( .A(n74742), .Z(n74744) );
  NOR U95013 ( .A(n74744), .B(n74743), .Z(n75745) );
  NOR U95014 ( .A(n74746), .B(n74745), .Z(n75754) );
  NOR U95015 ( .A(n75745), .B(n75754), .Z(n74747) );
  XOR U95016 ( .A(n75755), .B(n74747), .Z(n74757) );
  IV U95017 ( .A(n74757), .Z(n74748) );
  NOR U95018 ( .A(n74749), .B(n74748), .Z(n80159) );
  IV U95019 ( .A(n74750), .Z(n74752) );
  NOR U95020 ( .A(n74752), .B(n74751), .Z(n75746) );
  IV U95021 ( .A(n75746), .Z(n74753) );
  NOR U95022 ( .A(n74753), .B(n75755), .Z(n85841) );
  NOR U95023 ( .A(n74754), .B(n75746), .Z(n74755) );
  IV U95024 ( .A(n74755), .Z(n74756) );
  NOR U95025 ( .A(n74757), .B(n74756), .Z(n74758) );
  NOR U95026 ( .A(n85841), .B(n74758), .Z(n74759) );
  IV U95027 ( .A(n74759), .Z(n80156) );
  NOR U95028 ( .A(n80159), .B(n80156), .Z(n74760) );
  IV U95029 ( .A(n74760), .Z(n75740) );
  IV U95030 ( .A(n74761), .Z(n74763) );
  NOR U95031 ( .A(n74763), .B(n74762), .Z(n80155) );
  NOR U95032 ( .A(n74764), .B(n75741), .Z(n74765) );
  NOR U95033 ( .A(n80155), .B(n74765), .Z(n74766) );
  XOR U95034 ( .A(n75740), .B(n74766), .Z(n75735) );
  XOR U95035 ( .A(n75732), .B(n75735), .Z(n80166) );
  XOR U95036 ( .A(n74767), .B(n80166), .Z(n80162) );
  XOR U95037 ( .A(n80163), .B(n80162), .Z(n75728) );
  IV U95038 ( .A(n74768), .Z(n74771) );
  IV U95039 ( .A(n74769), .Z(n74770) );
  NOR U95040 ( .A(n74771), .B(n74770), .Z(n75722) );
  NOR U95041 ( .A(n75727), .B(n75722), .Z(n74772) );
  XOR U95042 ( .A(n75728), .B(n74772), .Z(n75720) );
  XOR U95043 ( .A(n74773), .B(n75720), .Z(n75718) );
  IV U95044 ( .A(n74774), .Z(n74776) );
  NOR U95045 ( .A(n74776), .B(n74775), .Z(n75716) );
  XOR U95046 ( .A(n75718), .B(n75716), .Z(n80174) );
  IV U95047 ( .A(n74777), .Z(n74778) );
  NOR U95048 ( .A(n74779), .B(n74778), .Z(n80172) );
  XOR U95049 ( .A(n80174), .B(n80172), .Z(n80179) );
  XOR U95050 ( .A(n80175), .B(n80179), .Z(n75713) );
  IV U95051 ( .A(n74780), .Z(n74782) );
  NOR U95052 ( .A(n74782), .B(n74781), .Z(n80178) );
  IV U95053 ( .A(n74783), .Z(n74785) );
  NOR U95054 ( .A(n74785), .B(n74784), .Z(n75712) );
  NOR U95055 ( .A(n80178), .B(n75712), .Z(n74786) );
  XOR U95056 ( .A(n75713), .B(n74786), .Z(n75708) );
  XOR U95057 ( .A(n75706), .B(n75708), .Z(n75711) );
  XOR U95058 ( .A(n75709), .B(n75711), .Z(n80186) );
  XOR U95059 ( .A(n80184), .B(n80186), .Z(n75704) );
  XOR U95060 ( .A(n75705), .B(n75704), .Z(n74787) );
  IV U95061 ( .A(n74787), .Z(n80205) );
  IV U95062 ( .A(n74788), .Z(n75701) );
  NOR U95063 ( .A(n74789), .B(n75701), .Z(n74790) );
  XOR U95064 ( .A(n80205), .B(n74790), .Z(n75698) );
  IV U95065 ( .A(n75698), .Z(n74798) );
  IV U95066 ( .A(n74791), .Z(n74793) );
  NOR U95067 ( .A(n74793), .B(n74792), .Z(n80204) );
  IV U95068 ( .A(n74794), .Z(n74795) );
  NOR U95069 ( .A(n74796), .B(n74795), .Z(n75697) );
  NOR U95070 ( .A(n80204), .B(n75697), .Z(n74797) );
  XOR U95071 ( .A(n74798), .B(n74797), .Z(n75696) );
  XOR U95072 ( .A(n75695), .B(n75696), .Z(n74809) );
  IV U95073 ( .A(n74809), .Z(n74799) );
  NOR U95074 ( .A(n74800), .B(n74799), .Z(n75694) );
  IV U95075 ( .A(n74801), .Z(n74802) );
  NOR U95076 ( .A(n74803), .B(n74802), .Z(n74806) );
  IV U95077 ( .A(n74806), .Z(n74804) );
  NOR U95078 ( .A(n75696), .B(n74804), .Z(n81139) );
  NOR U95079 ( .A(n74806), .B(n74805), .Z(n74807) );
  IV U95080 ( .A(n74807), .Z(n74808) );
  NOR U95081 ( .A(n74809), .B(n74808), .Z(n74810) );
  NOR U95082 ( .A(n81139), .B(n74810), .Z(n74811) );
  IV U95083 ( .A(n74811), .Z(n75685) );
  NOR U95084 ( .A(n75694), .B(n75685), .Z(n74812) );
  IV U95085 ( .A(n74812), .Z(n75682) );
  NOR U95086 ( .A(n74813), .B(n75686), .Z(n74817) );
  IV U95087 ( .A(n74814), .Z(n74815) );
  NOR U95088 ( .A(n74816), .B(n74815), .Z(n75681) );
  NOR U95089 ( .A(n74817), .B(n75681), .Z(n74818) );
  XOR U95090 ( .A(n75682), .B(n74818), .Z(n74829) );
  IV U95091 ( .A(n74829), .Z(n80218) );
  XOR U95092 ( .A(n80213), .B(n80218), .Z(n74819) );
  NOR U95093 ( .A(n74820), .B(n74819), .Z(n81121) );
  IV U95094 ( .A(n74821), .Z(n74823) );
  NOR U95095 ( .A(n74823), .B(n74822), .Z(n74824) );
  IV U95096 ( .A(n74824), .Z(n80220) );
  IV U95097 ( .A(n74825), .Z(n74827) );
  NOR U95098 ( .A(n74827), .B(n74826), .Z(n80216) );
  NOR U95099 ( .A(n80216), .B(n80213), .Z(n74828) );
  XOR U95100 ( .A(n74829), .B(n74828), .Z(n80219) );
  XOR U95101 ( .A(n80220), .B(n80219), .Z(n74830) );
  NOR U95102 ( .A(n74831), .B(n74830), .Z(n74832) );
  NOR U95103 ( .A(n81121), .B(n74832), .Z(n74839) );
  IV U95104 ( .A(n74839), .Z(n80223) );
  XOR U95105 ( .A(n74838), .B(n80223), .Z(n74833) );
  NOR U95106 ( .A(n74834), .B(n74833), .Z(n81110) );
  IV U95107 ( .A(n74835), .Z(n74836) );
  NOR U95108 ( .A(n74837), .B(n74836), .Z(n75679) );
  NOR U95109 ( .A(n74838), .B(n75679), .Z(n74840) );
  XOR U95110 ( .A(n74840), .B(n74839), .Z(n74845) );
  IV U95111 ( .A(n74845), .Z(n74841) );
  NOR U95112 ( .A(n74842), .B(n74841), .Z(n74843) );
  NOR U95113 ( .A(n81110), .B(n74843), .Z(n74862) );
  NOR U95114 ( .A(n74844), .B(n74862), .Z(n74847) );
  IV U95115 ( .A(n74844), .Z(n74846) );
  NOR U95116 ( .A(n74846), .B(n74845), .Z(n85917) );
  NOR U95117 ( .A(n74847), .B(n85917), .Z(n74858) );
  IV U95118 ( .A(n74850), .Z(n74849) );
  NOR U95119 ( .A(n74849), .B(n74848), .Z(n74857) );
  NOR U95120 ( .A(n74851), .B(n74850), .Z(n74854) );
  IV U95121 ( .A(n74852), .Z(n74853) );
  NOR U95122 ( .A(n74854), .B(n74853), .Z(n74861) );
  NOR U95123 ( .A(n74857), .B(n74861), .Z(n74855) );
  IV U95124 ( .A(n74855), .Z(n74856) );
  NOR U95125 ( .A(n74858), .B(n74856), .Z(n74866) );
  IV U95126 ( .A(n74857), .Z(n74860) );
  IV U95127 ( .A(n74858), .Z(n74859) );
  NOR U95128 ( .A(n74860), .B(n74859), .Z(n85915) );
  IV U95129 ( .A(n74861), .Z(n74864) );
  IV U95130 ( .A(n74862), .Z(n74863) );
  NOR U95131 ( .A(n74864), .B(n74863), .Z(n85921) );
  NOR U95132 ( .A(n85915), .B(n85921), .Z(n74865) );
  IV U95133 ( .A(n74865), .Z(n80238) );
  NOR U95134 ( .A(n74866), .B(n80238), .Z(n74867) );
  IV U95135 ( .A(n74867), .Z(n80235) );
  XOR U95136 ( .A(n80234), .B(n80235), .Z(n75674) );
  XOR U95137 ( .A(n75673), .B(n75674), .Z(n75677) );
  XOR U95138 ( .A(n75676), .B(n75677), .Z(n80245) );
  NOR U95139 ( .A(n74868), .B(n75670), .Z(n74872) );
  IV U95140 ( .A(n74869), .Z(n74871) );
  IV U95141 ( .A(n74870), .Z(n74875) );
  NOR U95142 ( .A(n74871), .B(n74875), .Z(n80243) );
  NOR U95143 ( .A(n74872), .B(n80243), .Z(n74873) );
  XOR U95144 ( .A(n80245), .B(n74873), .Z(n75663) );
  IV U95145 ( .A(n74874), .Z(n74876) );
  NOR U95146 ( .A(n74876), .B(n74875), .Z(n74877) );
  IV U95147 ( .A(n74877), .Z(n75664) );
  XOR U95148 ( .A(n75663), .B(n75664), .Z(n75668) );
  XOR U95149 ( .A(n75666), .B(n75668), .Z(n81093) );
  XOR U95150 ( .A(n75658), .B(n81093), .Z(n75656) );
  IV U95151 ( .A(n74878), .Z(n74880) );
  NOR U95152 ( .A(n74880), .B(n74879), .Z(n75659) );
  NOR U95153 ( .A(n75655), .B(n75659), .Z(n74881) );
  XOR U95154 ( .A(n75656), .B(n74881), .Z(n75651) );
  IV U95155 ( .A(n74882), .Z(n74884) );
  NOR U95156 ( .A(n74884), .B(n74883), .Z(n75649) );
  XOR U95157 ( .A(n75651), .B(n75649), .Z(n75654) );
  XOR U95158 ( .A(n75652), .B(n75654), .Z(n80255) );
  XOR U95159 ( .A(n74885), .B(n80255), .Z(n74886) );
  IV U95160 ( .A(n74886), .Z(n75645) );
  XOR U95161 ( .A(n74887), .B(n75645), .Z(n74890) );
  IV U95162 ( .A(n74890), .Z(n74888) );
  NOR U95163 ( .A(n74889), .B(n74888), .Z(n85944) );
  NOR U95164 ( .A(n74891), .B(n74890), .Z(n80259) );
  NOR U95165 ( .A(n85944), .B(n80259), .Z(n75637) );
  XOR U95166 ( .A(n74892), .B(n75637), .Z(n80263) );
  XOR U95167 ( .A(n80261), .B(n80263), .Z(n80266) );
  IV U95168 ( .A(n74893), .Z(n74894) );
  NOR U95169 ( .A(n74895), .B(n74894), .Z(n80264) );
  XOR U95170 ( .A(n80266), .B(n80264), .Z(n75634) );
  IV U95171 ( .A(n74896), .Z(n74897) );
  NOR U95172 ( .A(n74898), .B(n74897), .Z(n75633) );
  NOR U95173 ( .A(n74899), .B(n75621), .Z(n74900) );
  NOR U95174 ( .A(n75633), .B(n74900), .Z(n74901) );
  XOR U95175 ( .A(n75634), .B(n74901), .Z(n74902) );
  IV U95176 ( .A(n74902), .Z(n75626) );
  XOR U95177 ( .A(n75614), .B(n75626), .Z(n85971) );
  XOR U95178 ( .A(n80274), .B(n85971), .Z(n80279) );
  XOR U95179 ( .A(n80280), .B(n80279), .Z(n80277) );
  XOR U95180 ( .A(n80275), .B(n80277), .Z(n75609) );
  XOR U95181 ( .A(n75608), .B(n75609), .Z(n80288) );
  XOR U95182 ( .A(n75611), .B(n80288), .Z(n75603) );
  XOR U95183 ( .A(n74903), .B(n75603), .Z(n75598) );
  XOR U95184 ( .A(n74904), .B(n75598), .Z(n75596) );
  XOR U95185 ( .A(n74905), .B(n75596), .Z(n74906) );
  IV U95186 ( .A(n74906), .Z(n80297) );
  XOR U95187 ( .A(n80296), .B(n80297), .Z(n75590) );
  IV U95188 ( .A(n74907), .Z(n74908) );
  NOR U95189 ( .A(n74909), .B(n74908), .Z(n75589) );
  NOR U95190 ( .A(n74910), .B(n75585), .Z(n74911) );
  NOR U95191 ( .A(n75589), .B(n74911), .Z(n74912) );
  XOR U95192 ( .A(n75590), .B(n74912), .Z(n74913) );
  IV U95193 ( .A(n74913), .Z(n80311) );
  IV U95194 ( .A(n74914), .Z(n74916) );
  NOR U95195 ( .A(n74916), .B(n74915), .Z(n74917) );
  IV U95196 ( .A(n74917), .Z(n74924) );
  NOR U95197 ( .A(n80311), .B(n74924), .Z(n81007) );
  IV U95198 ( .A(n74918), .Z(n74920) );
  IV U95199 ( .A(n74919), .Z(n74922) );
  NOR U95200 ( .A(n74920), .B(n74922), .Z(n80312) );
  IV U95201 ( .A(n74921), .Z(n74923) );
  NOR U95202 ( .A(n74923), .B(n74922), .Z(n80309) );
  XOR U95203 ( .A(n80309), .B(n80311), .Z(n80313) );
  IV U95204 ( .A(n80313), .Z(n74925) );
  XOR U95205 ( .A(n80312), .B(n74925), .Z(n74927) );
  NOR U95206 ( .A(n74925), .B(n74924), .Z(n74926) );
  NOR U95207 ( .A(n74927), .B(n74926), .Z(n74928) );
  NOR U95208 ( .A(n81007), .B(n74928), .Z(n74929) );
  IV U95209 ( .A(n74929), .Z(n80318) );
  IV U95210 ( .A(n74930), .Z(n74931) );
  NOR U95211 ( .A(n74932), .B(n74931), .Z(n80316) );
  XOR U95212 ( .A(n80318), .B(n80316), .Z(n80328) );
  XOR U95213 ( .A(n80320), .B(n80328), .Z(n80323) );
  XOR U95214 ( .A(n74933), .B(n80323), .Z(n74934) );
  IV U95215 ( .A(n74934), .Z(n80331) );
  XOR U95216 ( .A(n80329), .B(n80331), .Z(n80333) );
  XOR U95217 ( .A(n80332), .B(n80333), .Z(n75582) );
  XOR U95218 ( .A(n75581), .B(n75582), .Z(n75578) );
  IV U95219 ( .A(n74935), .Z(n74937) );
  NOR U95220 ( .A(n74937), .B(n74936), .Z(n75575) );
  NOR U95221 ( .A(n75577), .B(n75575), .Z(n74938) );
  XOR U95222 ( .A(n75578), .B(n74938), .Z(n75564) );
  XOR U95223 ( .A(n74939), .B(n75564), .Z(n80345) );
  XOR U95224 ( .A(n74940), .B(n80345), .Z(n80347) );
  XOR U95225 ( .A(n80348), .B(n80347), .Z(n80355) );
  IV U95226 ( .A(n74941), .Z(n74942) );
  NOR U95227 ( .A(n74943), .B(n74942), .Z(n80354) );
  NOR U95228 ( .A(n80349), .B(n80354), .Z(n74944) );
  XOR U95229 ( .A(n80355), .B(n74944), .Z(n74945) );
  IV U95230 ( .A(n74945), .Z(n75557) );
  NOR U95231 ( .A(n74946), .B(n75556), .Z(n74950) );
  IV U95232 ( .A(n74947), .Z(n74949) );
  IV U95233 ( .A(n74948), .Z(n74953) );
  NOR U95234 ( .A(n74949), .B(n74953), .Z(n75553) );
  NOR U95235 ( .A(n74950), .B(n75553), .Z(n74951) );
  XOR U95236 ( .A(n75557), .B(n74951), .Z(n75548) );
  IV U95237 ( .A(n74952), .Z(n74954) );
  NOR U95238 ( .A(n74954), .B(n74953), .Z(n75550) );
  IV U95239 ( .A(n74955), .Z(n74956) );
  NOR U95240 ( .A(n74956), .B(n74959), .Z(n75547) );
  NOR U95241 ( .A(n75550), .B(n75547), .Z(n74957) );
  XOR U95242 ( .A(n75548), .B(n74957), .Z(n75543) );
  IV U95243 ( .A(n74958), .Z(n74960) );
  NOR U95244 ( .A(n74960), .B(n74959), .Z(n75541) );
  XOR U95245 ( .A(n75543), .B(n75541), .Z(n75546) );
  XOR U95246 ( .A(n75544), .B(n75546), .Z(n75538) );
  XOR U95247 ( .A(n74961), .B(n75538), .Z(n74962) );
  IV U95248 ( .A(n74962), .Z(n75529) );
  XOR U95249 ( .A(n74963), .B(n75529), .Z(n75515) );
  XOR U95250 ( .A(n74964), .B(n75515), .Z(n75510) );
  IV U95251 ( .A(n74965), .Z(n74967) );
  NOR U95252 ( .A(n74967), .B(n74966), .Z(n75513) );
  IV U95253 ( .A(n74968), .Z(n74969) );
  NOR U95254 ( .A(n74969), .B(n74972), .Z(n75508) );
  NOR U95255 ( .A(n75513), .B(n75508), .Z(n74970) );
  XOR U95256 ( .A(n75510), .B(n74970), .Z(n80362) );
  IV U95257 ( .A(n74971), .Z(n74973) );
  NOR U95258 ( .A(n74973), .B(n74972), .Z(n74974) );
  IV U95259 ( .A(n74974), .Z(n80363) );
  XOR U95260 ( .A(n80362), .B(n80363), .Z(n75507) );
  XOR U95261 ( .A(n75505), .B(n75507), .Z(n74978) );
  IV U95262 ( .A(n74975), .Z(n74976) );
  NOR U95263 ( .A(n74981), .B(n74976), .Z(n74984) );
  IV U95264 ( .A(n74984), .Z(n74977) );
  NOR U95265 ( .A(n74978), .B(n74977), .Z(n80942) );
  IV U95266 ( .A(n74979), .Z(n74980) );
  NOR U95267 ( .A(n74981), .B(n74980), .Z(n75502) );
  NOR U95268 ( .A(n75505), .B(n75502), .Z(n74982) );
  XOR U95269 ( .A(n75507), .B(n74982), .Z(n74983) );
  NOR U95270 ( .A(n74984), .B(n74983), .Z(n74985) );
  NOR U95271 ( .A(n80942), .B(n74985), .Z(n80373) );
  XOR U95272 ( .A(n74986), .B(n80373), .Z(n80384) );
  XOR U95273 ( .A(n80376), .B(n80384), .Z(n75500) );
  IV U95274 ( .A(n75500), .Z(n74993) );
  IV U95275 ( .A(n74987), .Z(n74988) );
  NOR U95276 ( .A(n74989), .B(n74988), .Z(n74991) );
  NOR U95277 ( .A(n74991), .B(n74990), .Z(n74992) );
  XOR U95278 ( .A(n74993), .B(n74992), .Z(n80390) );
  IV U95279 ( .A(n74994), .Z(n74996) );
  IV U95280 ( .A(n74995), .Z(n75493) );
  NOR U95281 ( .A(n74996), .B(n75493), .Z(n80388) );
  XOR U95282 ( .A(n80390), .B(n80388), .Z(n80392) );
  NOR U95283 ( .A(n75003), .B(n80392), .Z(n86080) );
  IV U95284 ( .A(n74997), .Z(n74999) );
  NOR U95285 ( .A(n74999), .B(n74998), .Z(n75485) );
  IV U95286 ( .A(n75000), .Z(n75001) );
  NOR U95287 ( .A(n75002), .B(n75001), .Z(n80391) );
  XOR U95288 ( .A(n80391), .B(n80392), .Z(n75486) );
  IV U95289 ( .A(n75486), .Z(n75004) );
  XOR U95290 ( .A(n75485), .B(n75004), .Z(n75006) );
  NOR U95291 ( .A(n75004), .B(n75003), .Z(n75005) );
  NOR U95292 ( .A(n75006), .B(n75005), .Z(n75007) );
  NOR U95293 ( .A(n86080), .B(n75007), .Z(n75489) );
  XOR U95294 ( .A(n75488), .B(n75489), .Z(n75482) );
  IV U95295 ( .A(n75008), .Z(n75010) );
  NOR U95296 ( .A(n75010), .B(n75009), .Z(n80397) );
  IV U95297 ( .A(n75015), .Z(n75011) );
  NOR U95298 ( .A(n75011), .B(n75014), .Z(n75481) );
  NOR U95299 ( .A(n80397), .B(n75481), .Z(n75012) );
  XOR U95300 ( .A(n75482), .B(n75012), .Z(n75480) );
  IV U95301 ( .A(n75013), .Z(n75016) );
  NOR U95302 ( .A(n75016), .B(n75014), .Z(n75027) );
  XOR U95303 ( .A(n75015), .B(n75017), .Z(n75019) );
  NOR U95304 ( .A(n75017), .B(n75016), .Z(n75018) );
  NOR U95305 ( .A(n75019), .B(n75018), .Z(n75025) );
  IV U95306 ( .A(n75020), .Z(n75021) );
  NOR U95307 ( .A(n75022), .B(n75021), .Z(n75023) );
  IV U95308 ( .A(n75023), .Z(n75024) );
  NOR U95309 ( .A(n75025), .B(n75024), .Z(n75026) );
  NOR U95310 ( .A(n75027), .B(n75026), .Z(n75479) );
  XOR U95311 ( .A(n75480), .B(n75479), .Z(n75028) );
  NOR U95312 ( .A(n75033), .B(n75028), .Z(n75035) );
  IV U95313 ( .A(n75029), .Z(n75031) );
  NOR U95314 ( .A(n75031), .B(n75030), .Z(n75036) );
  IV U95315 ( .A(n75036), .Z(n75032) );
  NOR U95316 ( .A(n75035), .B(n75032), .Z(n80911) );
  IV U95317 ( .A(n75033), .Z(n75034) );
  NOR U95318 ( .A(n75480), .B(n75034), .Z(n80918) );
  NOR U95319 ( .A(n80918), .B(n75035), .Z(n75039) );
  NOR U95320 ( .A(n75036), .B(n75039), .Z(n75037) );
  NOR U95321 ( .A(n80911), .B(n75037), .Z(n75038) );
  NOR U95322 ( .A(n75040), .B(n75038), .Z(n75043) );
  IV U95323 ( .A(n75039), .Z(n75042) );
  IV U95324 ( .A(n75040), .Z(n75041) );
  NOR U95325 ( .A(n75042), .B(n75041), .Z(n80909) );
  NOR U95326 ( .A(n75043), .B(n80909), .Z(n75471) );
  XOR U95327 ( .A(n75044), .B(n75471), .Z(n75474) );
  XOR U95328 ( .A(n75473), .B(n75474), .Z(n86107) );
  IV U95329 ( .A(n86107), .Z(n75051) );
  IV U95330 ( .A(n75045), .Z(n75047) );
  NOR U95331 ( .A(n75047), .B(n75046), .Z(n86105) );
  IV U95332 ( .A(n75048), .Z(n75050) );
  NOR U95333 ( .A(n75050), .B(n75049), .Z(n86110) );
  NOR U95334 ( .A(n86105), .B(n86110), .Z(n80403) );
  XOR U95335 ( .A(n75051), .B(n80403), .Z(n80408) );
  XOR U95336 ( .A(n80404), .B(n80408), .Z(n86115) );
  XOR U95337 ( .A(n86116), .B(n86115), .Z(n75052) );
  IV U95338 ( .A(n75052), .Z(n80415) );
  XOR U95339 ( .A(n80414), .B(n80415), .Z(n80419) );
  IV U95340 ( .A(n75053), .Z(n75055) );
  NOR U95341 ( .A(n75055), .B(n75054), .Z(n80417) );
  XOR U95342 ( .A(n80419), .B(n80417), .Z(n75463) );
  XOR U95343 ( .A(n75464), .B(n75463), .Z(n75465) );
  IV U95344 ( .A(n75056), .Z(n75066) );
  IV U95345 ( .A(n75058), .Z(n75057) );
  NOR U95346 ( .A(n75066), .B(n75057), .Z(n86132) );
  XOR U95347 ( .A(n75066), .B(n75058), .Z(n75061) );
  IV U95348 ( .A(n75059), .Z(n75060) );
  NOR U95349 ( .A(n75061), .B(n75060), .Z(n86141) );
  NOR U95350 ( .A(n86132), .B(n86141), .Z(n75466) );
  XOR U95351 ( .A(n75465), .B(n75466), .Z(n86138) );
  IV U95352 ( .A(n75062), .Z(n75063) );
  NOR U95353 ( .A(n75063), .B(n75068), .Z(n75457) );
  IV U95354 ( .A(n75064), .Z(n75065) );
  NOR U95355 ( .A(n75066), .B(n75065), .Z(n86137) );
  IV U95356 ( .A(n75067), .Z(n75069) );
  NOR U95357 ( .A(n75069), .B(n75068), .Z(n86148) );
  NOR U95358 ( .A(n86137), .B(n86148), .Z(n75461) );
  IV U95359 ( .A(n75461), .Z(n75073) );
  NOR U95360 ( .A(n75457), .B(n75073), .Z(n75070) );
  XOR U95361 ( .A(n86138), .B(n75070), .Z(n75079) );
  NOR U95362 ( .A(n75071), .B(n75079), .Z(n75087) );
  IV U95363 ( .A(n75072), .Z(n75075) );
  XOR U95364 ( .A(n86138), .B(n75073), .Z(n75074) );
  NOR U95365 ( .A(n75075), .B(n75074), .Z(n75076) );
  IV U95366 ( .A(n75076), .Z(n75077) );
  NOR U95367 ( .A(n75081), .B(n75077), .Z(n75459) );
  IV U95368 ( .A(n75078), .Z(n75084) );
  IV U95369 ( .A(n75079), .Z(n75080) );
  NOR U95370 ( .A(n75081), .B(n75080), .Z(n75082) );
  IV U95371 ( .A(n75082), .Z(n75083) );
  NOR U95372 ( .A(n75084), .B(n75083), .Z(n75456) );
  NOR U95373 ( .A(n75459), .B(n75456), .Z(n75085) );
  IV U95374 ( .A(n75085), .Z(n75086) );
  NOR U95375 ( .A(n75087), .B(n75086), .Z(n80423) );
  XOR U95376 ( .A(n80424), .B(n80423), .Z(n80433) );
  IV U95377 ( .A(n75088), .Z(n75089) );
  NOR U95378 ( .A(n75090), .B(n75089), .Z(n80425) );
  NOR U95379 ( .A(n75092), .B(n75091), .Z(n80432) );
  NOR U95380 ( .A(n80425), .B(n80432), .Z(n75093) );
  XOR U95381 ( .A(n80433), .B(n75093), .Z(n75094) );
  IV U95382 ( .A(n75094), .Z(n80431) );
  XOR U95383 ( .A(n80429), .B(n80431), .Z(n75454) );
  XOR U95384 ( .A(n75095), .B(n75454), .Z(n80439) );
  IV U95385 ( .A(n75096), .Z(n75098) );
  NOR U95386 ( .A(n75098), .B(n75097), .Z(n75449) );
  IV U95387 ( .A(n75099), .Z(n75101) );
  NOR U95388 ( .A(n75101), .B(n75100), .Z(n80438) );
  NOR U95389 ( .A(n75449), .B(n80438), .Z(n75102) );
  XOR U95390 ( .A(n80439), .B(n75102), .Z(n75447) );
  XOR U95391 ( .A(n75442), .B(n75447), .Z(n75103) );
  XOR U95392 ( .A(n75104), .B(n75103), .Z(n75441) );
  XOR U95393 ( .A(n75440), .B(n75441), .Z(n75431) );
  IV U95394 ( .A(n75105), .Z(n75107) );
  NOR U95395 ( .A(n75107), .B(n75106), .Z(n75438) );
  IV U95396 ( .A(n75108), .Z(n75109) );
  NOR U95397 ( .A(n75110), .B(n75109), .Z(n75430) );
  NOR U95398 ( .A(n75438), .B(n75430), .Z(n75111) );
  XOR U95399 ( .A(n75431), .B(n75111), .Z(n80445) );
  XOR U95400 ( .A(n75119), .B(n80445), .Z(n75115) );
  IV U95401 ( .A(n75112), .Z(n75113) );
  NOR U95402 ( .A(n75113), .B(n75128), .Z(n75122) );
  IV U95403 ( .A(n75122), .Z(n75114) );
  NOR U95404 ( .A(n75115), .B(n75114), .Z(n86198) );
  IV U95405 ( .A(n75116), .Z(n75118) );
  NOR U95406 ( .A(n75118), .B(n75117), .Z(n80443) );
  NOR U95407 ( .A(n75119), .B(n80443), .Z(n75120) );
  XOR U95408 ( .A(n80445), .B(n75120), .Z(n75121) );
  NOR U95409 ( .A(n75122), .B(n75121), .Z(n75123) );
  NOR U95410 ( .A(n86198), .B(n75123), .Z(n75420) );
  IV U95411 ( .A(n75124), .Z(n75125) );
  NOR U95412 ( .A(n75125), .B(n75128), .Z(n75126) );
  IV U95413 ( .A(n75126), .Z(n75421) );
  XOR U95414 ( .A(n75420), .B(n75421), .Z(n75425) );
  IV U95415 ( .A(n75127), .Z(n75129) );
  NOR U95416 ( .A(n75129), .B(n75128), .Z(n75423) );
  XOR U95417 ( .A(n75425), .B(n75423), .Z(n75135) );
  IV U95418 ( .A(n75135), .Z(n75130) );
  NOR U95419 ( .A(n75131), .B(n75130), .Z(n75138) );
  IV U95420 ( .A(n75132), .Z(n75133) );
  NOR U95421 ( .A(n75133), .B(n75425), .Z(n80847) );
  IV U95422 ( .A(n75134), .Z(n75136) );
  NOR U95423 ( .A(n75136), .B(n75135), .Z(n80844) );
  NOR U95424 ( .A(n80847), .B(n80844), .Z(n75137) );
  IV U95425 ( .A(n75137), .Z(n75419) );
  NOR U95426 ( .A(n75138), .B(n75419), .Z(n75139) );
  IV U95427 ( .A(n75139), .Z(n75417) );
  IV U95428 ( .A(n75140), .Z(n75142) );
  NOR U95429 ( .A(n75142), .B(n75141), .Z(n75416) );
  NOR U95430 ( .A(n75416), .B(n75414), .Z(n75143) );
  XOR U95431 ( .A(n75417), .B(n75143), .Z(n75149) );
  IV U95432 ( .A(n75149), .Z(n75148) );
  IV U95433 ( .A(n75144), .Z(n75146) );
  NOR U95434 ( .A(n75146), .B(n75145), .Z(n75150) );
  IV U95435 ( .A(n75150), .Z(n75147) );
  NOR U95436 ( .A(n75148), .B(n75147), .Z(n86201) );
  NOR U95437 ( .A(n75150), .B(n75149), .Z(n80454) );
  IV U95438 ( .A(n75151), .Z(n75153) );
  NOR U95439 ( .A(n75153), .B(n75152), .Z(n80452) );
  XOR U95440 ( .A(n80454), .B(n80452), .Z(n75154) );
  NOR U95441 ( .A(n86201), .B(n75154), .Z(n80450) );
  IV U95442 ( .A(n75155), .Z(n75157) );
  NOR U95443 ( .A(n75157), .B(n75156), .Z(n80449) );
  IV U95444 ( .A(n75158), .Z(n75159) );
  NOR U95445 ( .A(n75160), .B(n75159), .Z(n80460) );
  NOR U95446 ( .A(n80449), .B(n80460), .Z(n75161) );
  XOR U95447 ( .A(n80450), .B(n75161), .Z(n80466) );
  IV U95448 ( .A(n75162), .Z(n75163) );
  NOR U95449 ( .A(n75164), .B(n75163), .Z(n80458) );
  IV U95450 ( .A(n75165), .Z(n75166) );
  NOR U95451 ( .A(n75167), .B(n75166), .Z(n80464) );
  NOR U95452 ( .A(n80458), .B(n80464), .Z(n75168) );
  XOR U95453 ( .A(n80466), .B(n75168), .Z(n75169) );
  IV U95454 ( .A(n75169), .Z(n80471) );
  IV U95455 ( .A(n75170), .Z(n75172) );
  NOR U95456 ( .A(n75172), .B(n75171), .Z(n80467) );
  NOR U95457 ( .A(n75173), .B(n80472), .Z(n75174) );
  NOR U95458 ( .A(n80467), .B(n75174), .Z(n75175) );
  XOR U95459 ( .A(n80471), .B(n75175), .Z(n75408) );
  IV U95460 ( .A(n75176), .Z(n75177) );
  NOR U95461 ( .A(n75179), .B(n75177), .Z(n75411) );
  IV U95462 ( .A(n75178), .Z(n75182) );
  NOR U95463 ( .A(n75180), .B(n75179), .Z(n75181) );
  IV U95464 ( .A(n75181), .Z(n75185) );
  NOR U95465 ( .A(n75182), .B(n75185), .Z(n75409) );
  NOR U95466 ( .A(n75411), .B(n75409), .Z(n75183) );
  XOR U95467 ( .A(n75408), .B(n75183), .Z(n80483) );
  IV U95468 ( .A(n75184), .Z(n75186) );
  NOR U95469 ( .A(n75186), .B(n75185), .Z(n80481) );
  XOR U95470 ( .A(n80483), .B(n80481), .Z(n80495) );
  IV U95471 ( .A(n75187), .Z(n75189) );
  NOR U95472 ( .A(n75189), .B(n75188), .Z(n75190) );
  IV U95473 ( .A(n75190), .Z(n80493) );
  XOR U95474 ( .A(n80495), .B(n80493), .Z(n75191) );
  XOR U95475 ( .A(n75192), .B(n75191), .Z(n75403) );
  IV U95476 ( .A(n75193), .Z(n75194) );
  NOR U95477 ( .A(n75194), .B(n75199), .Z(n75402) );
  IV U95478 ( .A(n75195), .Z(n75196) );
  NOR U95479 ( .A(n80496), .B(n75196), .Z(n75405) );
  NOR U95480 ( .A(n75402), .B(n75405), .Z(n75197) );
  XOR U95481 ( .A(n75403), .B(n75197), .Z(n75401) );
  IV U95482 ( .A(n75198), .Z(n75200) );
  NOR U95483 ( .A(n75200), .B(n75199), .Z(n75399) );
  XOR U95484 ( .A(n75401), .B(n75399), .Z(n75395) );
  XOR U95485 ( .A(n75393), .B(n75395), .Z(n75398) );
  XOR U95486 ( .A(n75396), .B(n75398), .Z(n75389) );
  XOR U95487 ( .A(n75388), .B(n75389), .Z(n80507) );
  XOR U95488 ( .A(n75201), .B(n80507), .Z(n80510) );
  IV U95489 ( .A(n75202), .Z(n75203) );
  NOR U95490 ( .A(n75203), .B(n75206), .Z(n80513) );
  IV U95491 ( .A(n75204), .Z(n75205) );
  NOR U95492 ( .A(n75206), .B(n75205), .Z(n80509) );
  NOR U95493 ( .A(n80513), .B(n80509), .Z(n75207) );
  XOR U95494 ( .A(n80510), .B(n75207), .Z(n75384) );
  IV U95495 ( .A(n75208), .Z(n75210) );
  NOR U95496 ( .A(n75210), .B(n75209), .Z(n75380) );
  NOR U95497 ( .A(n75382), .B(n75380), .Z(n75211) );
  XOR U95498 ( .A(n75384), .B(n75211), .Z(n75375) );
  IV U95499 ( .A(n75212), .Z(n75214) );
  NOR U95500 ( .A(n75214), .B(n75213), .Z(n75377) );
  IV U95501 ( .A(n75215), .Z(n75217) );
  NOR U95502 ( .A(n75217), .B(n75216), .Z(n75374) );
  NOR U95503 ( .A(n75377), .B(n75374), .Z(n75218) );
  XOR U95504 ( .A(n75375), .B(n75218), .Z(n80523) );
  XOR U95505 ( .A(n75219), .B(n80523), .Z(n75220) );
  IV U95506 ( .A(n75220), .Z(n80521) );
  XOR U95507 ( .A(n75221), .B(n80521), .Z(n75228) );
  IV U95508 ( .A(n75228), .Z(n75222) );
  NOR U95509 ( .A(n75223), .B(n75222), .Z(n80776) );
  IV U95510 ( .A(n75224), .Z(n75226) );
  NOR U95511 ( .A(n75226), .B(n75225), .Z(n75229) );
  IV U95512 ( .A(n75229), .Z(n75227) );
  NOR U95513 ( .A(n80521), .B(n75227), .Z(n86274) );
  NOR U95514 ( .A(n75229), .B(n75228), .Z(n75230) );
  NOR U95515 ( .A(n86274), .B(n75230), .Z(n75231) );
  NOR U95516 ( .A(n75232), .B(n75231), .Z(n75233) );
  NOR U95517 ( .A(n80776), .B(n75233), .Z(n75234) );
  IV U95518 ( .A(n75234), .Z(n80771) );
  XOR U95519 ( .A(n80770), .B(n80771), .Z(n75365) );
  XOR U95520 ( .A(n75235), .B(n75365), .Z(n75363) );
  IV U95521 ( .A(n75236), .Z(n75238) );
  NOR U95522 ( .A(n75238), .B(n75237), .Z(n75361) );
  IV U95523 ( .A(n75239), .Z(n75240) );
  NOR U95524 ( .A(n75241), .B(n75240), .Z(n75356) );
  NOR U95525 ( .A(n75361), .B(n75356), .Z(n75242) );
  XOR U95526 ( .A(n75363), .B(n75242), .Z(n75354) );
  NOR U95527 ( .A(n86472), .B(n80756), .Z(n75358) );
  IV U95528 ( .A(n75243), .Z(n75244) );
  NOR U95529 ( .A(n75245), .B(n75244), .Z(n75353) );
  NOR U95530 ( .A(n75358), .B(n75353), .Z(n75246) );
  XOR U95531 ( .A(n75354), .B(n75246), .Z(n80535) );
  XOR U95532 ( .A(n75247), .B(n80535), .Z(n75248) );
  XOR U95533 ( .A(n80533), .B(n75248), .Z(n80736) );
  XOR U95534 ( .A(n80546), .B(n80736), .Z(n80547) );
  IV U95535 ( .A(n75249), .Z(n75250) );
  NOR U95536 ( .A(n75251), .B(n75250), .Z(n75256) );
  IV U95537 ( .A(n75252), .Z(n75254) );
  NOR U95538 ( .A(n75254), .B(n75253), .Z(n75255) );
  NOR U95539 ( .A(n75256), .B(n75255), .Z(n80549) );
  XOR U95540 ( .A(n80547), .B(n80549), .Z(n80555) );
  IV U95541 ( .A(n75257), .Z(n75258) );
  NOR U95542 ( .A(n75259), .B(n75258), .Z(n80554) );
  IV U95543 ( .A(n75260), .Z(n75261) );
  NOR U95544 ( .A(n75262), .B(n75261), .Z(n80552) );
  NOR U95545 ( .A(n80554), .B(n80552), .Z(n75263) );
  XOR U95546 ( .A(n80555), .B(n75263), .Z(n75264) );
  NOR U95547 ( .A(n75265), .B(n75264), .Z(n75268) );
  XOR U95548 ( .A(n80554), .B(n80555), .Z(n75267) );
  IV U95549 ( .A(n75265), .Z(n75266) );
  NOR U95550 ( .A(n75267), .B(n75266), .Z(n86290) );
  NOR U95551 ( .A(n75268), .B(n86290), .Z(n80558) );
  IV U95552 ( .A(n75269), .Z(n75278) );
  IV U95553 ( .A(n75270), .Z(n75271) );
  NOR U95554 ( .A(n75278), .B(n75271), .Z(n80562) );
  IV U95555 ( .A(n75272), .Z(n75274) );
  NOR U95556 ( .A(n75274), .B(n75273), .Z(n80559) );
  NOR U95557 ( .A(n80562), .B(n80559), .Z(n75275) );
  XOR U95558 ( .A(n80558), .B(n75275), .Z(n80569) );
  IV U95559 ( .A(n75276), .Z(n75277) );
  NOR U95560 ( .A(n75278), .B(n75277), .Z(n75279) );
  IV U95561 ( .A(n75279), .Z(n80568) );
  XOR U95562 ( .A(n80569), .B(n80568), .Z(n75287) );
  XOR U95563 ( .A(n75346), .B(n75287), .Z(n75285) );
  IV U95564 ( .A(n75280), .Z(n75282) );
  NOR U95565 ( .A(n75282), .B(n75281), .Z(n75283) );
  IV U95566 ( .A(n75283), .Z(n75288) );
  NOR U95567 ( .A(n75287), .B(n75288), .Z(n75284) );
  NOR U95568 ( .A(n75285), .B(n75284), .Z(n80703) );
  NOR U95569 ( .A(n75286), .B(n80703), .Z(n80577) );
  IV U95570 ( .A(n75287), .Z(n75347) );
  NOR U95571 ( .A(n75288), .B(n75347), .Z(n80718) );
  NOR U95572 ( .A(n80718), .B(n80703), .Z(n75293) );
  NOR U95573 ( .A(n75289), .B(n75293), .Z(n75290) );
  NOR U95574 ( .A(n80577), .B(n75290), .Z(n75291) );
  NOR U95575 ( .A(n75292), .B(n75291), .Z(n75298) );
  IV U95576 ( .A(n75293), .Z(n75294) );
  NOR U95577 ( .A(n75295), .B(n75294), .Z(n75296) );
  IV U95578 ( .A(n75296), .Z(n80585) );
  NOR U95579 ( .A(n75297), .B(n80585), .Z(n80579) );
  NOR U95580 ( .A(n75298), .B(n80579), .Z(n80591) );
  IV U95581 ( .A(n75299), .Z(n75301) );
  NOR U95582 ( .A(n75301), .B(n75300), .Z(n86307) );
  IV U95583 ( .A(n75302), .Z(n75304) );
  NOR U95584 ( .A(n75304), .B(n75303), .Z(n80697) );
  NOR U95585 ( .A(n86307), .B(n80697), .Z(n80592) );
  XOR U95586 ( .A(n80591), .B(n80592), .Z(n80594) );
  XOR U95587 ( .A(n75305), .B(n80594), .Z(n80599) );
  XOR U95588 ( .A(n75306), .B(n80599), .Z(n80622) );
  NOR U95589 ( .A(n75307), .B(n80622), .Z(n80686) );
  IV U95590 ( .A(n75308), .Z(n75309) );
  NOR U95591 ( .A(n75312), .B(n75309), .Z(n80618) );
  IV U95592 ( .A(n75310), .Z(n75311) );
  NOR U95593 ( .A(n75312), .B(n75311), .Z(n80621) );
  XOR U95594 ( .A(n80621), .B(n80622), .Z(n80619) );
  XOR U95595 ( .A(n80618), .B(n80619), .Z(n80629) );
  IV U95596 ( .A(n80629), .Z(n75313) );
  NOR U95597 ( .A(n75314), .B(n75313), .Z(n75315) );
  NOR U95598 ( .A(n80686), .B(n75315), .Z(n75340) );
  XOR U95599 ( .A(n75316), .B(n75340), .Z(n80637) );
  XOR U95600 ( .A(n75317), .B(n80637), .Z(n80666) );
  XOR U95601 ( .A(n80664), .B(n80666), .Z(n80661) );
  XOR U95602 ( .A(n75319), .B(n75318), .Z(n86361) );
  IV U95603 ( .A(n75320), .Z(n75322) );
  NOR U95604 ( .A(n75322), .B(n75321), .Z(n80649) );
  IV U95605 ( .A(n80649), .Z(n75323) );
  NOR U95606 ( .A(n75324), .B(n75323), .Z(n80644) );
  IV U95607 ( .A(n80644), .Z(n75329) );
  NOR U95608 ( .A(n75326), .B(n75325), .Z(n75328) );
  XOR U95609 ( .A(n75328), .B(n75327), .Z(n80643) );
  NOR U95610 ( .A(n75329), .B(n80643), .Z(n86359) );
  IV U95611 ( .A(n86359), .Z(n75330) );
  NOR U95612 ( .A(n86361), .B(n75330), .Z(n80639) );
  IV U95613 ( .A(n80639), .Z(n75331) );
  NOR U95614 ( .A(n75332), .B(n75331), .Z(n80662) );
  IV U95615 ( .A(n80662), .Z(n75333) );
  NOR U95616 ( .A(n80661), .B(n75333), .Z(n86352) );
  IV U95617 ( .A(n86352), .Z(n80667) );
  IV U95618 ( .A(n75334), .Z(n75337) );
  NOR U95619 ( .A(n80637), .B(n75335), .Z(n75336) );
  IV U95620 ( .A(n75336), .Z(n80633) );
  NOR U95621 ( .A(n75337), .B(n80633), .Z(n75338) );
  IV U95622 ( .A(n75338), .Z(n80675) );
  IV U95623 ( .A(n75339), .Z(n75342) );
  IV U95624 ( .A(n75340), .Z(n75341) );
  NOR U95625 ( .A(n75342), .B(n75341), .Z(n75343) );
  IV U95626 ( .A(n75343), .Z(n86342) );
  IV U95627 ( .A(n75344), .Z(n75345) );
  NOR U95628 ( .A(n75345), .B(n80594), .Z(n80694) );
  IV U95629 ( .A(n75346), .Z(n75348) );
  NOR U95630 ( .A(n75348), .B(n75347), .Z(n80574) );
  IV U95631 ( .A(n80574), .Z(n80567) );
  IV U95632 ( .A(n75349), .Z(n75352) );
  NOR U95633 ( .A(n75350), .B(n80535), .Z(n75351) );
  IV U95634 ( .A(n75351), .Z(n80538) );
  NOR U95635 ( .A(n75352), .B(n80538), .Z(n80740) );
  IV U95636 ( .A(n75353), .Z(n75355) );
  IV U95637 ( .A(n75354), .Z(n80753) );
  NOR U95638 ( .A(n75355), .B(n80753), .Z(n80744) );
  IV U95639 ( .A(n75356), .Z(n75357) );
  NOR U95640 ( .A(n75363), .B(n75357), .Z(n80761) );
  IV U95641 ( .A(n75358), .Z(n75359) );
  NOR U95642 ( .A(n75359), .B(n80753), .Z(n75360) );
  NOR U95643 ( .A(n80761), .B(n75360), .Z(n80532) );
  IV U95644 ( .A(n75361), .Z(n75362) );
  NOR U95645 ( .A(n75363), .B(n75362), .Z(n80764) );
  IV U95646 ( .A(n75364), .Z(n75366) );
  NOR U95647 ( .A(n75366), .B(n75365), .Z(n75367) );
  NOR U95648 ( .A(n80764), .B(n75367), .Z(n80531) );
  NOR U95649 ( .A(n80770), .B(n75368), .Z(n75369) );
  NOR U95650 ( .A(n80771), .B(n75369), .Z(n80530) );
  IV U95651 ( .A(n75370), .Z(n75371) );
  NOR U95652 ( .A(n80521), .B(n75371), .Z(n86262) );
  NOR U95653 ( .A(n80776), .B(n86262), .Z(n80528) );
  IV U95654 ( .A(n75372), .Z(n75373) );
  NOR U95655 ( .A(n75373), .B(n80523), .Z(n80781) );
  IV U95656 ( .A(n75374), .Z(n75376) );
  IV U95657 ( .A(n75375), .Z(n75378) );
  NOR U95658 ( .A(n75376), .B(n75378), .Z(n80778) );
  IV U95659 ( .A(n75377), .Z(n75379) );
  NOR U95660 ( .A(n75379), .B(n75378), .Z(n80786) );
  IV U95661 ( .A(n75380), .Z(n75381) );
  NOR U95662 ( .A(n75384), .B(n75381), .Z(n80788) );
  NOR U95663 ( .A(n80786), .B(n80788), .Z(n80517) );
  IV U95664 ( .A(n75382), .Z(n75383) );
  NOR U95665 ( .A(n75384), .B(n75383), .Z(n86255) );
  XOR U95666 ( .A(n75391), .B(n80507), .Z(n75387) );
  IV U95667 ( .A(n75385), .Z(n75386) );
  NOR U95668 ( .A(n75387), .B(n75386), .Z(n80797) );
  IV U95669 ( .A(n75388), .Z(n75390) );
  NOR U95670 ( .A(n75390), .B(n75389), .Z(n80807) );
  IV U95671 ( .A(n75391), .Z(n75392) );
  NOR U95672 ( .A(n80507), .B(n75392), .Z(n80803) );
  NOR U95673 ( .A(n80807), .B(n80803), .Z(n80505) );
  IV U95674 ( .A(n75393), .Z(n75394) );
  NOR U95675 ( .A(n75395), .B(n75394), .Z(n86234) );
  IV U95676 ( .A(n75396), .Z(n75397) );
  NOR U95677 ( .A(n75398), .B(n75397), .Z(n80809) );
  NOR U95678 ( .A(n86234), .B(n80809), .Z(n80504) );
  IV U95679 ( .A(n75399), .Z(n75400) );
  NOR U95680 ( .A(n75401), .B(n75400), .Z(n80811) );
  IV U95681 ( .A(n75402), .Z(n75404) );
  IV U95682 ( .A(n75403), .Z(n75406) );
  NOR U95683 ( .A(n75404), .B(n75406), .Z(n86230) );
  NOR U95684 ( .A(n80811), .B(n86230), .Z(n80503) );
  IV U95685 ( .A(n75405), .Z(n75407) );
  NOR U95686 ( .A(n75407), .B(n75406), .Z(n80814) );
  IV U95687 ( .A(n75408), .Z(n75413) );
  IV U95688 ( .A(n75409), .Z(n75410) );
  NOR U95689 ( .A(n75413), .B(n75410), .Z(n80485) );
  IV U95690 ( .A(n75411), .Z(n75412) );
  NOR U95691 ( .A(n75413), .B(n75412), .Z(n80816) );
  IV U95692 ( .A(n75414), .Z(n75415) );
  NOR U95693 ( .A(n75415), .B(n75417), .Z(n86206) );
  IV U95694 ( .A(n75416), .Z(n75418) );
  NOR U95695 ( .A(n75418), .B(n75417), .Z(n80841) );
  NOR U95696 ( .A(n75419), .B(n80841), .Z(n80448) );
  IV U95697 ( .A(n75420), .Z(n75422) );
  NOR U95698 ( .A(n75422), .B(n75421), .Z(n80851) );
  IV U95699 ( .A(n75423), .Z(n75424) );
  NOR U95700 ( .A(n75425), .B(n75424), .Z(n80849) );
  NOR U95701 ( .A(n80851), .B(n80849), .Z(n80447) );
  IV U95702 ( .A(n75426), .Z(n75429) );
  NOR U95703 ( .A(n80445), .B(n75427), .Z(n75428) );
  IV U95704 ( .A(n75428), .Z(n75435) );
  NOR U95705 ( .A(n75429), .B(n75435), .Z(n86189) );
  IV U95706 ( .A(n75430), .Z(n75433) );
  IV U95707 ( .A(n75431), .Z(n75432) );
  NOR U95708 ( .A(n75433), .B(n75432), .Z(n80855) );
  IV U95709 ( .A(n75434), .Z(n75436) );
  NOR U95710 ( .A(n75436), .B(n75435), .Z(n80856) );
  XOR U95711 ( .A(n80855), .B(n80856), .Z(n75437) );
  NOR U95712 ( .A(n86189), .B(n75437), .Z(n80442) );
  IV U95713 ( .A(n75438), .Z(n75439) );
  NOR U95714 ( .A(n75441), .B(n75439), .Z(n86172) );
  NOR U95715 ( .A(n75441), .B(n75440), .Z(n86169) );
  NOR U95716 ( .A(n75447), .B(n75442), .Z(n80861) );
  IV U95717 ( .A(n75443), .Z(n75444) );
  NOR U95718 ( .A(n75447), .B(n75444), .Z(n80867) );
  IV U95719 ( .A(n75445), .Z(n75446) );
  NOR U95720 ( .A(n75447), .B(n75446), .Z(n80864) );
  IV U95721 ( .A(n75450), .Z(n75448) );
  NOR U95722 ( .A(n75448), .B(n75454), .Z(n80873) );
  IV U95723 ( .A(n75449), .Z(n75452) );
  XOR U95724 ( .A(n75450), .B(n75454), .Z(n75451) );
  NOR U95725 ( .A(n75452), .B(n75451), .Z(n86162) );
  NOR U95726 ( .A(n80873), .B(n86162), .Z(n80437) );
  IV U95727 ( .A(n75453), .Z(n75455) );
  NOR U95728 ( .A(n75455), .B(n75454), .Z(n86161) );
  IV U95729 ( .A(n75456), .Z(n80889) );
  IV U95730 ( .A(n75457), .Z(n75458) );
  NOR U95731 ( .A(n75458), .B(n86138), .Z(n75460) );
  NOR U95732 ( .A(n75460), .B(n75459), .Z(n80896) );
  NOR U95733 ( .A(n75461), .B(n86138), .Z(n75462) );
  IV U95734 ( .A(n75462), .Z(n86150) );
  NOR U95735 ( .A(n75464), .B(n75463), .Z(n80897) );
  IV U95736 ( .A(n75465), .Z(n86142) );
  NOR U95737 ( .A(n75466), .B(n86142), .Z(n75467) );
  NOR U95738 ( .A(n80897), .B(n75467), .Z(n80422) );
  IV U95739 ( .A(n75468), .Z(n75469) );
  NOR U95740 ( .A(n75469), .B(n86115), .Z(n80413) );
  IV U95741 ( .A(n75470), .Z(n75472) );
  IV U95742 ( .A(n75471), .Z(n75477) );
  NOR U95743 ( .A(n75472), .B(n75477), .Z(n80905) );
  IV U95744 ( .A(n75473), .Z(n75475) );
  NOR U95745 ( .A(n75475), .B(n75474), .Z(n80903) );
  NOR U95746 ( .A(n80905), .B(n80903), .Z(n80402) );
  IV U95747 ( .A(n75476), .Z(n75478) );
  NOR U95748 ( .A(n75478), .B(n75477), .Z(n86102) );
  NOR U95749 ( .A(n80909), .B(n86102), .Z(n80401) );
  NOR U95750 ( .A(n80918), .B(n80911), .Z(n80400) );
  NOR U95751 ( .A(n75480), .B(n75479), .Z(n80917) );
  IV U95752 ( .A(n80917), .Z(n80915) );
  IV U95753 ( .A(n75481), .Z(n75483) );
  IV U95754 ( .A(n75482), .Z(n80398) );
  NOR U95755 ( .A(n75483), .B(n80398), .Z(n75484) );
  IV U95756 ( .A(n75484), .Z(n86100) );
  IV U95757 ( .A(n75485), .Z(n75487) );
  NOR U95758 ( .A(n75487), .B(n75486), .Z(n80924) );
  IV U95759 ( .A(n75488), .Z(n75491) );
  IV U95760 ( .A(n75489), .Z(n75490) );
  NOR U95761 ( .A(n75491), .B(n75490), .Z(n86093) );
  NOR U95762 ( .A(n80924), .B(n86093), .Z(n80396) );
  IV U95763 ( .A(n75492), .Z(n75498) );
  NOR U95764 ( .A(n75493), .B(n75500), .Z(n75494) );
  IV U95765 ( .A(n75494), .Z(n75495) );
  NOR U95766 ( .A(n75496), .B(n75495), .Z(n75497) );
  IV U95767 ( .A(n75497), .Z(n80386) );
  NOR U95768 ( .A(n75498), .B(n80386), .Z(n80930) );
  IV U95769 ( .A(n75499), .Z(n75501) );
  NOR U95770 ( .A(n75501), .B(n75500), .Z(n86060) );
  IV U95771 ( .A(n75502), .Z(n75503) );
  NOR U95772 ( .A(n75507), .B(n75503), .Z(n75504) );
  IV U95773 ( .A(n75504), .Z(n80948) );
  IV U95774 ( .A(n75505), .Z(n75506) );
  NOR U95775 ( .A(n75507), .B(n75506), .Z(n80369) );
  IV U95776 ( .A(n80369), .Z(n80361) );
  IV U95777 ( .A(n75508), .Z(n75509) );
  NOR U95778 ( .A(n75510), .B(n75509), .Z(n75511) );
  IV U95779 ( .A(n75511), .Z(n80952) );
  IV U95780 ( .A(n75512), .Z(n75514) );
  IV U95781 ( .A(n75515), .Z(n75523) );
  NOR U95782 ( .A(n75514), .B(n75523), .Z(n75521) );
  IV U95783 ( .A(n75513), .Z(n75519) );
  XOR U95784 ( .A(n75522), .B(n75515), .Z(n75517) );
  NOR U95785 ( .A(n75515), .B(n75514), .Z(n75516) );
  NOR U95786 ( .A(n75517), .B(n75516), .Z(n75518) );
  NOR U95787 ( .A(n75519), .B(n75518), .Z(n75520) );
  NOR U95788 ( .A(n75521), .B(n75520), .Z(n80950) );
  IV U95789 ( .A(n75522), .Z(n75524) );
  NOR U95790 ( .A(n75524), .B(n75523), .Z(n86052) );
  IV U95791 ( .A(n75525), .Z(n75526) );
  NOR U95792 ( .A(n75529), .B(n75526), .Z(n80956) );
  NOR U95793 ( .A(n86052), .B(n80956), .Z(n80359) );
  IV U95794 ( .A(n75527), .Z(n75531) );
  NOR U95795 ( .A(n75529), .B(n75528), .Z(n75530) );
  IV U95796 ( .A(n75530), .Z(n75533) );
  NOR U95797 ( .A(n75531), .B(n75533), .Z(n86047) );
  IV U95798 ( .A(n75532), .Z(n75534) );
  NOR U95799 ( .A(n75534), .B(n75533), .Z(n86044) );
  IV U95800 ( .A(n75535), .Z(n75536) );
  NOR U95801 ( .A(n75538), .B(n75536), .Z(n86040) );
  IV U95802 ( .A(n75537), .Z(n75539) );
  NOR U95803 ( .A(n75539), .B(n75538), .Z(n86039) );
  XOR U95804 ( .A(n86040), .B(n86039), .Z(n75540) );
  NOR U95805 ( .A(n86044), .B(n75540), .Z(n80358) );
  IV U95806 ( .A(n75541), .Z(n75542) );
  NOR U95807 ( .A(n75543), .B(n75542), .Z(n80958) );
  IV U95808 ( .A(n75544), .Z(n75545) );
  NOR U95809 ( .A(n75546), .B(n75545), .Z(n86034) );
  NOR U95810 ( .A(n80958), .B(n86034), .Z(n80357) );
  IV U95811 ( .A(n75547), .Z(n75549) );
  IV U95812 ( .A(n75548), .Z(n75551) );
  NOR U95813 ( .A(n75549), .B(n75551), .Z(n80960) );
  IV U95814 ( .A(n75550), .Z(n75552) );
  NOR U95815 ( .A(n75552), .B(n75551), .Z(n86018) );
  IV U95816 ( .A(n75553), .Z(n75554) );
  NOR U95817 ( .A(n75557), .B(n75554), .Z(n86015) );
  IV U95818 ( .A(n75555), .Z(n75559) );
  NOR U95819 ( .A(n75557), .B(n75556), .Z(n75558) );
  IV U95820 ( .A(n75558), .Z(n75561) );
  NOR U95821 ( .A(n75559), .B(n75561), .Z(n80963) );
  IV U95822 ( .A(n75560), .Z(n75562) );
  NOR U95823 ( .A(n75562), .B(n75561), .Z(n86010) );
  IV U95824 ( .A(n75563), .Z(n75567) );
  IV U95825 ( .A(n75564), .Z(n75570) );
  NOR U95826 ( .A(n75570), .B(n75565), .Z(n75566) );
  IV U95827 ( .A(n75566), .Z(n75572) );
  NOR U95828 ( .A(n75567), .B(n75572), .Z(n80974) );
  IV U95829 ( .A(n75568), .Z(n75569) );
  NOR U95830 ( .A(n75570), .B(n75569), .Z(n85999) );
  IV U95831 ( .A(n75571), .Z(n75573) );
  NOR U95832 ( .A(n75573), .B(n75572), .Z(n80977) );
  NOR U95833 ( .A(n85999), .B(n80977), .Z(n75574) );
  IV U95834 ( .A(n75574), .Z(n80341) );
  IV U95835 ( .A(n75575), .Z(n75576) );
  NOR U95836 ( .A(n75576), .B(n75578), .Z(n80980) );
  IV U95837 ( .A(n75577), .Z(n75579) );
  NOR U95838 ( .A(n75579), .B(n75578), .Z(n75580) );
  IV U95839 ( .A(n75580), .Z(n80984) );
  IV U95840 ( .A(n75581), .Z(n75583) );
  NOR U95841 ( .A(n75583), .B(n75582), .Z(n80337) );
  IV U95842 ( .A(n75584), .Z(n75587) );
  NOR U95843 ( .A(n75585), .B(n75590), .Z(n75586) );
  IV U95844 ( .A(n75586), .Z(n80306) );
  NOR U95845 ( .A(n75587), .B(n80306), .Z(n75588) );
  IV U95846 ( .A(n75588), .Z(n81016) );
  IV U95847 ( .A(n75589), .Z(n75591) );
  NOR U95848 ( .A(n75591), .B(n75590), .Z(n80303) );
  IV U95849 ( .A(n80303), .Z(n80295) );
  IV U95850 ( .A(n75592), .Z(n75593) );
  NOR U95851 ( .A(n75593), .B(n75596), .Z(n75594) );
  IV U95852 ( .A(n75594), .Z(n81023) );
  IV U95853 ( .A(n75595), .Z(n75597) );
  NOR U95854 ( .A(n75597), .B(n75596), .Z(n81028) );
  IV U95855 ( .A(n75598), .Z(n75607) );
  IV U95856 ( .A(n75599), .Z(n75600) );
  NOR U95857 ( .A(n75607), .B(n75600), .Z(n75601) );
  IV U95858 ( .A(n75601), .Z(n81026) );
  IV U95859 ( .A(n75602), .Z(n75604) );
  NOR U95860 ( .A(n75604), .B(n75603), .Z(n81033) );
  IV U95861 ( .A(n75605), .Z(n75606) );
  NOR U95862 ( .A(n75607), .B(n75606), .Z(n81031) );
  NOR U95863 ( .A(n81033), .B(n81031), .Z(n80293) );
  IV U95864 ( .A(n75608), .Z(n75610) );
  NOR U95865 ( .A(n75610), .B(n75609), .Z(n81041) );
  IV U95866 ( .A(n75611), .Z(n75612) );
  NOR U95867 ( .A(n75612), .B(n80288), .Z(n81038) );
  NOR U95868 ( .A(n81041), .B(n81038), .Z(n80292) );
  IV U95869 ( .A(n75613), .Z(n75618) );
  IV U95870 ( .A(n75614), .Z(n75615) );
  NOR U95871 ( .A(n75626), .B(n75615), .Z(n75616) );
  IV U95872 ( .A(n75616), .Z(n75617) );
  NOR U95873 ( .A(n75618), .B(n75617), .Z(n75619) );
  IV U95874 ( .A(n75619), .Z(n85978) );
  IV U95875 ( .A(n75620), .Z(n75623) );
  NOR U95876 ( .A(n75621), .B(n75634), .Z(n75622) );
  IV U95877 ( .A(n75622), .Z(n75631) );
  NOR U95878 ( .A(n75623), .B(n75631), .Z(n81055) );
  IV U95879 ( .A(n75624), .Z(n75629) );
  NOR U95880 ( .A(n75626), .B(n75625), .Z(n75627) );
  IV U95881 ( .A(n75627), .Z(n75628) );
  NOR U95882 ( .A(n75629), .B(n75628), .Z(n81048) );
  NOR U95883 ( .A(n81055), .B(n81048), .Z(n80273) );
  IV U95884 ( .A(n75630), .Z(n75632) );
  NOR U95885 ( .A(n75632), .B(n75631), .Z(n81054) );
  IV U95886 ( .A(n81054), .Z(n81052) );
  IV U95887 ( .A(n75633), .Z(n75635) );
  NOR U95888 ( .A(n75635), .B(n75634), .Z(n80269) );
  IV U95889 ( .A(n75636), .Z(n75639) );
  IV U95890 ( .A(n75637), .Z(n75638) );
  NOR U95891 ( .A(n75639), .B(n75638), .Z(n75640) );
  IV U95892 ( .A(n75640), .Z(n85952) );
  IV U95893 ( .A(n75641), .Z(n75642) );
  NOR U95894 ( .A(n75645), .B(n75642), .Z(n81066) );
  IV U95895 ( .A(n75643), .Z(n75644) );
  NOR U95896 ( .A(n75645), .B(n75644), .Z(n81072) );
  IV U95897 ( .A(n75646), .Z(n75647) );
  NOR U95898 ( .A(n75647), .B(n75654), .Z(n75648) );
  IV U95899 ( .A(n75648), .Z(n81078) );
  IV U95900 ( .A(n75649), .Z(n75650) );
  NOR U95901 ( .A(n75651), .B(n75650), .Z(n81080) );
  IV U95902 ( .A(n75652), .Z(n75653) );
  NOR U95903 ( .A(n75654), .B(n75653), .Z(n81086) );
  NOR U95904 ( .A(n81080), .B(n81086), .Z(n80253) );
  IV U95905 ( .A(n75655), .Z(n75657) );
  IV U95906 ( .A(n75656), .Z(n75660) );
  NOR U95907 ( .A(n75657), .B(n75660), .Z(n81083) );
  NOR U95908 ( .A(n75658), .B(n81093), .Z(n75662) );
  IV U95909 ( .A(n75659), .Z(n75661) );
  NOR U95910 ( .A(n75661), .B(n75660), .Z(n81090) );
  NOR U95911 ( .A(n75662), .B(n81090), .Z(n80252) );
  IV U95912 ( .A(n75663), .Z(n75665) );
  NOR U95913 ( .A(n75665), .B(n75664), .Z(n85931) );
  IV U95914 ( .A(n75666), .Z(n75667) );
  NOR U95915 ( .A(n75668), .B(n75667), .Z(n85934) );
  NOR U95916 ( .A(n85931), .B(n85934), .Z(n80251) );
  IV U95917 ( .A(n75669), .Z(n75672) );
  NOR U95918 ( .A(n75670), .B(n75674), .Z(n75671) );
  IV U95919 ( .A(n75671), .Z(n80248) );
  NOR U95920 ( .A(n75672), .B(n80248), .Z(n81098) );
  IV U95921 ( .A(n75673), .Z(n75675) );
  NOR U95922 ( .A(n75675), .B(n75674), .Z(n81107) );
  IV U95923 ( .A(n75676), .Z(n75678) );
  NOR U95924 ( .A(n75678), .B(n75677), .Z(n81102) );
  NOR U95925 ( .A(n81107), .B(n81102), .Z(n80242) );
  IV U95926 ( .A(n75679), .Z(n75680) );
  NOR U95927 ( .A(n75680), .B(n80223), .Z(n81117) );
  IV U95928 ( .A(n75681), .Z(n75683) );
  NOR U95929 ( .A(n75683), .B(n75682), .Z(n80212) );
  IV U95930 ( .A(n80212), .Z(n80210) );
  IV U95931 ( .A(n75684), .Z(n75688) );
  NOR U95932 ( .A(n75686), .B(n75685), .Z(n75687) );
  IV U95933 ( .A(n75687), .Z(n75691) );
  NOR U95934 ( .A(n75688), .B(n75691), .Z(n75689) );
  IV U95935 ( .A(n75689), .Z(n81138) );
  IV U95936 ( .A(n75690), .Z(n75692) );
  NOR U95937 ( .A(n75692), .B(n75691), .Z(n75693) );
  NOR U95938 ( .A(n75694), .B(n75693), .Z(n81136) );
  NOR U95939 ( .A(n75696), .B(n75695), .Z(n81147) );
  NOR U95940 ( .A(n81147), .B(n81139), .Z(n80208) );
  IV U95941 ( .A(n75697), .Z(n75699) );
  NOR U95942 ( .A(n75699), .B(n75698), .Z(n81142) );
  IV U95943 ( .A(n81142), .Z(n81144) );
  IV U95944 ( .A(n75700), .Z(n75703) );
  NOR U95945 ( .A(n75701), .B(n80205), .Z(n75702) );
  IV U95946 ( .A(n75702), .Z(n80202) );
  NOR U95947 ( .A(n75703), .B(n80202), .Z(n80195) );
  NOR U95948 ( .A(n75705), .B(n75704), .Z(n80192) );
  IV U95949 ( .A(n80192), .Z(n80183) );
  IV U95950 ( .A(n75706), .Z(n75707) );
  NOR U95951 ( .A(n75708), .B(n75707), .Z(n85892) );
  IV U95952 ( .A(n75709), .Z(n75710) );
  NOR U95953 ( .A(n75711), .B(n75710), .Z(n85893) );
  NOR U95954 ( .A(n85892), .B(n85893), .Z(n80181) );
  IV U95955 ( .A(n75712), .Z(n75715) );
  IV U95956 ( .A(n75713), .Z(n75714) );
  NOR U95957 ( .A(n75715), .B(n75714), .Z(n81152) );
  IV U95958 ( .A(n75716), .Z(n75717) );
  NOR U95959 ( .A(n75718), .B(n75717), .Z(n86925) );
  IV U95960 ( .A(n86925), .Z(n81159) );
  IV U95961 ( .A(n75719), .Z(n75721) );
  IV U95962 ( .A(n75720), .Z(n75725) );
  NOR U95963 ( .A(n75721), .B(n75725), .Z(n81155) );
  IV U95964 ( .A(n75722), .Z(n75723) );
  NOR U95965 ( .A(n75723), .B(n75728), .Z(n81165) );
  IV U95966 ( .A(n75724), .Z(n75726) );
  NOR U95967 ( .A(n75726), .B(n75725), .Z(n81156) );
  NOR U95968 ( .A(n81165), .B(n81156), .Z(n80170) );
  IV U95969 ( .A(n75727), .Z(n75729) );
  NOR U95970 ( .A(n75729), .B(n75728), .Z(n81163) );
  IV U95971 ( .A(n75735), .Z(n75733) );
  IV U95972 ( .A(n75730), .Z(n75731) );
  NOR U95973 ( .A(n75733), .B(n75731), .Z(n85861) );
  NOR U95974 ( .A(n75733), .B(n75732), .Z(n85864) );
  IV U95975 ( .A(n75734), .Z(n75738) );
  NOR U95976 ( .A(n75741), .B(n75735), .Z(n75736) );
  IV U95977 ( .A(n75736), .Z(n75737) );
  NOR U95978 ( .A(n75738), .B(n75737), .Z(n85850) );
  NOR U95979 ( .A(n85864), .B(n85850), .Z(n80160) );
  IV U95980 ( .A(n75739), .Z(n75744) );
  NOR U95981 ( .A(n75741), .B(n75740), .Z(n75742) );
  IV U95982 ( .A(n75742), .Z(n75743) );
  NOR U95983 ( .A(n75744), .B(n75743), .Z(n81177) );
  IV U95984 ( .A(n75745), .Z(n85845) );
  XOR U95985 ( .A(n75746), .B(n85845), .Z(n75747) );
  NOR U95986 ( .A(n75755), .B(n75747), .Z(n75753) );
  IV U95987 ( .A(n75748), .Z(n75750) );
  NOR U95988 ( .A(n75750), .B(n75749), .Z(n75751) );
  IV U95989 ( .A(n75751), .Z(n85835) );
  NOR U95990 ( .A(n85845), .B(n75755), .Z(n81181) );
  NOR U95991 ( .A(n85835), .B(n81181), .Z(n75752) );
  NOR U95992 ( .A(n75753), .B(n75752), .Z(n80154) );
  IV U95993 ( .A(n75754), .Z(n75756) );
  NOR U95994 ( .A(n75756), .B(n75755), .Z(n81180) );
  IV U95995 ( .A(n75757), .Z(n75758) );
  NOR U95996 ( .A(n80147), .B(n75758), .Z(n85832) );
  IV U95997 ( .A(n75759), .Z(n75760) );
  NOR U95998 ( .A(n75760), .B(n80131), .Z(n81192) );
  IV U95999 ( .A(n75761), .Z(n75763) );
  IV U96000 ( .A(n75762), .Z(n75770) );
  NOR U96001 ( .A(n75763), .B(n75770), .Z(n75768) );
  IV U96002 ( .A(n75764), .Z(n75766) );
  NOR U96003 ( .A(n75766), .B(n75765), .Z(n75767) );
  NOR U96004 ( .A(n75768), .B(n75767), .Z(n81191) );
  IV U96005 ( .A(n75769), .Z(n75771) );
  NOR U96006 ( .A(n75771), .B(n75770), .Z(n81198) );
  IV U96007 ( .A(n75772), .Z(n75774) );
  NOR U96008 ( .A(n75774), .B(n75773), .Z(n75775) );
  IV U96009 ( .A(n75775), .Z(n80120) );
  IV U96010 ( .A(n75776), .Z(n75777) );
  NOR U96011 ( .A(n80112), .B(n75777), .Z(n81209) );
  IV U96012 ( .A(n75778), .Z(n75779) );
  NOR U96013 ( .A(n75779), .B(n80112), .Z(n81206) );
  IV U96014 ( .A(n75780), .Z(n75781) );
  NOR U96015 ( .A(n75782), .B(n75781), .Z(n75783) );
  IV U96016 ( .A(n75783), .Z(n81231) );
  IV U96017 ( .A(n75784), .Z(n75785) );
  NOR U96018 ( .A(n81242), .B(n75785), .Z(n81251) );
  NOR U96019 ( .A(n75786), .B(n81235), .Z(n75787) );
  NOR U96020 ( .A(n81251), .B(n75787), .Z(n80090) );
  IV U96021 ( .A(n75788), .Z(n75789) );
  NOR U96022 ( .A(n75789), .B(n80087), .Z(n81246) );
  IV U96023 ( .A(n81246), .Z(n81249) );
  IV U96024 ( .A(n80077), .Z(n80068) );
  IV U96025 ( .A(n75790), .Z(n75794) );
  IV U96026 ( .A(n75791), .Z(n75796) );
  NOR U96027 ( .A(n75792), .B(n75796), .Z(n75793) );
  IV U96028 ( .A(n75793), .Z(n80061) );
  NOR U96029 ( .A(n75794), .B(n80061), .Z(n80051) );
  IV U96030 ( .A(n75795), .Z(n75797) );
  NOR U96031 ( .A(n75797), .B(n75796), .Z(n80049) );
  IV U96032 ( .A(n80049), .Z(n80043) );
  IV U96033 ( .A(n75798), .Z(n75800) );
  IV U96034 ( .A(n75799), .Z(n75802) );
  NOR U96035 ( .A(n75800), .B(n75802), .Z(n85758) );
  IV U96036 ( .A(n75801), .Z(n75803) );
  NOR U96037 ( .A(n75803), .B(n75802), .Z(n81266) );
  IV U96038 ( .A(n75804), .Z(n75805) );
  NOR U96039 ( .A(n80040), .B(n75805), .Z(n80034) );
  IV U96040 ( .A(n75806), .Z(n75807) );
  NOR U96041 ( .A(n75807), .B(n75813), .Z(n85737) );
  NOR U96042 ( .A(n75809), .B(n75808), .Z(n81277) );
  NOR U96043 ( .A(n85737), .B(n81277), .Z(n80027) );
  IV U96044 ( .A(n75810), .Z(n81283) );
  NOR U96045 ( .A(n81283), .B(n75811), .Z(n75815) );
  IV U96046 ( .A(n75812), .Z(n75814) );
  NOR U96047 ( .A(n75814), .B(n75813), .Z(n85740) );
  NOR U96048 ( .A(n75815), .B(n85740), .Z(n80026) );
  IV U96049 ( .A(n75816), .Z(n75817) );
  NOR U96050 ( .A(n75817), .B(n80012), .Z(n75818) );
  IV U96051 ( .A(n75818), .Z(n81280) );
  NOR U96052 ( .A(n80005), .B(n75819), .Z(n75820) );
  IV U96053 ( .A(n75820), .Z(n75825) );
  NOR U96054 ( .A(n75822), .B(n75821), .Z(n75823) );
  IV U96055 ( .A(n75823), .Z(n75824) );
  NOR U96056 ( .A(n75825), .B(n75824), .Z(n75826) );
  IV U96057 ( .A(n75826), .Z(n75827) );
  NOR U96058 ( .A(n75828), .B(n75827), .Z(n85721) );
  IV U96059 ( .A(n75829), .Z(n75830) );
  NOR U96060 ( .A(n80005), .B(n75830), .Z(n85714) );
  IV U96061 ( .A(n75831), .Z(n80007) );
  IV U96062 ( .A(n75832), .Z(n75833) );
  NOR U96063 ( .A(n80007), .B(n75833), .Z(n85704) );
  NOR U96064 ( .A(n75835), .B(n75834), .Z(n81291) );
  IV U96065 ( .A(n75836), .Z(n75837) );
  NOR U96066 ( .A(n75837), .B(n80001), .Z(n75838) );
  IV U96067 ( .A(n75838), .Z(n81298) );
  NOR U96068 ( .A(n80001), .B(n75839), .Z(n81300) );
  IV U96069 ( .A(n75840), .Z(n75841) );
  NOR U96070 ( .A(n75844), .B(n75841), .Z(n81307) );
  NOR U96071 ( .A(n81300), .B(n81307), .Z(n79999) );
  IV U96072 ( .A(n75842), .Z(n75843) );
  NOR U96073 ( .A(n75844), .B(n75843), .Z(n81304) );
  IV U96074 ( .A(n75845), .Z(n75849) );
  NOR U96075 ( .A(n75847), .B(n75846), .Z(n75848) );
  IV U96076 ( .A(n75848), .Z(n75851) );
  NOR U96077 ( .A(n75849), .B(n75851), .Z(n85694) );
  IV U96078 ( .A(n75850), .Z(n75852) );
  NOR U96079 ( .A(n75852), .B(n75851), .Z(n81313) );
  IV U96080 ( .A(n75853), .Z(n75855) );
  IV U96081 ( .A(n75854), .Z(n79988) );
  NOR U96082 ( .A(n75855), .B(n79988), .Z(n81310) );
  IV U96083 ( .A(n75856), .Z(n75858) );
  XOR U96084 ( .A(n79992), .B(n79994), .Z(n75857) );
  NOR U96085 ( .A(n75858), .B(n75857), .Z(n85686) );
  IV U96086 ( .A(n75859), .Z(n75860) );
  NOR U96087 ( .A(n75860), .B(n75865), .Z(n85679) );
  IV U96088 ( .A(n75861), .Z(n75869) );
  IV U96089 ( .A(n75862), .Z(n75863) );
  NOR U96090 ( .A(n75869), .B(n75863), .Z(n85674) );
  IV U96091 ( .A(n75864), .Z(n75866) );
  NOR U96092 ( .A(n75866), .B(n75865), .Z(n81320) );
  NOR U96093 ( .A(n85674), .B(n81320), .Z(n79986) );
  IV U96094 ( .A(n75867), .Z(n75868) );
  NOR U96095 ( .A(n75869), .B(n75868), .Z(n81325) );
  IV U96096 ( .A(n75870), .Z(n75871) );
  NOR U96097 ( .A(n75872), .B(n75871), .Z(n81322) );
  NOR U96098 ( .A(n75874), .B(n75873), .Z(n75880) );
  NOR U96099 ( .A(n75876), .B(n75875), .Z(n75877) );
  NOR U96100 ( .A(n75878), .B(n75877), .Z(n75879) );
  NOR U96101 ( .A(n75880), .B(n75879), .Z(n81333) );
  IV U96102 ( .A(n75881), .Z(n75888) );
  NOR U96103 ( .A(n75883), .B(n75882), .Z(n75884) );
  IV U96104 ( .A(n75884), .Z(n75885) );
  NOR U96105 ( .A(n75886), .B(n75885), .Z(n75887) );
  IV U96106 ( .A(n75887), .Z(n75890) );
  NOR U96107 ( .A(n75888), .B(n75890), .Z(n81330) );
  IV U96108 ( .A(n75889), .Z(n75891) );
  NOR U96109 ( .A(n75891), .B(n75890), .Z(n81339) );
  NOR U96110 ( .A(n75892), .B(n79953), .Z(n75893) );
  IV U96111 ( .A(n75893), .Z(n75900) );
  XOR U96112 ( .A(n75895), .B(n75894), .Z(n75897) );
  NOR U96113 ( .A(n75897), .B(n75896), .Z(n75898) );
  IV U96114 ( .A(n75898), .Z(n75899) );
  NOR U96115 ( .A(n75900), .B(n75899), .Z(n75901) );
  IV U96116 ( .A(n75901), .Z(n75902) );
  NOR U96117 ( .A(n79950), .B(n75902), .Z(n75903) );
  IV U96118 ( .A(n75903), .Z(n75904) );
  NOR U96119 ( .A(n75905), .B(n75904), .Z(n81365) );
  IV U96120 ( .A(n75906), .Z(n79918) );
  IV U96121 ( .A(n75907), .Z(n75908) );
  NOR U96122 ( .A(n79918), .B(n75908), .Z(n85661) );
  IV U96123 ( .A(n75909), .Z(n75912) );
  NOR U96124 ( .A(n75910), .B(n79920), .Z(n75911) );
  IV U96125 ( .A(n75911), .Z(n75917) );
  NOR U96126 ( .A(n75912), .B(n75917), .Z(n81380) );
  IV U96127 ( .A(n75913), .Z(n75915) );
  NOR U96128 ( .A(n75915), .B(n75914), .Z(n85656) );
  IV U96129 ( .A(n75916), .Z(n75918) );
  NOR U96130 ( .A(n75918), .B(n75917), .Z(n81389) );
  NOR U96131 ( .A(n85656), .B(n81389), .Z(n79915) );
  IV U96132 ( .A(n75919), .Z(n75920) );
  NOR U96133 ( .A(n75920), .B(n79902), .Z(n75921) );
  IV U96134 ( .A(n75921), .Z(n85652) );
  IV U96135 ( .A(n75922), .Z(n75923) );
  NOR U96136 ( .A(n75924), .B(n75923), .Z(n81400) );
  IV U96137 ( .A(n75925), .Z(n75926) );
  NOR U96138 ( .A(n79892), .B(n75926), .Z(n81398) );
  NOR U96139 ( .A(n81400), .B(n81398), .Z(n79897) );
  IV U96140 ( .A(n75927), .Z(n75928) );
  NOR U96141 ( .A(n75928), .B(n79875), .Z(n75929) );
  IV U96142 ( .A(n75929), .Z(n81405) );
  IV U96143 ( .A(n75930), .Z(n75931) );
  NOR U96144 ( .A(n75932), .B(n75931), .Z(n81407) );
  IV U96145 ( .A(n75933), .Z(n79871) );
  IV U96146 ( .A(n75934), .Z(n75935) );
  NOR U96147 ( .A(n79871), .B(n75935), .Z(n81411) );
  NOR U96148 ( .A(n81407), .B(n81411), .Z(n79873) );
  IV U96149 ( .A(n75936), .Z(n75938) );
  NOR U96150 ( .A(n75938), .B(n75937), .Z(n81413) );
  IV U96151 ( .A(n75939), .Z(n75940) );
  NOR U96152 ( .A(n75940), .B(n75942), .Z(n81424) );
  IV U96153 ( .A(n75941), .Z(n75943) );
  NOR U96154 ( .A(n75943), .B(n75942), .Z(n75944) );
  IV U96155 ( .A(n75944), .Z(n81422) );
  IV U96156 ( .A(n75945), .Z(n75946) );
  NOR U96157 ( .A(n75946), .B(n75949), .Z(n75947) );
  IV U96158 ( .A(n75947), .Z(n81435) );
  IV U96159 ( .A(n75948), .Z(n75950) );
  NOR U96160 ( .A(n75950), .B(n75949), .Z(n85642) );
  IV U96161 ( .A(n75951), .Z(n75953) );
  NOR U96162 ( .A(n75953), .B(n75952), .Z(n81437) );
  NOR U96163 ( .A(n85642), .B(n81437), .Z(n79861) );
  IV U96164 ( .A(n75954), .Z(n75956) );
  IV U96165 ( .A(n75955), .Z(n75960) );
  NOR U96166 ( .A(n75956), .B(n75960), .Z(n85636) );
  IV U96167 ( .A(n75957), .Z(n75958) );
  NOR U96168 ( .A(n75958), .B(n75966), .Z(n81442) );
  IV U96169 ( .A(n75959), .Z(n75961) );
  NOR U96170 ( .A(n75961), .B(n75960), .Z(n81440) );
  NOR U96171 ( .A(n81442), .B(n81440), .Z(n79860) );
  IV U96172 ( .A(n75962), .Z(n75963) );
  NOR U96173 ( .A(n75964), .B(n75963), .Z(n85628) );
  IV U96174 ( .A(n75965), .Z(n75967) );
  NOR U96175 ( .A(n75967), .B(n75966), .Z(n85632) );
  NOR U96176 ( .A(n85628), .B(n85632), .Z(n79859) );
  IV U96177 ( .A(n75968), .Z(n75969) );
  NOR U96178 ( .A(n75970), .B(n75969), .Z(n85626) );
  IV U96179 ( .A(n75971), .Z(n75972) );
  NOR U96180 ( .A(n75972), .B(n79854), .Z(n81446) );
  IV U96181 ( .A(n75973), .Z(n75974) );
  NOR U96182 ( .A(n75975), .B(n75974), .Z(n75980) );
  IV U96183 ( .A(n75976), .Z(n75978) );
  NOR U96184 ( .A(n75978), .B(n75977), .Z(n75979) );
  NOR U96185 ( .A(n75980), .B(n75979), .Z(n81454) );
  IV U96186 ( .A(n75981), .Z(n75986) );
  IV U96187 ( .A(n75982), .Z(n75983) );
  NOR U96188 ( .A(n75986), .B(n75983), .Z(n85607) );
  IV U96189 ( .A(n75984), .Z(n75985) );
  NOR U96190 ( .A(n75986), .B(n75985), .Z(n81462) );
  IV U96191 ( .A(n75987), .Z(n75988) );
  NOR U96192 ( .A(n75988), .B(n75990), .Z(n81459) );
  IV U96193 ( .A(n75989), .Z(n75991) );
  NOR U96194 ( .A(n75991), .B(n75990), .Z(n81467) );
  IV U96195 ( .A(n75992), .Z(n75993) );
  NOR U96196 ( .A(n75994), .B(n75993), .Z(n85599) );
  IV U96197 ( .A(n75995), .Z(n75997) );
  IV U96198 ( .A(n75996), .Z(n79823) );
  NOR U96199 ( .A(n75997), .B(n79823), .Z(n81470) );
  NOR U96200 ( .A(n85599), .B(n81470), .Z(n79833) );
  IV U96201 ( .A(n75998), .Z(n76004) );
  NOR U96202 ( .A(n76007), .B(n75999), .Z(n76000) );
  IV U96203 ( .A(n76000), .Z(n79829) );
  NOR U96204 ( .A(n76001), .B(n79829), .Z(n76002) );
  IV U96205 ( .A(n76002), .Z(n76003) );
  NOR U96206 ( .A(n76004), .B(n76003), .Z(n81477) );
  IV U96207 ( .A(n76005), .Z(n76006) );
  NOR U96208 ( .A(n76007), .B(n76006), .Z(n81474) );
  IV U96209 ( .A(n76008), .Z(n76010) );
  NOR U96210 ( .A(n76010), .B(n76009), .Z(n81485) );
  IV U96211 ( .A(n76011), .Z(n76013) );
  IV U96212 ( .A(n76012), .Z(n85587) );
  NOR U96213 ( .A(n76013), .B(n85587), .Z(n76018) );
  IV U96214 ( .A(n76014), .Z(n76016) );
  XOR U96215 ( .A(n76020), .B(n85587), .Z(n76015) );
  NOR U96216 ( .A(n76016), .B(n76015), .Z(n76017) );
  NOR U96217 ( .A(n76018), .B(n76017), .Z(n81483) );
  NOR U96218 ( .A(n76019), .B(n85579), .Z(n76023) );
  IV U96219 ( .A(n76020), .Z(n76021) );
  NOR U96220 ( .A(n76021), .B(n85587), .Z(n76022) );
  NOR U96221 ( .A(n76023), .B(n76022), .Z(n79821) );
  IV U96222 ( .A(n76024), .Z(n76029) );
  IV U96223 ( .A(n76025), .Z(n76026) );
  NOR U96224 ( .A(n76029), .B(n76026), .Z(n85575) );
  IV U96225 ( .A(n85575), .Z(n85573) );
  IV U96226 ( .A(n76027), .Z(n76028) );
  NOR U96227 ( .A(n76029), .B(n76028), .Z(n76030) );
  IV U96228 ( .A(n76030), .Z(n85570) );
  IV U96229 ( .A(n76031), .Z(n76032) );
  NOR U96230 ( .A(n76032), .B(n79809), .Z(n85566) );
  IV U96231 ( .A(n76033), .Z(n76034) );
  NOR U96232 ( .A(n76035), .B(n76034), .Z(n85558) );
  IV U96233 ( .A(n76036), .Z(n76037) );
  NOR U96234 ( .A(n76037), .B(n79816), .Z(n85561) );
  NOR U96235 ( .A(n85558), .B(n85561), .Z(n79806) );
  IV U96236 ( .A(n76038), .Z(n85548) );
  NOR U96237 ( .A(n85548), .B(n76039), .Z(n85553) );
  IV U96238 ( .A(n76040), .Z(n76041) );
  NOR U96239 ( .A(n76044), .B(n76041), .Z(n81498) );
  IV U96240 ( .A(n76042), .Z(n76043) );
  NOR U96241 ( .A(n76044), .B(n76043), .Z(n81496) );
  IV U96242 ( .A(n76045), .Z(n76046) );
  NOR U96243 ( .A(n76046), .B(n79787), .Z(n81510) );
  IV U96244 ( .A(n76047), .Z(n76051) );
  NOR U96245 ( .A(n76049), .B(n76048), .Z(n76050) );
  IV U96246 ( .A(n76050), .Z(n79754) );
  NOR U96247 ( .A(n76051), .B(n79754), .Z(n76052) );
  NOR U96248 ( .A(n76053), .B(n76052), .Z(n81533) );
  IV U96249 ( .A(n76054), .Z(n76058) );
  NOR U96250 ( .A(n76056), .B(n76055), .Z(n76057) );
  IV U96251 ( .A(n76057), .Z(n76063) );
  NOR U96252 ( .A(n76058), .B(n76063), .Z(n81529) );
  IV U96253 ( .A(n76059), .Z(n76060) );
  NOR U96254 ( .A(n76061), .B(n76060), .Z(n76065) );
  IV U96255 ( .A(n76062), .Z(n76064) );
  NOR U96256 ( .A(n76064), .B(n76063), .Z(n81534) );
  NOR U96257 ( .A(n76065), .B(n81534), .Z(n79751) );
  IV U96258 ( .A(n76066), .Z(n76067) );
  NOR U96259 ( .A(n76068), .B(n76067), .Z(n76069) );
  IV U96260 ( .A(n76069), .Z(n76071) );
  NOR U96261 ( .A(n76071), .B(n76070), .Z(n81553) );
  IV U96262 ( .A(n79738), .Z(n76072) );
  IV U96263 ( .A(n79740), .Z(n79737) );
  NOR U96264 ( .A(n76072), .B(n79737), .Z(n81560) );
  IV U96265 ( .A(n76073), .Z(n76074) );
  NOR U96266 ( .A(n76075), .B(n76074), .Z(n81569) );
  NOR U96267 ( .A(n76076), .B(n81566), .Z(n76077) );
  NOR U96268 ( .A(n81569), .B(n76077), .Z(n79734) );
  IV U96269 ( .A(n76078), .Z(n76080) );
  NOR U96270 ( .A(n76080), .B(n76079), .Z(n76081) );
  NOR U96271 ( .A(n76082), .B(n76081), .Z(n85527) );
  IV U96272 ( .A(n85529), .Z(n76089) );
  IV U96273 ( .A(n76086), .Z(n76087) );
  NOR U96274 ( .A(n76088), .B(n76087), .Z(n81573) );
  NOR U96275 ( .A(n76089), .B(n81573), .Z(n79733) );
  IV U96276 ( .A(n76090), .Z(n76092) );
  IV U96277 ( .A(n76091), .Z(n76094) );
  NOR U96278 ( .A(n76092), .B(n76094), .Z(n81572) );
  IV U96279 ( .A(n76093), .Z(n76095) );
  NOR U96280 ( .A(n76095), .B(n76094), .Z(n81580) );
  IV U96281 ( .A(n76096), .Z(n76097) );
  NOR U96282 ( .A(n76100), .B(n76097), .Z(n81577) );
  IV U96283 ( .A(n76098), .Z(n76099) );
  NOR U96284 ( .A(n76100), .B(n76099), .Z(n81583) );
  IV U96285 ( .A(n76101), .Z(n76106) );
  NOR U96286 ( .A(n76103), .B(n76102), .Z(n76104) );
  IV U96287 ( .A(n76104), .Z(n76105) );
  NOR U96288 ( .A(n76106), .B(n76105), .Z(n76107) );
  IV U96289 ( .A(n76107), .Z(n81588) );
  IV U96290 ( .A(n76108), .Z(n76110) );
  IV U96291 ( .A(n76109), .Z(n79722) );
  NOR U96292 ( .A(n76110), .B(n79722), .Z(n76111) );
  IV U96293 ( .A(n76111), .Z(n81586) );
  IV U96294 ( .A(n76112), .Z(n76114) );
  NOR U96295 ( .A(n76114), .B(n76113), .Z(n79719) );
  IV U96296 ( .A(n79719), .Z(n79714) );
  IV U96297 ( .A(n76115), .Z(n81605) );
  IV U96298 ( .A(n76116), .Z(n76118) );
  NOR U96299 ( .A(n76118), .B(n76117), .Z(n81602) );
  IV U96300 ( .A(n76119), .Z(n76121) );
  NOR U96301 ( .A(n76121), .B(n76120), .Z(n85501) );
  IV U96302 ( .A(n76122), .Z(n76123) );
  NOR U96303 ( .A(n76123), .B(n85504), .Z(n76124) );
  NOR U96304 ( .A(n85501), .B(n76124), .Z(n79701) );
  IV U96305 ( .A(n76125), .Z(n76127) );
  NOR U96306 ( .A(n76127), .B(n76126), .Z(n85496) );
  IV U96307 ( .A(n76128), .Z(n76129) );
  NOR U96308 ( .A(n76129), .B(n85504), .Z(n76130) );
  NOR U96309 ( .A(n85496), .B(n76130), .Z(n79700) );
  IV U96310 ( .A(n76131), .Z(n81610) );
  NOR U96311 ( .A(n81610), .B(n76132), .Z(n76136) );
  IV U96312 ( .A(n76133), .Z(n76135) );
  NOR U96313 ( .A(n76135), .B(n76134), .Z(n81606) );
  NOR U96314 ( .A(n76136), .B(n81606), .Z(n79699) );
  IV U96315 ( .A(n76137), .Z(n76138) );
  NOR U96316 ( .A(n76138), .B(n76140), .Z(n81613) );
  IV U96317 ( .A(n76139), .Z(n76141) );
  NOR U96318 ( .A(n76141), .B(n76140), .Z(n81622) );
  IV U96319 ( .A(n76142), .Z(n76146) );
  IV U96320 ( .A(n76143), .Z(n79693) );
  NOR U96321 ( .A(n79693), .B(n76144), .Z(n76145) );
  IV U96322 ( .A(n76145), .Z(n79697) );
  NOR U96323 ( .A(n76146), .B(n79697), .Z(n81619) );
  IV U96324 ( .A(n76147), .Z(n76150) );
  NOR U96325 ( .A(n76148), .B(n79689), .Z(n76149) );
  IV U96326 ( .A(n76149), .Z(n76152) );
  NOR U96327 ( .A(n76150), .B(n76152), .Z(n81626) );
  IV U96328 ( .A(n81626), .Z(n81628) );
  IV U96329 ( .A(n76151), .Z(n76153) );
  NOR U96330 ( .A(n76153), .B(n76152), .Z(n81637) );
  IV U96331 ( .A(n76154), .Z(n76156) );
  IV U96332 ( .A(n76155), .Z(n76158) );
  NOR U96333 ( .A(n76156), .B(n76158), .Z(n81634) );
  IV U96334 ( .A(n76157), .Z(n76159) );
  NOR U96335 ( .A(n76159), .B(n76158), .Z(n81640) );
  IV U96336 ( .A(n76160), .Z(n76161) );
  NOR U96337 ( .A(n85467), .B(n76161), .Z(n81643) );
  NOR U96338 ( .A(n81640), .B(n81643), .Z(n79687) );
  IV U96339 ( .A(n76162), .Z(n76163) );
  NOR U96340 ( .A(n76163), .B(n85467), .Z(n79686) );
  IV U96341 ( .A(n76164), .Z(n76169) );
  IV U96342 ( .A(n76165), .Z(n76166) );
  NOR U96343 ( .A(n76167), .B(n76166), .Z(n76168) );
  IV U96344 ( .A(n76168), .Z(n76171) );
  NOR U96345 ( .A(n76169), .B(n76171), .Z(n81647) );
  IV U96346 ( .A(n76170), .Z(n76172) );
  NOR U96347 ( .A(n76172), .B(n76171), .Z(n81653) );
  IV U96348 ( .A(n76173), .Z(n76174) );
  NOR U96349 ( .A(n79664), .B(n76174), .Z(n79669) );
  IV U96350 ( .A(n79669), .Z(n79667) );
  NOR U96351 ( .A(n76176), .B(n76175), .Z(n85443) );
  IV U96352 ( .A(n76177), .Z(n76178) );
  NOR U96353 ( .A(n76178), .B(n79648), .Z(n81673) );
  NOR U96354 ( .A(n81673), .B(n81668), .Z(n79660) );
  IV U96355 ( .A(n76179), .Z(n76180) );
  NOR U96356 ( .A(n76180), .B(n76182), .Z(n81683) );
  IV U96357 ( .A(n76181), .Z(n76183) );
  NOR U96358 ( .A(n76183), .B(n76182), .Z(n85426) );
  IV U96359 ( .A(n76184), .Z(n76186) );
  NOR U96360 ( .A(n76186), .B(n76185), .Z(n81686) );
  IV U96361 ( .A(n76187), .Z(n76189) );
  NOR U96362 ( .A(n76189), .B(n76188), .Z(n85429) );
  NOR U96363 ( .A(n81686), .B(n85429), .Z(n79642) );
  IV U96364 ( .A(n76190), .Z(n76191) );
  NOR U96365 ( .A(n76191), .B(n79639), .Z(n81689) );
  IV U96366 ( .A(n79633), .Z(n79631) );
  IV U96367 ( .A(n76192), .Z(n76193) );
  NOR U96368 ( .A(n76194), .B(n76193), .Z(n81699) );
  IV U96369 ( .A(n76195), .Z(n76198) );
  NOR U96370 ( .A(n76196), .B(n79622), .Z(n76197) );
  IV U96371 ( .A(n76197), .Z(n79628) );
  NOR U96372 ( .A(n76198), .B(n79628), .Z(n81704) );
  IV U96373 ( .A(n79601), .Z(n76199) );
  NOR U96374 ( .A(n76199), .B(n79604), .Z(n79598) );
  IV U96375 ( .A(n79598), .Z(n79591) );
  IV U96376 ( .A(n76200), .Z(n76201) );
  NOR U96377 ( .A(n76202), .B(n76201), .Z(n76207) );
  IV U96378 ( .A(n76203), .Z(n76205) );
  NOR U96379 ( .A(n76205), .B(n76204), .Z(n76206) );
  NOR U96380 ( .A(n76207), .B(n76206), .Z(n81721) );
  IV U96381 ( .A(n76208), .Z(n76209) );
  NOR U96382 ( .A(n76210), .B(n76209), .Z(n81726) );
  IV U96383 ( .A(n76211), .Z(n76212) );
  NOR U96384 ( .A(n76213), .B(n76212), .Z(n76214) );
  IV U96385 ( .A(n76214), .Z(n81746) );
  IV U96386 ( .A(n76215), .Z(n76217) );
  NOR U96387 ( .A(n76217), .B(n76216), .Z(n81750) );
  IV U96388 ( .A(n76218), .Z(n76219) );
  NOR U96389 ( .A(n76219), .B(n81738), .Z(n81748) );
  NOR U96390 ( .A(n81750), .B(n81748), .Z(n79588) );
  IV U96391 ( .A(n76220), .Z(n76222) );
  NOR U96392 ( .A(n76222), .B(n76221), .Z(n81758) );
  IV U96393 ( .A(n76223), .Z(n76224) );
  NOR U96394 ( .A(n76225), .B(n76224), .Z(n81753) );
  NOR U96395 ( .A(n81758), .B(n81753), .Z(n91165) );
  IV U96396 ( .A(n76226), .Z(n76227) );
  NOR U96397 ( .A(n76228), .B(n76227), .Z(n76229) );
  IV U96398 ( .A(n76229), .Z(n79584) );
  IV U96399 ( .A(n76230), .Z(n76231) );
  NOR U96400 ( .A(n76231), .B(n79579), .Z(n79573) );
  IV U96401 ( .A(n76232), .Z(n76234) );
  NOR U96402 ( .A(n76234), .B(n76233), .Z(n79570) );
  IV U96403 ( .A(n79570), .Z(n79565) );
  IV U96404 ( .A(n76235), .Z(n76236) );
  NOR U96405 ( .A(n76236), .B(n79567), .Z(n81772) );
  IV U96406 ( .A(n76237), .Z(n76239) );
  NOR U96407 ( .A(n76239), .B(n76238), .Z(n76244) );
  IV U96408 ( .A(n76240), .Z(n76242) );
  NOR U96409 ( .A(n76242), .B(n76241), .Z(n76243) );
  NOR U96410 ( .A(n76244), .B(n76243), .Z(n81771) );
  IV U96411 ( .A(n76245), .Z(n76246) );
  NOR U96412 ( .A(n76247), .B(n76246), .Z(n76252) );
  IV U96413 ( .A(n76248), .Z(n76250) );
  NOR U96414 ( .A(n76250), .B(n76249), .Z(n76251) );
  NOR U96415 ( .A(n76252), .B(n76251), .Z(n85362) );
  IV U96416 ( .A(n76253), .Z(n76256) );
  NOR U96417 ( .A(n76254), .B(n76261), .Z(n76255) );
  IV U96418 ( .A(n76255), .Z(n76258) );
  NOR U96419 ( .A(n76256), .B(n76258), .Z(n85363) );
  IV U96420 ( .A(n76257), .Z(n76259) );
  NOR U96421 ( .A(n76259), .B(n76258), .Z(n81780) );
  IV U96422 ( .A(n76260), .Z(n76264) );
  NOR U96423 ( .A(n76262), .B(n76261), .Z(n76263) );
  IV U96424 ( .A(n76263), .Z(n76266) );
  NOR U96425 ( .A(n76264), .B(n76266), .Z(n81777) );
  IV U96426 ( .A(n76265), .Z(n76267) );
  NOR U96427 ( .A(n76267), .B(n76266), .Z(n85352) );
  IV U96428 ( .A(n76268), .Z(n76269) );
  NOR U96429 ( .A(n76270), .B(n76269), .Z(n85355) );
  IV U96430 ( .A(n76271), .Z(n76274) );
  NOR U96431 ( .A(n76277), .B(n76280), .Z(n76272) );
  IV U96432 ( .A(n76272), .Z(n76273) );
  NOR U96433 ( .A(n76274), .B(n76273), .Z(n81783) );
  NOR U96434 ( .A(n85355), .B(n81783), .Z(n76275) );
  IV U96435 ( .A(n76275), .Z(n79563) );
  NOR U96436 ( .A(n76276), .B(n76280), .Z(n81787) );
  NOR U96437 ( .A(n76278), .B(n76277), .Z(n76279) );
  IV U96438 ( .A(n76279), .Z(n76281) );
  NOR U96439 ( .A(n76281), .B(n76280), .Z(n85349) );
  NOR U96440 ( .A(n81787), .B(n85349), .Z(n79562) );
  IV U96441 ( .A(n76282), .Z(n76283) );
  NOR U96442 ( .A(n76284), .B(n76283), .Z(n79560) );
  IV U96443 ( .A(n79560), .Z(n79555) );
  IV U96444 ( .A(n76285), .Z(n76287) );
  IV U96445 ( .A(n76286), .Z(n79557) );
  NOR U96446 ( .A(n76287), .B(n79557), .Z(n85342) );
  IV U96447 ( .A(n76288), .Z(n76289) );
  NOR U96448 ( .A(n76289), .B(n85329), .Z(n79542) );
  IV U96449 ( .A(n76290), .Z(n76292) );
  IV U96450 ( .A(n76291), .Z(n79534) );
  NOR U96451 ( .A(n76292), .B(n79534), .Z(n81796) );
  IV U96452 ( .A(n76293), .Z(n79518) );
  IV U96453 ( .A(n79517), .Z(n76295) );
  NOR U96454 ( .A(n79518), .B(n76295), .Z(n81814) );
  IV U96455 ( .A(n76294), .Z(n76298) );
  NOR U96456 ( .A(n76296), .B(n76295), .Z(n76297) );
  IV U96457 ( .A(n76297), .Z(n79514) );
  NOR U96458 ( .A(n76298), .B(n79514), .Z(n85299) );
  NOR U96459 ( .A(n81814), .B(n85299), .Z(n79512) );
  IV U96460 ( .A(n76299), .Z(n76300) );
  NOR U96461 ( .A(n76301), .B(n76300), .Z(n81811) );
  IV U96462 ( .A(n81811), .Z(n81812) );
  IV U96463 ( .A(n76302), .Z(n76306) );
  IV U96464 ( .A(n76303), .Z(n79502) );
  NOR U96465 ( .A(n76304), .B(n79502), .Z(n76305) );
  IV U96466 ( .A(n76305), .Z(n79506) );
  NOR U96467 ( .A(n76306), .B(n79506), .Z(n85288) );
  IV U96468 ( .A(n76307), .Z(n79479) );
  IV U96469 ( .A(n76308), .Z(n76309) );
  NOR U96470 ( .A(n79479), .B(n76309), .Z(n81839) );
  IV U96471 ( .A(n76310), .Z(n76312) );
  NOR U96472 ( .A(n76312), .B(n76311), .Z(n79473) );
  IV U96473 ( .A(n76313), .Z(n76314) );
  NOR U96474 ( .A(n76314), .B(n79462), .Z(n79470) );
  IV U96475 ( .A(n79470), .Z(n79460) );
  IV U96476 ( .A(n76315), .Z(n76316) );
  NOR U96477 ( .A(n79439), .B(n76316), .Z(n81855) );
  IV U96478 ( .A(n76317), .Z(n76318) );
  NOR U96479 ( .A(n76319), .B(n76318), .Z(n85258) );
  NOR U96480 ( .A(n81855), .B(n85258), .Z(n79436) );
  IV U96481 ( .A(n76320), .Z(n76322) );
  IV U96482 ( .A(n76321), .Z(n79428) );
  NOR U96483 ( .A(n76322), .B(n79428), .Z(n81854) );
  IV U96484 ( .A(n81854), .Z(n81852) );
  IV U96485 ( .A(n76323), .Z(n76326) );
  NOR U96486 ( .A(n79411), .B(n76324), .Z(n76325) );
  IV U96487 ( .A(n76325), .Z(n76328) );
  NOR U96488 ( .A(n76326), .B(n76328), .Z(n81866) );
  IV U96489 ( .A(n76327), .Z(n76329) );
  NOR U96490 ( .A(n76329), .B(n76328), .Z(n81863) );
  IV U96491 ( .A(n76330), .Z(n76331) );
  NOR U96492 ( .A(n76332), .B(n76331), .Z(n81882) );
  IV U96493 ( .A(n76333), .Z(n76334) );
  NOR U96494 ( .A(n76334), .B(n79398), .Z(n85246) );
  NOR U96495 ( .A(n81882), .B(n85246), .Z(n79396) );
  IV U96496 ( .A(n76335), .Z(n76337) );
  NOR U96497 ( .A(n76337), .B(n76336), .Z(n85239) );
  IV U96498 ( .A(n76338), .Z(n76339) );
  NOR U96499 ( .A(n76340), .B(n76339), .Z(n81900) );
  IV U96500 ( .A(n76341), .Z(n76342) );
  NOR U96501 ( .A(n79387), .B(n76342), .Z(n81897) );
  NOR U96502 ( .A(n81900), .B(n81897), .Z(n76343) );
  IV U96503 ( .A(n76343), .Z(n79390) );
  IV U96504 ( .A(n76344), .Z(n81905) );
  NOR U96505 ( .A(n81905), .B(n76345), .Z(n79385) );
  IV U96506 ( .A(n76346), .Z(n76347) );
  NOR U96507 ( .A(n76350), .B(n76347), .Z(n76348) );
  IV U96508 ( .A(n76348), .Z(n81912) );
  IV U96509 ( .A(n76349), .Z(n76351) );
  NOR U96510 ( .A(n76351), .B(n76350), .Z(n79381) );
  NOR U96511 ( .A(n76352), .B(n81923), .Z(n79371) );
  IV U96512 ( .A(n76353), .Z(n76354) );
  NOR U96513 ( .A(n79369), .B(n76354), .Z(n85216) );
  IV U96514 ( .A(n76355), .Z(n76357) );
  NOR U96515 ( .A(n76357), .B(n76356), .Z(n85203) );
  IV U96516 ( .A(n76358), .Z(n76360) );
  IV U96517 ( .A(n76359), .Z(n79365) );
  NOR U96518 ( .A(n76360), .B(n79365), .Z(n81930) );
  NOR U96519 ( .A(n85203), .B(n81930), .Z(n79363) );
  IV U96520 ( .A(n76361), .Z(n76363) );
  NOR U96521 ( .A(n76363), .B(n76362), .Z(n76365) );
  NOR U96522 ( .A(n76365), .B(n76364), .Z(n85207) );
  IV U96523 ( .A(n76366), .Z(n76367) );
  NOR U96524 ( .A(n76367), .B(n76371), .Z(n85200) );
  NOR U96525 ( .A(n85209), .B(n85200), .Z(n79362) );
  IV U96526 ( .A(n76368), .Z(n76369) );
  NOR U96527 ( .A(n76369), .B(n76371), .Z(n81935) );
  IV U96528 ( .A(n76370), .Z(n76372) );
  NOR U96529 ( .A(n76372), .B(n76371), .Z(n85187) );
  IV U96530 ( .A(n76373), .Z(n76375) );
  NOR U96531 ( .A(n76375), .B(n76374), .Z(n85191) );
  IV U96532 ( .A(n76376), .Z(n76378) );
  NOR U96533 ( .A(n76378), .B(n76377), .Z(n76383) );
  IV U96534 ( .A(n76379), .Z(n76381) );
  NOR U96535 ( .A(n76381), .B(n76380), .Z(n76382) );
  NOR U96536 ( .A(n76383), .B(n76382), .Z(n85180) );
  IV U96537 ( .A(n76384), .Z(n76386) );
  IV U96538 ( .A(n76385), .Z(n76389) );
  NOR U96539 ( .A(n76386), .B(n76389), .Z(n81950) );
  NOR U96540 ( .A(n76387), .B(n81963), .Z(n76391) );
  IV U96541 ( .A(n76388), .Z(n76390) );
  NOR U96542 ( .A(n76390), .B(n76389), .Z(n81958) );
  NOR U96543 ( .A(n76391), .B(n81958), .Z(n79340) );
  IV U96544 ( .A(n76392), .Z(n81989) );
  IV U96545 ( .A(n76393), .Z(n76394) );
  NOR U96546 ( .A(n76397), .B(n76394), .Z(n81993) );
  IV U96547 ( .A(n76395), .Z(n76396) );
  NOR U96548 ( .A(n76397), .B(n76396), .Z(n81990) );
  IV U96549 ( .A(n76398), .Z(n76399) );
  NOR U96550 ( .A(n76399), .B(n79310), .Z(n79317) );
  IV U96551 ( .A(n76400), .Z(n76403) );
  NOR U96552 ( .A(n76406), .B(n76401), .Z(n76402) );
  IV U96553 ( .A(n76402), .Z(n79313) );
  NOR U96554 ( .A(n76403), .B(n79313), .Z(n85162) );
  IV U96555 ( .A(n76404), .Z(n76405) );
  NOR U96556 ( .A(n76406), .B(n76405), .Z(n85159) );
  IV U96557 ( .A(n76407), .Z(n76410) );
  IV U96558 ( .A(n76408), .Z(n76409) );
  NOR U96559 ( .A(n76410), .B(n76409), .Z(n82001) );
  IV U96560 ( .A(n76411), .Z(n76414) );
  IV U96561 ( .A(n76412), .Z(n76413) );
  NOR U96562 ( .A(n76414), .B(n76413), .Z(n85155) );
  IV U96563 ( .A(n76415), .Z(n76417) );
  IV U96564 ( .A(n76416), .Z(n79295) );
  NOR U96565 ( .A(n76417), .B(n79295), .Z(n82006) );
  IV U96566 ( .A(n76418), .Z(n76419) );
  NOR U96567 ( .A(n76419), .B(n76424), .Z(n82009) );
  IV U96568 ( .A(n76420), .Z(n76421) );
  NOR U96569 ( .A(n76422), .B(n76421), .Z(n85137) );
  IV U96570 ( .A(n76423), .Z(n76425) );
  NOR U96571 ( .A(n76425), .B(n76424), .Z(n82012) );
  NOR U96572 ( .A(n85137), .B(n82012), .Z(n76426) );
  IV U96573 ( .A(n76426), .Z(n79293) );
  IV U96574 ( .A(n76427), .Z(n82017) );
  NOR U96575 ( .A(n82017), .B(n76428), .Z(n85128) );
  IV U96576 ( .A(n76429), .Z(n76431) );
  NOR U96577 ( .A(n76431), .B(n76430), .Z(n82023) );
  IV U96578 ( .A(n76432), .Z(n76435) );
  NOR U96579 ( .A(n76433), .B(n76440), .Z(n76434) );
  IV U96580 ( .A(n76434), .Z(n76437) );
  NOR U96581 ( .A(n76435), .B(n76437), .Z(n82034) );
  IV U96582 ( .A(n76436), .Z(n76438) );
  NOR U96583 ( .A(n76438), .B(n76437), .Z(n82031) );
  IV U96584 ( .A(n76439), .Z(n76441) );
  NOR U96585 ( .A(n76441), .B(n76440), .Z(n82052) );
  IV U96586 ( .A(n76442), .Z(n76443) );
  NOR U96587 ( .A(n76443), .B(n82043), .Z(n76444) );
  NOR U96588 ( .A(n82052), .B(n76444), .Z(n76445) );
  IV U96589 ( .A(n76445), .Z(n79292) );
  IV U96590 ( .A(n76448), .Z(n82057) );
  NOR U96591 ( .A(n82057), .B(n76446), .Z(n76452) );
  IV U96592 ( .A(n76447), .Z(n76451) );
  NOR U96593 ( .A(n76454), .B(n76448), .Z(n76449) );
  IV U96594 ( .A(n76449), .Z(n76450) );
  NOR U96595 ( .A(n76451), .B(n76450), .Z(n82060) );
  NOR U96596 ( .A(n76452), .B(n82060), .Z(n79291) );
  IV U96597 ( .A(n76453), .Z(n76457) );
  NOR U96598 ( .A(n76454), .B(n79283), .Z(n76455) );
  IV U96599 ( .A(n76455), .Z(n76456) );
  NOR U96600 ( .A(n76457), .B(n76456), .Z(n79286) );
  IV U96601 ( .A(n76458), .Z(n76459) );
  NOR U96602 ( .A(n76459), .B(n76461), .Z(n79278) );
  IV U96603 ( .A(n76460), .Z(n76462) );
  NOR U96604 ( .A(n76462), .B(n76461), .Z(n79276) );
  IV U96605 ( .A(n79276), .Z(n79271) );
  IV U96606 ( .A(n76463), .Z(n76465) );
  IV U96607 ( .A(n76464), .Z(n76467) );
  NOR U96608 ( .A(n76465), .B(n76467), .Z(n85104) );
  IV U96609 ( .A(n76466), .Z(n76468) );
  NOR U96610 ( .A(n76468), .B(n76467), .Z(n85099) );
  IV U96611 ( .A(n76469), .Z(n76470) );
  NOR U96612 ( .A(n76472), .B(n76470), .Z(n82088) );
  IV U96613 ( .A(n76471), .Z(n76473) );
  NOR U96614 ( .A(n76473), .B(n76472), .Z(n82097) );
  IV U96615 ( .A(n76474), .Z(n79243) );
  IV U96616 ( .A(n76475), .Z(n76476) );
  NOR U96617 ( .A(n79243), .B(n76476), .Z(n82101) );
  IV U96618 ( .A(n76477), .Z(n76478) );
  NOR U96619 ( .A(n76478), .B(n76483), .Z(n82103) );
  NOR U96620 ( .A(n82101), .B(n82103), .Z(n79240) );
  IV U96621 ( .A(n76479), .Z(n76481) );
  NOR U96622 ( .A(n76481), .B(n76480), .Z(n82110) );
  IV U96623 ( .A(n76482), .Z(n76484) );
  NOR U96624 ( .A(n76484), .B(n76483), .Z(n82106) );
  NOR U96625 ( .A(n82110), .B(n82106), .Z(n79239) );
  IV U96626 ( .A(n76485), .Z(n76486) );
  NOR U96627 ( .A(n76486), .B(n76488), .Z(n82121) );
  IV U96628 ( .A(n76487), .Z(n76489) );
  NOR U96629 ( .A(n76489), .B(n76488), .Z(n82124) );
  NOR U96630 ( .A(n82121), .B(n82124), .Z(n82109) );
  IV U96631 ( .A(n82109), .Z(n76493) );
  IV U96632 ( .A(n76490), .Z(n82115) );
  NOR U96633 ( .A(n76491), .B(n82115), .Z(n76492) );
  NOR U96634 ( .A(n76493), .B(n76492), .Z(n79238) );
  IV U96635 ( .A(n76494), .Z(n76496) );
  NOR U96636 ( .A(n76496), .B(n76495), .Z(n79236) );
  IV U96637 ( .A(n79236), .Z(n79231) );
  IV U96638 ( .A(n76497), .Z(n82129) );
  IV U96639 ( .A(n76498), .Z(n76499) );
  NOR U96640 ( .A(n76499), .B(n76501), .Z(n85083) );
  IV U96641 ( .A(n76500), .Z(n76502) );
  NOR U96642 ( .A(n76502), .B(n76501), .Z(n85080) );
  IV U96643 ( .A(n76503), .Z(n76504) );
  NOR U96644 ( .A(n76504), .B(n79217), .Z(n85059) );
  IV U96645 ( .A(n76505), .Z(n76506) );
  NOR U96646 ( .A(n76507), .B(n76506), .Z(n82140) );
  NOR U96647 ( .A(n76508), .B(n82137), .Z(n76509) );
  NOR U96648 ( .A(n82140), .B(n76509), .Z(n79214) );
  IV U96649 ( .A(n76510), .Z(n76517) );
  IV U96650 ( .A(n76511), .Z(n76512) );
  NOR U96651 ( .A(n76517), .B(n76512), .Z(n85051) );
  IV U96652 ( .A(n76513), .Z(n76514) );
  NOR U96653 ( .A(n76519), .B(n76514), .Z(n85046) );
  IV U96654 ( .A(n76515), .Z(n76516) );
  NOR U96655 ( .A(n76517), .B(n76516), .Z(n85055) );
  NOR U96656 ( .A(n85046), .B(n85055), .Z(n90746) );
  IV U96657 ( .A(n76518), .Z(n76520) );
  NOR U96658 ( .A(n76520), .B(n76519), .Z(n76521) );
  IV U96659 ( .A(n76521), .Z(n79210) );
  IV U96660 ( .A(n76522), .Z(n79206) );
  IV U96661 ( .A(n76523), .Z(n76524) );
  NOR U96662 ( .A(n79206), .B(n76524), .Z(n76525) );
  IV U96663 ( .A(n76525), .Z(n85033) );
  IV U96664 ( .A(n76526), .Z(n76528) );
  NOR U96665 ( .A(n76528), .B(n76527), .Z(n85023) );
  IV U96666 ( .A(n76529), .Z(n76530) );
  NOR U96667 ( .A(n76530), .B(n79200), .Z(n85030) );
  NOR U96668 ( .A(n85023), .B(n85030), .Z(n79203) );
  IV U96669 ( .A(n76531), .Z(n76532) );
  NOR U96670 ( .A(n79196), .B(n76532), .Z(n79192) );
  IV U96671 ( .A(n79192), .Z(n79180) );
  NOR U96672 ( .A(n76533), .B(n82159), .Z(n79184) );
  IV U96673 ( .A(n76534), .Z(n76537) );
  NOR U96674 ( .A(n76542), .B(n76535), .Z(n76536) );
  IV U96675 ( .A(n76536), .Z(n79168) );
  NOR U96676 ( .A(n76537), .B(n79168), .Z(n84995) );
  IV U96677 ( .A(n76538), .Z(n76539) );
  NOR U96678 ( .A(n76539), .B(n79153), .Z(n84991) );
  IV U96679 ( .A(n76540), .Z(n76541) );
  NOR U96680 ( .A(n76542), .B(n76541), .Z(n82162) );
  NOR U96681 ( .A(n84991), .B(n82162), .Z(n79163) );
  IV U96682 ( .A(n76543), .Z(n76545) );
  NOR U96683 ( .A(n76545), .B(n76544), .Z(n82168) );
  IV U96684 ( .A(n76546), .Z(n76548) );
  IV U96685 ( .A(n76547), .Z(n76550) );
  NOR U96686 ( .A(n76548), .B(n76550), .Z(n84983) );
  IV U96687 ( .A(n76549), .Z(n76551) );
  NOR U96688 ( .A(n76551), .B(n76550), .Z(n82171) );
  IV U96689 ( .A(n76552), .Z(n76553) );
  NOR U96690 ( .A(n76554), .B(n76553), .Z(n84976) );
  IV U96691 ( .A(n76555), .Z(n76558) );
  NOR U96692 ( .A(n79141), .B(n76556), .Z(n76557) );
  IV U96693 ( .A(n76557), .Z(n76560) );
  NOR U96694 ( .A(n76558), .B(n76560), .Z(n84973) );
  IV U96695 ( .A(n76559), .Z(n76561) );
  NOR U96696 ( .A(n76561), .B(n76560), .Z(n82177) );
  XOR U96697 ( .A(n82186), .B(n76562), .Z(n76565) );
  IV U96698 ( .A(n76563), .Z(n76564) );
  NOR U96699 ( .A(n76565), .B(n76564), .Z(n84945) );
  IV U96700 ( .A(n76566), .Z(n76567) );
  NOR U96701 ( .A(n76568), .B(n76567), .Z(n82204) );
  IV U96702 ( .A(n76569), .Z(n76570) );
  NOR U96703 ( .A(n76571), .B(n76570), .Z(n82201) );
  NOR U96704 ( .A(n82204), .B(n82201), .Z(n79123) );
  IV U96705 ( .A(n76572), .Z(n76573) );
  NOR U96706 ( .A(n76574), .B(n76573), .Z(n82209) );
  IV U96707 ( .A(n76575), .Z(n76577) );
  NOR U96708 ( .A(n76577), .B(n76576), .Z(n84900) );
  IV U96709 ( .A(n76578), .Z(n76580) );
  NOR U96710 ( .A(n76580), .B(n76579), .Z(n79084) );
  IV U96711 ( .A(n76581), .Z(n76583) );
  NOR U96712 ( .A(n76583), .B(n76582), .Z(n84852) );
  IV U96713 ( .A(n76584), .Z(n76586) );
  NOR U96714 ( .A(n76586), .B(n76585), .Z(n82238) );
  IV U96715 ( .A(n76587), .Z(n76588) );
  NOR U96716 ( .A(n76588), .B(n76597), .Z(n82250) );
  IV U96717 ( .A(n76589), .Z(n76590) );
  NOR U96718 ( .A(n76591), .B(n76590), .Z(n82243) );
  NOR U96719 ( .A(n82250), .B(n82243), .Z(n76592) );
  IV U96720 ( .A(n76592), .Z(n79061) );
  IV U96721 ( .A(n76593), .Z(n76595) );
  NOR U96722 ( .A(n76595), .B(n76594), .Z(n82254) );
  IV U96723 ( .A(n76596), .Z(n76598) );
  NOR U96724 ( .A(n76598), .B(n76597), .Z(n82248) );
  NOR U96725 ( .A(n82254), .B(n82248), .Z(n79060) );
  IV U96726 ( .A(n76599), .Z(n76601) );
  NOR U96727 ( .A(n76601), .B(n76600), .Z(n82260) );
  IV U96728 ( .A(n76602), .Z(n76604) );
  NOR U96729 ( .A(n76604), .B(n76603), .Z(n82257) );
  NOR U96730 ( .A(n82260), .B(n82257), .Z(n79059) );
  IV U96731 ( .A(n76605), .Z(n84824) );
  NOR U96732 ( .A(n84824), .B(n76606), .Z(n79058) );
  IV U96733 ( .A(n76607), .Z(n76608) );
  NOR U96734 ( .A(n76608), .B(n76610), .Z(n84817) );
  IV U96735 ( .A(n76609), .Z(n76613) );
  NOR U96736 ( .A(n76611), .B(n76610), .Z(n76612) );
  IV U96737 ( .A(n76612), .Z(n79051) );
  NOR U96738 ( .A(n76613), .B(n79051), .Z(n79055) );
  IV U96739 ( .A(n79055), .Z(n79044) );
  IV U96740 ( .A(n76614), .Z(n76619) );
  IV U96741 ( .A(n76615), .Z(n76616) );
  NOR U96742 ( .A(n76619), .B(n76616), .Z(n82269) );
  IV U96743 ( .A(n76617), .Z(n76618) );
  NOR U96744 ( .A(n76619), .B(n76618), .Z(n76620) );
  IV U96745 ( .A(n76620), .Z(n82277) );
  IV U96746 ( .A(n76621), .Z(n76622) );
  NOR U96747 ( .A(n76622), .B(n79021), .Z(n84799) );
  IV U96748 ( .A(n76623), .Z(n76628) );
  IV U96749 ( .A(n76624), .Z(n76625) );
  NOR U96750 ( .A(n76625), .B(n79021), .Z(n76626) );
  IV U96751 ( .A(n76626), .Z(n76627) );
  NOR U96752 ( .A(n76628), .B(n76627), .Z(n84796) );
  IV U96753 ( .A(n76629), .Z(n76630) );
  NOR U96754 ( .A(n76630), .B(n76633), .Z(n82288) );
  IV U96755 ( .A(n76631), .Z(n76632) );
  NOR U96756 ( .A(n76633), .B(n76632), .Z(n82296) );
  IV U96757 ( .A(n76634), .Z(n76635) );
  NOR U96758 ( .A(n76636), .B(n76635), .Z(n76637) );
  IV U96759 ( .A(n76637), .Z(n76641) );
  NOR U96760 ( .A(n76645), .B(n76638), .Z(n76639) );
  IV U96761 ( .A(n76639), .Z(n76640) );
  NOR U96762 ( .A(n76641), .B(n76640), .Z(n82300) );
  IV U96763 ( .A(n76642), .Z(n76648) );
  IV U96764 ( .A(n76643), .Z(n76644) );
  NOR U96765 ( .A(n76645), .B(n76644), .Z(n76646) );
  IV U96766 ( .A(n76646), .Z(n76647) );
  NOR U96767 ( .A(n76648), .B(n76647), .Z(n84792) );
  IV U96768 ( .A(n76649), .Z(n76650) );
  NOR U96769 ( .A(n76655), .B(n76650), .Z(n84780) );
  IV U96770 ( .A(n76651), .Z(n84772) );
  NOR U96771 ( .A(n76652), .B(n84772), .Z(n76656) );
  IV U96772 ( .A(n76653), .Z(n76654) );
  NOR U96773 ( .A(n76655), .B(n76654), .Z(n84783) );
  NOR U96774 ( .A(n76656), .B(n84783), .Z(n76657) );
  IV U96775 ( .A(n76657), .Z(n79018) );
  IV U96776 ( .A(n76658), .Z(n76659) );
  NOR U96777 ( .A(n76659), .B(n76668), .Z(n76663) );
  IV U96778 ( .A(n76660), .Z(n76661) );
  NOR U96779 ( .A(n76661), .B(n84772), .Z(n76662) );
  NOR U96780 ( .A(n76663), .B(n76662), .Z(n84769) );
  IV U96781 ( .A(n76664), .Z(n76665) );
  NOR U96782 ( .A(n76666), .B(n76665), .Z(n84761) );
  IV U96783 ( .A(n76667), .Z(n76669) );
  NOR U96784 ( .A(n76669), .B(n76668), .Z(n84765) );
  NOR U96785 ( .A(n84761), .B(n84765), .Z(n79017) );
  NOR U96786 ( .A(n76670), .B(n82303), .Z(n79016) );
  IV U96787 ( .A(n76671), .Z(n76673) );
  IV U96788 ( .A(n76672), .Z(n79015) );
  NOR U96789 ( .A(n76673), .B(n79015), .Z(n79009) );
  IV U96790 ( .A(n79009), .Z(n79007) );
  NOR U96791 ( .A(n76675), .B(n76674), .Z(n84736) );
  IV U96792 ( .A(n76676), .Z(n76678) );
  IV U96793 ( .A(n76677), .Z(n76680) );
  NOR U96794 ( .A(n76678), .B(n76680), .Z(n84733) );
  IV U96795 ( .A(n76679), .Z(n76681) );
  NOR U96796 ( .A(n76681), .B(n76680), .Z(n84729) );
  IV U96797 ( .A(n76682), .Z(n76683) );
  NOR U96798 ( .A(n76683), .B(n76689), .Z(n76684) );
  IV U96799 ( .A(n76684), .Z(n84728) );
  IV U96800 ( .A(n76685), .Z(n76686) );
  NOR U96801 ( .A(n76687), .B(n76686), .Z(n88111) );
  IV U96802 ( .A(n76688), .Z(n76690) );
  NOR U96803 ( .A(n76690), .B(n76689), .Z(n88136) );
  NOR U96804 ( .A(n88111), .B(n88136), .Z(n82308) );
  NOR U96805 ( .A(n76691), .B(n82319), .Z(n82309) );
  IV U96806 ( .A(n76692), .Z(n76697) );
  IV U96807 ( .A(n76693), .Z(n76694) );
  NOR U96808 ( .A(n76697), .B(n76694), .Z(n84709) );
  IV U96809 ( .A(n76695), .Z(n76699) );
  NOR U96810 ( .A(n76697), .B(n76696), .Z(n76698) );
  IV U96811 ( .A(n76698), .Z(n78983) );
  NOR U96812 ( .A(n76699), .B(n78983), .Z(n82326) );
  NOR U96813 ( .A(n84709), .B(n82326), .Z(n78987) );
  IV U96814 ( .A(n76700), .Z(n76701) );
  NOR U96815 ( .A(n76704), .B(n76701), .Z(n82336) );
  IV U96816 ( .A(n82336), .Z(n82334) );
  IV U96817 ( .A(n76702), .Z(n76703) );
  NOR U96818 ( .A(n76704), .B(n76703), .Z(n76705) );
  IV U96819 ( .A(n76705), .Z(n84706) );
  IV U96820 ( .A(n76706), .Z(n76711) );
  IV U96821 ( .A(n76707), .Z(n76708) );
  NOR U96822 ( .A(n76711), .B(n76708), .Z(n84696) );
  IV U96823 ( .A(n76709), .Z(n76710) );
  NOR U96824 ( .A(n76711), .B(n76710), .Z(n82349) );
  IV U96825 ( .A(n76712), .Z(n76714) );
  NOR U96826 ( .A(n76714), .B(n76713), .Z(n82346) );
  IV U96827 ( .A(n76715), .Z(n76717) );
  IV U96828 ( .A(n76716), .Z(n76718) );
  NOR U96829 ( .A(n76717), .B(n76718), .Z(n82343) );
  NOR U96830 ( .A(n76719), .B(n76718), .Z(n84690) );
  IV U96831 ( .A(n76720), .Z(n76721) );
  NOR U96832 ( .A(n76721), .B(n76726), .Z(n84687) );
  IV U96833 ( .A(n76722), .Z(n76724) );
  NOR U96834 ( .A(n76724), .B(n76723), .Z(n84684) );
  IV U96835 ( .A(n76725), .Z(n76727) );
  NOR U96836 ( .A(n76727), .B(n76726), .Z(n82357) );
  NOR U96837 ( .A(n84684), .B(n82357), .Z(n78967) );
  IV U96838 ( .A(n76728), .Z(n76729) );
  NOR U96839 ( .A(n76732), .B(n76729), .Z(n82362) );
  IV U96840 ( .A(n76730), .Z(n76731) );
  NOR U96841 ( .A(n76732), .B(n76731), .Z(n82360) );
  IV U96842 ( .A(n76733), .Z(n76734) );
  NOR U96843 ( .A(n76734), .B(n76739), .Z(n84668) );
  IV U96844 ( .A(n76735), .Z(n76737) );
  NOR U96845 ( .A(n76737), .B(n76736), .Z(n82383) );
  IV U96846 ( .A(n76738), .Z(n76740) );
  NOR U96847 ( .A(n76740), .B(n76739), .Z(n82379) );
  NOR U96848 ( .A(n82383), .B(n82379), .Z(n78955) );
  IV U96849 ( .A(n76741), .Z(n76742) );
  NOR U96850 ( .A(n76743), .B(n76742), .Z(n76744) );
  IV U96851 ( .A(n76744), .Z(n82385) );
  NOR U96852 ( .A(n76745), .B(n84657), .Z(n82393) );
  IV U96853 ( .A(n76746), .Z(n76747) );
  NOR U96854 ( .A(n76748), .B(n76747), .Z(n82392) );
  NOR U96855 ( .A(n82393), .B(n82392), .Z(n78947) );
  IV U96856 ( .A(n76749), .Z(n76750) );
  NOR U96857 ( .A(n76751), .B(n76750), .Z(n78945) );
  IV U96858 ( .A(n78945), .Z(n78940) );
  IV U96859 ( .A(n76752), .Z(n76753) );
  NOR U96860 ( .A(n76754), .B(n76753), .Z(n84650) );
  IV U96861 ( .A(n76755), .Z(n76756) );
  NOR U96862 ( .A(n78930), .B(n76756), .Z(n82400) );
  IV U96863 ( .A(n76757), .Z(n78932) );
  IV U96864 ( .A(n76758), .Z(n76759) );
  NOR U96865 ( .A(n78932), .B(n76759), .Z(n82407) );
  NOR U96866 ( .A(n82400), .B(n82407), .Z(n78927) );
  IV U96867 ( .A(n76760), .Z(n76761) );
  NOR U96868 ( .A(n76764), .B(n76761), .Z(n82410) );
  IV U96869 ( .A(n76762), .Z(n76763) );
  NOR U96870 ( .A(n76764), .B(n76763), .Z(n84636) );
  IV U96871 ( .A(n76765), .Z(n76766) );
  NOR U96872 ( .A(n76768), .B(n76766), .Z(n78892) );
  IV U96873 ( .A(n76767), .Z(n76769) );
  NOR U96874 ( .A(n76769), .B(n76768), .Z(n78890) );
  IV U96875 ( .A(n78890), .Z(n78885) );
  IV U96876 ( .A(n76770), .Z(n76773) );
  NOR U96877 ( .A(n76782), .B(n76775), .Z(n76771) );
  IV U96878 ( .A(n76771), .Z(n76772) );
  NOR U96879 ( .A(n76773), .B(n76772), .Z(n82442) );
  IV U96880 ( .A(n76774), .Z(n76779) );
  XOR U96881 ( .A(n76780), .B(n76782), .Z(n76776) );
  NOR U96882 ( .A(n76776), .B(n76775), .Z(n76777) );
  IV U96883 ( .A(n76777), .Z(n76778) );
  NOR U96884 ( .A(n76779), .B(n76778), .Z(n84608) );
  IV U96885 ( .A(n76780), .Z(n76781) );
  NOR U96886 ( .A(n76782), .B(n76781), .Z(n76783) );
  IV U96887 ( .A(n76783), .Z(n76784) );
  NOR U96888 ( .A(n76785), .B(n76784), .Z(n84605) );
  NOR U96889 ( .A(n76787), .B(n76786), .Z(n76789) );
  NOR U96890 ( .A(n76789), .B(n76788), .Z(n76790) );
  NOR U96891 ( .A(n76791), .B(n76790), .Z(n82445) );
  IV U96892 ( .A(n76792), .Z(n76794) );
  NOR U96893 ( .A(n76794), .B(n76793), .Z(n78863) );
  IV U96894 ( .A(n78863), .Z(n78856) );
  IV U96895 ( .A(n76795), .Z(n76800) );
  IV U96896 ( .A(n76796), .Z(n76797) );
  NOR U96897 ( .A(n76800), .B(n76797), .Z(n82466) );
  IV U96898 ( .A(n76798), .Z(n76799) );
  NOR U96899 ( .A(n76800), .B(n76799), .Z(n76801) );
  IV U96900 ( .A(n76801), .Z(n82469) );
  IV U96901 ( .A(n76802), .Z(n76809) );
  IV U96902 ( .A(n76803), .Z(n76804) );
  NOR U96903 ( .A(n76809), .B(n76804), .Z(n82475) );
  IV U96904 ( .A(n76805), .Z(n76807) );
  NOR U96905 ( .A(n76807), .B(n76806), .Z(n82471) );
  NOR U96906 ( .A(n76809), .B(n76808), .Z(n82480) );
  NOR U96907 ( .A(n82471), .B(n82480), .Z(n76810) );
  IV U96908 ( .A(n76810), .Z(n76811) );
  NOR U96909 ( .A(n82475), .B(n76811), .Z(n78833) );
  IV U96910 ( .A(n76812), .Z(n76814) );
  NOR U96911 ( .A(n76814), .B(n76813), .Z(n82482) );
  IV U96912 ( .A(n82482), .Z(n82479) );
  IV U96913 ( .A(n78829), .Z(n78817) );
  IV U96914 ( .A(n76815), .Z(n78830) );
  NOR U96915 ( .A(n78817), .B(n78830), .Z(n76816) );
  IV U96916 ( .A(n76816), .Z(n78823) );
  IV U96917 ( .A(n76820), .Z(n76818) );
  NOR U96918 ( .A(n76818), .B(n76817), .Z(n90391) );
  NOR U96919 ( .A(n76820), .B(n76819), .Z(n76823) );
  IV U96920 ( .A(n76821), .Z(n76822) );
  NOR U96921 ( .A(n76823), .B(n76822), .Z(n76824) );
  NOR U96922 ( .A(n90391), .B(n76824), .Z(n84573) );
  IV U96923 ( .A(n76825), .Z(n76826) );
  NOR U96924 ( .A(n76826), .B(n76828), .Z(n84569) );
  IV U96925 ( .A(n76827), .Z(n76829) );
  NOR U96926 ( .A(n76829), .B(n76828), .Z(n84566) );
  IV U96927 ( .A(n76830), .Z(n82498) );
  NOR U96928 ( .A(n82498), .B(n76831), .Z(n76834) );
  IV U96929 ( .A(n76832), .Z(n76833) );
  NOR U96930 ( .A(n76833), .B(n76836), .Z(n84558) );
  NOR U96931 ( .A(n76834), .B(n84558), .Z(n78815) );
  IV U96932 ( .A(n76835), .Z(n76837) );
  NOR U96933 ( .A(n76837), .B(n76836), .Z(n78811) );
  IV U96934 ( .A(n76838), .Z(n78808) );
  IV U96935 ( .A(n76839), .Z(n76840) );
  NOR U96936 ( .A(n78808), .B(n76840), .Z(n84551) );
  IV U96937 ( .A(n76841), .Z(n76843) );
  NOR U96938 ( .A(n76843), .B(n76842), .Z(n76844) );
  IV U96939 ( .A(n76844), .Z(n82504) );
  IV U96940 ( .A(n76845), .Z(n76846) );
  NOR U96941 ( .A(n76846), .B(n76848), .Z(n82507) );
  IV U96942 ( .A(n76847), .Z(n76849) );
  NOR U96943 ( .A(n76849), .B(n76848), .Z(n84518) );
  IV U96944 ( .A(n76850), .Z(n76851) );
  NOR U96945 ( .A(n76852), .B(n76851), .Z(n82509) );
  NOR U96946 ( .A(n84518), .B(n82509), .Z(n76853) );
  IV U96947 ( .A(n76853), .Z(n76854) );
  NOR U96948 ( .A(n82507), .B(n76854), .Z(n78789) );
  IV U96949 ( .A(n76855), .Z(n76857) );
  NOR U96950 ( .A(n76857), .B(n76856), .Z(n82511) );
  IV U96951 ( .A(n76858), .Z(n76859) );
  NOR U96952 ( .A(n76859), .B(n78784), .Z(n82518) );
  IV U96953 ( .A(n76860), .Z(n76865) );
  IV U96954 ( .A(n76861), .Z(n76862) );
  NOR U96955 ( .A(n76862), .B(n78784), .Z(n76863) );
  IV U96956 ( .A(n76863), .Z(n76864) );
  NOR U96957 ( .A(n76865), .B(n76864), .Z(n82515) );
  IV U96958 ( .A(n76866), .Z(n76867) );
  NOR U96959 ( .A(n76867), .B(n76869), .Z(n82532) );
  IV U96960 ( .A(n82532), .Z(n82530) );
  IV U96961 ( .A(n76868), .Z(n76870) );
  NOR U96962 ( .A(n76870), .B(n76869), .Z(n84507) );
  IV U96963 ( .A(n76871), .Z(n76872) );
  NOR U96964 ( .A(n76872), .B(n78767), .Z(n82543) );
  IV U96965 ( .A(n76873), .Z(n76874) );
  NOR U96966 ( .A(n76875), .B(n76874), .Z(n84510) );
  NOR U96967 ( .A(n82543), .B(n84510), .Z(n78774) );
  IV U96968 ( .A(n76876), .Z(n76878) );
  NOR U96969 ( .A(n76878), .B(n76877), .Z(n82538) );
  IV U96970 ( .A(n76879), .Z(n78771) );
  IV U96971 ( .A(n76880), .Z(n76881) );
  NOR U96972 ( .A(n78771), .B(n76881), .Z(n82548) );
  IV U96973 ( .A(n76882), .Z(n76883) );
  NOR U96974 ( .A(n76883), .B(n76885), .Z(n82552) );
  NOR U96975 ( .A(n82548), .B(n82552), .Z(n78765) );
  IV U96976 ( .A(n76884), .Z(n76886) );
  NOR U96977 ( .A(n76886), .B(n76885), .Z(n78763) );
  IV U96978 ( .A(n78763), .Z(n78749) );
  IV U96979 ( .A(n76887), .Z(n76888) );
  NOR U96980 ( .A(n76889), .B(n76888), .Z(n78731) );
  IV U96981 ( .A(n78731), .Z(n78726) );
  IV U96982 ( .A(n76890), .Z(n76891) );
  NOR U96983 ( .A(n76892), .B(n76891), .Z(n82563) );
  IV U96984 ( .A(n76893), .Z(n76896) );
  IV U96985 ( .A(n76894), .Z(n76895) );
  NOR U96986 ( .A(n76896), .B(n76895), .Z(n82569) );
  IV U96987 ( .A(n76897), .Z(n76900) );
  IV U96988 ( .A(n76898), .Z(n76899) );
  NOR U96989 ( .A(n76900), .B(n76899), .Z(n82566) );
  IV U96990 ( .A(n76901), .Z(n78719) );
  IV U96991 ( .A(n76902), .Z(n76904) );
  IV U96992 ( .A(n76903), .Z(n76906) );
  NOR U96993 ( .A(n76904), .B(n76906), .Z(n82577) );
  IV U96994 ( .A(n76905), .Z(n76907) );
  NOR U96995 ( .A(n76907), .B(n76906), .Z(n82588) );
  IV U96996 ( .A(n76908), .Z(n76910) );
  NOR U96997 ( .A(n76910), .B(n76909), .Z(n82585) );
  IV U96998 ( .A(n76911), .Z(n76912) );
  NOR U96999 ( .A(n76913), .B(n76912), .Z(n76914) );
  IV U97000 ( .A(n76914), .Z(n84493) );
  IV U97001 ( .A(n76915), .Z(n76916) );
  NOR U97002 ( .A(n76916), .B(n78708), .Z(n82601) );
  IV U97003 ( .A(n76917), .Z(n76918) );
  NOR U97004 ( .A(n76919), .B(n76918), .Z(n82599) );
  IV U97005 ( .A(n76920), .Z(n76923) );
  NOR U97006 ( .A(n76921), .B(n76928), .Z(n76922) );
  IV U97007 ( .A(n76922), .Z(n76925) );
  NOR U97008 ( .A(n76923), .B(n76925), .Z(n84476) );
  NOR U97009 ( .A(n82599), .B(n84476), .Z(n78705) );
  IV U97010 ( .A(n76924), .Z(n76926) );
  NOR U97011 ( .A(n76926), .B(n76925), .Z(n84479) );
  IV U97012 ( .A(n76927), .Z(n76931) );
  NOR U97013 ( .A(n76929), .B(n76928), .Z(n76930) );
  IV U97014 ( .A(n76930), .Z(n76933) );
  NOR U97015 ( .A(n76931), .B(n76933), .Z(n82609) );
  IV U97016 ( .A(n76932), .Z(n76934) );
  NOR U97017 ( .A(n76934), .B(n76933), .Z(n82606) );
  IV U97018 ( .A(n76935), .Z(n76936) );
  NOR U97019 ( .A(n76936), .B(n76941), .Z(n78700) );
  IV U97020 ( .A(n76937), .Z(n78692) );
  IV U97021 ( .A(n76938), .Z(n76939) );
  NOR U97022 ( .A(n78692), .B(n76939), .Z(n82638) );
  IV U97023 ( .A(n76940), .Z(n76942) );
  NOR U97024 ( .A(n76942), .B(n76941), .Z(n84472) );
  NOR U97025 ( .A(n82638), .B(n84472), .Z(n78698) );
  IV U97026 ( .A(n76943), .Z(n76947) );
  NOR U97027 ( .A(n76945), .B(n76944), .Z(n76946) );
  IV U97028 ( .A(n76946), .Z(n78676) );
  NOR U97029 ( .A(n76947), .B(n78676), .Z(n82652) );
  IV U97030 ( .A(n82652), .Z(n82650) );
  NOR U97031 ( .A(n76949), .B(n76948), .Z(n76951) );
  NOR U97032 ( .A(n76951), .B(n76950), .Z(n76952) );
  IV U97033 ( .A(n76952), .Z(n82665) );
  IV U97034 ( .A(n76953), .Z(n78667) );
  IV U97035 ( .A(n76954), .Z(n76955) );
  NOR U97036 ( .A(n78667), .B(n76955), .Z(n82661) );
  IV U97037 ( .A(n76956), .Z(n76958) );
  IV U97038 ( .A(n76957), .Z(n78669) );
  NOR U97039 ( .A(n76958), .B(n78669), .Z(n84456) );
  IV U97040 ( .A(n76959), .Z(n76960) );
  NOR U97041 ( .A(n76960), .B(n76963), .Z(n82669) );
  NOR U97042 ( .A(n76961), .B(n78669), .Z(n84448) );
  NOR U97043 ( .A(n82669), .B(n84448), .Z(n78664) );
  IV U97044 ( .A(n76962), .Z(n76964) );
  NOR U97045 ( .A(n76964), .B(n76963), .Z(n82666) );
  IV U97046 ( .A(n76965), .Z(n76970) );
  IV U97047 ( .A(n76966), .Z(n76967) );
  NOR U97048 ( .A(n76970), .B(n76967), .Z(n82671) );
  IV U97049 ( .A(n76968), .Z(n76969) );
  NOR U97050 ( .A(n76970), .B(n76969), .Z(n84441) );
  IV U97051 ( .A(n76971), .Z(n76973) );
  NOR U97052 ( .A(n76973), .B(n76972), .Z(n84438) );
  NOR U97053 ( .A(n76975), .B(n76974), .Z(n76977) );
  NOR U97054 ( .A(n76977), .B(n76976), .Z(n82675) );
  IV U97055 ( .A(n76978), .Z(n76983) );
  IV U97056 ( .A(n76979), .Z(n76980) );
  NOR U97057 ( .A(n76983), .B(n76980), .Z(n84434) );
  IV U97058 ( .A(n76981), .Z(n76982) );
  NOR U97059 ( .A(n76983), .B(n76982), .Z(n84431) );
  IV U97060 ( .A(n76984), .Z(n76985) );
  NOR U97061 ( .A(n76985), .B(n82688), .Z(n82678) );
  NOR U97062 ( .A(n76986), .B(n82688), .Z(n84421) );
  IV U97063 ( .A(n76987), .Z(n76989) );
  IV U97064 ( .A(n76988), .Z(n76992) );
  NOR U97065 ( .A(n76989), .B(n76992), .Z(n82685) );
  IV U97066 ( .A(n76990), .Z(n76991) );
  NOR U97067 ( .A(n76992), .B(n76991), .Z(n76993) );
  IV U97068 ( .A(n76993), .Z(n82698) );
  IV U97069 ( .A(n76994), .Z(n76995) );
  NOR U97070 ( .A(n76995), .B(n76997), .Z(n82694) );
  IV U97071 ( .A(n76996), .Z(n76998) );
  NOR U97072 ( .A(n76998), .B(n76997), .Z(n82703) );
  IV U97073 ( .A(n76999), .Z(n77000) );
  NOR U97074 ( .A(n77001), .B(n77000), .Z(n82708) );
  IV U97075 ( .A(n77002), .Z(n77004) );
  NOR U97076 ( .A(n77004), .B(n77003), .Z(n82701) );
  NOR U97077 ( .A(n82708), .B(n82701), .Z(n77005) );
  IV U97078 ( .A(n77005), .Z(n78663) );
  IV U97079 ( .A(n77006), .Z(n77014) );
  IV U97080 ( .A(n77007), .Z(n77008) );
  NOR U97081 ( .A(n77014), .B(n77008), .Z(n84416) );
  IV U97082 ( .A(n77009), .Z(n77010) );
  NOR U97083 ( .A(n77011), .B(n77010), .Z(n82712) );
  NOR U97084 ( .A(n84416), .B(n82712), .Z(n78662) );
  IV U97085 ( .A(n77012), .Z(n77013) );
  NOR U97086 ( .A(n77014), .B(n77013), .Z(n77015) );
  IV U97087 ( .A(n77015), .Z(n82711) );
  IV U97088 ( .A(n77019), .Z(n77016) );
  NOR U97089 ( .A(n77017), .B(n77016), .Z(n77024) );
  IV U97090 ( .A(n77017), .Z(n77018) );
  NOR U97091 ( .A(n77019), .B(n77018), .Z(n77022) );
  IV U97092 ( .A(n77020), .Z(n77021) );
  NOR U97093 ( .A(n77022), .B(n77021), .Z(n77023) );
  NOR U97094 ( .A(n77024), .B(n77023), .Z(n82719) );
  IV U97095 ( .A(n77025), .Z(n77032) );
  IV U97096 ( .A(n77026), .Z(n77027) );
  NOR U97097 ( .A(n77032), .B(n77027), .Z(n82715) );
  IV U97098 ( .A(n77028), .Z(n77029) );
  NOR U97099 ( .A(n77035), .B(n77029), .Z(n84409) );
  IV U97100 ( .A(n77030), .Z(n77031) );
  NOR U97101 ( .A(n77032), .B(n77031), .Z(n82722) );
  NOR U97102 ( .A(n84409), .B(n82722), .Z(n78659) );
  IV U97103 ( .A(n77033), .Z(n77034) );
  NOR U97104 ( .A(n77035), .B(n77034), .Z(n84412) );
  IV U97105 ( .A(n77036), .Z(n77038) );
  IV U97106 ( .A(n77037), .Z(n77041) );
  NOR U97107 ( .A(n77038), .B(n77041), .Z(n84402) );
  NOR U97108 ( .A(n84412), .B(n84402), .Z(n77045) );
  NOR U97109 ( .A(n77039), .B(n82725), .Z(n77043) );
  IV U97110 ( .A(n77040), .Z(n77042) );
  NOR U97111 ( .A(n77042), .B(n77041), .Z(n84398) );
  NOR U97112 ( .A(n77043), .B(n84398), .Z(n77044) );
  XOR U97113 ( .A(n77045), .B(n77044), .Z(n78658) );
  IV U97114 ( .A(n77046), .Z(n77051) );
  IV U97115 ( .A(n77047), .Z(n77048) );
  NOR U97116 ( .A(n77051), .B(n77048), .Z(n84382) );
  IV U97117 ( .A(n77049), .Z(n77050) );
  NOR U97118 ( .A(n77051), .B(n77050), .Z(n84385) );
  IV U97119 ( .A(n77052), .Z(n77054) );
  NOR U97120 ( .A(n77054), .B(n77053), .Z(n82731) );
  NOR U97121 ( .A(n77055), .B(n77056), .Z(n77062) );
  IV U97122 ( .A(n77056), .Z(n77058) );
  NOR U97123 ( .A(n77058), .B(n77057), .Z(n77060) );
  NOR U97124 ( .A(n77060), .B(n77059), .Z(n77061) );
  NOR U97125 ( .A(n77062), .B(n77061), .Z(n82734) );
  IV U97126 ( .A(n77063), .Z(n77065) );
  NOR U97127 ( .A(n77065), .B(n77064), .Z(n84368) );
  IV U97128 ( .A(n77066), .Z(n77067) );
  NOR U97129 ( .A(n77070), .B(n77067), .Z(n82740) );
  IV U97130 ( .A(n77068), .Z(n77069) );
  NOR U97131 ( .A(n77070), .B(n77069), .Z(n88468) );
  IV U97132 ( .A(n77071), .Z(n77072) );
  NOR U97133 ( .A(n77072), .B(n77077), .Z(n88506) );
  NOR U97134 ( .A(n88468), .B(n88506), .Z(n82739) );
  IV U97135 ( .A(n77073), .Z(n77074) );
  NOR U97136 ( .A(n77075), .B(n77074), .Z(n82746) );
  IV U97137 ( .A(n77076), .Z(n77078) );
  NOR U97138 ( .A(n77078), .B(n77077), .Z(n82743) );
  NOR U97139 ( .A(n82746), .B(n82743), .Z(n78657) );
  IV U97140 ( .A(n77079), .Z(n77080) );
  NOR U97141 ( .A(n78654), .B(n77080), .Z(n84355) );
  IV U97142 ( .A(n77081), .Z(n77083) );
  NOR U97143 ( .A(n77083), .B(n77082), .Z(n78636) );
  IV U97144 ( .A(n78636), .Z(n78631) );
  IV U97145 ( .A(n77084), .Z(n77085) );
  NOR U97146 ( .A(n77086), .B(n77085), .Z(n77087) );
  IV U97147 ( .A(n77087), .Z(n78615) );
  IV U97148 ( .A(n77088), .Z(n77090) );
  IV U97149 ( .A(n77089), .Z(n78613) );
  NOR U97150 ( .A(n77090), .B(n78613), .Z(n84330) );
  NOR U97151 ( .A(n77092), .B(n77091), .Z(n82771) );
  IV U97152 ( .A(n77093), .Z(n77096) );
  IV U97153 ( .A(n77094), .Z(n77095) );
  NOR U97154 ( .A(n77096), .B(n77095), .Z(n82773) );
  NOR U97155 ( .A(n82771), .B(n82773), .Z(n78608) );
  IV U97156 ( .A(n77097), .Z(n77100) );
  NOR U97157 ( .A(n77100), .B(n77104), .Z(n82787) );
  IV U97158 ( .A(n77098), .Z(n77102) );
  XOR U97159 ( .A(n77100), .B(n77099), .Z(n77101) );
  NOR U97160 ( .A(n77102), .B(n77101), .Z(n82776) );
  NOR U97161 ( .A(n82787), .B(n82776), .Z(n78607) );
  IV U97162 ( .A(n77103), .Z(n77105) );
  NOR U97163 ( .A(n77105), .B(n77104), .Z(n82779) );
  IV U97164 ( .A(n77106), .Z(n77107) );
  NOR U97165 ( .A(n77110), .B(n77107), .Z(n82782) );
  IV U97166 ( .A(n82782), .Z(n82785) );
  IV U97167 ( .A(n77108), .Z(n77109) );
  NOR U97168 ( .A(n77110), .B(n77109), .Z(n77111) );
  IV U97169 ( .A(n77111), .Z(n82791) );
  IV U97170 ( .A(n77112), .Z(n77115) );
  IV U97171 ( .A(n77113), .Z(n77114) );
  NOR U97172 ( .A(n77115), .B(n77114), .Z(n82795) );
  IV U97173 ( .A(n77116), .Z(n77118) );
  XOR U97174 ( .A(n77125), .B(n77126), .Z(n77117) );
  NOR U97175 ( .A(n77118), .B(n77117), .Z(n82792) );
  IV U97176 ( .A(n77119), .Z(n77120) );
  NOR U97177 ( .A(n77120), .B(n77126), .Z(n77121) );
  IV U97178 ( .A(n77121), .Z(n82802) );
  IV U97179 ( .A(n77122), .Z(n77124) );
  NOR U97180 ( .A(n77124), .B(n77123), .Z(n82807) );
  IV U97181 ( .A(n77125), .Z(n77127) );
  NOR U97182 ( .A(n77127), .B(n77126), .Z(n82803) );
  NOR U97183 ( .A(n82807), .B(n82803), .Z(n78606) );
  IV U97184 ( .A(n77128), .Z(n77129) );
  NOR U97185 ( .A(n77130), .B(n77129), .Z(n82814) );
  IV U97186 ( .A(n77131), .Z(n77133) );
  NOR U97187 ( .A(n77133), .B(n77132), .Z(n82810) );
  NOR U97188 ( .A(n82814), .B(n82810), .Z(n78605) );
  IV U97189 ( .A(n77134), .Z(n77138) );
  IV U97190 ( .A(n77135), .Z(n78590) );
  NOR U97191 ( .A(n77136), .B(n78590), .Z(n77137) );
  IV U97192 ( .A(n77137), .Z(n78596) );
  NOR U97193 ( .A(n77138), .B(n78596), .Z(n82822) );
  IV U97194 ( .A(n77139), .Z(n77140) );
  NOR U97195 ( .A(n77140), .B(n78590), .Z(n77141) );
  IV U97196 ( .A(n77141), .Z(n77142) );
  NOR U97197 ( .A(n77143), .B(n77142), .Z(n82833) );
  NOR U97198 ( .A(n77145), .B(n77144), .Z(n82836) );
  IV U97199 ( .A(n77146), .Z(n77147) );
  NOR U97200 ( .A(n78577), .B(n77147), .Z(n82841) );
  NOR U97201 ( .A(n82841), .B(n82839), .Z(n77148) );
  IV U97202 ( .A(n77148), .Z(n78588) );
  IV U97203 ( .A(n77149), .Z(n77150) );
  NOR U97204 ( .A(n78577), .B(n77150), .Z(n84322) );
  IV U97205 ( .A(n77151), .Z(n77152) );
  NOR U97206 ( .A(n77153), .B(n77152), .Z(n77156) );
  NOR U97207 ( .A(n77154), .B(n78581), .Z(n77155) );
  NOR U97208 ( .A(n77156), .B(n77155), .Z(n82845) );
  IV U97209 ( .A(n82845), .Z(n78572) );
  IV U97210 ( .A(n77157), .Z(n77160) );
  IV U97211 ( .A(n77158), .Z(n77159) );
  NOR U97212 ( .A(n77160), .B(n77159), .Z(n84310) );
  IV U97213 ( .A(n77161), .Z(n77164) );
  IV U97214 ( .A(n77162), .Z(n77163) );
  NOR U97215 ( .A(n77164), .B(n77163), .Z(n84307) );
  IV U97216 ( .A(n77165), .Z(n77167) );
  NOR U97217 ( .A(n77167), .B(n77166), .Z(n82870) );
  IV U97218 ( .A(n77168), .Z(n77170) );
  NOR U97219 ( .A(n77170), .B(n77169), .Z(n82866) );
  NOR U97220 ( .A(n82870), .B(n82866), .Z(n78555) );
  IV U97221 ( .A(n77171), .Z(n77175) );
  XOR U97222 ( .A(n77188), .B(n77189), .Z(n77172) );
  NOR U97223 ( .A(n77173), .B(n77172), .Z(n77174) );
  IV U97224 ( .A(n77174), .Z(n77178) );
  NOR U97225 ( .A(n77175), .B(n77178), .Z(n77176) );
  IV U97226 ( .A(n77176), .Z(n82875) );
  IV U97227 ( .A(n77177), .Z(n77179) );
  NOR U97228 ( .A(n77179), .B(n77178), .Z(n77180) );
  IV U97229 ( .A(n77180), .Z(n82881) );
  IV U97230 ( .A(n77181), .Z(n77182) );
  NOR U97231 ( .A(n77182), .B(n77189), .Z(n77187) );
  IV U97232 ( .A(n77183), .Z(n77185) );
  NOR U97233 ( .A(n77185), .B(n77184), .Z(n77186) );
  NOR U97234 ( .A(n77187), .B(n77186), .Z(n82878) );
  IV U97235 ( .A(n77188), .Z(n77190) );
  NOR U97236 ( .A(n77190), .B(n77189), .Z(n82886) );
  NOR U97237 ( .A(n77192), .B(n77191), .Z(n82894) );
  IV U97238 ( .A(n77193), .Z(n77194) );
  NOR U97239 ( .A(n77195), .B(n77194), .Z(n84270) );
  IV U97240 ( .A(n77196), .Z(n77198) );
  IV U97241 ( .A(n77197), .Z(n78487) );
  NOR U97242 ( .A(n77198), .B(n78487), .Z(n77202) );
  IV U97243 ( .A(n77199), .Z(n77200) );
  NOR U97244 ( .A(n77200), .B(n78492), .Z(n77201) );
  NOR U97245 ( .A(n77202), .B(n77201), .Z(n84251) );
  IV U97246 ( .A(n77203), .Z(n77204) );
  NOR U97247 ( .A(n78484), .B(n77204), .Z(n84245) );
  IV U97248 ( .A(n77205), .Z(n77206) );
  NOR U97249 ( .A(n77206), .B(n77211), .Z(n82917) );
  IV U97250 ( .A(n77207), .Z(n77208) );
  NOR U97251 ( .A(n77209), .B(n77208), .Z(n82913) );
  NOR U97252 ( .A(n82917), .B(n82913), .Z(n78482) );
  IV U97253 ( .A(n77210), .Z(n77212) );
  NOR U97254 ( .A(n77212), .B(n77211), .Z(n78480) );
  IV U97255 ( .A(n78480), .Z(n78471) );
  IV U97256 ( .A(n77213), .Z(n77215) );
  NOR U97257 ( .A(n77215), .B(n77214), .Z(n77216) );
  IV U97258 ( .A(n77216), .Z(n82925) );
  IV U97259 ( .A(n77217), .Z(n77218) );
  NOR U97260 ( .A(n77218), .B(n77223), .Z(n82921) );
  IV U97261 ( .A(n77219), .Z(n77220) );
  NOR U97262 ( .A(n77221), .B(n77220), .Z(n82930) );
  IV U97263 ( .A(n77222), .Z(n77224) );
  NOR U97264 ( .A(n77224), .B(n77223), .Z(n82927) );
  NOR U97265 ( .A(n82930), .B(n82927), .Z(n78470) );
  NOR U97266 ( .A(n77225), .B(n82935), .Z(n77229) );
  IV U97267 ( .A(n77226), .Z(n77231) );
  IV U97268 ( .A(n77227), .Z(n77228) );
  NOR U97269 ( .A(n77231), .B(n77228), .Z(n84228) );
  NOR U97270 ( .A(n77229), .B(n84228), .Z(n78469) );
  IV U97271 ( .A(n77230), .Z(n77232) );
  NOR U97272 ( .A(n77232), .B(n77231), .Z(n82941) );
  IV U97273 ( .A(n77233), .Z(n77235) );
  NOR U97274 ( .A(n77235), .B(n77234), .Z(n82938) );
  IV U97275 ( .A(n77236), .Z(n77238) );
  NOR U97276 ( .A(n77238), .B(n77237), .Z(n84209) );
  IV U97277 ( .A(n77239), .Z(n77241) );
  NOR U97278 ( .A(n77241), .B(n77240), .Z(n84218) );
  NOR U97279 ( .A(n84209), .B(n84218), .Z(n77242) );
  IV U97280 ( .A(n77242), .Z(n78468) );
  IV U97281 ( .A(n77243), .Z(n77244) );
  NOR U97282 ( .A(n77244), .B(n77246), .Z(n84192) );
  IV U97283 ( .A(n77245), .Z(n77247) );
  NOR U97284 ( .A(n77247), .B(n77246), .Z(n82961) );
  IV U97285 ( .A(n77248), .Z(n77251) );
  IV U97286 ( .A(n77249), .Z(n77250) );
  NOR U97287 ( .A(n77251), .B(n77250), .Z(n78424) );
  XOR U97288 ( .A(n77252), .B(n78414), .Z(n77255) );
  IV U97289 ( .A(n77253), .Z(n77254) );
  NOR U97290 ( .A(n77255), .B(n77254), .Z(n78421) );
  IV U97291 ( .A(n78421), .Z(n78412) );
  IV U97292 ( .A(n77256), .Z(n77258) );
  NOR U97293 ( .A(n77258), .B(n77257), .Z(n82972) );
  IV U97294 ( .A(n77259), .Z(n77261) );
  NOR U97295 ( .A(n77261), .B(n77260), .Z(n78371) );
  IV U97296 ( .A(n78371), .Z(n78362) );
  IV U97297 ( .A(n77262), .Z(n77264) );
  NOR U97298 ( .A(n77264), .B(n77263), .Z(n82993) );
  IV U97299 ( .A(n77265), .Z(n77266) );
  NOR U97300 ( .A(n77266), .B(n78352), .Z(n82991) );
  NOR U97301 ( .A(n82993), .B(n82991), .Z(n78349) );
  IV U97302 ( .A(n77267), .Z(n77268) );
  NOR U97303 ( .A(n77268), .B(n78345), .Z(n84154) );
  IV U97304 ( .A(n77269), .Z(n77271) );
  NOR U97305 ( .A(n77271), .B(n77270), .Z(n83002) );
  NOR U97306 ( .A(n77273), .B(n77272), .Z(n78334) );
  IV U97307 ( .A(n78334), .Z(n78326) );
  IV U97308 ( .A(n77274), .Z(n77275) );
  NOR U97309 ( .A(n78330), .B(n77275), .Z(n83015) );
  IV U97310 ( .A(n77276), .Z(n83026) );
  NOR U97311 ( .A(n77277), .B(n83026), .Z(n83017) );
  IV U97312 ( .A(n77278), .Z(n77279) );
  NOR U97313 ( .A(n77282), .B(n77279), .Z(n83035) );
  IV U97314 ( .A(n77280), .Z(n77281) );
  NOR U97315 ( .A(n77282), .B(n77281), .Z(n83032) );
  XOR U97316 ( .A(n83035), .B(n83032), .Z(n77283) );
  NOR U97317 ( .A(n83017), .B(n77283), .Z(n78324) );
  IV U97318 ( .A(n77284), .Z(n77287) );
  IV U97319 ( .A(n77285), .Z(n77286) );
  NOR U97320 ( .A(n77287), .B(n77286), .Z(n83051) );
  IV U97321 ( .A(n77288), .Z(n77290) );
  NOR U97322 ( .A(n77290), .B(n77289), .Z(n83046) );
  IV U97323 ( .A(n77291), .Z(n77292) );
  NOR U97324 ( .A(n77292), .B(n77297), .Z(n83043) );
  IV U97325 ( .A(n77293), .Z(n77295) );
  NOR U97326 ( .A(n77295), .B(n77294), .Z(n83057) );
  IV U97327 ( .A(n77296), .Z(n77298) );
  NOR U97328 ( .A(n77298), .B(n77297), .Z(n83055) );
  NOR U97329 ( .A(n83057), .B(n83055), .Z(n77299) );
  IV U97330 ( .A(n77299), .Z(n78323) );
  IV U97331 ( .A(n77300), .Z(n77301) );
  NOR U97332 ( .A(n77302), .B(n77301), .Z(n83067) );
  IV U97333 ( .A(n77303), .Z(n77304) );
  NOR U97334 ( .A(n77305), .B(n77304), .Z(n83060) );
  NOR U97335 ( .A(n83067), .B(n83060), .Z(n78322) );
  IV U97336 ( .A(n77306), .Z(n77307) );
  NOR U97337 ( .A(n78316), .B(n77307), .Z(n83070) );
  IV U97338 ( .A(n77308), .Z(n78302) );
  IV U97339 ( .A(n77311), .Z(n77309) );
  NOR U97340 ( .A(n78302), .B(n77309), .Z(n83088) );
  IV U97341 ( .A(n77310), .Z(n77313) );
  XOR U97342 ( .A(n77311), .B(n78302), .Z(n77312) );
  NOR U97343 ( .A(n77313), .B(n77312), .Z(n84113) );
  NOR U97344 ( .A(n83088), .B(n84113), .Z(n78299) );
  IV U97345 ( .A(n77314), .Z(n77315) );
  NOR U97346 ( .A(n78263), .B(n77315), .Z(n78269) );
  IV U97347 ( .A(n78269), .Z(n78260) );
  IV U97348 ( .A(n77316), .Z(n77317) );
  NOR U97349 ( .A(n77318), .B(n77317), .Z(n83107) );
  IV U97350 ( .A(n77319), .Z(n77320) );
  NOR U97351 ( .A(n77321), .B(n77320), .Z(n83105) );
  NOR U97352 ( .A(n83107), .B(n83105), .Z(n78258) );
  IV U97353 ( .A(n77322), .Z(n77323) );
  NOR U97354 ( .A(n77324), .B(n77323), .Z(n84094) );
  IV U97355 ( .A(n77325), .Z(n77326) );
  NOR U97356 ( .A(n77326), .B(n78251), .Z(n84087) );
  NOR U97357 ( .A(n84094), .B(n84087), .Z(n78257) );
  IV U97358 ( .A(n77327), .Z(n78245) );
  NOR U97359 ( .A(n78245), .B(n77328), .Z(n77329) );
  NOR U97360 ( .A(n77330), .B(n77329), .Z(n84080) );
  IV U97361 ( .A(n77331), .Z(n77333) );
  NOR U97362 ( .A(n77333), .B(n77332), .Z(n84065) );
  IV U97363 ( .A(n77334), .Z(n77335) );
  NOR U97364 ( .A(n77336), .B(n77335), .Z(n84062) );
  NOR U97365 ( .A(n84065), .B(n84062), .Z(n78242) );
  IV U97366 ( .A(n77337), .Z(n77338) );
  NOR U97367 ( .A(n77339), .B(n77338), .Z(n83114) );
  IV U97368 ( .A(n77340), .Z(n77341) );
  NOR U97369 ( .A(n77342), .B(n77341), .Z(n84068) );
  NOR U97370 ( .A(n83114), .B(n84068), .Z(n78241) );
  IV U97371 ( .A(n77343), .Z(n77345) );
  IV U97372 ( .A(n77344), .Z(n78232) );
  NOR U97373 ( .A(n77345), .B(n78232), .Z(n78239) );
  IV U97374 ( .A(n78239), .Z(n78230) );
  IV U97375 ( .A(n77346), .Z(n77347) );
  NOR U97376 ( .A(n77347), .B(n77349), .Z(n83119) );
  IV U97377 ( .A(n77348), .Z(n77350) );
  NOR U97378 ( .A(n77350), .B(n77349), .Z(n83121) );
  NOR U97379 ( .A(n83119), .B(n83121), .Z(n78228) );
  IV U97380 ( .A(n77351), .Z(n77353) );
  NOR U97381 ( .A(n77353), .B(n77352), .Z(n83124) );
  NOR U97382 ( .A(n84051), .B(n83124), .Z(n78226) );
  IV U97383 ( .A(n77354), .Z(n77355) );
  NOR U97384 ( .A(n77358), .B(n77355), .Z(n84046) );
  IV U97385 ( .A(n84046), .Z(n84049) );
  IV U97386 ( .A(n77356), .Z(n77357) );
  NOR U97387 ( .A(n77358), .B(n77357), .Z(n77359) );
  IV U97388 ( .A(n77359), .Z(n83130) );
  IV U97389 ( .A(n77360), .Z(n77362) );
  NOR U97390 ( .A(n77362), .B(n77361), .Z(n84036) );
  IV U97391 ( .A(n77363), .Z(n77364) );
  NOR U97392 ( .A(n78218), .B(n77364), .Z(n84033) );
  IV U97393 ( .A(n77365), .Z(n77367) );
  NOR U97394 ( .A(n77367), .B(n77366), .Z(n77368) );
  IV U97395 ( .A(n77368), .Z(n84027) );
  IV U97396 ( .A(n77369), .Z(n77375) );
  IV U97397 ( .A(n77370), .Z(n77372) );
  NOR U97398 ( .A(n77372), .B(n77371), .Z(n77373) );
  IV U97399 ( .A(n77373), .Z(n77374) );
  NOR U97400 ( .A(n77375), .B(n77374), .Z(n84014) );
  IV U97401 ( .A(n77376), .Z(n77377) );
  NOR U97402 ( .A(n77377), .B(n77384), .Z(n77378) );
  IV U97403 ( .A(n77378), .Z(n77379) );
  NOR U97404 ( .A(n77380), .B(n77379), .Z(n83139) );
  NOR U97405 ( .A(n77381), .B(n83998), .Z(n77385) );
  IV U97406 ( .A(n77382), .Z(n77383) );
  NOR U97407 ( .A(n77384), .B(n77383), .Z(n84007) );
  NOR U97408 ( .A(n77385), .B(n84007), .Z(n78205) );
  IV U97409 ( .A(n77386), .Z(n77387) );
  NOR U97410 ( .A(n77388), .B(n77387), .Z(n77393) );
  IV U97411 ( .A(n77389), .Z(n77391) );
  NOR U97412 ( .A(n77391), .B(n77390), .Z(n77392) );
  NOR U97413 ( .A(n77393), .B(n77392), .Z(n84003) );
  IV U97414 ( .A(n77394), .Z(n77396) );
  NOR U97415 ( .A(n77396), .B(n77395), .Z(n77397) );
  IV U97416 ( .A(n77397), .Z(n83990) );
  IV U97417 ( .A(n77398), .Z(n77400) );
  NOR U97418 ( .A(n77400), .B(n77399), .Z(n83992) );
  IV U97419 ( .A(n77401), .Z(n77403) );
  NOR U97420 ( .A(n77403), .B(n77402), .Z(n83143) );
  NOR U97421 ( .A(n83143), .B(n83975), .Z(n77404) );
  IV U97422 ( .A(n77404), .Z(n77405) );
  NOR U97423 ( .A(n83992), .B(n77405), .Z(n78204) );
  IV U97424 ( .A(n77406), .Z(n77408) );
  NOR U97425 ( .A(n77408), .B(n77407), .Z(n83145) );
  IV U97426 ( .A(n77409), .Z(n77411) );
  NOR U97427 ( .A(n77411), .B(n77410), .Z(n83175) );
  IV U97428 ( .A(n77412), .Z(n77413) );
  NOR U97429 ( .A(n77414), .B(n77413), .Z(n83173) );
  NOR U97430 ( .A(n83175), .B(n83173), .Z(n78180) );
  IV U97431 ( .A(n77415), .Z(n77416) );
  NOR U97432 ( .A(n77416), .B(n78182), .Z(n83171) );
  NOR U97433 ( .A(n78161), .B(n77417), .Z(n77418) );
  IV U97434 ( .A(n77418), .Z(n78167) );
  NOR U97435 ( .A(n77419), .B(n78167), .Z(n77420) );
  IV U97436 ( .A(n77420), .Z(n77421) );
  NOR U97437 ( .A(n78166), .B(n77421), .Z(n77422) );
  IV U97438 ( .A(n77422), .Z(n83963) );
  IV U97439 ( .A(n77423), .Z(n77425) );
  IV U97440 ( .A(n77424), .Z(n78153) );
  NOR U97441 ( .A(n77425), .B(n78153), .Z(n78151) );
  IV U97442 ( .A(n78151), .Z(n78146) );
  XOR U97443 ( .A(n78142), .B(n78148), .Z(n77428) );
  IV U97444 ( .A(n77426), .Z(n77427) );
  NOR U97445 ( .A(n77428), .B(n77427), .Z(n83948) );
  IV U97446 ( .A(n77429), .Z(n77431) );
  IV U97447 ( .A(n77430), .Z(n78137) );
  NOR U97448 ( .A(n77431), .B(n78137), .Z(n83192) );
  IV U97449 ( .A(n77432), .Z(n77433) );
  NOR U97450 ( .A(n77433), .B(n77438), .Z(n83199) );
  IV U97451 ( .A(n77434), .Z(n77435) );
  NOR U97452 ( .A(n77436), .B(n77435), .Z(n83938) );
  IV U97453 ( .A(n77437), .Z(n77439) );
  NOR U97454 ( .A(n77439), .B(n77438), .Z(n83205) );
  NOR U97455 ( .A(n83938), .B(n83205), .Z(n78134) );
  NOR U97456 ( .A(n78117), .B(n77440), .Z(n83929) );
  IV U97457 ( .A(n77441), .Z(n77442) );
  NOR U97458 ( .A(n78109), .B(n77442), .Z(n78102) );
  IV U97459 ( .A(n77443), .Z(n77445) );
  NOR U97460 ( .A(n77445), .B(n77444), .Z(n78098) );
  IV U97461 ( .A(n77446), .Z(n77447) );
  NOR U97462 ( .A(n77447), .B(n78095), .Z(n83910) );
  NOR U97463 ( .A(n77448), .B(n83236), .Z(n77452) );
  IV U97464 ( .A(n77449), .Z(n77451) );
  NOR U97465 ( .A(n77451), .B(n77450), .Z(n83906) );
  NOR U97466 ( .A(n77452), .B(n83906), .Z(n78093) );
  IV U97467 ( .A(n77453), .Z(n77455) );
  IV U97468 ( .A(n77454), .Z(n78081) );
  NOR U97469 ( .A(n77455), .B(n78081), .Z(n78089) );
  NOR U97470 ( .A(n77456), .B(n83248), .Z(n78079) );
  IV U97471 ( .A(n77457), .Z(n77458) );
  NOR U97472 ( .A(n77461), .B(n77458), .Z(n83259) );
  IV U97473 ( .A(n77459), .Z(n77460) );
  NOR U97474 ( .A(n77461), .B(n77460), .Z(n83891) );
  NOR U97475 ( .A(n83259), .B(n83891), .Z(n77462) );
  IV U97476 ( .A(n77462), .Z(n77463) );
  NOR U97477 ( .A(n83257), .B(n77463), .Z(n77464) );
  IV U97478 ( .A(n77464), .Z(n78073) );
  NOR U97479 ( .A(n77465), .B(n83870), .Z(n77466) );
  IV U97480 ( .A(n77466), .Z(n83268) );
  IV U97481 ( .A(n77467), .Z(n77469) );
  NOR U97482 ( .A(n77469), .B(n77468), .Z(n83279) );
  IV U97483 ( .A(n77470), .Z(n77472) );
  NOR U97484 ( .A(n77472), .B(n77471), .Z(n83272) );
  NOR U97485 ( .A(n83279), .B(n83272), .Z(n78056) );
  IV U97486 ( .A(n77473), .Z(n77474) );
  NOR U97487 ( .A(n77474), .B(n77480), .Z(n83277) );
  IV U97488 ( .A(n83277), .Z(n83275) );
  IV U97489 ( .A(n77475), .Z(n77477) );
  IV U97490 ( .A(n77476), .Z(n77487) );
  NOR U97491 ( .A(n77477), .B(n77487), .Z(n89593) );
  IV U97492 ( .A(n77478), .Z(n77479) );
  NOR U97493 ( .A(n77480), .B(n77479), .Z(n89018) );
  NOR U97494 ( .A(n89593), .B(n89018), .Z(n83860) );
  IV U97495 ( .A(n77481), .Z(n77484) );
  IV U97496 ( .A(n77482), .Z(n77483) );
  NOR U97497 ( .A(n77484), .B(n77483), .Z(n83857) );
  IV U97498 ( .A(n77485), .Z(n77486) );
  NOR U97499 ( .A(n77487), .B(n77486), .Z(n89592) );
  NOR U97500 ( .A(n83857), .B(n89592), .Z(n78055) );
  IV U97501 ( .A(n77488), .Z(n77489) );
  NOR U97502 ( .A(n77490), .B(n77489), .Z(n83296) );
  IV U97503 ( .A(n77491), .Z(n77492) );
  NOR U97504 ( .A(n77492), .B(n77494), .Z(n83298) );
  NOR U97505 ( .A(n83296), .B(n83298), .Z(n78038) );
  IV U97506 ( .A(n77493), .Z(n77495) );
  NOR U97507 ( .A(n77495), .B(n77494), .Z(n83846) );
  IV U97508 ( .A(n77496), .Z(n77497) );
  NOR U97509 ( .A(n77504), .B(n77497), .Z(n83302) );
  IV U97510 ( .A(n77498), .Z(n77499) );
  NOR U97511 ( .A(n77500), .B(n77499), .Z(n83850) );
  NOR U97512 ( .A(n83302), .B(n83850), .Z(n78037) );
  IV U97513 ( .A(n77501), .Z(n83841) );
  NOR U97514 ( .A(n77502), .B(n83841), .Z(n77506) );
  IV U97515 ( .A(n77503), .Z(n77505) );
  NOR U97516 ( .A(n77505), .B(n77504), .Z(n83304) );
  NOR U97517 ( .A(n77506), .B(n83304), .Z(n78036) );
  IV U97518 ( .A(n77507), .Z(n77511) );
  NOR U97519 ( .A(n77509), .B(n77508), .Z(n77510) );
  IV U97520 ( .A(n77510), .Z(n77513) );
  NOR U97521 ( .A(n77511), .B(n77513), .Z(n83308) );
  IV U97522 ( .A(n83308), .Z(n83306) );
  IV U97523 ( .A(n77512), .Z(n77514) );
  NOR U97524 ( .A(n77514), .B(n77513), .Z(n77515) );
  IV U97525 ( .A(n77515), .Z(n83835) );
  NOR U97526 ( .A(n78018), .B(n77516), .Z(n77517) );
  IV U97527 ( .A(n77517), .Z(n77522) );
  NOR U97528 ( .A(n77519), .B(n77518), .Z(n77520) );
  IV U97529 ( .A(n77520), .Z(n77521) );
  NOR U97530 ( .A(n77522), .B(n77521), .Z(n78011) );
  IV U97531 ( .A(n77523), .Z(n77526) );
  NOR U97532 ( .A(n77997), .B(n77524), .Z(n77525) );
  IV U97533 ( .A(n77525), .Z(n77999) );
  NOR U97534 ( .A(n77526), .B(n77999), .Z(n77527) );
  IV U97535 ( .A(n77527), .Z(n83323) );
  IV U97536 ( .A(n77528), .Z(n77530) );
  NOR U97537 ( .A(n77530), .B(n77529), .Z(n77531) );
  IV U97538 ( .A(n77531), .Z(n83322) );
  IV U97539 ( .A(n77532), .Z(n77533) );
  NOR U97540 ( .A(n77992), .B(n77533), .Z(n77534) );
  IV U97541 ( .A(n77534), .Z(n77986) );
  IV U97542 ( .A(n77535), .Z(n77536) );
  NOR U97543 ( .A(n77537), .B(n77536), .Z(n83815) );
  IV U97544 ( .A(n77538), .Z(n77539) );
  NOR U97545 ( .A(n77540), .B(n77539), .Z(n77928) );
  IV U97546 ( .A(n77928), .Z(n77923) );
  IV U97547 ( .A(n77541), .Z(n77918) );
  IV U97548 ( .A(n77542), .Z(n77543) );
  NOR U97549 ( .A(n77918), .B(n77543), .Z(n83794) );
  IV U97550 ( .A(n77544), .Z(n77545) );
  NOR U97551 ( .A(n77546), .B(n77545), .Z(n83783) );
  IV U97552 ( .A(n77547), .Z(n77548) );
  NOR U97553 ( .A(n77548), .B(n77906), .Z(n83787) );
  NOR U97554 ( .A(n83783), .B(n83787), .Z(n77903) );
  IV U97555 ( .A(n77549), .Z(n77902) );
  IV U97556 ( .A(n77550), .Z(n77551) );
  NOR U97557 ( .A(n77902), .B(n77551), .Z(n83369) );
  IV U97558 ( .A(n77552), .Z(n77554) );
  NOR U97559 ( .A(n77554), .B(n77553), .Z(n83398) );
  IV U97560 ( .A(n77555), .Z(n77556) );
  NOR U97561 ( .A(n77559), .B(n77556), .Z(n83405) );
  IV U97562 ( .A(n77557), .Z(n77558) );
  NOR U97563 ( .A(n77559), .B(n77558), .Z(n83408) );
  IV U97564 ( .A(n77560), .Z(n77562) );
  IV U97565 ( .A(n77561), .Z(n77564) );
  NOR U97566 ( .A(n77562), .B(n77564), .Z(n83411) );
  NOR U97567 ( .A(n83408), .B(n83411), .Z(n77876) );
  IV U97568 ( .A(n77563), .Z(n77567) );
  NOR U97569 ( .A(n77565), .B(n77564), .Z(n77566) );
  IV U97570 ( .A(n77566), .Z(n77569) );
  NOR U97571 ( .A(n77567), .B(n77569), .Z(n83766) );
  IV U97572 ( .A(n77568), .Z(n77570) );
  NOR U97573 ( .A(n77570), .B(n77569), .Z(n83763) );
  IV U97574 ( .A(n77571), .Z(n77573) );
  NOR U97575 ( .A(n77573), .B(n77572), .Z(n83416) );
  IV U97576 ( .A(n77574), .Z(n77576) );
  NOR U97577 ( .A(n77576), .B(n77575), .Z(n83424) );
  IV U97578 ( .A(n77577), .Z(n77579) );
  NOR U97579 ( .A(n77579), .B(n77578), .Z(n83422) );
  NOR U97580 ( .A(n83424), .B(n83422), .Z(n77875) );
  IV U97581 ( .A(n77580), .Z(n77581) );
  NOR U97582 ( .A(n77872), .B(n77581), .Z(n83748) );
  IV U97583 ( .A(n77582), .Z(n77583) );
  NOR U97584 ( .A(n77859), .B(n77583), .Z(n83743) );
  IV U97585 ( .A(n77584), .Z(n77586) );
  IV U97586 ( .A(n77585), .Z(n77589) );
  NOR U97587 ( .A(n77586), .B(n77589), .Z(n77587) );
  IV U97588 ( .A(n77587), .Z(n83741) );
  IV U97589 ( .A(n77588), .Z(n77590) );
  NOR U97590 ( .A(n77590), .B(n77589), .Z(n83726) );
  NOR U97591 ( .A(n77591), .B(n83726), .Z(n77856) );
  IV U97592 ( .A(n77592), .Z(n77594) );
  NOR U97593 ( .A(n77594), .B(n77593), .Z(n83451) );
  IV U97594 ( .A(n83451), .Z(n83448) );
  IV U97595 ( .A(n77595), .Z(n77596) );
  NOR U97596 ( .A(n77599), .B(n77596), .Z(n83467) );
  IV U97597 ( .A(n77597), .Z(n77598) );
  NOR U97598 ( .A(n77599), .B(n77598), .Z(n83464) );
  IV U97599 ( .A(n77600), .Z(n77601) );
  NOR U97600 ( .A(n77604), .B(n77601), .Z(n83474) );
  IV U97601 ( .A(n77602), .Z(n77603) );
  NOR U97602 ( .A(n77604), .B(n77603), .Z(n83476) );
  IV U97603 ( .A(n77605), .Z(n77607) );
  NOR U97604 ( .A(n77607), .B(n77606), .Z(n83470) );
  NOR U97605 ( .A(n83476), .B(n83470), .Z(n77850) );
  IV U97606 ( .A(n77608), .Z(n77611) );
  IV U97607 ( .A(n77609), .Z(n77610) );
  NOR U97608 ( .A(n77611), .B(n77610), .Z(n77612) );
  IV U97609 ( .A(n77612), .Z(n83707) );
  IV U97610 ( .A(n77613), .Z(n77616) );
  IV U97611 ( .A(n77614), .Z(n77615) );
  NOR U97612 ( .A(n77616), .B(n77615), .Z(n83704) );
  IV U97613 ( .A(n77617), .Z(n77619) );
  NOR U97614 ( .A(n77619), .B(n77618), .Z(n77624) );
  IV U97615 ( .A(n77620), .Z(n77622) );
  NOR U97616 ( .A(n77622), .B(n77621), .Z(n77623) );
  NOR U97617 ( .A(n77624), .B(n77623), .Z(n83481) );
  IV U97618 ( .A(n83481), .Z(n77849) );
  IV U97619 ( .A(n77628), .Z(n77625) );
  NOR U97620 ( .A(n77625), .B(n77626), .Z(n83483) );
  IV U97621 ( .A(n77626), .Z(n77627) );
  NOR U97622 ( .A(n77628), .B(n77627), .Z(n77633) );
  XOR U97623 ( .A(n77630), .B(n77629), .Z(n77631) );
  IV U97624 ( .A(n77631), .Z(n77632) );
  NOR U97625 ( .A(n77633), .B(n77632), .Z(n77634) );
  NOR U97626 ( .A(n83483), .B(n77634), .Z(n77848) );
  IV U97627 ( .A(n77635), .Z(n77637) );
  NOR U97628 ( .A(n77637), .B(n77636), .Z(n77846) );
  IV U97629 ( .A(n77846), .Z(n77837) );
  IV U97630 ( .A(n77638), .Z(n77639) );
  NOR U97631 ( .A(n77639), .B(n77645), .Z(n77640) );
  IV U97632 ( .A(n77640), .Z(n83488) );
  IV U97633 ( .A(n77641), .Z(n77642) );
  NOR U97634 ( .A(n77643), .B(n77642), .Z(n83495) );
  IV U97635 ( .A(n77644), .Z(n77646) );
  NOR U97636 ( .A(n77646), .B(n77645), .Z(n83493) );
  NOR U97637 ( .A(n83495), .B(n83493), .Z(n77836) );
  IV U97638 ( .A(n77647), .Z(n77652) );
  IV U97639 ( .A(n77648), .Z(n77649) );
  NOR U97640 ( .A(n77652), .B(n77649), .Z(n83502) );
  IV U97641 ( .A(n77650), .Z(n77651) );
  NOR U97642 ( .A(n77652), .B(n77651), .Z(n83509) );
  NOR U97643 ( .A(n83502), .B(n83509), .Z(n77827) );
  IV U97644 ( .A(n77653), .Z(n77654) );
  NOR U97645 ( .A(n77654), .B(n77823), .Z(n83515) );
  IV U97646 ( .A(n77655), .Z(n77658) );
  NOR U97647 ( .A(n77656), .B(n77807), .Z(n77657) );
  IV U97648 ( .A(n77657), .Z(n77813) );
  NOR U97649 ( .A(n77658), .B(n77813), .Z(n83680) );
  IV U97650 ( .A(n77659), .Z(n77800) );
  IV U97651 ( .A(n77660), .Z(n77661) );
  NOR U97652 ( .A(n77800), .B(n77661), .Z(n83527) );
  IV U97653 ( .A(n77662), .Z(n77663) );
  NOR U97654 ( .A(n77663), .B(n77773), .Z(n77664) );
  IV U97655 ( .A(n77664), .Z(n77778) );
  IV U97656 ( .A(n77665), .Z(n77673) );
  IV U97657 ( .A(n77666), .Z(n77667) );
  NOR U97658 ( .A(n77673), .B(n77667), .Z(n83546) );
  IV U97659 ( .A(n77668), .Z(n77669) );
  NOR U97660 ( .A(n77670), .B(n77669), .Z(n83547) );
  NOR U97661 ( .A(n83546), .B(n83547), .Z(n77754) );
  IV U97662 ( .A(n77671), .Z(n77672) );
  NOR U97663 ( .A(n77673), .B(n77672), .Z(n83648) );
  IV U97664 ( .A(n77674), .Z(n77675) );
  NOR U97665 ( .A(n77675), .B(n77749), .Z(n83645) );
  NOR U97666 ( .A(n77676), .B(n83561), .Z(n77753) );
  IV U97667 ( .A(n77677), .Z(n77678) );
  NOR U97668 ( .A(n77678), .B(n77684), .Z(n77679) );
  IV U97669 ( .A(n77679), .Z(n83628) );
  IV U97670 ( .A(n77680), .Z(n77681) );
  NOR U97671 ( .A(n77682), .B(n77681), .Z(n83567) );
  IV U97672 ( .A(n77683), .Z(n77685) );
  NOR U97673 ( .A(n77685), .B(n77684), .Z(n83564) );
  NOR U97674 ( .A(n83567), .B(n83564), .Z(n77745) );
  IV U97675 ( .A(n77686), .Z(n77689) );
  IV U97676 ( .A(n77687), .Z(n77688) );
  NOR U97677 ( .A(n77689), .B(n77688), .Z(n83617) );
  IV U97678 ( .A(n77690), .Z(n77692) );
  XOR U97679 ( .A(n77739), .B(n77742), .Z(n77691) );
  NOR U97680 ( .A(n77692), .B(n77691), .Z(n83614) );
  IV U97681 ( .A(n77693), .Z(n77695) );
  IV U97682 ( .A(n77694), .Z(n77697) );
  NOR U97683 ( .A(n77695), .B(n77697), .Z(n83606) );
  IV U97684 ( .A(n77696), .Z(n77698) );
  NOR U97685 ( .A(n77698), .B(n77697), .Z(n83586) );
  NOR U97686 ( .A(n83581), .B(n83586), .Z(n77722) );
  IV U97687 ( .A(n77701), .Z(n77699) );
  NOR U97688 ( .A(n77700), .B(n77699), .Z(n77706) );
  NOR U97689 ( .A(n77702), .B(n77701), .Z(n77704) );
  NOR U97690 ( .A(n77704), .B(n77703), .Z(n77705) );
  NOR U97691 ( .A(n77706), .B(n77705), .Z(n83576) );
  IV U97692 ( .A(n77707), .Z(n77708) );
  NOR U97693 ( .A(n77709), .B(n77708), .Z(n77714) );
  IV U97694 ( .A(n77710), .Z(n77711) );
  NOR U97695 ( .A(n77712), .B(n77711), .Z(n77713) );
  NOR U97696 ( .A(n77714), .B(n77713), .Z(n83578) );
  XOR U97697 ( .A(n83576), .B(n83578), .Z(n83590) );
  IV U97698 ( .A(n77715), .Z(n77716) );
  NOR U97699 ( .A(n77717), .B(n77716), .Z(n77721) );
  NOR U97700 ( .A(n77719), .B(n77718), .Z(n77720) );
  NOR U97701 ( .A(n77721), .B(n77720), .Z(n83591) );
  IV U97702 ( .A(n83591), .Z(n83579) );
  XOR U97703 ( .A(n83590), .B(n83579), .Z(n83587) );
  XOR U97704 ( .A(n77722), .B(n83587), .Z(n83605) );
  IV U97705 ( .A(n83605), .Z(n83608) );
  XOR U97706 ( .A(n83606), .B(n83608), .Z(n83601) );
  IV U97707 ( .A(n77723), .Z(n77725) );
  NOR U97708 ( .A(n77725), .B(n77724), .Z(n83610) );
  IV U97709 ( .A(n77726), .Z(n77727) );
  NOR U97710 ( .A(n77728), .B(n77727), .Z(n83600) );
  NOR U97711 ( .A(n83610), .B(n83600), .Z(n77729) );
  XOR U97712 ( .A(n83601), .B(n77729), .Z(n77730) );
  IV U97713 ( .A(n77730), .Z(n83599) );
  IV U97714 ( .A(n77731), .Z(n77732) );
  NOR U97715 ( .A(n77733), .B(n77732), .Z(n77738) );
  IV U97716 ( .A(n77734), .Z(n77735) );
  NOR U97717 ( .A(n77736), .B(n77735), .Z(n77737) );
  NOR U97718 ( .A(n77738), .B(n77737), .Z(n83598) );
  XOR U97719 ( .A(n83599), .B(n83598), .Z(n83571) );
  IV U97720 ( .A(n77739), .Z(n77740) );
  NOR U97721 ( .A(n77740), .B(n77742), .Z(n83573) );
  IV U97722 ( .A(n77741), .Z(n77743) );
  NOR U97723 ( .A(n77743), .B(n77742), .Z(n83570) );
  NOR U97724 ( .A(n83573), .B(n83570), .Z(n77744) );
  XOR U97725 ( .A(n83571), .B(n77744), .Z(n83616) );
  XOR U97726 ( .A(n83614), .B(n83616), .Z(n83618) );
  XOR U97727 ( .A(n83617), .B(n83618), .Z(n83568) );
  XOR U97728 ( .A(n77745), .B(n83568), .Z(n83560) );
  XOR U97729 ( .A(n83628), .B(n83560), .Z(n83639) );
  XOR U97730 ( .A(n77753), .B(n83639), .Z(n83553) );
  IV U97731 ( .A(n77746), .Z(n77747) );
  NOR U97732 ( .A(n77749), .B(n77747), .Z(n83549) );
  IV U97733 ( .A(n77748), .Z(n77750) );
  NOR U97734 ( .A(n77750), .B(n77749), .Z(n83551) );
  IV U97735 ( .A(n77751), .Z(n83643) );
  NOR U97736 ( .A(n77752), .B(n83643), .Z(n83554) );
  XOR U97737 ( .A(n83645), .B(n83647), .Z(n83649) );
  XOR U97738 ( .A(n83648), .B(n83649), .Z(n83548) );
  XOR U97739 ( .A(n77754), .B(n83548), .Z(n83655) );
  IV U97740 ( .A(n77755), .Z(n77756) );
  NOR U97741 ( .A(n77756), .B(n77762), .Z(n77757) );
  IV U97742 ( .A(n77757), .Z(n83656) );
  XOR U97743 ( .A(n83655), .B(n83656), .Z(n83663) );
  IV U97744 ( .A(n77758), .Z(n77759) );
  NOR U97745 ( .A(n77760), .B(n77759), .Z(n83543) );
  IV U97746 ( .A(n77761), .Z(n77763) );
  NOR U97747 ( .A(n77763), .B(n77762), .Z(n83661) );
  NOR U97748 ( .A(n83543), .B(n83661), .Z(n77764) );
  XOR U97749 ( .A(n83663), .B(n77764), .Z(n77765) );
  IV U97750 ( .A(n77765), .Z(n83537) );
  IV U97751 ( .A(n77766), .Z(n77771) );
  IV U97752 ( .A(n77767), .Z(n77768) );
  NOR U97753 ( .A(n77771), .B(n77768), .Z(n83535) );
  XOR U97754 ( .A(n83537), .B(n83535), .Z(n83540) );
  NOR U97755 ( .A(n77778), .B(n83540), .Z(n89242) );
  IV U97756 ( .A(n77769), .Z(n77770) );
  NOR U97757 ( .A(n77771), .B(n77770), .Z(n83538) );
  XOR U97758 ( .A(n83540), .B(n83538), .Z(n83668) );
  IV U97759 ( .A(n77772), .Z(n77777) );
  NOR U97760 ( .A(n77774), .B(n77773), .Z(n77775) );
  IV U97761 ( .A(n77775), .Z(n77776) );
  NOR U97762 ( .A(n77777), .B(n77776), .Z(n77779) );
  IV U97763 ( .A(n77779), .Z(n83667) );
  XOR U97764 ( .A(n83668), .B(n83667), .Z(n77781) );
  NOR U97765 ( .A(n77779), .B(n77778), .Z(n77780) );
  NOR U97766 ( .A(n77781), .B(n77780), .Z(n77782) );
  NOR U97767 ( .A(n89242), .B(n77782), .Z(n77794) );
  IV U97768 ( .A(n77794), .Z(n83534) );
  IV U97769 ( .A(n77783), .Z(n77784) );
  NOR U97770 ( .A(n77784), .B(n77788), .Z(n77796) );
  IV U97771 ( .A(n77796), .Z(n77785) );
  NOR U97772 ( .A(n83534), .B(n77785), .Z(n89245) );
  IV U97773 ( .A(n77786), .Z(n77792) );
  IV U97774 ( .A(n77787), .Z(n77789) );
  NOR U97775 ( .A(n77789), .B(n77788), .Z(n77790) );
  IV U97776 ( .A(n77790), .Z(n77791) );
  NOR U97777 ( .A(n77792), .B(n77791), .Z(n77793) );
  IV U97778 ( .A(n77793), .Z(n83533) );
  XOR U97779 ( .A(n77794), .B(n83533), .Z(n83531) );
  IV U97780 ( .A(n83531), .Z(n77795) );
  NOR U97781 ( .A(n77796), .B(n77795), .Z(n77797) );
  NOR U97782 ( .A(n89245), .B(n77797), .Z(n83528) );
  IV U97783 ( .A(n77798), .Z(n77799) );
  NOR U97784 ( .A(n77800), .B(n77799), .Z(n83674) );
  IV U97785 ( .A(n77801), .Z(n77803) );
  NOR U97786 ( .A(n77803), .B(n77802), .Z(n83530) );
  NOR U97787 ( .A(n83674), .B(n83530), .Z(n77804) );
  XOR U97788 ( .A(n83528), .B(n77804), .Z(n83679) );
  XOR U97789 ( .A(n83527), .B(n83679), .Z(n83526) );
  IV U97790 ( .A(n77805), .Z(n77806) );
  NOR U97791 ( .A(n77807), .B(n77806), .Z(n83677) );
  IV U97792 ( .A(n77808), .Z(n77809) );
  NOR U97793 ( .A(n77810), .B(n77809), .Z(n83524) );
  NOR U97794 ( .A(n83677), .B(n83524), .Z(n77811) );
  XOR U97795 ( .A(n83526), .B(n77811), .Z(n83521) );
  IV U97796 ( .A(n77812), .Z(n77814) );
  NOR U97797 ( .A(n77814), .B(n77813), .Z(n77815) );
  IV U97798 ( .A(n77815), .Z(n83522) );
  XOR U97799 ( .A(n83521), .B(n83522), .Z(n83681) );
  XOR U97800 ( .A(n83680), .B(n83681), .Z(n83685) );
  IV U97801 ( .A(n77816), .Z(n77817) );
  NOR U97802 ( .A(n77818), .B(n77817), .Z(n83683) );
  XOR U97803 ( .A(n83685), .B(n83683), .Z(n83519) );
  IV U97804 ( .A(n77819), .Z(n77820) );
  NOR U97805 ( .A(n77821), .B(n77820), .Z(n83518) );
  IV U97806 ( .A(n77822), .Z(n77824) );
  NOR U97807 ( .A(n77824), .B(n77823), .Z(n83513) );
  NOR U97808 ( .A(n83518), .B(n83513), .Z(n77825) );
  XOR U97809 ( .A(n83519), .B(n77825), .Z(n77826) );
  IV U97810 ( .A(n77826), .Z(n83517) );
  XOR U97811 ( .A(n83515), .B(n83517), .Z(n83511) );
  XOR U97812 ( .A(n77827), .B(n83511), .Z(n77835) );
  IV U97813 ( .A(n77828), .Z(n77830) );
  NOR U97814 ( .A(n77830), .B(n77829), .Z(n83504) );
  IV U97815 ( .A(n77831), .Z(n77832) );
  NOR U97816 ( .A(n77833), .B(n77832), .Z(n83499) );
  NOR U97817 ( .A(n83504), .B(n83499), .Z(n77834) );
  XOR U97818 ( .A(n77835), .B(n77834), .Z(n83497) );
  XOR U97819 ( .A(n77836), .B(n83497), .Z(n83487) );
  XOR U97820 ( .A(n83488), .B(n83487), .Z(n83492) );
  NOR U97821 ( .A(n77837), .B(n83492), .Z(n89177) );
  IV U97822 ( .A(n77838), .Z(n77843) );
  IV U97823 ( .A(n77839), .Z(n77840) );
  NOR U97824 ( .A(n77843), .B(n77840), .Z(n83490) );
  XOR U97825 ( .A(n83492), .B(n83490), .Z(n83486) );
  IV U97826 ( .A(n77841), .Z(n77842) );
  NOR U97827 ( .A(n77843), .B(n77842), .Z(n77844) );
  IV U97828 ( .A(n77844), .Z(n83485) );
  XOR U97829 ( .A(n83486), .B(n83485), .Z(n77845) );
  NOR U97830 ( .A(n77846), .B(n77845), .Z(n77847) );
  NOR U97831 ( .A(n89177), .B(n77847), .Z(n83694) );
  XOR U97832 ( .A(n77848), .B(n83694), .Z(n83482) );
  XOR U97833 ( .A(n77849), .B(n83482), .Z(n83698) );
  XOR U97834 ( .A(n83697), .B(n83698), .Z(n83701) );
  XOR U97835 ( .A(n83700), .B(n83701), .Z(n83706) );
  XOR U97836 ( .A(n83704), .B(n83706), .Z(n83708) );
  XOR U97837 ( .A(n83707), .B(n83708), .Z(n83475) );
  XOR U97838 ( .A(n77850), .B(n83475), .Z(n77851) );
  XOR U97839 ( .A(n83474), .B(n77851), .Z(n83465) );
  XOR U97840 ( .A(n83464), .B(n83465), .Z(n83468) );
  XOR U97841 ( .A(n83467), .B(n83468), .Z(n83712) );
  IV U97842 ( .A(n77852), .Z(n83458) );
  NOR U97843 ( .A(n77853), .B(n83458), .Z(n77854) );
  NOR U97844 ( .A(n83711), .B(n77854), .Z(n77855) );
  XOR U97845 ( .A(n83712), .B(n77855), .Z(n83450) );
  XOR U97846 ( .A(n83448), .B(n83450), .Z(n83728) );
  XOR U97847 ( .A(n77856), .B(n83728), .Z(n83740) );
  XOR U97848 ( .A(n83741), .B(n83740), .Z(n83744) );
  XOR U97849 ( .A(n83743), .B(n83744), .Z(n83443) );
  IV U97850 ( .A(n77857), .Z(n77858) );
  NOR U97851 ( .A(n77859), .B(n77858), .Z(n83444) );
  IV U97852 ( .A(n77860), .Z(n77862) );
  IV U97853 ( .A(n77861), .Z(n77865) );
  NOR U97854 ( .A(n77862), .B(n77865), .Z(n83441) );
  NOR U97855 ( .A(n83444), .B(n83441), .Z(n77863) );
  XOR U97856 ( .A(n83443), .B(n77863), .Z(n83438) );
  IV U97857 ( .A(n77864), .Z(n77866) );
  NOR U97858 ( .A(n77866), .B(n77865), .Z(n77867) );
  IV U97859 ( .A(n77867), .Z(n83439) );
  XOR U97860 ( .A(n83438), .B(n83439), .Z(n83749) );
  XOR U97861 ( .A(n83748), .B(n83749), .Z(n83436) );
  IV U97862 ( .A(n77868), .Z(n83428) );
  NOR U97863 ( .A(n77869), .B(n83428), .Z(n77873) );
  IV U97864 ( .A(n77870), .Z(n77871) );
  NOR U97865 ( .A(n77872), .B(n77871), .Z(n83434) );
  NOR U97866 ( .A(n77873), .B(n83434), .Z(n77874) );
  XOR U97867 ( .A(n83436), .B(n77874), .Z(n83421) );
  XOR U97868 ( .A(n77875), .B(n83421), .Z(n83414) );
  XOR U97869 ( .A(n83413), .B(n83414), .Z(n83417) );
  XOR U97870 ( .A(n83416), .B(n83417), .Z(n83764) );
  XOR U97871 ( .A(n83763), .B(n83764), .Z(n83768) );
  XOR U97872 ( .A(n83766), .B(n83768), .Z(n83410) );
  XOR U97873 ( .A(n77876), .B(n83410), .Z(n77877) );
  IV U97874 ( .A(n77877), .Z(n83407) );
  XOR U97875 ( .A(n83405), .B(n83407), .Z(n83399) );
  XOR U97876 ( .A(n83398), .B(n83399), .Z(n83386) );
  NOR U97877 ( .A(n77878), .B(n83395), .Z(n77882) );
  IV U97878 ( .A(n77879), .Z(n83387) );
  NOR U97879 ( .A(n77880), .B(n83387), .Z(n77881) );
  NOR U97880 ( .A(n77882), .B(n77881), .Z(n77883) );
  XOR U97881 ( .A(n83386), .B(n77883), .Z(n83378) );
  IV U97882 ( .A(n77884), .Z(n77885) );
  NOR U97883 ( .A(n77887), .B(n77885), .Z(n83776) );
  IV U97884 ( .A(n77886), .Z(n77890) );
  NOR U97885 ( .A(n77888), .B(n77887), .Z(n77889) );
  IV U97886 ( .A(n77889), .Z(n77896) );
  NOR U97887 ( .A(n77890), .B(n77896), .Z(n83379) );
  NOR U97888 ( .A(n83776), .B(n83379), .Z(n77891) );
  XOR U97889 ( .A(n83378), .B(n77891), .Z(n83376) );
  IV U97890 ( .A(n83376), .Z(n77899) );
  IV U97891 ( .A(n77892), .Z(n77893) );
  NOR U97892 ( .A(n77894), .B(n77893), .Z(n83374) );
  IV U97893 ( .A(n77895), .Z(n77897) );
  NOR U97894 ( .A(n77897), .B(n77896), .Z(n83381) );
  NOR U97895 ( .A(n83374), .B(n83381), .Z(n77898) );
  XOR U97896 ( .A(n77899), .B(n77898), .Z(n83368) );
  IV U97897 ( .A(n77900), .Z(n77901) );
  NOR U97898 ( .A(n77902), .B(n77901), .Z(n83366) );
  XOR U97899 ( .A(n83368), .B(n83366), .Z(n83371) );
  XOR U97900 ( .A(n83369), .B(n83371), .Z(n83788) );
  XOR U97901 ( .A(n77903), .B(n83788), .Z(n77904) );
  IV U97902 ( .A(n77904), .Z(n83793) );
  IV U97903 ( .A(n77905), .Z(n77909) );
  NOR U97904 ( .A(n77907), .B(n77906), .Z(n77908) );
  IV U97905 ( .A(n77908), .Z(n77912) );
  NOR U97906 ( .A(n77909), .B(n77912), .Z(n77910) );
  IV U97907 ( .A(n77910), .Z(n83786) );
  IV U97908 ( .A(n77911), .Z(n77913) );
  NOR U97909 ( .A(n77913), .B(n77912), .Z(n77914) );
  IV U97910 ( .A(n77914), .Z(n83792) );
  XOR U97911 ( .A(n83786), .B(n83792), .Z(n77915) );
  XOR U97912 ( .A(n83793), .B(n77915), .Z(n89493) );
  IV U97913 ( .A(n77916), .Z(n77917) );
  NOR U97914 ( .A(n77918), .B(n77917), .Z(n89491) );
  IV U97915 ( .A(n77919), .Z(n77921) );
  NOR U97916 ( .A(n77921), .B(n77920), .Z(n89492) );
  NOR U97917 ( .A(n89491), .B(n89492), .Z(n83796) );
  XOR U97918 ( .A(n89493), .B(n83796), .Z(n77926) );
  IV U97919 ( .A(n77926), .Z(n89103) );
  XOR U97920 ( .A(n83794), .B(n89103), .Z(n77922) );
  NOR U97921 ( .A(n77923), .B(n77922), .Z(n89098) );
  NOR U97922 ( .A(n77924), .B(n89106), .Z(n83364) );
  NOR U97923 ( .A(n83794), .B(n83364), .Z(n77925) );
  XOR U97924 ( .A(n77926), .B(n77925), .Z(n77938) );
  IV U97925 ( .A(n77938), .Z(n77927) );
  NOR U97926 ( .A(n77928), .B(n77927), .Z(n77929) );
  NOR U97927 ( .A(n89098), .B(n77929), .Z(n83356) );
  IV U97928 ( .A(n77930), .Z(n77934) );
  NOR U97929 ( .A(n77932), .B(n77931), .Z(n77933) );
  IV U97930 ( .A(n77933), .Z(n77954) );
  NOR U97931 ( .A(n77934), .B(n77954), .Z(n77950) );
  IV U97932 ( .A(n77950), .Z(n83357) );
  NOR U97933 ( .A(n83356), .B(n83357), .Z(n77952) );
  NOR U97934 ( .A(n77935), .B(n77939), .Z(n77936) );
  NOR U97935 ( .A(n83356), .B(n77936), .Z(n77947) );
  IV U97936 ( .A(n77937), .Z(n77941) );
  NOR U97937 ( .A(n77939), .B(n77938), .Z(n77940) );
  IV U97938 ( .A(n77940), .Z(n77943) );
  NOR U97939 ( .A(n77941), .B(n77943), .Z(n89078) );
  IV U97940 ( .A(n77942), .Z(n77944) );
  NOR U97941 ( .A(n77944), .B(n77943), .Z(n89081) );
  NOR U97942 ( .A(n89078), .B(n89081), .Z(n77945) );
  IV U97943 ( .A(n77945), .Z(n77946) );
  NOR U97944 ( .A(n77947), .B(n77946), .Z(n77948) );
  IV U97945 ( .A(n77948), .Z(n77949) );
  NOR U97946 ( .A(n77950), .B(n77949), .Z(n77951) );
  NOR U97947 ( .A(n77952), .B(n77951), .Z(n83361) );
  IV U97948 ( .A(n77953), .Z(n77955) );
  NOR U97949 ( .A(n77955), .B(n77954), .Z(n83359) );
  XOR U97950 ( .A(n83361), .B(n83359), .Z(n83353) );
  IV U97951 ( .A(n77956), .Z(n77966) );
  IV U97952 ( .A(n77957), .Z(n77958) );
  NOR U97953 ( .A(n77966), .B(n77958), .Z(n83347) );
  NOR U97954 ( .A(n83347), .B(n77959), .Z(n77960) );
  XOR U97955 ( .A(n83353), .B(n77960), .Z(n77961) );
  IV U97956 ( .A(n77961), .Z(n83805) );
  IV U97957 ( .A(n77962), .Z(n77963) );
  NOR U97958 ( .A(n77964), .B(n77963), .Z(n83344) );
  IV U97959 ( .A(n77965), .Z(n77967) );
  NOR U97960 ( .A(n77967), .B(n77966), .Z(n83803) );
  NOR U97961 ( .A(n83344), .B(n83803), .Z(n77968) );
  XOR U97962 ( .A(n83805), .B(n77968), .Z(n83342) );
  IV U97963 ( .A(n77969), .Z(n77970) );
  NOR U97964 ( .A(n77970), .B(n77972), .Z(n83341) );
  IV U97965 ( .A(n77971), .Z(n77975) );
  NOR U97966 ( .A(n77973), .B(n77972), .Z(n77974) );
  IV U97967 ( .A(n77974), .Z(n77978) );
  NOR U97968 ( .A(n77975), .B(n77978), .Z(n83809) );
  NOR U97969 ( .A(n83341), .B(n83809), .Z(n77976) );
  XOR U97970 ( .A(n83342), .B(n77976), .Z(n83814) );
  IV U97971 ( .A(n77977), .Z(n77979) );
  NOR U97972 ( .A(n77979), .B(n77978), .Z(n83812) );
  XOR U97973 ( .A(n83814), .B(n83812), .Z(n83816) );
  XOR U97974 ( .A(n83815), .B(n83816), .Z(n83339) );
  NOR U97975 ( .A(n77986), .B(n83339), .Z(n89539) );
  IV U97976 ( .A(n77980), .Z(n77982) );
  NOR U97977 ( .A(n77982), .B(n77981), .Z(n83338) );
  XOR U97978 ( .A(n83338), .B(n83339), .Z(n83337) );
  IV U97979 ( .A(n77983), .Z(n77984) );
  NOR U97980 ( .A(n77985), .B(n77984), .Z(n77987) );
  IV U97981 ( .A(n77987), .Z(n83336) );
  XOR U97982 ( .A(n83337), .B(n83336), .Z(n77989) );
  NOR U97983 ( .A(n77987), .B(n77986), .Z(n77988) );
  NOR U97984 ( .A(n77989), .B(n77988), .Z(n77990) );
  NOR U97985 ( .A(n89539), .B(n77990), .Z(n83333) );
  IV U97986 ( .A(n77991), .Z(n77993) );
  NOR U97987 ( .A(n77993), .B(n77992), .Z(n77994) );
  IV U97988 ( .A(n77994), .Z(n83334) );
  XOR U97989 ( .A(n83333), .B(n83334), .Z(n83327) );
  IV U97990 ( .A(n83327), .Z(n83325) );
  IV U97991 ( .A(n77995), .Z(n77996) );
  NOR U97992 ( .A(n77997), .B(n77996), .Z(n83326) );
  IV U97993 ( .A(n77998), .Z(n78000) );
  NOR U97994 ( .A(n78000), .B(n77999), .Z(n83330) );
  NOR U97995 ( .A(n83326), .B(n83330), .Z(n78001) );
  XOR U97996 ( .A(n83325), .B(n78001), .Z(n83324) );
  XOR U97997 ( .A(n83322), .B(n83324), .Z(n78002) );
  XOR U97998 ( .A(n83323), .B(n78002), .Z(n83821) );
  IV U97999 ( .A(n78003), .Z(n78005) );
  NOR U98000 ( .A(n78005), .B(n78004), .Z(n83319) );
  IV U98001 ( .A(n78006), .Z(n78008) );
  NOR U98002 ( .A(n78008), .B(n78007), .Z(n83820) );
  NOR U98003 ( .A(n83319), .B(n83820), .Z(n78009) );
  XOR U98004 ( .A(n83821), .B(n78009), .Z(n78010) );
  NOR U98005 ( .A(n78011), .B(n78010), .Z(n78014) );
  IV U98006 ( .A(n78011), .Z(n78013) );
  XOR U98007 ( .A(n83319), .B(n83821), .Z(n78012) );
  NOR U98008 ( .A(n78013), .B(n78012), .Z(n83827) );
  NOR U98009 ( .A(n78014), .B(n83827), .Z(n78015) );
  IV U98010 ( .A(n78015), .Z(n83825) );
  IV U98011 ( .A(n78016), .Z(n78017) );
  NOR U98012 ( .A(n78018), .B(n78017), .Z(n83823) );
  XOR U98013 ( .A(n83825), .B(n83823), .Z(n83830) );
  IV U98014 ( .A(n78019), .Z(n78021) );
  NOR U98015 ( .A(n78021), .B(n78020), .Z(n83317) );
  IV U98016 ( .A(n78022), .Z(n78023) );
  NOR U98017 ( .A(n78023), .B(n78027), .Z(n83829) );
  NOR U98018 ( .A(n83317), .B(n83829), .Z(n78024) );
  XOR U98019 ( .A(n83830), .B(n78024), .Z(n78025) );
  IV U98020 ( .A(n78025), .Z(n83834) );
  NOR U98021 ( .A(n78027), .B(n78026), .Z(n78028) );
  IV U98022 ( .A(n78028), .Z(n78035) );
  XOR U98023 ( .A(n78030), .B(n78029), .Z(n78032) );
  NOR U98024 ( .A(n78032), .B(n78031), .Z(n78033) );
  IV U98025 ( .A(n78033), .Z(n78034) );
  NOR U98026 ( .A(n78035), .B(n78034), .Z(n83832) );
  XOR U98027 ( .A(n83834), .B(n83832), .Z(n83836) );
  XOR U98028 ( .A(n83835), .B(n83836), .Z(n83309) );
  XOR U98029 ( .A(n83306), .B(n83309), .Z(n83840) );
  XOR U98030 ( .A(n78036), .B(n83840), .Z(n83849) );
  XOR U98031 ( .A(n78037), .B(n83849), .Z(n83848) );
  XOR U98032 ( .A(n83846), .B(n83848), .Z(n83300) );
  XOR U98033 ( .A(n78038), .B(n83300), .Z(n83291) );
  IV U98034 ( .A(n78039), .Z(n78040) );
  NOR U98035 ( .A(n78041), .B(n78040), .Z(n83293) );
  IV U98036 ( .A(n78042), .Z(n78044) );
  NOR U98037 ( .A(n78044), .B(n78043), .Z(n83290) );
  NOR U98038 ( .A(n83293), .B(n83290), .Z(n78045) );
  XOR U98039 ( .A(n83291), .B(n78045), .Z(n83286) );
  IV U98040 ( .A(n78046), .Z(n78050) );
  NOR U98041 ( .A(n83286), .B(n78050), .Z(n89002) );
  IV U98042 ( .A(n78047), .Z(n78049) );
  NOR U98043 ( .A(n78049), .B(n78048), .Z(n83284) );
  XOR U98044 ( .A(n83284), .B(n83286), .Z(n83288) );
  IV U98045 ( .A(n83288), .Z(n78051) );
  XOR U98046 ( .A(n83287), .B(n78051), .Z(n78053) );
  NOR U98047 ( .A(n78051), .B(n78050), .Z(n78052) );
  NOR U98048 ( .A(n78053), .B(n78052), .Z(n78054) );
  NOR U98049 ( .A(n89002), .B(n78054), .Z(n83858) );
  XOR U98050 ( .A(n78055), .B(n83858), .Z(n83861) );
  XOR U98051 ( .A(n83860), .B(n83861), .Z(n83278) );
  XOR U98052 ( .A(n83275), .B(n83278), .Z(n83273) );
  XOR U98053 ( .A(n78056), .B(n83273), .Z(n83267) );
  XOR U98054 ( .A(n83268), .B(n83267), .Z(n83881) );
  IV U98055 ( .A(n78057), .Z(n78058) );
  NOR U98056 ( .A(n78058), .B(n78060), .Z(n83877) );
  IV U98057 ( .A(n78059), .Z(n78063) );
  NOR U98058 ( .A(n78061), .B(n78060), .Z(n78062) );
  IV U98059 ( .A(n78062), .Z(n78069) );
  NOR U98060 ( .A(n78063), .B(n78069), .Z(n83880) );
  NOR U98061 ( .A(n83877), .B(n83880), .Z(n78064) );
  XOR U98062 ( .A(n83881), .B(n78064), .Z(n83262) );
  IV U98063 ( .A(n78065), .Z(n78066) );
  NOR U98064 ( .A(n78067), .B(n78066), .Z(n83261) );
  IV U98065 ( .A(n78068), .Z(n78070) );
  NOR U98066 ( .A(n78070), .B(n78069), .Z(n78071) );
  IV U98067 ( .A(n78071), .Z(n83264) );
  XOR U98068 ( .A(n83261), .B(n83264), .Z(n78072) );
  XOR U98069 ( .A(n83262), .B(n78072), .Z(n83892) );
  XOR U98070 ( .A(n78073), .B(n83892), .Z(n83896) );
  XOR U98071 ( .A(n83894), .B(n83896), .Z(n83898) );
  XOR U98072 ( .A(n83897), .B(n83898), .Z(n83902) );
  IV U98073 ( .A(n83902), .Z(n78078) );
  IV U98074 ( .A(n78074), .Z(n78075) );
  NOR U98075 ( .A(n78076), .B(n78075), .Z(n83255) );
  NOR U98076 ( .A(n83901), .B(n83255), .Z(n78077) );
  XOR U98077 ( .A(n78078), .B(n78077), .Z(n83249) );
  XOR U98078 ( .A(n78079), .B(n83249), .Z(n83246) );
  IV U98079 ( .A(n78080), .Z(n78082) );
  NOR U98080 ( .A(n78082), .B(n78081), .Z(n78087) );
  IV U98081 ( .A(n78087), .Z(n78083) );
  NOR U98082 ( .A(n83246), .B(n78083), .Z(n83243) );
  IV U98083 ( .A(n78084), .Z(n78085) );
  NOR U98084 ( .A(n78085), .B(n83248), .Z(n83244) );
  XOR U98085 ( .A(n83244), .B(n83246), .Z(n83235) );
  IV U98086 ( .A(n83235), .Z(n78086) );
  NOR U98087 ( .A(n78087), .B(n78086), .Z(n78091) );
  NOR U98088 ( .A(n83243), .B(n78091), .Z(n78088) );
  NOR U98089 ( .A(n78089), .B(n78088), .Z(n78092) );
  IV U98090 ( .A(n78089), .Z(n78090) );
  NOR U98091 ( .A(n78091), .B(n78090), .Z(n83242) );
  NOR U98092 ( .A(n78092), .B(n83242), .Z(n83907) );
  XOR U98093 ( .A(n78093), .B(n83907), .Z(n83912) );
  XOR U98094 ( .A(n83910), .B(n83912), .Z(n83233) );
  IV U98095 ( .A(n78094), .Z(n78096) );
  NOR U98096 ( .A(n78096), .B(n78095), .Z(n83231) );
  XOR U98097 ( .A(n83233), .B(n83231), .Z(n78103) );
  IV U98098 ( .A(n78103), .Z(n78097) );
  NOR U98099 ( .A(n78098), .B(n78097), .Z(n78100) );
  IV U98100 ( .A(n78098), .Z(n78099) );
  NOR U98101 ( .A(n83912), .B(n78099), .Z(n88965) );
  NOR U98102 ( .A(n78100), .B(n88965), .Z(n78101) );
  NOR U98103 ( .A(n78102), .B(n78101), .Z(n83922) );
  IV U98104 ( .A(n78102), .Z(n78104) );
  NOR U98105 ( .A(n78104), .B(n78103), .Z(n83919) );
  NOR U98106 ( .A(n83922), .B(n83919), .Z(n83229) );
  IV U98107 ( .A(n78105), .Z(n78114) );
  NOR U98108 ( .A(n78106), .B(n78114), .Z(n83923) );
  IV U98109 ( .A(n78107), .Z(n78108) );
  NOR U98110 ( .A(n78109), .B(n78108), .Z(n83920) );
  NOR U98111 ( .A(n83228), .B(n83920), .Z(n78110) );
  IV U98112 ( .A(n78110), .Z(n78111) );
  NOR U98113 ( .A(n83923), .B(n78111), .Z(n78112) );
  XOR U98114 ( .A(n83229), .B(n78112), .Z(n83928) );
  IV U98115 ( .A(n78113), .Z(n78115) );
  NOR U98116 ( .A(n78115), .B(n78114), .Z(n83926) );
  XOR U98117 ( .A(n83928), .B(n83926), .Z(n83930) );
  XOR U98118 ( .A(n83929), .B(n83930), .Z(n83224) );
  IV U98119 ( .A(n78116), .Z(n78118) );
  NOR U98120 ( .A(n78118), .B(n78117), .Z(n83222) );
  XOR U98121 ( .A(n83224), .B(n83222), .Z(n83226) );
  IV U98122 ( .A(n83226), .Z(n78125) );
  IV U98123 ( .A(n78119), .Z(n78120) );
  NOR U98124 ( .A(n78121), .B(n78120), .Z(n83225) );
  NOR U98125 ( .A(n78122), .B(n83216), .Z(n78123) );
  NOR U98126 ( .A(n83225), .B(n78123), .Z(n78124) );
  XOR U98127 ( .A(n78125), .B(n78124), .Z(n83209) );
  IV U98128 ( .A(n78126), .Z(n78132) );
  NOR U98129 ( .A(n78127), .B(n78132), .Z(n78128) );
  IV U98130 ( .A(n78128), .Z(n83208) );
  NOR U98131 ( .A(n78129), .B(n83208), .Z(n78130) );
  XOR U98132 ( .A(n83209), .B(n78130), .Z(n83937) );
  IV U98133 ( .A(n78131), .Z(n78133) );
  NOR U98134 ( .A(n78133), .B(n78132), .Z(n83935) );
  XOR U98135 ( .A(n83937), .B(n83935), .Z(n83939) );
  XOR U98136 ( .A(n78134), .B(n83939), .Z(n78135) );
  IV U98137 ( .A(n78135), .Z(n83200) );
  XOR U98138 ( .A(n83199), .B(n83200), .Z(n83204) );
  IV U98139 ( .A(n78136), .Z(n78138) );
  NOR U98140 ( .A(n78138), .B(n78137), .Z(n83202) );
  XOR U98141 ( .A(n83204), .B(n83202), .Z(n83193) );
  XOR U98142 ( .A(n83192), .B(n83193), .Z(n83946) );
  IV U98143 ( .A(n83946), .Z(n78145) );
  IV U98144 ( .A(n78139), .Z(n78140) );
  NOR U98145 ( .A(n78141), .B(n78140), .Z(n83196) );
  IV U98146 ( .A(n78142), .Z(n78143) );
  NOR U98147 ( .A(n78148), .B(n78143), .Z(n83945) );
  NOR U98148 ( .A(n83196), .B(n83945), .Z(n78144) );
  XOR U98149 ( .A(n78145), .B(n78144), .Z(n83950) );
  XOR U98150 ( .A(n83948), .B(n83950), .Z(n83952) );
  NOR U98151 ( .A(n78146), .B(n83952), .Z(n83190) );
  IV U98152 ( .A(n78147), .Z(n78149) );
  NOR U98153 ( .A(n78149), .B(n78148), .Z(n83951) );
  XOR U98154 ( .A(n83951), .B(n83952), .Z(n83958) );
  IV U98155 ( .A(n83958), .Z(n78150) );
  NOR U98156 ( .A(n78151), .B(n78150), .Z(n83188) );
  NOR U98157 ( .A(n83190), .B(n83188), .Z(n78158) );
  IV U98158 ( .A(n78152), .Z(n78154) );
  NOR U98159 ( .A(n78154), .B(n78153), .Z(n83186) );
  IV U98160 ( .A(n78155), .Z(n78156) );
  NOR U98161 ( .A(n78156), .B(n78163), .Z(n83956) );
  NOR U98162 ( .A(n83186), .B(n83956), .Z(n78157) );
  XOR U98163 ( .A(n78158), .B(n78157), .Z(n83961) );
  IV U98164 ( .A(n78159), .Z(n78160) );
  NOR U98165 ( .A(n78161), .B(n78160), .Z(n83959) );
  IV U98166 ( .A(n78162), .Z(n78164) );
  NOR U98167 ( .A(n78164), .B(n78163), .Z(n83184) );
  NOR U98168 ( .A(n83959), .B(n83184), .Z(n78165) );
  XOR U98169 ( .A(n83961), .B(n78165), .Z(n83181) );
  IV U98170 ( .A(n78166), .Z(n78171) );
  NOR U98171 ( .A(n78168), .B(n78167), .Z(n78169) );
  IV U98172 ( .A(n78169), .Z(n78170) );
  NOR U98173 ( .A(n78171), .B(n78170), .Z(n78172) );
  IV U98174 ( .A(n78172), .Z(n83182) );
  XOR U98175 ( .A(n83181), .B(n83182), .Z(n83962) );
  XOR U98176 ( .A(n83963), .B(n83962), .Z(n83179) );
  IV U98177 ( .A(n78173), .Z(n78174) );
  NOR U98178 ( .A(n78175), .B(n78174), .Z(n83178) );
  NOR U98179 ( .A(n83966), .B(n78176), .Z(n78177) );
  NOR U98180 ( .A(n83178), .B(n78177), .Z(n78178) );
  XOR U98181 ( .A(n83179), .B(n78178), .Z(n83177) );
  XOR U98182 ( .A(n83171), .B(n83177), .Z(n78179) );
  XOR U98183 ( .A(n78180), .B(n78179), .Z(n83165) );
  IV U98184 ( .A(n78181), .Z(n78183) );
  NOR U98185 ( .A(n78183), .B(n78182), .Z(n83168) );
  IV U98186 ( .A(n78184), .Z(n78186) );
  IV U98187 ( .A(n78185), .Z(n78189) );
  NOR U98188 ( .A(n78186), .B(n78189), .Z(n83166) );
  NOR U98189 ( .A(n83168), .B(n83166), .Z(n78187) );
  XOR U98190 ( .A(n83165), .B(n78187), .Z(n83164) );
  IV U98191 ( .A(n78188), .Z(n78192) );
  NOR U98192 ( .A(n78190), .B(n78189), .Z(n78191) );
  IV U98193 ( .A(n78191), .Z(n78194) );
  NOR U98194 ( .A(n78192), .B(n78194), .Z(n83162) );
  XOR U98195 ( .A(n83164), .B(n83162), .Z(n83157) );
  IV U98196 ( .A(n83157), .Z(n83155) );
  IV U98197 ( .A(n78193), .Z(n78195) );
  NOR U98198 ( .A(n78195), .B(n78194), .Z(n83154) );
  IV U98199 ( .A(n83154), .Z(n83156) );
  XOR U98200 ( .A(n83155), .B(n83156), .Z(n83152) );
  IV U98201 ( .A(n78196), .Z(n78197) );
  NOR U98202 ( .A(n78198), .B(n78197), .Z(n83159) );
  IV U98203 ( .A(n78199), .Z(n78201) );
  NOR U98204 ( .A(n78201), .B(n78200), .Z(n83151) );
  NOR U98205 ( .A(n83159), .B(n83151), .Z(n78202) );
  XOR U98206 ( .A(n83152), .B(n78202), .Z(n78203) );
  IV U98207 ( .A(n78203), .Z(n83147) );
  XOR U98208 ( .A(n83145), .B(n83147), .Z(n83149) );
  XOR U98209 ( .A(n83148), .B(n83149), .Z(n83978) );
  XOR U98210 ( .A(n83977), .B(n83978), .Z(n83993) );
  XOR U98211 ( .A(n78204), .B(n83993), .Z(n83989) );
  XOR U98212 ( .A(n83990), .B(n83989), .Z(n84002) );
  XOR U98213 ( .A(n84003), .B(n84002), .Z(n83997) );
  XOR U98214 ( .A(n78205), .B(n83997), .Z(n83141) );
  XOR U98215 ( .A(n83139), .B(n83141), .Z(n84015) );
  XOR U98216 ( .A(n84014), .B(n84015), .Z(n84018) );
  XOR U98217 ( .A(n84017), .B(n84018), .Z(n84026) );
  XOR U98218 ( .A(n84027), .B(n84026), .Z(n83135) );
  NOR U98219 ( .A(n78221), .B(n78206), .Z(n78207) );
  IV U98220 ( .A(n78207), .Z(n78211) );
  IV U98221 ( .A(n78208), .Z(n78213) );
  NOR U98222 ( .A(n78209), .B(n78213), .Z(n78210) );
  IV U98223 ( .A(n78210), .Z(n78220) );
  NOR U98224 ( .A(n78211), .B(n78220), .Z(n83137) );
  IV U98225 ( .A(n78212), .Z(n78214) );
  NOR U98226 ( .A(n78214), .B(n78213), .Z(n84029) );
  NOR U98227 ( .A(n83137), .B(n84029), .Z(n78215) );
  XOR U98228 ( .A(n83135), .B(n78215), .Z(n83133) );
  IV U98229 ( .A(n78216), .Z(n78217) );
  NOR U98230 ( .A(n78218), .B(n78217), .Z(n83131) );
  IV U98231 ( .A(n78219), .Z(n78224) );
  NOR U98232 ( .A(n78221), .B(n78220), .Z(n78222) );
  IV U98233 ( .A(n78222), .Z(n78223) );
  NOR U98234 ( .A(n78224), .B(n78223), .Z(n83134) );
  XOR U98235 ( .A(n83131), .B(n83134), .Z(n78225) );
  XOR U98236 ( .A(n83133), .B(n78225), .Z(n84035) );
  XOR U98237 ( .A(n84033), .B(n84035), .Z(n84038) );
  XOR U98238 ( .A(n84036), .B(n84038), .Z(n83129) );
  XOR U98239 ( .A(n83130), .B(n83129), .Z(n84047) );
  XOR U98240 ( .A(n84049), .B(n84047), .Z(n83126) );
  XOR U98241 ( .A(n78226), .B(n83126), .Z(n78227) );
  IV U98242 ( .A(n78227), .Z(n83123) );
  XOR U98243 ( .A(n78228), .B(n83123), .Z(n78236) );
  IV U98244 ( .A(n78236), .Z(n78229) );
  NOR U98245 ( .A(n78230), .B(n78229), .Z(n88789) );
  IV U98246 ( .A(n78231), .Z(n78233) );
  NOR U98247 ( .A(n78233), .B(n78232), .Z(n78237) );
  IV U98248 ( .A(n78237), .Z(n78235) );
  XOR U98249 ( .A(n83121), .B(n83123), .Z(n78234) );
  NOR U98250 ( .A(n78235), .B(n78234), .Z(n88792) );
  NOR U98251 ( .A(n78237), .B(n78236), .Z(n78238) );
  NOR U98252 ( .A(n88792), .B(n78238), .Z(n83115) );
  NOR U98253 ( .A(n78239), .B(n83115), .Z(n78240) );
  NOR U98254 ( .A(n88789), .B(n78240), .Z(n84069) );
  XOR U98255 ( .A(n78241), .B(n84069), .Z(n84067) );
  XOR U98256 ( .A(n78242), .B(n84067), .Z(n78243) );
  IV U98257 ( .A(n78243), .Z(n84076) );
  XOR U98258 ( .A(n84075), .B(n84076), .Z(n84079) );
  XOR U98259 ( .A(n84080), .B(n84079), .Z(n84081) );
  IV U98260 ( .A(n78244), .Z(n78248) );
  NOR U98261 ( .A(n78246), .B(n78245), .Z(n78247) );
  IV U98262 ( .A(n78247), .Z(n78254) );
  NOR U98263 ( .A(n78248), .B(n78254), .Z(n78249) );
  IV U98264 ( .A(n78249), .Z(n84082) );
  XOR U98265 ( .A(n84081), .B(n84082), .Z(n84085) );
  IV U98266 ( .A(n78250), .Z(n78252) );
  NOR U98267 ( .A(n78252), .B(n78251), .Z(n83110) );
  IV U98268 ( .A(n78253), .Z(n78255) );
  NOR U98269 ( .A(n78255), .B(n78254), .Z(n84086) );
  NOR U98270 ( .A(n83110), .B(n84086), .Z(n78256) );
  XOR U98271 ( .A(n84085), .B(n78256), .Z(n84095) );
  XOR U98272 ( .A(n78257), .B(n84095), .Z(n83109) );
  XOR U98273 ( .A(n78258), .B(n83109), .Z(n78266) );
  IV U98274 ( .A(n78266), .Z(n78259) );
  NOR U98275 ( .A(n78260), .B(n78259), .Z(n89805) );
  IV U98276 ( .A(n78261), .Z(n78262) );
  NOR U98277 ( .A(n78263), .B(n78262), .Z(n78267) );
  IV U98278 ( .A(n78267), .Z(n78265) );
  XOR U98279 ( .A(n83107), .B(n83109), .Z(n78264) );
  NOR U98280 ( .A(n78265), .B(n78264), .Z(n89802) );
  NOR U98281 ( .A(n78267), .B(n78266), .Z(n78268) );
  NOR U98282 ( .A(n89802), .B(n78268), .Z(n83103) );
  NOR U98283 ( .A(n78269), .B(n83103), .Z(n78270) );
  NOR U98284 ( .A(n89805), .B(n78270), .Z(n84103) );
  IV U98285 ( .A(n78271), .Z(n78275) );
  IV U98286 ( .A(n78272), .Z(n78287) );
  NOR U98287 ( .A(n78273), .B(n78287), .Z(n78274) );
  IV U98288 ( .A(n78274), .Z(n84105) );
  NOR U98289 ( .A(n78275), .B(n84105), .Z(n78277) );
  NOR U98290 ( .A(n78277), .B(n78276), .Z(n78278) );
  XOR U98291 ( .A(n84103), .B(n78278), .Z(n78282) );
  IV U98292 ( .A(n78279), .Z(n78280) );
  NOR U98293 ( .A(n84105), .B(n78280), .Z(n78281) );
  XOR U98294 ( .A(n78282), .B(n78281), .Z(n83101) );
  IV U98295 ( .A(n78283), .Z(n78284) );
  NOR U98296 ( .A(n78285), .B(n78284), .Z(n83097) );
  IV U98297 ( .A(n78286), .Z(n78288) );
  NOR U98298 ( .A(n78288), .B(n78287), .Z(n83099) );
  NOR U98299 ( .A(n83097), .B(n83099), .Z(n78289) );
  XOR U98300 ( .A(n83101), .B(n78289), .Z(n83095) );
  IV U98301 ( .A(n78290), .Z(n78291) );
  NOR U98302 ( .A(n78292), .B(n78291), .Z(n83094) );
  IV U98303 ( .A(n78293), .Z(n78294) );
  NOR U98304 ( .A(n78294), .B(n78297), .Z(n84109) );
  NOR U98305 ( .A(n83094), .B(n84109), .Z(n78295) );
  XOR U98306 ( .A(n83095), .B(n78295), .Z(n83092) );
  IV U98307 ( .A(n78296), .Z(n78298) );
  NOR U98308 ( .A(n78298), .B(n78297), .Z(n83090) );
  XOR U98309 ( .A(n83092), .B(n83090), .Z(n84114) );
  XOR U98310 ( .A(n78299), .B(n84114), .Z(n83080) );
  IV U98311 ( .A(n78300), .Z(n78301) );
  NOR U98312 ( .A(n78302), .B(n78301), .Z(n83085) );
  IV U98313 ( .A(n78303), .Z(n78304) );
  NOR U98314 ( .A(n78305), .B(n78304), .Z(n83082) );
  NOR U98315 ( .A(n83085), .B(n83082), .Z(n78306) );
  XOR U98316 ( .A(n83080), .B(n78306), .Z(n83078) );
  IV U98317 ( .A(n83078), .Z(n78314) );
  IV U98318 ( .A(n78307), .Z(n78308) );
  NOR U98319 ( .A(n78309), .B(n78308), .Z(n83079) );
  IV U98320 ( .A(n78310), .Z(n78312) );
  NOR U98321 ( .A(n78312), .B(n78311), .Z(n83076) );
  NOR U98322 ( .A(n83079), .B(n83076), .Z(n78313) );
  XOR U98323 ( .A(n78314), .B(n78313), .Z(n83071) );
  XOR U98324 ( .A(n83070), .B(n83071), .Z(n83074) );
  IV U98325 ( .A(n78315), .Z(n78317) );
  NOR U98326 ( .A(n78317), .B(n78316), .Z(n83073) );
  IV U98327 ( .A(n78318), .Z(n78320) );
  NOR U98328 ( .A(n78320), .B(n78319), .Z(n83065) );
  NOR U98329 ( .A(n83073), .B(n83065), .Z(n78321) );
  XOR U98330 ( .A(n83074), .B(n78321), .Z(n83061) );
  XOR U98331 ( .A(n78322), .B(n83061), .Z(n83058) );
  XOR U98332 ( .A(n78323), .B(n83058), .Z(n83045) );
  XOR U98333 ( .A(n83043), .B(n83045), .Z(n83047) );
  XOR U98334 ( .A(n83046), .B(n83047), .Z(n83053) );
  XOR U98335 ( .A(n83051), .B(n83053), .Z(n83036) );
  XOR U98336 ( .A(n78324), .B(n83036), .Z(n78331) );
  IV U98337 ( .A(n78331), .Z(n84146) );
  XOR U98338 ( .A(n83015), .B(n84146), .Z(n78325) );
  NOR U98339 ( .A(n78326), .B(n78325), .Z(n83014) );
  IV U98340 ( .A(n78327), .Z(n84149) );
  IV U98341 ( .A(n78328), .Z(n78329) );
  NOR U98342 ( .A(n78330), .B(n78329), .Z(n84145) );
  NOR U98343 ( .A(n84145), .B(n83015), .Z(n78332) );
  XOR U98344 ( .A(n78332), .B(n78331), .Z(n84148) );
  XOR U98345 ( .A(n84149), .B(n84148), .Z(n78333) );
  NOR U98346 ( .A(n78334), .B(n78333), .Z(n78335) );
  NOR U98347 ( .A(n83014), .B(n78335), .Z(n78336) );
  IV U98348 ( .A(n78336), .Z(n83011) );
  XOR U98349 ( .A(n83010), .B(n83011), .Z(n83003) );
  XOR U98350 ( .A(n83002), .B(n83003), .Z(n83007) );
  IV U98351 ( .A(n78337), .Z(n78340) );
  IV U98352 ( .A(n78338), .Z(n78339) );
  NOR U98353 ( .A(n78340), .B(n78339), .Z(n83005) );
  XOR U98354 ( .A(n83007), .B(n83005), .Z(n82997) );
  IV U98355 ( .A(n82997), .Z(n78348) );
  IV U98356 ( .A(n78341), .Z(n78342) );
  NOR U98357 ( .A(n78343), .B(n78342), .Z(n82999) );
  IV U98358 ( .A(n78344), .Z(n78346) );
  NOR U98359 ( .A(n78346), .B(n78345), .Z(n82996) );
  NOR U98360 ( .A(n82999), .B(n82996), .Z(n78347) );
  XOR U98361 ( .A(n78348), .B(n78347), .Z(n84156) );
  XOR U98362 ( .A(n84154), .B(n84156), .Z(n82994) );
  XOR U98363 ( .A(n78349), .B(n82994), .Z(n84161) );
  IV U98364 ( .A(n78350), .Z(n78351) );
  NOR U98365 ( .A(n78352), .B(n78351), .Z(n78353) );
  IV U98366 ( .A(n78353), .Z(n84162) );
  XOR U98367 ( .A(n84161), .B(n84162), .Z(n84166) );
  IV U98368 ( .A(n78354), .Z(n78359) );
  IV U98369 ( .A(n78355), .Z(n78356) );
  NOR U98370 ( .A(n78359), .B(n78356), .Z(n82988) );
  IV U98371 ( .A(n78357), .Z(n78358) );
  NOR U98372 ( .A(n78359), .B(n78358), .Z(n84164) );
  NOR U98373 ( .A(n82988), .B(n84164), .Z(n78360) );
  XOR U98374 ( .A(n84166), .B(n78360), .Z(n78368) );
  IV U98375 ( .A(n78368), .Z(n78361) );
  NOR U98376 ( .A(n78362), .B(n78361), .Z(n82987) );
  IV U98377 ( .A(n78363), .Z(n78365) );
  NOR U98378 ( .A(n78365), .B(n78364), .Z(n78369) );
  IV U98379 ( .A(n78369), .Z(n78367) );
  XOR U98380 ( .A(n84164), .B(n84166), .Z(n78366) );
  NOR U98381 ( .A(n78367), .B(n78366), .Z(n88714) );
  NOR U98382 ( .A(n78369), .B(n78368), .Z(n78370) );
  NOR U98383 ( .A(n88714), .B(n78370), .Z(n82982) );
  NOR U98384 ( .A(n78371), .B(n82982), .Z(n78372) );
  NOR U98385 ( .A(n82987), .B(n78372), .Z(n82977) );
  IV U98386 ( .A(n78373), .Z(n78375) );
  NOR U98387 ( .A(n78375), .B(n78374), .Z(n82983) );
  NOR U98388 ( .A(n78376), .B(n82979), .Z(n78377) );
  NOR U98389 ( .A(n82983), .B(n78377), .Z(n78378) );
  XOR U98390 ( .A(n82977), .B(n78378), .Z(n84172) );
  XOR U98391 ( .A(n82972), .B(n84172), .Z(n78386) );
  IV U98392 ( .A(n78379), .Z(n78381) );
  NOR U98393 ( .A(n78381), .B(n78380), .Z(n84170) );
  IV U98394 ( .A(n78382), .Z(n78384) );
  NOR U98395 ( .A(n78384), .B(n78383), .Z(n82974) );
  NOR U98396 ( .A(n84170), .B(n82974), .Z(n78385) );
  XOR U98397 ( .A(n78386), .B(n78385), .Z(n78400) );
  IV U98398 ( .A(n78400), .Z(n82971) );
  IV U98399 ( .A(n78387), .Z(n78388) );
  NOR U98400 ( .A(n78389), .B(n78388), .Z(n78399) );
  IV U98401 ( .A(n78390), .Z(n78391) );
  NOR U98402 ( .A(n78392), .B(n78391), .Z(n82968) );
  NOR U98403 ( .A(n78399), .B(n82968), .Z(n78393) );
  XOR U98404 ( .A(n82971), .B(n78393), .Z(n84179) );
  IV U98405 ( .A(n78394), .Z(n78395) );
  NOR U98406 ( .A(n78395), .B(n78397), .Z(n78407) );
  IV U98407 ( .A(n78407), .Z(n84181) );
  NOR U98408 ( .A(n84179), .B(n84181), .Z(n78409) );
  IV U98409 ( .A(n78396), .Z(n78398) );
  NOR U98410 ( .A(n78398), .B(n78397), .Z(n78403) );
  IV U98411 ( .A(n78403), .Z(n78402) );
  IV U98412 ( .A(n78399), .Z(n82970) );
  XOR U98413 ( .A(n82970), .B(n78400), .Z(n78401) );
  NOR U98414 ( .A(n78402), .B(n78401), .Z(n88703) );
  NOR U98415 ( .A(n84179), .B(n78403), .Z(n78404) );
  NOR U98416 ( .A(n88703), .B(n78404), .Z(n78405) );
  IV U98417 ( .A(n78405), .Z(n78406) );
  NOR U98418 ( .A(n78407), .B(n78406), .Z(n78408) );
  NOR U98419 ( .A(n78409), .B(n78408), .Z(n84184) );
  IV U98420 ( .A(n78410), .Z(n78411) );
  NOR U98421 ( .A(n78411), .B(n78414), .Z(n84182) );
  XOR U98422 ( .A(n84184), .B(n84182), .Z(n78417) );
  NOR U98423 ( .A(n78412), .B(n78417), .Z(n89960) );
  IV U98424 ( .A(n78413), .Z(n78415) );
  NOR U98425 ( .A(n78415), .B(n78414), .Z(n78419) );
  IV U98426 ( .A(n78419), .Z(n78416) );
  NOR U98427 ( .A(n78416), .B(n84184), .Z(n89971) );
  IV U98428 ( .A(n78417), .Z(n78418) );
  NOR U98429 ( .A(n78419), .B(n78418), .Z(n78420) );
  NOR U98430 ( .A(n89971), .B(n78420), .Z(n78425) );
  NOR U98431 ( .A(n78421), .B(n78425), .Z(n78422) );
  NOR U98432 ( .A(n89960), .B(n78422), .Z(n78423) );
  NOR U98433 ( .A(n78424), .B(n78423), .Z(n82966) );
  IV U98434 ( .A(n78424), .Z(n78427) );
  IV U98435 ( .A(n78425), .Z(n78426) );
  NOR U98436 ( .A(n78427), .B(n78426), .Z(n89990) );
  NOR U98437 ( .A(n82966), .B(n89990), .Z(n84189) );
  IV U98438 ( .A(n78428), .Z(n78429) );
  NOR U98439 ( .A(n78430), .B(n78429), .Z(n82964) );
  IV U98440 ( .A(n78431), .Z(n78432) );
  NOR U98441 ( .A(n78433), .B(n78432), .Z(n84188) );
  NOR U98442 ( .A(n82964), .B(n84188), .Z(n78434) );
  XOR U98443 ( .A(n84189), .B(n78434), .Z(n82963) );
  XOR U98444 ( .A(n82961), .B(n82963), .Z(n84194) );
  XOR U98445 ( .A(n84192), .B(n84194), .Z(n78439) );
  IV U98446 ( .A(n78435), .Z(n78437) );
  IV U98447 ( .A(n78436), .Z(n78443) );
  NOR U98448 ( .A(n78437), .B(n78443), .Z(n78447) );
  IV U98449 ( .A(n78447), .Z(n78438) );
  NOR U98450 ( .A(n78439), .B(n78438), .Z(n78440) );
  IV U98451 ( .A(n78440), .Z(n78441) );
  NOR U98452 ( .A(n78442), .B(n78441), .Z(n89999) );
  IV U98453 ( .A(n78442), .Z(n78444) );
  NOR U98454 ( .A(n78444), .B(n78443), .Z(n84193) );
  NOR U98455 ( .A(n84192), .B(n84193), .Z(n78445) );
  XOR U98456 ( .A(n84194), .B(n78445), .Z(n78446) );
  NOR U98457 ( .A(n78447), .B(n78446), .Z(n78448) );
  NOR U98458 ( .A(n89999), .B(n78448), .Z(n82958) );
  IV U98459 ( .A(n78449), .Z(n78450) );
  NOR U98460 ( .A(n78454), .B(n78450), .Z(n78451) );
  IV U98461 ( .A(n78451), .Z(n82959) );
  XOR U98462 ( .A(n82958), .B(n82959), .Z(n82950) );
  IV U98463 ( .A(n82950), .Z(n82952) );
  IV U98464 ( .A(n78452), .Z(n78453) );
  NOR U98465 ( .A(n78454), .B(n78453), .Z(n82951) );
  IV U98466 ( .A(n82951), .Z(n82949) );
  XOR U98467 ( .A(n82952), .B(n82949), .Z(n82948) );
  IV U98468 ( .A(n78455), .Z(n78457) );
  NOR U98469 ( .A(n78457), .B(n78456), .Z(n82953) );
  IV U98470 ( .A(n78458), .Z(n78459) );
  NOR U98471 ( .A(n78464), .B(n78459), .Z(n82946) );
  NOR U98472 ( .A(n82953), .B(n82946), .Z(n78460) );
  XOR U98473 ( .A(n82948), .B(n78460), .Z(n82944) );
  IV U98474 ( .A(n78461), .Z(n84197) );
  NOR U98475 ( .A(n78462), .B(n84197), .Z(n78466) );
  IV U98476 ( .A(n78463), .Z(n78465) );
  NOR U98477 ( .A(n78465), .B(n78464), .Z(n84211) );
  NOR U98478 ( .A(n78466), .B(n84211), .Z(n78467) );
  XOR U98479 ( .A(n82944), .B(n78467), .Z(n84220) );
  XOR U98480 ( .A(n78468), .B(n84220), .Z(n84216) );
  XOR U98481 ( .A(n84215), .B(n84216), .Z(n82940) );
  XOR U98482 ( .A(n82938), .B(n82940), .Z(n82942) );
  XOR U98483 ( .A(n82941), .B(n82942), .Z(n84229) );
  XOR U98484 ( .A(n78469), .B(n84229), .Z(n82926) );
  XOR U98485 ( .A(n78470), .B(n82926), .Z(n82923) );
  XOR U98486 ( .A(n82921), .B(n82923), .Z(n82924) );
  XOR U98487 ( .A(n82925), .B(n82924), .Z(n78476) );
  IV U98488 ( .A(n78476), .Z(n82918) );
  NOR U98489 ( .A(n78471), .B(n82918), .Z(n88664) );
  IV U98490 ( .A(n78472), .Z(n78473) );
  NOR U98491 ( .A(n78474), .B(n78473), .Z(n78477) );
  IV U98492 ( .A(n78477), .Z(n78475) );
  NOR U98493 ( .A(n78475), .B(n82924), .Z(n82920) );
  NOR U98494 ( .A(n78477), .B(n78476), .Z(n78478) );
  NOR U98495 ( .A(n82920), .B(n78478), .Z(n78479) );
  NOR U98496 ( .A(n78480), .B(n78479), .Z(n78481) );
  NOR U98497 ( .A(n88664), .B(n78481), .Z(n82914) );
  XOR U98498 ( .A(n78482), .B(n82914), .Z(n84243) );
  XOR U98499 ( .A(n84245), .B(n84243), .Z(n88654) );
  IV U98500 ( .A(n78483), .Z(n78485) );
  NOR U98501 ( .A(n78485), .B(n78484), .Z(n78490) );
  IV U98502 ( .A(n78486), .Z(n78488) );
  NOR U98503 ( .A(n78488), .B(n78487), .Z(n78489) );
  NOR U98504 ( .A(n78490), .B(n78489), .Z(n88655) );
  XOR U98505 ( .A(n88654), .B(n88655), .Z(n84249) );
  XOR U98506 ( .A(n84251), .B(n84249), .Z(n84254) );
  IV U98507 ( .A(n78491), .Z(n78493) );
  NOR U98508 ( .A(n78493), .B(n78492), .Z(n84252) );
  XOR U98509 ( .A(n84254), .B(n84252), .Z(n84256) );
  IV U98510 ( .A(n78494), .Z(n78495) );
  NOR U98511 ( .A(n78496), .B(n78495), .Z(n82910) );
  NOR U98512 ( .A(n82910), .B(n78497), .Z(n78498) );
  XOR U98513 ( .A(n84256), .B(n78498), .Z(n84260) );
  IV U98514 ( .A(n78499), .Z(n78500) );
  NOR U98515 ( .A(n78500), .B(n78504), .Z(n84261) );
  NOR U98516 ( .A(n78501), .B(n84261), .Z(n78502) );
  XOR U98517 ( .A(n84260), .B(n78502), .Z(n82909) );
  IV U98518 ( .A(n78503), .Z(n78505) );
  NOR U98519 ( .A(n78505), .B(n78504), .Z(n82907) );
  XOR U98520 ( .A(n82909), .B(n82907), .Z(n84271) );
  XOR U98521 ( .A(n84270), .B(n84271), .Z(n82906) );
  NOR U98522 ( .A(n78506), .B(n78507), .Z(n78513) );
  IV U98523 ( .A(n78507), .Z(n78509) );
  NOR U98524 ( .A(n78509), .B(n78508), .Z(n78510) );
  NOR U98525 ( .A(n78511), .B(n78510), .Z(n78512) );
  NOR U98526 ( .A(n78513), .B(n78512), .Z(n82904) );
  XOR U98527 ( .A(n82906), .B(n82904), .Z(n84279) );
  IV U98528 ( .A(n78514), .Z(n78516) );
  NOR U98529 ( .A(n78516), .B(n78515), .Z(n82902) );
  IV U98530 ( .A(n78517), .Z(n78518) );
  NOR U98531 ( .A(n78519), .B(n78518), .Z(n84277) );
  NOR U98532 ( .A(n82902), .B(n84277), .Z(n78520) );
  XOR U98533 ( .A(n84279), .B(n78520), .Z(n82897) );
  NOR U98534 ( .A(n78522), .B(n78521), .Z(n82899) );
  NOR U98535 ( .A(n78523), .B(n82899), .Z(n78524) );
  XOR U98536 ( .A(n82897), .B(n78524), .Z(n82895) );
  XOR U98537 ( .A(n82894), .B(n82895), .Z(n82890) );
  IV U98538 ( .A(n78525), .Z(n78527) );
  NOR U98539 ( .A(n78527), .B(n78526), .Z(n82889) );
  NOR U98540 ( .A(n82892), .B(n82889), .Z(n78528) );
  XOR U98541 ( .A(n82890), .B(n78528), .Z(n82885) );
  XOR U98542 ( .A(n82886), .B(n82885), .Z(n82880) );
  XOR U98543 ( .A(n82878), .B(n82880), .Z(n82876) );
  XOR U98544 ( .A(n82881), .B(n82876), .Z(n78529) );
  XOR U98545 ( .A(n82875), .B(n78529), .Z(n84287) );
  IV U98546 ( .A(n78530), .Z(n78532) );
  NOR U98547 ( .A(n78532), .B(n78531), .Z(n84285) );
  XOR U98548 ( .A(n84287), .B(n84285), .Z(n84289) );
  IV U98549 ( .A(n78533), .Z(n78534) );
  NOR U98550 ( .A(n78535), .B(n78534), .Z(n84288) );
  NOR U98551 ( .A(n78536), .B(n84282), .Z(n78537) );
  NOR U98552 ( .A(n84288), .B(n78537), .Z(n78538) );
  XOR U98553 ( .A(n84289), .B(n78538), .Z(n78548) );
  IV U98554 ( .A(n78548), .Z(n78540) );
  IV U98555 ( .A(n78553), .Z(n78539) );
  NOR U98556 ( .A(n78540), .B(n78539), .Z(n82874) );
  IV U98557 ( .A(n78541), .Z(n78542) );
  NOR U98558 ( .A(n78542), .B(n78544), .Z(n84299) );
  IV U98559 ( .A(n78543), .Z(n78545) );
  NOR U98560 ( .A(n78545), .B(n78544), .Z(n78549) );
  IV U98561 ( .A(n78549), .Z(n78547) );
  XOR U98562 ( .A(n84288), .B(n84289), .Z(n78546) );
  NOR U98563 ( .A(n78547), .B(n78546), .Z(n88613) );
  NOR U98564 ( .A(n78549), .B(n78548), .Z(n78550) );
  NOR U98565 ( .A(n88613), .B(n78550), .Z(n78551) );
  IV U98566 ( .A(n78551), .Z(n84300) );
  XOR U98567 ( .A(n84299), .B(n84300), .Z(n82872) );
  IV U98568 ( .A(n82872), .Z(n78552) );
  NOR U98569 ( .A(n78553), .B(n78552), .Z(n78554) );
  NOR U98570 ( .A(n82874), .B(n78554), .Z(n82867) );
  XOR U98571 ( .A(n78555), .B(n82867), .Z(n82856) );
  NOR U98572 ( .A(n78556), .B(n82855), .Z(n78557) );
  XOR U98573 ( .A(n82856), .B(n78557), .Z(n84304) );
  IV U98574 ( .A(n84304), .Z(n78571) );
  IV U98575 ( .A(n78558), .Z(n78559) );
  NOR U98576 ( .A(n78559), .B(n78565), .Z(n78560) );
  IV U98577 ( .A(n78560), .Z(n78561) );
  NOR U98578 ( .A(n78562), .B(n78561), .Z(n84303) );
  NOR U98579 ( .A(n78564), .B(n78563), .Z(n78569) );
  NOR U98580 ( .A(n78566), .B(n78565), .Z(n78567) );
  IV U98581 ( .A(n78567), .Z(n78568) );
  NOR U98582 ( .A(n78569), .B(n78568), .Z(n82859) );
  NOR U98583 ( .A(n84303), .B(n82859), .Z(n78570) );
  XOR U98584 ( .A(n78571), .B(n78570), .Z(n82853) );
  XOR U98585 ( .A(n82851), .B(n82853), .Z(n84309) );
  XOR U98586 ( .A(n84307), .B(n84309), .Z(n84311) );
  XOR U98587 ( .A(n84310), .B(n84311), .Z(n82844) );
  XOR U98588 ( .A(n78572), .B(n82844), .Z(n82848) );
  IV U98589 ( .A(n78573), .Z(n78574) );
  NOR U98590 ( .A(n78574), .B(n78581), .Z(n82846) );
  XOR U98591 ( .A(n82848), .B(n82846), .Z(n84318) );
  IV U98592 ( .A(n78575), .Z(n78579) );
  NOR U98593 ( .A(n78577), .B(n78576), .Z(n78578) );
  IV U98594 ( .A(n78578), .Z(n78586) );
  NOR U98595 ( .A(n78579), .B(n78586), .Z(n84316) );
  IV U98596 ( .A(n78580), .Z(n78582) );
  NOR U98597 ( .A(n78582), .B(n78581), .Z(n84314) );
  NOR U98598 ( .A(n84316), .B(n84314), .Z(n78583) );
  XOR U98599 ( .A(n84318), .B(n78583), .Z(n78584) );
  IV U98600 ( .A(n78584), .Z(n84321) );
  IV U98601 ( .A(n78585), .Z(n78587) );
  NOR U98602 ( .A(n78587), .B(n78586), .Z(n84319) );
  XOR U98603 ( .A(n84321), .B(n84319), .Z(n84323) );
  XOR U98604 ( .A(n84322), .B(n84323), .Z(n82842) );
  XOR U98605 ( .A(n78588), .B(n82842), .Z(n82838) );
  XOR U98606 ( .A(n82836), .B(n82838), .Z(n82832) );
  IV U98607 ( .A(n78589), .Z(n78594) );
  NOR U98608 ( .A(n78591), .B(n78590), .Z(n78592) );
  IV U98609 ( .A(n78592), .Z(n78593) );
  NOR U98610 ( .A(n78594), .B(n78593), .Z(n82830) );
  XOR U98611 ( .A(n82832), .B(n82830), .Z(n82834) );
  XOR U98612 ( .A(n82833), .B(n82834), .Z(n82823) );
  XOR U98613 ( .A(n82822), .B(n82823), .Z(n82827) );
  IV U98614 ( .A(n78595), .Z(n78597) );
  NOR U98615 ( .A(n78597), .B(n78596), .Z(n82825) );
  XOR U98616 ( .A(n82827), .B(n82825), .Z(n82818) );
  IV U98617 ( .A(n78598), .Z(n78599) );
  NOR U98618 ( .A(n78600), .B(n78599), .Z(n82820) );
  IV U98619 ( .A(n78601), .Z(n78602) );
  NOR U98620 ( .A(n78603), .B(n78602), .Z(n82817) );
  NOR U98621 ( .A(n82820), .B(n82817), .Z(n78604) );
  XOR U98622 ( .A(n82818), .B(n78604), .Z(n82811) );
  XOR U98623 ( .A(n78605), .B(n82811), .Z(n82809) );
  XOR U98624 ( .A(n78606), .B(n82809), .Z(n82800) );
  XOR U98625 ( .A(n82802), .B(n82800), .Z(n82793) );
  XOR U98626 ( .A(n82792), .B(n82793), .Z(n82797) );
  XOR U98627 ( .A(n82795), .B(n82797), .Z(n82790) );
  XOR U98628 ( .A(n82791), .B(n82790), .Z(n82783) );
  XOR U98629 ( .A(n82785), .B(n82783), .Z(n82780) );
  XOR U98630 ( .A(n82779), .B(n82780), .Z(n82778) );
  XOR U98631 ( .A(n78607), .B(n82778), .Z(n82770) );
  XOR U98632 ( .A(n78608), .B(n82770), .Z(n84332) );
  XOR U98633 ( .A(n84330), .B(n84332), .Z(n84335) );
  NOR U98634 ( .A(n78615), .B(n84335), .Z(n90176) );
  IV U98635 ( .A(n78609), .Z(n78611) );
  NOR U98636 ( .A(n78611), .B(n78610), .Z(n82762) );
  IV U98637 ( .A(n78612), .Z(n78614) );
  NOR U98638 ( .A(n78614), .B(n78613), .Z(n84333) );
  XOR U98639 ( .A(n84335), .B(n84333), .Z(n82763) );
  IV U98640 ( .A(n82763), .Z(n78616) );
  XOR U98641 ( .A(n82762), .B(n78616), .Z(n78618) );
  NOR U98642 ( .A(n78616), .B(n78615), .Z(n78617) );
  NOR U98643 ( .A(n78618), .B(n78617), .Z(n78619) );
  NOR U98644 ( .A(n90176), .B(n78619), .Z(n82766) );
  IV U98645 ( .A(n78620), .Z(n78622) );
  NOR U98646 ( .A(n78622), .B(n78621), .Z(n78623) );
  NOR U98647 ( .A(n78624), .B(n78623), .Z(n84340) );
  IV U98648 ( .A(n84340), .Z(n78625) );
  NOR U98649 ( .A(n82765), .B(n78625), .Z(n78626) );
  XOR U98650 ( .A(n82766), .B(n78626), .Z(n84349) );
  IV U98651 ( .A(n78627), .Z(n78630) );
  IV U98652 ( .A(n78628), .Z(n78629) );
  NOR U98653 ( .A(n78630), .B(n78629), .Z(n84341) );
  XOR U98654 ( .A(n84349), .B(n84341), .Z(n78634) );
  NOR U98655 ( .A(n78631), .B(n78634), .Z(n90208) );
  NOR U98656 ( .A(n84348), .B(n84343), .Z(n78632) );
  NOR U98657 ( .A(n78632), .B(n84350), .Z(n78633) );
  XOR U98658 ( .A(n78634), .B(n78633), .Z(n82760) );
  IV U98659 ( .A(n82760), .Z(n78635) );
  NOR U98660 ( .A(n78636), .B(n78635), .Z(n78637) );
  NOR U98661 ( .A(n90208), .B(n78637), .Z(n82756) );
  IV U98662 ( .A(n78638), .Z(n78639) );
  NOR U98663 ( .A(n78640), .B(n78639), .Z(n82759) );
  IV U98664 ( .A(n78641), .Z(n78643) );
  NOR U98665 ( .A(n78643), .B(n78642), .Z(n82755) );
  NOR U98666 ( .A(n82759), .B(n82755), .Z(n78644) );
  XOR U98667 ( .A(n82756), .B(n78644), .Z(n82753) );
  IV U98668 ( .A(n78645), .Z(n78647) );
  IV U98669 ( .A(n78646), .Z(n78651) );
  NOR U98670 ( .A(n78647), .B(n78651), .Z(n82750) );
  NOR U98671 ( .A(n82750), .B(n78648), .Z(n78649) );
  XOR U98672 ( .A(n82753), .B(n78649), .Z(n84359) );
  IV U98673 ( .A(n78650), .Z(n78652) );
  NOR U98674 ( .A(n78652), .B(n78651), .Z(n82748) );
  IV U98675 ( .A(n78653), .Z(n78655) );
  NOR U98676 ( .A(n78655), .B(n78654), .Z(n84358) );
  NOR U98677 ( .A(n82748), .B(n84358), .Z(n78656) );
  XOR U98678 ( .A(n84359), .B(n78656), .Z(n84357) );
  XOR U98679 ( .A(n84355), .B(n84357), .Z(n82745) );
  XOR U98680 ( .A(n78657), .B(n82745), .Z(n82738) );
  XOR U98681 ( .A(n82739), .B(n82738), .Z(n82742) );
  XOR U98682 ( .A(n82740), .B(n82742), .Z(n84370) );
  XOR U98683 ( .A(n84368), .B(n84370), .Z(n82736) );
  XOR U98684 ( .A(n82734), .B(n82736), .Z(n82733) );
  XOR U98685 ( .A(n82731), .B(n82733), .Z(n84386) );
  XOR U98686 ( .A(n84385), .B(n84386), .Z(n84383) );
  XOR U98687 ( .A(n84382), .B(n84383), .Z(n84403) );
  XOR U98688 ( .A(n78658), .B(n84403), .Z(n84410) );
  IV U98689 ( .A(n84410), .Z(n84414) );
  XOR U98690 ( .A(n78659), .B(n84414), .Z(n82717) );
  XOR U98691 ( .A(n82715), .B(n82717), .Z(n82718) );
  XOR U98692 ( .A(n82719), .B(n82718), .Z(n78660) );
  IV U98693 ( .A(n78660), .Z(n84417) );
  XOR U98694 ( .A(n82711), .B(n84417), .Z(n78661) );
  XOR U98695 ( .A(n78662), .B(n78661), .Z(n82710) );
  XOR U98696 ( .A(n78663), .B(n82710), .Z(n82704) );
  XOR U98697 ( .A(n82703), .B(n82704), .Z(n82695) );
  XOR U98698 ( .A(n82694), .B(n82695), .Z(n82697) );
  XOR U98699 ( .A(n82698), .B(n82697), .Z(n82684) );
  IV U98700 ( .A(n82684), .Z(n82682) );
  XOR U98701 ( .A(n82685), .B(n82682), .Z(n84422) );
  XOR U98702 ( .A(n84421), .B(n84422), .Z(n82680) );
  XOR U98703 ( .A(n82678), .B(n82680), .Z(n84433) );
  XOR U98704 ( .A(n84431), .B(n84433), .Z(n84435) );
  XOR U98705 ( .A(n84434), .B(n84435), .Z(n82676) );
  XOR U98706 ( .A(n82675), .B(n82676), .Z(n84439) );
  XOR U98707 ( .A(n84438), .B(n84439), .Z(n84442) );
  XOR U98708 ( .A(n84441), .B(n84442), .Z(n82672) );
  XOR U98709 ( .A(n82671), .B(n82672), .Z(n82667) );
  XOR U98710 ( .A(n82666), .B(n82667), .Z(n84449) );
  XOR U98711 ( .A(n78664), .B(n84449), .Z(n84455) );
  IV U98712 ( .A(n84455), .Z(n84454) );
  XOR U98713 ( .A(n84456), .B(n84454), .Z(n84452) );
  IV U98714 ( .A(n78665), .Z(n78666) );
  NOR U98715 ( .A(n78667), .B(n78666), .Z(n84451) );
  IV U98716 ( .A(n78668), .Z(n78670) );
  NOR U98717 ( .A(n78670), .B(n78669), .Z(n84457) );
  NOR U98718 ( .A(n84451), .B(n84457), .Z(n78671) );
  XOR U98719 ( .A(n84452), .B(n78671), .Z(n78672) );
  IV U98720 ( .A(n78672), .Z(n82663) );
  XOR U98721 ( .A(n82661), .B(n82663), .Z(n82664) );
  XOR U98722 ( .A(n82665), .B(n82664), .Z(n82653) );
  IV U98723 ( .A(n82653), .Z(n82651) );
  XOR U98724 ( .A(n82650), .B(n82651), .Z(n78679) );
  NOR U98725 ( .A(n78674), .B(n78673), .Z(n82654) );
  IV U98726 ( .A(n78675), .Z(n78677) );
  NOR U98727 ( .A(n78677), .B(n78676), .Z(n82659) );
  NOR U98728 ( .A(n82654), .B(n82659), .Z(n78678) );
  XOR U98729 ( .A(n78679), .B(n78678), .Z(n84463) );
  IV U98730 ( .A(n78680), .Z(n84462) );
  IV U98731 ( .A(n78681), .Z(n78683) );
  NOR U98732 ( .A(n78683), .B(n78682), .Z(n82628) );
  NOR U98733 ( .A(n78684), .B(n82629), .Z(n78685) );
  XOR U98734 ( .A(n82628), .B(n78685), .Z(n78686) );
  XOR U98735 ( .A(n84462), .B(n78686), .Z(n78687) );
  XOR U98736 ( .A(n84463), .B(n78687), .Z(n82639) );
  IV U98737 ( .A(n82639), .Z(n82630) );
  IV U98738 ( .A(n78688), .Z(n78689) );
  NOR U98739 ( .A(n78689), .B(n78694), .Z(n82626) );
  XOR U98740 ( .A(n82630), .B(n82626), .Z(n82634) );
  IV U98741 ( .A(n78690), .Z(n78691) );
  NOR U98742 ( .A(n78692), .B(n78691), .Z(n82637) );
  IV U98743 ( .A(n78693), .Z(n78695) );
  NOR U98744 ( .A(n78695), .B(n78694), .Z(n78696) );
  IV U98745 ( .A(n78696), .Z(n82636) );
  XOR U98746 ( .A(n82637), .B(n82636), .Z(n78697) );
  XOR U98747 ( .A(n82634), .B(n78697), .Z(n84473) );
  XOR U98748 ( .A(n78698), .B(n84473), .Z(n78699) );
  NOR U98749 ( .A(n78700), .B(n78699), .Z(n82625) );
  IV U98750 ( .A(n78700), .Z(n78701) );
  NOR U98751 ( .A(n78701), .B(n84473), .Z(n82623) );
  NOR U98752 ( .A(n82625), .B(n82623), .Z(n82613) );
  IV U98753 ( .A(n78702), .Z(n82621) );
  NOR U98754 ( .A(n78703), .B(n82621), .Z(n78704) );
  IV U98755 ( .A(n78704), .Z(n82615) );
  XOR U98756 ( .A(n82613), .B(n82615), .Z(n82607) );
  XOR U98757 ( .A(n82606), .B(n82607), .Z(n82610) );
  XOR U98758 ( .A(n82609), .B(n82610), .Z(n84480) );
  XOR U98759 ( .A(n84479), .B(n84480), .Z(n84477) );
  XOR U98760 ( .A(n78705), .B(n84477), .Z(n78706) );
  IV U98761 ( .A(n78706), .Z(n82602) );
  XOR U98762 ( .A(n82601), .B(n82602), .Z(n82598) );
  IV U98763 ( .A(n78707), .Z(n78709) );
  NOR U98764 ( .A(n78709), .B(n78708), .Z(n82596) );
  XOR U98765 ( .A(n82598), .B(n82596), .Z(n84492) );
  XOR U98766 ( .A(n84493), .B(n84492), .Z(n82594) );
  IV U98767 ( .A(n78710), .Z(n78711) );
  NOR U98768 ( .A(n78712), .B(n78711), .Z(n84494) );
  NOR U98769 ( .A(n84494), .B(n82593), .Z(n78713) );
  XOR U98770 ( .A(n82594), .B(n78713), .Z(n82586) );
  XOR U98771 ( .A(n82585), .B(n82586), .Z(n82590) );
  XOR U98772 ( .A(n82588), .B(n82590), .Z(n82579) );
  XOR U98773 ( .A(n82577), .B(n82579), .Z(n82581) );
  NOR U98774 ( .A(n78719), .B(n82581), .Z(n88368) );
  IV U98775 ( .A(n78714), .Z(n78715) );
  NOR U98776 ( .A(n78718), .B(n78715), .Z(n82574) );
  IV U98777 ( .A(n78716), .Z(n78717) );
  NOR U98778 ( .A(n78718), .B(n78717), .Z(n82580) );
  XOR U98779 ( .A(n82580), .B(n82581), .Z(n82575) );
  IV U98780 ( .A(n82575), .Z(n78720) );
  XOR U98781 ( .A(n82574), .B(n78720), .Z(n78722) );
  NOR U98782 ( .A(n78720), .B(n78719), .Z(n78721) );
  NOR U98783 ( .A(n78722), .B(n78721), .Z(n78723) );
  NOR U98784 ( .A(n88368), .B(n78723), .Z(n78724) );
  IV U98785 ( .A(n78724), .Z(n82567) );
  XOR U98786 ( .A(n82566), .B(n82567), .Z(n82571) );
  XOR U98787 ( .A(n82569), .B(n82571), .Z(n82564) );
  XOR U98788 ( .A(n82563), .B(n82564), .Z(n78725) );
  NOR U98789 ( .A(n78726), .B(n78725), .Z(n88320) );
  IV U98790 ( .A(n78727), .Z(n78728) );
  NOR U98791 ( .A(n78729), .B(n78728), .Z(n82561) );
  NOR U98792 ( .A(n82563), .B(n82561), .Z(n78730) );
  XOR U98793 ( .A(n78730), .B(n82564), .Z(n78740) );
  NOR U98794 ( .A(n78731), .B(n78740), .Z(n78732) );
  NOR U98795 ( .A(n88320), .B(n78732), .Z(n78743) );
  IV U98796 ( .A(n78743), .Z(n78737) );
  IV U98797 ( .A(n78733), .Z(n78735) );
  NOR U98798 ( .A(n78735), .B(n78734), .Z(n78746) );
  IV U98799 ( .A(n78746), .Z(n78736) );
  NOR U98800 ( .A(n78737), .B(n78736), .Z(n88313) );
  IV U98801 ( .A(n78738), .Z(n78739) );
  NOR U98802 ( .A(n78739), .B(n78755), .Z(n78744) );
  IV U98803 ( .A(n78744), .Z(n78742) );
  IV U98804 ( .A(n78740), .Z(n78741) );
  NOR U98805 ( .A(n78742), .B(n78741), .Z(n88323) );
  NOR U98806 ( .A(n78744), .B(n78743), .Z(n78745) );
  NOR U98807 ( .A(n88323), .B(n78745), .Z(n78756) );
  NOR U98808 ( .A(n78746), .B(n78756), .Z(n78747) );
  NOR U98809 ( .A(n88313), .B(n78747), .Z(n78759) );
  IV U98810 ( .A(n78759), .Z(n78748) );
  NOR U98811 ( .A(n78749), .B(n78748), .Z(n88333) );
  IV U98812 ( .A(n78750), .Z(n78751) );
  NOR U98813 ( .A(n78752), .B(n78751), .Z(n82555) );
  IV U98814 ( .A(n78753), .Z(n78754) );
  NOR U98815 ( .A(n78755), .B(n78754), .Z(n78760) );
  IV U98816 ( .A(n78760), .Z(n78758) );
  IV U98817 ( .A(n78756), .Z(n78757) );
  NOR U98818 ( .A(n78758), .B(n78757), .Z(n82560) );
  NOR U98819 ( .A(n78760), .B(n78759), .Z(n78761) );
  NOR U98820 ( .A(n82560), .B(n78761), .Z(n82556) );
  XOR U98821 ( .A(n82555), .B(n82556), .Z(n78762) );
  NOR U98822 ( .A(n78763), .B(n78762), .Z(n78764) );
  NOR U98823 ( .A(n88333), .B(n78764), .Z(n82549) );
  XOR U98824 ( .A(n78765), .B(n82549), .Z(n82547) );
  IV U98825 ( .A(n78766), .Z(n78768) );
  NOR U98826 ( .A(n78768), .B(n78767), .Z(n82541) );
  IV U98827 ( .A(n78769), .Z(n78770) );
  NOR U98828 ( .A(n78771), .B(n78770), .Z(n82545) );
  NOR U98829 ( .A(n82541), .B(n82545), .Z(n78772) );
  XOR U98830 ( .A(n82547), .B(n78772), .Z(n82539) );
  XOR U98831 ( .A(n82538), .B(n82539), .Z(n78773) );
  XOR U98832 ( .A(n78774), .B(n78773), .Z(n84509) );
  XOR U98833 ( .A(n84507), .B(n84509), .Z(n82529) );
  IV U98834 ( .A(n82529), .Z(n82531) );
  XOR U98835 ( .A(n82530), .B(n82531), .Z(n82526) );
  IV U98836 ( .A(n78775), .Z(n78777) );
  NOR U98837 ( .A(n78777), .B(n78776), .Z(n82533) );
  IV U98838 ( .A(n78778), .Z(n78779) );
  NOR U98839 ( .A(n78780), .B(n78779), .Z(n82524) );
  NOR U98840 ( .A(n82533), .B(n82524), .Z(n78781) );
  XOR U98841 ( .A(n82526), .B(n78781), .Z(n78782) );
  IV U98842 ( .A(n78782), .Z(n82523) );
  IV U98843 ( .A(n78783), .Z(n78788) );
  NOR U98844 ( .A(n78785), .B(n78784), .Z(n78786) );
  IV U98845 ( .A(n78786), .Z(n78787) );
  NOR U98846 ( .A(n78788), .B(n78787), .Z(n82521) );
  XOR U98847 ( .A(n82523), .B(n82521), .Z(n82516) );
  XOR U98848 ( .A(n82515), .B(n82516), .Z(n82519) );
  XOR U98849 ( .A(n82518), .B(n82519), .Z(n82513) );
  XOR U98850 ( .A(n82511), .B(n82513), .Z(n84519) );
  XOR U98851 ( .A(n78789), .B(n84519), .Z(n82503) );
  XOR U98852 ( .A(n82504), .B(n82503), .Z(n84536) );
  IV U98853 ( .A(n78790), .Z(n78797) );
  IV U98854 ( .A(n78791), .Z(n78792) );
  NOR U98855 ( .A(n78797), .B(n78792), .Z(n84534) );
  XOR U98856 ( .A(n84536), .B(n84534), .Z(n84549) );
  IV U98857 ( .A(n78793), .Z(n78794) );
  NOR U98858 ( .A(n78794), .B(n78800), .Z(n84547) );
  IV U98859 ( .A(n78795), .Z(n78796) );
  NOR U98860 ( .A(n78797), .B(n78796), .Z(n84530) );
  NOR U98861 ( .A(n84547), .B(n84530), .Z(n78798) );
  XOR U98862 ( .A(n84549), .B(n78798), .Z(n84544) );
  IV U98863 ( .A(n78799), .Z(n78801) );
  NOR U98864 ( .A(n78801), .B(n78800), .Z(n78802) );
  IV U98865 ( .A(n78802), .Z(n84545) );
  XOR U98866 ( .A(n84544), .B(n84545), .Z(n84553) );
  XOR U98867 ( .A(n84551), .B(n84553), .Z(n84556) );
  IV U98868 ( .A(n78803), .Z(n78804) );
  NOR U98869 ( .A(n78805), .B(n78804), .Z(n82501) );
  IV U98870 ( .A(n78806), .Z(n78807) );
  NOR U98871 ( .A(n78808), .B(n78807), .Z(n84554) );
  NOR U98872 ( .A(n82501), .B(n84554), .Z(n78809) );
  XOR U98873 ( .A(n84556), .B(n78809), .Z(n78810) );
  NOR U98874 ( .A(n78811), .B(n78810), .Z(n78814) );
  IV U98875 ( .A(n78811), .Z(n78813) );
  XOR U98876 ( .A(n84554), .B(n84556), .Z(n78812) );
  NOR U98877 ( .A(n78813), .B(n78812), .Z(n90360) );
  NOR U98878 ( .A(n78814), .B(n90360), .Z(n82497) );
  XOR U98879 ( .A(n78815), .B(n82497), .Z(n84568) );
  XOR U98880 ( .A(n84566), .B(n84568), .Z(n84570) );
  XOR U98881 ( .A(n84569), .B(n84570), .Z(n90393) );
  XOR U98882 ( .A(n84573), .B(n90393), .Z(n78822) );
  IV U98883 ( .A(n78822), .Z(n84574) );
  NOR U98884 ( .A(n78823), .B(n84574), .Z(n90429) );
  IV U98885 ( .A(n78816), .Z(n78818) );
  NOR U98886 ( .A(n78818), .B(n78817), .Z(n82487) );
  IV U98887 ( .A(n78819), .Z(n78820) );
  NOR U98888 ( .A(n90423), .B(n78820), .Z(n78821) );
  IV U98889 ( .A(n78821), .Z(n84575) );
  XOR U98890 ( .A(n84575), .B(n78822), .Z(n82488) );
  IV U98891 ( .A(n82488), .Z(n78824) );
  XOR U98892 ( .A(n82487), .B(n78824), .Z(n78826) );
  NOR U98893 ( .A(n78824), .B(n78823), .Z(n78825) );
  NOR U98894 ( .A(n78826), .B(n78825), .Z(n78827) );
  NOR U98895 ( .A(n90429), .B(n78827), .Z(n82490) );
  IV U98896 ( .A(n78828), .Z(n78832) );
  XOR U98897 ( .A(n78830), .B(n78829), .Z(n78831) );
  NOR U98898 ( .A(n78832), .B(n78831), .Z(n82491) );
  XOR U98899 ( .A(n82490), .B(n82491), .Z(n82481) );
  XOR U98900 ( .A(n82479), .B(n82481), .Z(n82477) );
  XOR U98901 ( .A(n78833), .B(n82477), .Z(n82459) );
  XOR U98902 ( .A(n82469), .B(n82459), .Z(n82467) );
  XOR U98903 ( .A(n82466), .B(n82467), .Z(n84582) );
  NOR U98904 ( .A(n78834), .B(n82460), .Z(n78838) );
  IV U98905 ( .A(n78835), .Z(n78837) );
  IV U98906 ( .A(n78836), .Z(n78843) );
  NOR U98907 ( .A(n78837), .B(n78843), .Z(n84581) );
  NOR U98908 ( .A(n78838), .B(n84581), .Z(n78839) );
  XOR U98909 ( .A(n84582), .B(n78839), .Z(n84584) );
  NOR U98910 ( .A(n78841), .B(n78840), .Z(n84586) );
  IV U98911 ( .A(n78842), .Z(n78844) );
  NOR U98912 ( .A(n78844), .B(n78843), .Z(n84591) );
  NOR U98913 ( .A(n84586), .B(n84591), .Z(n78845) );
  XOR U98914 ( .A(n84584), .B(n78845), .Z(n82456) );
  IV U98915 ( .A(n78846), .Z(n78847) );
  NOR U98916 ( .A(n78848), .B(n78847), .Z(n84590) );
  IV U98917 ( .A(n78849), .Z(n78850) );
  NOR U98918 ( .A(n78850), .B(n78854), .Z(n82455) );
  NOR U98919 ( .A(n84590), .B(n82455), .Z(n78851) );
  XOR U98920 ( .A(n82456), .B(n78851), .Z(n78861) );
  IV U98921 ( .A(n78861), .Z(n82453) );
  IV U98922 ( .A(n78852), .Z(n78853) );
  NOR U98923 ( .A(n78854), .B(n78853), .Z(n82451) );
  XOR U98924 ( .A(n82453), .B(n82451), .Z(n78855) );
  NOR U98925 ( .A(n78856), .B(n78855), .Z(n90482) );
  IV U98926 ( .A(n78857), .Z(n78858) );
  NOR U98927 ( .A(n78859), .B(n78858), .Z(n82449) );
  NOR U98928 ( .A(n82449), .B(n82451), .Z(n78860) );
  XOR U98929 ( .A(n78861), .B(n78860), .Z(n78872) );
  IV U98930 ( .A(n78872), .Z(n78862) );
  NOR U98931 ( .A(n78863), .B(n78862), .Z(n78864) );
  NOR U98932 ( .A(n90482), .B(n78864), .Z(n78874) );
  IV U98933 ( .A(n78874), .Z(n78868) );
  IV U98934 ( .A(n78865), .Z(n78866) );
  NOR U98935 ( .A(n78882), .B(n78866), .Z(n78878) );
  IV U98936 ( .A(n78878), .Z(n78867) );
  NOR U98937 ( .A(n78868), .B(n78867), .Z(n88251) );
  IV U98938 ( .A(n78869), .Z(n78870) );
  NOR U98939 ( .A(n78871), .B(n78870), .Z(n78875) );
  IV U98940 ( .A(n78875), .Z(n78873) );
  NOR U98941 ( .A(n78873), .B(n78872), .Z(n82448) );
  NOR U98942 ( .A(n78875), .B(n78874), .Z(n78876) );
  NOR U98943 ( .A(n82448), .B(n78876), .Z(n78877) );
  NOR U98944 ( .A(n78878), .B(n78877), .Z(n78879) );
  NOR U98945 ( .A(n88251), .B(n78879), .Z(n84600) );
  IV U98946 ( .A(n78880), .Z(n78881) );
  NOR U98947 ( .A(n78882), .B(n78881), .Z(n78883) );
  IV U98948 ( .A(n78883), .Z(n84601) );
  XOR U98949 ( .A(n84600), .B(n84601), .Z(n82446) );
  XOR U98950 ( .A(n82445), .B(n82446), .Z(n84607) );
  XOR U98951 ( .A(n84605), .B(n84607), .Z(n84610) );
  XOR U98952 ( .A(n84608), .B(n84610), .Z(n82444) );
  XOR U98953 ( .A(n82442), .B(n82444), .Z(n78884) );
  NOR U98954 ( .A(n78885), .B(n78884), .Z(n78886) );
  NOR U98955 ( .A(n78892), .B(n78886), .Z(n82429) );
  IV U98956 ( .A(n82429), .Z(n78891) );
  IV U98957 ( .A(n78887), .Z(n82438) );
  NOR U98958 ( .A(n78888), .B(n82438), .Z(n82432) );
  NOR U98959 ( .A(n82432), .B(n82442), .Z(n78889) );
  XOR U98960 ( .A(n78889), .B(n82444), .Z(n78894) );
  NOR U98961 ( .A(n78890), .B(n78894), .Z(n82430) );
  NOR U98962 ( .A(n78891), .B(n82430), .Z(n78896) );
  IV U98963 ( .A(n78892), .Z(n78893) );
  NOR U98964 ( .A(n78894), .B(n78893), .Z(n78895) );
  NOR U98965 ( .A(n78896), .B(n78895), .Z(n82423) );
  IV U98966 ( .A(n78897), .Z(n82422) );
  NOR U98967 ( .A(n78898), .B(n82422), .Z(n78902) );
  IV U98968 ( .A(n78899), .Z(n78900) );
  NOR U98969 ( .A(n78901), .B(n78900), .Z(n82419) );
  NOR U98970 ( .A(n78902), .B(n82419), .Z(n78903) );
  XOR U98971 ( .A(n82423), .B(n78903), .Z(n82414) );
  IV U98972 ( .A(n78904), .Z(n78905) );
  NOR U98973 ( .A(n78906), .B(n78905), .Z(n82416) );
  IV U98974 ( .A(n78907), .Z(n78909) );
  NOR U98975 ( .A(n78909), .B(n78908), .Z(n82413) );
  NOR U98976 ( .A(n82416), .B(n82413), .Z(n78910) );
  XOR U98977 ( .A(n82414), .B(n78910), .Z(n84620) );
  IV U98978 ( .A(n78911), .Z(n78913) );
  IV U98979 ( .A(n78912), .Z(n78924) );
  NOR U98980 ( .A(n78913), .B(n78924), .Z(n78914) );
  IV U98981 ( .A(n78914), .Z(n78918) );
  NOR U98982 ( .A(n84620), .B(n78918), .Z(n88227) );
  IV U98983 ( .A(n78915), .Z(n78917) );
  NOR U98984 ( .A(n78917), .B(n78916), .Z(n84618) );
  XOR U98985 ( .A(n84618), .B(n84620), .Z(n84616) );
  IV U98986 ( .A(n84616), .Z(n78919) );
  XOR U98987 ( .A(n84615), .B(n78919), .Z(n78921) );
  NOR U98988 ( .A(n78919), .B(n78918), .Z(n78920) );
  NOR U98989 ( .A(n78921), .B(n78920), .Z(n78922) );
  NOR U98990 ( .A(n88227), .B(n78922), .Z(n84630) );
  IV U98991 ( .A(n78923), .Z(n78925) );
  NOR U98992 ( .A(n78925), .B(n78924), .Z(n78926) );
  IV U98993 ( .A(n78926), .Z(n84631) );
  XOR U98994 ( .A(n84630), .B(n84631), .Z(n84637) );
  XOR U98995 ( .A(n84636), .B(n84637), .Z(n82411) );
  XOR U98996 ( .A(n82410), .B(n82411), .Z(n82406) );
  XOR U98997 ( .A(n78927), .B(n82406), .Z(n78935) );
  IV U98998 ( .A(n78928), .Z(n78929) );
  NOR U98999 ( .A(n78930), .B(n78929), .Z(n82402) );
  IV U99000 ( .A(n78931), .Z(n78933) );
  NOR U99001 ( .A(n78933), .B(n78932), .Z(n82405) );
  NOR U99002 ( .A(n82402), .B(n82405), .Z(n78934) );
  XOR U99003 ( .A(n78935), .B(n78934), .Z(n84649) );
  IV U99004 ( .A(n78936), .Z(n78938) );
  NOR U99005 ( .A(n78938), .B(n78937), .Z(n84647) );
  XOR U99006 ( .A(n84649), .B(n84647), .Z(n84651) );
  XOR U99007 ( .A(n84650), .B(n84651), .Z(n78939) );
  NOR U99008 ( .A(n78940), .B(n78939), .Z(n84664) );
  IV U99009 ( .A(n78941), .Z(n78942) );
  NOR U99010 ( .A(n78943), .B(n78942), .Z(n82398) );
  NOR U99011 ( .A(n84650), .B(n82398), .Z(n78944) );
  XOR U99012 ( .A(n78944), .B(n84651), .Z(n84655) );
  NOR U99013 ( .A(n78945), .B(n84655), .Z(n78946) );
  NOR U99014 ( .A(n84664), .B(n78946), .Z(n82394) );
  XOR U99015 ( .A(n78947), .B(n82394), .Z(n82388) );
  IV U99016 ( .A(n78948), .Z(n78950) );
  NOR U99017 ( .A(n78950), .B(n78949), .Z(n82391) );
  IV U99018 ( .A(n78951), .Z(n78952) );
  NOR U99019 ( .A(n78953), .B(n78952), .Z(n82387) );
  NOR U99020 ( .A(n82391), .B(n82387), .Z(n78954) );
  XOR U99021 ( .A(n82388), .B(n78954), .Z(n82382) );
  XOR U99022 ( .A(n82385), .B(n82382), .Z(n82380) );
  XOR U99023 ( .A(n78955), .B(n82380), .Z(n78956) );
  IV U99024 ( .A(n78956), .Z(n84670) );
  XOR U99025 ( .A(n84668), .B(n84670), .Z(n82376) );
  XOR U99026 ( .A(n82373), .B(n82376), .Z(n82372) );
  IV U99027 ( .A(n78957), .Z(n78960) );
  IV U99028 ( .A(n78958), .Z(n78959) );
  NOR U99029 ( .A(n78960), .B(n78959), .Z(n82370) );
  NOR U99030 ( .A(n82375), .B(n82370), .Z(n78961) );
  XOR U99031 ( .A(n82372), .B(n78961), .Z(n82367) );
  IV U99032 ( .A(n78962), .Z(n78965) );
  IV U99033 ( .A(n78963), .Z(n78964) );
  NOR U99034 ( .A(n78965), .B(n78964), .Z(n78966) );
  IV U99035 ( .A(n78966), .Z(n82368) );
  XOR U99036 ( .A(n82367), .B(n82368), .Z(n84685) );
  XOR U99037 ( .A(n82360), .B(n84685), .Z(n82364) );
  XOR U99038 ( .A(n82362), .B(n82364), .Z(n82358) );
  XOR U99039 ( .A(n78967), .B(n82358), .Z(n78968) );
  IV U99040 ( .A(n78968), .Z(n84689) );
  XOR U99041 ( .A(n84687), .B(n84689), .Z(n84691) );
  XOR U99042 ( .A(n84690), .B(n84691), .Z(n82344) );
  XOR U99043 ( .A(n82343), .B(n82344), .Z(n82347) );
  XOR U99044 ( .A(n82346), .B(n82347), .Z(n82350) );
  XOR U99045 ( .A(n82349), .B(n82350), .Z(n84697) );
  XOR U99046 ( .A(n84696), .B(n84697), .Z(n84700) );
  IV U99047 ( .A(n78969), .Z(n78970) );
  NOR U99048 ( .A(n78971), .B(n78970), .Z(n84695) );
  IV U99049 ( .A(n78972), .Z(n78973) );
  NOR U99050 ( .A(n78976), .B(n78973), .Z(n84699) );
  NOR U99051 ( .A(n84695), .B(n84699), .Z(n78974) );
  XOR U99052 ( .A(n84700), .B(n78974), .Z(n84702) );
  IV U99053 ( .A(n78975), .Z(n78977) );
  NOR U99054 ( .A(n78977), .B(n78976), .Z(n78978) );
  IV U99055 ( .A(n78978), .Z(n84703) );
  XOR U99056 ( .A(n84702), .B(n84703), .Z(n84705) );
  XOR U99057 ( .A(n84706), .B(n84705), .Z(n82337) );
  XOR U99058 ( .A(n82334), .B(n82337), .Z(n82332) );
  IV U99059 ( .A(n78979), .Z(n78981) );
  NOR U99060 ( .A(n78981), .B(n78980), .Z(n82338) );
  IV U99061 ( .A(n78982), .Z(n78984) );
  NOR U99062 ( .A(n78984), .B(n78983), .Z(n78985) );
  IV U99063 ( .A(n78985), .Z(n82331) );
  XOR U99064 ( .A(n82338), .B(n82331), .Z(n78986) );
  XOR U99065 ( .A(n82332), .B(n78986), .Z(n82329) );
  XOR U99066 ( .A(n78987), .B(n82329), .Z(n84713) );
  IV U99067 ( .A(n78988), .Z(n78989) );
  NOR U99068 ( .A(n78991), .B(n78989), .Z(n84712) );
  IV U99069 ( .A(n78990), .Z(n78992) );
  NOR U99070 ( .A(n78992), .B(n78991), .Z(n78993) );
  IV U99071 ( .A(n78993), .Z(n82328) );
  XOR U99072 ( .A(n84712), .B(n82328), .Z(n78994) );
  XOR U99073 ( .A(n84713), .B(n78994), .Z(n78995) );
  IV U99074 ( .A(n78995), .Z(n84722) );
  IV U99075 ( .A(n78996), .Z(n78997) );
  NOR U99076 ( .A(n78998), .B(n78997), .Z(n84721) );
  NOR U99077 ( .A(n82323), .B(n84721), .Z(n78999) );
  XOR U99078 ( .A(n84722), .B(n78999), .Z(n82314) );
  IV U99079 ( .A(n79000), .Z(n79002) );
  NOR U99080 ( .A(n79002), .B(n79001), .Z(n84718) );
  IV U99081 ( .A(n79003), .Z(n79005) );
  NOR U99082 ( .A(n79005), .B(n79004), .Z(n82315) );
  NOR U99083 ( .A(n84718), .B(n82315), .Z(n79006) );
  XOR U99084 ( .A(n82314), .B(n79006), .Z(n88113) );
  XOR U99085 ( .A(n82309), .B(n88113), .Z(n82307) );
  XOR U99086 ( .A(n82308), .B(n82307), .Z(n84726) );
  XOR U99087 ( .A(n84728), .B(n84726), .Z(n84730) );
  XOR U99088 ( .A(n84729), .B(n84730), .Z(n84734) );
  XOR U99089 ( .A(n84733), .B(n84734), .Z(n84741) );
  XOR U99090 ( .A(n84736), .B(n84741), .Z(n84744) );
  NOR U99091 ( .A(n79007), .B(n84744), .Z(n84747) );
  XOR U99092 ( .A(n79008), .B(n84744), .Z(n82304) );
  IV U99093 ( .A(n82304), .Z(n79010) );
  NOR U99094 ( .A(n79010), .B(n79009), .Z(n79011) );
  NOR U99095 ( .A(n84747), .B(n79011), .Z(n79012) );
  IV U99096 ( .A(n79012), .Z(n84750) );
  IV U99097 ( .A(n79013), .Z(n79014) );
  NOR U99098 ( .A(n79015), .B(n79014), .Z(n84749) );
  XOR U99099 ( .A(n84750), .B(n84749), .Z(n84762) );
  XOR U99100 ( .A(n79016), .B(n84762), .Z(n84766) );
  XOR U99101 ( .A(n79017), .B(n84766), .Z(n84768) );
  XOR U99102 ( .A(n84769), .B(n84768), .Z(n84785) );
  XOR U99103 ( .A(n79018), .B(n84785), .Z(n84782) );
  XOR U99104 ( .A(n84780), .B(n84782), .Z(n84793) );
  XOR U99105 ( .A(n84792), .B(n84793), .Z(n79019) );
  XOR U99106 ( .A(n82300), .B(n79019), .Z(n82297) );
  XOR U99107 ( .A(n82296), .B(n82297), .Z(n82289) );
  XOR U99108 ( .A(n82288), .B(n82289), .Z(n82293) );
  IV U99109 ( .A(n79020), .Z(n79025) );
  NOR U99110 ( .A(n79022), .B(n79021), .Z(n79023) );
  IV U99111 ( .A(n79023), .Z(n79024) );
  NOR U99112 ( .A(n79025), .B(n79024), .Z(n82291) );
  XOR U99113 ( .A(n82293), .B(n82291), .Z(n84797) );
  XOR U99114 ( .A(n84796), .B(n84797), .Z(n84800) );
  XOR U99115 ( .A(n84799), .B(n84800), .Z(n82281) );
  XOR U99116 ( .A(n82280), .B(n82281), .Z(n82285) );
  IV U99117 ( .A(n79026), .Z(n79028) );
  NOR U99118 ( .A(n79028), .B(n79027), .Z(n82283) );
  XOR U99119 ( .A(n82285), .B(n82283), .Z(n84807) );
  IV U99120 ( .A(n79029), .Z(n79032) );
  IV U99121 ( .A(n79030), .Z(n79031) );
  NOR U99122 ( .A(n79032), .B(n79031), .Z(n84805) );
  XOR U99123 ( .A(n84807), .B(n84805), .Z(n84814) );
  IV U99124 ( .A(n79033), .Z(n79034) );
  NOR U99125 ( .A(n79035), .B(n79034), .Z(n84809) );
  IV U99126 ( .A(n79036), .Z(n79037) );
  NOR U99127 ( .A(n79037), .B(n79041), .Z(n84812) );
  NOR U99128 ( .A(n84809), .B(n84812), .Z(n79038) );
  XOR U99129 ( .A(n84814), .B(n79038), .Z(n79039) );
  IV U99130 ( .A(n79039), .Z(n82275) );
  IV U99131 ( .A(n79040), .Z(n79042) );
  NOR U99132 ( .A(n79042), .B(n79041), .Z(n82273) );
  XOR U99133 ( .A(n82275), .B(n82273), .Z(n82276) );
  XOR U99134 ( .A(n82277), .B(n82276), .Z(n79048) );
  IV U99135 ( .A(n79048), .Z(n82270) );
  XOR U99136 ( .A(n82269), .B(n82270), .Z(n79043) );
  NOR U99137 ( .A(n79044), .B(n79043), .Z(n90704) );
  IV U99138 ( .A(n79045), .Z(n79047) );
  NOR U99139 ( .A(n79047), .B(n79046), .Z(n82263) );
  NOR U99140 ( .A(n82269), .B(n82263), .Z(n79049) );
  XOR U99141 ( .A(n79049), .B(n79048), .Z(n82266) );
  IV U99142 ( .A(n79050), .Z(n79052) );
  NOR U99143 ( .A(n79052), .B(n79051), .Z(n79053) );
  IV U99144 ( .A(n79053), .Z(n82265) );
  XOR U99145 ( .A(n82266), .B(n82265), .Z(n79054) );
  NOR U99146 ( .A(n79055), .B(n79054), .Z(n79056) );
  NOR U99147 ( .A(n90704), .B(n79056), .Z(n79057) );
  IV U99148 ( .A(n79057), .Z(n84823) );
  XOR U99149 ( .A(n84817), .B(n84823), .Z(n82261) );
  XOR U99150 ( .A(n79058), .B(n82261), .Z(n82258) );
  XOR U99151 ( .A(n79059), .B(n82258), .Z(n82247) );
  XOR U99152 ( .A(n79060), .B(n82247), .Z(n82251) );
  XOR U99153 ( .A(n79061), .B(n82251), .Z(n82242) );
  NOR U99154 ( .A(n79063), .B(n79062), .Z(n79065) );
  NOR U99155 ( .A(n79065), .B(n79064), .Z(n82240) );
  XOR U99156 ( .A(n82242), .B(n82240), .Z(n84841) );
  XOR U99157 ( .A(n82238), .B(n84841), .Z(n84847) );
  IV U99158 ( .A(n79066), .Z(n79067) );
  NOR U99159 ( .A(n79068), .B(n79067), .Z(n84840) );
  IV U99160 ( .A(n79069), .Z(n79070) );
  NOR U99161 ( .A(n79070), .B(n79073), .Z(n84846) );
  NOR U99162 ( .A(n84840), .B(n84846), .Z(n79071) );
  XOR U99163 ( .A(n84847), .B(n79071), .Z(n84849) );
  IV U99164 ( .A(n79072), .Z(n79074) );
  NOR U99165 ( .A(n79074), .B(n79073), .Z(n79075) );
  IV U99166 ( .A(n79075), .Z(n84850) );
  XOR U99167 ( .A(n84849), .B(n84850), .Z(n84853) );
  XOR U99168 ( .A(n84852), .B(n84853), .Z(n82235) );
  IV U99169 ( .A(n79076), .Z(n79077) );
  NOR U99170 ( .A(n79078), .B(n79077), .Z(n82234) );
  IV U99171 ( .A(n79079), .Z(n79080) );
  NOR U99172 ( .A(n79081), .B(n79080), .Z(n82232) );
  NOR U99173 ( .A(n82234), .B(n82232), .Z(n79082) );
  XOR U99174 ( .A(n82235), .B(n79082), .Z(n79083) );
  NOR U99175 ( .A(n79084), .B(n79083), .Z(n82229) );
  IV U99176 ( .A(n79084), .Z(n79086) );
  XOR U99177 ( .A(n82234), .B(n82235), .Z(n79085) );
  NOR U99178 ( .A(n79086), .B(n79085), .Z(n82231) );
  NOR U99179 ( .A(n82229), .B(n82231), .Z(n82224) );
  IV U99180 ( .A(n79087), .Z(n79088) );
  NOR U99181 ( .A(n79089), .B(n79088), .Z(n82227) );
  IV U99182 ( .A(n79090), .Z(n79091) );
  NOR U99183 ( .A(n79094), .B(n79091), .Z(n82223) );
  NOR U99184 ( .A(n82227), .B(n82223), .Z(n79092) );
  XOR U99185 ( .A(n82224), .B(n79092), .Z(n84859) );
  IV U99186 ( .A(n79093), .Z(n79095) );
  NOR U99187 ( .A(n79095), .B(n79094), .Z(n84857) );
  IV U99188 ( .A(n79096), .Z(n79098) );
  NOR U99189 ( .A(n79098), .B(n79097), .Z(n82221) );
  NOR U99190 ( .A(n84857), .B(n82221), .Z(n79099) );
  XOR U99191 ( .A(n84859), .B(n79099), .Z(n79100) );
  IV U99192 ( .A(n79100), .Z(n84886) );
  IV U99193 ( .A(n79101), .Z(n79103) );
  NOR U99194 ( .A(n79103), .B(n79102), .Z(n84871) );
  IV U99195 ( .A(n79104), .Z(n79105) );
  NOR U99196 ( .A(n79105), .B(n84889), .Z(n84885) );
  NOR U99197 ( .A(n84871), .B(n84885), .Z(n79106) );
  XOR U99198 ( .A(n84886), .B(n79106), .Z(n82214) );
  IV U99199 ( .A(n79107), .Z(n79109) );
  NOR U99200 ( .A(n79109), .B(n79108), .Z(n82217) );
  NOR U99201 ( .A(n82217), .B(n82215), .Z(n79110) );
  IV U99202 ( .A(n79110), .Z(n79111) );
  NOR U99203 ( .A(n79112), .B(n79111), .Z(n79113) );
  XOR U99204 ( .A(n82214), .B(n79113), .Z(n84901) );
  XOR U99205 ( .A(n84900), .B(n84901), .Z(n84904) );
  IV U99206 ( .A(n84904), .Z(n79119) );
  IV U99207 ( .A(n79114), .Z(n79121) );
  NOR U99208 ( .A(n79115), .B(n79121), .Z(n84899) );
  IV U99209 ( .A(n79116), .Z(n79117) );
  NOR U99210 ( .A(n79117), .B(n79121), .Z(n84903) );
  NOR U99211 ( .A(n84899), .B(n84903), .Z(n79118) );
  XOR U99212 ( .A(n79119), .B(n79118), .Z(n82208) );
  IV U99213 ( .A(n79120), .Z(n79122) );
  NOR U99214 ( .A(n79122), .B(n79121), .Z(n82206) );
  XOR U99215 ( .A(n82208), .B(n82206), .Z(n82210) );
  XOR U99216 ( .A(n82209), .B(n82210), .Z(n82202) );
  XOR U99217 ( .A(n79123), .B(n82202), .Z(n79124) );
  IV U99218 ( .A(n79124), .Z(n84910) );
  IV U99219 ( .A(n79125), .Z(n79126) );
  NOR U99220 ( .A(n79127), .B(n79126), .Z(n84908) );
  NOR U99221 ( .A(n79128), .B(n82195), .Z(n79129) );
  NOR U99222 ( .A(n84908), .B(n79129), .Z(n79130) );
  XOR U99223 ( .A(n84910), .B(n79130), .Z(n82185) );
  IV U99224 ( .A(n79131), .Z(n82191) );
  NOR U99225 ( .A(n79132), .B(n82191), .Z(n79135) );
  NOR U99226 ( .A(n79133), .B(n82186), .Z(n79134) );
  NOR U99227 ( .A(n79135), .B(n79134), .Z(n79136) );
  XOR U99228 ( .A(n82185), .B(n79136), .Z(n84947) );
  XOR U99229 ( .A(n84945), .B(n84947), .Z(n84965) );
  IV U99230 ( .A(n79137), .Z(n79138) );
  NOR U99231 ( .A(n79138), .B(n79145), .Z(n84963) );
  XOR U99232 ( .A(n84965), .B(n84963), .Z(n84962) );
  IV U99233 ( .A(n79139), .Z(n79143) );
  NOR U99234 ( .A(n79141), .B(n79140), .Z(n79142) );
  IV U99235 ( .A(n79142), .Z(n79149) );
  NOR U99236 ( .A(n79143), .B(n79149), .Z(n84960) );
  IV U99237 ( .A(n79144), .Z(n79146) );
  NOR U99238 ( .A(n79146), .B(n79145), .Z(n82182) );
  NOR U99239 ( .A(n84960), .B(n82182), .Z(n79147) );
  XOR U99240 ( .A(n84962), .B(n79147), .Z(n82174) );
  IV U99241 ( .A(n79148), .Z(n79150) );
  NOR U99242 ( .A(n79150), .B(n79149), .Z(n79151) );
  IV U99243 ( .A(n79151), .Z(n82175) );
  XOR U99244 ( .A(n82174), .B(n82175), .Z(n82179) );
  XOR U99245 ( .A(n82177), .B(n82179), .Z(n84974) );
  XOR U99246 ( .A(n84973), .B(n84974), .Z(n84978) );
  XOR U99247 ( .A(n84976), .B(n84978), .Z(n82172) );
  XOR U99248 ( .A(n82171), .B(n82172), .Z(n84984) );
  XOR U99249 ( .A(n84983), .B(n84984), .Z(n82169) );
  XOR U99250 ( .A(n82168), .B(n82169), .Z(n79156) );
  IV U99251 ( .A(n79152), .Z(n79154) );
  NOR U99252 ( .A(n79154), .B(n79153), .Z(n79161) );
  IV U99253 ( .A(n79161), .Z(n79155) );
  NOR U99254 ( .A(n79156), .B(n79155), .Z(n90725) );
  IV U99255 ( .A(n79157), .Z(n79159) );
  NOR U99256 ( .A(n79159), .B(n79158), .Z(n82166) );
  NOR U99257 ( .A(n82168), .B(n82166), .Z(n79160) );
  XOR U99258 ( .A(n79160), .B(n82169), .Z(n84992) );
  NOR U99259 ( .A(n79161), .B(n84992), .Z(n79162) );
  NOR U99260 ( .A(n90725), .B(n79162), .Z(n82163) );
  XOR U99261 ( .A(n79163), .B(n82163), .Z(n84997) );
  XOR U99262 ( .A(n84995), .B(n84997), .Z(n85002) );
  IV U99263 ( .A(n79164), .Z(n79166) );
  IV U99264 ( .A(n79165), .Z(n79172) );
  NOR U99265 ( .A(n79166), .B(n79172), .Z(n85001) );
  IV U99266 ( .A(n79167), .Z(n79169) );
  NOR U99267 ( .A(n79169), .B(n79168), .Z(n84998) );
  XOR U99268 ( .A(n85001), .B(n84998), .Z(n79170) );
  XOR U99269 ( .A(n85002), .B(n79170), .Z(n85009) );
  IV U99270 ( .A(n79171), .Z(n79173) );
  NOR U99271 ( .A(n79173), .B(n79172), .Z(n79178) );
  IV U99272 ( .A(n79174), .Z(n79175) );
  NOR U99273 ( .A(n79176), .B(n79175), .Z(n79177) );
  NOR U99274 ( .A(n79178), .B(n79177), .Z(n85010) );
  XOR U99275 ( .A(n85009), .B(n85010), .Z(n79185) );
  IV U99276 ( .A(n79185), .Z(n82158) );
  XOR U99277 ( .A(n79184), .B(n82158), .Z(n79179) );
  NOR U99278 ( .A(n79180), .B(n79179), .Z(n87909) );
  IV U99279 ( .A(n79181), .Z(n79183) );
  IV U99280 ( .A(n79182), .Z(n79189) );
  NOR U99281 ( .A(n79183), .B(n79189), .Z(n82151) );
  NOR U99282 ( .A(n79184), .B(n82151), .Z(n79186) );
  XOR U99283 ( .A(n79186), .B(n79185), .Z(n82154) );
  IV U99284 ( .A(n79187), .Z(n79188) );
  NOR U99285 ( .A(n79189), .B(n79188), .Z(n79190) );
  IV U99286 ( .A(n79190), .Z(n82153) );
  XOR U99287 ( .A(n82154), .B(n82153), .Z(n79191) );
  NOR U99288 ( .A(n79192), .B(n79191), .Z(n79193) );
  NOR U99289 ( .A(n87909), .B(n79193), .Z(n85020) );
  IV U99290 ( .A(n79194), .Z(n79195) );
  NOR U99291 ( .A(n79196), .B(n79195), .Z(n85019) );
  IV U99292 ( .A(n85019), .Z(n85022) );
  XOR U99293 ( .A(n85024), .B(n85022), .Z(n79197) );
  XOR U99294 ( .A(n85020), .B(n79197), .Z(n85031) );
  IV U99295 ( .A(n79198), .Z(n79199) );
  NOR U99296 ( .A(n79200), .B(n79199), .Z(n79201) );
  IV U99297 ( .A(n79201), .Z(n82150) );
  XOR U99298 ( .A(n85031), .B(n82150), .Z(n79202) );
  XOR U99299 ( .A(n79203), .B(n79202), .Z(n82149) );
  IV U99300 ( .A(n79204), .Z(n79205) );
  NOR U99301 ( .A(n79206), .B(n79205), .Z(n82147) );
  XOR U99302 ( .A(n82149), .B(n82147), .Z(n85034) );
  XOR U99303 ( .A(n85033), .B(n85034), .Z(n79211) );
  IV U99304 ( .A(n79211), .Z(n82144) );
  NOR U99305 ( .A(n79210), .B(n82144), .Z(n90748) );
  IV U99306 ( .A(n79207), .Z(n79209) );
  NOR U99307 ( .A(n79209), .B(n79208), .Z(n82143) );
  XOR U99308 ( .A(n82143), .B(n79211), .Z(n79213) );
  NOR U99309 ( .A(n79211), .B(n79210), .Z(n79212) );
  NOR U99310 ( .A(n79213), .B(n79212), .Z(n85047) );
  NOR U99311 ( .A(n90748), .B(n85047), .Z(n85054) );
  XOR U99312 ( .A(n90746), .B(n85054), .Z(n85052) );
  XOR U99313 ( .A(n85051), .B(n85052), .Z(n82141) );
  XOR U99314 ( .A(n79214), .B(n82141), .Z(n79215) );
  IV U99315 ( .A(n79215), .Z(n85061) );
  XOR U99316 ( .A(n85059), .B(n85061), .Z(n82135) );
  IV U99317 ( .A(n79216), .Z(n79218) );
  NOR U99318 ( .A(n79218), .B(n79217), .Z(n82133) );
  XOR U99319 ( .A(n82135), .B(n82133), .Z(n85072) );
  IV U99320 ( .A(n85072), .Z(n85074) );
  IV U99321 ( .A(n79219), .Z(n79220) );
  NOR U99322 ( .A(n79221), .B(n79220), .Z(n85073) );
  IV U99323 ( .A(n85073), .Z(n85071) );
  XOR U99324 ( .A(n85074), .B(n85071), .Z(n82131) );
  IV U99325 ( .A(n79222), .Z(n79223) );
  NOR U99326 ( .A(n79224), .B(n79223), .Z(n85075) );
  IV U99327 ( .A(n79225), .Z(n79227) );
  NOR U99328 ( .A(n79227), .B(n79226), .Z(n82130) );
  NOR U99329 ( .A(n85075), .B(n82130), .Z(n79228) );
  XOR U99330 ( .A(n82131), .B(n79228), .Z(n79229) );
  IV U99331 ( .A(n79229), .Z(n85082) );
  XOR U99332 ( .A(n85080), .B(n85082), .Z(n85084) );
  XOR U99333 ( .A(n85083), .B(n85084), .Z(n82128) );
  XOR U99334 ( .A(n82129), .B(n82128), .Z(n79233) );
  IV U99335 ( .A(n79233), .Z(n79230) );
  NOR U99336 ( .A(n79231), .B(n79230), .Z(n87846) );
  IV U99337 ( .A(n79234), .Z(n79232) );
  NOR U99338 ( .A(n79232), .B(n85084), .Z(n87824) );
  NOR U99339 ( .A(n79234), .B(n79233), .Z(n79235) );
  NOR U99340 ( .A(n87824), .B(n79235), .Z(n82125) );
  NOR U99341 ( .A(n79236), .B(n82125), .Z(n79237) );
  NOR U99342 ( .A(n87846), .B(n79237), .Z(n82114) );
  XOR U99343 ( .A(n79238), .B(n82114), .Z(n82108) );
  XOR U99344 ( .A(n79239), .B(n82108), .Z(n82100) );
  XOR U99345 ( .A(n79240), .B(n82100), .Z(n82096) );
  IV U99346 ( .A(n79241), .Z(n79242) );
  NOR U99347 ( .A(n79243), .B(n79242), .Z(n82094) );
  XOR U99348 ( .A(n82096), .B(n82094), .Z(n82098) );
  XOR U99349 ( .A(n82097), .B(n82098), .Z(n82086) );
  XOR U99350 ( .A(n82088), .B(n82086), .Z(n82084) );
  IV U99351 ( .A(n79244), .Z(n79249) );
  IV U99352 ( .A(n79245), .Z(n79247) );
  NOR U99353 ( .A(n79247), .B(n79246), .Z(n79248) );
  IV U99354 ( .A(n79248), .Z(n79252) );
  NOR U99355 ( .A(n79249), .B(n79252), .Z(n82082) );
  NOR U99356 ( .A(n82089), .B(n82082), .Z(n79250) );
  XOR U99357 ( .A(n82084), .B(n79250), .Z(n82078) );
  IV U99358 ( .A(n79251), .Z(n79253) );
  NOR U99359 ( .A(n79253), .B(n79252), .Z(n82079) );
  IV U99360 ( .A(n79254), .Z(n79257) );
  NOR U99361 ( .A(n79255), .B(n79264), .Z(n79256) );
  IV U99362 ( .A(n79256), .Z(n79260) );
  NOR U99363 ( .A(n79257), .B(n79260), .Z(n85091) );
  NOR U99364 ( .A(n82079), .B(n85091), .Z(n79258) );
  XOR U99365 ( .A(n82078), .B(n79258), .Z(n82077) );
  IV U99366 ( .A(n79259), .Z(n79261) );
  NOR U99367 ( .A(n79261), .B(n79260), .Z(n82075) );
  XOR U99368 ( .A(n82077), .B(n82075), .Z(n85098) );
  IV U99369 ( .A(n79262), .Z(n79263) );
  NOR U99370 ( .A(n79264), .B(n79263), .Z(n85096) );
  XOR U99371 ( .A(n85098), .B(n85096), .Z(n85100) );
  XOR U99372 ( .A(n85099), .B(n85100), .Z(n85105) );
  IV U99373 ( .A(n85105), .Z(n79273) );
  XOR U99374 ( .A(n85104), .B(n79273), .Z(n79269) );
  IV U99375 ( .A(n79265), .Z(n79266) );
  NOR U99376 ( .A(n79267), .B(n79266), .Z(n79272) );
  IV U99377 ( .A(n79272), .Z(n82072) );
  NOR U99378 ( .A(n79273), .B(n82072), .Z(n79268) );
  NOR U99379 ( .A(n79269), .B(n79268), .Z(n79270) );
  NOR U99380 ( .A(n79271), .B(n79270), .Z(n82073) );
  NOR U99381 ( .A(n85104), .B(n79272), .Z(n79274) );
  XOR U99382 ( .A(n79274), .B(n79273), .Z(n79279) );
  IV U99383 ( .A(n79279), .Z(n79275) );
  NOR U99384 ( .A(n79276), .B(n79275), .Z(n79277) );
  NOR U99385 ( .A(n82073), .B(n79277), .Z(n79287) );
  NOR U99386 ( .A(n79278), .B(n79287), .Z(n79281) );
  IV U99387 ( .A(n79278), .Z(n79280) );
  NOR U99388 ( .A(n79280), .B(n79279), .Z(n82071) );
  NOR U99389 ( .A(n79281), .B(n82071), .Z(n82063) );
  IV U99390 ( .A(n79282), .Z(n79284) );
  NOR U99391 ( .A(n79284), .B(n79283), .Z(n82064) );
  XOR U99392 ( .A(n82063), .B(n82064), .Z(n79285) );
  NOR U99393 ( .A(n79286), .B(n79285), .Z(n79290) );
  IV U99394 ( .A(n79286), .Z(n79289) );
  IV U99395 ( .A(n79287), .Z(n79288) );
  NOR U99396 ( .A(n79289), .B(n79288), .Z(n82067) );
  NOR U99397 ( .A(n79290), .B(n82067), .Z(n82056) );
  XOR U99398 ( .A(n79291), .B(n82056), .Z(n82054) );
  XOR U99399 ( .A(n79292), .B(n82054), .Z(n82033) );
  XOR U99400 ( .A(n82031), .B(n82033), .Z(n82036) );
  XOR U99401 ( .A(n82034), .B(n82036), .Z(n82025) );
  XOR U99402 ( .A(n82023), .B(n82025), .Z(n85138) );
  XOR U99403 ( .A(n85128), .B(n85138), .Z(n82013) );
  XOR U99404 ( .A(n79293), .B(n82013), .Z(n82011) );
  XOR U99405 ( .A(n82009), .B(n82011), .Z(n82007) );
  XOR U99406 ( .A(n82006), .B(n82007), .Z(n85143) );
  IV U99407 ( .A(n79294), .Z(n79296) );
  NOR U99408 ( .A(n79296), .B(n79295), .Z(n85142) );
  IV U99409 ( .A(n79297), .Z(n79299) );
  NOR U99410 ( .A(n79299), .B(n79298), .Z(n79300) );
  IV U99411 ( .A(n79300), .Z(n79301) );
  NOR U99412 ( .A(n79301), .B(n79304), .Z(n82004) );
  NOR U99413 ( .A(n85142), .B(n82004), .Z(n79302) );
  XOR U99414 ( .A(n85143), .B(n79302), .Z(n85145) );
  IV U99415 ( .A(n79303), .Z(n79308) );
  NOR U99416 ( .A(n79305), .B(n79304), .Z(n79306) );
  IV U99417 ( .A(n79306), .Z(n79307) );
  NOR U99418 ( .A(n79308), .B(n79307), .Z(n79309) );
  IV U99419 ( .A(n79309), .Z(n85146) );
  XOR U99420 ( .A(n85145), .B(n85146), .Z(n85149) );
  XOR U99421 ( .A(n85148), .B(n85149), .Z(n85153) );
  XOR U99422 ( .A(n85152), .B(n85153), .Z(n85157) );
  XOR U99423 ( .A(n85155), .B(n85157), .Z(n82002) );
  XOR U99424 ( .A(n82001), .B(n82002), .Z(n85161) );
  XOR U99425 ( .A(n85159), .B(n85161), .Z(n85164) );
  XOR U99426 ( .A(n85162), .B(n85164), .Z(n82000) );
  NOR U99427 ( .A(n79311), .B(n79310), .Z(n81996) );
  IV U99428 ( .A(n79312), .Z(n79314) );
  NOR U99429 ( .A(n79314), .B(n79313), .Z(n81998) );
  NOR U99430 ( .A(n81996), .B(n81998), .Z(n79315) );
  XOR U99431 ( .A(n82000), .B(n79315), .Z(n79316) );
  NOR U99432 ( .A(n79317), .B(n79316), .Z(n79320) );
  IV U99433 ( .A(n79317), .Z(n79319) );
  XOR U99434 ( .A(n81998), .B(n82000), .Z(n79318) );
  NOR U99435 ( .A(n79319), .B(n79318), .Z(n90848) );
  NOR U99436 ( .A(n79320), .B(n90848), .Z(n85166) );
  IV U99437 ( .A(n79321), .Z(n79324) );
  IV U99438 ( .A(n79322), .Z(n79323) );
  NOR U99439 ( .A(n79324), .B(n79323), .Z(n79325) );
  IV U99440 ( .A(n79325), .Z(n85167) );
  XOR U99441 ( .A(n85166), .B(n85167), .Z(n81991) );
  XOR U99442 ( .A(n81990), .B(n81991), .Z(n81994) );
  XOR U99443 ( .A(n81993), .B(n81994), .Z(n81988) );
  XOR U99444 ( .A(n81989), .B(n81988), .Z(n81983) );
  IV U99445 ( .A(n79326), .Z(n79327) );
  NOR U99446 ( .A(n79327), .B(n79331), .Z(n81982) );
  NOR U99447 ( .A(n81986), .B(n81982), .Z(n79328) );
  XOR U99448 ( .A(n81983), .B(n79328), .Z(n81981) );
  IV U99449 ( .A(n79329), .Z(n79330) );
  NOR U99450 ( .A(n79331), .B(n79330), .Z(n79332) );
  XOR U99451 ( .A(n81981), .B(n79332), .Z(n81971) );
  IV U99452 ( .A(n79333), .Z(n81970) );
  NOR U99453 ( .A(n79334), .B(n81970), .Z(n79338) );
  IV U99454 ( .A(n79335), .Z(n79336) );
  NOR U99455 ( .A(n81977), .B(n79336), .Z(n79337) );
  NOR U99456 ( .A(n79338), .B(n79337), .Z(n79339) );
  XOR U99457 ( .A(n81971), .B(n79339), .Z(n81959) );
  XOR U99458 ( .A(n79340), .B(n81959), .Z(n81952) );
  XOR U99459 ( .A(n81950), .B(n81952), .Z(n81941) );
  NOR U99460 ( .A(n79341), .B(n81944), .Z(n79350) );
  IV U99461 ( .A(n79342), .Z(n79344) );
  NOR U99462 ( .A(n79344), .B(n79343), .Z(n81940) );
  NOR U99463 ( .A(n79350), .B(n81940), .Z(n79345) );
  XOR U99464 ( .A(n81941), .B(n79345), .Z(n79353) );
  IV U99465 ( .A(n79353), .Z(n79346) );
  NOR U99466 ( .A(n79347), .B(n79346), .Z(n87656) );
  NOR U99467 ( .A(n79349), .B(n79348), .Z(n79354) );
  IV U99468 ( .A(n79354), .Z(n79352) );
  XOR U99469 ( .A(n79350), .B(n81941), .Z(n79351) );
  NOR U99470 ( .A(n79352), .B(n79351), .Z(n90877) );
  NOR U99471 ( .A(n79354), .B(n79353), .Z(n79355) );
  NOR U99472 ( .A(n90877), .B(n79355), .Z(n79357) );
  NOR U99473 ( .A(n79357), .B(n79356), .Z(n79358) );
  NOR U99474 ( .A(n87656), .B(n79358), .Z(n85178) );
  XOR U99475 ( .A(n85180), .B(n85178), .Z(n85174) );
  IV U99476 ( .A(n85174), .Z(n90906) );
  IV U99477 ( .A(n79359), .Z(n79360) );
  NOR U99478 ( .A(n90894), .B(n79360), .Z(n90907) );
  NOR U99479 ( .A(n90907), .B(n81938), .Z(n79361) );
  XOR U99480 ( .A(n90906), .B(n79361), .Z(n85192) );
  XOR U99481 ( .A(n85191), .B(n85192), .Z(n85189) );
  XOR U99482 ( .A(n85187), .B(n85189), .Z(n81937) );
  XOR U99483 ( .A(n81935), .B(n81937), .Z(n85211) );
  XOR U99484 ( .A(n79362), .B(n85211), .Z(n85206) );
  XOR U99485 ( .A(n85207), .B(n85206), .Z(n85204) );
  XOR U99486 ( .A(n79363), .B(n85204), .Z(n81926) );
  IV U99487 ( .A(n79364), .Z(n79366) );
  NOR U99488 ( .A(n79366), .B(n79365), .Z(n81932) );
  IV U99489 ( .A(n79367), .Z(n79368) );
  NOR U99490 ( .A(n79369), .B(n79368), .Z(n81927) );
  NOR U99491 ( .A(n81932), .B(n81927), .Z(n79370) );
  XOR U99492 ( .A(n81926), .B(n79370), .Z(n85218) );
  XOR U99493 ( .A(n85216), .B(n85218), .Z(n81916) );
  XOR U99494 ( .A(n79371), .B(n81916), .Z(n81920) );
  XOR U99495 ( .A(n79372), .B(n81920), .Z(n85230) );
  IV U99496 ( .A(n79373), .Z(n79374) );
  NOR U99497 ( .A(n79375), .B(n79374), .Z(n81913) );
  IV U99498 ( .A(n79376), .Z(n79378) );
  NOR U99499 ( .A(n79378), .B(n79377), .Z(n85228) );
  NOR U99500 ( .A(n81913), .B(n85228), .Z(n79379) );
  XOR U99501 ( .A(n85230), .B(n79379), .Z(n79380) );
  NOR U99502 ( .A(n79381), .B(n79380), .Z(n79384) );
  IV U99503 ( .A(n79381), .Z(n79383) );
  XOR U99504 ( .A(n81913), .B(n85230), .Z(n79382) );
  NOR U99505 ( .A(n79383), .B(n79382), .Z(n85227) );
  NOR U99506 ( .A(n79384), .B(n85227), .Z(n81904) );
  XOR U99507 ( .A(n81912), .B(n81904), .Z(n81901) );
  XOR U99508 ( .A(n79385), .B(n81901), .Z(n81898) );
  IV U99509 ( .A(n79386), .Z(n79388) );
  NOR U99510 ( .A(n79388), .B(n79387), .Z(n81895) );
  XOR U99511 ( .A(n81898), .B(n81895), .Z(n79389) );
  XOR U99512 ( .A(n79390), .B(n79389), .Z(n81888) );
  IV U99513 ( .A(n79391), .Z(n81889) );
  NOR U99514 ( .A(n81889), .B(n79392), .Z(n79393) );
  XOR U99515 ( .A(n81888), .B(n79393), .Z(n81886) );
  IV U99516 ( .A(n79394), .Z(n79395) );
  NOR U99517 ( .A(n81889), .B(n79395), .Z(n81884) );
  XOR U99518 ( .A(n81886), .B(n81884), .Z(n85240) );
  XOR U99519 ( .A(n85239), .B(n85240), .Z(n85247) );
  XOR U99520 ( .A(n79396), .B(n85247), .Z(n81877) );
  IV U99521 ( .A(n79397), .Z(n79399) );
  NOR U99522 ( .A(n79399), .B(n79398), .Z(n81879) );
  IV U99523 ( .A(n79400), .Z(n79402) );
  IV U99524 ( .A(n79401), .Z(n79406) );
  NOR U99525 ( .A(n79402), .B(n79406), .Z(n81876) );
  NOR U99526 ( .A(n81879), .B(n81876), .Z(n79403) );
  XOR U99527 ( .A(n81877), .B(n79403), .Z(n81875) );
  IV U99528 ( .A(n81875), .Z(n79409) );
  IV U99529 ( .A(n79412), .Z(n79404) );
  NOR U99530 ( .A(n79411), .B(n79404), .Z(n81871) );
  IV U99531 ( .A(n79405), .Z(n79407) );
  NOR U99532 ( .A(n79407), .B(n79406), .Z(n81873) );
  NOR U99533 ( .A(n81871), .B(n81873), .Z(n79408) );
  XOR U99534 ( .A(n79409), .B(n79408), .Z(n81864) );
  XOR U99535 ( .A(n81863), .B(n81864), .Z(n81867) );
  XOR U99536 ( .A(n81866), .B(n81867), .Z(n81862) );
  IV U99537 ( .A(n79410), .Z(n79414) );
  XOR U99538 ( .A(n79412), .B(n79411), .Z(n79413) );
  NOR U99539 ( .A(n79414), .B(n79413), .Z(n81860) );
  XOR U99540 ( .A(n81862), .B(n81860), .Z(n85253) );
  IV U99541 ( .A(n79415), .Z(n79416) );
  NOR U99542 ( .A(n79417), .B(n79416), .Z(n85251) );
  XOR U99543 ( .A(n85253), .B(n85251), .Z(n85256) );
  XOR U99544 ( .A(n79419), .B(n79418), .Z(n79434) );
  XOR U99545 ( .A(n79421), .B(n79420), .Z(n79425) );
  XOR U99546 ( .A(n79423), .B(n79422), .Z(n79424) );
  NOR U99547 ( .A(n79425), .B(n79424), .Z(n79426) );
  IV U99548 ( .A(n79426), .Z(n79431) );
  NOR U99549 ( .A(n79428), .B(n79427), .Z(n79429) );
  IV U99550 ( .A(n79429), .Z(n79430) );
  NOR U99551 ( .A(n79431), .B(n79430), .Z(n79432) );
  IV U99552 ( .A(n79432), .Z(n79433) );
  NOR U99553 ( .A(n79434), .B(n79433), .Z(n85254) );
  XOR U99554 ( .A(n85256), .B(n85254), .Z(n85259) );
  XOR U99555 ( .A(n81852), .B(n85259), .Z(n79435) );
  XOR U99556 ( .A(n79436), .B(n79435), .Z(n81850) );
  IV U99557 ( .A(n79437), .Z(n79438) );
  NOR U99558 ( .A(n79439), .B(n79438), .Z(n81848) );
  XOR U99559 ( .A(n81850), .B(n81848), .Z(n85269) );
  IV U99560 ( .A(n85269), .Z(n79447) );
  IV U99561 ( .A(n79440), .Z(n79441) );
  NOR U99562 ( .A(n79442), .B(n79441), .Z(n85268) );
  IV U99563 ( .A(n79443), .Z(n79445) );
  NOR U99564 ( .A(n79445), .B(n79444), .Z(n81846) );
  NOR U99565 ( .A(n85268), .B(n81846), .Z(n79446) );
  XOR U99566 ( .A(n79447), .B(n79446), .Z(n87602) );
  IV U99567 ( .A(n79448), .Z(n79449) );
  NOR U99568 ( .A(n79449), .B(n79451), .Z(n85271) );
  IV U99569 ( .A(n79450), .Z(n79452) );
  NOR U99570 ( .A(n79452), .B(n79451), .Z(n85264) );
  NOR U99571 ( .A(n85271), .B(n85264), .Z(n87601) );
  XOR U99572 ( .A(n87602), .B(n87601), .Z(n81844) );
  IV U99573 ( .A(n79453), .Z(n79455) );
  NOR U99574 ( .A(n79455), .B(n79454), .Z(n85276) );
  IV U99575 ( .A(n79456), .Z(n79458) );
  NOR U99576 ( .A(n79458), .B(n79457), .Z(n85277) );
  NOR U99577 ( .A(n85276), .B(n85277), .Z(n79459) );
  XOR U99578 ( .A(n81844), .B(n79459), .Z(n79465) );
  NOR U99579 ( .A(n79460), .B(n79465), .Z(n87553) );
  XOR U99580 ( .A(n81844), .B(n85277), .Z(n79464) );
  IV U99581 ( .A(n79461), .Z(n79463) );
  NOR U99582 ( .A(n79463), .B(n79462), .Z(n79466) );
  IV U99583 ( .A(n79466), .Z(n81845) );
  NOR U99584 ( .A(n79464), .B(n81845), .Z(n79468) );
  NOR U99585 ( .A(n79466), .B(n79465), .Z(n79467) );
  NOR U99586 ( .A(n79468), .B(n79467), .Z(n79474) );
  IV U99587 ( .A(n79474), .Z(n79469) );
  NOR U99588 ( .A(n79470), .B(n79469), .Z(n79471) );
  NOR U99589 ( .A(n87553), .B(n79471), .Z(n79472) );
  NOR U99590 ( .A(n79473), .B(n79472), .Z(n79476) );
  IV U99591 ( .A(n79473), .Z(n79475) );
  NOR U99592 ( .A(n79475), .B(n79474), .Z(n87543) );
  NOR U99593 ( .A(n79476), .B(n87543), .Z(n81836) );
  IV U99594 ( .A(n79477), .Z(n79478) );
  NOR U99595 ( .A(n79479), .B(n79478), .Z(n79480) );
  IV U99596 ( .A(n79480), .Z(n81838) );
  XOR U99597 ( .A(n81836), .B(n81838), .Z(n81840) );
  XOR U99598 ( .A(n81839), .B(n81840), .Z(n87539) );
  IV U99599 ( .A(n79481), .Z(n79482) );
  NOR U99600 ( .A(n79487), .B(n79482), .Z(n81833) );
  IV U99601 ( .A(n79483), .Z(n79485) );
  NOR U99602 ( .A(n79485), .B(n79484), .Z(n87541) );
  IV U99603 ( .A(n79486), .Z(n79488) );
  NOR U99604 ( .A(n79488), .B(n79487), .Z(n91008) );
  NOR U99605 ( .A(n87541), .B(n91008), .Z(n81835) );
  IV U99606 ( .A(n81835), .Z(n81830) );
  NOR U99607 ( .A(n81833), .B(n81830), .Z(n79489) );
  XOR U99608 ( .A(n87539), .B(n79489), .Z(n81825) );
  IV U99609 ( .A(n79490), .Z(n79491) );
  NOR U99610 ( .A(n79492), .B(n79491), .Z(n81829) );
  IV U99611 ( .A(n79493), .Z(n79494) );
  NOR U99612 ( .A(n79494), .B(n79496), .Z(n81826) );
  NOR U99613 ( .A(n81829), .B(n81826), .Z(n79495) );
  XOR U99614 ( .A(n81825), .B(n79495), .Z(n81824) );
  NOR U99615 ( .A(n79497), .B(n79496), .Z(n79498) );
  IV U99616 ( .A(n79498), .Z(n79499) );
  NOR U99617 ( .A(n79500), .B(n79499), .Z(n81822) );
  IV U99618 ( .A(n79501), .Z(n79503) );
  NOR U99619 ( .A(n79503), .B(n79502), .Z(n81820) );
  NOR U99620 ( .A(n81822), .B(n81820), .Z(n79504) );
  XOR U99621 ( .A(n81824), .B(n79504), .Z(n81817) );
  IV U99622 ( .A(n79505), .Z(n79507) );
  NOR U99623 ( .A(n79507), .B(n79506), .Z(n79508) );
  IV U99624 ( .A(n79508), .Z(n81818) );
  XOR U99625 ( .A(n81817), .B(n81818), .Z(n85289) );
  XOR U99626 ( .A(n85288), .B(n85289), .Z(n85282) );
  NOR U99627 ( .A(n85295), .B(n85281), .Z(n79509) );
  NOR U99628 ( .A(n79509), .B(n85283), .Z(n79510) );
  XOR U99629 ( .A(n85282), .B(n79510), .Z(n85301) );
  IV U99630 ( .A(n85301), .Z(n81810) );
  XOR U99631 ( .A(n81812), .B(n81810), .Z(n79511) );
  XOR U99632 ( .A(n79512), .B(n79511), .Z(n81807) );
  IV U99633 ( .A(n79513), .Z(n79515) );
  NOR U99634 ( .A(n79515), .B(n79514), .Z(n81808) );
  IV U99635 ( .A(n79516), .Z(n79522) );
  XOR U99636 ( .A(n79518), .B(n79517), .Z(n79519) );
  NOR U99637 ( .A(n79520), .B(n79519), .Z(n79521) );
  IV U99638 ( .A(n79521), .Z(n79525) );
  NOR U99639 ( .A(n79522), .B(n79525), .Z(n85307) );
  NOR U99640 ( .A(n81808), .B(n85307), .Z(n79523) );
  XOR U99641 ( .A(n81807), .B(n79523), .Z(n85306) );
  IV U99642 ( .A(n79524), .Z(n79526) );
  NOR U99643 ( .A(n79526), .B(n79525), .Z(n85304) );
  XOR U99644 ( .A(n85306), .B(n85304), .Z(n81801) );
  IV U99645 ( .A(n79527), .Z(n79528) );
  NOR U99646 ( .A(n79529), .B(n79528), .Z(n81799) );
  XOR U99647 ( .A(n81801), .B(n81799), .Z(n81804) );
  IV U99648 ( .A(n79530), .Z(n79531) );
  NOR U99649 ( .A(n79532), .B(n79531), .Z(n81802) );
  XOR U99650 ( .A(n81804), .B(n81802), .Z(n81797) );
  XOR U99651 ( .A(n81796), .B(n81797), .Z(n85322) );
  IV U99652 ( .A(n79533), .Z(n79535) );
  NOR U99653 ( .A(n79535), .B(n79534), .Z(n85320) );
  XOR U99654 ( .A(n85322), .B(n85320), .Z(n85324) );
  IV U99655 ( .A(n85324), .Z(n79541) );
  IV U99656 ( .A(n79536), .Z(n79537) );
  NOR U99657 ( .A(n79538), .B(n79537), .Z(n85323) );
  IV U99658 ( .A(n79543), .Z(n79539) );
  NOR U99659 ( .A(n85329), .B(n79539), .Z(n81794) );
  NOR U99660 ( .A(n85323), .B(n81794), .Z(n79540) );
  XOR U99661 ( .A(n79541), .B(n79540), .Z(n85330) );
  XOR U99662 ( .A(n79542), .B(n85330), .Z(n85341) );
  XOR U99663 ( .A(n79543), .B(n85329), .Z(n79547) );
  XOR U99664 ( .A(n79545), .B(n79544), .Z(n79546) );
  NOR U99665 ( .A(n79547), .B(n79546), .Z(n79548) );
  IV U99666 ( .A(n79548), .Z(n79553) );
  NOR U99667 ( .A(n79550), .B(n79549), .Z(n79551) );
  IV U99668 ( .A(n79551), .Z(n79552) );
  NOR U99669 ( .A(n79553), .B(n79552), .Z(n85339) );
  XOR U99670 ( .A(n85341), .B(n85339), .Z(n85344) );
  XOR U99671 ( .A(n85342), .B(n85344), .Z(n79554) );
  NOR U99672 ( .A(n79555), .B(n79554), .Z(n81791) );
  IV U99673 ( .A(n79556), .Z(n79558) );
  NOR U99674 ( .A(n79558), .B(n79557), .Z(n81792) );
  NOR U99675 ( .A(n81792), .B(n85342), .Z(n79559) );
  XOR U99676 ( .A(n79559), .B(n85344), .Z(n81786) );
  NOR U99677 ( .A(n79560), .B(n81786), .Z(n79561) );
  NOR U99678 ( .A(n81791), .B(n79561), .Z(n85348) );
  XOR U99679 ( .A(n79562), .B(n85348), .Z(n85357) );
  XOR U99680 ( .A(n79563), .B(n85357), .Z(n85354) );
  XOR U99681 ( .A(n85352), .B(n85354), .Z(n81778) );
  XOR U99682 ( .A(n81777), .B(n81778), .Z(n81781) );
  XOR U99683 ( .A(n81780), .B(n81781), .Z(n85364) );
  XOR U99684 ( .A(n85363), .B(n85364), .Z(n85361) );
  XOR U99685 ( .A(n85362), .B(n85361), .Z(n81769) );
  XOR U99686 ( .A(n81771), .B(n81769), .Z(n81773) );
  XOR U99687 ( .A(n81772), .B(n81773), .Z(n79564) );
  NOR U99688 ( .A(n79565), .B(n79564), .Z(n87516) );
  IV U99689 ( .A(n79566), .Z(n79568) );
  NOR U99690 ( .A(n79568), .B(n79567), .Z(n81766) );
  NOR U99691 ( .A(n81766), .B(n81772), .Z(n79569) );
  XOR U99692 ( .A(n79569), .B(n81773), .Z(n79574) );
  NOR U99693 ( .A(n79570), .B(n79574), .Z(n79571) );
  NOR U99694 ( .A(n87516), .B(n79571), .Z(n79572) );
  NOR U99695 ( .A(n79573), .B(n79572), .Z(n79577) );
  IV U99696 ( .A(n79573), .Z(n79576) );
  IV U99697 ( .A(n79574), .Z(n79575) );
  NOR U99698 ( .A(n79576), .B(n79575), .Z(n81765) );
  NOR U99699 ( .A(n79577), .B(n81765), .Z(n85378) );
  IV U99700 ( .A(n79578), .Z(n79580) );
  NOR U99701 ( .A(n79580), .B(n79579), .Z(n85377) );
  XOR U99702 ( .A(n85378), .B(n85377), .Z(n79585) );
  IV U99703 ( .A(n79585), .Z(n81763) );
  NOR U99704 ( .A(n79584), .B(n81763), .Z(n91134) );
  IV U99705 ( .A(n79581), .Z(n79582) );
  NOR U99706 ( .A(n79583), .B(n79582), .Z(n81762) );
  XOR U99707 ( .A(n81762), .B(n79585), .Z(n79587) );
  NOR U99708 ( .A(n79585), .B(n79584), .Z(n79586) );
  NOR U99709 ( .A(n79587), .B(n79586), .Z(n81759) );
  NOR U99710 ( .A(n91134), .B(n81759), .Z(n81754) );
  XOR U99711 ( .A(n91165), .B(n81754), .Z(n81751) );
  XOR U99712 ( .A(n79588), .B(n81751), .Z(n81737) );
  XOR U99713 ( .A(n81746), .B(n81737), .Z(n81731) );
  IV U99714 ( .A(n79589), .Z(n79590) );
  NOR U99715 ( .A(n79590), .B(n81738), .Z(n81729) );
  XOR U99716 ( .A(n81731), .B(n81729), .Z(n81727) );
  XOR U99717 ( .A(n81726), .B(n81727), .Z(n81720) );
  XOR U99718 ( .A(n81721), .B(n81720), .Z(n79596) );
  IV U99719 ( .A(n79596), .Z(n81722) );
  NOR U99720 ( .A(n79591), .B(n81722), .Z(n81719) );
  IV U99721 ( .A(n79592), .Z(n79593) );
  NOR U99722 ( .A(n79594), .B(n79593), .Z(n79595) );
  IV U99723 ( .A(n79595), .Z(n81723) );
  XOR U99724 ( .A(n81723), .B(n79596), .Z(n85395) );
  IV U99725 ( .A(n85395), .Z(n79597) );
  NOR U99726 ( .A(n79598), .B(n79597), .Z(n79599) );
  NOR U99727 ( .A(n81719), .B(n79599), .Z(n79612) );
  IV U99728 ( .A(n79600), .Z(n79603) );
  XOR U99729 ( .A(n79601), .B(n79604), .Z(n79602) );
  NOR U99730 ( .A(n79603), .B(n79602), .Z(n81717) );
  NOR U99731 ( .A(n79605), .B(n79604), .Z(n79606) );
  IV U99732 ( .A(n79606), .Z(n79617) );
  NOR U99733 ( .A(n79607), .B(n79617), .Z(n79608) );
  IV U99734 ( .A(n79608), .Z(n79609) );
  NOR U99735 ( .A(n79610), .B(n79609), .Z(n85393) );
  NOR U99736 ( .A(n81717), .B(n85393), .Z(n79611) );
  XOR U99737 ( .A(n79612), .B(n79611), .Z(n85399) );
  IV U99738 ( .A(n79613), .Z(n79625) );
  IV U99739 ( .A(n79614), .Z(n79615) );
  NOR U99740 ( .A(n79625), .B(n79615), .Z(n81715) );
  IV U99741 ( .A(n79616), .Z(n79618) );
  NOR U99742 ( .A(n79618), .B(n79617), .Z(n85397) );
  NOR U99743 ( .A(n81715), .B(n85397), .Z(n79619) );
  XOR U99744 ( .A(n85399), .B(n79619), .Z(n81710) );
  IV U99745 ( .A(n79620), .Z(n79621) );
  NOR U99746 ( .A(n79622), .B(n79621), .Z(n81709) );
  IV U99747 ( .A(n79623), .Z(n79624) );
  NOR U99748 ( .A(n79625), .B(n79624), .Z(n81712) );
  NOR U99749 ( .A(n81709), .B(n81712), .Z(n79626) );
  XOR U99750 ( .A(n81710), .B(n79626), .Z(n81703) );
  IV U99751 ( .A(n79627), .Z(n79629) );
  NOR U99752 ( .A(n79629), .B(n79628), .Z(n81701) );
  XOR U99753 ( .A(n81703), .B(n81701), .Z(n81705) );
  XOR U99754 ( .A(n81704), .B(n81705), .Z(n85403) );
  XOR U99755 ( .A(n85402), .B(n85403), .Z(n81697) );
  XOR U99756 ( .A(n81699), .B(n81697), .Z(n79630) );
  NOR U99757 ( .A(n79631), .B(n79630), .Z(n85423) );
  NOR U99758 ( .A(n81696), .B(n81699), .Z(n79632) );
  XOR U99759 ( .A(n79632), .B(n81697), .Z(n85419) );
  NOR U99760 ( .A(n79633), .B(n85419), .Z(n79634) );
  NOR U99761 ( .A(n85423), .B(n79634), .Z(n81693) );
  IV U99762 ( .A(n79635), .Z(n79637) );
  NOR U99763 ( .A(n79637), .B(n79636), .Z(n85418) );
  IV U99764 ( .A(n79638), .Z(n79640) );
  NOR U99765 ( .A(n79640), .B(n79639), .Z(n81692) );
  NOR U99766 ( .A(n85418), .B(n81692), .Z(n79641) );
  XOR U99767 ( .A(n81693), .B(n79641), .Z(n81691) );
  XOR U99768 ( .A(n81689), .B(n81691), .Z(n85431) );
  XOR U99769 ( .A(n79642), .B(n85431), .Z(n79643) );
  IV U99770 ( .A(n79643), .Z(n85428) );
  XOR U99771 ( .A(n85426), .B(n85428), .Z(n81684) );
  XOR U99772 ( .A(n81683), .B(n81684), .Z(n81680) );
  XOR U99773 ( .A(n81679), .B(n81680), .Z(n79656) );
  IV U99774 ( .A(n79656), .Z(n79652) );
  IV U99775 ( .A(n79644), .Z(n79645) );
  NOR U99776 ( .A(n79646), .B(n79645), .Z(n79653) );
  IV U99777 ( .A(n79647), .Z(n79649) );
  NOR U99778 ( .A(n79649), .B(n79648), .Z(n79655) );
  NOR U99779 ( .A(n79653), .B(n79655), .Z(n79650) );
  IV U99780 ( .A(n79650), .Z(n79651) );
  NOR U99781 ( .A(n79652), .B(n79651), .Z(n79658) );
  IV U99782 ( .A(n79653), .Z(n79654) );
  NOR U99783 ( .A(n79654), .B(n81680), .Z(n81682) );
  IV U99784 ( .A(n79655), .Z(n79657) );
  NOR U99785 ( .A(n79657), .B(n79656), .Z(n85438) );
  NOR U99786 ( .A(n81682), .B(n85438), .Z(n91227) );
  IV U99787 ( .A(n91227), .Z(n91229) );
  NOR U99788 ( .A(n79658), .B(n91229), .Z(n81672) );
  XOR U99789 ( .A(n81674), .B(n81672), .Z(n79659) );
  XOR U99790 ( .A(n79660), .B(n79659), .Z(n85444) );
  XOR U99791 ( .A(n85443), .B(n85444), .Z(n85447) );
  XOR U99792 ( .A(n79661), .B(n85447), .Z(n81667) );
  IV U99793 ( .A(n79662), .Z(n79663) );
  NOR U99794 ( .A(n79664), .B(n79663), .Z(n79665) );
  IV U99795 ( .A(n79665), .Z(n81666) );
  XOR U99796 ( .A(n81667), .B(n81666), .Z(n79668) );
  IV U99797 ( .A(n79668), .Z(n79666) );
  NOR U99798 ( .A(n79667), .B(n79666), .Z(n91240) );
  NOR U99799 ( .A(n79669), .B(n79668), .Z(n85457) );
  IV U99800 ( .A(n79670), .Z(n79672) );
  IV U99801 ( .A(n79671), .Z(n79677) );
  NOR U99802 ( .A(n79672), .B(n79677), .Z(n85455) );
  XOR U99803 ( .A(n85457), .B(n85455), .Z(n79673) );
  NOR U99804 ( .A(n91240), .B(n79673), .Z(n81664) );
  NOR U99805 ( .A(n79675), .B(n79674), .Z(n81663) );
  IV U99806 ( .A(n79676), .Z(n79678) );
  NOR U99807 ( .A(n79678), .B(n79677), .Z(n85452) );
  NOR U99808 ( .A(n81663), .B(n85452), .Z(n79679) );
  XOR U99809 ( .A(n81664), .B(n79679), .Z(n81658) );
  XOR U99810 ( .A(n81657), .B(n81658), .Z(n81661) );
  XOR U99811 ( .A(n81660), .B(n81661), .Z(n81655) );
  XOR U99812 ( .A(n81653), .B(n81655), .Z(n81649) );
  XOR U99813 ( .A(n81647), .B(n81649), .Z(n85466) );
  IV U99814 ( .A(n79680), .Z(n79683) );
  IV U99815 ( .A(n79681), .Z(n79682) );
  NOR U99816 ( .A(n79683), .B(n79682), .Z(n79684) );
  IV U99817 ( .A(n79684), .Z(n81650) );
  XOR U99818 ( .A(n85466), .B(n81650), .Z(n79685) );
  XOR U99819 ( .A(n79686), .B(n79685), .Z(n81641) );
  XOR U99820 ( .A(n79687), .B(n81641), .Z(n81635) );
  XOR U99821 ( .A(n81634), .B(n81635), .Z(n81638) );
  XOR U99822 ( .A(n81637), .B(n81638), .Z(n81627) );
  IV U99823 ( .A(n81627), .Z(n81625) );
  XOR U99824 ( .A(n81628), .B(n81625), .Z(n85489) );
  IV U99825 ( .A(n79688), .Z(n79690) );
  NOR U99826 ( .A(n79690), .B(n79689), .Z(n81629) );
  IV U99827 ( .A(n79691), .Z(n79692) );
  NOR U99828 ( .A(n79693), .B(n79692), .Z(n85487) );
  NOR U99829 ( .A(n81629), .B(n85487), .Z(n79694) );
  XOR U99830 ( .A(n85489), .B(n79694), .Z(n79695) );
  IV U99831 ( .A(n79695), .Z(n85486) );
  IV U99832 ( .A(n79696), .Z(n79698) );
  NOR U99833 ( .A(n79698), .B(n79697), .Z(n85484) );
  XOR U99834 ( .A(n85486), .B(n85484), .Z(n81621) );
  XOR U99835 ( .A(n81619), .B(n81621), .Z(n81624) );
  XOR U99836 ( .A(n81622), .B(n81624), .Z(n81615) );
  XOR U99837 ( .A(n81613), .B(n81615), .Z(n81607) );
  XOR U99838 ( .A(n79699), .B(n81607), .Z(n85495) );
  XOR U99839 ( .A(n79700), .B(n85495), .Z(n85502) );
  XOR U99840 ( .A(n79701), .B(n85502), .Z(n79702) );
  IV U99841 ( .A(n79702), .Z(n81604) );
  XOR U99842 ( .A(n81602), .B(n81604), .Z(n85513) );
  XOR U99843 ( .A(n81605), .B(n85513), .Z(n81598) );
  IV U99844 ( .A(n79703), .Z(n79705) );
  NOR U99845 ( .A(n79705), .B(n79704), .Z(n85512) );
  IV U99846 ( .A(n79706), .Z(n79707) );
  NOR U99847 ( .A(n79707), .B(n79711), .Z(n81599) );
  NOR U99848 ( .A(n85512), .B(n81599), .Z(n79708) );
  XOR U99849 ( .A(n81598), .B(n79708), .Z(n85522) );
  IV U99850 ( .A(n79709), .Z(n79710) );
  NOR U99851 ( .A(n79711), .B(n79710), .Z(n79712) );
  IV U99852 ( .A(n79712), .Z(n85521) );
  XOR U99853 ( .A(n85522), .B(n85521), .Z(n79716) );
  IV U99854 ( .A(n79716), .Z(n79713) );
  NOR U99855 ( .A(n79714), .B(n79713), .Z(n87341) );
  IV U99856 ( .A(n79717), .Z(n79715) );
  NOR U99857 ( .A(n85522), .B(n79715), .Z(n87338) );
  NOR U99858 ( .A(n79717), .B(n79716), .Z(n79718) );
  NOR U99859 ( .A(n87338), .B(n79718), .Z(n81595) );
  NOR U99860 ( .A(n79719), .B(n81595), .Z(n79720) );
  NOR U99861 ( .A(n87341), .B(n79720), .Z(n81590) );
  NOR U99862 ( .A(n79722), .B(n79721), .Z(n79723) );
  IV U99863 ( .A(n79723), .Z(n79730) );
  XOR U99864 ( .A(n79725), .B(n79724), .Z(n79726) );
  NOR U99865 ( .A(n79727), .B(n79726), .Z(n79728) );
  IV U99866 ( .A(n79728), .Z(n79729) );
  NOR U99867 ( .A(n79730), .B(n79729), .Z(n81591) );
  NOR U99868 ( .A(n81594), .B(n81591), .Z(n79731) );
  XOR U99869 ( .A(n81590), .B(n79731), .Z(n81589) );
  XOR U99870 ( .A(n81586), .B(n81589), .Z(n79732) );
  XOR U99871 ( .A(n81588), .B(n79732), .Z(n81584) );
  XOR U99872 ( .A(n81583), .B(n81584), .Z(n81579) );
  XOR U99873 ( .A(n81577), .B(n81579), .Z(n81582) );
  XOR U99874 ( .A(n81580), .B(n81582), .Z(n81574) );
  XOR U99875 ( .A(n81572), .B(n81574), .Z(n85528) );
  XOR U99876 ( .A(n79733), .B(n85528), .Z(n85525) );
  XOR U99877 ( .A(n85527), .B(n85525), .Z(n81570) );
  XOR U99878 ( .A(n79734), .B(n81570), .Z(n79735) );
  IV U99879 ( .A(n79735), .Z(n81562) );
  XOR U99880 ( .A(n81560), .B(n81562), .Z(n81563) );
  IV U99881 ( .A(n79736), .Z(n79739) );
  NOR U99882 ( .A(n79737), .B(n79739), .Z(n79750) );
  XOR U99883 ( .A(n79738), .B(n79740), .Z(n79742) );
  NOR U99884 ( .A(n79740), .B(n79739), .Z(n79741) );
  NOR U99885 ( .A(n79742), .B(n79741), .Z(n79748) );
  IV U99886 ( .A(n79743), .Z(n79745) );
  NOR U99887 ( .A(n79745), .B(n79744), .Z(n79746) );
  IV U99888 ( .A(n79746), .Z(n79747) );
  NOR U99889 ( .A(n79748), .B(n79747), .Z(n79749) );
  NOR U99890 ( .A(n79750), .B(n79749), .Z(n81564) );
  XOR U99891 ( .A(n81563), .B(n81564), .Z(n81554) );
  IV U99892 ( .A(n81554), .Z(n81552) );
  XOR U99893 ( .A(n81553), .B(n81552), .Z(n81549) );
  XOR U99894 ( .A(n81538), .B(n81549), .Z(n81536) );
  XOR U99895 ( .A(n79751), .B(n81536), .Z(n79752) );
  IV U99896 ( .A(n79752), .Z(n81530) );
  XOR U99897 ( .A(n81529), .B(n81530), .Z(n81532) );
  XOR U99898 ( .A(n81533), .B(n81532), .Z(n81521) );
  IV U99899 ( .A(n79753), .Z(n79755) );
  NOR U99900 ( .A(n79755), .B(n79754), .Z(n79756) );
  IV U99901 ( .A(n79756), .Z(n81522) );
  XOR U99902 ( .A(n81521), .B(n81522), .Z(n81525) );
  IV U99903 ( .A(n79757), .Z(n79758) );
  NOR U99904 ( .A(n79759), .B(n79758), .Z(n81524) );
  IV U99905 ( .A(n79760), .Z(n79762) );
  NOR U99906 ( .A(n79762), .B(n79761), .Z(n81519) );
  NOR U99907 ( .A(n81519), .B(n81517), .Z(n79763) );
  IV U99908 ( .A(n79763), .Z(n79764) );
  NOR U99909 ( .A(n81524), .B(n79764), .Z(n79765) );
  XOR U99910 ( .A(n81525), .B(n79765), .Z(n79779) );
  IV U99911 ( .A(n79779), .Z(n79770) );
  IV U99912 ( .A(n79766), .Z(n79767) );
  NOR U99913 ( .A(n79768), .B(n79767), .Z(n79783) );
  IV U99914 ( .A(n79783), .Z(n79769) );
  NOR U99915 ( .A(n79770), .B(n79769), .Z(n87299) );
  IV U99916 ( .A(n79771), .Z(n79772) );
  NOR U99917 ( .A(n79773), .B(n79772), .Z(n81513) );
  IV U99918 ( .A(n79774), .Z(n79776) );
  NOR U99919 ( .A(n79776), .B(n79775), .Z(n79780) );
  IV U99920 ( .A(n79780), .Z(n79778) );
  XOR U99921 ( .A(n81524), .B(n81525), .Z(n79777) );
  NOR U99922 ( .A(n79778), .B(n79777), .Z(n91357) );
  NOR U99923 ( .A(n79780), .B(n79779), .Z(n79781) );
  NOR U99924 ( .A(n91357), .B(n79781), .Z(n81514) );
  XOR U99925 ( .A(n81513), .B(n81514), .Z(n79782) );
  NOR U99926 ( .A(n79783), .B(n79782), .Z(n79784) );
  NOR U99927 ( .A(n87299), .B(n79784), .Z(n79785) );
  IV U99928 ( .A(n79785), .Z(n81511) );
  XOR U99929 ( .A(n81510), .B(n81511), .Z(n81507) );
  IV U99930 ( .A(n79786), .Z(n79788) );
  NOR U99931 ( .A(n79788), .B(n79787), .Z(n81509) );
  IV U99932 ( .A(n79789), .Z(n79804) );
  NOR U99933 ( .A(n79804), .B(n79790), .Z(n79791) );
  IV U99934 ( .A(n79791), .Z(n79797) );
  IV U99935 ( .A(n79792), .Z(n79793) );
  NOR U99936 ( .A(n79794), .B(n79793), .Z(n79795) );
  IV U99937 ( .A(n79795), .Z(n79796) );
  NOR U99938 ( .A(n79797), .B(n79796), .Z(n79798) );
  IV U99939 ( .A(n79798), .Z(n79799) );
  NOR U99940 ( .A(n79800), .B(n79799), .Z(n81506) );
  NOR U99941 ( .A(n81509), .B(n81506), .Z(n79801) );
  XOR U99942 ( .A(n81507), .B(n79801), .Z(n79802) );
  IV U99943 ( .A(n79802), .Z(n81505) );
  IV U99944 ( .A(n79803), .Z(n79805) );
  NOR U99945 ( .A(n79805), .B(n79804), .Z(n81503) );
  XOR U99946 ( .A(n81505), .B(n81503), .Z(n85547) );
  XOR U99947 ( .A(n81496), .B(n85547), .Z(n81500) );
  XOR U99948 ( .A(n81498), .B(n81500), .Z(n85559) );
  XOR U99949 ( .A(n85553), .B(n85559), .Z(n85563) );
  XOR U99950 ( .A(n79806), .B(n85563), .Z(n79807) );
  IV U99951 ( .A(n79807), .Z(n85565) );
  IV U99952 ( .A(n79808), .Z(n79810) );
  NOR U99953 ( .A(n79810), .B(n79809), .Z(n79811) );
  IV U99954 ( .A(n79811), .Z(n85564) );
  IV U99955 ( .A(n79812), .Z(n79814) );
  NOR U99956 ( .A(n79814), .B(n79813), .Z(n79819) );
  IV U99957 ( .A(n79815), .Z(n79817) );
  NOR U99958 ( .A(n79817), .B(n79816), .Z(n79818) );
  NOR U99959 ( .A(n79819), .B(n79818), .Z(n81495) );
  XOR U99960 ( .A(n85564), .B(n81495), .Z(n79820) );
  XOR U99961 ( .A(n85565), .B(n79820), .Z(n85568) );
  XOR U99962 ( .A(n85566), .B(n85568), .Z(n85569) );
  XOR U99963 ( .A(n85570), .B(n85569), .Z(n85576) );
  XOR U99964 ( .A(n85573), .B(n85576), .Z(n85586) );
  XOR U99965 ( .A(n79821), .B(n85586), .Z(n81482) );
  XOR U99966 ( .A(n81483), .B(n81482), .Z(n81487) );
  XOR U99967 ( .A(n81485), .B(n81487), .Z(n81475) );
  XOR U99968 ( .A(n81474), .B(n81475), .Z(n81479) );
  XOR U99969 ( .A(n81477), .B(n81479), .Z(n85597) );
  IV U99970 ( .A(n79822), .Z(n79824) );
  NOR U99971 ( .A(n79824), .B(n79823), .Z(n85596) );
  IV U99972 ( .A(n79825), .Z(n79827) );
  NOR U99973 ( .A(n79827), .B(n79826), .Z(n79828) );
  IV U99974 ( .A(n79828), .Z(n79830) );
  NOR U99975 ( .A(n79830), .B(n79829), .Z(n79831) );
  IV U99976 ( .A(n79831), .Z(n81473) );
  XOR U99977 ( .A(n85596), .B(n81473), .Z(n79832) );
  XOR U99978 ( .A(n85597), .B(n79832), .Z(n81471) );
  XOR U99979 ( .A(n79833), .B(n81471), .Z(n81469) );
  XOR U99980 ( .A(n81467), .B(n81469), .Z(n81460) );
  XOR U99981 ( .A(n81459), .B(n81460), .Z(n81463) );
  XOR U99982 ( .A(n81462), .B(n81463), .Z(n85608) );
  XOR U99983 ( .A(n85607), .B(n85608), .Z(n85610) );
  IV U99984 ( .A(n79834), .Z(n79835) );
  NOR U99985 ( .A(n79836), .B(n79835), .Z(n79841) );
  IV U99986 ( .A(n79837), .Z(n79839) );
  NOR U99987 ( .A(n79839), .B(n79838), .Z(n79840) );
  NOR U99988 ( .A(n79841), .B(n79840), .Z(n85611) );
  XOR U99989 ( .A(n85610), .B(n85611), .Z(n81452) );
  XOR U99990 ( .A(n81454), .B(n81452), .Z(n85617) );
  IV U99991 ( .A(n85617), .Z(n79851) );
  IV U99992 ( .A(n79842), .Z(n79844) );
  NOR U99993 ( .A(n79844), .B(n79843), .Z(n81455) );
  IV U99994 ( .A(n79845), .Z(n79849) );
  NOR U99995 ( .A(n79846), .B(n79854), .Z(n79847) );
  IV U99996 ( .A(n79847), .Z(n79848) );
  NOR U99997 ( .A(n79849), .B(n79848), .Z(n85615) );
  NOR U99998 ( .A(n81455), .B(n85615), .Z(n79850) );
  XOR U99999 ( .A(n79851), .B(n79850), .Z(n81451) );
  IV U100000 ( .A(n79852), .Z(n79858) );
  IV U100001 ( .A(n79853), .Z(n79855) );
  NOR U100002 ( .A(n79855), .B(n79854), .Z(n79856) );
  IV U100003 ( .A(n79856), .Z(n79857) );
  NOR U100004 ( .A(n79858), .B(n79857), .Z(n81449) );
  XOR U100005 ( .A(n81451), .B(n81449), .Z(n85621) );
  XOR U100006 ( .A(n85620), .B(n85621), .Z(n81448) );
  XOR U100007 ( .A(n81446), .B(n81448), .Z(n85633) );
  XOR U100008 ( .A(n85626), .B(n85633), .Z(n85629) );
  XOR U100009 ( .A(n79859), .B(n85629), .Z(n81439) );
  XOR U100010 ( .A(n79860), .B(n81439), .Z(n85637) );
  XOR U100011 ( .A(n85636), .B(n85637), .Z(n85643) );
  XOR U100012 ( .A(n79861), .B(n85643), .Z(n81432) );
  XOR U100013 ( .A(n81435), .B(n81432), .Z(n81430) );
  IV U100014 ( .A(n79862), .Z(n79864) );
  NOR U100015 ( .A(n79864), .B(n79863), .Z(n81429) );
  IV U100016 ( .A(n79865), .Z(n79867) );
  NOR U100017 ( .A(n79867), .B(n79866), .Z(n81433) );
  NOR U100018 ( .A(n81429), .B(n81433), .Z(n79868) );
  XOR U100019 ( .A(n81430), .B(n79868), .Z(n81421) );
  XOR U100020 ( .A(n81422), .B(n81421), .Z(n81426) );
  XOR U100021 ( .A(n81424), .B(n81426), .Z(n81415) );
  XOR U100022 ( .A(n81413), .B(n81415), .Z(n81418) );
  IV U100023 ( .A(n79869), .Z(n79870) );
  NOR U100024 ( .A(n79871), .B(n79870), .Z(n81416) );
  XOR U100025 ( .A(n81418), .B(n81416), .Z(n79872) );
  XOR U100026 ( .A(n79873), .B(n79872), .Z(n81404) );
  XOR U100027 ( .A(n81405), .B(n81404), .Z(n85648) );
  IV U100028 ( .A(n85648), .Z(n79887) );
  IV U100029 ( .A(n79874), .Z(n79876) );
  NOR U100030 ( .A(n79876), .B(n79875), .Z(n85646) );
  NOR U100031 ( .A(n79887), .B(n85646), .Z(n79885) );
  IV U100032 ( .A(n79877), .Z(n79879) );
  NOR U100033 ( .A(n79879), .B(n79878), .Z(n79884) );
  IV U100034 ( .A(n79880), .Z(n79882) );
  NOR U100035 ( .A(n79882), .B(n79881), .Z(n79883) );
  NOR U100036 ( .A(n79884), .B(n79883), .Z(n79886) );
  NOR U100037 ( .A(n79885), .B(n79886), .Z(n85649) );
  IV U100038 ( .A(n79886), .Z(n79889) );
  XOR U100039 ( .A(n85646), .B(n79887), .Z(n79888) );
  NOR U100040 ( .A(n79889), .B(n79888), .Z(n79890) );
  NOR U100041 ( .A(n85649), .B(n79890), .Z(n81392) );
  IV U100042 ( .A(n79891), .Z(n79895) );
  NOR U100043 ( .A(n79893), .B(n79892), .Z(n79894) );
  IV U100044 ( .A(n79894), .Z(n79899) );
  NOR U100045 ( .A(n79895), .B(n79899), .Z(n81393) );
  XOR U100046 ( .A(n81392), .B(n81393), .Z(n79896) );
  XOR U100047 ( .A(n79897), .B(n79896), .Z(n81397) );
  IV U100048 ( .A(n79898), .Z(n79900) );
  NOR U100049 ( .A(n79900), .B(n79899), .Z(n81395) );
  XOR U100050 ( .A(n81397), .B(n81395), .Z(n85653) );
  XOR U100051 ( .A(n85652), .B(n85653), .Z(n79911) );
  IV U100052 ( .A(n79911), .Z(n79905) );
  IV U100053 ( .A(n79901), .Z(n79903) );
  NOR U100054 ( .A(n79903), .B(n79902), .Z(n79913) );
  IV U100055 ( .A(n79913), .Z(n79904) );
  NOR U100056 ( .A(n79905), .B(n79904), .Z(n87155) );
  IV U100057 ( .A(n79906), .Z(n79908) );
  NOR U100058 ( .A(n79908), .B(n79907), .Z(n79910) );
  IV U100059 ( .A(n79910), .Z(n79909) );
  NOR U100060 ( .A(n81397), .B(n79909), .Z(n87151) );
  NOR U100061 ( .A(n79911), .B(n79910), .Z(n79912) );
  NOR U100062 ( .A(n87151), .B(n79912), .Z(n85657) );
  NOR U100063 ( .A(n79913), .B(n85657), .Z(n79914) );
  NOR U100064 ( .A(n87155), .B(n79914), .Z(n81388) );
  XOR U100065 ( .A(n79915), .B(n81388), .Z(n81382) );
  XOR U100066 ( .A(n81380), .B(n81382), .Z(n81385) );
  IV U100067 ( .A(n79916), .Z(n79917) );
  NOR U100068 ( .A(n79918), .B(n79917), .Z(n85660) );
  IV U100069 ( .A(n79919), .Z(n79921) );
  NOR U100070 ( .A(n79921), .B(n79920), .Z(n81383) );
  NOR U100071 ( .A(n85660), .B(n81383), .Z(n79922) );
  XOR U100072 ( .A(n81385), .B(n79922), .Z(n79927) );
  XOR U100073 ( .A(n85661), .B(n79927), .Z(n85662) );
  IV U100074 ( .A(n85662), .Z(n79926) );
  IV U100075 ( .A(n79923), .Z(n79924) );
  NOR U100076 ( .A(n79924), .B(n79929), .Z(n79935) );
  IV U100077 ( .A(n79935), .Z(n79925) );
  NOR U100078 ( .A(n79926), .B(n79925), .Z(n85669) );
  IV U100079 ( .A(n79927), .Z(n79932) );
  IV U100080 ( .A(n79928), .Z(n79930) );
  NOR U100081 ( .A(n79930), .B(n79929), .Z(n79933) );
  IV U100082 ( .A(n79933), .Z(n79931) );
  NOR U100083 ( .A(n79932), .B(n79931), .Z(n87160) );
  NOR U100084 ( .A(n79933), .B(n85662), .Z(n79934) );
  NOR U100085 ( .A(n87160), .B(n79934), .Z(n81378) );
  NOR U100086 ( .A(n79935), .B(n81378), .Z(n79936) );
  NOR U100087 ( .A(n85669), .B(n79936), .Z(n79945) );
  IV U100088 ( .A(n79937), .Z(n79940) );
  IV U100089 ( .A(n79938), .Z(n79939) );
  NOR U100090 ( .A(n79940), .B(n79939), .Z(n85665) );
  IV U100091 ( .A(n79941), .Z(n79943) );
  IV U100092 ( .A(n79942), .Z(n79947) );
  NOR U100093 ( .A(n79943), .B(n79947), .Z(n81377) );
  NOR U100094 ( .A(n85665), .B(n81377), .Z(n79944) );
  XOR U100095 ( .A(n79945), .B(n79944), .Z(n81373) );
  IV U100096 ( .A(n79946), .Z(n79948) );
  NOR U100097 ( .A(n79948), .B(n79947), .Z(n81371) );
  XOR U100098 ( .A(n81373), .B(n81371), .Z(n81376) );
  IV U100099 ( .A(n79949), .Z(n79951) );
  NOR U100100 ( .A(n79951), .B(n79950), .Z(n79952) );
  IV U100101 ( .A(n79952), .Z(n79954) );
  NOR U100102 ( .A(n79954), .B(n79953), .Z(n81374) );
  XOR U100103 ( .A(n81376), .B(n81374), .Z(n81366) );
  XOR U100104 ( .A(n81365), .B(n81366), .Z(n81369) );
  IV U100105 ( .A(n79955), .Z(n79956) );
  NOR U100106 ( .A(n79956), .B(n79960), .Z(n81363) );
  XOR U100107 ( .A(n81369), .B(n81363), .Z(n81361) );
  IV U100108 ( .A(n79957), .Z(n79958) );
  NOR U100109 ( .A(n79958), .B(n79960), .Z(n81360) );
  IV U100110 ( .A(n79959), .Z(n79961) );
  NOR U100111 ( .A(n79961), .B(n79960), .Z(n81368) );
  NOR U100112 ( .A(n81360), .B(n81368), .Z(n79962) );
  XOR U100113 ( .A(n81361), .B(n79962), .Z(n79973) );
  IV U100114 ( .A(n79973), .Z(n81352) );
  IV U100115 ( .A(n79963), .Z(n79964) );
  NOR U100116 ( .A(n79964), .B(n79969), .Z(n79975) );
  IV U100117 ( .A(n79975), .Z(n79965) );
  NOR U100118 ( .A(n81352), .B(n79965), .Z(n91539) );
  IV U100119 ( .A(n79966), .Z(n81354) );
  NOR U100120 ( .A(n81354), .B(n79967), .Z(n79971) );
  IV U100121 ( .A(n79968), .Z(n79970) );
  NOR U100122 ( .A(n79970), .B(n79969), .Z(n81350) );
  NOR U100123 ( .A(n79971), .B(n81350), .Z(n79972) );
  XOR U100124 ( .A(n79973), .B(n79972), .Z(n81348) );
  IV U100125 ( .A(n81348), .Z(n79974) );
  NOR U100126 ( .A(n79975), .B(n79974), .Z(n79976) );
  NOR U100127 ( .A(n91539), .B(n79976), .Z(n81343) );
  IV U100128 ( .A(n79977), .Z(n79985) );
  NOR U100129 ( .A(n79985), .B(n79978), .Z(n81342) );
  IV U100130 ( .A(n79979), .Z(n79980) );
  NOR U100131 ( .A(n79981), .B(n79980), .Z(n81346) );
  NOR U100132 ( .A(n81342), .B(n81346), .Z(n79982) );
  XOR U100133 ( .A(n81343), .B(n79982), .Z(n81338) );
  IV U100134 ( .A(n79983), .Z(n79984) );
  NOR U100135 ( .A(n79985), .B(n79984), .Z(n81336) );
  XOR U100136 ( .A(n81338), .B(n81336), .Z(n81340) );
  XOR U100137 ( .A(n81339), .B(n81340), .Z(n81331) );
  XOR U100138 ( .A(n81330), .B(n81331), .Z(n81335) );
  XOR U100139 ( .A(n81333), .B(n81335), .Z(n81324) );
  XOR U100140 ( .A(n81322), .B(n81324), .Z(n81326) );
  XOR U100141 ( .A(n81325), .B(n81326), .Z(n85675) );
  XOR U100142 ( .A(n79986), .B(n85675), .Z(n85678) );
  IV U100143 ( .A(n85678), .Z(n85681) );
  XOR U100144 ( .A(n85679), .B(n85681), .Z(n85690) );
  IV U100145 ( .A(n79987), .Z(n79989) );
  NOR U100146 ( .A(n79989), .B(n79988), .Z(n85689) );
  IV U100147 ( .A(n79990), .Z(n79991) );
  NOR U100148 ( .A(n79994), .B(n79991), .Z(n81318) );
  IV U100149 ( .A(n79992), .Z(n79993) );
  NOR U100150 ( .A(n79994), .B(n79993), .Z(n85683) );
  NOR U100151 ( .A(n81318), .B(n85683), .Z(n79995) );
  IV U100152 ( .A(n79995), .Z(n79996) );
  NOR U100153 ( .A(n85689), .B(n79996), .Z(n79997) );
  XOR U100154 ( .A(n85690), .B(n79997), .Z(n79998) );
  IV U100155 ( .A(n79998), .Z(n85688) );
  XOR U100156 ( .A(n85686), .B(n85688), .Z(n81312) );
  XOR U100157 ( .A(n81310), .B(n81312), .Z(n81314) );
  XOR U100158 ( .A(n81313), .B(n81314), .Z(n85696) );
  XOR U100159 ( .A(n85694), .B(n85696), .Z(n81306) );
  XOR U100160 ( .A(n81304), .B(n81306), .Z(n81309) );
  XOR U100161 ( .A(n79999), .B(n81309), .Z(n81297) );
  XOR U100162 ( .A(n81298), .B(n81297), .Z(n81296) );
  IV U100163 ( .A(n80000), .Z(n80002) );
  NOR U100164 ( .A(n80002), .B(n80001), .Z(n81294) );
  XOR U100165 ( .A(n81296), .B(n81294), .Z(n81292) );
  XOR U100166 ( .A(n81291), .B(n81292), .Z(n85705) );
  XOR U100167 ( .A(n85704), .B(n85705), .Z(n85712) );
  IV U100168 ( .A(n80003), .Z(n80004) );
  NOR U100169 ( .A(n80005), .B(n80004), .Z(n85711) );
  IV U100170 ( .A(n80006), .Z(n80008) );
  NOR U100171 ( .A(n80008), .B(n80007), .Z(n85707) );
  NOR U100172 ( .A(n85711), .B(n85707), .Z(n80009) );
  XOR U100173 ( .A(n85712), .B(n80009), .Z(n80010) );
  IV U100174 ( .A(n80010), .Z(n85715) );
  XOR U100175 ( .A(n85714), .B(n85715), .Z(n85723) );
  XOR U100176 ( .A(n85721), .B(n85723), .Z(n85720) );
  IV U100177 ( .A(n80011), .Z(n80013) );
  NOR U100178 ( .A(n80013), .B(n80012), .Z(n80014) );
  IV U100179 ( .A(n80014), .Z(n80021) );
  NOR U100180 ( .A(n85720), .B(n80021), .Z(n87070) );
  IV U100181 ( .A(n80015), .Z(n80020) );
  IV U100182 ( .A(n80016), .Z(n80017) );
  NOR U100183 ( .A(n80020), .B(n80017), .Z(n81288) );
  IV U100184 ( .A(n80018), .Z(n80019) );
  NOR U100185 ( .A(n80020), .B(n80019), .Z(n85718) );
  XOR U100186 ( .A(n85720), .B(n85718), .Z(n81289) );
  IV U100187 ( .A(n81289), .Z(n80022) );
  XOR U100188 ( .A(n81288), .B(n80022), .Z(n80024) );
  NOR U100189 ( .A(n80022), .B(n80021), .Z(n80023) );
  NOR U100190 ( .A(n80024), .B(n80023), .Z(n80025) );
  NOR U100191 ( .A(n87070), .B(n80025), .Z(n81279) );
  XOR U100192 ( .A(n81280), .B(n81279), .Z(n85742) );
  XOR U100193 ( .A(n80026), .B(n85742), .Z(n81276) );
  XOR U100194 ( .A(n80027), .B(n81276), .Z(n81273) );
  IV U100195 ( .A(n80028), .Z(n80029) );
  NOR U100196 ( .A(n80030), .B(n80029), .Z(n81268) );
  NOR U100197 ( .A(n81268), .B(n80033), .Z(n80031) );
  XOR U100198 ( .A(n81273), .B(n80031), .Z(n80032) );
  NOR U100199 ( .A(n80034), .B(n80032), .Z(n80037) );
  XOR U100200 ( .A(n80033), .B(n81273), .Z(n80036) );
  IV U100201 ( .A(n80034), .Z(n80035) );
  NOR U100202 ( .A(n80036), .B(n80035), .Z(n85753) );
  NOR U100203 ( .A(n80037), .B(n85753), .Z(n80038) );
  IV U100204 ( .A(n80038), .Z(n85751) );
  IV U100205 ( .A(n80039), .Z(n80041) );
  NOR U100206 ( .A(n80041), .B(n80040), .Z(n85750) );
  XOR U100207 ( .A(n85751), .B(n85750), .Z(n85762) );
  XOR U100208 ( .A(n81266), .B(n85762), .Z(n85759) );
  XOR U100209 ( .A(n85758), .B(n85759), .Z(n80042) );
  NOR U100210 ( .A(n80043), .B(n80042), .Z(n80044) );
  NOR U100211 ( .A(n80051), .B(n80044), .Z(n85771) );
  IV U100212 ( .A(n85771), .Z(n80050) );
  NOR U100213 ( .A(n80045), .B(n85763), .Z(n80047) );
  XOR U100214 ( .A(n85758), .B(n81266), .Z(n80046) );
  NOR U100215 ( .A(n80047), .B(n80046), .Z(n80048) );
  XOR U100216 ( .A(n80048), .B(n85762), .Z(n80053) );
  NOR U100217 ( .A(n80049), .B(n80053), .Z(n85772) );
  NOR U100218 ( .A(n80050), .B(n85772), .Z(n80055) );
  IV U100219 ( .A(n80051), .Z(n80052) );
  NOR U100220 ( .A(n80053), .B(n80052), .Z(n80054) );
  NOR U100221 ( .A(n80055), .B(n80054), .Z(n81265) );
  IV U100222 ( .A(n80056), .Z(n80057) );
  NOR U100223 ( .A(n80058), .B(n80057), .Z(n80059) );
  IV U100224 ( .A(n80059), .Z(n80063) );
  NOR U100225 ( .A(n81265), .B(n80063), .Z(n87016) );
  IV U100226 ( .A(n80060), .Z(n80062) );
  NOR U100227 ( .A(n80062), .B(n80061), .Z(n80064) );
  IV U100228 ( .A(n80064), .Z(n81264) );
  XOR U100229 ( .A(n81265), .B(n81264), .Z(n80066) );
  NOR U100230 ( .A(n80064), .B(n80063), .Z(n80065) );
  NOR U100231 ( .A(n80066), .B(n80065), .Z(n85774) );
  NOR U100232 ( .A(n87016), .B(n85774), .Z(n85780) );
  XOR U100233 ( .A(n87015), .B(n85780), .Z(n80067) );
  NOR U100234 ( .A(n80068), .B(n80067), .Z(n85790) );
  IV U100235 ( .A(n80069), .Z(n80070) );
  NOR U100236 ( .A(n80070), .B(n80072), .Z(n81260) );
  IV U100237 ( .A(n80071), .Z(n80073) );
  NOR U100238 ( .A(n80073), .B(n80072), .Z(n85779) );
  NOR U100239 ( .A(n85779), .B(n80074), .Z(n80075) );
  XOR U100240 ( .A(n85780), .B(n80075), .Z(n81261) );
  XOR U100241 ( .A(n81260), .B(n81261), .Z(n85788) );
  IV U100242 ( .A(n85788), .Z(n80076) );
  NOR U100243 ( .A(n80077), .B(n80076), .Z(n80078) );
  NOR U100244 ( .A(n85790), .B(n80078), .Z(n81257) );
  IV U100245 ( .A(n80079), .Z(n80080) );
  NOR U100246 ( .A(n80081), .B(n80080), .Z(n85786) );
  IV U100247 ( .A(n80082), .Z(n80083) );
  NOR U100248 ( .A(n80084), .B(n80083), .Z(n81256) );
  NOR U100249 ( .A(n85786), .B(n81256), .Z(n80085) );
  XOR U100250 ( .A(n81257), .B(n80085), .Z(n81255) );
  IV U100251 ( .A(n80086), .Z(n80088) );
  NOR U100252 ( .A(n80088), .B(n80087), .Z(n80089) );
  IV U100253 ( .A(n80089), .Z(n81254) );
  XOR U100254 ( .A(n81255), .B(n81254), .Z(n81247) );
  XOR U100255 ( .A(n81249), .B(n81247), .Z(n81238) );
  XOR U100256 ( .A(n80090), .B(n81238), .Z(n81227) );
  XOR U100257 ( .A(n81231), .B(n81227), .Z(n85796) );
  NOR U100258 ( .A(n80091), .B(n81228), .Z(n80095) );
  IV U100259 ( .A(n80092), .Z(n80094) );
  NOR U100260 ( .A(n80094), .B(n80093), .Z(n85795) );
  NOR U100261 ( .A(n80095), .B(n85795), .Z(n80096) );
  XOR U100262 ( .A(n85796), .B(n80096), .Z(n80097) );
  IV U100263 ( .A(n80097), .Z(n85809) );
  IV U100264 ( .A(n85803), .Z(n80098) );
  NOR U100265 ( .A(n80098), .B(n85799), .Z(n80100) );
  NOR U100266 ( .A(n85798), .B(n85802), .Z(n80099) );
  NOR U100267 ( .A(n80099), .B(n85799), .Z(n80105) );
  XOR U100268 ( .A(n80100), .B(n80105), .Z(n80107) );
  IV U100269 ( .A(n80101), .Z(n80103) );
  NOR U100270 ( .A(n80103), .B(n80102), .Z(n80104) );
  IV U100271 ( .A(n80104), .Z(n85808) );
  NOR U100272 ( .A(n80105), .B(n85808), .Z(n80106) );
  NOR U100273 ( .A(n80107), .B(n80106), .Z(n80108) );
  XOR U100274 ( .A(n85809), .B(n80108), .Z(n81219) );
  IV U100275 ( .A(n80109), .Z(n80111) );
  NOR U100276 ( .A(n80111), .B(n80110), .Z(n81222) );
  NOR U100277 ( .A(n80113), .B(n80112), .Z(n81220) );
  NOR U100278 ( .A(n81222), .B(n81220), .Z(n80114) );
  XOR U100279 ( .A(n81219), .B(n80114), .Z(n81208) );
  XOR U100280 ( .A(n81206), .B(n81208), .Z(n81211) );
  XOR U100281 ( .A(n81209), .B(n81211), .Z(n81216) );
  NOR U100282 ( .A(n80120), .B(n81216), .Z(n86989) );
  IV U100283 ( .A(n80115), .Z(n80116) );
  NOR U100284 ( .A(n80116), .B(n80126), .Z(n81203) );
  IV U100285 ( .A(n80117), .Z(n80118) );
  NOR U100286 ( .A(n80119), .B(n80118), .Z(n81215) );
  XOR U100287 ( .A(n81215), .B(n81216), .Z(n81204) );
  IV U100288 ( .A(n81204), .Z(n80121) );
  XOR U100289 ( .A(n81203), .B(n80121), .Z(n80123) );
  NOR U100290 ( .A(n80121), .B(n80120), .Z(n80122) );
  NOR U100291 ( .A(n80123), .B(n80122), .Z(n80124) );
  NOR U100292 ( .A(n86989), .B(n80124), .Z(n81195) );
  IV U100293 ( .A(n80125), .Z(n80127) );
  NOR U100294 ( .A(n80127), .B(n80126), .Z(n80128) );
  IV U100295 ( .A(n80128), .Z(n81197) );
  XOR U100296 ( .A(n81195), .B(n81197), .Z(n81199) );
  XOR U100297 ( .A(n81198), .B(n81199), .Z(n81190) );
  XOR U100298 ( .A(n81191), .B(n81190), .Z(n80129) );
  IV U100299 ( .A(n80129), .Z(n81193) );
  XOR U100300 ( .A(n81192), .B(n81193), .Z(n85817) );
  IV U100301 ( .A(n80130), .Z(n80132) );
  NOR U100302 ( .A(n80132), .B(n80131), .Z(n85816) );
  IV U100303 ( .A(n80133), .Z(n80135) );
  NOR U100304 ( .A(n80135), .B(n80134), .Z(n85814) );
  NOR U100305 ( .A(n85816), .B(n85814), .Z(n80136) );
  IV U100306 ( .A(n80136), .Z(n80137) );
  NOR U100307 ( .A(n81188), .B(n80137), .Z(n80138) );
  XOR U100308 ( .A(n85817), .B(n80138), .Z(n80139) );
  IV U100309 ( .A(n80139), .Z(n81184) );
  IV U100310 ( .A(n80140), .Z(n80142) );
  NOR U100311 ( .A(n80142), .B(n80141), .Z(n80143) );
  NOR U100312 ( .A(n80144), .B(n80143), .Z(n81183) );
  XOR U100313 ( .A(n81184), .B(n81183), .Z(n81185) );
  IV U100314 ( .A(n80145), .Z(n80146) );
  NOR U100315 ( .A(n80147), .B(n80146), .Z(n85829) );
  IV U100316 ( .A(n80148), .Z(n80151) );
  IV U100317 ( .A(n80149), .Z(n80150) );
  NOR U100318 ( .A(n80151), .B(n80150), .Z(n81186) );
  NOR U100319 ( .A(n85829), .B(n81186), .Z(n80152) );
  XOR U100320 ( .A(n81185), .B(n80152), .Z(n85834) );
  XOR U100321 ( .A(n85832), .B(n85834), .Z(n85842) );
  XOR U100322 ( .A(n81180), .B(n85842), .Z(n80153) );
  XOR U100323 ( .A(n80154), .B(n80153), .Z(n85838) );
  IV U100324 ( .A(n80155), .Z(n80157) );
  NOR U100325 ( .A(n80157), .B(n80156), .Z(n80158) );
  NOR U100326 ( .A(n80159), .B(n80158), .Z(n85840) );
  XOR U100327 ( .A(n85838), .B(n85840), .Z(n81178) );
  XOR U100328 ( .A(n81177), .B(n81178), .Z(n85866) );
  XOR U100329 ( .A(n80160), .B(n85866), .Z(n80161) );
  IV U100330 ( .A(n80161), .Z(n85863) );
  XOR U100331 ( .A(n85861), .B(n85863), .Z(n81171) );
  IV U100332 ( .A(n81171), .Z(n81168) );
  IV U100333 ( .A(n80162), .Z(n80164) );
  NOR U100334 ( .A(n80164), .B(n80163), .Z(n81173) );
  IV U100335 ( .A(n80165), .Z(n80167) );
  NOR U100336 ( .A(n80167), .B(n80166), .Z(n81169) );
  NOR U100337 ( .A(n81173), .B(n81169), .Z(n80168) );
  XOR U100338 ( .A(n81168), .B(n80168), .Z(n81167) );
  XOR U100339 ( .A(n81163), .B(n81167), .Z(n80169) );
  XOR U100340 ( .A(n80170), .B(n80169), .Z(n80171) );
  XOR U100341 ( .A(n81155), .B(n80171), .Z(n81158) );
  XOR U100342 ( .A(n81159), .B(n81158), .Z(n85889) );
  IV U100343 ( .A(n80172), .Z(n80173) );
  NOR U100344 ( .A(n80174), .B(n80173), .Z(n81160) );
  NOR U100345 ( .A(n80175), .B(n80179), .Z(n85887) );
  NOR U100346 ( .A(n81160), .B(n85887), .Z(n80176) );
  XOR U100347 ( .A(n85889), .B(n80176), .Z(n80177) );
  IV U100348 ( .A(n80177), .Z(n85886) );
  IV U100349 ( .A(n80178), .Z(n80180) );
  NOR U100350 ( .A(n80180), .B(n80179), .Z(n85884) );
  XOR U100351 ( .A(n85886), .B(n85884), .Z(n81153) );
  XOR U100352 ( .A(n81152), .B(n81153), .Z(n85894) );
  XOR U100353 ( .A(n80181), .B(n85894), .Z(n80189) );
  IV U100354 ( .A(n80189), .Z(n80182) );
  NOR U100355 ( .A(n80183), .B(n80182), .Z(n91707) );
  IV U100356 ( .A(n80184), .Z(n80185) );
  NOR U100357 ( .A(n80186), .B(n80185), .Z(n80190) );
  IV U100358 ( .A(n80190), .Z(n80188) );
  XOR U100359 ( .A(n85892), .B(n85894), .Z(n80187) );
  NOR U100360 ( .A(n80188), .B(n80187), .Z(n91702) );
  NOR U100361 ( .A(n80190), .B(n80189), .Z(n80191) );
  NOR U100362 ( .A(n91702), .B(n80191), .Z(n80196) );
  NOR U100363 ( .A(n80192), .B(n80196), .Z(n80193) );
  NOR U100364 ( .A(n91707), .B(n80193), .Z(n80194) );
  NOR U100365 ( .A(n80195), .B(n80194), .Z(n80199) );
  IV U100366 ( .A(n80195), .Z(n80198) );
  IV U100367 ( .A(n80196), .Z(n80197) );
  NOR U100368 ( .A(n80198), .B(n80197), .Z(n91706) );
  NOR U100369 ( .A(n80199), .B(n91706), .Z(n80200) );
  IV U100370 ( .A(n80200), .Z(n85905) );
  IV U100371 ( .A(n80201), .Z(n80203) );
  NOR U100372 ( .A(n80203), .B(n80202), .Z(n85904) );
  IV U100373 ( .A(n80204), .Z(n80206) );
  NOR U100374 ( .A(n80206), .B(n80205), .Z(n81150) );
  NOR U100375 ( .A(n85904), .B(n81150), .Z(n80207) );
  XOR U100376 ( .A(n85905), .B(n80207), .Z(n81143) );
  XOR U100377 ( .A(n81144), .B(n81143), .Z(n81140) );
  XOR U100378 ( .A(n80208), .B(n81140), .Z(n81134) );
  XOR U100379 ( .A(n81136), .B(n81134), .Z(n81137) );
  XOR U100380 ( .A(n81138), .B(n81137), .Z(n80211) );
  IV U100381 ( .A(n80211), .Z(n80209) );
  NOR U100382 ( .A(n80210), .B(n80209), .Z(n86888) );
  NOR U100383 ( .A(n80212), .B(n80211), .Z(n81130) );
  IV U100384 ( .A(n80213), .Z(n80214) );
  NOR U100385 ( .A(n80218), .B(n80214), .Z(n81128) );
  XOR U100386 ( .A(n81130), .B(n81128), .Z(n80215) );
  NOR U100387 ( .A(n86888), .B(n80215), .Z(n81126) );
  IV U100388 ( .A(n80216), .Z(n80217) );
  NOR U100389 ( .A(n80218), .B(n80217), .Z(n81131) );
  NOR U100390 ( .A(n80220), .B(n80219), .Z(n81125) );
  NOR U100391 ( .A(n81131), .B(n81125), .Z(n80221) );
  XOR U100392 ( .A(n81126), .B(n80221), .Z(n81123) );
  IV U100393 ( .A(n80222), .Z(n80226) );
  NOR U100394 ( .A(n80224), .B(n80223), .Z(n80225) );
  IV U100395 ( .A(n80225), .Z(n80230) );
  NOR U100396 ( .A(n80226), .B(n80230), .Z(n81119) );
  NOR U100397 ( .A(n81121), .B(n81119), .Z(n80227) );
  XOR U100398 ( .A(n81123), .B(n80227), .Z(n80228) );
  IV U100399 ( .A(n80228), .Z(n81116) );
  IV U100400 ( .A(n80229), .Z(n80231) );
  NOR U100401 ( .A(n80231), .B(n80230), .Z(n81114) );
  XOR U100402 ( .A(n81116), .B(n81114), .Z(n85918) );
  XOR U100403 ( .A(n81117), .B(n85918), .Z(n81111) );
  NOR U100404 ( .A(n81110), .B(n85917), .Z(n80232) );
  XOR U100405 ( .A(n81111), .B(n80232), .Z(n80233) );
  IV U100406 ( .A(n80233), .Z(n85923) );
  IV U100407 ( .A(n80234), .Z(n80236) );
  NOR U100408 ( .A(n80236), .B(n80235), .Z(n80240) );
  IV U100409 ( .A(n80240), .Z(n80237) );
  NOR U100410 ( .A(n85923), .B(n80237), .Z(n86857) );
  XOR U100411 ( .A(n80238), .B(n85923), .Z(n81108) );
  IV U100412 ( .A(n81108), .Z(n80239) );
  NOR U100413 ( .A(n80240), .B(n80239), .Z(n80241) );
  NOR U100414 ( .A(n86857), .B(n80241), .Z(n81101) );
  XOR U100415 ( .A(n80242), .B(n81101), .Z(n81100) );
  XOR U100416 ( .A(n81098), .B(n81100), .Z(n85928) );
  IV U100417 ( .A(n80243), .Z(n80244) );
  NOR U100418 ( .A(n80245), .B(n80244), .Z(n80250) );
  IV U100419 ( .A(n80246), .Z(n80247) );
  NOR U100420 ( .A(n80248), .B(n80247), .Z(n80249) );
  NOR U100421 ( .A(n80250), .B(n80249), .Z(n85929) );
  IV U100422 ( .A(n85929), .Z(n85926) );
  XOR U100423 ( .A(n85928), .B(n85926), .Z(n85935) );
  XOR U100424 ( .A(n80251), .B(n85935), .Z(n81089) );
  XOR U100425 ( .A(n80252), .B(n81089), .Z(n81085) );
  XOR U100426 ( .A(n81083), .B(n81085), .Z(n81087) );
  XOR U100427 ( .A(n80253), .B(n81087), .Z(n81077) );
  XOR U100428 ( .A(n81078), .B(n81077), .Z(n81071) );
  IV U100429 ( .A(n80254), .Z(n80256) );
  NOR U100430 ( .A(n80256), .B(n80255), .Z(n81069) );
  XOR U100431 ( .A(n81071), .B(n81069), .Z(n81073) );
  XOR U100432 ( .A(n81072), .B(n81073), .Z(n85945) );
  XOR U100433 ( .A(n81066), .B(n85945), .Z(n81062) );
  IV U100434 ( .A(n80257), .Z(n80258) );
  NOR U100435 ( .A(n80259), .B(n80258), .Z(n80260) );
  NOR U100436 ( .A(n85944), .B(n80260), .Z(n81063) );
  XOR U100437 ( .A(n81062), .B(n81063), .Z(n85951) );
  XOR U100438 ( .A(n85952), .B(n85951), .Z(n85955) );
  IV U100439 ( .A(n80261), .Z(n80262) );
  NOR U100440 ( .A(n80263), .B(n80262), .Z(n85954) );
  IV U100441 ( .A(n80264), .Z(n80265) );
  NOR U100442 ( .A(n80266), .B(n80265), .Z(n81060) );
  NOR U100443 ( .A(n85954), .B(n81060), .Z(n80267) );
  XOR U100444 ( .A(n85955), .B(n80267), .Z(n80268) );
  NOR U100445 ( .A(n80269), .B(n80268), .Z(n80272) );
  IV U100446 ( .A(n80269), .Z(n80271) );
  XOR U100447 ( .A(n85954), .B(n85955), .Z(n80270) );
  NOR U100448 ( .A(n80271), .B(n80270), .Z(n86752) );
  NOR U100449 ( .A(n80272), .B(n86752), .Z(n81053) );
  XOR U100450 ( .A(n81052), .B(n81053), .Z(n81050) );
  XOR U100451 ( .A(n80273), .B(n81050), .Z(n85970) );
  XOR U100452 ( .A(n85978), .B(n85970), .Z(n85964) );
  NOR U100453 ( .A(n80274), .B(n85971), .Z(n80278) );
  IV U100454 ( .A(n80275), .Z(n80276) );
  NOR U100455 ( .A(n80277), .B(n80276), .Z(n81044) );
  XOR U100456 ( .A(n80278), .B(n81044), .Z(n80284) );
  IV U100457 ( .A(n80279), .Z(n85965) );
  NOR U100458 ( .A(n80280), .B(n85965), .Z(n80281) );
  IV U100459 ( .A(n80281), .Z(n80282) );
  NOR U100460 ( .A(n81044), .B(n80282), .Z(n80283) );
  NOR U100461 ( .A(n80284), .B(n80283), .Z(n80285) );
  XOR U100462 ( .A(n85964), .B(n80285), .Z(n80286) );
  IV U100463 ( .A(n80286), .Z(n81042) );
  IV U100464 ( .A(n80287), .Z(n80289) );
  NOR U100465 ( .A(n80289), .B(n80288), .Z(n80290) );
  IV U100466 ( .A(n80290), .Z(n81037) );
  XOR U100467 ( .A(n81042), .B(n81037), .Z(n80291) );
  XOR U100468 ( .A(n80292), .B(n80291), .Z(n81035) );
  XOR U100469 ( .A(n80293), .B(n81035), .Z(n81025) );
  XOR U100470 ( .A(n81026), .B(n81025), .Z(n81029) );
  XOR U100471 ( .A(n81028), .B(n81029), .Z(n81022) );
  XOR U100472 ( .A(n81023), .B(n81022), .Z(n80300) );
  IV U100473 ( .A(n80300), .Z(n80294) );
  NOR U100474 ( .A(n80295), .B(n80294), .Z(n81021) );
  IV U100475 ( .A(n80296), .Z(n80298) );
  NOR U100476 ( .A(n80298), .B(n80297), .Z(n80301) );
  IV U100477 ( .A(n80301), .Z(n80299) );
  NOR U100478 ( .A(n80299), .B(n81029), .Z(n91752) );
  NOR U100479 ( .A(n80301), .B(n80300), .Z(n80302) );
  NOR U100480 ( .A(n91752), .B(n80302), .Z(n81014) );
  NOR U100481 ( .A(n80303), .B(n81014), .Z(n80304) );
  NOR U100482 ( .A(n81021), .B(n80304), .Z(n81017) );
  IV U100483 ( .A(n80305), .Z(n80307) );
  NOR U100484 ( .A(n80307), .B(n80306), .Z(n80308) );
  IV U100485 ( .A(n80308), .Z(n81018) );
  XOR U100486 ( .A(n81017), .B(n81018), .Z(n85991) );
  XOR U100487 ( .A(n81016), .B(n85991), .Z(n81011) );
  IV U100488 ( .A(n80309), .Z(n80310) );
  NOR U100489 ( .A(n80311), .B(n80310), .Z(n85990) );
  IV U100490 ( .A(n80312), .Z(n80314) );
  NOR U100491 ( .A(n80314), .B(n80313), .Z(n81010) );
  NOR U100492 ( .A(n85990), .B(n81010), .Z(n80315) );
  XOR U100493 ( .A(n81011), .B(n80315), .Z(n81009) );
  IV U100494 ( .A(n80316), .Z(n80317) );
  NOR U100495 ( .A(n80318), .B(n80317), .Z(n81001) );
  NOR U100496 ( .A(n81007), .B(n81001), .Z(n80319) );
  XOR U100497 ( .A(n81009), .B(n80319), .Z(n81004) );
  IV U100498 ( .A(n80320), .Z(n80321) );
  NOR U100499 ( .A(n80321), .B(n80328), .Z(n81003) );
  IV U100500 ( .A(n80322), .Z(n80324) );
  NOR U100501 ( .A(n80324), .B(n80323), .Z(n80997) );
  NOR U100502 ( .A(n81003), .B(n80997), .Z(n80325) );
  XOR U100503 ( .A(n81004), .B(n80325), .Z(n80991) );
  IV U100504 ( .A(n80326), .Z(n80327) );
  NOR U100505 ( .A(n80328), .B(n80327), .Z(n80989) );
  XOR U100506 ( .A(n80991), .B(n80989), .Z(n80993) );
  IV U100507 ( .A(n80329), .Z(n80330) );
  NOR U100508 ( .A(n80331), .B(n80330), .Z(n80992) );
  IV U100509 ( .A(n80332), .Z(n80334) );
  NOR U100510 ( .A(n80334), .B(n80333), .Z(n80987) );
  NOR U100511 ( .A(n80992), .B(n80987), .Z(n80335) );
  XOR U100512 ( .A(n80993), .B(n80335), .Z(n80336) );
  NOR U100513 ( .A(n80337), .B(n80336), .Z(n80340) );
  IV U100514 ( .A(n80337), .Z(n80339) );
  XOR U100515 ( .A(n80992), .B(n80993), .Z(n80338) );
  NOR U100516 ( .A(n80339), .B(n80338), .Z(n80986) );
  NOR U100517 ( .A(n80340), .B(n80986), .Z(n80983) );
  XOR U100518 ( .A(n80984), .B(n80983), .Z(n80982) );
  XOR U100519 ( .A(n80980), .B(n80982), .Z(n80979) );
  XOR U100520 ( .A(n80341), .B(n80979), .Z(n80976) );
  XOR U100521 ( .A(n80974), .B(n80976), .Z(n80971) );
  IV U100522 ( .A(n80342), .Z(n80343) );
  NOR U100523 ( .A(n80343), .B(n80345), .Z(n80969) );
  XOR U100524 ( .A(n80971), .B(n80969), .Z(n86005) );
  IV U100525 ( .A(n80344), .Z(n80346) );
  NOR U100526 ( .A(n80346), .B(n80345), .Z(n80972) );
  XOR U100527 ( .A(n86005), .B(n80972), .Z(n80968) );
  IV U100528 ( .A(n80347), .Z(n80351) );
  NOR U100529 ( .A(n80351), .B(n80348), .Z(n86004) );
  IV U100530 ( .A(n80349), .Z(n80350) );
  NOR U100531 ( .A(n80351), .B(n80350), .Z(n80966) );
  NOR U100532 ( .A(n86004), .B(n80966), .Z(n80352) );
  XOR U100533 ( .A(n80968), .B(n80352), .Z(n80353) );
  IV U100534 ( .A(n80353), .Z(n86009) );
  IV U100535 ( .A(n80354), .Z(n80356) );
  NOR U100536 ( .A(n80356), .B(n80355), .Z(n86007) );
  XOR U100537 ( .A(n86009), .B(n86007), .Z(n86012) );
  XOR U100538 ( .A(n86010), .B(n86012), .Z(n80964) );
  XOR U100539 ( .A(n80963), .B(n80964), .Z(n86017) );
  XOR U100540 ( .A(n86015), .B(n86017), .Z(n86020) );
  XOR U100541 ( .A(n86018), .B(n86020), .Z(n80961) );
  XOR U100542 ( .A(n80960), .B(n80961), .Z(n86035) );
  XOR U100543 ( .A(n80357), .B(n86035), .Z(n86037) );
  XOR U100544 ( .A(n80358), .B(n86037), .Z(n86049) );
  XOR U100545 ( .A(n86047), .B(n86049), .Z(n86053) );
  XOR U100546 ( .A(n80359), .B(n86053), .Z(n80949) );
  XOR U100547 ( .A(n80950), .B(n80949), .Z(n80953) );
  XOR U100548 ( .A(n80952), .B(n80953), .Z(n80366) );
  IV U100549 ( .A(n80366), .Z(n80360) );
  NOR U100550 ( .A(n80361), .B(n80360), .Z(n91851) );
  IV U100551 ( .A(n80362), .Z(n80364) );
  NOR U100552 ( .A(n80364), .B(n80363), .Z(n80367) );
  IV U100553 ( .A(n80367), .Z(n80365) );
  NOR U100554 ( .A(n80365), .B(n80953), .Z(n91848) );
  NOR U100555 ( .A(n80367), .B(n80366), .Z(n80368) );
  NOR U100556 ( .A(n91848), .B(n80368), .Z(n80946) );
  NOR U100557 ( .A(n80369), .B(n80946), .Z(n80370) );
  NOR U100558 ( .A(n91851), .B(n80370), .Z(n80371) );
  XOR U100559 ( .A(n80948), .B(n80371), .Z(n80943) );
  IV U100560 ( .A(n80372), .Z(n80374) );
  IV U100561 ( .A(n80373), .Z(n80379) );
  NOR U100562 ( .A(n80374), .B(n80379), .Z(n80940) );
  NOR U100563 ( .A(n80942), .B(n80940), .Z(n80375) );
  XOR U100564 ( .A(n80943), .B(n80375), .Z(n80933) );
  IV U100565 ( .A(n80376), .Z(n80377) );
  NOR U100566 ( .A(n80384), .B(n80377), .Z(n80934) );
  IV U100567 ( .A(n80378), .Z(n80380) );
  NOR U100568 ( .A(n80380), .B(n80379), .Z(n80937) );
  NOR U100569 ( .A(n80934), .B(n80937), .Z(n80381) );
  XOR U100570 ( .A(n80933), .B(n80381), .Z(n86059) );
  IV U100571 ( .A(n80382), .Z(n80383) );
  NOR U100572 ( .A(n80384), .B(n80383), .Z(n86057) );
  XOR U100573 ( .A(n86059), .B(n86057), .Z(n86061) );
  XOR U100574 ( .A(n86060), .B(n86061), .Z(n80931) );
  XOR U100575 ( .A(n80930), .B(n80931), .Z(n86070) );
  IV U100576 ( .A(n86070), .Z(n86072) );
  IV U100577 ( .A(n80385), .Z(n80387) );
  NOR U100578 ( .A(n80387), .B(n80386), .Z(n86071) );
  IV U100579 ( .A(n86071), .Z(n86069) );
  XOR U100580 ( .A(n86072), .B(n86069), .Z(n80928) );
  IV U100581 ( .A(n80388), .Z(n80389) );
  NOR U100582 ( .A(n80390), .B(n80389), .Z(n86073) );
  IV U100583 ( .A(n80391), .Z(n80393) );
  NOR U100584 ( .A(n80393), .B(n80392), .Z(n80927) );
  NOR U100585 ( .A(n86073), .B(n80927), .Z(n80394) );
  XOR U100586 ( .A(n80928), .B(n80394), .Z(n80923) );
  XOR U100587 ( .A(n86080), .B(n80923), .Z(n80395) );
  XOR U100588 ( .A(n80396), .B(n80395), .Z(n86098) );
  IV U100589 ( .A(n80397), .Z(n80399) );
  NOR U100590 ( .A(n80399), .B(n80398), .Z(n86096) );
  XOR U100591 ( .A(n86098), .B(n86096), .Z(n86099) );
  XOR U100592 ( .A(n86100), .B(n86099), .Z(n80916) );
  XOR U100593 ( .A(n80915), .B(n80916), .Z(n80912) );
  XOR U100594 ( .A(n80400), .B(n80912), .Z(n80908) );
  XOR U100595 ( .A(n80401), .B(n80908), .Z(n80906) );
  XOR U100596 ( .A(n80402), .B(n80906), .Z(n86106) );
  NOR U100597 ( .A(n80403), .B(n86107), .Z(n86119) );
  IV U100598 ( .A(n80404), .Z(n80405) );
  NOR U100599 ( .A(n80408), .B(n80405), .Z(n86113) );
  IV U100600 ( .A(n80406), .Z(n80407) );
  NOR U100601 ( .A(n80408), .B(n80407), .Z(n80409) );
  NOR U100602 ( .A(n86113), .B(n80409), .Z(n80410) );
  IV U100603 ( .A(n80410), .Z(n80411) );
  NOR U100604 ( .A(n86119), .B(n80411), .Z(n80412) );
  XOR U100605 ( .A(n86106), .B(n80412), .Z(n80901) );
  XOR U100606 ( .A(n80413), .B(n80901), .Z(n86129) );
  IV U100607 ( .A(n86129), .Z(n80421) );
  IV U100608 ( .A(n80414), .Z(n80416) );
  NOR U100609 ( .A(n80416), .B(n80415), .Z(n80900) );
  IV U100610 ( .A(n80417), .Z(n80418) );
  NOR U100611 ( .A(n80419), .B(n80418), .Z(n86128) );
  NOR U100612 ( .A(n80900), .B(n86128), .Z(n80420) );
  XOR U100613 ( .A(n80421), .B(n80420), .Z(n86133) );
  XOR U100614 ( .A(n80422), .B(n86133), .Z(n86145) );
  XOR U100615 ( .A(n86150), .B(n86145), .Z(n80895) );
  XOR U100616 ( .A(n80896), .B(n80895), .Z(n80884) );
  XOR U100617 ( .A(n80889), .B(n80884), .Z(n80882) );
  IV U100618 ( .A(n80423), .Z(n80885) );
  NOR U100619 ( .A(n80424), .B(n80885), .Z(n80427) );
  IV U100620 ( .A(n80425), .Z(n80426) );
  NOR U100621 ( .A(n80426), .B(n80433), .Z(n80880) );
  NOR U100622 ( .A(n80427), .B(n80880), .Z(n80428) );
  XOR U100623 ( .A(n80882), .B(n80428), .Z(n80870) );
  IV U100624 ( .A(n80429), .Z(n80430) );
  NOR U100625 ( .A(n80431), .B(n80430), .Z(n80871) );
  IV U100626 ( .A(n80432), .Z(n80434) );
  NOR U100627 ( .A(n80434), .B(n80433), .Z(n80877) );
  NOR U100628 ( .A(n80871), .B(n80877), .Z(n80435) );
  XOR U100629 ( .A(n80870), .B(n80435), .Z(n86158) );
  IV U100630 ( .A(n86158), .Z(n86160) );
  XOR U100631 ( .A(n86161), .B(n86160), .Z(n80436) );
  XOR U100632 ( .A(n80437), .B(n80436), .Z(n86157) );
  IV U100633 ( .A(n80438), .Z(n80441) );
  IV U100634 ( .A(n80439), .Z(n80440) );
  NOR U100635 ( .A(n80441), .B(n80440), .Z(n86155) );
  XOR U100636 ( .A(n86157), .B(n86155), .Z(n80866) );
  XOR U100637 ( .A(n80864), .B(n80866), .Z(n80868) );
  XOR U100638 ( .A(n80867), .B(n80868), .Z(n80862) );
  XOR U100639 ( .A(n80861), .B(n80862), .Z(n86170) );
  XOR U100640 ( .A(n86169), .B(n86170), .Z(n86173) );
  XOR U100641 ( .A(n86172), .B(n86173), .Z(n86190) );
  XOR U100642 ( .A(n80442), .B(n86190), .Z(n86193) );
  IV U100643 ( .A(n80443), .Z(n80444) );
  NOR U100644 ( .A(n80445), .B(n80444), .Z(n86192) );
  NOR U100645 ( .A(n86198), .B(n86192), .Z(n80446) );
  XOR U100646 ( .A(n86193), .B(n80446), .Z(n80853) );
  XOR U100647 ( .A(n80447), .B(n80853), .Z(n80842) );
  XOR U100648 ( .A(n80448), .B(n80842), .Z(n86208) );
  XOR U100649 ( .A(n86206), .B(n86208), .Z(n86202) );
  IV U100650 ( .A(n80449), .Z(n80451) );
  IV U100651 ( .A(n80450), .Z(n80461) );
  NOR U100652 ( .A(n80451), .B(n80461), .Z(n80837) );
  IV U100653 ( .A(n80452), .Z(n80453) );
  NOR U100654 ( .A(n80454), .B(n80453), .Z(n80839) );
  NOR U100655 ( .A(n86201), .B(n80839), .Z(n80455) );
  IV U100656 ( .A(n80455), .Z(n80456) );
  NOR U100657 ( .A(n80837), .B(n80456), .Z(n80457) );
  XOR U100658 ( .A(n86202), .B(n80457), .Z(n80831) );
  IV U100659 ( .A(n80458), .Z(n80459) );
  NOR U100660 ( .A(n80466), .B(n80459), .Z(n80832) );
  IV U100661 ( .A(n80460), .Z(n80462) );
  NOR U100662 ( .A(n80462), .B(n80461), .Z(n80835) );
  NOR U100663 ( .A(n80832), .B(n80835), .Z(n80463) );
  XOR U100664 ( .A(n80831), .B(n80463), .Z(n80829) );
  IV U100665 ( .A(n80464), .Z(n80465) );
  NOR U100666 ( .A(n80466), .B(n80465), .Z(n80828) );
  IV U100667 ( .A(n80467), .Z(n80468) );
  NOR U100668 ( .A(n80468), .B(n80471), .Z(n80824) );
  NOR U100669 ( .A(n80828), .B(n80824), .Z(n80469) );
  XOR U100670 ( .A(n80829), .B(n80469), .Z(n80819) );
  IV U100671 ( .A(n80470), .Z(n80474) );
  NOR U100672 ( .A(n80472), .B(n80471), .Z(n80473) );
  IV U100673 ( .A(n80473), .Z(n80476) );
  NOR U100674 ( .A(n80474), .B(n80476), .Z(n80821) );
  IV U100675 ( .A(n80475), .Z(n80477) );
  NOR U100676 ( .A(n80477), .B(n80476), .Z(n80478) );
  IV U100677 ( .A(n80478), .Z(n80820) );
  XOR U100678 ( .A(n80821), .B(n80820), .Z(n80479) );
  XOR U100679 ( .A(n80819), .B(n80479), .Z(n80817) );
  XOR U100680 ( .A(n80816), .B(n80817), .Z(n80486) );
  IV U100681 ( .A(n80486), .Z(n80480) );
  NOR U100682 ( .A(n80485), .B(n80480), .Z(n80490) );
  IV U100683 ( .A(n80490), .Z(n80484) );
  IV U100684 ( .A(n80481), .Z(n80482) );
  NOR U100685 ( .A(n80483), .B(n80482), .Z(n80488) );
  NOR U100686 ( .A(n80484), .B(n80488), .Z(n80492) );
  IV U100687 ( .A(n80485), .Z(n80487) );
  NOR U100688 ( .A(n80487), .B(n80486), .Z(n86520) );
  IV U100689 ( .A(n80488), .Z(n80489) );
  NOR U100690 ( .A(n80490), .B(n80489), .Z(n86489) );
  NOR U100691 ( .A(n86520), .B(n86489), .Z(n80491) );
  IV U100692 ( .A(n80491), .Z(n91944) );
  NOR U100693 ( .A(n80492), .B(n91944), .Z(n86216) );
  NOR U100694 ( .A(n80495), .B(n80493), .Z(n86215) );
  IV U100695 ( .A(n80494), .Z(n80498) );
  NOR U100696 ( .A(n80496), .B(n80495), .Z(n80497) );
  IV U100697 ( .A(n80497), .Z(n80501) );
  NOR U100698 ( .A(n80498), .B(n80501), .Z(n86223) );
  NOR U100699 ( .A(n86215), .B(n86223), .Z(n80499) );
  XOR U100700 ( .A(n86216), .B(n80499), .Z(n86222) );
  IV U100701 ( .A(n80500), .Z(n80502) );
  NOR U100702 ( .A(n80502), .B(n80501), .Z(n86220) );
  XOR U100703 ( .A(n86222), .B(n86220), .Z(n86232) );
  XOR U100704 ( .A(n80814), .B(n86232), .Z(n80812) );
  XOR U100705 ( .A(n80503), .B(n80812), .Z(n80806) );
  XOR U100706 ( .A(n80504), .B(n80806), .Z(n80804) );
  XOR U100707 ( .A(n80505), .B(n80804), .Z(n80796) );
  IV U100708 ( .A(n80796), .Z(n80795) );
  XOR U100709 ( .A(n80797), .B(n80795), .Z(n80793) );
  IV U100710 ( .A(n80506), .Z(n80508) );
  NOR U100711 ( .A(n80508), .B(n80507), .Z(n80798) );
  IV U100712 ( .A(n80509), .Z(n80511) );
  IV U100713 ( .A(n80510), .Z(n80514) );
  NOR U100714 ( .A(n80511), .B(n80514), .Z(n80791) );
  NOR U100715 ( .A(n80798), .B(n80791), .Z(n80512) );
  XOR U100716 ( .A(n80793), .B(n80512), .Z(n86252) );
  IV U100717 ( .A(n80513), .Z(n80515) );
  NOR U100718 ( .A(n80515), .B(n80514), .Z(n80516) );
  IV U100719 ( .A(n80516), .Z(n86253) );
  XOR U100720 ( .A(n86252), .B(n86253), .Z(n86257) );
  XOR U100721 ( .A(n86255), .B(n86257), .Z(n80789) );
  XOR U100722 ( .A(n80517), .B(n80789), .Z(n80518) );
  IV U100723 ( .A(n80518), .Z(n80779) );
  XOR U100724 ( .A(n80778), .B(n80779), .Z(n80782) );
  XOR U100725 ( .A(n80781), .B(n80782), .Z(n86265) );
  IV U100726 ( .A(n86265), .Z(n80526) );
  IV U100727 ( .A(n80519), .Z(n80520) );
  NOR U100728 ( .A(n80521), .B(n80520), .Z(n86264) );
  IV U100729 ( .A(n80522), .Z(n80524) );
  NOR U100730 ( .A(n80524), .B(n80523), .Z(n86260) );
  NOR U100731 ( .A(n86264), .B(n86260), .Z(n80525) );
  XOR U100732 ( .A(n80526), .B(n80525), .Z(n86276) );
  XOR U100733 ( .A(n86274), .B(n86276), .Z(n80527) );
  XOR U100734 ( .A(n80528), .B(n80527), .Z(n80529) );
  IV U100735 ( .A(n80529), .Z(n80775) );
  XOR U100736 ( .A(n80530), .B(n80775), .Z(n80766) );
  XOR U100737 ( .A(n80531), .B(n80766), .Z(n80752) );
  XOR U100738 ( .A(n80532), .B(n80752), .Z(n80746) );
  XOR U100739 ( .A(n80744), .B(n80746), .Z(n80747) );
  IV U100740 ( .A(n80533), .Z(n80534) );
  NOR U100741 ( .A(n80535), .B(n80534), .Z(n80542) );
  IV U100742 ( .A(n80542), .Z(n80748) );
  XOR U100743 ( .A(n80747), .B(n80748), .Z(n80536) );
  NOR U100744 ( .A(n80740), .B(n80536), .Z(n80541) );
  IV U100745 ( .A(n80537), .Z(n80539) );
  NOR U100746 ( .A(n80539), .B(n80538), .Z(n80544) );
  IV U100747 ( .A(n80544), .Z(n80540) );
  NOR U100748 ( .A(n80541), .B(n80540), .Z(n80742) );
  NOR U100749 ( .A(n80542), .B(n80740), .Z(n80543) );
  XOR U100750 ( .A(n80543), .B(n80747), .Z(n80734) );
  NOR U100751 ( .A(n80544), .B(n80734), .Z(n80545) );
  NOR U100752 ( .A(n80742), .B(n80545), .Z(n80730) );
  NOR U100753 ( .A(n80546), .B(n80736), .Z(n80550) );
  IV U100754 ( .A(n80547), .Z(n80548) );
  NOR U100755 ( .A(n80549), .B(n80548), .Z(n80729) );
  NOR U100756 ( .A(n80550), .B(n80729), .Z(n80551) );
  XOR U100757 ( .A(n80730), .B(n80551), .Z(n80728) );
  IV U100758 ( .A(n80552), .Z(n80553) );
  NOR U100759 ( .A(n80553), .B(n80555), .Z(n80724) );
  IV U100760 ( .A(n80554), .Z(n80556) );
  NOR U100761 ( .A(n80556), .B(n80555), .Z(n80726) );
  NOR U100762 ( .A(n80724), .B(n80726), .Z(n80557) );
  XOR U100763 ( .A(n80728), .B(n80557), .Z(n80722) );
  IV U100764 ( .A(n80558), .Z(n80564) );
  IV U100765 ( .A(n80559), .Z(n80560) );
  NOR U100766 ( .A(n80564), .B(n80560), .Z(n80721) );
  NOR U100767 ( .A(n86290), .B(n80721), .Z(n80561) );
  XOR U100768 ( .A(n80722), .B(n80561), .Z(n86296) );
  IV U100769 ( .A(n80562), .Z(n80563) );
  NOR U100770 ( .A(n80564), .B(n80563), .Z(n80565) );
  IV U100771 ( .A(n80565), .Z(n86295) );
  XOR U100772 ( .A(n86296), .B(n86295), .Z(n80571) );
  IV U100773 ( .A(n80571), .Z(n80566) );
  NOR U100774 ( .A(n80567), .B(n80566), .Z(n86432) );
  NOR U100775 ( .A(n80569), .B(n80568), .Z(n80572) );
  IV U100776 ( .A(n80572), .Z(n80570) );
  NOR U100777 ( .A(n86296), .B(n80570), .Z(n86428) );
  NOR U100778 ( .A(n80572), .B(n80571), .Z(n80573) );
  NOR U100779 ( .A(n86428), .B(n80573), .Z(n80711) );
  NOR U100780 ( .A(n80574), .B(n80711), .Z(n80575) );
  NOR U100781 ( .A(n86432), .B(n80575), .Z(n80576) );
  IV U100782 ( .A(n80576), .Z(n80719) );
  XOR U100783 ( .A(n80718), .B(n80719), .Z(n80706) );
  XOR U100784 ( .A(n80577), .B(n80706), .Z(n80698) );
  IV U100785 ( .A(n80698), .Z(n80578) );
  NOR U100786 ( .A(n80579), .B(n80578), .Z(n80590) );
  IV U100787 ( .A(n80580), .Z(n80583) );
  NOR U100788 ( .A(n80585), .B(n80706), .Z(n80581) );
  IV U100789 ( .A(n80581), .Z(n80582) );
  NOR U100790 ( .A(n80583), .B(n80582), .Z(n86420) );
  IV U100791 ( .A(n80584), .Z(n80588) );
  NOR U100792 ( .A(n80585), .B(n80698), .Z(n80586) );
  IV U100793 ( .A(n80586), .Z(n80587) );
  NOR U100794 ( .A(n80588), .B(n80587), .Z(n92064) );
  NOR U100795 ( .A(n86420), .B(n92064), .Z(n80589) );
  IV U100796 ( .A(n80589), .Z(n86305) );
  NOR U100797 ( .A(n80590), .B(n86305), .Z(n86313) );
  IV U100798 ( .A(n80591), .Z(n80699) );
  NOR U100799 ( .A(n80592), .B(n80699), .Z(n80596) );
  IV U100800 ( .A(n80593), .Z(n80595) );
  NOR U100801 ( .A(n80595), .B(n80594), .Z(n86314) );
  NOR U100802 ( .A(n80596), .B(n86314), .Z(n80597) );
  XOR U100803 ( .A(n86313), .B(n80597), .Z(n80696) );
  XOR U100804 ( .A(n80694), .B(n80696), .Z(n86334) );
  IV U100805 ( .A(n86334), .Z(n80609) );
  IV U100806 ( .A(n80598), .Z(n80602) );
  IV U100807 ( .A(n80599), .Z(n80606) );
  NOR U100808 ( .A(n80606), .B(n80600), .Z(n80601) );
  IV U100809 ( .A(n80601), .Z(n86333) );
  NOR U100810 ( .A(n80602), .B(n86333), .Z(n80613) );
  IV U100811 ( .A(n80613), .Z(n80603) );
  NOR U100812 ( .A(n80609), .B(n80603), .Z(n80615) );
  IV U100813 ( .A(n80604), .Z(n80605) );
  NOR U100814 ( .A(n80606), .B(n80605), .Z(n80608) );
  IV U100815 ( .A(n80608), .Z(n80607) );
  NOR U100816 ( .A(n80696), .B(n80607), .Z(n86322) );
  NOR U100817 ( .A(n80609), .B(n80608), .Z(n80610) );
  NOR U100818 ( .A(n86322), .B(n80610), .Z(n80611) );
  IV U100819 ( .A(n80611), .Z(n80612) );
  NOR U100820 ( .A(n80613), .B(n80612), .Z(n80614) );
  NOR U100821 ( .A(n80615), .B(n80614), .Z(n80692) );
  IV U100822 ( .A(n80616), .Z(n80617) );
  NOR U100823 ( .A(n80617), .B(n86333), .Z(n80626) );
  IV U100824 ( .A(n80618), .Z(n80620) );
  NOR U100825 ( .A(n80620), .B(n80619), .Z(n80689) );
  IV U100826 ( .A(n80621), .Z(n80623) );
  NOR U100827 ( .A(n80623), .B(n80622), .Z(n80691) );
  NOR U100828 ( .A(n80689), .B(n80691), .Z(n80624) );
  IV U100829 ( .A(n80624), .Z(n80625) );
  NOR U100830 ( .A(n80626), .B(n80625), .Z(n80627) );
  XOR U100831 ( .A(n80692), .B(n80627), .Z(n80683) );
  IV U100832 ( .A(n80628), .Z(n80630) );
  NOR U100833 ( .A(n80630), .B(n80629), .Z(n80684) );
  NOR U100834 ( .A(n80686), .B(n80684), .Z(n80631) );
  XOR U100835 ( .A(n80683), .B(n80631), .Z(n86341) );
  XOR U100836 ( .A(n86342), .B(n86341), .Z(n80680) );
  IV U100837 ( .A(n80632), .Z(n80634) );
  NOR U100838 ( .A(n80634), .B(n80633), .Z(n86348) );
  IV U100839 ( .A(n80635), .Z(n80636) );
  NOR U100840 ( .A(n80637), .B(n80636), .Z(n80681) );
  NOR U100841 ( .A(n86348), .B(n80681), .Z(n80638) );
  XOR U100842 ( .A(n80680), .B(n80638), .Z(n80674) );
  XOR U100843 ( .A(n80675), .B(n80674), .Z(n86355) );
  IV U100844 ( .A(n86355), .Z(n80676) );
  NOR U100845 ( .A(n80667), .B(n80676), .Z(n80673) );
  NOR U100846 ( .A(n80640), .B(n80639), .Z(n80641) );
  XOR U100847 ( .A(n80642), .B(n80641), .Z(n86357) );
  XOR U100848 ( .A(n80644), .B(n80643), .Z(n86362) );
  NOR U100849 ( .A(n80646), .B(n80645), .Z(n80648) );
  XOR U100850 ( .A(n80648), .B(n80647), .Z(n92112) );
  NOR U100851 ( .A(n80650), .B(n80649), .Z(n86387) );
  NOR U100852 ( .A(n80651), .B(n86387), .Z(n80653) );
  XOR U100853 ( .A(n80653), .B(n80652), .Z(n92113) );
  NOR U100854 ( .A(n92112), .B(n92113), .Z(n80654) );
  IV U100855 ( .A(n80654), .Z(n86370) );
  XOR U100856 ( .A(n86386), .B(n86387), .Z(n92121) );
  IV U100857 ( .A(n92121), .Z(n86368) );
  IV U100858 ( .A(n80655), .Z(n80657) );
  NOR U100859 ( .A(n80657), .B(n80656), .Z(n92119) );
  IV U100860 ( .A(n92119), .Z(n86391) );
  NOR U100861 ( .A(n86368), .B(n86391), .Z(n86388) );
  IV U100862 ( .A(n86388), .Z(n92111) );
  NOR U100863 ( .A(n86370), .B(n92111), .Z(n86363) );
  IV U100864 ( .A(n86363), .Z(n80658) );
  NOR U100865 ( .A(n86362), .B(n80658), .Z(n86358) );
  IV U100866 ( .A(n86358), .Z(n80659) );
  NOR U100867 ( .A(n86361), .B(n80659), .Z(n86356) );
  IV U100868 ( .A(n86356), .Z(n80660) );
  NOR U100869 ( .A(n86357), .B(n80660), .Z(n86405) );
  IV U100870 ( .A(n86405), .Z(n80663) );
  XOR U100871 ( .A(n80662), .B(n80661), .Z(n86404) );
  NOR U100872 ( .A(n80663), .B(n86404), .Z(n86379) );
  IV U100873 ( .A(n86379), .Z(n80671) );
  IV U100874 ( .A(n80664), .Z(n80665) );
  NOR U100875 ( .A(n80666), .B(n80665), .Z(n86353) );
  XOR U100876 ( .A(n86353), .B(n86355), .Z(n80669) );
  NOR U100877 ( .A(n86355), .B(n80667), .Z(n80668) );
  NOR U100878 ( .A(n80669), .B(n80668), .Z(n80670) );
  NOR U100879 ( .A(n80671), .B(n80670), .Z(n80672) );
  NOR U100880 ( .A(n80673), .B(n80672), .Z(n92307) );
  NOR U100881 ( .A(n80675), .B(n80674), .Z(n80679) );
  IV U100882 ( .A(n86353), .Z(n80677) );
  NOR U100883 ( .A(n80677), .B(n80676), .Z(n80678) );
  NOR U100884 ( .A(n80679), .B(n80678), .Z(n92312) );
  IV U100885 ( .A(n92312), .Z(n86351) );
  IV U100886 ( .A(n80680), .Z(n86349) );
  IV U100887 ( .A(n80681), .Z(n80682) );
  NOR U100888 ( .A(n86349), .B(n80682), .Z(n86345) );
  IV U100889 ( .A(n86345), .Z(n86340) );
  IV U100890 ( .A(n80683), .Z(n80688) );
  IV U100891 ( .A(n80684), .Z(n80685) );
  NOR U100892 ( .A(n80688), .B(n80685), .Z(n92090) );
  IV U100893 ( .A(n80686), .Z(n80687) );
  NOR U100894 ( .A(n80688), .B(n80687), .Z(n92087) );
  IV U100895 ( .A(n80689), .Z(n80690) );
  NOR U100896 ( .A(n80690), .B(n80692), .Z(n92080) );
  IV U100897 ( .A(n80691), .Z(n80693) );
  NOR U100898 ( .A(n80693), .B(n80692), .Z(n92077) );
  IV U100899 ( .A(n80694), .Z(n80695) );
  NOR U100900 ( .A(n80696), .B(n80695), .Z(n86326) );
  IV U100901 ( .A(n80697), .Z(n80701) );
  NOR U100902 ( .A(n80699), .B(n80698), .Z(n80700) );
  IV U100903 ( .A(n80700), .Z(n86308) );
  NOR U100904 ( .A(n80701), .B(n86308), .Z(n86312) );
  IV U100905 ( .A(n86312), .Z(n92050) );
  IV U100906 ( .A(n80702), .Z(n80709) );
  NOR U100907 ( .A(n80704), .B(n80703), .Z(n80705) );
  IV U100908 ( .A(n80705), .Z(n80712) );
  NOR U100909 ( .A(n80706), .B(n80712), .Z(n80707) );
  IV U100910 ( .A(n80707), .Z(n80708) );
  NOR U100911 ( .A(n80709), .B(n80708), .Z(n92059) );
  IV U100912 ( .A(n92059), .Z(n92061) );
  IV U100913 ( .A(n80710), .Z(n80716) );
  IV U100914 ( .A(n80711), .Z(n80713) );
  NOR U100915 ( .A(n80713), .B(n80712), .Z(n80714) );
  IV U100916 ( .A(n80714), .Z(n80715) );
  NOR U100917 ( .A(n80716), .B(n80715), .Z(n80717) );
  IV U100918 ( .A(n80717), .Z(n86418) );
  IV U100919 ( .A(n80718), .Z(n80720) );
  NOR U100920 ( .A(n80720), .B(n80719), .Z(n86414) );
  NOR U100921 ( .A(n86432), .B(n86414), .Z(n86304) );
  IV U100922 ( .A(n80721), .Z(n80723) );
  IV U100923 ( .A(n80722), .Z(n86291) );
  NOR U100924 ( .A(n80723), .B(n86291), .Z(n86298) );
  IV U100925 ( .A(n80724), .Z(n80725) );
  NOR U100926 ( .A(n80728), .B(n80725), .Z(n92009) );
  IV U100927 ( .A(n80726), .Z(n80727) );
  NOR U100928 ( .A(n80728), .B(n80727), .Z(n92019) );
  IV U100929 ( .A(n80729), .Z(n80732) );
  IV U100930 ( .A(n80730), .Z(n80731) );
  NOR U100931 ( .A(n80732), .B(n80731), .Z(n92016) );
  IV U100932 ( .A(n80733), .Z(n80738) );
  IV U100933 ( .A(n80734), .Z(n80735) );
  NOR U100934 ( .A(n80736), .B(n80735), .Z(n80737) );
  IV U100935 ( .A(n80737), .Z(n86288) );
  NOR U100936 ( .A(n80738), .B(n86288), .Z(n80739) );
  IV U100937 ( .A(n80739), .Z(n92028) );
  IV U100938 ( .A(n80740), .Z(n80741) );
  NOR U100939 ( .A(n80747), .B(n80741), .Z(n80743) );
  NOR U100940 ( .A(n80743), .B(n80742), .Z(n86466) );
  IV U100941 ( .A(n80744), .Z(n80745) );
  NOR U100942 ( .A(n80746), .B(n80745), .Z(n80750) );
  NOR U100943 ( .A(n80748), .B(n80747), .Z(n80749) );
  NOR U100944 ( .A(n80750), .B(n80749), .Z(n86464) );
  IV U100945 ( .A(n80751), .Z(n80758) );
  IV U100946 ( .A(n80752), .Z(n80762) );
  NOR U100947 ( .A(n80753), .B(n80762), .Z(n80754) );
  IV U100948 ( .A(n80754), .Z(n80755) );
  NOR U100949 ( .A(n80756), .B(n80755), .Z(n80757) );
  IV U100950 ( .A(n80757), .Z(n86473) );
  NOR U100951 ( .A(n80758), .B(n86473), .Z(n86286) );
  IV U100952 ( .A(n80759), .Z(n80760) );
  NOR U100953 ( .A(n80760), .B(n86473), .Z(n86280) );
  IV U100954 ( .A(n80761), .Z(n80763) );
  NOR U100955 ( .A(n80763), .B(n80762), .Z(n86480) );
  IV U100956 ( .A(n80764), .Z(n80765) );
  NOR U100957 ( .A(n80766), .B(n80765), .Z(n86469) );
  NOR U100958 ( .A(n86480), .B(n86469), .Z(n86278) );
  NOR U100959 ( .A(n80775), .B(n80771), .Z(n80767) );
  IV U100960 ( .A(n80767), .Z(n80768) );
  NOR U100961 ( .A(n80769), .B(n80768), .Z(n92002) );
  IV U100962 ( .A(n80770), .Z(n80772) );
  NOR U100963 ( .A(n80772), .B(n80771), .Z(n80773) );
  IV U100964 ( .A(n80773), .Z(n80774) );
  NOR U100965 ( .A(n80775), .B(n80774), .Z(n91999) );
  IV U100966 ( .A(n80776), .Z(n80777) );
  NOR U100967 ( .A(n86276), .B(n80777), .Z(n86455) );
  IV U100968 ( .A(n80778), .Z(n80780) );
  NOR U100969 ( .A(n80780), .B(n80779), .Z(n80785) );
  IV U100970 ( .A(n80781), .Z(n80783) );
  NOR U100971 ( .A(n80783), .B(n80782), .Z(n80784) );
  NOR U100972 ( .A(n80785), .B(n80784), .Z(n86438) );
  IV U100973 ( .A(n80786), .Z(n80787) );
  NOR U100974 ( .A(n80787), .B(n80789), .Z(n86440) );
  IV U100975 ( .A(n80788), .Z(n80790) );
  NOR U100976 ( .A(n80790), .B(n80789), .Z(n91963) );
  NOR U100977 ( .A(n86440), .B(n91963), .Z(n86259) );
  IV U100978 ( .A(n80791), .Z(n80792) );
  NOR U100979 ( .A(n80793), .B(n80792), .Z(n91981) );
  IV U100980 ( .A(n80797), .Z(n80794) );
  NOR U100981 ( .A(n80795), .B(n80794), .Z(n80802) );
  NOR U100982 ( .A(n80797), .B(n80796), .Z(n80800) );
  IV U100983 ( .A(n80798), .Z(n80799) );
  NOR U100984 ( .A(n80800), .B(n80799), .Z(n80801) );
  NOR U100985 ( .A(n80802), .B(n80801), .Z(n91972) );
  IV U100986 ( .A(n80803), .Z(n80805) );
  NOR U100987 ( .A(n80805), .B(n80804), .Z(n91978) );
  IV U100988 ( .A(n80806), .Z(n86236) );
  IV U100989 ( .A(n80807), .Z(n80808) );
  NOR U100990 ( .A(n86236), .B(n80808), .Z(n86247) );
  IV U100991 ( .A(n80809), .Z(n80810) );
  NOR U100992 ( .A(n86236), .B(n80810), .Z(n86243) );
  IV U100993 ( .A(n80811), .Z(n80813) );
  NOR U100994 ( .A(n80813), .B(n80812), .Z(n91936) );
  IV U100995 ( .A(n80814), .Z(n80815) );
  NOR U100996 ( .A(n86232), .B(n80815), .Z(n91952) );
  IV U100997 ( .A(n80816), .Z(n80818) );
  NOR U100998 ( .A(n80818), .B(n80817), .Z(n86491) );
  IV U100999 ( .A(n80819), .Z(n80822) );
  NOR U101000 ( .A(n80822), .B(n80820), .Z(n86493) );
  IV U101001 ( .A(n80821), .Z(n80823) );
  NOR U101002 ( .A(n80823), .B(n80822), .Z(n80827) );
  IV U101003 ( .A(n80824), .Z(n80825) );
  NOR U101004 ( .A(n80825), .B(n80829), .Z(n80826) );
  NOR U101005 ( .A(n80827), .B(n80826), .Z(n86519) );
  IV U101006 ( .A(n80828), .Z(n80830) );
  NOR U101007 ( .A(n80830), .B(n80829), .Z(n86544) );
  IV U101008 ( .A(n80831), .Z(n80834) );
  IV U101009 ( .A(n80832), .Z(n80833) );
  NOR U101010 ( .A(n80834), .B(n80833), .Z(n86541) );
  IV U101011 ( .A(n80835), .Z(n80836) );
  NOR U101012 ( .A(n80836), .B(n86202), .Z(n86525) );
  IV U101013 ( .A(n80837), .Z(n80838) );
  NOR U101014 ( .A(n86202), .B(n80838), .Z(n86531) );
  IV U101015 ( .A(n80839), .Z(n80840) );
  NOR U101016 ( .A(n86208), .B(n80840), .Z(n86528) );
  IV U101017 ( .A(n80841), .Z(n80843) );
  IV U101018 ( .A(n80842), .Z(n80845) );
  NOR U101019 ( .A(n80843), .B(n80845), .Z(n86514) );
  IV U101020 ( .A(n80844), .Z(n80846) );
  NOR U101021 ( .A(n80846), .B(n80845), .Z(n86503) );
  IV U101022 ( .A(n80847), .Z(n80848) );
  NOR U101023 ( .A(n80853), .B(n80848), .Z(n86501) );
  IV U101024 ( .A(n80849), .Z(n80850) );
  NOR U101025 ( .A(n80853), .B(n80850), .Z(n86505) );
  IV U101026 ( .A(n80851), .Z(n80852) );
  NOR U101027 ( .A(n80853), .B(n80852), .Z(n86510) );
  IV U101028 ( .A(n80855), .Z(n80854) );
  NOR U101029 ( .A(n80854), .B(n86190), .Z(n80860) );
  XOR U101030 ( .A(n80855), .B(n86190), .Z(n80858) );
  IV U101031 ( .A(n80856), .Z(n80857) );
  NOR U101032 ( .A(n80858), .B(n80857), .Z(n80859) );
  NOR U101033 ( .A(n80860), .B(n80859), .Z(n86576) );
  IV U101034 ( .A(n80861), .Z(n80863) );
  NOR U101035 ( .A(n80863), .B(n80862), .Z(n86181) );
  IV U101036 ( .A(n80864), .Z(n80865) );
  NOR U101037 ( .A(n80866), .B(n80865), .Z(n86558) );
  IV U101038 ( .A(n80867), .Z(n80869) );
  NOR U101039 ( .A(n80869), .B(n80868), .Z(n86564) );
  NOR U101040 ( .A(n86558), .B(n86564), .Z(n86168) );
  IV U101041 ( .A(n80870), .Z(n80879) );
  IV U101042 ( .A(n80871), .Z(n80872) );
  NOR U101043 ( .A(n80879), .B(n80872), .Z(n80876) );
  IV U101044 ( .A(n80873), .Z(n80874) );
  NOR U101045 ( .A(n80874), .B(n86158), .Z(n80875) );
  NOR U101046 ( .A(n80876), .B(n80875), .Z(n86570) );
  IV U101047 ( .A(n80877), .Z(n80878) );
  NOR U101048 ( .A(n80879), .B(n80878), .Z(n86591) );
  IV U101049 ( .A(n80880), .Z(n80881) );
  NOR U101050 ( .A(n80882), .B(n80881), .Z(n86588) );
  IV U101051 ( .A(n80883), .Z(n80887) );
  IV U101052 ( .A(n80884), .Z(n80888) );
  NOR U101053 ( .A(n80885), .B(n80888), .Z(n80886) );
  IV U101054 ( .A(n80886), .Z(n80891) );
  NOR U101055 ( .A(n80887), .B(n80891), .Z(n91909) );
  NOR U101056 ( .A(n80889), .B(n80888), .Z(n80894) );
  IV U101057 ( .A(n80890), .Z(n80892) );
  NOR U101058 ( .A(n80892), .B(n80891), .Z(n80893) );
  NOR U101059 ( .A(n80894), .B(n80893), .Z(n91908) );
  NOR U101060 ( .A(n80896), .B(n80895), .Z(n91917) );
  IV U101061 ( .A(n80897), .Z(n80898) );
  NOR U101062 ( .A(n86133), .B(n80898), .Z(n80899) );
  IV U101063 ( .A(n80899), .Z(n86615) );
  IV U101064 ( .A(n80900), .Z(n80902) );
  NOR U101065 ( .A(n80902), .B(n80901), .Z(n86127) );
  IV U101066 ( .A(n86127), .Z(n86125) );
  IV U101067 ( .A(n80903), .Z(n80904) );
  NOR U101068 ( .A(n80904), .B(n80906), .Z(n91881) );
  IV U101069 ( .A(n80905), .Z(n80907) );
  NOR U101070 ( .A(n80907), .B(n80906), .Z(n91884) );
  IV U101071 ( .A(n80908), .Z(n86104) );
  IV U101072 ( .A(n80909), .Z(n80910) );
  NOR U101073 ( .A(n86104), .B(n80910), .Z(n86632) );
  IV U101074 ( .A(n80911), .Z(n80913) );
  NOR U101075 ( .A(n80913), .B(n80912), .Z(n86629) );
  IV U101076 ( .A(n80916), .Z(n80914) );
  NOR U101077 ( .A(n80915), .B(n80914), .Z(n80922) );
  NOR U101078 ( .A(n80917), .B(n80916), .Z(n80920) );
  IV U101079 ( .A(n80918), .Z(n80919) );
  NOR U101080 ( .A(n80920), .B(n80919), .Z(n80921) );
  NOR U101081 ( .A(n80922), .B(n80921), .Z(n86642) );
  IV U101082 ( .A(n80923), .Z(n86095) );
  IV U101083 ( .A(n80924), .Z(n80925) );
  NOR U101084 ( .A(n86095), .B(n80925), .Z(n80926) );
  IV U101085 ( .A(n80926), .Z(n91860) );
  IV U101086 ( .A(n80927), .Z(n80929) );
  NOR U101087 ( .A(n80929), .B(n80928), .Z(n86083) );
  IV U101088 ( .A(n80930), .Z(n80932) );
  NOR U101089 ( .A(n80932), .B(n80931), .Z(n86065) );
  IV U101090 ( .A(n80933), .Z(n80939) );
  IV U101091 ( .A(n80934), .Z(n80935) );
  NOR U101092 ( .A(n80939), .B(n80935), .Z(n80936) );
  IV U101093 ( .A(n80936), .Z(n86647) );
  IV U101094 ( .A(n80937), .Z(n80938) );
  NOR U101095 ( .A(n80939), .B(n80938), .Z(n86643) );
  IV U101096 ( .A(n80940), .Z(n80941) );
  NOR U101097 ( .A(n80941), .B(n80943), .Z(n91832) );
  IV U101098 ( .A(n80942), .Z(n80944) );
  NOR U101099 ( .A(n80944), .B(n80943), .Z(n91838) );
  XOR U101100 ( .A(n91832), .B(n91838), .Z(n80945) );
  NOR U101101 ( .A(n86643), .B(n80945), .Z(n86056) );
  IV U101102 ( .A(n80946), .Z(n80947) );
  NOR U101103 ( .A(n80948), .B(n80947), .Z(n91835) );
  IV U101104 ( .A(n80949), .Z(n80951) );
  NOR U101105 ( .A(n80951), .B(n80950), .Z(n80955) );
  NOR U101106 ( .A(n80953), .B(n80952), .Z(n80954) );
  NOR U101107 ( .A(n80955), .B(n80954), .Z(n86659) );
  IV U101108 ( .A(n80956), .Z(n80957) );
  NOR U101109 ( .A(n86049), .B(n80957), .Z(n86663) );
  IV U101110 ( .A(n80958), .Z(n80959) );
  NOR U101111 ( .A(n80959), .B(n86020), .Z(n91815) );
  IV U101112 ( .A(n80960), .Z(n80962) );
  NOR U101113 ( .A(n80962), .B(n80961), .Z(n91812) );
  IV U101114 ( .A(n80963), .Z(n80965) );
  NOR U101115 ( .A(n80965), .B(n80964), .Z(n86024) );
  IV U101116 ( .A(n80966), .Z(n80967) );
  NOR U101117 ( .A(n80968), .B(n80967), .Z(n91771) );
  IV U101118 ( .A(n80969), .Z(n80970) );
  NOR U101119 ( .A(n80971), .B(n80970), .Z(n86708) );
  IV U101120 ( .A(n80972), .Z(n80973) );
  NOR U101121 ( .A(n86005), .B(n80973), .Z(n91780) );
  NOR U101122 ( .A(n86708), .B(n91780), .Z(n86003) );
  IV U101123 ( .A(n80974), .Z(n80975) );
  NOR U101124 ( .A(n80976), .B(n80975), .Z(n91784) );
  IV U101125 ( .A(n80977), .Z(n80978) );
  NOR U101126 ( .A(n80979), .B(n80978), .Z(n91787) );
  IV U101127 ( .A(n80980), .Z(n80981) );
  NOR U101128 ( .A(n80982), .B(n80981), .Z(n91797) );
  IV U101129 ( .A(n80983), .Z(n86001) );
  NOR U101130 ( .A(n80984), .B(n86001), .Z(n80985) );
  NOR U101131 ( .A(n80986), .B(n80985), .Z(n91796) );
  IV U101132 ( .A(n80987), .Z(n80988) );
  NOR U101133 ( .A(n80988), .B(n80993), .Z(n86713) );
  IV U101134 ( .A(n80989), .Z(n80990) );
  NOR U101135 ( .A(n80991), .B(n80990), .Z(n80996) );
  IV U101136 ( .A(n80992), .Z(n80994) );
  NOR U101137 ( .A(n80994), .B(n80993), .Z(n80995) );
  NOR U101138 ( .A(n80996), .B(n80995), .Z(n86712) );
  XOR U101139 ( .A(n81007), .B(n81009), .Z(n80999) );
  IV U101140 ( .A(n80997), .Z(n80998) );
  NOR U101141 ( .A(n80999), .B(n80998), .Z(n81000) );
  IV U101142 ( .A(n81000), .Z(n86669) );
  IV U101143 ( .A(n81001), .Z(n81002) );
  NOR U101144 ( .A(n81009), .B(n81002), .Z(n86678) );
  IV U101145 ( .A(n81003), .Z(n81006) );
  IV U101146 ( .A(n81004), .Z(n81005) );
  NOR U101147 ( .A(n81006), .B(n81005), .Z(n86671) );
  NOR U101148 ( .A(n86678), .B(n86671), .Z(n85996) );
  IV U101149 ( .A(n81007), .Z(n81008) );
  NOR U101150 ( .A(n81009), .B(n81008), .Z(n86680) );
  IV U101151 ( .A(n86680), .Z(n86677) );
  IV U101152 ( .A(n81010), .Z(n81013) );
  IV U101153 ( .A(n81011), .Z(n81012) );
  NOR U101154 ( .A(n81013), .B(n81012), .Z(n86687) );
  IV U101155 ( .A(n81014), .Z(n81015) );
  NOR U101156 ( .A(n81016), .B(n81015), .Z(n85989) );
  IV U101157 ( .A(n85989), .Z(n86694) );
  IV U101158 ( .A(n81017), .Z(n81019) );
  NOR U101159 ( .A(n81019), .B(n81018), .Z(n81020) );
  NOR U101160 ( .A(n81021), .B(n81020), .Z(n91756) );
  NOR U101161 ( .A(n81023), .B(n81022), .Z(n81024) );
  IV U101162 ( .A(n81024), .Z(n91735) );
  IV U101163 ( .A(n81025), .Z(n81027) );
  NOR U101164 ( .A(n81027), .B(n81026), .Z(n91747) );
  IV U101165 ( .A(n81028), .Z(n81030) );
  NOR U101166 ( .A(n81030), .B(n81029), .Z(n91737) );
  NOR U101167 ( .A(n91747), .B(n91737), .Z(n85987) );
  IV U101168 ( .A(n81031), .Z(n81032) );
  NOR U101169 ( .A(n81035), .B(n81032), .Z(n91742) );
  IV U101170 ( .A(n91742), .Z(n91745) );
  IV U101171 ( .A(n81033), .Z(n81034) );
  NOR U101172 ( .A(n81035), .B(n81034), .Z(n81036) );
  IV U101173 ( .A(n81036), .Z(n86733) );
  NOR U101174 ( .A(n81042), .B(n81037), .Z(n86741) );
  IV U101175 ( .A(n81038), .Z(n81039) );
  NOR U101176 ( .A(n81039), .B(n81042), .Z(n81040) );
  IV U101177 ( .A(n81040), .Z(n86739) );
  IV U101178 ( .A(n81041), .Z(n81043) );
  NOR U101179 ( .A(n81043), .B(n81042), .Z(n81047) );
  IV U101180 ( .A(n81044), .Z(n81045) );
  NOR U101181 ( .A(n81045), .B(n85964), .Z(n81046) );
  NOR U101182 ( .A(n81047), .B(n81046), .Z(n86726) );
  IV U101183 ( .A(n81048), .Z(n81049) );
  NOR U101184 ( .A(n81050), .B(n81049), .Z(n86822) );
  IV U101185 ( .A(n81053), .Z(n81051) );
  NOR U101186 ( .A(n81052), .B(n81051), .Z(n81059) );
  NOR U101187 ( .A(n81054), .B(n81053), .Z(n81057) );
  IV U101188 ( .A(n81055), .Z(n81056) );
  NOR U101189 ( .A(n81057), .B(n81056), .Z(n81058) );
  NOR U101190 ( .A(n81059), .B(n81058), .Z(n86760) );
  IV U101191 ( .A(n81060), .Z(n81061) );
  NOR U101192 ( .A(n81061), .B(n85955), .Z(n85961) );
  IV U101193 ( .A(n85961), .Z(n85959) );
  NOR U101194 ( .A(n81063), .B(n81062), .Z(n81064) );
  IV U101195 ( .A(n81064), .Z(n81065) );
  NOR U101196 ( .A(n85944), .B(n81065), .Z(n85949) );
  IV U101197 ( .A(n85949), .Z(n85943) );
  IV U101198 ( .A(n81066), .Z(n81067) );
  NOR U101199 ( .A(n81067), .B(n85945), .Z(n81068) );
  IV U101200 ( .A(n81068), .Z(n86801) );
  IV U101201 ( .A(n81069), .Z(n81070) );
  NOR U101202 ( .A(n81071), .B(n81070), .Z(n81076) );
  IV U101203 ( .A(n81072), .Z(n81074) );
  NOR U101204 ( .A(n81074), .B(n81073), .Z(n81075) );
  NOR U101205 ( .A(n81076), .B(n81075), .Z(n86806) );
  IV U101206 ( .A(n81077), .Z(n81079) );
  NOR U101207 ( .A(n81079), .B(n81078), .Z(n86802) );
  IV U101208 ( .A(n81080), .Z(n81081) );
  NOR U101209 ( .A(n81081), .B(n81085), .Z(n81082) );
  IV U101210 ( .A(n81082), .Z(n86766) );
  IV U101211 ( .A(n81083), .Z(n81084) );
  NOR U101212 ( .A(n81085), .B(n81084), .Z(n86787) );
  IV U101213 ( .A(n81086), .Z(n81088) );
  NOR U101214 ( .A(n81088), .B(n81087), .Z(n86768) );
  NOR U101215 ( .A(n86787), .B(n86768), .Z(n85942) );
  IV U101216 ( .A(n81089), .Z(n81094) );
  IV U101217 ( .A(n81090), .Z(n81091) );
  NOR U101218 ( .A(n81094), .B(n81091), .Z(n86782) );
  IV U101219 ( .A(n86782), .Z(n86784) );
  IV U101220 ( .A(n81092), .Z(n81096) );
  NOR U101221 ( .A(n81094), .B(n81093), .Z(n81095) );
  IV U101222 ( .A(n81095), .Z(n85938) );
  NOR U101223 ( .A(n81096), .B(n85938), .Z(n81097) );
  IV U101224 ( .A(n81097), .Z(n86773) );
  IV U101225 ( .A(n81098), .Z(n81099) );
  NOR U101226 ( .A(n81100), .B(n81099), .Z(n81106) );
  IV U101227 ( .A(n81101), .Z(n81104) );
  IV U101228 ( .A(n81102), .Z(n81103) );
  NOR U101229 ( .A(n81104), .B(n81103), .Z(n81105) );
  NOR U101230 ( .A(n81106), .B(n81105), .Z(n86851) );
  IV U101231 ( .A(n81107), .Z(n81109) );
  NOR U101232 ( .A(n81109), .B(n81108), .Z(n86847) );
  IV U101233 ( .A(n81110), .Z(n81112) );
  NOR U101234 ( .A(n81112), .B(n81111), .Z(n81113) );
  IV U101235 ( .A(n81113), .Z(n86838) );
  IV U101236 ( .A(n81114), .Z(n81115) );
  NOR U101237 ( .A(n81116), .B(n81115), .Z(n86897) );
  IV U101238 ( .A(n81117), .Z(n81118) );
  NOR U101239 ( .A(n81118), .B(n85918), .Z(n86840) );
  NOR U101240 ( .A(n86897), .B(n86840), .Z(n85914) );
  IV U101241 ( .A(n81119), .Z(n81120) );
  NOR U101242 ( .A(n81123), .B(n81120), .Z(n86892) );
  IV U101243 ( .A(n86892), .Z(n86894) );
  IV U101244 ( .A(n81121), .Z(n81122) );
  NOR U101245 ( .A(n81123), .B(n81122), .Z(n81124) );
  IV U101246 ( .A(n81124), .Z(n86880) );
  IV U101247 ( .A(n81125), .Z(n81127) );
  IV U101248 ( .A(n81126), .Z(n81132) );
  NOR U101249 ( .A(n81127), .B(n81132), .Z(n86876) );
  IV U101250 ( .A(n81128), .Z(n81129) );
  NOR U101251 ( .A(n81130), .B(n81129), .Z(n86887) );
  IV U101252 ( .A(n81131), .Z(n81133) );
  NOR U101253 ( .A(n81133), .B(n81132), .Z(n86872) );
  NOR U101254 ( .A(n86887), .B(n86872), .Z(n85913) );
  IV U101255 ( .A(n81134), .Z(n81135) );
  NOR U101256 ( .A(n81136), .B(n81135), .Z(n86889) );
  NOR U101257 ( .A(n81138), .B(n81137), .Z(n86890) );
  NOR U101258 ( .A(n86889), .B(n86890), .Z(n85908) );
  IV U101259 ( .A(n81139), .Z(n81141) );
  NOR U101260 ( .A(n81141), .B(n81140), .Z(n86905) );
  NOR U101261 ( .A(n81143), .B(n81142), .Z(n81149) );
  IV U101262 ( .A(n81143), .Z(n81145) );
  NOR U101263 ( .A(n81145), .B(n81144), .Z(n81146) );
  NOR U101264 ( .A(n81147), .B(n81146), .Z(n81148) );
  NOR U101265 ( .A(n81149), .B(n81148), .Z(n86902) );
  IV U101266 ( .A(n81150), .Z(n81151) );
  NOR U101267 ( .A(n81151), .B(n85905), .Z(n86913) );
  IV U101268 ( .A(n91707), .Z(n91711) );
  IV U101269 ( .A(n81152), .Z(n81154) );
  NOR U101270 ( .A(n81154), .B(n81153), .Z(n86936) );
  NOR U101271 ( .A(n81156), .B(n81155), .Z(n81157) );
  NOR U101272 ( .A(n81157), .B(n81158), .Z(n86920) );
  IV U101273 ( .A(n81158), .Z(n81162) );
  NOR U101274 ( .A(n81162), .B(n81159), .Z(n86921) );
  IV U101275 ( .A(n81160), .Z(n81161) );
  NOR U101276 ( .A(n81162), .B(n81161), .Z(n86923) );
  NOR U101277 ( .A(n86921), .B(n86923), .Z(n85882) );
  IV U101278 ( .A(n81163), .Z(n81164) );
  NOR U101279 ( .A(n81167), .B(n81164), .Z(n85877) );
  IV U101280 ( .A(n81165), .Z(n81166) );
  NOR U101281 ( .A(n81167), .B(n81166), .Z(n85880) );
  IV U101282 ( .A(n85880), .Z(n85871) );
  XOR U101283 ( .A(n85877), .B(n85871), .Z(n85870) );
  NOR U101284 ( .A(n81168), .B(n81169), .Z(n81175) );
  IV U101285 ( .A(n81169), .Z(n81170) );
  NOR U101286 ( .A(n81171), .B(n81170), .Z(n81172) );
  NOR U101287 ( .A(n81173), .B(n81172), .Z(n81174) );
  NOR U101288 ( .A(n81175), .B(n81174), .Z(n81176) );
  IV U101289 ( .A(n81176), .Z(n86971) );
  IV U101290 ( .A(n81177), .Z(n81179) );
  NOR U101291 ( .A(n81179), .B(n81178), .Z(n85852) );
  IV U101292 ( .A(n81180), .Z(n85843) );
  NOR U101293 ( .A(n85843), .B(n85842), .Z(n91685) );
  IV U101294 ( .A(n81181), .Z(n81182) );
  NOR U101295 ( .A(n81182), .B(n85842), .Z(n86950) );
  NOR U101296 ( .A(n81184), .B(n81183), .Z(n86945) );
  IV U101297 ( .A(n81185), .Z(n85830) );
  IV U101298 ( .A(n81186), .Z(n81187) );
  NOR U101299 ( .A(n85830), .B(n81187), .Z(n86955) );
  NOR U101300 ( .A(n86945), .B(n86955), .Z(n85828) );
  IV U101301 ( .A(n81188), .Z(n81189) );
  NOR U101302 ( .A(n81189), .B(n85817), .Z(n91657) );
  NOR U101303 ( .A(n81191), .B(n81190), .Z(n91672) );
  IV U101304 ( .A(n81192), .Z(n81194) );
  NOR U101305 ( .A(n81194), .B(n81193), .Z(n91655) );
  NOR U101306 ( .A(n91672), .B(n91655), .Z(n85813) );
  IV U101307 ( .A(n81195), .Z(n81196) );
  NOR U101308 ( .A(n81197), .B(n81196), .Z(n81202) );
  IV U101309 ( .A(n81198), .Z(n81200) );
  NOR U101310 ( .A(n81200), .B(n81199), .Z(n81201) );
  NOR U101311 ( .A(n81202), .B(n81201), .Z(n91671) );
  IV U101312 ( .A(n81203), .Z(n81205) );
  NOR U101313 ( .A(n81205), .B(n81204), .Z(n86992) );
  IV U101314 ( .A(n81206), .Z(n81207) );
  NOR U101315 ( .A(n81208), .B(n81207), .Z(n81213) );
  IV U101316 ( .A(n81209), .Z(n81210) );
  NOR U101317 ( .A(n81211), .B(n81210), .Z(n81212) );
  NOR U101318 ( .A(n81213), .B(n81212), .Z(n81214) );
  IV U101319 ( .A(n81214), .Z(n86983) );
  IV U101320 ( .A(n81215), .Z(n81217) );
  NOR U101321 ( .A(n81217), .B(n81216), .Z(n86984) );
  NOR U101322 ( .A(n86983), .B(n86984), .Z(n81218) );
  IV U101323 ( .A(n81218), .Z(n85811) );
  IV U101324 ( .A(n81219), .Z(n81224) );
  IV U101325 ( .A(n81220), .Z(n81221) );
  NOR U101326 ( .A(n81224), .B(n81221), .Z(n86980) );
  IV U101327 ( .A(n81222), .Z(n81223) );
  NOR U101328 ( .A(n81224), .B(n81223), .Z(n81225) );
  IV U101329 ( .A(n81225), .Z(n87003) );
  IV U101330 ( .A(n81226), .Z(n81230) );
  IV U101331 ( .A(n81227), .Z(n81232) );
  NOR U101332 ( .A(n81232), .B(n81228), .Z(n81229) );
  IV U101333 ( .A(n81229), .Z(n85793) );
  NOR U101334 ( .A(n81230), .B(n85793), .Z(n91608) );
  NOR U101335 ( .A(n81232), .B(n81231), .Z(n81240) );
  IV U101336 ( .A(n81233), .Z(n81234) );
  NOR U101337 ( .A(n81235), .B(n81234), .Z(n81236) );
  IV U101338 ( .A(n81236), .Z(n81237) );
  NOR U101339 ( .A(n81238), .B(n81237), .Z(n81239) );
  NOR U101340 ( .A(n81240), .B(n81239), .Z(n91620) );
  IV U101341 ( .A(n81241), .Z(n81245) );
  NOR U101342 ( .A(n81242), .B(n81255), .Z(n81243) );
  IV U101343 ( .A(n81243), .Z(n81244) );
  NOR U101344 ( .A(n81245), .B(n81244), .Z(n91616) );
  NOR U101345 ( .A(n81246), .B(n81247), .Z(n81253) );
  IV U101346 ( .A(n81247), .Z(n81248) );
  NOR U101347 ( .A(n81249), .B(n81248), .Z(n81250) );
  NOR U101348 ( .A(n81251), .B(n81250), .Z(n81252) );
  NOR U101349 ( .A(n81253), .B(n81252), .Z(n91632) );
  NOR U101350 ( .A(n81255), .B(n81254), .Z(n91629) );
  IV U101351 ( .A(n81256), .Z(n81259) );
  IV U101352 ( .A(n81257), .Z(n81258) );
  NOR U101353 ( .A(n81259), .B(n81258), .Z(n87038) );
  IV U101354 ( .A(n81260), .Z(n81262) );
  NOR U101355 ( .A(n81262), .B(n81261), .Z(n81263) );
  IV U101356 ( .A(n81263), .Z(n87037) );
  NOR U101357 ( .A(n81265), .B(n81264), .Z(n87013) );
  IV U101358 ( .A(n87013), .Z(n87011) );
  IV U101359 ( .A(n81266), .Z(n81267) );
  NOR U101360 ( .A(n81267), .B(n85762), .Z(n85756) );
  IV U101361 ( .A(n85756), .Z(n85748) );
  IV U101362 ( .A(n85753), .Z(n91578) );
  IV U101363 ( .A(n81268), .Z(n81269) );
  NOR U101364 ( .A(n81269), .B(n81273), .Z(n91576) );
  IV U101365 ( .A(n81270), .Z(n81271) );
  NOR U101366 ( .A(n81271), .B(n81273), .Z(n91583) );
  IV U101367 ( .A(n81272), .Z(n81274) );
  NOR U101368 ( .A(n81274), .B(n81273), .Z(n91584) );
  XOR U101369 ( .A(n91583), .B(n91584), .Z(n81275) );
  NOR U101370 ( .A(n91576), .B(n81275), .Z(n85746) );
  IV U101371 ( .A(n81276), .Z(n85739) );
  IV U101372 ( .A(n81277), .Z(n81278) );
  NOR U101373 ( .A(n85739), .B(n81278), .Z(n87077) );
  IV U101374 ( .A(n81279), .Z(n81282) );
  NOR U101375 ( .A(n81282), .B(n81280), .Z(n81287) );
  IV U101376 ( .A(n81281), .Z(n81285) );
  NOR U101377 ( .A(n81283), .B(n81282), .Z(n81284) );
  IV U101378 ( .A(n81284), .Z(n85734) );
  NOR U101379 ( .A(n81285), .B(n85734), .Z(n81286) );
  NOR U101380 ( .A(n81287), .B(n81286), .Z(n91564) );
  IV U101381 ( .A(n81288), .Z(n81290) );
  NOR U101382 ( .A(n81290), .B(n81289), .Z(n87067) );
  IV U101383 ( .A(n81291), .Z(n81293) );
  NOR U101384 ( .A(n81293), .B(n81292), .Z(n87089) );
  IV U101385 ( .A(n81294), .Z(n81295) );
  NOR U101386 ( .A(n81296), .B(n81295), .Z(n87094) );
  IV U101387 ( .A(n81297), .Z(n81299) );
  NOR U101388 ( .A(n81299), .B(n81298), .Z(n81303) );
  IV U101389 ( .A(n81300), .Z(n81301) );
  NOR U101390 ( .A(n81309), .B(n81301), .Z(n81302) );
  NOR U101391 ( .A(n81303), .B(n81302), .Z(n87093) );
  IV U101392 ( .A(n87093), .Z(n85703) );
  IV U101393 ( .A(n81304), .Z(n81305) );
  NOR U101394 ( .A(n81306), .B(n81305), .Z(n87082) );
  IV U101395 ( .A(n81307), .Z(n81308) );
  NOR U101396 ( .A(n81309), .B(n81308), .Z(n87085) );
  IV U101397 ( .A(n81310), .Z(n81311) );
  NOR U101398 ( .A(n81312), .B(n81311), .Z(n81317) );
  IV U101399 ( .A(n81313), .Z(n81315) );
  NOR U101400 ( .A(n81315), .B(n81314), .Z(n81316) );
  NOR U101401 ( .A(n81317), .B(n81316), .Z(n87103) );
  IV U101402 ( .A(n81318), .Z(n81319) );
  NOR U101403 ( .A(n81319), .B(n85690), .Z(n87131) );
  IV U101404 ( .A(n81320), .Z(n81321) );
  NOR U101405 ( .A(n85675), .B(n81321), .Z(n87138) );
  IV U101406 ( .A(n81322), .Z(n81323) );
  NOR U101407 ( .A(n81324), .B(n81323), .Z(n81329) );
  IV U101408 ( .A(n81325), .Z(n81327) );
  NOR U101409 ( .A(n81327), .B(n81326), .Z(n81328) );
  NOR U101410 ( .A(n81329), .B(n81328), .Z(n87123) );
  IV U101411 ( .A(n81330), .Z(n81332) );
  NOR U101412 ( .A(n81332), .B(n81331), .Z(n87112) );
  IV U101413 ( .A(n81333), .Z(n81334) );
  NOR U101414 ( .A(n81335), .B(n81334), .Z(n87110) );
  NOR U101415 ( .A(n87112), .B(n87110), .Z(n85673) );
  IV U101416 ( .A(n81336), .Z(n81337) );
  NOR U101417 ( .A(n81338), .B(n81337), .Z(n91531) );
  IV U101418 ( .A(n81339), .Z(n81341) );
  NOR U101419 ( .A(n81341), .B(n81340), .Z(n87115) );
  NOR U101420 ( .A(n91531), .B(n87115), .Z(n85672) );
  IV U101421 ( .A(n81342), .Z(n81345) );
  IV U101422 ( .A(n81343), .Z(n81344) );
  NOR U101423 ( .A(n81345), .B(n81344), .Z(n91526) );
  IV U101424 ( .A(n91526), .Z(n91529) );
  IV U101425 ( .A(n81346), .Z(n81347) );
  NOR U101426 ( .A(n81348), .B(n81347), .Z(n81349) );
  IV U101427 ( .A(n81349), .Z(n91534) );
  IV U101428 ( .A(n81350), .Z(n81351) );
  NOR U101429 ( .A(n81352), .B(n81351), .Z(n91536) );
  IV U101430 ( .A(n81353), .Z(n81356) );
  NOR U101431 ( .A(n81354), .B(n81361), .Z(n81355) );
  IV U101432 ( .A(n81355), .Z(n81358) );
  NOR U101433 ( .A(n81356), .B(n81358), .Z(n91502) );
  IV U101434 ( .A(n81357), .Z(n81359) );
  NOR U101435 ( .A(n81359), .B(n81358), .Z(n91506) );
  IV U101436 ( .A(n81360), .Z(n81362) );
  NOR U101437 ( .A(n81362), .B(n81361), .Z(n91499) );
  IV U101438 ( .A(n81363), .Z(n81364) );
  NOR U101439 ( .A(n81369), .B(n81364), .Z(n91492) );
  IV U101440 ( .A(n81365), .Z(n81367) );
  NOR U101441 ( .A(n81367), .B(n81366), .Z(n87189) );
  IV U101442 ( .A(n81368), .Z(n81370) );
  NOR U101443 ( .A(n81370), .B(n81369), .Z(n91489) );
  NOR U101444 ( .A(n87189), .B(n91489), .Z(n85671) );
  IV U101445 ( .A(n81371), .Z(n81372) );
  NOR U101446 ( .A(n81373), .B(n81372), .Z(n91519) );
  IV U101447 ( .A(n81374), .Z(n81375) );
  NOR U101448 ( .A(n81376), .B(n81375), .Z(n87191) );
  NOR U101449 ( .A(n91519), .B(n87191), .Z(n85670) );
  IV U101450 ( .A(n81377), .Z(n81379) );
  IV U101451 ( .A(n81378), .Z(n85667) );
  NOR U101452 ( .A(n81379), .B(n85667), .Z(n91514) );
  IV U101453 ( .A(n91514), .Z(n91516) );
  IV U101454 ( .A(n81380), .Z(n81381) );
  NOR U101455 ( .A(n81382), .B(n81381), .Z(n81387) );
  IV U101456 ( .A(n81383), .Z(n81384) );
  NOR U101457 ( .A(n81385), .B(n81384), .Z(n81386) );
  NOR U101458 ( .A(n81387), .B(n81386), .Z(n87168) );
  IV U101459 ( .A(n81388), .Z(n81391) );
  IV U101460 ( .A(n81389), .Z(n81390) );
  NOR U101461 ( .A(n81391), .B(n81390), .Z(n87179) );
  IV U101462 ( .A(n87151), .Z(n87152) );
  IV U101463 ( .A(n81392), .Z(n81401) );
  IV U101464 ( .A(n81393), .Z(n81394) );
  NOR U101465 ( .A(n81401), .B(n81394), .Z(n91463) );
  IV U101466 ( .A(n81395), .Z(n81396) );
  NOR U101467 ( .A(n81397), .B(n81396), .Z(n87196) );
  NOR U101468 ( .A(n91463), .B(n87196), .Z(n85651) );
  IV U101469 ( .A(n81398), .Z(n81399) );
  NOR U101470 ( .A(n81399), .B(n81401), .Z(n91464) );
  IV U101471 ( .A(n91464), .Z(n91469) );
  IV U101472 ( .A(n81400), .Z(n81402) );
  NOR U101473 ( .A(n81402), .B(n81401), .Z(n81403) );
  IV U101474 ( .A(n81403), .Z(n91471) );
  IV U101475 ( .A(n81404), .Z(n81406) );
  NOR U101476 ( .A(n81406), .B(n81405), .Z(n81410) );
  IV U101477 ( .A(n81407), .Z(n81408) );
  NOR U101478 ( .A(n81408), .B(n81418), .Z(n81409) );
  NOR U101479 ( .A(n81410), .B(n81409), .Z(n91457) );
  IV U101480 ( .A(n81411), .Z(n81412) );
  NOR U101481 ( .A(n81418), .B(n81412), .Z(n91453) );
  IV U101482 ( .A(n81413), .Z(n81414) );
  NOR U101483 ( .A(n81415), .B(n81414), .Z(n81420) );
  IV U101484 ( .A(n81416), .Z(n81417) );
  NOR U101485 ( .A(n81418), .B(n81417), .Z(n81419) );
  NOR U101486 ( .A(n81420), .B(n81419), .Z(n87226) );
  IV U101487 ( .A(n81421), .Z(n81423) );
  NOR U101488 ( .A(n81423), .B(n81422), .Z(n81428) );
  IV U101489 ( .A(n81424), .Z(n81425) );
  NOR U101490 ( .A(n81426), .B(n81425), .Z(n81427) );
  NOR U101491 ( .A(n81428), .B(n81427), .Z(n87229) );
  IV U101492 ( .A(n81429), .Z(n81431) );
  NOR U101493 ( .A(n81431), .B(n81430), .Z(n87221) );
  IV U101494 ( .A(n81432), .Z(n81436) );
  IV U101495 ( .A(n81433), .Z(n81434) );
  NOR U101496 ( .A(n81436), .B(n81434), .Z(n87202) );
  NOR U101497 ( .A(n81436), .B(n81435), .Z(n87199) );
  IV U101498 ( .A(n81437), .Z(n81438) );
  NOR U101499 ( .A(n81438), .B(n85643), .Z(n87210) );
  IV U101500 ( .A(n81439), .Z(n81444) );
  IV U101501 ( .A(n81440), .Z(n81441) );
  NOR U101502 ( .A(n81444), .B(n81441), .Z(n87243) );
  IV U101503 ( .A(n87243), .Z(n87247) );
  IV U101504 ( .A(n81442), .Z(n81443) );
  NOR U101505 ( .A(n81444), .B(n81443), .Z(n81445) );
  IV U101506 ( .A(n81445), .Z(n87239) );
  IV U101507 ( .A(n81446), .Z(n81447) );
  NOR U101508 ( .A(n81448), .B(n81447), .Z(n85624) );
  IV U101509 ( .A(n85624), .Z(n85619) );
  IV U101510 ( .A(n81449), .Z(n81450) );
  NOR U101511 ( .A(n81451), .B(n81450), .Z(n87276) );
  IV U101512 ( .A(n81452), .Z(n81453) );
  NOR U101513 ( .A(n81454), .B(n81453), .Z(n81458) );
  IV U101514 ( .A(n81455), .Z(n81456) );
  NOR U101515 ( .A(n81456), .B(n85617), .Z(n81457) );
  NOR U101516 ( .A(n81458), .B(n81457), .Z(n87272) );
  IV U101517 ( .A(n81459), .Z(n81461) );
  NOR U101518 ( .A(n81461), .B(n81460), .Z(n81466) );
  IV U101519 ( .A(n81462), .Z(n81464) );
  NOR U101520 ( .A(n81464), .B(n81463), .Z(n81465) );
  NOR U101521 ( .A(n81466), .B(n81465), .Z(n87252) );
  IV U101522 ( .A(n81467), .Z(n81468) );
  NOR U101523 ( .A(n81469), .B(n81468), .Z(n85604) );
  IV U101524 ( .A(n81470), .Z(n81472) );
  IV U101525 ( .A(n81471), .Z(n85600) );
  NOR U101526 ( .A(n81472), .B(n85600), .Z(n87261) );
  NOR U101527 ( .A(n85597), .B(n81473), .Z(n91417) );
  IV U101528 ( .A(n81474), .Z(n81476) );
  NOR U101529 ( .A(n81476), .B(n81475), .Z(n81481) );
  IV U101530 ( .A(n81477), .Z(n81478) );
  NOR U101531 ( .A(n81479), .B(n81478), .Z(n81480) );
  NOR U101532 ( .A(n81481), .B(n81480), .Z(n91424) );
  IV U101533 ( .A(n81482), .Z(n81484) );
  NOR U101534 ( .A(n81484), .B(n81483), .Z(n81489) );
  IV U101535 ( .A(n81485), .Z(n81486) );
  NOR U101536 ( .A(n81487), .B(n81486), .Z(n81488) );
  NOR U101537 ( .A(n81489), .B(n81488), .Z(n91421) );
  IV U101538 ( .A(n81490), .Z(n81493) );
  NOR U101539 ( .A(n85579), .B(n85586), .Z(n81491) );
  IV U101540 ( .A(n81491), .Z(n81492) );
  NOR U101541 ( .A(n81493), .B(n81492), .Z(n81494) );
  IV U101542 ( .A(n81494), .Z(n91391) );
  NOR U101543 ( .A(n81495), .B(n85565), .Z(n87314) );
  IV U101544 ( .A(n81496), .Z(n81497) );
  NOR U101545 ( .A(n81497), .B(n85547), .Z(n81502) );
  IV U101546 ( .A(n81498), .Z(n81499) );
  NOR U101547 ( .A(n81500), .B(n81499), .Z(n81501) );
  NOR U101548 ( .A(n81502), .B(n81501), .Z(n91395) );
  IV U101549 ( .A(n81503), .Z(n81504) );
  NOR U101550 ( .A(n81505), .B(n81504), .Z(n87288) );
  IV U101551 ( .A(n81506), .Z(n81508) );
  NOR U101552 ( .A(n81508), .B(n81507), .Z(n87294) );
  NOR U101553 ( .A(n81510), .B(n81509), .Z(n81512) );
  NOR U101554 ( .A(n81512), .B(n81511), .Z(n87291) );
  IV U101555 ( .A(n81513), .Z(n81516) );
  IV U101556 ( .A(n81514), .Z(n81515) );
  NOR U101557 ( .A(n81516), .B(n81515), .Z(n87302) );
  IV U101558 ( .A(n81517), .Z(n81518) );
  NOR U101559 ( .A(n81518), .B(n81525), .Z(n91363) );
  IV U101560 ( .A(n81519), .Z(n81520) );
  NOR U101561 ( .A(n81520), .B(n81525), .Z(n91360) );
  IV U101562 ( .A(n81521), .Z(n81523) );
  NOR U101563 ( .A(n81523), .B(n81522), .Z(n81528) );
  IV U101564 ( .A(n81524), .Z(n81526) );
  NOR U101565 ( .A(n81526), .B(n81525), .Z(n81527) );
  NOR U101566 ( .A(n81528), .B(n81527), .Z(n91374) );
  IV U101567 ( .A(n81529), .Z(n81531) );
  NOR U101568 ( .A(n81531), .B(n81530), .Z(n91354) );
  NOR U101569 ( .A(n81533), .B(n81532), .Z(n91376) );
  NOR U101570 ( .A(n91354), .B(n91376), .Z(n85541) );
  IV U101571 ( .A(n81534), .Z(n81535) );
  NOR U101572 ( .A(n81536), .B(n81535), .Z(n91349) );
  IV U101573 ( .A(n91349), .Z(n91352) );
  IV U101574 ( .A(n81537), .Z(n81543) );
  NOR U101575 ( .A(n81538), .B(n81549), .Z(n81539) );
  IV U101576 ( .A(n81539), .Z(n81540) );
  NOR U101577 ( .A(n81541), .B(n81540), .Z(n81542) );
  IV U101578 ( .A(n81542), .Z(n81546) );
  NOR U101579 ( .A(n81543), .B(n81546), .Z(n81544) );
  IV U101580 ( .A(n81544), .Z(n91333) );
  IV U101581 ( .A(n81545), .Z(n81547) );
  NOR U101582 ( .A(n81547), .B(n81546), .Z(n91337) );
  IV U101583 ( .A(n81548), .Z(n81550) );
  NOR U101584 ( .A(n81550), .B(n81549), .Z(n91334) );
  IV U101585 ( .A(n81553), .Z(n81551) );
  NOR U101586 ( .A(n81552), .B(n81551), .Z(n81559) );
  NOR U101587 ( .A(n81554), .B(n81553), .Z(n81557) );
  IV U101588 ( .A(n81555), .Z(n81556) );
  NOR U101589 ( .A(n81557), .B(n81556), .Z(n81558) );
  NOR U101590 ( .A(n81559), .B(n81558), .Z(n91326) );
  IV U101591 ( .A(n81560), .Z(n81561) );
  NOR U101592 ( .A(n81562), .B(n81561), .Z(n91319) );
  NOR U101593 ( .A(n81564), .B(n81563), .Z(n91327) );
  NOR U101594 ( .A(n91319), .B(n91327), .Z(n85540) );
  IV U101595 ( .A(n81565), .Z(n81568) );
  NOR U101596 ( .A(n81566), .B(n81570), .Z(n81567) );
  IV U101597 ( .A(n81567), .Z(n85535) );
  NOR U101598 ( .A(n81568), .B(n85535), .Z(n91314) );
  IV U101599 ( .A(n91314), .Z(n91317) );
  IV U101600 ( .A(n81569), .Z(n81571) );
  NOR U101601 ( .A(n81571), .B(n81570), .Z(n85533) );
  IV U101602 ( .A(n85533), .Z(n87361) );
  NOR U101603 ( .A(n81573), .B(n81572), .Z(n81575) );
  NOR U101604 ( .A(n81575), .B(n81574), .Z(n81576) );
  IV U101605 ( .A(n81576), .Z(n87386) );
  IV U101606 ( .A(n81577), .Z(n81578) );
  NOR U101607 ( .A(n81579), .B(n81578), .Z(n87367) );
  IV U101608 ( .A(n81580), .Z(n81581) );
  NOR U101609 ( .A(n81582), .B(n81581), .Z(n87380) );
  NOR U101610 ( .A(n87367), .B(n87380), .Z(n85524) );
  IV U101611 ( .A(n81583), .Z(n81585) );
  NOR U101612 ( .A(n81585), .B(n81584), .Z(n87369) );
  IV U101613 ( .A(n87369), .Z(n87366) );
  NOR U101614 ( .A(n81589), .B(n81586), .Z(n81587) );
  IV U101615 ( .A(n81587), .Z(n87334) );
  NOR U101616 ( .A(n81589), .B(n81588), .Z(n87331) );
  IV U101617 ( .A(n81590), .Z(n81593) );
  IV U101618 ( .A(n81591), .Z(n81592) );
  NOR U101619 ( .A(n81593), .B(n81592), .Z(n87351) );
  IV U101620 ( .A(n81594), .Z(n81597) );
  IV U101621 ( .A(n81595), .Z(n81596) );
  NOR U101622 ( .A(n81597), .B(n81596), .Z(n87348) );
  IV U101623 ( .A(n81598), .Z(n81601) );
  IV U101624 ( .A(n81599), .Z(n81600) );
  NOR U101625 ( .A(n81601), .B(n81600), .Z(n85517) );
  IV U101626 ( .A(n81602), .Z(n81603) );
  NOR U101627 ( .A(n81604), .B(n81603), .Z(n91293) );
  NOR U101628 ( .A(n81605), .B(n85513), .Z(n91299) );
  NOR U101629 ( .A(n91293), .B(n91299), .Z(n85510) );
  IV U101630 ( .A(n81606), .Z(n81608) );
  NOR U101631 ( .A(n81608), .B(n81607), .Z(n85494) );
  IV U101632 ( .A(n85494), .Z(n87438) );
  IV U101633 ( .A(n81609), .Z(n81612) );
  NOR U101634 ( .A(n81610), .B(n81624), .Z(n81611) );
  IV U101635 ( .A(n81611), .Z(n81617) );
  NOR U101636 ( .A(n81612), .B(n81617), .Z(n87422) );
  IV U101637 ( .A(n81613), .Z(n81614) );
  NOR U101638 ( .A(n81615), .B(n81614), .Z(n87414) );
  IV U101639 ( .A(n81616), .Z(n81618) );
  NOR U101640 ( .A(n81618), .B(n81617), .Z(n87425) );
  NOR U101641 ( .A(n87414), .B(n87425), .Z(n85492) );
  IV U101642 ( .A(n81619), .Z(n81620) );
  NOR U101643 ( .A(n81621), .B(n81620), .Z(n87407) );
  IV U101644 ( .A(n81622), .Z(n81623) );
  NOR U101645 ( .A(n81624), .B(n81623), .Z(n87416) );
  NOR U101646 ( .A(n87407), .B(n87416), .Z(n85491) );
  NOR U101647 ( .A(n81626), .B(n81625), .Z(n81632) );
  NOR U101648 ( .A(n81628), .B(n81627), .Z(n81630) );
  NOR U101649 ( .A(n81630), .B(n81629), .Z(n81631) );
  NOR U101650 ( .A(n81632), .B(n81631), .Z(n81633) );
  IV U101651 ( .A(n81633), .Z(n87395) );
  IV U101652 ( .A(n81634), .Z(n81636) );
  NOR U101653 ( .A(n81636), .B(n81635), .Z(n87454) );
  IV U101654 ( .A(n81637), .Z(n81639) );
  NOR U101655 ( .A(n81639), .B(n81638), .Z(n87397) );
  NOR U101656 ( .A(n87454), .B(n87397), .Z(n85483) );
  IV U101657 ( .A(n81640), .Z(n81642) );
  IV U101658 ( .A(n81641), .Z(n81645) );
  NOR U101659 ( .A(n81642), .B(n81645), .Z(n87449) );
  IV U101660 ( .A(n87449), .Z(n87452) );
  IV U101661 ( .A(n81643), .Z(n81644) );
  NOR U101662 ( .A(n81645), .B(n81644), .Z(n81646) );
  IV U101663 ( .A(n81646), .Z(n91272) );
  IV U101664 ( .A(n81647), .Z(n81648) );
  NOR U101665 ( .A(n81649), .B(n81648), .Z(n81652) );
  NOR U101666 ( .A(n85466), .B(n81650), .Z(n81651) );
  NOR U101667 ( .A(n81652), .B(n81651), .Z(n85474) );
  IV U101668 ( .A(n85474), .Z(n85464) );
  IV U101669 ( .A(n81653), .Z(n81654) );
  NOR U101670 ( .A(n81655), .B(n81654), .Z(n81656) );
  IV U101671 ( .A(n81656), .Z(n87461) );
  IV U101672 ( .A(n81657), .Z(n81659) );
  NOR U101673 ( .A(n81659), .B(n81658), .Z(n87468) );
  IV U101674 ( .A(n81660), .Z(n81662) );
  NOR U101675 ( .A(n81662), .B(n81661), .Z(n87463) );
  NOR U101676 ( .A(n87468), .B(n87463), .Z(n85461) );
  IV U101677 ( .A(n81663), .Z(n81665) );
  IV U101678 ( .A(n81664), .Z(n85454) );
  NOR U101679 ( .A(n81665), .B(n85454), .Z(n87469) );
  NOR U101680 ( .A(n81667), .B(n81666), .Z(n87479) );
  IV U101681 ( .A(n87479), .Z(n87477) );
  IV U101682 ( .A(n81668), .Z(n81669) );
  IV U101683 ( .A(n81672), .Z(n81670) );
  NOR U101684 ( .A(n81669), .B(n81670), .Z(n91253) );
  IV U101685 ( .A(n91253), .Z(n91250) );
  IV U101686 ( .A(n81673), .Z(n81671) );
  NOR U101687 ( .A(n81671), .B(n81670), .Z(n81678) );
  NOR U101688 ( .A(n81673), .B(n81672), .Z(n81676) );
  IV U101689 ( .A(n81674), .Z(n81675) );
  NOR U101690 ( .A(n81676), .B(n81675), .Z(n81677) );
  NOR U101691 ( .A(n81678), .B(n81677), .Z(n91239) );
  IV U101692 ( .A(n81679), .Z(n81681) );
  NOR U101693 ( .A(n81681), .B(n81680), .Z(n91228) );
  NOR U101694 ( .A(n91228), .B(n81682), .Z(n85436) );
  IV U101695 ( .A(n81683), .Z(n81685) );
  NOR U101696 ( .A(n81685), .B(n81684), .Z(n91231) );
  IV U101697 ( .A(n81686), .Z(n81687) );
  NOR U101698 ( .A(n81691), .B(n81687), .Z(n81688) );
  IV U101699 ( .A(n81688), .Z(n91218) );
  IV U101700 ( .A(n81689), .Z(n81690) );
  NOR U101701 ( .A(n81691), .B(n81690), .Z(n87496) );
  IV U101702 ( .A(n81692), .Z(n81695) );
  IV U101703 ( .A(n81693), .Z(n81694) );
  NOR U101704 ( .A(n81695), .B(n81694), .Z(n87492) );
  NOR U101705 ( .A(n87496), .B(n87492), .Z(n85425) );
  IV U101706 ( .A(n81696), .Z(n81698) );
  NOR U101707 ( .A(n81698), .B(n81697), .Z(n87487) );
  IV U101708 ( .A(n81699), .Z(n81700) );
  NOR U101709 ( .A(n81705), .B(n81700), .Z(n85406) );
  IV U101710 ( .A(n81701), .Z(n81702) );
  NOR U101711 ( .A(n81703), .B(n81702), .Z(n81708) );
  IV U101712 ( .A(n81704), .Z(n81706) );
  NOR U101713 ( .A(n81706), .B(n81705), .Z(n81707) );
  NOR U101714 ( .A(n81708), .B(n81707), .Z(n91190) );
  IV U101715 ( .A(n81709), .Z(n81711) );
  IV U101716 ( .A(n81710), .Z(n81713) );
  NOR U101717 ( .A(n81711), .B(n81713), .Z(n91186) );
  IV U101718 ( .A(n81712), .Z(n81714) );
  NOR U101719 ( .A(n81714), .B(n81713), .Z(n91193) );
  IV U101720 ( .A(n81715), .Z(n81716) );
  NOR U101721 ( .A(n85399), .B(n81716), .Z(n91199) );
  IV U101722 ( .A(n81717), .Z(n81718) );
  NOR U101723 ( .A(n81718), .B(n85395), .Z(n85392) );
  IV U101724 ( .A(n85392), .Z(n85390) );
  IV U101725 ( .A(n81719), .Z(n91181) );
  NOR U101726 ( .A(n81721), .B(n81720), .Z(n81725) );
  NOR U101727 ( .A(n81723), .B(n81722), .Z(n81724) );
  NOR U101728 ( .A(n81725), .B(n81724), .Z(n91159) );
  IV U101729 ( .A(n81726), .Z(n81728) );
  NOR U101730 ( .A(n81728), .B(n81727), .Z(n81736) );
  IV U101731 ( .A(n81729), .Z(n81730) );
  NOR U101732 ( .A(n81731), .B(n81730), .Z(n81732) );
  IV U101733 ( .A(n81732), .Z(n81734) );
  NOR U101734 ( .A(n81734), .B(n81733), .Z(n81735) );
  NOR U101735 ( .A(n81736), .B(n81735), .Z(n91179) );
  IV U101736 ( .A(n81737), .Z(n81747) );
  NOR U101737 ( .A(n81747), .B(n81738), .Z(n81739) );
  IV U101738 ( .A(n81739), .Z(n81745) );
  IV U101739 ( .A(n81740), .Z(n81742) );
  NOR U101740 ( .A(n81742), .B(n81741), .Z(n81743) );
  IV U101741 ( .A(n81743), .Z(n81744) );
  NOR U101742 ( .A(n81745), .B(n81744), .Z(n91175) );
  NOR U101743 ( .A(n81747), .B(n81746), .Z(n91145) );
  IV U101744 ( .A(n81748), .Z(n81749) );
  NOR U101745 ( .A(n81749), .B(n81751), .Z(n91160) );
  IV U101746 ( .A(n81750), .Z(n81752) );
  NOR U101747 ( .A(n81752), .B(n81751), .Z(n91148) );
  IV U101748 ( .A(n81753), .Z(n81755) );
  IV U101749 ( .A(n81754), .Z(n91164) );
  NOR U101750 ( .A(n81755), .B(n91164), .Z(n81756) );
  NOR U101751 ( .A(n91148), .B(n81756), .Z(n81757) );
  IV U101752 ( .A(n81757), .Z(n85388) );
  IV U101753 ( .A(n81758), .Z(n81760) );
  NOR U101754 ( .A(n81760), .B(n81759), .Z(n81761) );
  NOR U101755 ( .A(n91134), .B(n81761), .Z(n85387) );
  IV U101756 ( .A(n81762), .Z(n81764) );
  NOR U101757 ( .A(n81764), .B(n81763), .Z(n85385) );
  IV U101758 ( .A(n85385), .Z(n85376) );
  IV U101759 ( .A(n81765), .Z(n91144) );
  IV U101760 ( .A(n81766), .Z(n81767) );
  NOR U101761 ( .A(n81767), .B(n81773), .Z(n81768) );
  IV U101762 ( .A(n81768), .Z(n87515) );
  IV U101763 ( .A(n81769), .Z(n81770) );
  NOR U101764 ( .A(n81771), .B(n81770), .Z(n81776) );
  IV U101765 ( .A(n81772), .Z(n81774) );
  NOR U101766 ( .A(n81774), .B(n81773), .Z(n81775) );
  NOR U101767 ( .A(n81776), .B(n81775), .Z(n91117) );
  IV U101768 ( .A(n81777), .Z(n81779) );
  NOR U101769 ( .A(n81779), .B(n81778), .Z(n91120) );
  IV U101770 ( .A(n81780), .Z(n81782) );
  NOR U101771 ( .A(n81782), .B(n81781), .Z(n91098) );
  NOR U101772 ( .A(n91120), .B(n91098), .Z(n85360) );
  IV U101773 ( .A(n81783), .Z(n81784) );
  NOR U101774 ( .A(n85357), .B(n81784), .Z(n81785) );
  IV U101775 ( .A(n81785), .Z(n91101) );
  IV U101776 ( .A(n81786), .Z(n81789) );
  IV U101777 ( .A(n81787), .Z(n81788) );
  NOR U101778 ( .A(n81789), .B(n81788), .Z(n81790) );
  NOR U101779 ( .A(n81791), .B(n81790), .Z(n87522) );
  IV U101780 ( .A(n81792), .Z(n81793) );
  NOR U101781 ( .A(n85344), .B(n81793), .Z(n91090) );
  IV U101782 ( .A(n81794), .Z(n81795) );
  NOR U101783 ( .A(n81795), .B(n85324), .Z(n91076) );
  IV U101784 ( .A(n81796), .Z(n81798) );
  NOR U101785 ( .A(n81798), .B(n81797), .Z(n87531) );
  IV U101786 ( .A(n81799), .Z(n81800) );
  NOR U101787 ( .A(n81801), .B(n81800), .Z(n81806) );
  IV U101788 ( .A(n81802), .Z(n81803) );
  NOR U101789 ( .A(n81804), .B(n81803), .Z(n81805) );
  NOR U101790 ( .A(n81806), .B(n81805), .Z(n91049) );
  IV U101791 ( .A(n81807), .Z(n85309) );
  IV U101792 ( .A(n81808), .Z(n81809) );
  NOR U101793 ( .A(n85309), .B(n81809), .Z(n85313) );
  NOR U101794 ( .A(n81811), .B(n81810), .Z(n81816) );
  NOR U101795 ( .A(n81812), .B(n85301), .Z(n81813) );
  NOR U101796 ( .A(n81814), .B(n81813), .Z(n81815) );
  NOR U101797 ( .A(n81816), .B(n81815), .Z(n91039) );
  IV U101798 ( .A(n81817), .Z(n81819) );
  NOR U101799 ( .A(n81819), .B(n81818), .Z(n91059) );
  IV U101800 ( .A(n81820), .Z(n81821) );
  NOR U101801 ( .A(n81824), .B(n81821), .Z(n91056) );
  IV U101802 ( .A(n81822), .Z(n81823) );
  NOR U101803 ( .A(n81824), .B(n81823), .Z(n91003) );
  IV U101804 ( .A(n81825), .Z(n81828) );
  IV U101805 ( .A(n81826), .Z(n81827) );
  NOR U101806 ( .A(n81828), .B(n81827), .Z(n91000) );
  IV U101807 ( .A(n81829), .Z(n81832) );
  XOR U101808 ( .A(n81830), .B(n87539), .Z(n81831) );
  NOR U101809 ( .A(n81832), .B(n81831), .Z(n91014) );
  IV U101810 ( .A(n81833), .Z(n81834) );
  NOR U101811 ( .A(n81834), .B(n87539), .Z(n91011) );
  NOR U101812 ( .A(n81835), .B(n87539), .Z(n85280) );
  IV U101813 ( .A(n81836), .Z(n81837) );
  NOR U101814 ( .A(n81838), .B(n81837), .Z(n81843) );
  IV U101815 ( .A(n81839), .Z(n81841) );
  NOR U101816 ( .A(n81841), .B(n81840), .Z(n81842) );
  NOR U101817 ( .A(n81843), .B(n81842), .Z(n87547) );
  IV U101818 ( .A(n87547), .Z(n85279) );
  IV U101819 ( .A(n81844), .Z(n85278) );
  NOR U101820 ( .A(n81845), .B(n85278), .Z(n87550) );
  IV U101821 ( .A(n81846), .Z(n81847) );
  NOR U101822 ( .A(n85269), .B(n81847), .Z(n85262) );
  IV U101823 ( .A(n81848), .Z(n81849) );
  NOR U101824 ( .A(n81850), .B(n81849), .Z(n81851) );
  IV U101825 ( .A(n81851), .Z(n87564) );
  NOR U101826 ( .A(n81852), .B(n85259), .Z(n81859) );
  IV U101827 ( .A(n85259), .Z(n81853) );
  NOR U101828 ( .A(n81854), .B(n81853), .Z(n81857) );
  IV U101829 ( .A(n81855), .Z(n81856) );
  NOR U101830 ( .A(n81857), .B(n81856), .Z(n81858) );
  NOR U101831 ( .A(n81859), .B(n81858), .Z(n87577) );
  IV U101832 ( .A(n81860), .Z(n81861) );
  NOR U101833 ( .A(n81862), .B(n81861), .Z(n87570) );
  IV U101834 ( .A(n81863), .Z(n81865) );
  NOR U101835 ( .A(n81865), .B(n81864), .Z(n81870) );
  IV U101836 ( .A(n81866), .Z(n81868) );
  NOR U101837 ( .A(n81868), .B(n81867), .Z(n81869) );
  NOR U101838 ( .A(n81870), .B(n81869), .Z(n87568) );
  IV U101839 ( .A(n87568), .Z(n85250) );
  IV U101840 ( .A(n81871), .Z(n81872) );
  NOR U101841 ( .A(n81875), .B(n81872), .Z(n87588) );
  IV U101842 ( .A(n81873), .Z(n81874) );
  NOR U101843 ( .A(n81875), .B(n81874), .Z(n87585) );
  IV U101844 ( .A(n81876), .Z(n81878) );
  IV U101845 ( .A(n81877), .Z(n81880) );
  NOR U101846 ( .A(n81878), .B(n81880), .Z(n87615) );
  IV U101847 ( .A(n81879), .Z(n81881) );
  NOR U101848 ( .A(n81881), .B(n81880), .Z(n87612) );
  IV U101849 ( .A(n81882), .Z(n81883) );
  NOR U101850 ( .A(n81883), .B(n85247), .Z(n85244) );
  IV U101851 ( .A(n85244), .Z(n85238) );
  IV U101852 ( .A(n81884), .Z(n81885) );
  NOR U101853 ( .A(n81886), .B(n81885), .Z(n90975) );
  IV U101854 ( .A(n81887), .Z(n81891) );
  NOR U101855 ( .A(n81889), .B(n81888), .Z(n81890) );
  IV U101856 ( .A(n81890), .Z(n81893) );
  NOR U101857 ( .A(n81891), .B(n81893), .Z(n90972) );
  IV U101858 ( .A(n81892), .Z(n81894) );
  NOR U101859 ( .A(n81894), .B(n81893), .Z(n87623) );
  IV U101860 ( .A(n81895), .Z(n81896) );
  NOR U101861 ( .A(n81898), .B(n81896), .Z(n87620) );
  IV U101862 ( .A(n81897), .Z(n81899) );
  NOR U101863 ( .A(n81899), .B(n81898), .Z(n90953) );
  IV U101864 ( .A(n81900), .Z(n81902) );
  NOR U101865 ( .A(n81902), .B(n81901), .Z(n90950) );
  IV U101866 ( .A(n81903), .Z(n81907) );
  IV U101867 ( .A(n81904), .Z(n81911) );
  NOR U101868 ( .A(n81905), .B(n81911), .Z(n81906) );
  IV U101869 ( .A(n81906), .Z(n81909) );
  NOR U101870 ( .A(n81907), .B(n81909), .Z(n90961) );
  IV U101871 ( .A(n81908), .Z(n81910) );
  NOR U101872 ( .A(n81910), .B(n81909), .Z(n90958) );
  NOR U101873 ( .A(n81912), .B(n81911), .Z(n85234) );
  IV U101874 ( .A(n85234), .Z(n85226) );
  IV U101875 ( .A(n81913), .Z(n81914) );
  NOR U101876 ( .A(n85230), .B(n81914), .Z(n87631) );
  IV U101877 ( .A(n81915), .Z(n81917) );
  NOR U101878 ( .A(n81917), .B(n81916), .Z(n81918) );
  IV U101879 ( .A(n81918), .Z(n87628) );
  IV U101880 ( .A(n81919), .Z(n81921) );
  NOR U101881 ( .A(n81921), .B(n81920), .Z(n90935) );
  IV U101882 ( .A(n81922), .Z(n81925) );
  NOR U101883 ( .A(n85218), .B(n81923), .Z(n81924) );
  IV U101884 ( .A(n81924), .Z(n85220) );
  NOR U101885 ( .A(n81925), .B(n85220), .Z(n90932) );
  IV U101886 ( .A(n81926), .Z(n81934) );
  IV U101887 ( .A(n81927), .Z(n81928) );
  NOR U101888 ( .A(n81934), .B(n81928), .Z(n81929) );
  IV U101889 ( .A(n81929), .Z(n87653) );
  IV U101890 ( .A(n81930), .Z(n81931) );
  NOR U101891 ( .A(n81931), .B(n85204), .Z(n87643) );
  IV U101892 ( .A(n81932), .Z(n81933) );
  NOR U101893 ( .A(n81934), .B(n81933), .Z(n87638) );
  NOR U101894 ( .A(n87643), .B(n87638), .Z(n85215) );
  IV U101895 ( .A(n81935), .Z(n81936) );
  NOR U101896 ( .A(n81937), .B(n81936), .Z(n85198) );
  IV U101897 ( .A(n85198), .Z(n85186) );
  IV U101898 ( .A(n81938), .Z(n81939) );
  NOR U101899 ( .A(n81939), .B(n85174), .Z(n85194) );
  IV U101900 ( .A(n81940), .Z(n81942) );
  NOR U101901 ( .A(n81942), .B(n81941), .Z(n90874) );
  IV U101902 ( .A(n81943), .Z(n81948) );
  NOR U101903 ( .A(n81952), .B(n81944), .Z(n81945) );
  IV U101904 ( .A(n81945), .Z(n81954) );
  NOR U101905 ( .A(n81946), .B(n81954), .Z(n81947) );
  IV U101906 ( .A(n81947), .Z(n85172) );
  NOR U101907 ( .A(n81948), .B(n85172), .Z(n81949) );
  IV U101908 ( .A(n81949), .Z(n90884) );
  IV U101909 ( .A(n81950), .Z(n81951) );
  NOR U101910 ( .A(n81952), .B(n81951), .Z(n81957) );
  IV U101911 ( .A(n81953), .Z(n81955) );
  NOR U101912 ( .A(n81955), .B(n81954), .Z(n81956) );
  NOR U101913 ( .A(n81957), .B(n81956), .Z(n87670) );
  IV U101914 ( .A(n81958), .Z(n81960) );
  IV U101915 ( .A(n81959), .Z(n81962) );
  NOR U101916 ( .A(n81960), .B(n81962), .Z(n87694) );
  IV U101917 ( .A(n81961), .Z(n81965) );
  NOR U101918 ( .A(n81963), .B(n81962), .Z(n81964) );
  IV U101919 ( .A(n81964), .Z(n81967) );
  NOR U101920 ( .A(n81965), .B(n81967), .Z(n87691) );
  IV U101921 ( .A(n81966), .Z(n81968) );
  NOR U101922 ( .A(n81968), .B(n81967), .Z(n87664) );
  IV U101923 ( .A(n81969), .Z(n81973) );
  NOR U101924 ( .A(n81971), .B(n81970), .Z(n81972) );
  IV U101925 ( .A(n81972), .Z(n81975) );
  NOR U101926 ( .A(n81973), .B(n81975), .Z(n87661) );
  IV U101927 ( .A(n81974), .Z(n81976) );
  NOR U101928 ( .A(n81976), .B(n81975), .Z(n87702) );
  NOR U101929 ( .A(n81978), .B(n81977), .Z(n81979) );
  IV U101930 ( .A(n81979), .Z(n81980) );
  NOR U101931 ( .A(n81981), .B(n81980), .Z(n87699) );
  IV U101932 ( .A(n81982), .Z(n81985) );
  IV U101933 ( .A(n81983), .Z(n81984) );
  NOR U101934 ( .A(n81985), .B(n81984), .Z(n87676) );
  IV U101935 ( .A(n81986), .Z(n81987) );
  NOR U101936 ( .A(n81987), .B(n81994), .Z(n87673) );
  NOR U101937 ( .A(n81989), .B(n81988), .Z(n87684) );
  IV U101938 ( .A(n81990), .Z(n81992) );
  NOR U101939 ( .A(n81992), .B(n81991), .Z(n87707) );
  IV U101940 ( .A(n81993), .Z(n81995) );
  NOR U101941 ( .A(n81995), .B(n81994), .Z(n87682) );
  NOR U101942 ( .A(n87707), .B(n87682), .Z(n85170) );
  IV U101943 ( .A(n81996), .Z(n81997) );
  NOR U101944 ( .A(n81997), .B(n82000), .Z(n90843) );
  IV U101945 ( .A(n90843), .Z(n90846) );
  IV U101946 ( .A(n81998), .Z(n81999) );
  NOR U101947 ( .A(n82000), .B(n81999), .Z(n90852) );
  IV U101948 ( .A(n82001), .Z(n82003) );
  NOR U101949 ( .A(n82003), .B(n82002), .Z(n87717) );
  IV U101950 ( .A(n82004), .Z(n82005) );
  NOR U101951 ( .A(n85143), .B(n82005), .Z(n90821) );
  IV U101952 ( .A(n82006), .Z(n82008) );
  NOR U101953 ( .A(n82008), .B(n82007), .Z(n87739) );
  IV U101954 ( .A(n82009), .Z(n82010) );
  NOR U101955 ( .A(n82011), .B(n82010), .Z(n90830) );
  IV U101956 ( .A(n82012), .Z(n82014) );
  NOR U101957 ( .A(n82014), .B(n82013), .Z(n90832) );
  XOR U101958 ( .A(n90830), .B(n90832), .Z(n82015) );
  NOR U101959 ( .A(n87739), .B(n82015), .Z(n85140) );
  IV U101960 ( .A(n82016), .Z(n82022) );
  NOR U101961 ( .A(n82017), .B(n82025), .Z(n82018) );
  IV U101962 ( .A(n82018), .Z(n82019) );
  NOR U101963 ( .A(n82020), .B(n82019), .Z(n82021) );
  IV U101964 ( .A(n82021), .Z(n82027) );
  NOR U101965 ( .A(n82022), .B(n82027), .Z(n85127) );
  IV U101966 ( .A(n85127), .Z(n90804) );
  IV U101967 ( .A(n82023), .Z(n82024) );
  NOR U101968 ( .A(n82025), .B(n82024), .Z(n82030) );
  IV U101969 ( .A(n82026), .Z(n82028) );
  NOR U101970 ( .A(n82028), .B(n82027), .Z(n82029) );
  NOR U101971 ( .A(n82030), .B(n82029), .Z(n90797) );
  IV U101972 ( .A(n82031), .Z(n82032) );
  NOR U101973 ( .A(n82033), .B(n82032), .Z(n82038) );
  IV U101974 ( .A(n82034), .Z(n82035) );
  NOR U101975 ( .A(n82036), .B(n82035), .Z(n82037) );
  NOR U101976 ( .A(n82038), .B(n82037), .Z(n87736) );
  IV U101977 ( .A(n82039), .Z(n82048) );
  NOR U101978 ( .A(n82054), .B(n82040), .Z(n82041) );
  IV U101979 ( .A(n82041), .Z(n82046) );
  NOR U101980 ( .A(n82043), .B(n82042), .Z(n82044) );
  IV U101981 ( .A(n82044), .Z(n82045) );
  NOR U101982 ( .A(n82046), .B(n82045), .Z(n82047) );
  IV U101983 ( .A(n82047), .Z(n82050) );
  NOR U101984 ( .A(n82048), .B(n82050), .Z(n87732) );
  IV U101985 ( .A(n82049), .Z(n82051) );
  NOR U101986 ( .A(n82051), .B(n82050), .Z(n87792) );
  IV U101987 ( .A(n82052), .Z(n82053) );
  NOR U101988 ( .A(n82054), .B(n82053), .Z(n87789) );
  IV U101989 ( .A(n82055), .Z(n82059) );
  IV U101990 ( .A(n82056), .Z(n82062) );
  NOR U101991 ( .A(n82057), .B(n82062), .Z(n82058) );
  IV U101992 ( .A(n82058), .Z(n85110) );
  NOR U101993 ( .A(n82059), .B(n85110), .Z(n87746) );
  IV U101994 ( .A(n82060), .Z(n82061) );
  NOR U101995 ( .A(n82062), .B(n82061), .Z(n85113) );
  IV U101996 ( .A(n82063), .Z(n82066) );
  IV U101997 ( .A(n82064), .Z(n82065) );
  NOR U101998 ( .A(n82066), .B(n82065), .Z(n82068) );
  NOR U101999 ( .A(n82068), .B(n82067), .Z(n82069) );
  IV U102000 ( .A(n82069), .Z(n82070) );
  NOR U102001 ( .A(n82071), .B(n82070), .Z(n87788) );
  NOR U102002 ( .A(n82072), .B(n85105), .Z(n82074) );
  NOR U102003 ( .A(n82074), .B(n82073), .Z(n87755) );
  IV U102004 ( .A(n87755), .Z(n85107) );
  IV U102005 ( .A(n82075), .Z(n82076) );
  NOR U102006 ( .A(n82077), .B(n82076), .Z(n85095) );
  IV U102007 ( .A(n85095), .Z(n85090) );
  IV U102008 ( .A(n82078), .Z(n85093) );
  IV U102009 ( .A(n82079), .Z(n82080) );
  NOR U102010 ( .A(n85093), .B(n82080), .Z(n82081) );
  IV U102011 ( .A(n82081), .Z(n87762) );
  IV U102012 ( .A(n82082), .Z(n82083) );
  NOR U102013 ( .A(n82084), .B(n82083), .Z(n87758) );
  IV U102014 ( .A(n82088), .Z(n82085) );
  NOR U102015 ( .A(n82085), .B(n82086), .Z(n82093) );
  IV U102016 ( .A(n82086), .Z(n82087) );
  NOR U102017 ( .A(n82088), .B(n82087), .Z(n82091) );
  IV U102018 ( .A(n82089), .Z(n82090) );
  NOR U102019 ( .A(n82091), .B(n82090), .Z(n82092) );
  NOR U102020 ( .A(n82093), .B(n82092), .Z(n87803) );
  IV U102021 ( .A(n82094), .Z(n82095) );
  NOR U102022 ( .A(n82096), .B(n82095), .Z(n87816) );
  IV U102023 ( .A(n82097), .Z(n82099) );
  NOR U102024 ( .A(n82099), .B(n82098), .Z(n87804) );
  NOR U102025 ( .A(n87816), .B(n87804), .Z(n85089) );
  IV U102026 ( .A(n82100), .Z(n82105) );
  IV U102027 ( .A(n82101), .Z(n82102) );
  NOR U102028 ( .A(n82105), .B(n82102), .Z(n87811) );
  IV U102029 ( .A(n82103), .Z(n82104) );
  NOR U102030 ( .A(n82105), .B(n82104), .Z(n87808) );
  IV U102031 ( .A(n82106), .Z(n82107) );
  NOR U102032 ( .A(n82108), .B(n82107), .Z(n87841) );
  XOR U102033 ( .A(n82109), .B(n82114), .Z(n82112) );
  IV U102034 ( .A(n82110), .Z(n82111) );
  NOR U102035 ( .A(n82112), .B(n82111), .Z(n87838) );
  IV U102036 ( .A(n82113), .Z(n82117) );
  IV U102037 ( .A(n82114), .Z(n82122) );
  NOR U102038 ( .A(n82115), .B(n82122), .Z(n82116) );
  IV U102039 ( .A(n82116), .Z(n82119) );
  NOR U102040 ( .A(n82117), .B(n82119), .Z(n90775) );
  IV U102041 ( .A(n82118), .Z(n82120) );
  NOR U102042 ( .A(n82120), .B(n82119), .Z(n90781) );
  IV U102043 ( .A(n82121), .Z(n82123) );
  NOR U102044 ( .A(n82123), .B(n82122), .Z(n90778) );
  IV U102045 ( .A(n82124), .Z(n82127) );
  IV U102046 ( .A(n82125), .Z(n82126) );
  NOR U102047 ( .A(n82127), .B(n82126), .Z(n87849) );
  NOR U102048 ( .A(n82129), .B(n82128), .Z(n87821) );
  IV U102049 ( .A(n82130), .Z(n82132) );
  NOR U102050 ( .A(n82132), .B(n82131), .Z(n87829) );
  IV U102051 ( .A(n82133), .Z(n82134) );
  NOR U102052 ( .A(n82135), .B(n82134), .Z(n85067) );
  IV U102053 ( .A(n82136), .Z(n82139) );
  NOR U102054 ( .A(n82137), .B(n82141), .Z(n82138) );
  IV U102055 ( .A(n82138), .Z(n85063) );
  NOR U102056 ( .A(n82139), .B(n85063), .Z(n87865) );
  IV U102057 ( .A(n82140), .Z(n82142) );
  NOR U102058 ( .A(n82142), .B(n82141), .Z(n87854) );
  IV U102059 ( .A(n82143), .Z(n82145) );
  NOR U102060 ( .A(n82145), .B(n82144), .Z(n82146) );
  IV U102061 ( .A(n82146), .Z(n85042) );
  IV U102062 ( .A(n82147), .Z(n82148) );
  NOR U102063 ( .A(n82149), .B(n82148), .Z(n90756) );
  NOR U102064 ( .A(n85031), .B(n82150), .Z(n90753) );
  IV U102065 ( .A(n82151), .Z(n82152) );
  NOR U102066 ( .A(n82158), .B(n82152), .Z(n82156) );
  NOR U102067 ( .A(n82154), .B(n82153), .Z(n82155) );
  NOR U102068 ( .A(n82156), .B(n82155), .Z(n87908) );
  IV U102069 ( .A(n82157), .Z(n82161) );
  NOR U102070 ( .A(n82159), .B(n82158), .Z(n82160) );
  IV U102071 ( .A(n82160), .Z(n85006) );
  NOR U102072 ( .A(n82161), .B(n85006), .Z(n85015) );
  IV U102073 ( .A(n82162), .Z(n82165) );
  IV U102074 ( .A(n82163), .Z(n82164) );
  NOR U102075 ( .A(n82165), .B(n82164), .Z(n87889) );
  IV U102076 ( .A(n82166), .Z(n82167) );
  NOR U102077 ( .A(n82167), .B(n82169), .Z(n90733) );
  IV U102078 ( .A(n82168), .Z(n82170) );
  NOR U102079 ( .A(n82170), .B(n82169), .Z(n84988) );
  IV U102080 ( .A(n84988), .Z(n84982) );
  IV U102081 ( .A(n82171), .Z(n82173) );
  NOR U102082 ( .A(n82173), .B(n82172), .Z(n90738) );
  IV U102083 ( .A(n82174), .Z(n82176) );
  NOR U102084 ( .A(n82176), .B(n82175), .Z(n82181) );
  IV U102085 ( .A(n82177), .Z(n82178) );
  NOR U102086 ( .A(n82179), .B(n82178), .Z(n82180) );
  NOR U102087 ( .A(n82181), .B(n82180), .Z(n87956) );
  IV U102088 ( .A(n82182), .Z(n82183) );
  NOR U102089 ( .A(n84962), .B(n82183), .Z(n87972) );
  IV U102090 ( .A(n82184), .Z(n82188) );
  IV U102091 ( .A(n82185), .Z(n82190) );
  NOR U102092 ( .A(n82186), .B(n82190), .Z(n82187) );
  IV U102093 ( .A(n82187), .Z(n84931) );
  NOR U102094 ( .A(n82188), .B(n84931), .Z(n84949) );
  IV U102095 ( .A(n82189), .Z(n82193) );
  NOR U102096 ( .A(n82191), .B(n82190), .Z(n82192) );
  IV U102097 ( .A(n82192), .Z(n84918) );
  NOR U102098 ( .A(n82193), .B(n84918), .Z(n84938) );
  IV U102099 ( .A(n82194), .Z(n82197) );
  NOR U102100 ( .A(n84910), .B(n82195), .Z(n82196) );
  IV U102101 ( .A(n82196), .Z(n82199) );
  NOR U102102 ( .A(n82197), .B(n82199), .Z(n84921) );
  IV U102103 ( .A(n82198), .Z(n82200) );
  NOR U102104 ( .A(n82200), .B(n82199), .Z(n87942) );
  IV U102105 ( .A(n82201), .Z(n82203) );
  NOR U102106 ( .A(n82203), .B(n82202), .Z(n84907) );
  IV U102107 ( .A(n84907), .Z(n87948) );
  IV U102108 ( .A(n82204), .Z(n82205) );
  NOR U102109 ( .A(n82205), .B(n82210), .Z(n87930) );
  IV U102110 ( .A(n82206), .Z(n82207) );
  NOR U102111 ( .A(n82208), .B(n82207), .Z(n82213) );
  IV U102112 ( .A(n82209), .Z(n82211) );
  NOR U102113 ( .A(n82211), .B(n82210), .Z(n82212) );
  NOR U102114 ( .A(n82213), .B(n82212), .Z(n88009) );
  IV U102115 ( .A(n82214), .Z(n84890) );
  IV U102116 ( .A(n82215), .Z(n82216) );
  NOR U102117 ( .A(n84890), .B(n82216), .Z(n88015) );
  IV U102118 ( .A(n82217), .Z(n82218) );
  NOR U102119 ( .A(n84890), .B(n82218), .Z(n88012) );
  IV U102120 ( .A(n82219), .Z(n82220) );
  NOR U102121 ( .A(n84890), .B(n82220), .Z(n87982) );
  IV U102122 ( .A(n82221), .Z(n82222) );
  NOR U102123 ( .A(n84859), .B(n82222), .Z(n84878) );
  IV U102124 ( .A(n82223), .Z(n82226) );
  IV U102125 ( .A(n82224), .Z(n82225) );
  NOR U102126 ( .A(n82226), .B(n82225), .Z(n84861) );
  IV U102127 ( .A(n82227), .Z(n82228) );
  NOR U102128 ( .A(n82229), .B(n82228), .Z(n82230) );
  NOR U102129 ( .A(n82231), .B(n82230), .Z(n88063) );
  IV U102130 ( .A(n82232), .Z(n82233) );
  NOR U102131 ( .A(n82233), .B(n82235), .Z(n88059) );
  IV U102132 ( .A(n82234), .Z(n82236) );
  NOR U102133 ( .A(n82236), .B(n82235), .Z(n82237) );
  IV U102134 ( .A(n82237), .Z(n88025) );
  IV U102135 ( .A(n82238), .Z(n82239) );
  NOR U102136 ( .A(n82239), .B(n84841), .Z(n88033) );
  IV U102137 ( .A(n88033), .Z(n88037) );
  IV U102138 ( .A(n82240), .Z(n82241) );
  NOR U102139 ( .A(n82242), .B(n82241), .Z(n82246) );
  IV U102140 ( .A(n82243), .Z(n82244) );
  NOR U102141 ( .A(n82251), .B(n82244), .Z(n82245) );
  NOR U102142 ( .A(n82246), .B(n82245), .Z(n88040) );
  IV U102143 ( .A(n82247), .Z(n82256) );
  IV U102144 ( .A(n82248), .Z(n82249) );
  NOR U102145 ( .A(n82256), .B(n82249), .Z(n88054) );
  IV U102146 ( .A(n82250), .Z(n82252) );
  NOR U102147 ( .A(n82252), .B(n82251), .Z(n88042) );
  NOR U102148 ( .A(n88054), .B(n88042), .Z(n82253) );
  IV U102149 ( .A(n82253), .Z(n84838) );
  IV U102150 ( .A(n82254), .Z(n82255) );
  NOR U102151 ( .A(n82256), .B(n82255), .Z(n88049) );
  IV U102152 ( .A(n88049), .Z(n88052) );
  IV U102153 ( .A(n82257), .Z(n82259) );
  NOR U102154 ( .A(n82259), .B(n82258), .Z(n90709) );
  IV U102155 ( .A(n82260), .Z(n82262) );
  NOR U102156 ( .A(n82262), .B(n82261), .Z(n84836) );
  IV U102157 ( .A(n84836), .Z(n84821) );
  IV U102158 ( .A(n82263), .Z(n82264) );
  NOR U102159 ( .A(n82264), .B(n82270), .Z(n82268) );
  NOR U102160 ( .A(n82266), .B(n82265), .Z(n82267) );
  NOR U102161 ( .A(n82268), .B(n82267), .Z(n90671) );
  IV U102162 ( .A(n82269), .Z(n82271) );
  NOR U102163 ( .A(n82271), .B(n82270), .Z(n82272) );
  IV U102164 ( .A(n82272), .Z(n90668) );
  IV U102165 ( .A(n82273), .Z(n82274) );
  NOR U102166 ( .A(n82275), .B(n82274), .Z(n82279) );
  NOR U102167 ( .A(n82277), .B(n82276), .Z(n82278) );
  NOR U102168 ( .A(n82279), .B(n82278), .Z(n90688) );
  IV U102169 ( .A(n82280), .Z(n82282) );
  NOR U102170 ( .A(n82282), .B(n82281), .Z(n82287) );
  IV U102171 ( .A(n82283), .Z(n82284) );
  NOR U102172 ( .A(n82285), .B(n82284), .Z(n82286) );
  NOR U102173 ( .A(n82287), .B(n82286), .Z(n90676) );
  IV U102174 ( .A(n82288), .Z(n82290) );
  NOR U102175 ( .A(n82290), .B(n82289), .Z(n82295) );
  IV U102176 ( .A(n82291), .Z(n82292) );
  NOR U102177 ( .A(n82293), .B(n82292), .Z(n82294) );
  NOR U102178 ( .A(n82295), .B(n82294), .Z(n90656) );
  IV U102179 ( .A(n82296), .Z(n82298) );
  NOR U102180 ( .A(n82298), .B(n82297), .Z(n82299) );
  IV U102181 ( .A(n82299), .Z(n88082) );
  IV U102182 ( .A(n82300), .Z(n82301) );
  NOR U102183 ( .A(n84793), .B(n82301), .Z(n84788) );
  IV U102184 ( .A(n82302), .Z(n82306) );
  NOR U102185 ( .A(n82304), .B(n82303), .Z(n82305) );
  IV U102186 ( .A(n82305), .Z(n84753) );
  NOR U102187 ( .A(n82306), .B(n84753), .Z(n84760) );
  IV U102188 ( .A(n84760), .Z(n84757) );
  NOR U102189 ( .A(n82308), .B(n82307), .Z(n88137) );
  IV U102190 ( .A(n82309), .Z(n82310) );
  NOR U102191 ( .A(n82310), .B(n88113), .Z(n82311) );
  IV U102192 ( .A(n82311), .Z(n82312) );
  NOR U102193 ( .A(n82313), .B(n82312), .Z(n88110) );
  IV U102194 ( .A(n82314), .Z(n84720) );
  IV U102195 ( .A(n82315), .Z(n82316) );
  NOR U102196 ( .A(n84720), .B(n82316), .Z(n88104) );
  IV U102197 ( .A(n82317), .Z(n82322) );
  XOR U102198 ( .A(n84718), .B(n84720), .Z(n82318) );
  NOR U102199 ( .A(n82319), .B(n82318), .Z(n82320) );
  IV U102200 ( .A(n82320), .Z(n82321) );
  NOR U102201 ( .A(n82322), .B(n82321), .Z(n88123) );
  NOR U102202 ( .A(n88104), .B(n88123), .Z(n84725) );
  IV U102203 ( .A(n82323), .Z(n82324) );
  NOR U102204 ( .A(n82324), .B(n84722), .Z(n82325) );
  IV U102205 ( .A(n82325), .Z(n90592) );
  IV U102206 ( .A(n82326), .Z(n82330) );
  XOR U102207 ( .A(n82330), .B(n82329), .Z(n82327) );
  NOR U102208 ( .A(n82328), .B(n82327), .Z(n90588) );
  IV U102209 ( .A(n82329), .Z(n84710) );
  NOR U102210 ( .A(n84710), .B(n82330), .Z(n90595) );
  NOR U102211 ( .A(n82332), .B(n82331), .Z(n82333) );
  IV U102212 ( .A(n82333), .Z(n90608) );
  IV U102213 ( .A(n82337), .Z(n82335) );
  NOR U102214 ( .A(n82335), .B(n82334), .Z(n82342) );
  NOR U102215 ( .A(n82337), .B(n82336), .Z(n82340) );
  IV U102216 ( .A(n82338), .Z(n82339) );
  NOR U102217 ( .A(n82340), .B(n82339), .Z(n82341) );
  NOR U102218 ( .A(n82342), .B(n82341), .Z(n90605) );
  IV U102219 ( .A(n82343), .Z(n82345) );
  NOR U102220 ( .A(n82345), .B(n82344), .Z(n82356) );
  IV U102221 ( .A(n82346), .Z(n82348) );
  NOR U102222 ( .A(n82348), .B(n82347), .Z(n82353) );
  IV U102223 ( .A(n82349), .Z(n82351) );
  NOR U102224 ( .A(n82351), .B(n82350), .Z(n82352) );
  NOR U102225 ( .A(n82353), .B(n82352), .Z(n82354) );
  IV U102226 ( .A(n82354), .Z(n82355) );
  NOR U102227 ( .A(n82356), .B(n82355), .Z(n90576) );
  IV U102228 ( .A(n82357), .Z(n82359) );
  NOR U102229 ( .A(n82359), .B(n82358), .Z(n88162) );
  IV U102230 ( .A(n82360), .Z(n82361) );
  NOR U102231 ( .A(n82361), .B(n84685), .Z(n82366) );
  IV U102232 ( .A(n82362), .Z(n82363) );
  NOR U102233 ( .A(n82364), .B(n82363), .Z(n82365) );
  NOR U102234 ( .A(n82366), .B(n82365), .Z(n88170) );
  IV U102235 ( .A(n88170), .Z(n84683) );
  IV U102236 ( .A(n82367), .Z(n82369) );
  NOR U102237 ( .A(n82369), .B(n82368), .Z(n88179) );
  IV U102238 ( .A(n82370), .Z(n82371) );
  NOR U102239 ( .A(n82372), .B(n82371), .Z(n88176) );
  IV U102240 ( .A(n82373), .Z(n82374) );
  NOR U102241 ( .A(n82374), .B(n82376), .Z(n90552) );
  IV U102242 ( .A(n82375), .Z(n82377) );
  NOR U102243 ( .A(n82377), .B(n82376), .Z(n82378) );
  IV U102244 ( .A(n82378), .Z(n90551) );
  IV U102245 ( .A(n82379), .Z(n82381) );
  NOR U102246 ( .A(n82381), .B(n82380), .Z(n84672) );
  IV U102247 ( .A(n82382), .Z(n82386) );
  IV U102248 ( .A(n82383), .Z(n82384) );
  NOR U102249 ( .A(n82386), .B(n82384), .Z(n88189) );
  NOR U102250 ( .A(n82386), .B(n82385), .Z(n88194) );
  IV U102251 ( .A(n82387), .Z(n82389) );
  NOR U102252 ( .A(n82389), .B(n82388), .Z(n88196) );
  XOR U102253 ( .A(n88194), .B(n88196), .Z(n82390) );
  NOR U102254 ( .A(n88189), .B(n82390), .Z(n84666) );
  NOR U102255 ( .A(n82392), .B(n82391), .Z(n82397) );
  IV U102256 ( .A(n82393), .Z(n82395) );
  XOR U102257 ( .A(n82395), .B(n82394), .Z(n82396) );
  NOR U102258 ( .A(n82397), .B(n82396), .Z(n88186) );
  IV U102259 ( .A(n82398), .Z(n82399) );
  NOR U102260 ( .A(n82399), .B(n84651), .Z(n90535) );
  IV U102261 ( .A(n82400), .Z(n82401) );
  NOR U102262 ( .A(n82406), .B(n82401), .Z(n88206) );
  IV U102263 ( .A(n82402), .Z(n82403) );
  NOR U102264 ( .A(n82403), .B(n82406), .Z(n90506) );
  IV U102265 ( .A(n82407), .Z(n82404) );
  NOR U102266 ( .A(n82406), .B(n82404), .Z(n90516) );
  IV U102267 ( .A(n82405), .Z(n82409) );
  XOR U102268 ( .A(n82407), .B(n82406), .Z(n82408) );
  NOR U102269 ( .A(n82409), .B(n82408), .Z(n90509) );
  NOR U102270 ( .A(n90516), .B(n90509), .Z(n84646) );
  IV U102271 ( .A(n82410), .Z(n82412) );
  NOR U102272 ( .A(n82412), .B(n82411), .Z(n84644) );
  IV U102273 ( .A(n84644), .Z(n84635) );
  IV U102274 ( .A(n82413), .Z(n82415) );
  IV U102275 ( .A(n82414), .Z(n82417) );
  NOR U102276 ( .A(n82415), .B(n82417), .Z(n88220) );
  IV U102277 ( .A(n82416), .Z(n82418) );
  NOR U102278 ( .A(n82418), .B(n82417), .Z(n88223) );
  NOR U102279 ( .A(n88220), .B(n88223), .Z(n84614) );
  IV U102280 ( .A(n82419), .Z(n82420) );
  NOR U102281 ( .A(n82423), .B(n82420), .Z(n88221) );
  IV U102282 ( .A(n82421), .Z(n82425) );
  NOR U102283 ( .A(n82423), .B(n82422), .Z(n82424) );
  IV U102284 ( .A(n82424), .Z(n82427) );
  NOR U102285 ( .A(n82425), .B(n82427), .Z(n88214) );
  IV U102286 ( .A(n82426), .Z(n82428) );
  NOR U102287 ( .A(n82428), .B(n82427), .Z(n88212) );
  NOR U102288 ( .A(n82430), .B(n82429), .Z(n88218) );
  IV U102289 ( .A(n82431), .Z(n82436) );
  IV U102290 ( .A(n82432), .Z(n82433) );
  NOR U102291 ( .A(n82433), .B(n82444), .Z(n82434) );
  IV U102292 ( .A(n82434), .Z(n82435) );
  NOR U102293 ( .A(n82436), .B(n82435), .Z(n88216) );
  IV U102294 ( .A(n82437), .Z(n82441) );
  NOR U102295 ( .A(n82438), .B(n82444), .Z(n82439) );
  IV U102296 ( .A(n82439), .Z(n82440) );
  NOR U102297 ( .A(n82441), .B(n82440), .Z(n88245) );
  IV U102298 ( .A(n82442), .Z(n82443) );
  NOR U102299 ( .A(n82444), .B(n82443), .Z(n88237) );
  IV U102300 ( .A(n82445), .Z(n82447) );
  NOR U102301 ( .A(n82447), .B(n82446), .Z(n88234) );
  IV U102302 ( .A(n82448), .Z(n90479) );
  IV U102303 ( .A(n82449), .Z(n82450) );
  NOR U102304 ( .A(n82453), .B(n82450), .Z(n84596) );
  IV U102305 ( .A(n84596), .Z(n90483) );
  IV U102306 ( .A(n82451), .Z(n82452) );
  NOR U102307 ( .A(n82453), .B(n82452), .Z(n82454) );
  IV U102308 ( .A(n82454), .Z(n88260) );
  IV U102309 ( .A(n82455), .Z(n82457) );
  NOR U102310 ( .A(n82457), .B(n82456), .Z(n88256) );
  IV U102311 ( .A(n82458), .Z(n82462) );
  IV U102312 ( .A(n82459), .Z(n82470) );
  NOR U102313 ( .A(n82470), .B(n82460), .Z(n82461) );
  IV U102314 ( .A(n82461), .Z(n82464) );
  NOR U102315 ( .A(n82462), .B(n82464), .Z(n90445) );
  IV U102316 ( .A(n82463), .Z(n82465) );
  NOR U102317 ( .A(n82465), .B(n82464), .Z(n90451) );
  IV U102318 ( .A(n82466), .Z(n82468) );
  NOR U102319 ( .A(n82468), .B(n82467), .Z(n90448) );
  NOR U102320 ( .A(n82470), .B(n82469), .Z(n82474) );
  IV U102321 ( .A(n82471), .Z(n82472) );
  NOR U102322 ( .A(n82472), .B(n82477), .Z(n82473) );
  NOR U102323 ( .A(n82474), .B(n82473), .Z(n90465) );
  IV U102324 ( .A(n82475), .Z(n82476) );
  NOR U102325 ( .A(n82477), .B(n82476), .Z(n90461) );
  IV U102326 ( .A(n82481), .Z(n82478) );
  NOR U102327 ( .A(n82479), .B(n82478), .Z(n82486) );
  IV U102328 ( .A(n82480), .Z(n82484) );
  NOR U102329 ( .A(n82482), .B(n82481), .Z(n82483) );
  NOR U102330 ( .A(n82484), .B(n82483), .Z(n82485) );
  NOR U102331 ( .A(n82486), .B(n82485), .Z(n88272) );
  IV U102332 ( .A(n82487), .Z(n82489) );
  NOR U102333 ( .A(n82489), .B(n82488), .Z(n82495) );
  IV U102334 ( .A(n82490), .Z(n82493) );
  IV U102335 ( .A(n82491), .Z(n82492) );
  NOR U102336 ( .A(n82493), .B(n82492), .Z(n82494) );
  NOR U102337 ( .A(n82495), .B(n82494), .Z(n88269) );
  IV U102338 ( .A(n82496), .Z(n82500) );
  IV U102339 ( .A(n82497), .Z(n84560) );
  NOR U102340 ( .A(n82498), .B(n84560), .Z(n82499) );
  IV U102341 ( .A(n82499), .Z(n84563) );
  NOR U102342 ( .A(n82500), .B(n84563), .Z(n90415) );
  IV U102343 ( .A(n90415), .Z(n90412) );
  IV U102344 ( .A(n82501), .Z(n82502) );
  NOR U102345 ( .A(n82502), .B(n84556), .Z(n90359) );
  IV U102346 ( .A(n90359), .Z(n90357) );
  IV U102347 ( .A(n82503), .Z(n82505) );
  NOR U102348 ( .A(n82505), .B(n82504), .Z(n82506) );
  IV U102349 ( .A(n82506), .Z(n88285) );
  IV U102350 ( .A(n82507), .Z(n82508) );
  NOR U102351 ( .A(n84519), .B(n82508), .Z(n88287) );
  IV U102352 ( .A(n82509), .Z(n82510) );
  NOR U102353 ( .A(n82510), .B(n84519), .Z(n84521) );
  IV U102354 ( .A(n82511), .Z(n82512) );
  NOR U102355 ( .A(n82513), .B(n82512), .Z(n82514) );
  IV U102356 ( .A(n82514), .Z(n88277) );
  IV U102357 ( .A(n82515), .Z(n82517) );
  NOR U102358 ( .A(n82517), .B(n82516), .Z(n88308) );
  IV U102359 ( .A(n82518), .Z(n82520) );
  NOR U102360 ( .A(n82520), .B(n82519), .Z(n88279) );
  NOR U102361 ( .A(n88308), .B(n88279), .Z(n84515) );
  IV U102362 ( .A(n82521), .Z(n82522) );
  NOR U102363 ( .A(n82523), .B(n82522), .Z(n82528) );
  IV U102364 ( .A(n82524), .Z(n82525) );
  NOR U102365 ( .A(n82526), .B(n82525), .Z(n82527) );
  NOR U102366 ( .A(n82528), .B(n82527), .Z(n88304) );
  IV U102367 ( .A(n88304), .Z(n88306) );
  NOR U102368 ( .A(n82530), .B(n82529), .Z(n82537) );
  NOR U102369 ( .A(n82532), .B(n82531), .Z(n82535) );
  IV U102370 ( .A(n82533), .Z(n82534) );
  NOR U102371 ( .A(n82535), .B(n82534), .Z(n82536) );
  NOR U102372 ( .A(n82537), .B(n82536), .Z(n88301) );
  IV U102373 ( .A(n82538), .Z(n82540) );
  IV U102374 ( .A(n82539), .Z(n84512) );
  NOR U102375 ( .A(n82540), .B(n84512), .Z(n88339) );
  IV U102376 ( .A(n82541), .Z(n82542) );
  NOR U102377 ( .A(n82542), .B(n82547), .Z(n88348) );
  IV U102378 ( .A(n82543), .Z(n82544) );
  NOR U102379 ( .A(n82544), .B(n84512), .Z(n88342) );
  NOR U102380 ( .A(n88348), .B(n88342), .Z(n84506) );
  IV U102381 ( .A(n82545), .Z(n82546) );
  NOR U102382 ( .A(n82547), .B(n82546), .Z(n84502) );
  IV U102383 ( .A(n82548), .Z(n82550) );
  IV U102384 ( .A(n82549), .Z(n82554) );
  NOR U102385 ( .A(n82550), .B(n82554), .Z(n82551) );
  IV U102386 ( .A(n82551), .Z(n88331) );
  IV U102387 ( .A(n82552), .Z(n82553) );
  NOR U102388 ( .A(n82554), .B(n82553), .Z(n88332) );
  NOR U102389 ( .A(n88333), .B(n88332), .Z(n84500) );
  IV U102390 ( .A(n82555), .Z(n82558) );
  IV U102391 ( .A(n82556), .Z(n82557) );
  NOR U102392 ( .A(n82558), .B(n82557), .Z(n82559) );
  NOR U102393 ( .A(n82560), .B(n82559), .Z(n88317) );
  IV U102394 ( .A(n82561), .Z(n82562) );
  NOR U102395 ( .A(n82562), .B(n82564), .Z(n88360) );
  IV U102396 ( .A(n82563), .Z(n82565) );
  NOR U102397 ( .A(n82565), .B(n82564), .Z(n88357) );
  IV U102398 ( .A(n82566), .Z(n82568) );
  NOR U102399 ( .A(n82568), .B(n82567), .Z(n82573) );
  IV U102400 ( .A(n82569), .Z(n82570) );
  NOR U102401 ( .A(n82571), .B(n82570), .Z(n82572) );
  NOR U102402 ( .A(n82573), .B(n82572), .Z(n88374) );
  IV U102403 ( .A(n82574), .Z(n82576) );
  NOR U102404 ( .A(n82576), .B(n82575), .Z(n88365) );
  IV U102405 ( .A(n82577), .Z(n82578) );
  NOR U102406 ( .A(n82579), .B(n82578), .Z(n82584) );
  IV U102407 ( .A(n82580), .Z(n82582) );
  NOR U102408 ( .A(n82582), .B(n82581), .Z(n82583) );
  NOR U102409 ( .A(n82584), .B(n82583), .Z(n88379) );
  IV U102410 ( .A(n82585), .Z(n82587) );
  NOR U102411 ( .A(n82587), .B(n82586), .Z(n82592) );
  IV U102412 ( .A(n82588), .Z(n82589) );
  NOR U102413 ( .A(n82590), .B(n82589), .Z(n82591) );
  NOR U102414 ( .A(n82592), .B(n82591), .Z(n88389) );
  IV U102415 ( .A(n82593), .Z(n82595) );
  IV U102416 ( .A(n82594), .Z(n84495) );
  NOR U102417 ( .A(n82595), .B(n84495), .Z(n88385) );
  IV U102418 ( .A(n82596), .Z(n82597) );
  NOR U102419 ( .A(n82598), .B(n82597), .Z(n88393) );
  IV U102420 ( .A(n82599), .Z(n82600) );
  NOR U102421 ( .A(n82600), .B(n84477), .Z(n82605) );
  IV U102422 ( .A(n82601), .Z(n82603) );
  NOR U102423 ( .A(n82603), .B(n82602), .Z(n82604) );
  NOR U102424 ( .A(n82605), .B(n82604), .Z(n90326) );
  IV U102425 ( .A(n82606), .Z(n82608) );
  NOR U102426 ( .A(n82608), .B(n82607), .Z(n88399) );
  IV U102427 ( .A(n82609), .Z(n82611) );
  NOR U102428 ( .A(n82611), .B(n82610), .Z(n90329) );
  NOR U102429 ( .A(n88399), .B(n90329), .Z(n84475) );
  IV U102430 ( .A(n82612), .Z(n82618) );
  IV U102431 ( .A(n82613), .Z(n82614) );
  NOR U102432 ( .A(n82615), .B(n82614), .Z(n82616) );
  IV U102433 ( .A(n82616), .Z(n82617) );
  NOR U102434 ( .A(n82618), .B(n82617), .Z(n88396) );
  IV U102435 ( .A(n82619), .Z(n82620) );
  NOR U102436 ( .A(n82621), .B(n82620), .Z(n82622) );
  NOR U102437 ( .A(n82623), .B(n82622), .Z(n82624) );
  NOR U102438 ( .A(n82625), .B(n82624), .Z(n88406) );
  IV U102439 ( .A(n82626), .Z(n82627) );
  NOR U102440 ( .A(n82639), .B(n82627), .Z(n82633) );
  NOR U102441 ( .A(n82629), .B(n82628), .Z(n82631) );
  NOR U102442 ( .A(n82631), .B(n82630), .Z(n82632) );
  NOR U102443 ( .A(n82633), .B(n82632), .Z(n90315) );
  IV U102444 ( .A(n90315), .Z(n90311) );
  IV U102445 ( .A(n82634), .Z(n82635) );
  NOR U102446 ( .A(n82636), .B(n82635), .Z(n82642) );
  NOR U102447 ( .A(n82638), .B(n82637), .Z(n82640) );
  NOR U102448 ( .A(n82640), .B(n82639), .Z(n82641) );
  NOR U102449 ( .A(n82642), .B(n82641), .Z(n90312) );
  IV U102450 ( .A(n82643), .Z(n82649) );
  NOR U102451 ( .A(n84463), .B(n82644), .Z(n82645) );
  IV U102452 ( .A(n82645), .Z(n82646) );
  NOR U102453 ( .A(n82647), .B(n82646), .Z(n82648) );
  IV U102454 ( .A(n82648), .Z(n84468) );
  NOR U102455 ( .A(n82649), .B(n84468), .Z(n84466) );
  IV U102456 ( .A(n84466), .Z(n84461) );
  NOR U102457 ( .A(n82651), .B(n82650), .Z(n82658) );
  NOR U102458 ( .A(n82653), .B(n82652), .Z(n82656) );
  IV U102459 ( .A(n82654), .Z(n82655) );
  NOR U102460 ( .A(n82656), .B(n82655), .Z(n82657) );
  NOR U102461 ( .A(n82658), .B(n82657), .Z(n88420) );
  IV U102462 ( .A(n82659), .Z(n82660) );
  NOR U102463 ( .A(n82664), .B(n82660), .Z(n88416) );
  IV U102464 ( .A(n82661), .Z(n82662) );
  NOR U102465 ( .A(n82663), .B(n82662), .Z(n90264) );
  NOR U102466 ( .A(n82665), .B(n82664), .Z(n90275) );
  NOR U102467 ( .A(n90264), .B(n90275), .Z(n84459) );
  IV U102468 ( .A(n82666), .Z(n82668) );
  NOR U102469 ( .A(n82668), .B(n82667), .Z(n90278) );
  IV U102470 ( .A(n82669), .Z(n82670) );
  NOR U102471 ( .A(n82670), .B(n84449), .Z(n90258) );
  NOR U102472 ( .A(n90278), .B(n90258), .Z(n84447) );
  IV U102473 ( .A(n82671), .Z(n82673) );
  NOR U102474 ( .A(n82673), .B(n82672), .Z(n82674) );
  IV U102475 ( .A(n82674), .Z(n90284) );
  IV U102476 ( .A(n82675), .Z(n82677) );
  NOR U102477 ( .A(n82677), .B(n82676), .Z(n88425) );
  IV U102478 ( .A(n82678), .Z(n82679) );
  NOR U102479 ( .A(n82680), .B(n82679), .Z(n82681) );
  IV U102480 ( .A(n82681), .Z(n84427) );
  IV U102481 ( .A(n82685), .Z(n82683) );
  NOR U102482 ( .A(n82683), .B(n82682), .Z(n82693) );
  NOR U102483 ( .A(n82685), .B(n82684), .Z(n82691) );
  IV U102484 ( .A(n82686), .Z(n82687) );
  NOR U102485 ( .A(n82688), .B(n82687), .Z(n82689) );
  IV U102486 ( .A(n82689), .Z(n82690) );
  NOR U102487 ( .A(n82691), .B(n82690), .Z(n82692) );
  NOR U102488 ( .A(n82693), .B(n82692), .Z(n90245) );
  IV U102489 ( .A(n82694), .Z(n82696) );
  NOR U102490 ( .A(n82696), .B(n82695), .Z(n82700) );
  NOR U102491 ( .A(n82698), .B(n82697), .Z(n82699) );
  NOR U102492 ( .A(n82700), .B(n82699), .Z(n90243) );
  IV U102493 ( .A(n82701), .Z(n82702) );
  NOR U102494 ( .A(n82710), .B(n82702), .Z(n82707) );
  IV U102495 ( .A(n82703), .Z(n82705) );
  NOR U102496 ( .A(n82705), .B(n82704), .Z(n82706) );
  NOR U102497 ( .A(n82707), .B(n82706), .Z(n88464) );
  IV U102498 ( .A(n82708), .Z(n82709) );
  NOR U102499 ( .A(n82710), .B(n82709), .Z(n88439) );
  NOR U102500 ( .A(n82711), .B(n84417), .Z(n88456) );
  IV U102501 ( .A(n82712), .Z(n82713) );
  NOR U102502 ( .A(n82713), .B(n84417), .Z(n82714) );
  IV U102503 ( .A(n82714), .Z(n88455) );
  IV U102504 ( .A(n82715), .Z(n82716) );
  NOR U102505 ( .A(n82717), .B(n82716), .Z(n82721) );
  NOR U102506 ( .A(n82719), .B(n82718), .Z(n82720) );
  NOR U102507 ( .A(n82721), .B(n82720), .Z(n88448) );
  IV U102508 ( .A(n82722), .Z(n82723) );
  NOR U102509 ( .A(n82723), .B(n84410), .Z(n88444) );
  IV U102510 ( .A(n82724), .Z(n82727) );
  NOR U102511 ( .A(n82725), .B(n84386), .Z(n82726) );
  IV U102512 ( .A(n82726), .Z(n82729) );
  NOR U102513 ( .A(n82727), .B(n82729), .Z(n88487) );
  IV U102514 ( .A(n82728), .Z(n82730) );
  NOR U102515 ( .A(n82730), .B(n82729), .Z(n88484) );
  IV U102516 ( .A(n82731), .Z(n82732) );
  NOR U102517 ( .A(n82733), .B(n82732), .Z(n88473) );
  IV U102518 ( .A(n82734), .Z(n82735) );
  NOR U102519 ( .A(n82736), .B(n82735), .Z(n82737) );
  IV U102520 ( .A(n82737), .Z(n84378) );
  IV U102521 ( .A(n82738), .Z(n88469) );
  NOR U102522 ( .A(n88469), .B(n82739), .Z(n84367) );
  IV U102523 ( .A(n82740), .Z(n82741) );
  NOR U102524 ( .A(n82742), .B(n82741), .Z(n88465) );
  NOR U102525 ( .A(n84367), .B(n88465), .Z(n84365) );
  IV U102526 ( .A(n82743), .Z(n82744) );
  NOR U102527 ( .A(n82745), .B(n82744), .Z(n88498) );
  IV U102528 ( .A(n82746), .Z(n82747) );
  NOR U102529 ( .A(n84357), .B(n82747), .Z(n88495) );
  IV U102530 ( .A(n82748), .Z(n82749) );
  NOR U102531 ( .A(n82753), .B(n82749), .Z(n88533) );
  IV U102532 ( .A(n88533), .Z(n88531) );
  IV U102533 ( .A(n82750), .Z(n82751) );
  NOR U102534 ( .A(n82753), .B(n82751), .Z(n82752) );
  IV U102535 ( .A(n82752), .Z(n88515) );
  NOR U102536 ( .A(n82754), .B(n82753), .Z(n88511) );
  IV U102537 ( .A(n82755), .Z(n82758) );
  IV U102538 ( .A(n82756), .Z(n82757) );
  NOR U102539 ( .A(n82758), .B(n82757), .Z(n88521) );
  IV U102540 ( .A(n82759), .Z(n82761) );
  NOR U102541 ( .A(n82761), .B(n82760), .Z(n88518) );
  IV U102542 ( .A(n82762), .Z(n82764) );
  NOR U102543 ( .A(n82764), .B(n82763), .Z(n82769) );
  IV U102544 ( .A(n82765), .Z(n82767) );
  IV U102545 ( .A(n82766), .Z(n84339) );
  NOR U102546 ( .A(n82767), .B(n84339), .Z(n82768) );
  NOR U102547 ( .A(n82769), .B(n82768), .Z(n88539) );
  IV U102548 ( .A(n88539), .Z(n84338) );
  IV U102549 ( .A(n82770), .Z(n82775) );
  IV U102550 ( .A(n82771), .Z(n82772) );
  NOR U102551 ( .A(n82775), .B(n82772), .Z(n90188) );
  IV U102552 ( .A(n82773), .Z(n82774) );
  NOR U102553 ( .A(n82775), .B(n82774), .Z(n90195) );
  IV U102554 ( .A(n82776), .Z(n82777) );
  NOR U102555 ( .A(n82778), .B(n82777), .Z(n90198) );
  NOR U102556 ( .A(n90195), .B(n90198), .Z(n84329) );
  IV U102557 ( .A(n82779), .Z(n82781) );
  NOR U102558 ( .A(n82781), .B(n82780), .Z(n90199) );
  NOR U102559 ( .A(n82782), .B(n82783), .Z(n82789) );
  IV U102560 ( .A(n82783), .Z(n82784) );
  NOR U102561 ( .A(n82785), .B(n82784), .Z(n82786) );
  NOR U102562 ( .A(n82787), .B(n82786), .Z(n82788) );
  NOR U102563 ( .A(n82789), .B(n82788), .Z(n88548) );
  NOR U102564 ( .A(n82791), .B(n82790), .Z(n88545) );
  IV U102565 ( .A(n82792), .Z(n82794) );
  NOR U102566 ( .A(n82794), .B(n82793), .Z(n82799) );
  IV U102567 ( .A(n82795), .Z(n82796) );
  NOR U102568 ( .A(n82797), .B(n82796), .Z(n82798) );
  NOR U102569 ( .A(n82799), .B(n82798), .Z(n88557) );
  IV U102570 ( .A(n82800), .Z(n82801) );
  NOR U102571 ( .A(n82802), .B(n82801), .Z(n82806) );
  IV U102572 ( .A(n82803), .Z(n82804) );
  NOR U102573 ( .A(n82809), .B(n82804), .Z(n82805) );
  NOR U102574 ( .A(n82806), .B(n82805), .Z(n88554) );
  IV U102575 ( .A(n82807), .Z(n82808) );
  NOR U102576 ( .A(n82809), .B(n82808), .Z(n88563) );
  IV U102577 ( .A(n82810), .Z(n82813) );
  IV U102578 ( .A(n82811), .Z(n82812) );
  NOR U102579 ( .A(n82813), .B(n82812), .Z(n88560) );
  IV U102580 ( .A(n82814), .Z(n82816) );
  XOR U102581 ( .A(n82820), .B(n82818), .Z(n82815) );
  NOR U102582 ( .A(n82816), .B(n82815), .Z(n88594) );
  IV U102583 ( .A(n82817), .Z(n82819) );
  NOR U102584 ( .A(n82819), .B(n82818), .Z(n88587) );
  IV U102585 ( .A(n82820), .Z(n82821) );
  NOR U102586 ( .A(n82821), .B(n82827), .Z(n88584) );
  IV U102587 ( .A(n82822), .Z(n82824) );
  NOR U102588 ( .A(n82824), .B(n82823), .Z(n82829) );
  IV U102589 ( .A(n82825), .Z(n82826) );
  NOR U102590 ( .A(n82827), .B(n82826), .Z(n82828) );
  NOR U102591 ( .A(n82829), .B(n82828), .Z(n88571) );
  IV U102592 ( .A(n82830), .Z(n82831) );
  NOR U102593 ( .A(n82832), .B(n82831), .Z(n88578) );
  IV U102594 ( .A(n82833), .Z(n82835) );
  NOR U102595 ( .A(n82835), .B(n82834), .Z(n88573) );
  NOR U102596 ( .A(n88578), .B(n88573), .Z(n84328) );
  IV U102597 ( .A(n82836), .Z(n82837) );
  NOR U102598 ( .A(n82838), .B(n82837), .Z(n88579) );
  IV U102599 ( .A(n82839), .Z(n82840) );
  NOR U102600 ( .A(n82840), .B(n82842), .Z(n88600) );
  IV U102601 ( .A(n82841), .Z(n82843) );
  NOR U102602 ( .A(n82843), .B(n82842), .Z(n88597) );
  NOR U102603 ( .A(n82845), .B(n82844), .Z(n82850) );
  IV U102604 ( .A(n82846), .Z(n82847) );
  NOR U102605 ( .A(n82848), .B(n82847), .Z(n82849) );
  NOR U102606 ( .A(n82850), .B(n82849), .Z(n90156) );
  IV U102607 ( .A(n82851), .Z(n82852) );
  NOR U102608 ( .A(n82853), .B(n82852), .Z(n90142) );
  IV U102609 ( .A(n82854), .Z(n82858) );
  NOR U102610 ( .A(n82856), .B(n82855), .Z(n82857) );
  IV U102611 ( .A(n82857), .Z(n82864) );
  NOR U102612 ( .A(n82858), .B(n82864), .Z(n82862) );
  IV U102613 ( .A(n82859), .Z(n82860) );
  NOR U102614 ( .A(n82860), .B(n84304), .Z(n82861) );
  NOR U102615 ( .A(n82862), .B(n82861), .Z(n90126) );
  IV U102616 ( .A(n82863), .Z(n82865) );
  NOR U102617 ( .A(n82865), .B(n82864), .Z(n90118) );
  IV U102618 ( .A(n82866), .Z(n82869) );
  IV U102619 ( .A(n82867), .Z(n82868) );
  NOR U102620 ( .A(n82869), .B(n82868), .Z(n90115) );
  IV U102621 ( .A(n82870), .Z(n82871) );
  NOR U102622 ( .A(n82872), .B(n82871), .Z(n82873) );
  NOR U102623 ( .A(n82874), .B(n82873), .Z(n90108) );
  NOR U102624 ( .A(n82876), .B(n82875), .Z(n90096) );
  IV U102625 ( .A(n90096), .Z(n90094) );
  IV U102626 ( .A(n82880), .Z(n82877) );
  NOR U102627 ( .A(n82878), .B(n82877), .Z(n82884) );
  IV U102628 ( .A(n82878), .Z(n82879) );
  NOR U102629 ( .A(n82880), .B(n82879), .Z(n82882) );
  NOR U102630 ( .A(n82882), .B(n82881), .Z(n82883) );
  NOR U102631 ( .A(n82884), .B(n82883), .Z(n88636) );
  IV U102632 ( .A(n82885), .Z(n82888) );
  IV U102633 ( .A(n82886), .Z(n82887) );
  NOR U102634 ( .A(n82888), .B(n82887), .Z(n88608) );
  IV U102635 ( .A(n82889), .Z(n82891) );
  NOR U102636 ( .A(n82891), .B(n82890), .Z(n88605) );
  IV U102637 ( .A(n82892), .Z(n82893) );
  NOR U102638 ( .A(n82893), .B(n82895), .Z(n90070) );
  IV U102639 ( .A(n82894), .Z(n82896) );
  NOR U102640 ( .A(n82896), .B(n82895), .Z(n90067) );
  IV U102641 ( .A(n82897), .Z(n82901) );
  NOR U102642 ( .A(n82901), .B(n82898), .Z(n90078) );
  IV U102643 ( .A(n82899), .Z(n82900) );
  NOR U102644 ( .A(n82901), .B(n82900), .Z(n90075) );
  IV U102645 ( .A(n82902), .Z(n82903) );
  NOR U102646 ( .A(n82903), .B(n84279), .Z(n88630) );
  IV U102647 ( .A(n82904), .Z(n82905) );
  NOR U102648 ( .A(n82906), .B(n82905), .Z(n84275) );
  IV U102649 ( .A(n84275), .Z(n84269) );
  IV U102650 ( .A(n82907), .Z(n82908) );
  NOR U102651 ( .A(n82909), .B(n82908), .Z(n88641) );
  IV U102652 ( .A(n82910), .Z(n82911) );
  NOR U102653 ( .A(n82911), .B(n84254), .Z(n82912) );
  IV U102654 ( .A(n82912), .Z(n90058) );
  IV U102655 ( .A(n82913), .Z(n82916) );
  IV U102656 ( .A(n82914), .Z(n82915) );
  NOR U102657 ( .A(n82916), .B(n82915), .Z(n90040) );
  IV U102658 ( .A(n82917), .Z(n82919) );
  NOR U102659 ( .A(n82919), .B(n82918), .Z(n90037) );
  IV U102660 ( .A(n82920), .Z(n88662) );
  IV U102661 ( .A(n82921), .Z(n82922) );
  NOR U102662 ( .A(n82923), .B(n82922), .Z(n88692) );
  NOR U102663 ( .A(n82925), .B(n82924), .Z(n88693) );
  NOR U102664 ( .A(n88692), .B(n88693), .Z(n84241) );
  IV U102665 ( .A(n82926), .Z(n82929) );
  IV U102666 ( .A(n82927), .Z(n82928) );
  NOR U102667 ( .A(n82929), .B(n82928), .Z(n88688) );
  IV U102668 ( .A(n88688), .Z(n88690) );
  IV U102669 ( .A(n82930), .Z(n82932) );
  XOR U102670 ( .A(n84228), .B(n84229), .Z(n82931) );
  NOR U102671 ( .A(n82932), .B(n82931), .Z(n82933) );
  IV U102672 ( .A(n82933), .Z(n88683) );
  IV U102673 ( .A(n82934), .Z(n82937) );
  NOR U102674 ( .A(n82935), .B(n84229), .Z(n82936) );
  IV U102675 ( .A(n82936), .Z(n84226) );
  NOR U102676 ( .A(n82937), .B(n84226), .Z(n88679) );
  IV U102677 ( .A(n82938), .Z(n82939) );
  NOR U102678 ( .A(n82940), .B(n82939), .Z(n88669) );
  IV U102679 ( .A(n82941), .Z(n82943) );
  NOR U102680 ( .A(n82943), .B(n82942), .Z(n88672) );
  NOR U102681 ( .A(n88669), .B(n88672), .Z(n84224) );
  IV U102682 ( .A(n82944), .Z(n84210) );
  IV U102683 ( .A(n84211), .Z(n82945) );
  NOR U102684 ( .A(n84210), .B(n82945), .Z(n90026) );
  IV U102685 ( .A(n82946), .Z(n82947) );
  NOR U102686 ( .A(n82948), .B(n82947), .Z(n90023) );
  NOR U102687 ( .A(n82950), .B(n82949), .Z(n82957) );
  NOR U102688 ( .A(n82952), .B(n82951), .Z(n82955) );
  IV U102689 ( .A(n82953), .Z(n82954) );
  NOR U102690 ( .A(n82955), .B(n82954), .Z(n82956) );
  NOR U102691 ( .A(n82957), .B(n82956), .Z(n90010) );
  IV U102692 ( .A(n82958), .Z(n82960) );
  NOR U102693 ( .A(n82960), .B(n82959), .Z(n90012) );
  NOR U102694 ( .A(n89999), .B(n90012), .Z(n84195) );
  IV U102695 ( .A(n82961), .Z(n82962) );
  NOR U102696 ( .A(n82963), .B(n82962), .Z(n89982) );
  IV U102697 ( .A(n82964), .Z(n82965) );
  NOR U102698 ( .A(n82966), .B(n82965), .Z(n82967) );
  NOR U102699 ( .A(n89990), .B(n82967), .Z(n89988) );
  IV U102700 ( .A(n89988), .Z(n84187) );
  IV U102701 ( .A(n89960), .Z(n89963) );
  IV U102702 ( .A(n82968), .Z(n82969) );
  NOR U102703 ( .A(n82971), .B(n82969), .Z(n88700) );
  NOR U102704 ( .A(n82971), .B(n82970), .Z(n88723) );
  IV U102705 ( .A(n82972), .Z(n82973) );
  NOR U102706 ( .A(n84172), .B(n82973), .Z(n88729) );
  IV U102707 ( .A(n82974), .Z(n82975) );
  NOR U102708 ( .A(n84172), .B(n82975), .Z(n88726) );
  IV U102709 ( .A(n82976), .Z(n82981) );
  IV U102710 ( .A(n82977), .Z(n82978) );
  NOR U102711 ( .A(n82979), .B(n82978), .Z(n82980) );
  IV U102712 ( .A(n82980), .Z(n84174) );
  NOR U102713 ( .A(n82981), .B(n84174), .Z(n88708) );
  IV U102714 ( .A(n82982), .Z(n82985) );
  IV U102715 ( .A(n82983), .Z(n82984) );
  NOR U102716 ( .A(n82985), .B(n82984), .Z(n82986) );
  NOR U102717 ( .A(n82987), .B(n82986), .Z(n88718) );
  IV U102718 ( .A(n82988), .Z(n82989) );
  NOR U102719 ( .A(n84166), .B(n82989), .Z(n82990) );
  IV U102720 ( .A(n82990), .Z(n88740) );
  IV U102721 ( .A(n82991), .Z(n82992) );
  NOR U102722 ( .A(n82992), .B(n82994), .Z(n88741) );
  IV U102723 ( .A(n82993), .Z(n82995) );
  NOR U102724 ( .A(n82995), .B(n82994), .Z(n89940) );
  IV U102725 ( .A(n82996), .Z(n82998) );
  NOR U102726 ( .A(n82998), .B(n82997), .Z(n84153) );
  IV U102727 ( .A(n84153), .Z(n89935) );
  IV U102728 ( .A(n82999), .Z(n83000) );
  NOR U102729 ( .A(n83000), .B(n83007), .Z(n83001) );
  IV U102730 ( .A(n83001), .Z(n89928) );
  IV U102731 ( .A(n83002), .Z(n83004) );
  NOR U102732 ( .A(n83004), .B(n83003), .Z(n83009) );
  IV U102733 ( .A(n83005), .Z(n83006) );
  NOR U102734 ( .A(n83007), .B(n83006), .Z(n83008) );
  NOR U102735 ( .A(n83009), .B(n83008), .Z(n89927) );
  IV U102736 ( .A(n83010), .Z(n83012) );
  NOR U102737 ( .A(n83012), .B(n83011), .Z(n83013) );
  NOR U102738 ( .A(n83014), .B(n83013), .Z(n88752) );
  IV U102739 ( .A(n83015), .Z(n83016) );
  NOR U102740 ( .A(n83016), .B(n84146), .Z(n83024) );
  IV U102741 ( .A(n83017), .Z(n83018) );
  NOR U102742 ( .A(n83018), .B(n83036), .Z(n83019) );
  IV U102743 ( .A(n83019), .Z(n83022) );
  IV U102744 ( .A(n83020), .Z(n83021) );
  NOR U102745 ( .A(n83022), .B(n83021), .Z(n83023) );
  NOR U102746 ( .A(n83024), .B(n83023), .Z(n88761) );
  IV U102747 ( .A(n83025), .Z(n83028) );
  NOR U102748 ( .A(n83026), .B(n83036), .Z(n83027) );
  IV U102749 ( .A(n83027), .Z(n83030) );
  NOR U102750 ( .A(n83028), .B(n83030), .Z(n88757) );
  IV U102751 ( .A(n83029), .Z(n83031) );
  NOR U102752 ( .A(n83031), .B(n83030), .Z(n83042) );
  IV U102753 ( .A(n83032), .Z(n83034) );
  XOR U102754 ( .A(n83035), .B(n83036), .Z(n83033) );
  NOR U102755 ( .A(n83034), .B(n83033), .Z(n83039) );
  IV U102756 ( .A(n83035), .Z(n83037) );
  NOR U102757 ( .A(n83037), .B(n83036), .Z(n83038) );
  NOR U102758 ( .A(n83039), .B(n83038), .Z(n83040) );
  IV U102759 ( .A(n83040), .Z(n83041) );
  NOR U102760 ( .A(n83042), .B(n83041), .Z(n88755) );
  IV U102761 ( .A(n83043), .Z(n83044) );
  NOR U102762 ( .A(n83045), .B(n83044), .Z(n83050) );
  IV U102763 ( .A(n83046), .Z(n83048) );
  NOR U102764 ( .A(n83048), .B(n83047), .Z(n83049) );
  NOR U102765 ( .A(n83050), .B(n83049), .Z(n89911) );
  IV U102766 ( .A(n89911), .Z(n83054) );
  IV U102767 ( .A(n83051), .Z(n83052) );
  NOR U102768 ( .A(n83053), .B(n83052), .Z(n89903) );
  NOR U102769 ( .A(n83054), .B(n89903), .Z(n84143) );
  IV U102770 ( .A(n83055), .Z(n83056) );
  NOR U102771 ( .A(n83058), .B(n83056), .Z(n84141) );
  IV U102772 ( .A(n83057), .Z(n83059) );
  NOR U102773 ( .A(n83059), .B(n83058), .Z(n83064) );
  IV U102774 ( .A(n83060), .Z(n83062) );
  IV U102775 ( .A(n83061), .Z(n83068) );
  NOR U102776 ( .A(n83062), .B(n83068), .Z(n83063) );
  NOR U102777 ( .A(n83064), .B(n83063), .Z(n89902) );
  IV U102778 ( .A(n83065), .Z(n83066) );
  NOR U102779 ( .A(n83066), .B(n83074), .Z(n89889) );
  IV U102780 ( .A(n83067), .Z(n83069) );
  NOR U102781 ( .A(n83069), .B(n83068), .Z(n88764) );
  NOR U102782 ( .A(n89889), .B(n88764), .Z(n84138) );
  IV U102783 ( .A(n83070), .Z(n83072) );
  NOR U102784 ( .A(n83072), .B(n83071), .Z(n89894) );
  IV U102785 ( .A(n83073), .Z(n83075) );
  NOR U102786 ( .A(n83075), .B(n83074), .Z(n88766) );
  NOR U102787 ( .A(n89894), .B(n88766), .Z(n84137) );
  IV U102788 ( .A(n83076), .Z(n83077) );
  NOR U102789 ( .A(n83078), .B(n83077), .Z(n84131) );
  IV U102790 ( .A(n83079), .Z(n83081) );
  IV U102791 ( .A(n83080), .Z(n83083) );
  NOR U102792 ( .A(n83081), .B(n83083), .Z(n84128) );
  IV U102793 ( .A(n83082), .Z(n83084) );
  NOR U102794 ( .A(n83084), .B(n83083), .Z(n89876) );
  IV U102795 ( .A(n83085), .Z(n83087) );
  XOR U102796 ( .A(n83088), .B(n84114), .Z(n83086) );
  NOR U102797 ( .A(n83087), .B(n83086), .Z(n89879) );
  IV U102798 ( .A(n83088), .Z(n83089) );
  NOR U102799 ( .A(n83089), .B(n84114), .Z(n84116) );
  IV U102800 ( .A(n83090), .Z(n83091) );
  NOR U102801 ( .A(n83092), .B(n83091), .Z(n83093) );
  IV U102802 ( .A(n83093), .Z(n89849) );
  IV U102803 ( .A(n83094), .Z(n83096) );
  IV U102804 ( .A(n83095), .Z(n84110) );
  NOR U102805 ( .A(n83096), .B(n84110), .Z(n89855) );
  IV U102806 ( .A(n83097), .Z(n83098) );
  NOR U102807 ( .A(n83101), .B(n83098), .Z(n89852) );
  IV U102808 ( .A(n83099), .Z(n83100) );
  NOR U102809 ( .A(n83101), .B(n83100), .Z(n89869) );
  IV U102810 ( .A(n83102), .Z(n83104) );
  IV U102811 ( .A(n83103), .Z(n84101) );
  NOR U102812 ( .A(n83104), .B(n84101), .Z(n88775) );
  IV U102813 ( .A(n83105), .Z(n83106) );
  NOR U102814 ( .A(n83109), .B(n83106), .Z(n89813) );
  IV U102815 ( .A(n83107), .Z(n83108) );
  NOR U102816 ( .A(n83109), .B(n83108), .Z(n89810) );
  IV U102817 ( .A(n83110), .Z(n83111) );
  NOR U102818 ( .A(n83111), .B(n84085), .Z(n83112) );
  IV U102819 ( .A(n83112), .Z(n89835) );
  IV U102820 ( .A(n84086), .Z(n83113) );
  NOR U102821 ( .A(n83113), .B(n84085), .Z(n89831) );
  IV U102822 ( .A(n83114), .Z(n83117) );
  IV U102823 ( .A(n83115), .Z(n83116) );
  NOR U102824 ( .A(n83117), .B(n83116), .Z(n83118) );
  IV U102825 ( .A(n83118), .Z(n88791) );
  IV U102826 ( .A(n83119), .Z(n83120) );
  NOR U102827 ( .A(n83123), .B(n83120), .Z(n88795) );
  IV U102828 ( .A(n83121), .Z(n83122) );
  NOR U102829 ( .A(n83123), .B(n83122), .Z(n83128) );
  IV U102830 ( .A(n83124), .Z(n83125) );
  NOR U102831 ( .A(n83126), .B(n83125), .Z(n83127) );
  NOR U102832 ( .A(n83128), .B(n83127), .Z(n88781) );
  NOR U102833 ( .A(n83130), .B(n83129), .Z(n84041) );
  IV U102834 ( .A(n83131), .Z(n83132) );
  NOR U102835 ( .A(n83133), .B(n83132), .Z(n88808) );
  IV U102836 ( .A(n83134), .Z(n83136) );
  IV U102837 ( .A(n83135), .Z(n84031) );
  NOR U102838 ( .A(n83136), .B(n84031), .Z(n88805) );
  IV U102839 ( .A(n83137), .Z(n83138) );
  NOR U102840 ( .A(n84031), .B(n83138), .Z(n88816) );
  IV U102841 ( .A(n83139), .Z(n83140) );
  NOR U102842 ( .A(n83141), .B(n83140), .Z(n83142) );
  IV U102843 ( .A(n83142), .Z(n88837) );
  IV U102844 ( .A(n83143), .Z(n83144) );
  NOR U102845 ( .A(n83144), .B(n83993), .Z(n88855) );
  IV U102846 ( .A(n83145), .Z(n83146) );
  NOR U102847 ( .A(n83147), .B(n83146), .Z(n88861) );
  IV U102848 ( .A(n83148), .Z(n83150) );
  NOR U102849 ( .A(n83150), .B(n83149), .Z(n88876) );
  NOR U102850 ( .A(n88861), .B(n88876), .Z(n83974) );
  IV U102851 ( .A(n83151), .Z(n83153) );
  NOR U102852 ( .A(n83153), .B(n83152), .Z(n88866) );
  NOR U102853 ( .A(n83155), .B(n83154), .Z(n83161) );
  NOR U102854 ( .A(n83157), .B(n83156), .Z(n83158) );
  NOR U102855 ( .A(n83159), .B(n83158), .Z(n83160) );
  NOR U102856 ( .A(n83161), .B(n83160), .Z(n88863) );
  IV U102857 ( .A(n83162), .Z(n83163) );
  NOR U102858 ( .A(n83164), .B(n83163), .Z(n88919) );
  IV U102859 ( .A(n83165), .Z(n83170) );
  IV U102860 ( .A(n83166), .Z(n83167) );
  NOR U102861 ( .A(n83170), .B(n83167), .Z(n88916) );
  IV U102862 ( .A(n83168), .Z(n83169) );
  NOR U102863 ( .A(n83170), .B(n83169), .Z(n88927) );
  IV U102864 ( .A(n83171), .Z(n83172) );
  NOR U102865 ( .A(n83177), .B(n83172), .Z(n88924) );
  IV U102866 ( .A(n83173), .Z(n83174) );
  NOR U102867 ( .A(n83177), .B(n83174), .Z(n88889) );
  IV U102868 ( .A(n83175), .Z(n83176) );
  NOR U102869 ( .A(n83177), .B(n83176), .Z(n88909) );
  IV U102870 ( .A(n83178), .Z(n83180) );
  IV U102871 ( .A(n83179), .Z(n83965) );
  NOR U102872 ( .A(n83180), .B(n83965), .Z(n88906) );
  IV U102873 ( .A(n83181), .Z(n83183) );
  NOR U102874 ( .A(n83183), .B(n83182), .Z(n88893) );
  IV U102875 ( .A(n83184), .Z(n83185) );
  NOR U102876 ( .A(n83961), .B(n83185), .Z(n88939) );
  IV U102877 ( .A(n83186), .Z(n83187) );
  NOR U102878 ( .A(n83188), .B(n83187), .Z(n83189) );
  NOR U102879 ( .A(n83190), .B(n83189), .Z(n89765) );
  IV U102880 ( .A(n83193), .Z(n83191) );
  NOR U102881 ( .A(n83192), .B(n83191), .Z(n83198) );
  IV U102882 ( .A(n83192), .Z(n83194) );
  NOR U102883 ( .A(n83194), .B(n83193), .Z(n83195) );
  NOR U102884 ( .A(n83196), .B(n83195), .Z(n83197) );
  NOR U102885 ( .A(n83198), .B(n83197), .Z(n89753) );
  IV U102886 ( .A(n83199), .Z(n83201) );
  NOR U102887 ( .A(n83201), .B(n83200), .Z(n89742) );
  IV U102888 ( .A(n83202), .Z(n83203) );
  NOR U102889 ( .A(n83204), .B(n83203), .Z(n88950) );
  NOR U102890 ( .A(n89742), .B(n88950), .Z(n83943) );
  IV U102891 ( .A(n83205), .Z(n83206) );
  NOR U102892 ( .A(n83206), .B(n83939), .Z(n89735) );
  IV U102893 ( .A(n83207), .Z(n83211) );
  NOR U102894 ( .A(n83209), .B(n83208), .Z(n83210) );
  IV U102895 ( .A(n83210), .Z(n83213) );
  NOR U102896 ( .A(n83211), .B(n83213), .Z(n89713) );
  IV U102897 ( .A(n83212), .Z(n83214) );
  NOR U102898 ( .A(n83214), .B(n83213), .Z(n89722) );
  IV U102899 ( .A(n83215), .Z(n83218) );
  NOR U102900 ( .A(n83216), .B(n83226), .Z(n83217) );
  IV U102901 ( .A(n83217), .Z(n83220) );
  NOR U102902 ( .A(n83218), .B(n83220), .Z(n89719) );
  IV U102903 ( .A(n83219), .Z(n83221) );
  NOR U102904 ( .A(n83221), .B(n83220), .Z(n88956) );
  IV U102905 ( .A(n83222), .Z(n83223) );
  NOR U102906 ( .A(n83224), .B(n83223), .Z(n89689) );
  IV U102907 ( .A(n83225), .Z(n83227) );
  NOR U102908 ( .A(n83227), .B(n83226), .Z(n88953) );
  NOR U102909 ( .A(n89689), .B(n88953), .Z(n83934) );
  IV U102910 ( .A(n83228), .Z(n83230) );
  IV U102911 ( .A(n83229), .Z(n83924) );
  NOR U102912 ( .A(n83230), .B(n83924), .Z(n89702) );
  IV U102913 ( .A(n83231), .Z(n83232) );
  NOR U102914 ( .A(n83233), .B(n83232), .Z(n88964) );
  IV U102915 ( .A(n83234), .Z(n83238) );
  NOR U102916 ( .A(n83236), .B(n83235), .Z(n83237) );
  IV U102917 ( .A(n83237), .Z(n83240) );
  NOR U102918 ( .A(n83238), .B(n83240), .Z(n89678) );
  IV U102919 ( .A(n83239), .Z(n83241) );
  NOR U102920 ( .A(n83241), .B(n83240), .Z(n89675) );
  NOR U102921 ( .A(n83243), .B(n83242), .Z(n89650) );
  IV U102922 ( .A(n83244), .Z(n83245) );
  NOR U102923 ( .A(n83246), .B(n83245), .Z(n89646) );
  IV U102924 ( .A(n83247), .Z(n83251) );
  NOR U102925 ( .A(n83249), .B(n83248), .Z(n83250) );
  IV U102926 ( .A(n83250), .Z(n83253) );
  NOR U102927 ( .A(n83251), .B(n83253), .Z(n89656) );
  IV U102928 ( .A(n83252), .Z(n83254) );
  NOR U102929 ( .A(n83254), .B(n83253), .Z(n89653) );
  IV U102930 ( .A(n83255), .Z(n83256) );
  NOR U102931 ( .A(n83256), .B(n83898), .Z(n89638) );
  IV U102932 ( .A(n83257), .Z(n83258) );
  NOR U102933 ( .A(n83258), .B(n83892), .Z(n88978) );
  IV U102934 ( .A(n83259), .Z(n83260) );
  NOR U102935 ( .A(n83260), .B(n83892), .Z(n88973) );
  IV U102936 ( .A(n83261), .Z(n83263) );
  IV U102937 ( .A(n83262), .Z(n83265) );
  NOR U102938 ( .A(n83263), .B(n83265), .Z(n89621) );
  NOR U102939 ( .A(n83265), .B(n83264), .Z(n89605) );
  IV U102940 ( .A(n83266), .Z(n83271) );
  IV U102941 ( .A(n83267), .Z(n83871) );
  NOR U102942 ( .A(n83871), .B(n83268), .Z(n83269) );
  IV U102943 ( .A(n83269), .Z(n83270) );
  NOR U102944 ( .A(n83271), .B(n83270), .Z(n83883) );
  IV U102945 ( .A(n83272), .Z(n83274) );
  NOR U102946 ( .A(n83274), .B(n83273), .Z(n83868) );
  IV U102947 ( .A(n83868), .Z(n83865) );
  IV U102948 ( .A(n83278), .Z(n83276) );
  NOR U102949 ( .A(n83276), .B(n83275), .Z(n83283) );
  NOR U102950 ( .A(n83278), .B(n83277), .Z(n83281) );
  IV U102951 ( .A(n83279), .Z(n83280) );
  NOR U102952 ( .A(n83281), .B(n83280), .Z(n83282) );
  NOR U102953 ( .A(n83283), .B(n83282), .Z(n89015) );
  IV U102954 ( .A(n83284), .Z(n83285) );
  NOR U102955 ( .A(n83286), .B(n83285), .Z(n89028) );
  IV U102956 ( .A(n83287), .Z(n83289) );
  NOR U102957 ( .A(n83289), .B(n83288), .Z(n88999) );
  NOR U102958 ( .A(n89028), .B(n88999), .Z(n83855) );
  IV U102959 ( .A(n83290), .Z(n83292) );
  IV U102960 ( .A(n83291), .Z(n83294) );
  NOR U102961 ( .A(n83292), .B(n83294), .Z(n89027) );
  IV U102962 ( .A(n83293), .Z(n83295) );
  NOR U102963 ( .A(n83295), .B(n83294), .Z(n88985) );
  IV U102964 ( .A(n83296), .Z(n83297) );
  NOR U102965 ( .A(n83297), .B(n83300), .Z(n88982) );
  IV U102966 ( .A(n83298), .Z(n83299) );
  NOR U102967 ( .A(n83300), .B(n83299), .Z(n83301) );
  IV U102968 ( .A(n83301), .Z(n88994) );
  IV U102969 ( .A(n83302), .Z(n83303) );
  NOR U102970 ( .A(n83303), .B(n83840), .Z(n89038) );
  IV U102971 ( .A(n83304), .Z(n83305) );
  NOR U102972 ( .A(n83305), .B(n83840), .Z(n89042) );
  IV U102973 ( .A(n83309), .Z(n83307) );
  NOR U102974 ( .A(n83307), .B(n83306), .Z(n83316) );
  NOR U102975 ( .A(n83309), .B(n83308), .Z(n83314) );
  IV U102976 ( .A(n83310), .Z(n83311) );
  NOR U102977 ( .A(n83311), .B(n83841), .Z(n83312) );
  IV U102978 ( .A(n83312), .Z(n83313) );
  NOR U102979 ( .A(n83314), .B(n83313), .Z(n83315) );
  NOR U102980 ( .A(n83316), .B(n83315), .Z(n89035) );
  IV U102981 ( .A(n83317), .Z(n83318) );
  NOR U102982 ( .A(n83318), .B(n83825), .Z(n89047) );
  IV U102983 ( .A(n83319), .Z(n83320) );
  NOR U102984 ( .A(n83320), .B(n83821), .Z(n83321) );
  IV U102985 ( .A(n83321), .Z(n89557) );
  NOR U102986 ( .A(n83324), .B(n83322), .Z(n89553) );
  NOR U102987 ( .A(n83324), .B(n83323), .Z(n89563) );
  NOR U102988 ( .A(n83326), .B(n83325), .Z(n83332) );
  IV U102989 ( .A(n83326), .Z(n83328) );
  NOR U102990 ( .A(n83328), .B(n83327), .Z(n83329) );
  NOR U102991 ( .A(n83330), .B(n83329), .Z(n83331) );
  NOR U102992 ( .A(n83332), .B(n83331), .Z(n89560) );
  IV U102993 ( .A(n83333), .Z(n83335) );
  NOR U102994 ( .A(n83335), .B(n83334), .Z(n89058) );
  NOR U102995 ( .A(n83337), .B(n83336), .Z(n89055) );
  IV U102996 ( .A(n83338), .Z(n83340) );
  NOR U102997 ( .A(n83340), .B(n83339), .Z(n89536) );
  IV U102998 ( .A(n83341), .Z(n83343) );
  IV U102999 ( .A(n83342), .Z(n83810) );
  NOR U103000 ( .A(n83343), .B(n83810), .Z(n89066) );
  IV U103001 ( .A(n83344), .Z(n83345) );
  NOR U103002 ( .A(n83805), .B(n83345), .Z(n83346) );
  IV U103003 ( .A(n83346), .Z(n89065) );
  IV U103004 ( .A(n83347), .Z(n83348) );
  NOR U103005 ( .A(n83353), .B(n83348), .Z(n83802) );
  IV U103006 ( .A(n83802), .Z(n89074) );
  IV U103007 ( .A(n83349), .Z(n83350) );
  NOR U103008 ( .A(n83350), .B(n83361), .Z(n83351) );
  IV U103009 ( .A(n83351), .Z(n89087) );
  IV U103010 ( .A(n83352), .Z(n83354) );
  NOR U103011 ( .A(n83354), .B(n83353), .Z(n83355) );
  IV U103012 ( .A(n83355), .Z(n89090) );
  IV U103013 ( .A(n83356), .Z(n83358) );
  NOR U103014 ( .A(n83358), .B(n83357), .Z(n83363) );
  IV U103015 ( .A(n83359), .Z(n83360) );
  NOR U103016 ( .A(n83361), .B(n83360), .Z(n83362) );
  NOR U103017 ( .A(n83363), .B(n83362), .Z(n89092) );
  IV U103018 ( .A(n83364), .Z(n83365) );
  NOR U103019 ( .A(n89103), .B(n83365), .Z(n83800) );
  IV U103020 ( .A(n83366), .Z(n83367) );
  NOR U103021 ( .A(n83368), .B(n83367), .Z(n83373) );
  IV U103022 ( .A(n83369), .Z(n83370) );
  NOR U103023 ( .A(n83371), .B(n83370), .Z(n83372) );
  NOR U103024 ( .A(n83373), .B(n83372), .Z(n89473) );
  IV U103025 ( .A(n83374), .Z(n83375) );
  NOR U103026 ( .A(n83376), .B(n83375), .Z(n89469) );
  XOR U103027 ( .A(n83776), .B(n83378), .Z(n83377) );
  NOR U103028 ( .A(n83379), .B(n83377), .Z(n83384) );
  IV U103029 ( .A(n83378), .Z(n83778) );
  IV U103030 ( .A(n83379), .Z(n83380) );
  NOR U103031 ( .A(n83778), .B(n83380), .Z(n83382) );
  NOR U103032 ( .A(n83382), .B(n83381), .Z(n83383) );
  NOR U103033 ( .A(n83384), .B(n83383), .Z(n89122) );
  IV U103034 ( .A(n83385), .Z(n83389) );
  NOR U103035 ( .A(n83387), .B(n83386), .Z(n83388) );
  IV U103036 ( .A(n83388), .Z(n83391) );
  NOR U103037 ( .A(n83389), .B(n83391), .Z(n83775) );
  IV U103038 ( .A(n83775), .Z(n89117) );
  IV U103039 ( .A(n83390), .Z(n83392) );
  NOR U103040 ( .A(n83392), .B(n83391), .Z(n83393) );
  IV U103041 ( .A(n83393), .Z(n89480) );
  IV U103042 ( .A(n83394), .Z(n83397) );
  NOR U103043 ( .A(n83395), .B(n83399), .Z(n83396) );
  IV U103044 ( .A(n83396), .Z(n83402) );
  NOR U103045 ( .A(n83397), .B(n83402), .Z(n89476) );
  IV U103046 ( .A(n83398), .Z(n83400) );
  NOR U103047 ( .A(n83400), .B(n83399), .Z(n89456) );
  IV U103048 ( .A(n83401), .Z(n83403) );
  NOR U103049 ( .A(n83403), .B(n83402), .Z(n89127) );
  NOR U103050 ( .A(n89456), .B(n89127), .Z(n83404) );
  IV U103051 ( .A(n83404), .Z(n83773) );
  IV U103052 ( .A(n83405), .Z(n83406) );
  NOR U103053 ( .A(n83407), .B(n83406), .Z(n89457) );
  IV U103054 ( .A(n83408), .Z(n83409) );
  NOR U103055 ( .A(n83410), .B(n83409), .Z(n89459) );
  NOR U103056 ( .A(n89457), .B(n89459), .Z(n83772) );
  IV U103057 ( .A(n83411), .Z(n83412) );
  NOR U103058 ( .A(n83768), .B(n83412), .Z(n89453) );
  IV U103059 ( .A(n83413), .Z(n83415) );
  NOR U103060 ( .A(n83415), .B(n83414), .Z(n83420) );
  IV U103061 ( .A(n83416), .Z(n83418) );
  NOR U103062 ( .A(n83418), .B(n83417), .Z(n83419) );
  NOR U103063 ( .A(n83420), .B(n83419), .Z(n89137) );
  IV U103064 ( .A(n83421), .Z(n83426) );
  IV U103065 ( .A(n83422), .Z(n83423) );
  NOR U103066 ( .A(n83426), .B(n83423), .Z(n89130) );
  IV U103067 ( .A(n83424), .Z(n83425) );
  NOR U103068 ( .A(n83426), .B(n83425), .Z(n89143) );
  IV U103069 ( .A(n83427), .Z(n83430) );
  NOR U103070 ( .A(n83428), .B(n83749), .Z(n83429) );
  IV U103071 ( .A(n83429), .Z(n83432) );
  NOR U103072 ( .A(n83430), .B(n83432), .Z(n89149) );
  IV U103073 ( .A(n83431), .Z(n83433) );
  NOR U103074 ( .A(n83433), .B(n83432), .Z(n89146) );
  IV U103075 ( .A(n83434), .Z(n83435) );
  NOR U103076 ( .A(n83436), .B(n83435), .Z(n83437) );
  IV U103077 ( .A(n83437), .Z(n83758) );
  IV U103078 ( .A(n83438), .Z(n83440) );
  NOR U103079 ( .A(n83440), .B(n83439), .Z(n89157) );
  IV U103080 ( .A(n83441), .Z(n83442) );
  NOR U103081 ( .A(n83443), .B(n83442), .Z(n89154) );
  IV U103082 ( .A(n83444), .Z(n83445) );
  NOR U103083 ( .A(n83744), .B(n83445), .Z(n89165) );
  IV U103084 ( .A(n83450), .Z(n83449) );
  IV U103085 ( .A(n83446), .Z(n83447) );
  NOR U103086 ( .A(n83449), .B(n83447), .Z(n83730) );
  NOR U103087 ( .A(n83449), .B(n83448), .Z(n83456) );
  NOR U103088 ( .A(n83451), .B(n83450), .Z(n83454) );
  IV U103089 ( .A(n83452), .Z(n83453) );
  NOR U103090 ( .A(n83454), .B(n83453), .Z(n83455) );
  NOR U103091 ( .A(n83456), .B(n83455), .Z(n89174) );
  IV U103092 ( .A(n83457), .Z(n83460) );
  NOR U103093 ( .A(n83458), .B(n83712), .Z(n83459) );
  IV U103094 ( .A(n83459), .Z(n83462) );
  NOR U103095 ( .A(n83460), .B(n83462), .Z(n83720) );
  IV U103096 ( .A(n83461), .Z(n83463) );
  NOR U103097 ( .A(n83463), .B(n83462), .Z(n83717) );
  IV U103098 ( .A(n83464), .Z(n83466) );
  NOR U103099 ( .A(n83466), .B(n83465), .Z(n89403) );
  IV U103100 ( .A(n83467), .Z(n83469) );
  NOR U103101 ( .A(n83469), .B(n83468), .Z(n89415) );
  NOR U103102 ( .A(n89403), .B(n89415), .Z(n83710) );
  IV U103103 ( .A(n83475), .Z(n83472) );
  IV U103104 ( .A(n83470), .Z(n83471) );
  NOR U103105 ( .A(n83472), .B(n83471), .Z(n89398) );
  IV U103106 ( .A(n89398), .Z(n89401) );
  IV U103107 ( .A(n83476), .Z(n83473) );
  NOR U103108 ( .A(n83473), .B(n83472), .Z(n83480) );
  IV U103109 ( .A(n83474), .Z(n83478) );
  NOR U103110 ( .A(n83476), .B(n83475), .Z(n83477) );
  NOR U103111 ( .A(n83478), .B(n83477), .Z(n83479) );
  NOR U103112 ( .A(n83480), .B(n83479), .Z(n89423) );
  NOR U103113 ( .A(n83482), .B(n83481), .Z(n89196) );
  IV U103114 ( .A(n83483), .Z(n83484) );
  NOR U103115 ( .A(n83484), .B(n83486), .Z(n89180) );
  NOR U103116 ( .A(n83486), .B(n83485), .Z(n89185) );
  IV U103117 ( .A(n83487), .Z(n83489) );
  NOR U103118 ( .A(n83489), .B(n83488), .Z(n89204) );
  IV U103119 ( .A(n83490), .Z(n83491) );
  NOR U103120 ( .A(n83492), .B(n83491), .Z(n89188) );
  NOR U103121 ( .A(n89204), .B(n89188), .Z(n83689) );
  IV U103122 ( .A(n83493), .Z(n83494) );
  NOR U103123 ( .A(n83497), .B(n83494), .Z(n89206) );
  IV U103124 ( .A(n89206), .Z(n89202) );
  IV U103125 ( .A(n83495), .Z(n83496) );
  NOR U103126 ( .A(n83497), .B(n83496), .Z(n83498) );
  IV U103127 ( .A(n83498), .Z(n89373) );
  IV U103128 ( .A(n83499), .Z(n83500) );
  XOR U103129 ( .A(n83509), .B(n83511), .Z(n83506) );
  NOR U103130 ( .A(n83500), .B(n83506), .Z(n83501) );
  IV U103131 ( .A(n83501), .Z(n89370) );
  IV U103132 ( .A(n83502), .Z(n83503) );
  NOR U103133 ( .A(n83503), .B(n83511), .Z(n83508) );
  IV U103134 ( .A(n83504), .Z(n83505) );
  NOR U103135 ( .A(n83506), .B(n83505), .Z(n83507) );
  NOR U103136 ( .A(n83508), .B(n83507), .Z(n89380) );
  IV U103137 ( .A(n83509), .Z(n83510) );
  NOR U103138 ( .A(n83511), .B(n83510), .Z(n83512) );
  IV U103139 ( .A(n83512), .Z(n89377) );
  IV U103140 ( .A(n83513), .Z(n83514) );
  NOR U103141 ( .A(n83519), .B(n83514), .Z(n89212) );
  IV U103142 ( .A(n83515), .Z(n83516) );
  NOR U103143 ( .A(n83517), .B(n83516), .Z(n89219) );
  NOR U103144 ( .A(n89212), .B(n89219), .Z(n83688) );
  IV U103145 ( .A(n83518), .Z(n83520) );
  NOR U103146 ( .A(n83520), .B(n83519), .Z(n89214) );
  IV U103147 ( .A(n89214), .Z(n89210) );
  IV U103148 ( .A(n83521), .Z(n83523) );
  NOR U103149 ( .A(n83523), .B(n83522), .Z(n89227) );
  IV U103150 ( .A(n83524), .Z(n83525) );
  NOR U103151 ( .A(n83526), .B(n83525), .Z(n89224) );
  IV U103152 ( .A(n83527), .Z(n83529) );
  IV U103153 ( .A(n83528), .Z(n83675) );
  NOR U103154 ( .A(n83529), .B(n83675), .Z(n89257) );
  IV U103155 ( .A(n83530), .Z(n83532) );
  NOR U103156 ( .A(n83532), .B(n83531), .Z(n89264) );
  NOR U103157 ( .A(n83534), .B(n83533), .Z(n83671) );
  IV U103158 ( .A(n83671), .Z(n83666) );
  IV U103159 ( .A(n83535), .Z(n83536) );
  NOR U103160 ( .A(n83537), .B(n83536), .Z(n83542) );
  IV U103161 ( .A(n83538), .Z(n83539) );
  NOR U103162 ( .A(n83540), .B(n83539), .Z(n83541) );
  NOR U103163 ( .A(n83542), .B(n83541), .Z(n89239) );
  IV U103164 ( .A(n83543), .Z(n83545) );
  XOR U103165 ( .A(n83546), .B(n83548), .Z(n83544) );
  NOR U103166 ( .A(n83545), .B(n83544), .Z(n83654) );
  IV U103167 ( .A(n83654), .Z(n89276) );
  IV U103168 ( .A(n83549), .Z(n83550) );
  NOR U103169 ( .A(n83550), .B(n83553), .Z(n89327) );
  IV U103170 ( .A(n83551), .Z(n83552) );
  NOR U103171 ( .A(n83553), .B(n83552), .Z(n89350) );
  NOR U103172 ( .A(n89327), .B(n89350), .Z(n83644) );
  IV U103173 ( .A(n83554), .Z(n83555) );
  NOR U103174 ( .A(n83555), .B(n83639), .Z(n83556) );
  IV U103175 ( .A(n83556), .Z(n83557) );
  NOR U103176 ( .A(n83558), .B(n83557), .Z(n89346) );
  IV U103177 ( .A(n83559), .Z(n83563) );
  IV U103178 ( .A(n83560), .Z(n83629) );
  NOR U103179 ( .A(n83629), .B(n83561), .Z(n83562) );
  IV U103180 ( .A(n83562), .Z(n83624) );
  NOR U103181 ( .A(n83563), .B(n83624), .Z(n89319) );
  IV U103182 ( .A(n83564), .Z(n83565) );
  NOR U103183 ( .A(n83565), .B(n83568), .Z(n83566) );
  IV U103184 ( .A(n83566), .Z(n89332) );
  IV U103185 ( .A(n83567), .Z(n83569) );
  NOR U103186 ( .A(n83569), .B(n83568), .Z(n89304) );
  IV U103187 ( .A(n83570), .Z(n83572) );
  IV U103188 ( .A(n83571), .Z(n83574) );
  NOR U103189 ( .A(n83572), .B(n83574), .Z(n89307) );
  IV U103190 ( .A(n83573), .Z(n83575) );
  NOR U103191 ( .A(n83575), .B(n83574), .Z(n89294) );
  IV U103192 ( .A(n83576), .Z(n83577) );
  NOR U103193 ( .A(n83578), .B(n83577), .Z(n83585) );
  IV U103194 ( .A(n83590), .Z(n83580) );
  NOR U103195 ( .A(n83580), .B(n83579), .Z(n83583) );
  IV U103196 ( .A(n83581), .Z(n83582) );
  NOR U103197 ( .A(n83583), .B(n83582), .Z(n83584) );
  NOR U103198 ( .A(n83585), .B(n83584), .Z(n83592) );
  IV U103199 ( .A(n83586), .Z(n83588) );
  NOR U103200 ( .A(n83588), .B(n83587), .Z(n83594) );
  IV U103201 ( .A(n83594), .Z(n83589) );
  NOR U103202 ( .A(n83592), .B(n83589), .Z(n89291) );
  NOR U103203 ( .A(n83591), .B(n83590), .Z(n83597) );
  IV U103204 ( .A(n83592), .Z(n83593) );
  NOR U103205 ( .A(n83594), .B(n83593), .Z(n83595) );
  IV U103206 ( .A(n83595), .Z(n83596) );
  NOR U103207 ( .A(n83597), .B(n83596), .Z(n89293) );
  NOR U103208 ( .A(n89291), .B(n89293), .Z(n83604) );
  NOR U103209 ( .A(n83599), .B(n83598), .Z(n89297) );
  IV U103210 ( .A(n83600), .Z(n83602) );
  NOR U103211 ( .A(n83602), .B(n83601), .Z(n89288) );
  NOR U103212 ( .A(n89297), .B(n89288), .Z(n83603) );
  XOR U103213 ( .A(n83604), .B(n83603), .Z(n83613) );
  NOR U103214 ( .A(n83606), .B(n83605), .Z(n83612) );
  IV U103215 ( .A(n83606), .Z(n83607) );
  NOR U103216 ( .A(n83608), .B(n83607), .Z(n83609) );
  NOR U103217 ( .A(n83610), .B(n83609), .Z(n83611) );
  NOR U103218 ( .A(n83612), .B(n83611), .Z(n89287) );
  XOR U103219 ( .A(n83613), .B(n89287), .Z(n89296) );
  XOR U103220 ( .A(n89294), .B(n89296), .Z(n89308) );
  XOR U103221 ( .A(n89307), .B(n89308), .Z(n89310) );
  IV U103222 ( .A(n83614), .Z(n83615) );
  NOR U103223 ( .A(n83616), .B(n83615), .Z(n83621) );
  IV U103224 ( .A(n83617), .Z(n83619) );
  NOR U103225 ( .A(n83619), .B(n83618), .Z(n83620) );
  NOR U103226 ( .A(n83621), .B(n83620), .Z(n89311) );
  XOR U103227 ( .A(n89310), .B(n89311), .Z(n83622) );
  IV U103228 ( .A(n83622), .Z(n89305) );
  XOR U103229 ( .A(n89304), .B(n89305), .Z(n89333) );
  XOR U103230 ( .A(n89332), .B(n89333), .Z(n83631) );
  IV U103231 ( .A(n83631), .Z(n83627) );
  IV U103232 ( .A(n83623), .Z(n83625) );
  NOR U103233 ( .A(n83625), .B(n83624), .Z(n83635) );
  IV U103234 ( .A(n83635), .Z(n83626) );
  NOR U103235 ( .A(n83627), .B(n83626), .Z(n89334) );
  NOR U103236 ( .A(n83629), .B(n83628), .Z(n83632) );
  IV U103237 ( .A(n83632), .Z(n83630) );
  NOR U103238 ( .A(n83630), .B(n89305), .Z(n89338) );
  NOR U103239 ( .A(n83632), .B(n83631), .Z(n83633) );
  NOR U103240 ( .A(n89338), .B(n83633), .Z(n83634) );
  NOR U103241 ( .A(n83635), .B(n83634), .Z(n83636) );
  NOR U103242 ( .A(n89334), .B(n83636), .Z(n83637) );
  IV U103243 ( .A(n83637), .Z(n89320) );
  XOR U103244 ( .A(n89319), .B(n89320), .Z(n89324) );
  IV U103245 ( .A(n83638), .Z(n83640) );
  NOR U103246 ( .A(n83640), .B(n83639), .Z(n83641) );
  IV U103247 ( .A(n83641), .Z(n83642) );
  NOR U103248 ( .A(n83643), .B(n83642), .Z(n89322) );
  XOR U103249 ( .A(n89324), .B(n89322), .Z(n89347) );
  XOR U103250 ( .A(n89346), .B(n89347), .Z(n89329) );
  XOR U103251 ( .A(n83644), .B(n89329), .Z(n89280) );
  IV U103252 ( .A(n83645), .Z(n83646) );
  NOR U103253 ( .A(n83647), .B(n83646), .Z(n83652) );
  IV U103254 ( .A(n83648), .Z(n83650) );
  NOR U103255 ( .A(n83650), .B(n83649), .Z(n83651) );
  NOR U103256 ( .A(n83652), .B(n83651), .Z(n89281) );
  XOR U103257 ( .A(n89280), .B(n89281), .Z(n89283) );
  XOR U103258 ( .A(n89284), .B(n89283), .Z(n83653) );
  IV U103259 ( .A(n83653), .Z(n89273) );
  NOR U103260 ( .A(n89276), .B(n89273), .Z(n83660) );
  NOR U103261 ( .A(n83654), .B(n83653), .Z(n83658) );
  IV U103262 ( .A(n83655), .Z(n83657) );
  NOR U103263 ( .A(n83657), .B(n83656), .Z(n89275) );
  XOR U103264 ( .A(n83658), .B(n89275), .Z(n83659) );
  NOR U103265 ( .A(n83660), .B(n83659), .Z(n89235) );
  IV U103266 ( .A(n83661), .Z(n83662) );
  NOR U103267 ( .A(n83663), .B(n83662), .Z(n83664) );
  IV U103268 ( .A(n83664), .Z(n89236) );
  XOR U103269 ( .A(n89235), .B(n89236), .Z(n89238) );
  XOR U103270 ( .A(n89239), .B(n89238), .Z(n83665) );
  IV U103271 ( .A(n83665), .Z(n89243) );
  XOR U103272 ( .A(n89242), .B(n89243), .Z(n89262) );
  NOR U103273 ( .A(n83666), .B(n89262), .Z(n89248) );
  NOR U103274 ( .A(n83668), .B(n83667), .Z(n83669) );
  IV U103275 ( .A(n83669), .Z(n89263) );
  XOR U103276 ( .A(n89263), .B(n89262), .Z(n83670) );
  NOR U103277 ( .A(n83671), .B(n83670), .Z(n89246) );
  XOR U103278 ( .A(n89246), .B(n89245), .Z(n83672) );
  NOR U103279 ( .A(n89248), .B(n83672), .Z(n83673) );
  IV U103280 ( .A(n83673), .Z(n89265) );
  XOR U103281 ( .A(n89264), .B(n89265), .Z(n89256) );
  IV U103282 ( .A(n83674), .Z(n83676) );
  NOR U103283 ( .A(n83676), .B(n83675), .Z(n89254) );
  XOR U103284 ( .A(n89256), .B(n89254), .Z(n89258) );
  XOR U103285 ( .A(n89257), .B(n89258), .Z(n89234) );
  IV U103286 ( .A(n83677), .Z(n83678) );
  NOR U103287 ( .A(n83679), .B(n83678), .Z(n89232) );
  XOR U103288 ( .A(n89234), .B(n89232), .Z(n89225) );
  XOR U103289 ( .A(n89224), .B(n89225), .Z(n89228) );
  XOR U103290 ( .A(n89227), .B(n89228), .Z(n89217) );
  IV U103291 ( .A(n83680), .Z(n83682) );
  NOR U103292 ( .A(n83682), .B(n83681), .Z(n83687) );
  IV U103293 ( .A(n83683), .Z(n83684) );
  NOR U103294 ( .A(n83685), .B(n83684), .Z(n83686) );
  NOR U103295 ( .A(n83687), .B(n83686), .Z(n89218) );
  XOR U103296 ( .A(n89217), .B(n89218), .Z(n89213) );
  XOR U103297 ( .A(n89210), .B(n89213), .Z(n89220) );
  XOR U103298 ( .A(n83688), .B(n89220), .Z(n89376) );
  XOR U103299 ( .A(n89377), .B(n89376), .Z(n89379) );
  XOR U103300 ( .A(n89380), .B(n89379), .Z(n89369) );
  XOR U103301 ( .A(n89370), .B(n89369), .Z(n89372) );
  XOR U103302 ( .A(n89373), .B(n89372), .Z(n89205) );
  XOR U103303 ( .A(n89202), .B(n89205), .Z(n89189) );
  XOR U103304 ( .A(n83689), .B(n89189), .Z(n83690) );
  IV U103305 ( .A(n83690), .Z(n89187) );
  XOR U103306 ( .A(n89185), .B(n89187), .Z(n89178) );
  XOR U103307 ( .A(n89177), .B(n89178), .Z(n89181) );
  XOR U103308 ( .A(n89180), .B(n89181), .Z(n89195) );
  NOR U103309 ( .A(n83692), .B(n83691), .Z(n83693) );
  IV U103310 ( .A(n83693), .Z(n83696) );
  IV U103311 ( .A(n83694), .Z(n83695) );
  NOR U103312 ( .A(n83696), .B(n83695), .Z(n89193) );
  XOR U103313 ( .A(n89195), .B(n89193), .Z(n89197) );
  XOR U103314 ( .A(n89196), .B(n89197), .Z(n89425) );
  IV U103315 ( .A(n83697), .Z(n83699) );
  NOR U103316 ( .A(n83699), .B(n83698), .Z(n89424) );
  IV U103317 ( .A(n83700), .Z(n83702) );
  NOR U103318 ( .A(n83702), .B(n83701), .Z(n89394) );
  NOR U103319 ( .A(n89424), .B(n89394), .Z(n83703) );
  XOR U103320 ( .A(n89425), .B(n83703), .Z(n89392) );
  IV U103321 ( .A(n83704), .Z(n83705) );
  NOR U103322 ( .A(n83706), .B(n83705), .Z(n89391) );
  NOR U103323 ( .A(n83708), .B(n83707), .Z(n89428) );
  NOR U103324 ( .A(n89391), .B(n89428), .Z(n83709) );
  XOR U103325 ( .A(n89392), .B(n83709), .Z(n89422) );
  XOR U103326 ( .A(n89423), .B(n89422), .Z(n89399) );
  XOR U103327 ( .A(n89401), .B(n89399), .Z(n89417) );
  XOR U103328 ( .A(n83710), .B(n89417), .Z(n83716) );
  IV U103329 ( .A(n83711), .Z(n83713) );
  NOR U103330 ( .A(n83713), .B(n83712), .Z(n89412) );
  XOR U103331 ( .A(n83716), .B(n89412), .Z(n83714) );
  NOR U103332 ( .A(n83717), .B(n83714), .Z(n83722) );
  IV U103333 ( .A(n83722), .Z(n83715) );
  NOR U103334 ( .A(n83720), .B(n83715), .Z(n83723) );
  IV U103335 ( .A(n83716), .Z(n89414) );
  IV U103336 ( .A(n83717), .Z(n83718) );
  NOR U103337 ( .A(n89414), .B(n83718), .Z(n83719) );
  NOR U103338 ( .A(n83720), .B(n83719), .Z(n83721) );
  NOR U103339 ( .A(n83722), .B(n83721), .Z(n89176) );
  NOR U103340 ( .A(n83723), .B(n89176), .Z(n89172) );
  XOR U103341 ( .A(n89174), .B(n89172), .Z(n83731) );
  IV U103342 ( .A(n83731), .Z(n83724) );
  NOR U103343 ( .A(n83730), .B(n83724), .Z(n83725) );
  IV U103344 ( .A(n83725), .Z(n83729) );
  IV U103345 ( .A(n83726), .Z(n83727) );
  NOR U103346 ( .A(n83728), .B(n83727), .Z(n83733) );
  NOR U103347 ( .A(n83729), .B(n83733), .Z(n83739) );
  IV U103348 ( .A(n83730), .Z(n83734) );
  XOR U103349 ( .A(n83733), .B(n83734), .Z(n83732) );
  NOR U103350 ( .A(n83732), .B(n83731), .Z(n83737) );
  IV U103351 ( .A(n83733), .Z(n83735) );
  NOR U103352 ( .A(n83735), .B(n83734), .Z(n83736) );
  NOR U103353 ( .A(n83737), .B(n83736), .Z(n89421) );
  IV U103354 ( .A(n89421), .Z(n83738) );
  NOR U103355 ( .A(n83739), .B(n83738), .Z(n89162) );
  IV U103356 ( .A(n83740), .Z(n83742) );
  NOR U103357 ( .A(n83742), .B(n83741), .Z(n83747) );
  IV U103358 ( .A(n83743), .Z(n83745) );
  NOR U103359 ( .A(n83745), .B(n83744), .Z(n83746) );
  NOR U103360 ( .A(n83747), .B(n83746), .Z(n89164) );
  XOR U103361 ( .A(n89162), .B(n89164), .Z(n89166) );
  XOR U103362 ( .A(n89165), .B(n89166), .Z(n89155) );
  XOR U103363 ( .A(n89154), .B(n89155), .Z(n89158) );
  XOR U103364 ( .A(n89157), .B(n89158), .Z(n83755) );
  NOR U103365 ( .A(n83758), .B(n83755), .Z(n83753) );
  IV U103366 ( .A(n83748), .Z(n83750) );
  NOR U103367 ( .A(n83750), .B(n83749), .Z(n83756) );
  IV U103368 ( .A(n83756), .Z(n83751) );
  NOR U103369 ( .A(n89158), .B(n83751), .Z(n83752) );
  NOR U103370 ( .A(n83753), .B(n83752), .Z(n83754) );
  IV U103371 ( .A(n83754), .Z(n89441) );
  IV U103372 ( .A(n83755), .Z(n83759) );
  NOR U103373 ( .A(n83756), .B(n83759), .Z(n83757) );
  NOR U103374 ( .A(n89441), .B(n83757), .Z(n83761) );
  NOR U103375 ( .A(n83759), .B(n83758), .Z(n83760) );
  NOR U103376 ( .A(n83761), .B(n83760), .Z(n89148) );
  XOR U103377 ( .A(n89146), .B(n89148), .Z(n89150) );
  XOR U103378 ( .A(n89149), .B(n89150), .Z(n89144) );
  XOR U103379 ( .A(n89143), .B(n89144), .Z(n89132) );
  XOR U103380 ( .A(n89130), .B(n89132), .Z(n89136) );
  XOR U103381 ( .A(n89137), .B(n89136), .Z(n83762) );
  IV U103382 ( .A(n83762), .Z(n89133) );
  IV U103383 ( .A(n83763), .Z(n83765) );
  NOR U103384 ( .A(n83765), .B(n83764), .Z(n83770) );
  IV U103385 ( .A(n83766), .Z(n83767) );
  NOR U103386 ( .A(n83768), .B(n83767), .Z(n83769) );
  NOR U103387 ( .A(n83770), .B(n83769), .Z(n89134) );
  XOR U103388 ( .A(n89133), .B(n89134), .Z(n89452) );
  XOR U103389 ( .A(n89453), .B(n89452), .Z(n83771) );
  XOR U103390 ( .A(n83772), .B(n83771), .Z(n89128) );
  XOR U103391 ( .A(n83773), .B(n89128), .Z(n89478) );
  XOR U103392 ( .A(n89476), .B(n89478), .Z(n89479) );
  XOR U103393 ( .A(n89480), .B(n89479), .Z(n83774) );
  IV U103394 ( .A(n83774), .Z(n89114) );
  NOR U103395 ( .A(n89117), .B(n89114), .Z(n83781) );
  NOR U103396 ( .A(n83775), .B(n83774), .Z(n83779) );
  IV U103397 ( .A(n83776), .Z(n83777) );
  NOR U103398 ( .A(n83778), .B(n83777), .Z(n89116) );
  XOR U103399 ( .A(n83779), .B(n89116), .Z(n83780) );
  NOR U103400 ( .A(n83781), .B(n83780), .Z(n83782) );
  IV U103401 ( .A(n83782), .Z(n89123) );
  XOR U103402 ( .A(n89122), .B(n89123), .Z(n89471) );
  XOR U103403 ( .A(n89469), .B(n89471), .Z(n89472) );
  XOR U103404 ( .A(n89473), .B(n89472), .Z(n89507) );
  IV U103405 ( .A(n83783), .Z(n83784) );
  NOR U103406 ( .A(n83784), .B(n83788), .Z(n83785) );
  IV U103407 ( .A(n83785), .Z(n89508) );
  XOR U103408 ( .A(n89507), .B(n89508), .Z(n89510) );
  NOR U103409 ( .A(n83786), .B(n83793), .Z(n83791) );
  IV U103410 ( .A(n83787), .Z(n83789) );
  NOR U103411 ( .A(n83789), .B(n83788), .Z(n83790) );
  NOR U103412 ( .A(n83791), .B(n83790), .Z(n89511) );
  XOR U103413 ( .A(n89510), .B(n89511), .Z(n89498) );
  IV U103414 ( .A(n89498), .Z(n89489) );
  NOR U103415 ( .A(n83793), .B(n83792), .Z(n89499) );
  IV U103416 ( .A(n89499), .Z(n89490) );
  IV U103417 ( .A(n83794), .Z(n83795) );
  NOR U103418 ( .A(n89103), .B(n83795), .Z(n83798) );
  NOR U103419 ( .A(n89493), .B(n83796), .Z(n83797) );
  NOR U103420 ( .A(n83798), .B(n83797), .Z(n89500) );
  XOR U103421 ( .A(n89490), .B(n89500), .Z(n83799) );
  XOR U103422 ( .A(n89489), .B(n83799), .Z(n89102) );
  XOR U103423 ( .A(n83800), .B(n89102), .Z(n89100) );
  XOR U103424 ( .A(n89098), .B(n89100), .Z(n89079) );
  XOR U103425 ( .A(n89078), .B(n89079), .Z(n89082) );
  XOR U103426 ( .A(n89081), .B(n89082), .Z(n89091) );
  XOR U103427 ( .A(n89092), .B(n89091), .Z(n89088) );
  XOR U103428 ( .A(n89090), .B(n89088), .Z(n89086) );
  XOR U103429 ( .A(n89087), .B(n89086), .Z(n83801) );
  IV U103430 ( .A(n83801), .Z(n89071) );
  NOR U103431 ( .A(n89074), .B(n89071), .Z(n83808) );
  NOR U103432 ( .A(n83802), .B(n83801), .Z(n83806) );
  IV U103433 ( .A(n83803), .Z(n83804) );
  NOR U103434 ( .A(n83805), .B(n83804), .Z(n89073) );
  XOR U103435 ( .A(n83806), .B(n89073), .Z(n83807) );
  NOR U103436 ( .A(n83808), .B(n83807), .Z(n89063) );
  XOR U103437 ( .A(n89065), .B(n89063), .Z(n89067) );
  XOR U103438 ( .A(n89066), .B(n89067), .Z(n89528) );
  IV U103439 ( .A(n83809), .Z(n83811) );
  NOR U103440 ( .A(n83811), .B(n83810), .Z(n89526) );
  XOR U103441 ( .A(n89528), .B(n89526), .Z(n89545) );
  IV U103442 ( .A(n89545), .Z(n83819) );
  IV U103443 ( .A(n83812), .Z(n83813) );
  NOR U103444 ( .A(n83814), .B(n83813), .Z(n89527) );
  IV U103445 ( .A(n83815), .Z(n83817) );
  NOR U103446 ( .A(n83817), .B(n83816), .Z(n89544) );
  NOR U103447 ( .A(n89527), .B(n89544), .Z(n83818) );
  XOR U103448 ( .A(n83819), .B(n83818), .Z(n89538) );
  XOR U103449 ( .A(n89536), .B(n89538), .Z(n89540) );
  XOR U103450 ( .A(n89539), .B(n89540), .Z(n89056) );
  XOR U103451 ( .A(n89055), .B(n89056), .Z(n89059) );
  XOR U103452 ( .A(n89058), .B(n89059), .Z(n89561) );
  XOR U103453 ( .A(n89560), .B(n89561), .Z(n89564) );
  XOR U103454 ( .A(n89563), .B(n89564), .Z(n89555) );
  XOR U103455 ( .A(n89553), .B(n89555), .Z(n89556) );
  XOR U103456 ( .A(n89557), .B(n89556), .Z(n89572) );
  IV U103457 ( .A(n83820), .Z(n83822) );
  NOR U103458 ( .A(n83822), .B(n83821), .Z(n89573) );
  IV U103459 ( .A(n83823), .Z(n83824) );
  NOR U103460 ( .A(n83825), .B(n83824), .Z(n83826) );
  NOR U103461 ( .A(n83827), .B(n83826), .Z(n89574) );
  XOR U103462 ( .A(n89573), .B(n89574), .Z(n83828) );
  XOR U103463 ( .A(n89572), .B(n83828), .Z(n89049) );
  XOR U103464 ( .A(n89047), .B(n89049), .Z(n89052) );
  IV U103465 ( .A(n83829), .Z(n83831) );
  NOR U103466 ( .A(n83831), .B(n83830), .Z(n89050) );
  XOR U103467 ( .A(n89052), .B(n89050), .Z(n89031) );
  IV U103468 ( .A(n83832), .Z(n83833) );
  NOR U103469 ( .A(n83834), .B(n83833), .Z(n83838) );
  NOR U103470 ( .A(n83836), .B(n83835), .Z(n83837) );
  NOR U103471 ( .A(n83838), .B(n83837), .Z(n89032) );
  XOR U103472 ( .A(n89031), .B(n89032), .Z(n89033) );
  XOR U103473 ( .A(n89035), .B(n89033), .Z(n89044) );
  IV U103474 ( .A(n83839), .Z(n83844) );
  NOR U103475 ( .A(n83841), .B(n83840), .Z(n83842) );
  IV U103476 ( .A(n83842), .Z(n83843) );
  NOR U103477 ( .A(n83844), .B(n83843), .Z(n89041) );
  XOR U103478 ( .A(n89044), .B(n89041), .Z(n89040) );
  XOR U103479 ( .A(n89042), .B(n89040), .Z(n83845) );
  XOR U103480 ( .A(n89038), .B(n83845), .Z(n88990) );
  IV U103481 ( .A(n83846), .Z(n83847) );
  NOR U103482 ( .A(n83848), .B(n83847), .Z(n83854) );
  IV U103483 ( .A(n83849), .Z(n83852) );
  IV U103484 ( .A(n83850), .Z(n83851) );
  NOR U103485 ( .A(n83852), .B(n83851), .Z(n83853) );
  NOR U103486 ( .A(n83854), .B(n83853), .Z(n88991) );
  XOR U103487 ( .A(n88990), .B(n88991), .Z(n88992) );
  XOR U103488 ( .A(n88994), .B(n88992), .Z(n88983) );
  XOR U103489 ( .A(n88982), .B(n88983), .Z(n88986) );
  XOR U103490 ( .A(n88985), .B(n88986), .Z(n89029) );
  XOR U103491 ( .A(n89027), .B(n89029), .Z(n89001) );
  XOR U103492 ( .A(n83855), .B(n89001), .Z(n83856) );
  IV U103493 ( .A(n83856), .Z(n89004) );
  XOR U103494 ( .A(n89002), .B(n89004), .Z(n89007) );
  IV U103495 ( .A(n83857), .Z(n83859) );
  IV U103496 ( .A(n83858), .Z(n89598) );
  NOR U103497 ( .A(n83859), .B(n89598), .Z(n89005) );
  XOR U103498 ( .A(n89007), .B(n89005), .Z(n89594) );
  NOR U103499 ( .A(n83861), .B(n83860), .Z(n83864) );
  IV U103500 ( .A(n89592), .Z(n83862) );
  NOR U103501 ( .A(n83862), .B(n89598), .Z(n83863) );
  NOR U103502 ( .A(n83864), .B(n83863), .Z(n89016) );
  XOR U103503 ( .A(n89594), .B(n89016), .Z(n89013) );
  XOR U103504 ( .A(n89015), .B(n89013), .Z(n83866) );
  NOR U103505 ( .A(n83865), .B(n83866), .Z(n89619) );
  IV U103506 ( .A(n83866), .Z(n83867) );
  NOR U103507 ( .A(n83868), .B(n83867), .Z(n89617) );
  IV U103508 ( .A(n83869), .Z(n83874) );
  NOR U103509 ( .A(n83871), .B(n83870), .Z(n83872) );
  IV U103510 ( .A(n83872), .Z(n83873) );
  NOR U103511 ( .A(n83874), .B(n83873), .Z(n89616) );
  XOR U103512 ( .A(n89617), .B(n89616), .Z(n83875) );
  NOR U103513 ( .A(n89619), .B(n83875), .Z(n83876) );
  NOR U103514 ( .A(n83883), .B(n83876), .Z(n83885) );
  IV U103515 ( .A(n83877), .Z(n83878) );
  NOR U103516 ( .A(n83878), .B(n83881), .Z(n83879) );
  IV U103517 ( .A(n83879), .Z(n83886) );
  NOR U103518 ( .A(n83885), .B(n83886), .Z(n89610) );
  IV U103519 ( .A(n83880), .Z(n83882) );
  NOR U103520 ( .A(n83882), .B(n83881), .Z(n89601) );
  IV U103521 ( .A(n83883), .Z(n83884) );
  NOR U103522 ( .A(n89617), .B(n83884), .Z(n89611) );
  NOR U103523 ( .A(n83885), .B(n89611), .Z(n89602) );
  XOR U103524 ( .A(n89601), .B(n89602), .Z(n83888) );
  NOR U103525 ( .A(n89602), .B(n83886), .Z(n83887) );
  NOR U103526 ( .A(n83888), .B(n83887), .Z(n83889) );
  NOR U103527 ( .A(n89610), .B(n83889), .Z(n83890) );
  IV U103528 ( .A(n83890), .Z(n89606) );
  XOR U103529 ( .A(n89605), .B(n89606), .Z(n89622) );
  XOR U103530 ( .A(n89621), .B(n89622), .Z(n88972) );
  IV U103531 ( .A(n83891), .Z(n83893) );
  NOR U103532 ( .A(n83893), .B(n83892), .Z(n88970) );
  XOR U103533 ( .A(n88972), .B(n88970), .Z(n88974) );
  XOR U103534 ( .A(n88973), .B(n88974), .Z(n88980) );
  XOR U103535 ( .A(n88978), .B(n88980), .Z(n89634) );
  IV U103536 ( .A(n83894), .Z(n83895) );
  NOR U103537 ( .A(n83896), .B(n83895), .Z(n88979) );
  IV U103538 ( .A(n83897), .Z(n83899) );
  NOR U103539 ( .A(n83899), .B(n83898), .Z(n89632) );
  NOR U103540 ( .A(n88979), .B(n89632), .Z(n83900) );
  XOR U103541 ( .A(n89634), .B(n83900), .Z(n89635) );
  IV U103542 ( .A(n83901), .Z(n83903) );
  NOR U103543 ( .A(n83903), .B(n83902), .Z(n83904) );
  IV U103544 ( .A(n83904), .Z(n89636) );
  XOR U103545 ( .A(n89635), .B(n89636), .Z(n89639) );
  XOR U103546 ( .A(n89638), .B(n89639), .Z(n89655) );
  XOR U103547 ( .A(n89653), .B(n89655), .Z(n89657) );
  XOR U103548 ( .A(n89656), .B(n89657), .Z(n89647) );
  XOR U103549 ( .A(n89646), .B(n89647), .Z(n89649) );
  XOR U103550 ( .A(n89650), .B(n89649), .Z(n83905) );
  IV U103551 ( .A(n83905), .Z(n89676) );
  XOR U103552 ( .A(n89675), .B(n89676), .Z(n89679) );
  XOR U103553 ( .A(n89678), .B(n89679), .Z(n89669) );
  IV U103554 ( .A(n83906), .Z(n83909) );
  IV U103555 ( .A(n83907), .Z(n83908) );
  NOR U103556 ( .A(n83909), .B(n83908), .Z(n89667) );
  XOR U103557 ( .A(n89669), .B(n89667), .Z(n89671) );
  XOR U103558 ( .A(n88965), .B(n89671), .Z(n83913) );
  IV U103559 ( .A(n83910), .Z(n83911) );
  NOR U103560 ( .A(n83912), .B(n83911), .Z(n89670) );
  XOR U103561 ( .A(n83913), .B(n89670), .Z(n83914) );
  NOR U103562 ( .A(n88964), .B(n83914), .Z(n83918) );
  IV U103563 ( .A(n88964), .Z(n88961) );
  IV U103564 ( .A(n89671), .Z(n88962) );
  NOR U103565 ( .A(n88965), .B(n88962), .Z(n83915) );
  IV U103566 ( .A(n83915), .Z(n83916) );
  NOR U103567 ( .A(n88961), .B(n83916), .Z(n83917) );
  NOR U103568 ( .A(n83918), .B(n83917), .Z(n89701) );
  NOR U103569 ( .A(n83920), .B(n83919), .Z(n83921) );
  NOR U103570 ( .A(n83922), .B(n83921), .Z(n89699) );
  XOR U103571 ( .A(n89701), .B(n89699), .Z(n89703) );
  XOR U103572 ( .A(n89702), .B(n89703), .Z(n89694) );
  IV U103573 ( .A(n83923), .Z(n83925) );
  NOR U103574 ( .A(n83925), .B(n83924), .Z(n89692) );
  XOR U103575 ( .A(n89694), .B(n89692), .Z(n89695) );
  IV U103576 ( .A(n83926), .Z(n83927) );
  NOR U103577 ( .A(n83928), .B(n83927), .Z(n83933) );
  IV U103578 ( .A(n83929), .Z(n83931) );
  NOR U103579 ( .A(n83931), .B(n83930), .Z(n83932) );
  NOR U103580 ( .A(n83933), .B(n83932), .Z(n89696) );
  XOR U103581 ( .A(n89695), .B(n89696), .Z(n88954) );
  XOR U103582 ( .A(n83934), .B(n88954), .Z(n88957) );
  XOR U103583 ( .A(n88956), .B(n88957), .Z(n89720) );
  XOR U103584 ( .A(n89719), .B(n89720), .Z(n89723) );
  XOR U103585 ( .A(n89722), .B(n89723), .Z(n89714) );
  XOR U103586 ( .A(n89713), .B(n89714), .Z(n89740) );
  IV U103587 ( .A(n83935), .Z(n83936) );
  NOR U103588 ( .A(n83937), .B(n83936), .Z(n89741) );
  IV U103589 ( .A(n83938), .Z(n83940) );
  NOR U103590 ( .A(n83940), .B(n83939), .Z(n89733) );
  NOR U103591 ( .A(n89741), .B(n89733), .Z(n83941) );
  XOR U103592 ( .A(n89740), .B(n83941), .Z(n83942) );
  IV U103593 ( .A(n83942), .Z(n89736) );
  XOR U103594 ( .A(n89735), .B(n89736), .Z(n88951) );
  XOR U103595 ( .A(n83943), .B(n88951), .Z(n83944) );
  IV U103596 ( .A(n83944), .Z(n89755) );
  XOR U103597 ( .A(n89753), .B(n89755), .Z(n89758) );
  IV U103598 ( .A(n83945), .Z(n83947) );
  NOR U103599 ( .A(n83947), .B(n83946), .Z(n89756) );
  XOR U103600 ( .A(n89758), .B(n89756), .Z(n89761) );
  IV U103601 ( .A(n83948), .Z(n83949) );
  NOR U103602 ( .A(n83950), .B(n83949), .Z(n83955) );
  IV U103603 ( .A(n83951), .Z(n83953) );
  NOR U103604 ( .A(n83953), .B(n83952), .Z(n83954) );
  NOR U103605 ( .A(n83955), .B(n83954), .Z(n89762) );
  XOR U103606 ( .A(n89761), .B(n89762), .Z(n89763) );
  XOR U103607 ( .A(n89765), .B(n89763), .Z(n88944) );
  IV U103608 ( .A(n83956), .Z(n83957) );
  NOR U103609 ( .A(n83958), .B(n83957), .Z(n88942) );
  XOR U103610 ( .A(n88944), .B(n88942), .Z(n88940) );
  XOR U103611 ( .A(n88939), .B(n88940), .Z(n88938) );
  IV U103612 ( .A(n83959), .Z(n83960) );
  NOR U103613 ( .A(n83961), .B(n83960), .Z(n88936) );
  XOR U103614 ( .A(n88938), .B(n88936), .Z(n88894) );
  XOR U103615 ( .A(n88893), .B(n88894), .Z(n88901) );
  NOR U103616 ( .A(n83963), .B(n83962), .Z(n88892) );
  IV U103617 ( .A(n83964), .Z(n83968) );
  NOR U103618 ( .A(n83966), .B(n83965), .Z(n83967) );
  IV U103619 ( .A(n83967), .Z(n83971) );
  NOR U103620 ( .A(n83968), .B(n83971), .Z(n88899) );
  NOR U103621 ( .A(n88892), .B(n88899), .Z(n83969) );
  XOR U103622 ( .A(n88901), .B(n83969), .Z(n88896) );
  IV U103623 ( .A(n83970), .Z(n83972) );
  NOR U103624 ( .A(n83972), .B(n83971), .Z(n83973) );
  IV U103625 ( .A(n83973), .Z(n88897) );
  XOR U103626 ( .A(n88896), .B(n88897), .Z(n88907) );
  XOR U103627 ( .A(n88906), .B(n88907), .Z(n88910) );
  XOR U103628 ( .A(n88909), .B(n88910), .Z(n88891) );
  XOR U103629 ( .A(n88889), .B(n88891), .Z(n88925) );
  XOR U103630 ( .A(n88924), .B(n88925), .Z(n88928) );
  XOR U103631 ( .A(n88927), .B(n88928), .Z(n88917) );
  XOR U103632 ( .A(n88916), .B(n88917), .Z(n88920) );
  XOR U103633 ( .A(n88919), .B(n88920), .Z(n88865) );
  XOR U103634 ( .A(n88863), .B(n88865), .Z(n88867) );
  XOR U103635 ( .A(n88866), .B(n88867), .Z(n88877) );
  XOR U103636 ( .A(n83974), .B(n88877), .Z(n88879) );
  IV U103637 ( .A(n83975), .Z(n83976) );
  NOR U103638 ( .A(n83976), .B(n83993), .Z(n83986) );
  IV U103639 ( .A(n83986), .Z(n88880) );
  NOR U103640 ( .A(n88879), .B(n88880), .Z(n83988) );
  IV U103641 ( .A(n83977), .Z(n83979) );
  NOR U103642 ( .A(n83979), .B(n83978), .Z(n83982) );
  IV U103643 ( .A(n83982), .Z(n83981) );
  XOR U103644 ( .A(n88861), .B(n88877), .Z(n83980) );
  NOR U103645 ( .A(n83981), .B(n83980), .Z(n88886) );
  NOR U103646 ( .A(n88879), .B(n83982), .Z(n83983) );
  NOR U103647 ( .A(n88886), .B(n83983), .Z(n83984) );
  IV U103648 ( .A(n83984), .Z(n83985) );
  NOR U103649 ( .A(n83986), .B(n83985), .Z(n83987) );
  NOR U103650 ( .A(n83988), .B(n83987), .Z(n88853) );
  XOR U103651 ( .A(n88855), .B(n88853), .Z(n88832) );
  IV U103652 ( .A(n83989), .Z(n83991) );
  NOR U103653 ( .A(n83991), .B(n83990), .Z(n88830) );
  IV U103654 ( .A(n83992), .Z(n83994) );
  NOR U103655 ( .A(n83994), .B(n83993), .Z(n88856) );
  NOR U103656 ( .A(n88830), .B(n88856), .Z(n83995) );
  XOR U103657 ( .A(n88832), .B(n83995), .Z(n84004) );
  IV U103658 ( .A(n84004), .Z(n88829) );
  IV U103659 ( .A(n83996), .Z(n84000) );
  IV U103660 ( .A(n83997), .Z(n84008) );
  NOR U103661 ( .A(n83998), .B(n84008), .Z(n83999) );
  IV U103662 ( .A(n83999), .Z(n84011) );
  NOR U103663 ( .A(n84000), .B(n84011), .Z(n84006) );
  IV U103664 ( .A(n84006), .Z(n84001) );
  NOR U103665 ( .A(n88829), .B(n84001), .Z(n88824) );
  NOR U103666 ( .A(n84003), .B(n84002), .Z(n88827) );
  XOR U103667 ( .A(n84004), .B(n88827), .Z(n84005) );
  NOR U103668 ( .A(n84006), .B(n84005), .Z(n88826) );
  NOR U103669 ( .A(n88824), .B(n88826), .Z(n88840) );
  IV U103670 ( .A(n84007), .Z(n84009) );
  NOR U103671 ( .A(n84009), .B(n84008), .Z(n88839) );
  IV U103672 ( .A(n84010), .Z(n84012) );
  NOR U103673 ( .A(n84012), .B(n84011), .Z(n88823) );
  NOR U103674 ( .A(n88839), .B(n88823), .Z(n84013) );
  XOR U103675 ( .A(n88840), .B(n84013), .Z(n88838) );
  XOR U103676 ( .A(n88837), .B(n88838), .Z(n84025) );
  IV U103677 ( .A(n84025), .Z(n84022) );
  IV U103678 ( .A(n84014), .Z(n84016) );
  NOR U103679 ( .A(n84016), .B(n84015), .Z(n84021) );
  IV U103680 ( .A(n84017), .Z(n84019) );
  NOR U103681 ( .A(n84019), .B(n84018), .Z(n84020) );
  NOR U103682 ( .A(n84021), .B(n84020), .Z(n84023) );
  NOR U103683 ( .A(n84022), .B(n84023), .Z(n88851) );
  IV U103684 ( .A(n84023), .Z(n84024) );
  NOR U103685 ( .A(n84025), .B(n84024), .Z(n88848) );
  NOR U103686 ( .A(n84027), .B(n84026), .Z(n88847) );
  XOR U103687 ( .A(n88848), .B(n88847), .Z(n84028) );
  NOR U103688 ( .A(n88851), .B(n84028), .Z(n88813) );
  IV U103689 ( .A(n84029), .Z(n84030) );
  NOR U103690 ( .A(n84031), .B(n84030), .Z(n84032) );
  IV U103691 ( .A(n84032), .Z(n88814) );
  XOR U103692 ( .A(n88813), .B(n88814), .Z(n88818) );
  XOR U103693 ( .A(n88816), .B(n88818), .Z(n88806) );
  XOR U103694 ( .A(n88805), .B(n88806), .Z(n88809) );
  XOR U103695 ( .A(n88808), .B(n88809), .Z(n88784) );
  IV U103696 ( .A(n84033), .Z(n84034) );
  NOR U103697 ( .A(n84035), .B(n84034), .Z(n88782) );
  IV U103698 ( .A(n84036), .Z(n84037) );
  NOR U103699 ( .A(n84038), .B(n84037), .Z(n88783) );
  NOR U103700 ( .A(n88782), .B(n88783), .Z(n84039) );
  XOR U103701 ( .A(n88784), .B(n84039), .Z(n84040) );
  NOR U103702 ( .A(n84041), .B(n84040), .Z(n84044) );
  IV U103703 ( .A(n84041), .Z(n84043) );
  XOR U103704 ( .A(n88782), .B(n88784), .Z(n84042) );
  NOR U103705 ( .A(n84043), .B(n84042), .Z(n88804) );
  NOR U103706 ( .A(n84044), .B(n88804), .Z(n84045) );
  IV U103707 ( .A(n84045), .Z(n88802) );
  NOR U103708 ( .A(n84046), .B(n84047), .Z(n84053) );
  IV U103709 ( .A(n84047), .Z(n84048) );
  NOR U103710 ( .A(n84049), .B(n84048), .Z(n84050) );
  NOR U103711 ( .A(n84051), .B(n84050), .Z(n84052) );
  NOR U103712 ( .A(n84053), .B(n84052), .Z(n88800) );
  XOR U103713 ( .A(n88802), .B(n88800), .Z(n88780) );
  XOR U103714 ( .A(n88781), .B(n88780), .Z(n84059) );
  IV U103715 ( .A(n84059), .Z(n88793) );
  NOR U103716 ( .A(n88795), .B(n88793), .Z(n84054) );
  IV U103717 ( .A(n84054), .Z(n84057) );
  XOR U103718 ( .A(n88795), .B(n88792), .Z(n84055) );
  NOR U103719 ( .A(n88789), .B(n84055), .Z(n84058) );
  IV U103720 ( .A(n84058), .Z(n84056) );
  NOR U103721 ( .A(n84057), .B(n84056), .Z(n84061) );
  NOR U103722 ( .A(n84059), .B(n84058), .Z(n84060) );
  NOR U103723 ( .A(n84061), .B(n84060), .Z(n88790) );
  XOR U103724 ( .A(n88791), .B(n88790), .Z(n88785) );
  IV U103725 ( .A(n88785), .Z(n88787) );
  IV U103726 ( .A(n84062), .Z(n84063) );
  NOR U103727 ( .A(n84067), .B(n84063), .Z(n84074) );
  IV U103728 ( .A(n84074), .Z(n84064) );
  NOR U103729 ( .A(n88787), .B(n84064), .Z(n89795) );
  IV U103730 ( .A(n84065), .Z(n84066) );
  NOR U103731 ( .A(n84067), .B(n84066), .Z(n88788) );
  IV U103732 ( .A(n84068), .Z(n84071) );
  IV U103733 ( .A(n84069), .Z(n84070) );
  NOR U103734 ( .A(n84071), .B(n84070), .Z(n88786) );
  NOR U103735 ( .A(n88788), .B(n88786), .Z(n84072) );
  XOR U103736 ( .A(n88787), .B(n84072), .Z(n84073) );
  NOR U103737 ( .A(n84074), .B(n84073), .Z(n89793) );
  IV U103738 ( .A(n84075), .Z(n84077) );
  NOR U103739 ( .A(n84077), .B(n84076), .Z(n89792) );
  XOR U103740 ( .A(n89793), .B(n89792), .Z(n84078) );
  NOR U103741 ( .A(n89795), .B(n84078), .Z(n89827) );
  NOR U103742 ( .A(n84080), .B(n84079), .Z(n89790) );
  IV U103743 ( .A(n84081), .Z(n84083) );
  NOR U103744 ( .A(n84083), .B(n84082), .Z(n89828) );
  NOR U103745 ( .A(n89790), .B(n89828), .Z(n84084) );
  XOR U103746 ( .A(n89827), .B(n84084), .Z(n89833) );
  XOR U103747 ( .A(n89831), .B(n89833), .Z(n89834) );
  XOR U103748 ( .A(n89835), .B(n89834), .Z(n84093) );
  IV U103749 ( .A(n84093), .Z(n84091) );
  XOR U103750 ( .A(n84086), .B(n84085), .Z(n84089) );
  IV U103751 ( .A(n84087), .Z(n84088) );
  NOR U103752 ( .A(n84089), .B(n84088), .Z(n84092) );
  IV U103753 ( .A(n84092), .Z(n84090) );
  NOR U103754 ( .A(n84091), .B(n84090), .Z(n89825) );
  NOR U103755 ( .A(n84093), .B(n84092), .Z(n89823) );
  IV U103756 ( .A(n84094), .Z(n84097) );
  IV U103757 ( .A(n84095), .Z(n84096) );
  NOR U103758 ( .A(n84097), .B(n84096), .Z(n89822) );
  XOR U103759 ( .A(n89823), .B(n89822), .Z(n84098) );
  NOR U103760 ( .A(n89825), .B(n84098), .Z(n84099) );
  IV U103761 ( .A(n84099), .Z(n89811) );
  XOR U103762 ( .A(n89810), .B(n89811), .Z(n89814) );
  XOR U103763 ( .A(n89813), .B(n89814), .Z(n89803) );
  XOR U103764 ( .A(n89802), .B(n89803), .Z(n89806) );
  XOR U103765 ( .A(n89805), .B(n89806), .Z(n88774) );
  IV U103766 ( .A(n84100), .Z(n84102) );
  NOR U103767 ( .A(n84102), .B(n84101), .Z(n88772) );
  XOR U103768 ( .A(n88774), .B(n88772), .Z(n88776) );
  XOR U103769 ( .A(n88775), .B(n88776), .Z(n89868) );
  IV U103770 ( .A(n84103), .Z(n84104) );
  NOR U103771 ( .A(n84105), .B(n84104), .Z(n84106) );
  IV U103772 ( .A(n84106), .Z(n84107) );
  NOR U103773 ( .A(n84108), .B(n84107), .Z(n89866) );
  XOR U103774 ( .A(n89868), .B(n89866), .Z(n89870) );
  XOR U103775 ( .A(n89869), .B(n89870), .Z(n89853) );
  XOR U103776 ( .A(n89852), .B(n89853), .Z(n89856) );
  XOR U103777 ( .A(n89855), .B(n89856), .Z(n89847) );
  IV U103778 ( .A(n84109), .Z(n84111) );
  NOR U103779 ( .A(n84111), .B(n84110), .Z(n89845) );
  XOR U103780 ( .A(n89847), .B(n89845), .Z(n89848) );
  XOR U103781 ( .A(n89849), .B(n89848), .Z(n84112) );
  NOR U103782 ( .A(n84116), .B(n84112), .Z(n84120) );
  IV U103783 ( .A(n84113), .Z(n84115) );
  NOR U103784 ( .A(n84115), .B(n84114), .Z(n84122) );
  IV U103785 ( .A(n84116), .Z(n84117) );
  NOR U103786 ( .A(n89848), .B(n84117), .Z(n84118) );
  NOR U103787 ( .A(n84122), .B(n84118), .Z(n84119) );
  NOR U103788 ( .A(n84120), .B(n84119), .Z(n89883) );
  IV U103789 ( .A(n84120), .Z(n84121) );
  NOR U103790 ( .A(n84122), .B(n84121), .Z(n84123) );
  NOR U103791 ( .A(n89883), .B(n84123), .Z(n84124) );
  IV U103792 ( .A(n84124), .Z(n89880) );
  XOR U103793 ( .A(n89879), .B(n89880), .Z(n89877) );
  XOR U103794 ( .A(n89876), .B(n89877), .Z(n84129) );
  IV U103795 ( .A(n84129), .Z(n84125) );
  NOR U103796 ( .A(n84128), .B(n84125), .Z(n84126) );
  IV U103797 ( .A(n84126), .Z(n84127) );
  NOR U103798 ( .A(n84131), .B(n84127), .Z(n89895) );
  IV U103799 ( .A(n84128), .Z(n84132) );
  XOR U103800 ( .A(n84131), .B(n84132), .Z(n84130) );
  NOR U103801 ( .A(n84130), .B(n84129), .Z(n84135) );
  IV U103802 ( .A(n84131), .Z(n84133) );
  NOR U103803 ( .A(n84133), .B(n84132), .Z(n84134) );
  NOR U103804 ( .A(n84135), .B(n84134), .Z(n84136) );
  IV U103805 ( .A(n84136), .Z(n89897) );
  NOR U103806 ( .A(n89895), .B(n89897), .Z(n88767) );
  XOR U103807 ( .A(n84137), .B(n88767), .Z(n89891) );
  XOR U103808 ( .A(n84138), .B(n89891), .Z(n84139) );
  IV U103809 ( .A(n84139), .Z(n89901) );
  XOR U103810 ( .A(n89902), .B(n89901), .Z(n84140) );
  NOR U103811 ( .A(n84141), .B(n84140), .Z(n89912) );
  IV U103812 ( .A(n84141), .Z(n84142) );
  NOR U103813 ( .A(n84142), .B(n89901), .Z(n89914) );
  NOR U103814 ( .A(n89912), .B(n89914), .Z(n89904) );
  XOR U103815 ( .A(n84143), .B(n89904), .Z(n88756) );
  XOR U103816 ( .A(n88755), .B(n88756), .Z(n84144) );
  IV U103817 ( .A(n84144), .Z(n88758) );
  XOR U103818 ( .A(n88757), .B(n88758), .Z(n88760) );
  XOR U103819 ( .A(n88761), .B(n88760), .Z(n88748) );
  IV U103820 ( .A(n84145), .Z(n84147) );
  NOR U103821 ( .A(n84147), .B(n84146), .Z(n84151) );
  NOR U103822 ( .A(n84149), .B(n84148), .Z(n84150) );
  NOR U103823 ( .A(n84151), .B(n84150), .Z(n88750) );
  XOR U103824 ( .A(n88748), .B(n88750), .Z(n88751) );
  XOR U103825 ( .A(n88752), .B(n88751), .Z(n89925) );
  XOR U103826 ( .A(n89927), .B(n89925), .Z(n89929) );
  XOR U103827 ( .A(n89928), .B(n89929), .Z(n84152) );
  IV U103828 ( .A(n84152), .Z(n89932) );
  NOR U103829 ( .A(n89935), .B(n89932), .Z(n84159) );
  NOR U103830 ( .A(n84153), .B(n84152), .Z(n84157) );
  IV U103831 ( .A(n84154), .Z(n84155) );
  NOR U103832 ( .A(n84156), .B(n84155), .Z(n89934) );
  XOR U103833 ( .A(n84157), .B(n89934), .Z(n84158) );
  NOR U103834 ( .A(n84159), .B(n84158), .Z(n84160) );
  IV U103835 ( .A(n84160), .Z(n89941) );
  XOR U103836 ( .A(n89940), .B(n89941), .Z(n88742) );
  XOR U103837 ( .A(n88741), .B(n88742), .Z(n88744) );
  IV U103838 ( .A(n84161), .Z(n84163) );
  NOR U103839 ( .A(n84163), .B(n84162), .Z(n84168) );
  IV U103840 ( .A(n84164), .Z(n84165) );
  NOR U103841 ( .A(n84166), .B(n84165), .Z(n84167) );
  NOR U103842 ( .A(n84168), .B(n84167), .Z(n88745) );
  XOR U103843 ( .A(n88744), .B(n88745), .Z(n88738) );
  XOR U103844 ( .A(n88740), .B(n88738), .Z(n88715) );
  XOR U103845 ( .A(n88714), .B(n88715), .Z(n88717) );
  XOR U103846 ( .A(n88718), .B(n88717), .Z(n84169) );
  IV U103847 ( .A(n84169), .Z(n89957) );
  XOR U103848 ( .A(n88708), .B(n89957), .Z(n88710) );
  IV U103849 ( .A(n84170), .Z(n84171) );
  NOR U103850 ( .A(n84172), .B(n84171), .Z(n89955) );
  IV U103851 ( .A(n84173), .Z(n84175) );
  NOR U103852 ( .A(n84175), .B(n84174), .Z(n84176) );
  IV U103853 ( .A(n84176), .Z(n88711) );
  XOR U103854 ( .A(n89955), .B(n88711), .Z(n84177) );
  XOR U103855 ( .A(n88710), .B(n84177), .Z(n84178) );
  IV U103856 ( .A(n84178), .Z(n88727) );
  XOR U103857 ( .A(n88726), .B(n88727), .Z(n88730) );
  XOR U103858 ( .A(n88729), .B(n88730), .Z(n88724) );
  XOR U103859 ( .A(n88723), .B(n88724), .Z(n88701) );
  XOR U103860 ( .A(n88700), .B(n88701), .Z(n88704) );
  XOR U103861 ( .A(n88703), .B(n88704), .Z(n89969) );
  IV U103862 ( .A(n84179), .Z(n84180) );
  NOR U103863 ( .A(n84181), .B(n84180), .Z(n84186) );
  IV U103864 ( .A(n84182), .Z(n84183) );
  NOR U103865 ( .A(n84184), .B(n84183), .Z(n84185) );
  NOR U103866 ( .A(n84186), .B(n84185), .Z(n89970) );
  XOR U103867 ( .A(n89969), .B(n89970), .Z(n89972) );
  XOR U103868 ( .A(n89971), .B(n89972), .Z(n89961) );
  XOR U103869 ( .A(n89963), .B(n89961), .Z(n89987) );
  XOR U103870 ( .A(n84187), .B(n89987), .Z(n89981) );
  IV U103871 ( .A(n84188), .Z(n84191) );
  IV U103872 ( .A(n84189), .Z(n84190) );
  NOR U103873 ( .A(n84191), .B(n84190), .Z(n89979) );
  XOR U103874 ( .A(n89981), .B(n89979), .Z(n89983) );
  XOR U103875 ( .A(n89982), .B(n89983), .Z(n90000) );
  IV U103876 ( .A(n89998), .Z(n90001) );
  XOR U103877 ( .A(n90000), .B(n90001), .Z(n90014) );
  XOR U103878 ( .A(n84195), .B(n90014), .Z(n90009) );
  XOR U103879 ( .A(n90010), .B(n90009), .Z(n90024) );
  XOR U103880 ( .A(n90023), .B(n90024), .Z(n90027) );
  XOR U103881 ( .A(n90026), .B(n90027), .Z(n84201) );
  IV U103882 ( .A(n84196), .Z(n84199) );
  NOR U103883 ( .A(n84197), .B(n84210), .Z(n84198) );
  IV U103884 ( .A(n84198), .Z(n84203) );
  NOR U103885 ( .A(n84199), .B(n84203), .Z(n84207) );
  IV U103886 ( .A(n84207), .Z(n84200) );
  NOR U103887 ( .A(n84201), .B(n84200), .Z(n90022) );
  IV U103888 ( .A(n84202), .Z(n84204) );
  NOR U103889 ( .A(n84204), .B(n84203), .Z(n90019) );
  NOR U103890 ( .A(n90026), .B(n90019), .Z(n84205) );
  XOR U103891 ( .A(n90027), .B(n84205), .Z(n84206) );
  NOR U103892 ( .A(n84207), .B(n84206), .Z(n84208) );
  NOR U103893 ( .A(n90022), .B(n84208), .Z(n88675) );
  IV U103894 ( .A(n84209), .Z(n84213) );
  XOR U103895 ( .A(n84211), .B(n84210), .Z(n84212) );
  NOR U103896 ( .A(n84213), .B(n84212), .Z(n84214) );
  IV U103897 ( .A(n84214), .Z(n88676) );
  XOR U103898 ( .A(n88675), .B(n88676), .Z(n88677) );
  IV U103899 ( .A(n88677), .Z(n84223) );
  IV U103900 ( .A(n84215), .Z(n84217) );
  NOR U103901 ( .A(n84217), .B(n84216), .Z(n84222) );
  IV U103902 ( .A(n84218), .Z(n84219) );
  NOR U103903 ( .A(n84220), .B(n84219), .Z(n84221) );
  NOR U103904 ( .A(n84222), .B(n84221), .Z(n88678) );
  XOR U103905 ( .A(n84223), .B(n88678), .Z(n88673) );
  XOR U103906 ( .A(n84224), .B(n88673), .Z(n88670) );
  IV U103907 ( .A(n84225), .Z(n84227) );
  NOR U103908 ( .A(n84227), .B(n84226), .Z(n84237) );
  IV U103909 ( .A(n84237), .Z(n88671) );
  NOR U103910 ( .A(n88670), .B(n88671), .Z(n84239) );
  IV U103911 ( .A(n84228), .Z(n84230) );
  NOR U103912 ( .A(n84230), .B(n84229), .Z(n84233) );
  IV U103913 ( .A(n84233), .Z(n84232) );
  XOR U103914 ( .A(n88669), .B(n88673), .Z(n84231) );
  NOR U103915 ( .A(n84232), .B(n84231), .Z(n88674) );
  NOR U103916 ( .A(n88670), .B(n84233), .Z(n84234) );
  NOR U103917 ( .A(n88674), .B(n84234), .Z(n84235) );
  IV U103918 ( .A(n84235), .Z(n84236) );
  NOR U103919 ( .A(n84237), .B(n84236), .Z(n84238) );
  NOR U103920 ( .A(n84239), .B(n84238), .Z(n88681) );
  XOR U103921 ( .A(n88679), .B(n88681), .Z(n88682) );
  XOR U103922 ( .A(n88683), .B(n88682), .Z(n88689) );
  XOR U103923 ( .A(n88690), .B(n88689), .Z(n84240) );
  XOR U103924 ( .A(n84241), .B(n84240), .Z(n88661) );
  XOR U103925 ( .A(n88662), .B(n88661), .Z(n88665) );
  XOR U103926 ( .A(n88664), .B(n88665), .Z(n90038) );
  XOR U103927 ( .A(n90037), .B(n90038), .Z(n90041) );
  XOR U103928 ( .A(n90040), .B(n90041), .Z(n90047) );
  IV U103929 ( .A(n84245), .Z(n84242) );
  NOR U103930 ( .A(n84243), .B(n84242), .Z(n90045) );
  IV U103931 ( .A(n84243), .Z(n84244) );
  NOR U103932 ( .A(n84245), .B(n84244), .Z(n84246) );
  NOR U103933 ( .A(n84246), .B(n88655), .Z(n84247) );
  NOR U103934 ( .A(n90045), .B(n84247), .Z(n84248) );
  XOR U103935 ( .A(n90047), .B(n84248), .Z(n88657) );
  IV U103936 ( .A(n84249), .Z(n84250) );
  NOR U103937 ( .A(n84251), .B(n84250), .Z(n88658) );
  IV U103938 ( .A(n84252), .Z(n84253) );
  NOR U103939 ( .A(n84254), .B(n84253), .Z(n90060) );
  NOR U103940 ( .A(n88658), .B(n90060), .Z(n84255) );
  XOR U103941 ( .A(n88657), .B(n84255), .Z(n90059) );
  XOR U103942 ( .A(n90058), .B(n90059), .Z(n84259) );
  IV U103943 ( .A(n84259), .Z(n88647) );
  NOR U103944 ( .A(n84257), .B(n84256), .Z(n84258) );
  IV U103945 ( .A(n84258), .Z(n88644) );
  NOR U103946 ( .A(n88647), .B(n88644), .Z(n84266) );
  NOR U103947 ( .A(n84259), .B(n84258), .Z(n84264) );
  IV U103948 ( .A(n84260), .Z(n84263) );
  IV U103949 ( .A(n84261), .Z(n84262) );
  NOR U103950 ( .A(n84263), .B(n84262), .Z(n88646) );
  XOR U103951 ( .A(n84264), .B(n88646), .Z(n84265) );
  NOR U103952 ( .A(n84266), .B(n84265), .Z(n84267) );
  IV U103953 ( .A(n84267), .Z(n88642) );
  XOR U103954 ( .A(n88641), .B(n88642), .Z(n84268) );
  NOR U103955 ( .A(n84269), .B(n84268), .Z(n88640) );
  IV U103956 ( .A(n84270), .Z(n84272) );
  NOR U103957 ( .A(n84272), .B(n84271), .Z(n88637) );
  NOR U103958 ( .A(n88641), .B(n88637), .Z(n84273) );
  XOR U103959 ( .A(n88642), .B(n84273), .Z(n84274) );
  NOR U103960 ( .A(n84275), .B(n84274), .Z(n84276) );
  NOR U103961 ( .A(n88640), .B(n84276), .Z(n88627) );
  IV U103962 ( .A(n84277), .Z(n84278) );
  NOR U103963 ( .A(n84279), .B(n84278), .Z(n84280) );
  IV U103964 ( .A(n84280), .Z(n88628) );
  XOR U103965 ( .A(n88627), .B(n88628), .Z(n88632) );
  XOR U103966 ( .A(n88630), .B(n88632), .Z(n90076) );
  XOR U103967 ( .A(n90075), .B(n90076), .Z(n90079) );
  XOR U103968 ( .A(n90078), .B(n90079), .Z(n90068) );
  XOR U103969 ( .A(n90067), .B(n90068), .Z(n90071) );
  XOR U103970 ( .A(n90070), .B(n90071), .Z(n88607) );
  XOR U103971 ( .A(n88605), .B(n88607), .Z(n88609) );
  XOR U103972 ( .A(n88608), .B(n88609), .Z(n88635) );
  XOR U103973 ( .A(n88636), .B(n88635), .Z(n90095) );
  XOR U103974 ( .A(n90094), .B(n90095), .Z(n88617) );
  IV U103975 ( .A(n84281), .Z(n84284) );
  NOR U103976 ( .A(n84282), .B(n84289), .Z(n84283) );
  IV U103977 ( .A(n84283), .Z(n84297) );
  NOR U103978 ( .A(n84284), .B(n84297), .Z(n88615) );
  IV U103979 ( .A(n84285), .Z(n84286) );
  NOR U103980 ( .A(n84287), .B(n84286), .Z(n84292) );
  IV U103981 ( .A(n84288), .Z(n84290) );
  NOR U103982 ( .A(n84290), .B(n84289), .Z(n84291) );
  NOR U103983 ( .A(n84292), .B(n84291), .Z(n90097) );
  IV U103984 ( .A(n90097), .Z(n84293) );
  NOR U103985 ( .A(n88615), .B(n84293), .Z(n84294) );
  XOR U103986 ( .A(n88617), .B(n84294), .Z(n84295) );
  IV U103987 ( .A(n84295), .Z(n88621) );
  IV U103988 ( .A(n84296), .Z(n84298) );
  NOR U103989 ( .A(n84298), .B(n84297), .Z(n88619) );
  XOR U103990 ( .A(n88621), .B(n88619), .Z(n90112) );
  IV U103991 ( .A(n84299), .Z(n84301) );
  NOR U103992 ( .A(n84301), .B(n84300), .Z(n90110) );
  NOR U103993 ( .A(n88613), .B(n90110), .Z(n84302) );
  XOR U103994 ( .A(n90112), .B(n84302), .Z(n90107) );
  XOR U103995 ( .A(n90108), .B(n90107), .Z(n90116) );
  XOR U103996 ( .A(n90115), .B(n90116), .Z(n90119) );
  XOR U103997 ( .A(n90118), .B(n90119), .Z(n90125) );
  XOR U103998 ( .A(n90126), .B(n90125), .Z(n90127) );
  IV U103999 ( .A(n84303), .Z(n84305) );
  NOR U104000 ( .A(n84305), .B(n84304), .Z(n84306) );
  IV U104001 ( .A(n84306), .Z(n90128) );
  XOR U104002 ( .A(n90127), .B(n90128), .Z(n90143) );
  XOR U104003 ( .A(n90142), .B(n90143), .Z(n90134) );
  IV U104004 ( .A(n84307), .Z(n84308) );
  NOR U104005 ( .A(n84309), .B(n84308), .Z(n90141) );
  IV U104006 ( .A(n84310), .Z(n84312) );
  NOR U104007 ( .A(n84312), .B(n84311), .Z(n90132) );
  NOR U104008 ( .A(n90141), .B(n90132), .Z(n84313) );
  XOR U104009 ( .A(n90134), .B(n84313), .Z(n90154) );
  XOR U104010 ( .A(n90156), .B(n90154), .Z(n90159) );
  IV U104011 ( .A(n84314), .Z(n84315) );
  NOR U104012 ( .A(n84318), .B(n84315), .Z(n90157) );
  XOR U104013 ( .A(n90159), .B(n90157), .Z(n90149) );
  IV U104014 ( .A(n84316), .Z(n84317) );
  NOR U104015 ( .A(n84318), .B(n84317), .Z(n90147) );
  XOR U104016 ( .A(n90149), .B(n90147), .Z(n90150) );
  IV U104017 ( .A(n84319), .Z(n84320) );
  NOR U104018 ( .A(n84321), .B(n84320), .Z(n84326) );
  IV U104019 ( .A(n84322), .Z(n84324) );
  NOR U104020 ( .A(n84324), .B(n84323), .Z(n84325) );
  NOR U104021 ( .A(n84326), .B(n84325), .Z(n90151) );
  XOR U104022 ( .A(n90150), .B(n90151), .Z(n84327) );
  IV U104023 ( .A(n84327), .Z(n88599) );
  XOR U104024 ( .A(n88597), .B(n88599), .Z(n88602) );
  XOR U104025 ( .A(n88600), .B(n88602), .Z(n88580) );
  XOR U104026 ( .A(n88579), .B(n88580), .Z(n88575) );
  XOR U104027 ( .A(n84328), .B(n88575), .Z(n88570) );
  XOR U104028 ( .A(n88571), .B(n88570), .Z(n88585) );
  XOR U104029 ( .A(n88584), .B(n88585), .Z(n88588) );
  XOR U104030 ( .A(n88587), .B(n88588), .Z(n88596) );
  XOR U104031 ( .A(n88594), .B(n88596), .Z(n88561) );
  XOR U104032 ( .A(n88560), .B(n88561), .Z(n88565) );
  XOR U104033 ( .A(n88563), .B(n88565), .Z(n88553) );
  XOR U104034 ( .A(n88554), .B(n88553), .Z(n88555) );
  XOR U104035 ( .A(n88557), .B(n88555), .Z(n88546) );
  XOR U104036 ( .A(n88545), .B(n88546), .Z(n88549) );
  XOR U104037 ( .A(n88548), .B(n88549), .Z(n90201) );
  XOR U104038 ( .A(n90199), .B(n90201), .Z(n90196) );
  XOR U104039 ( .A(n84329), .B(n90196), .Z(n90187) );
  IV U104040 ( .A(n90187), .Z(n90185) );
  XOR U104041 ( .A(n90188), .B(n90185), .Z(n90181) );
  IV U104042 ( .A(n90181), .Z(n84337) );
  IV U104043 ( .A(n84330), .Z(n84331) );
  NOR U104044 ( .A(n84332), .B(n84331), .Z(n90186) );
  IV U104045 ( .A(n84333), .Z(n84334) );
  NOR U104046 ( .A(n84335), .B(n84334), .Z(n90179) );
  NOR U104047 ( .A(n90186), .B(n90179), .Z(n84336) );
  XOR U104048 ( .A(n84337), .B(n84336), .Z(n90178) );
  XOR U104049 ( .A(n90176), .B(n90178), .Z(n88538) );
  XOR U104050 ( .A(n84338), .B(n88538), .Z(n88542) );
  NOR U104051 ( .A(n84340), .B(n84339), .Z(n88540) );
  XOR U104052 ( .A(n88542), .B(n88540), .Z(n90216) );
  IV U104053 ( .A(n84341), .Z(n84342) );
  NOR U104054 ( .A(n84349), .B(n84342), .Z(n90214) );
  IV U104055 ( .A(n84343), .Z(n84344) );
  NOR U104056 ( .A(n84350), .B(n84344), .Z(n84345) );
  IV U104057 ( .A(n84345), .Z(n84346) );
  NOR U104058 ( .A(n84349), .B(n84346), .Z(n88528) );
  NOR U104059 ( .A(n90214), .B(n88528), .Z(n84347) );
  XOR U104060 ( .A(n90216), .B(n84347), .Z(n90211) );
  IV U104061 ( .A(n84348), .Z(n84353) );
  NOR U104062 ( .A(n84350), .B(n84349), .Z(n84351) );
  IV U104063 ( .A(n84351), .Z(n84352) );
  NOR U104064 ( .A(n84353), .B(n84352), .Z(n84354) );
  IV U104065 ( .A(n84354), .Z(n90212) );
  XOR U104066 ( .A(n90211), .B(n90212), .Z(n90209) );
  XOR U104067 ( .A(n90208), .B(n90209), .Z(n88519) );
  XOR U104068 ( .A(n88518), .B(n88519), .Z(n88522) );
  XOR U104069 ( .A(n88521), .B(n88522), .Z(n88512) );
  XOR U104070 ( .A(n88511), .B(n88512), .Z(n88514) );
  XOR U104071 ( .A(n88515), .B(n88514), .Z(n88532) );
  XOR U104072 ( .A(n88531), .B(n88532), .Z(n88504) );
  IV U104073 ( .A(n84355), .Z(n84356) );
  NOR U104074 ( .A(n84357), .B(n84356), .Z(n88503) );
  IV U104075 ( .A(n84358), .Z(n84361) );
  IV U104076 ( .A(n84359), .Z(n84360) );
  NOR U104077 ( .A(n84361), .B(n84360), .Z(n84362) );
  IV U104078 ( .A(n84362), .Z(n88534) );
  XOR U104079 ( .A(n88503), .B(n88534), .Z(n84363) );
  XOR U104080 ( .A(n88504), .B(n84363), .Z(n84364) );
  IV U104081 ( .A(n84364), .Z(n88497) );
  XOR U104082 ( .A(n88495), .B(n88497), .Z(n88499) );
  XOR U104083 ( .A(n88498), .B(n88499), .Z(n88466) );
  XOR U104084 ( .A(n84365), .B(n88466), .Z(n84379) );
  IV U104085 ( .A(n84379), .Z(n84366) );
  NOR U104086 ( .A(n84378), .B(n84366), .Z(n84374) );
  XOR U104087 ( .A(n84367), .B(n88466), .Z(n84372) );
  IV U104088 ( .A(n84368), .Z(n84369) );
  NOR U104089 ( .A(n84370), .B(n84369), .Z(n84375) );
  IV U104090 ( .A(n84375), .Z(n84371) );
  NOR U104091 ( .A(n84372), .B(n84371), .Z(n84373) );
  NOR U104092 ( .A(n84374), .B(n84373), .Z(n88472) );
  IV U104093 ( .A(n88472), .Z(n84377) );
  NOR U104094 ( .A(n84375), .B(n84379), .Z(n84376) );
  NOR U104095 ( .A(n84377), .B(n84376), .Z(n84381) );
  NOR U104096 ( .A(n84379), .B(n84378), .Z(n84380) );
  NOR U104097 ( .A(n84381), .B(n84380), .Z(n88474) );
  XOR U104098 ( .A(n88473), .B(n88474), .Z(n88482) );
  IV U104099 ( .A(n88482), .Z(n84390) );
  IV U104100 ( .A(n84382), .Z(n84384) );
  NOR U104101 ( .A(n84384), .B(n84383), .Z(n84394) );
  IV U104102 ( .A(n84394), .Z(n88483) );
  NOR U104103 ( .A(n84390), .B(n88483), .Z(n84396) );
  IV U104104 ( .A(n84385), .Z(n84387) );
  NOR U104105 ( .A(n84387), .B(n84386), .Z(n84389) );
  IV U104106 ( .A(n84389), .Z(n84388) );
  NOR U104107 ( .A(n88474), .B(n84388), .Z(n88475) );
  NOR U104108 ( .A(n84390), .B(n84389), .Z(n84391) );
  NOR U104109 ( .A(n88475), .B(n84391), .Z(n84392) );
  IV U104110 ( .A(n84392), .Z(n84393) );
  NOR U104111 ( .A(n84394), .B(n84393), .Z(n84395) );
  NOR U104112 ( .A(n84396), .B(n84395), .Z(n88485) );
  XOR U104113 ( .A(n88484), .B(n88485), .Z(n88488) );
  IV U104114 ( .A(n88488), .Z(n84397) );
  NOR U104115 ( .A(n88487), .B(n84397), .Z(n84401) );
  IV U104116 ( .A(n84398), .Z(n84399) );
  NOR U104117 ( .A(n84399), .B(n84403), .Z(n84407) );
  IV U104118 ( .A(n84407), .Z(n84400) );
  NOR U104119 ( .A(n84401), .B(n84400), .Z(n88494) );
  IV U104120 ( .A(n84402), .Z(n84404) );
  NOR U104121 ( .A(n84404), .B(n84403), .Z(n84405) );
  IV U104122 ( .A(n84405), .Z(n88491) );
  XOR U104123 ( .A(n88487), .B(n88488), .Z(n88490) );
  XOR U104124 ( .A(n88491), .B(n88490), .Z(n84406) );
  NOR U104125 ( .A(n84407), .B(n84406), .Z(n84408) );
  NOR U104126 ( .A(n88494), .B(n84408), .Z(n88476) );
  IV U104127 ( .A(n84409), .Z(n84411) );
  NOR U104128 ( .A(n84411), .B(n84410), .Z(n88479) );
  IV U104129 ( .A(n84412), .Z(n84413) );
  NOR U104130 ( .A(n84414), .B(n84413), .Z(n88477) );
  NOR U104131 ( .A(n88479), .B(n88477), .Z(n84415) );
  XOR U104132 ( .A(n88476), .B(n84415), .Z(n88446) );
  XOR U104133 ( .A(n88444), .B(n88446), .Z(n88447) );
  XOR U104134 ( .A(n88448), .B(n88447), .Z(n88453) );
  XOR U104135 ( .A(n88455), .B(n88453), .Z(n88457) );
  XOR U104136 ( .A(n88456), .B(n88457), .Z(n88438) );
  IV U104137 ( .A(n84416), .Z(n84418) );
  NOR U104138 ( .A(n84418), .B(n84417), .Z(n88436) );
  XOR U104139 ( .A(n88438), .B(n88436), .Z(n88440) );
  XOR U104140 ( .A(n88439), .B(n88440), .Z(n88463) );
  XOR U104141 ( .A(n88464), .B(n88463), .Z(n90241) );
  XOR U104142 ( .A(n90243), .B(n90241), .Z(n90244) );
  XOR U104143 ( .A(n90245), .B(n90244), .Z(n84419) );
  IV U104144 ( .A(n84419), .Z(n88435) );
  NOR U104145 ( .A(n84427), .B(n88435), .Z(n90296) );
  IV U104146 ( .A(n84420), .Z(n84426) );
  IV U104147 ( .A(n84421), .Z(n84423) );
  NOR U104148 ( .A(n84423), .B(n84422), .Z(n84424) );
  IV U104149 ( .A(n84424), .Z(n84425) );
  NOR U104150 ( .A(n84426), .B(n84425), .Z(n84428) );
  IV U104151 ( .A(n84428), .Z(n88434) );
  XOR U104152 ( .A(n88435), .B(n88434), .Z(n84430) );
  NOR U104153 ( .A(n84428), .B(n84427), .Z(n84429) );
  NOR U104154 ( .A(n84430), .B(n84429), .Z(n90293) );
  NOR U104155 ( .A(n90296), .B(n90293), .Z(n88429) );
  IV U104156 ( .A(n84431), .Z(n84432) );
  NOR U104157 ( .A(n84433), .B(n84432), .Z(n90292) );
  IV U104158 ( .A(n84434), .Z(n84436) );
  NOR U104159 ( .A(n84436), .B(n84435), .Z(n88428) );
  NOR U104160 ( .A(n90292), .B(n88428), .Z(n84437) );
  XOR U104161 ( .A(n88429), .B(n84437), .Z(n88427) );
  XOR U104162 ( .A(n88425), .B(n88427), .Z(n90283) );
  XOR U104163 ( .A(n90284), .B(n90283), .Z(n90280) );
  IV U104164 ( .A(n90280), .Z(n90285) );
  IV U104165 ( .A(n84438), .Z(n84440) );
  NOR U104166 ( .A(n84440), .B(n84439), .Z(n84445) );
  IV U104167 ( .A(n84441), .Z(n84443) );
  NOR U104168 ( .A(n84443), .B(n84442), .Z(n84444) );
  NOR U104169 ( .A(n84445), .B(n84444), .Z(n90286) );
  XOR U104170 ( .A(n90285), .B(n90286), .Z(n84446) );
  XOR U104171 ( .A(n84447), .B(n84446), .Z(n90254) );
  IV U104172 ( .A(n84448), .Z(n84450) );
  NOR U104173 ( .A(n84450), .B(n84449), .Z(n90256) );
  XOR U104174 ( .A(n90254), .B(n90256), .Z(n90267) );
  IV U104175 ( .A(n84451), .Z(n84453) );
  NOR U104176 ( .A(n84453), .B(n84452), .Z(n90266) );
  NOR U104177 ( .A(n90266), .B(n90260), .Z(n84458) );
  XOR U104178 ( .A(n90267), .B(n84458), .Z(n90263) );
  XOR U104179 ( .A(n84459), .B(n90263), .Z(n88417) );
  XOR U104180 ( .A(n88416), .B(n88417), .Z(n88419) );
  XOR U104181 ( .A(n88420), .B(n88419), .Z(n84460) );
  IV U104182 ( .A(n84460), .Z(n88423) );
  NOR U104183 ( .A(n84461), .B(n88423), .Z(n88414) );
  NOR U104184 ( .A(n84463), .B(n84462), .Z(n84464) );
  IV U104185 ( .A(n84464), .Z(n88424) );
  XOR U104186 ( .A(n88424), .B(n88423), .Z(n84465) );
  NOR U104187 ( .A(n84466), .B(n84465), .Z(n88412) );
  IV U104188 ( .A(n84467), .Z(n84469) );
  NOR U104189 ( .A(n84469), .B(n84468), .Z(n88411) );
  XOR U104190 ( .A(n88412), .B(n88411), .Z(n84470) );
  NOR U104191 ( .A(n88414), .B(n84470), .Z(n90313) );
  XOR U104192 ( .A(n90312), .B(n90313), .Z(n84471) );
  XOR U104193 ( .A(n90311), .B(n84471), .Z(n88405) );
  IV U104194 ( .A(n84472), .Z(n84474) );
  NOR U104195 ( .A(n84474), .B(n84473), .Z(n88403) );
  XOR U104196 ( .A(n88405), .B(n88403), .Z(n88407) );
  XOR U104197 ( .A(n88406), .B(n88407), .Z(n88398) );
  XOR U104198 ( .A(n88396), .B(n88398), .Z(n90330) );
  XOR U104199 ( .A(n84475), .B(n90330), .Z(n90322) );
  IV U104200 ( .A(n84476), .Z(n84478) );
  NOR U104201 ( .A(n84478), .B(n84477), .Z(n84488) );
  IV U104202 ( .A(n84488), .Z(n90324) );
  NOR U104203 ( .A(n90322), .B(n90324), .Z(n84490) );
  IV U104204 ( .A(n84479), .Z(n84481) );
  NOR U104205 ( .A(n84481), .B(n84480), .Z(n84484) );
  IV U104206 ( .A(n84484), .Z(n84483) );
  XOR U104207 ( .A(n88399), .B(n90330), .Z(n84482) );
  NOR U104208 ( .A(n84483), .B(n84482), .Z(n90333) );
  NOR U104209 ( .A(n90322), .B(n84484), .Z(n84485) );
  NOR U104210 ( .A(n90333), .B(n84485), .Z(n84486) );
  IV U104211 ( .A(n84486), .Z(n84487) );
  NOR U104212 ( .A(n84488), .B(n84487), .Z(n84489) );
  NOR U104213 ( .A(n84490), .B(n84489), .Z(n90325) );
  XOR U104214 ( .A(n90326), .B(n90325), .Z(n84491) );
  IV U104215 ( .A(n84491), .Z(n88394) );
  XOR U104216 ( .A(n88393), .B(n88394), .Z(n88382) );
  NOR U104217 ( .A(n84493), .B(n84492), .Z(n88392) );
  IV U104218 ( .A(n84494), .Z(n84496) );
  NOR U104219 ( .A(n84496), .B(n84495), .Z(n88380) );
  NOR U104220 ( .A(n88392), .B(n88380), .Z(n84497) );
  XOR U104221 ( .A(n88382), .B(n84497), .Z(n84498) );
  IV U104222 ( .A(n84498), .Z(n88387) );
  XOR U104223 ( .A(n88385), .B(n88387), .Z(n88388) );
  XOR U104224 ( .A(n88389), .B(n88388), .Z(n88377) );
  XOR U104225 ( .A(n88379), .B(n88377), .Z(n88366) );
  XOR U104226 ( .A(n88365), .B(n88366), .Z(n88369) );
  XOR U104227 ( .A(n88368), .B(n88369), .Z(n88373) );
  XOR U104228 ( .A(n88374), .B(n88373), .Z(n84499) );
  IV U104229 ( .A(n84499), .Z(n88358) );
  XOR U104230 ( .A(n88357), .B(n88358), .Z(n88361) );
  XOR U104231 ( .A(n88360), .B(n88361), .Z(n88321) );
  XOR U104232 ( .A(n88320), .B(n88321), .Z(n88324) );
  XOR U104233 ( .A(n88323), .B(n88324), .Z(n88314) );
  XOR U104234 ( .A(n88313), .B(n88314), .Z(n88316) );
  XOR U104235 ( .A(n88317), .B(n88316), .Z(n84503) );
  XOR U104236 ( .A(n84500), .B(n84503), .Z(n88330) );
  XOR U104237 ( .A(n88331), .B(n88330), .Z(n84501) );
  NOR U104238 ( .A(n84502), .B(n84501), .Z(n88349) );
  IV U104239 ( .A(n84502), .Z(n84505) );
  IV U104240 ( .A(n84503), .Z(n88334) );
  XOR U104241 ( .A(n88333), .B(n88334), .Z(n84504) );
  NOR U104242 ( .A(n84505), .B(n84504), .Z(n88352) );
  NOR U104243 ( .A(n88349), .B(n88352), .Z(n88343) );
  XOR U104244 ( .A(n84506), .B(n88343), .Z(n88341) );
  XOR U104245 ( .A(n88339), .B(n88341), .Z(n88297) );
  IV U104246 ( .A(n84507), .Z(n84508) );
  NOR U104247 ( .A(n84509), .B(n84508), .Z(n84514) );
  IV U104248 ( .A(n84510), .Z(n84511) );
  NOR U104249 ( .A(n84512), .B(n84511), .Z(n84513) );
  NOR U104250 ( .A(n84514), .B(n84513), .Z(n88298) );
  XOR U104251 ( .A(n88297), .B(n88298), .Z(n88299) );
  XOR U104252 ( .A(n88301), .B(n88299), .Z(n88305) );
  XOR U104253 ( .A(n88306), .B(n88305), .Z(n88280) );
  XOR U104254 ( .A(n84515), .B(n88280), .Z(n84516) );
  IV U104255 ( .A(n84516), .Z(n88278) );
  XOR U104256 ( .A(n88277), .B(n88278), .Z(n84517) );
  NOR U104257 ( .A(n84521), .B(n84517), .Z(n84525) );
  IV U104258 ( .A(n84518), .Z(n84520) );
  NOR U104259 ( .A(n84520), .B(n84519), .Z(n84527) );
  IV U104260 ( .A(n84521), .Z(n84522) );
  NOR U104261 ( .A(n84522), .B(n88278), .Z(n84523) );
  NOR U104262 ( .A(n84527), .B(n84523), .Z(n84524) );
  NOR U104263 ( .A(n84525), .B(n84524), .Z(n88286) );
  IV U104264 ( .A(n84525), .Z(n84526) );
  NOR U104265 ( .A(n84527), .B(n84526), .Z(n84528) );
  NOR U104266 ( .A(n88286), .B(n84528), .Z(n84529) );
  IV U104267 ( .A(n84529), .Z(n88288) );
  XOR U104268 ( .A(n88287), .B(n88288), .Z(n88284) );
  XOR U104269 ( .A(n88285), .B(n88284), .Z(n84538) );
  IV U104270 ( .A(n84538), .Z(n84533) );
  IV U104271 ( .A(n84530), .Z(n84531) );
  NOR U104272 ( .A(n84549), .B(n84531), .Z(n84542) );
  IV U104273 ( .A(n84542), .Z(n84532) );
  NOR U104274 ( .A(n84533), .B(n84532), .Z(n88276) );
  IV U104275 ( .A(n84534), .Z(n84535) );
  NOR U104276 ( .A(n84536), .B(n84535), .Z(n84539) );
  IV U104277 ( .A(n84539), .Z(n84537) );
  NOR U104278 ( .A(n84537), .B(n88288), .Z(n88275) );
  NOR U104279 ( .A(n84539), .B(n84538), .Z(n84540) );
  NOR U104280 ( .A(n88275), .B(n84540), .Z(n84541) );
  NOR U104281 ( .A(n84542), .B(n84541), .Z(n84543) );
  NOR U104282 ( .A(n88276), .B(n84543), .Z(n90366) );
  IV U104283 ( .A(n84544), .Z(n84546) );
  NOR U104284 ( .A(n84546), .B(n84545), .Z(n90370) );
  IV U104285 ( .A(n84547), .Z(n84548) );
  NOR U104286 ( .A(n84549), .B(n84548), .Z(n90365) );
  NOR U104287 ( .A(n90370), .B(n90365), .Z(n84550) );
  XOR U104288 ( .A(n90366), .B(n84550), .Z(n90377) );
  IV U104289 ( .A(n84551), .Z(n84552) );
  NOR U104290 ( .A(n84553), .B(n84552), .Z(n90373) );
  IV U104291 ( .A(n84554), .Z(n84555) );
  NOR U104292 ( .A(n84556), .B(n84555), .Z(n90376) );
  NOR U104293 ( .A(n90373), .B(n90376), .Z(n84557) );
  XOR U104294 ( .A(n90377), .B(n84557), .Z(n90358) );
  IV U104295 ( .A(n90358), .Z(n90356) );
  XOR U104296 ( .A(n90357), .B(n90356), .Z(n90401) );
  IV U104297 ( .A(n84558), .Z(n84559) );
  NOR U104298 ( .A(n84560), .B(n84559), .Z(n90400) );
  NOR U104299 ( .A(n90360), .B(n90400), .Z(n84561) );
  XOR U104300 ( .A(n90401), .B(n84561), .Z(n90399) );
  IV U104301 ( .A(n84562), .Z(n84564) );
  NOR U104302 ( .A(n84564), .B(n84563), .Z(n84565) );
  IV U104303 ( .A(n84565), .Z(n90398) );
  XOR U104304 ( .A(n90399), .B(n90398), .Z(n90416) );
  XOR U104305 ( .A(n90412), .B(n90416), .Z(n90388) );
  IV U104306 ( .A(n84566), .Z(n84567) );
  NOR U104307 ( .A(n84568), .B(n84567), .Z(n90414) );
  IV U104308 ( .A(n84569), .Z(n84571) );
  NOR U104309 ( .A(n84571), .B(n84570), .Z(n90387) );
  NOR U104310 ( .A(n90414), .B(n90387), .Z(n84572) );
  XOR U104311 ( .A(n90388), .B(n84572), .Z(n90390) );
  NOR U104312 ( .A(n84573), .B(n90393), .Z(n84577) );
  NOR U104313 ( .A(n84575), .B(n84574), .Z(n84576) );
  NOR U104314 ( .A(n84577), .B(n84576), .Z(n90427) );
  IV U104315 ( .A(n90427), .Z(n84578) );
  NOR U104316 ( .A(n90429), .B(n84578), .Z(n84579) );
  XOR U104317 ( .A(n90390), .B(n84579), .Z(n88268) );
  XOR U104318 ( .A(n88269), .B(n88268), .Z(n88270) );
  XOR U104319 ( .A(n88272), .B(n88270), .Z(n90462) );
  XOR U104320 ( .A(n90461), .B(n90462), .Z(n90464) );
  XOR U104321 ( .A(n90465), .B(n90464), .Z(n84580) );
  IV U104322 ( .A(n84580), .Z(n90449) );
  XOR U104323 ( .A(n90448), .B(n90449), .Z(n90452) );
  XOR U104324 ( .A(n90451), .B(n90452), .Z(n90446) );
  XOR U104325 ( .A(n90445), .B(n90446), .Z(n90440) );
  IV U104326 ( .A(n84581), .Z(n84583) );
  NOR U104327 ( .A(n84583), .B(n84582), .Z(n90438) );
  XOR U104328 ( .A(n90440), .B(n90438), .Z(n88264) );
  IV U104329 ( .A(n84584), .Z(n84592) );
  IV U104330 ( .A(n84591), .Z(n84585) );
  NOR U104331 ( .A(n84592), .B(n84585), .Z(n90442) );
  IV U104332 ( .A(n84586), .Z(n84587) );
  NOR U104333 ( .A(n84592), .B(n84587), .Z(n88263) );
  NOR U104334 ( .A(n90442), .B(n88263), .Z(n84588) );
  XOR U104335 ( .A(n88264), .B(n84588), .Z(n84589) );
  IV U104336 ( .A(n84589), .Z(n88255) );
  IV U104337 ( .A(n84590), .Z(n84594) );
  XOR U104338 ( .A(n84592), .B(n84591), .Z(n84593) );
  NOR U104339 ( .A(n84594), .B(n84593), .Z(n88253) );
  XOR U104340 ( .A(n88255), .B(n88253), .Z(n88258) );
  XOR U104341 ( .A(n88256), .B(n88258), .Z(n88259) );
  XOR U104342 ( .A(n88260), .B(n88259), .Z(n84595) );
  IV U104343 ( .A(n84595), .Z(n90480) );
  NOR U104344 ( .A(n90483), .B(n90480), .Z(n84599) );
  NOR U104345 ( .A(n84596), .B(n84595), .Z(n84597) );
  XOR U104346 ( .A(n84597), .B(n90482), .Z(n84598) );
  NOR U104347 ( .A(n84599), .B(n84598), .Z(n88250) );
  XOR U104348 ( .A(n90479), .B(n88250), .Z(n88242) );
  IV U104349 ( .A(n84600), .Z(n84602) );
  NOR U104350 ( .A(n84602), .B(n84601), .Z(n88240) );
  NOR U104351 ( .A(n88251), .B(n88240), .Z(n84603) );
  XOR U104352 ( .A(n88242), .B(n84603), .Z(n84604) );
  IV U104353 ( .A(n84604), .Z(n88236) );
  XOR U104354 ( .A(n88234), .B(n88236), .Z(n88243) );
  IV U104355 ( .A(n84605), .Z(n84606) );
  NOR U104356 ( .A(n84607), .B(n84606), .Z(n84612) );
  IV U104357 ( .A(n84608), .Z(n84609) );
  NOR U104358 ( .A(n84610), .B(n84609), .Z(n84611) );
  NOR U104359 ( .A(n84612), .B(n84611), .Z(n88244) );
  XOR U104360 ( .A(n88243), .B(n88244), .Z(n84613) );
  IV U104361 ( .A(n84613), .Z(n88238) );
  XOR U104362 ( .A(n88237), .B(n88238), .Z(n88246) );
  XOR U104363 ( .A(n88245), .B(n88246), .Z(n88217) );
  XOR U104364 ( .A(n88216), .B(n88217), .Z(n88219) );
  XOR U104365 ( .A(n88218), .B(n88219), .Z(n88213) );
  XOR U104366 ( .A(n88212), .B(n88213), .Z(n88215) );
  XOR U104367 ( .A(n88214), .B(n88215), .Z(n88222) );
  XOR U104368 ( .A(n88221), .B(n88222), .Z(n88224) );
  XOR U104369 ( .A(n84614), .B(n88224), .Z(n88229) );
  IV U104370 ( .A(n84615), .Z(n84617) );
  NOR U104371 ( .A(n84617), .B(n84616), .Z(n84627) );
  IV U104372 ( .A(n84627), .Z(n88230) );
  NOR U104373 ( .A(n88229), .B(n88230), .Z(n84629) );
  IV U104374 ( .A(n84618), .Z(n84619) );
  NOR U104375 ( .A(n84620), .B(n84619), .Z(n84623) );
  IV U104376 ( .A(n84623), .Z(n84622) );
  XOR U104377 ( .A(n88223), .B(n88224), .Z(n84621) );
  NOR U104378 ( .A(n84622), .B(n84621), .Z(n88231) );
  NOR U104379 ( .A(n88229), .B(n84623), .Z(n84624) );
  NOR U104380 ( .A(n88231), .B(n84624), .Z(n84625) );
  IV U104381 ( .A(n84625), .Z(n84626) );
  NOR U104382 ( .A(n84627), .B(n84626), .Z(n84628) );
  NOR U104383 ( .A(n84629), .B(n84628), .Z(n88228) );
  IV U104384 ( .A(n84630), .Z(n84632) );
  NOR U104385 ( .A(n84632), .B(n84631), .Z(n88226) );
  NOR U104386 ( .A(n88227), .B(n88226), .Z(n84633) );
  XOR U104387 ( .A(n88228), .B(n84633), .Z(n84641) );
  IV U104388 ( .A(n84641), .Z(n84634) );
  NOR U104389 ( .A(n84635), .B(n84634), .Z(n88201) );
  IV U104390 ( .A(n84636), .Z(n84638) );
  NOR U104391 ( .A(n84638), .B(n84637), .Z(n84642) );
  IV U104392 ( .A(n84642), .Z(n84640) );
  XOR U104393 ( .A(n88227), .B(n88228), .Z(n84639) );
  NOR U104394 ( .A(n84640), .B(n84639), .Z(n88202) );
  NOR U104395 ( .A(n84642), .B(n84641), .Z(n84643) );
  NOR U104396 ( .A(n88202), .B(n84643), .Z(n90515) );
  NOR U104397 ( .A(n84644), .B(n90515), .Z(n84645) );
  NOR U104398 ( .A(n88201), .B(n84645), .Z(n90510) );
  XOR U104399 ( .A(n84646), .B(n90510), .Z(n90508) );
  XOR U104400 ( .A(n90506), .B(n90508), .Z(n88204) );
  XOR U104401 ( .A(n88206), .B(n88204), .Z(n90540) );
  IV U104402 ( .A(n84647), .Z(n84648) );
  NOR U104403 ( .A(n84649), .B(n84648), .Z(n88207) );
  IV U104404 ( .A(n84650), .Z(n84652) );
  NOR U104405 ( .A(n84652), .B(n84651), .Z(n90538) );
  NOR U104406 ( .A(n88207), .B(n90538), .Z(n84653) );
  XOR U104407 ( .A(n90540), .B(n84653), .Z(n90534) );
  XOR U104408 ( .A(n90535), .B(n90534), .Z(n90528) );
  IV U104409 ( .A(n84654), .Z(n84659) );
  IV U104410 ( .A(n84655), .Z(n84656) );
  NOR U104411 ( .A(n84657), .B(n84656), .Z(n84658) );
  IV U104412 ( .A(n84658), .Z(n84661) );
  NOR U104413 ( .A(n84659), .B(n84661), .Z(n90529) );
  IV U104414 ( .A(n84660), .Z(n84662) );
  NOR U104415 ( .A(n84662), .B(n84661), .Z(n84663) );
  NOR U104416 ( .A(n84664), .B(n84663), .Z(n90526) );
  XOR U104417 ( .A(n90529), .B(n90526), .Z(n84665) );
  XOR U104418 ( .A(n90528), .B(n84665), .Z(n88187) );
  XOR U104419 ( .A(n88186), .B(n88187), .Z(n88195) );
  XOR U104420 ( .A(n84666), .B(n88195), .Z(n84673) );
  NOR U104421 ( .A(n84672), .B(n84673), .Z(n84667) );
  IV U104422 ( .A(n84667), .Z(n84671) );
  IV U104423 ( .A(n84668), .Z(n84669) );
  NOR U104424 ( .A(n84670), .B(n84669), .Z(n84676) );
  NOR U104425 ( .A(n84671), .B(n84676), .Z(n84682) );
  IV U104426 ( .A(n84672), .Z(n84677) );
  XOR U104427 ( .A(n84676), .B(n84677), .Z(n84675) );
  IV U104428 ( .A(n84673), .Z(n84674) );
  NOR U104429 ( .A(n84675), .B(n84674), .Z(n84680) );
  IV U104430 ( .A(n84676), .Z(n84678) );
  NOR U104431 ( .A(n84678), .B(n84677), .Z(n84679) );
  NOR U104432 ( .A(n84680), .B(n84679), .Z(n90558) );
  IV U104433 ( .A(n90558), .Z(n84681) );
  NOR U104434 ( .A(n84682), .B(n84681), .Z(n90549) );
  XOR U104435 ( .A(n90551), .B(n90549), .Z(n90553) );
  XOR U104436 ( .A(n90552), .B(n90553), .Z(n88178) );
  XOR U104437 ( .A(n88176), .B(n88178), .Z(n88180) );
  XOR U104438 ( .A(n88179), .B(n88180), .Z(n88169) );
  XOR U104439 ( .A(n84683), .B(n88169), .Z(n88173) );
  IV U104440 ( .A(n84684), .Z(n84686) );
  NOR U104441 ( .A(n84686), .B(n84685), .Z(n88171) );
  XOR U104442 ( .A(n88173), .B(n88171), .Z(n88163) );
  XOR U104443 ( .A(n88162), .B(n88163), .Z(n88165) );
  IV U104444 ( .A(n84687), .Z(n84688) );
  NOR U104445 ( .A(n84689), .B(n84688), .Z(n84694) );
  IV U104446 ( .A(n84690), .Z(n84692) );
  NOR U104447 ( .A(n84692), .B(n84691), .Z(n84693) );
  NOR U104448 ( .A(n84694), .B(n84693), .Z(n88166) );
  XOR U104449 ( .A(n88165), .B(n88166), .Z(n90574) );
  XOR U104450 ( .A(n90576), .B(n90574), .Z(n90578) );
  NOR U104451 ( .A(n84696), .B(n84695), .Z(n84698) );
  NOR U104452 ( .A(n84698), .B(n84697), .Z(n90577) );
  XOR U104453 ( .A(n90578), .B(n90577), .Z(n90564) );
  IV U104454 ( .A(n90564), .Z(n90566) );
  IV U104455 ( .A(n84699), .Z(n84701) );
  NOR U104456 ( .A(n84701), .B(n84700), .Z(n90565) );
  XOR U104457 ( .A(n90566), .B(n90565), .Z(n84708) );
  IV U104458 ( .A(n84702), .Z(n84704) );
  NOR U104459 ( .A(n84704), .B(n84703), .Z(n90567) );
  NOR U104460 ( .A(n84706), .B(n84705), .Z(n90568) );
  NOR U104461 ( .A(n90567), .B(n90568), .Z(n84707) );
  XOR U104462 ( .A(n84708), .B(n84707), .Z(n90604) );
  XOR U104463 ( .A(n90605), .B(n90604), .Z(n90606) );
  XOR U104464 ( .A(n90608), .B(n90606), .Z(n90596) );
  XOR U104465 ( .A(n90595), .B(n90596), .Z(n90598) );
  IV U104466 ( .A(n84709), .Z(n84711) );
  NOR U104467 ( .A(n84711), .B(n84710), .Z(n84716) );
  IV U104468 ( .A(n84712), .Z(n84714) );
  NOR U104469 ( .A(n84714), .B(n84713), .Z(n84715) );
  NOR U104470 ( .A(n84716), .B(n84715), .Z(n90599) );
  XOR U104471 ( .A(n90598), .B(n90599), .Z(n84717) );
  IV U104472 ( .A(n84717), .Z(n90589) );
  XOR U104473 ( .A(n90588), .B(n90589), .Z(n90591) );
  XOR U104474 ( .A(n90592), .B(n90591), .Z(n88119) );
  IV U104475 ( .A(n88119), .Z(n88122) );
  IV U104476 ( .A(n84718), .Z(n84719) );
  NOR U104477 ( .A(n84720), .B(n84719), .Z(n88124) );
  IV U104478 ( .A(n84721), .Z(n84723) );
  NOR U104479 ( .A(n84723), .B(n84722), .Z(n88120) );
  XOR U104480 ( .A(n88124), .B(n88120), .Z(n84724) );
  XOR U104481 ( .A(n88122), .B(n84724), .Z(n88106) );
  XOR U104482 ( .A(n84725), .B(n88106), .Z(n88109) );
  IV U104483 ( .A(n88109), .Z(n88108) );
  XOR U104484 ( .A(n88110), .B(n88108), .Z(n88138) );
  XOR U104485 ( .A(n88137), .B(n88138), .Z(n90622) );
  IV U104486 ( .A(n84726), .Z(n84727) );
  NOR U104487 ( .A(n84728), .B(n84727), .Z(n88134) );
  IV U104488 ( .A(n84729), .Z(n84731) );
  NOR U104489 ( .A(n84731), .B(n84730), .Z(n90620) );
  NOR U104490 ( .A(n88134), .B(n90620), .Z(n84732) );
  XOR U104491 ( .A(n90622), .B(n84732), .Z(n90617) );
  IV U104492 ( .A(n84733), .Z(n84735) );
  NOR U104493 ( .A(n84735), .B(n84734), .Z(n84739) );
  IV U104494 ( .A(n84736), .Z(n84737) );
  NOR U104495 ( .A(n84737), .B(n84741), .Z(n84738) );
  NOR U104496 ( .A(n84739), .B(n84738), .Z(n90618) );
  XOR U104497 ( .A(n90617), .B(n90618), .Z(n88150) );
  IV U104498 ( .A(n84740), .Z(n84742) );
  NOR U104499 ( .A(n84742), .B(n84741), .Z(n88148) );
  XOR U104500 ( .A(n88150), .B(n88148), .Z(n88147) );
  IV U104501 ( .A(n84743), .Z(n84745) );
  NOR U104502 ( .A(n84745), .B(n84744), .Z(n88145) );
  XOR U104503 ( .A(n88147), .B(n88145), .Z(n88152) );
  IV U104504 ( .A(n88152), .Z(n84746) );
  NOR U104505 ( .A(n84747), .B(n84746), .Z(n90635) );
  IV U104506 ( .A(n84747), .Z(n84748) );
  NOR U104507 ( .A(n84748), .B(n88147), .Z(n90632) );
  NOR U104508 ( .A(n90635), .B(n90632), .Z(n84756) );
  IV U104509 ( .A(n84749), .Z(n84751) );
  NOR U104510 ( .A(n84751), .B(n84750), .Z(n88151) );
  IV U104511 ( .A(n84752), .Z(n84754) );
  NOR U104512 ( .A(n84754), .B(n84753), .Z(n90633) );
  NOR U104513 ( .A(n88151), .B(n90633), .Z(n84755) );
  XOR U104514 ( .A(n84756), .B(n84755), .Z(n84758) );
  NOR U104515 ( .A(n84757), .B(n84758), .Z(n90631) );
  IV U104516 ( .A(n84758), .Z(n84759) );
  NOR U104517 ( .A(n84760), .B(n84759), .Z(n90628) );
  IV U104518 ( .A(n84761), .Z(n84763) );
  NOR U104519 ( .A(n84763), .B(n84762), .Z(n90627) );
  XOR U104520 ( .A(n90628), .B(n90627), .Z(n84764) );
  NOR U104521 ( .A(n90631), .B(n84764), .Z(n90642) );
  IV U104522 ( .A(n84765), .Z(n84767) );
  NOR U104523 ( .A(n84767), .B(n84766), .Z(n90641) );
  IV U104524 ( .A(n90641), .Z(n90638) );
  XOR U104525 ( .A(n90642), .B(n90638), .Z(n88100) );
  IV U104526 ( .A(n84768), .Z(n84770) );
  NOR U104527 ( .A(n84770), .B(n84769), .Z(n90640) );
  IV U104528 ( .A(n84771), .Z(n84774) );
  NOR U104529 ( .A(n84772), .B(n84785), .Z(n84773) );
  IV U104530 ( .A(n84773), .Z(n84777) );
  NOR U104531 ( .A(n84774), .B(n84777), .Z(n88099) );
  NOR U104532 ( .A(n90640), .B(n88099), .Z(n84775) );
  XOR U104533 ( .A(n88100), .B(n84775), .Z(n88085) );
  IV U104534 ( .A(n84776), .Z(n84778) );
  NOR U104535 ( .A(n84778), .B(n84777), .Z(n84779) );
  IV U104536 ( .A(n84779), .Z(n88086) );
  XOR U104537 ( .A(n88085), .B(n88086), .Z(n88097) );
  IV U104538 ( .A(n84780), .Z(n84781) );
  NOR U104539 ( .A(n84782), .B(n84781), .Z(n88096) );
  IV U104540 ( .A(n84783), .Z(n84784) );
  NOR U104541 ( .A(n84785), .B(n84784), .Z(n88089) );
  NOR U104542 ( .A(n88096), .B(n88089), .Z(n84786) );
  XOR U104543 ( .A(n88097), .B(n84786), .Z(n84787) );
  NOR U104544 ( .A(n84788), .B(n84787), .Z(n84791) );
  IV U104545 ( .A(n84788), .Z(n84790) );
  XOR U104546 ( .A(n88089), .B(n88097), .Z(n84789) );
  NOR U104547 ( .A(n84790), .B(n84789), .Z(n88093) );
  NOR U104548 ( .A(n84791), .B(n88093), .Z(n88078) );
  IV U104549 ( .A(n84792), .Z(n84794) );
  NOR U104550 ( .A(n84794), .B(n84793), .Z(n84795) );
  IV U104551 ( .A(n84795), .Z(n88080) );
  XOR U104552 ( .A(n88078), .B(n88080), .Z(n88081) );
  XOR U104553 ( .A(n88082), .B(n88081), .Z(n90654) );
  XOR U104554 ( .A(n90656), .B(n90654), .Z(n84803) );
  IV U104555 ( .A(n84796), .Z(n84798) );
  NOR U104556 ( .A(n84798), .B(n84797), .Z(n90657) );
  IV U104557 ( .A(n84799), .Z(n84801) );
  NOR U104558 ( .A(n84801), .B(n84800), .Z(n90658) );
  NOR U104559 ( .A(n90657), .B(n90658), .Z(n84802) );
  XOR U104560 ( .A(n84803), .B(n84802), .Z(n90674) );
  XOR U104561 ( .A(n90676), .B(n90674), .Z(n90679) );
  IV U104562 ( .A(n84807), .Z(n84804) );
  NOR U104563 ( .A(n84804), .B(n84805), .Z(n84811) );
  IV U104564 ( .A(n84805), .Z(n84806) );
  NOR U104565 ( .A(n84807), .B(n84806), .Z(n84808) );
  NOR U104566 ( .A(n84809), .B(n84808), .Z(n84810) );
  NOR U104567 ( .A(n84811), .B(n84810), .Z(n90677) );
  XOR U104568 ( .A(n90679), .B(n90677), .Z(n90685) );
  IV U104569 ( .A(n84812), .Z(n84813) );
  NOR U104570 ( .A(n84814), .B(n84813), .Z(n90686) );
  XOR U104571 ( .A(n90685), .B(n90686), .Z(n84815) );
  XOR U104572 ( .A(n90688), .B(n84815), .Z(n90667) );
  XOR U104573 ( .A(n90668), .B(n90667), .Z(n90670) );
  XOR U104574 ( .A(n90671), .B(n90670), .Z(n84816) );
  IV U104575 ( .A(n84816), .Z(n90706) );
  IV U104576 ( .A(n84817), .Z(n84818) );
  NOR U104577 ( .A(n84823), .B(n84818), .Z(n90705) );
  NOR U104578 ( .A(n90704), .B(n90705), .Z(n84819) );
  XOR U104579 ( .A(n90706), .B(n84819), .Z(n84829) );
  IV U104580 ( .A(n84829), .Z(n84820) );
  NOR U104581 ( .A(n84821), .B(n84820), .Z(n90714) );
  XOR U104582 ( .A(n90704), .B(n90706), .Z(n84828) );
  IV U104583 ( .A(n84822), .Z(n84826) );
  NOR U104584 ( .A(n84824), .B(n84823), .Z(n84825) );
  IV U104585 ( .A(n84825), .Z(n84833) );
  NOR U104586 ( .A(n84826), .B(n84833), .Z(n84830) );
  IV U104587 ( .A(n84830), .Z(n84827) );
  NOR U104588 ( .A(n84828), .B(n84827), .Z(n90703) );
  NOR U104589 ( .A(n84830), .B(n84829), .Z(n84831) );
  NOR U104590 ( .A(n90703), .B(n84831), .Z(n90698) );
  IV U104591 ( .A(n84832), .Z(n84834) );
  NOR U104592 ( .A(n84834), .B(n84833), .Z(n90699) );
  XOR U104593 ( .A(n90698), .B(n90699), .Z(n84835) );
  NOR U104594 ( .A(n84836), .B(n84835), .Z(n84837) );
  NOR U104595 ( .A(n90714), .B(n84837), .Z(n90710) );
  XOR U104596 ( .A(n90709), .B(n90710), .Z(n88050) );
  XOR U104597 ( .A(n88052), .B(n88050), .Z(n88043) );
  XOR U104598 ( .A(n84838), .B(n88043), .Z(n88041) );
  XOR U104599 ( .A(n88040), .B(n88041), .Z(n84839) );
  IV U104600 ( .A(n84839), .Z(n88034) );
  NOR U104601 ( .A(n88037), .B(n88034), .Z(n84845) );
  NOR U104602 ( .A(n88033), .B(n84839), .Z(n84843) );
  IV U104603 ( .A(n84840), .Z(n84842) );
  NOR U104604 ( .A(n84842), .B(n84841), .Z(n88032) );
  XOR U104605 ( .A(n84843), .B(n88032), .Z(n84844) );
  NOR U104606 ( .A(n84845), .B(n84844), .Z(n88067) );
  IV U104607 ( .A(n84846), .Z(n84848) );
  NOR U104608 ( .A(n84848), .B(n84847), .Z(n88066) );
  IV U104609 ( .A(n88066), .Z(n88068) );
  XOR U104610 ( .A(n88067), .B(n88068), .Z(n88029) );
  IV U104611 ( .A(n84849), .Z(n84851) );
  NOR U104612 ( .A(n84851), .B(n84850), .Z(n88071) );
  IV U104613 ( .A(n84852), .Z(n84854) );
  NOR U104614 ( .A(n84854), .B(n84853), .Z(n88027) );
  NOR U104615 ( .A(n88071), .B(n88027), .Z(n84855) );
  XOR U104616 ( .A(n88029), .B(n84855), .Z(n88024) );
  XOR U104617 ( .A(n88025), .B(n88024), .Z(n88060) );
  XOR U104618 ( .A(n88059), .B(n88060), .Z(n88062) );
  XOR U104619 ( .A(n88063), .B(n88062), .Z(n84862) );
  NOR U104620 ( .A(n84861), .B(n84862), .Z(n84856) );
  IV U104621 ( .A(n84856), .Z(n84860) );
  IV U104622 ( .A(n84857), .Z(n84858) );
  NOR U104623 ( .A(n84859), .B(n84858), .Z(n84865) );
  NOR U104624 ( .A(n84860), .B(n84865), .Z(n84870) );
  IV U104625 ( .A(n84861), .Z(n84866) );
  XOR U104626 ( .A(n84865), .B(n84866), .Z(n84864) );
  IV U104627 ( .A(n84862), .Z(n84863) );
  NOR U104628 ( .A(n84864), .B(n84863), .Z(n84869) );
  IV U104629 ( .A(n84865), .Z(n84867) );
  NOR U104630 ( .A(n84867), .B(n84866), .Z(n84868) );
  NOR U104631 ( .A(n84869), .B(n84868), .Z(n88000) );
  IV U104632 ( .A(n88000), .Z(n87997) );
  NOR U104633 ( .A(n84870), .B(n87997), .Z(n84877) );
  NOR U104634 ( .A(n84878), .B(n84877), .Z(n84876) );
  IV U104635 ( .A(n84876), .Z(n84873) );
  IV U104636 ( .A(n84871), .Z(n84872) );
  NOR U104637 ( .A(n84872), .B(n84886), .Z(n84874) );
  NOR U104638 ( .A(n84873), .B(n84874), .Z(n84883) );
  IV U104639 ( .A(n84874), .Z(n84875) );
  NOR U104640 ( .A(n84876), .B(n84875), .Z(n87999) );
  IV U104641 ( .A(n84877), .Z(n84880) );
  IV U104642 ( .A(n84878), .Z(n84879) );
  NOR U104643 ( .A(n84880), .B(n84879), .Z(n84881) );
  NOR U104644 ( .A(n87999), .B(n84881), .Z(n87998) );
  IV U104645 ( .A(n87998), .Z(n84882) );
  NOR U104646 ( .A(n84883), .B(n84882), .Z(n84884) );
  IV U104647 ( .A(n84884), .Z(n87989) );
  IV U104648 ( .A(n84885), .Z(n84887) );
  NOR U104649 ( .A(n84887), .B(n84886), .Z(n87987) );
  XOR U104650 ( .A(n87989), .B(n87987), .Z(n87992) );
  IV U104651 ( .A(n84888), .Z(n84895) );
  NOR U104652 ( .A(n84890), .B(n84889), .Z(n84891) );
  IV U104653 ( .A(n84891), .Z(n84892) );
  NOR U104654 ( .A(n84893), .B(n84892), .Z(n84894) );
  IV U104655 ( .A(n84894), .Z(n84897) );
  NOR U104656 ( .A(n84895), .B(n84897), .Z(n87990) );
  XOR U104657 ( .A(n87992), .B(n87990), .Z(n87981) );
  IV U104658 ( .A(n84896), .Z(n84898) );
  NOR U104659 ( .A(n84898), .B(n84897), .Z(n87979) );
  XOR U104660 ( .A(n87981), .B(n87979), .Z(n87983) );
  XOR U104661 ( .A(n87982), .B(n87983), .Z(n88013) );
  XOR U104662 ( .A(n88012), .B(n88013), .Z(n88016) );
  XOR U104663 ( .A(n88015), .B(n88016), .Z(n87978) );
  NOR U104664 ( .A(n84900), .B(n84899), .Z(n84902) );
  NOR U104665 ( .A(n84902), .B(n84901), .Z(n87977) );
  XOR U104666 ( .A(n87978), .B(n87977), .Z(n88007) );
  IV U104667 ( .A(n84903), .Z(n84905) );
  NOR U104668 ( .A(n84905), .B(n84904), .Z(n88005) );
  XOR U104669 ( .A(n88007), .B(n88005), .Z(n88008) );
  XOR U104670 ( .A(n88009), .B(n88008), .Z(n87931) );
  XOR U104671 ( .A(n87930), .B(n87931), .Z(n84906) );
  IV U104672 ( .A(n84906), .Z(n87945) );
  NOR U104673 ( .A(n87948), .B(n87945), .Z(n84913) );
  NOR U104674 ( .A(n84907), .B(n84906), .Z(n84911) );
  IV U104675 ( .A(n84908), .Z(n84909) );
  NOR U104676 ( .A(n84910), .B(n84909), .Z(n87947) );
  XOR U104677 ( .A(n84911), .B(n87947), .Z(n84912) );
  NOR U104678 ( .A(n84913), .B(n84912), .Z(n84914) );
  IV U104679 ( .A(n84914), .Z(n87943) );
  XOR U104680 ( .A(n87942), .B(n87943), .Z(n84922) );
  IV U104681 ( .A(n84922), .Z(n84915) );
  NOR U104682 ( .A(n84921), .B(n84915), .Z(n84916) );
  IV U104683 ( .A(n84916), .Z(n84920) );
  IV U104684 ( .A(n84917), .Z(n84919) );
  NOR U104685 ( .A(n84919), .B(n84918), .Z(n84924) );
  NOR U104686 ( .A(n84920), .B(n84924), .Z(n84929) );
  IV U104687 ( .A(n84921), .Z(n84925) );
  XOR U104688 ( .A(n84924), .B(n84925), .Z(n84923) );
  NOR U104689 ( .A(n84923), .B(n84922), .Z(n84928) );
  IV U104690 ( .A(n84924), .Z(n84926) );
  NOR U104691 ( .A(n84926), .B(n84925), .Z(n84927) );
  NOR U104692 ( .A(n84928), .B(n84927), .Z(n87937) );
  IV U104693 ( .A(n87937), .Z(n87934) );
  NOR U104694 ( .A(n84929), .B(n87934), .Z(n84937) );
  NOR U104695 ( .A(n84938), .B(n84937), .Z(n84936) );
  IV U104696 ( .A(n84936), .Z(n84933) );
  IV U104697 ( .A(n84930), .Z(n84932) );
  NOR U104698 ( .A(n84932), .B(n84931), .Z(n84934) );
  NOR U104699 ( .A(n84933), .B(n84934), .Z(n84943) );
  IV U104700 ( .A(n84934), .Z(n84935) );
  NOR U104701 ( .A(n84936), .B(n84935), .Z(n87936) );
  IV U104702 ( .A(n84937), .Z(n84940) );
  IV U104703 ( .A(n84938), .Z(n84939) );
  NOR U104704 ( .A(n84940), .B(n84939), .Z(n84941) );
  NOR U104705 ( .A(n87936), .B(n84941), .Z(n87935) );
  IV U104706 ( .A(n87935), .Z(n84942) );
  NOR U104707 ( .A(n84943), .B(n84942), .Z(n84950) );
  NOR U104708 ( .A(n84949), .B(n84950), .Z(n84944) );
  IV U104709 ( .A(n84944), .Z(n84948) );
  IV U104710 ( .A(n84945), .Z(n84946) );
  NOR U104711 ( .A(n84947), .B(n84946), .Z(n84953) );
  NOR U104712 ( .A(n84948), .B(n84953), .Z(n84959) );
  IV U104713 ( .A(n84949), .Z(n84954) );
  XOR U104714 ( .A(n84953), .B(n84954), .Z(n84952) );
  IV U104715 ( .A(n84950), .Z(n84951) );
  NOR U104716 ( .A(n84952), .B(n84951), .Z(n84957) );
  IV U104717 ( .A(n84953), .Z(n84955) );
  NOR U104718 ( .A(n84955), .B(n84954), .Z(n84956) );
  NOR U104719 ( .A(n84957), .B(n84956), .Z(n84958) );
  IV U104720 ( .A(n84958), .Z(n87964) );
  NOR U104721 ( .A(n84959), .B(n87964), .Z(n87970) );
  IV U104722 ( .A(n84960), .Z(n84961) );
  NOR U104723 ( .A(n84962), .B(n84961), .Z(n84968) );
  IV U104724 ( .A(n84968), .Z(n87973) );
  XOR U104725 ( .A(n87970), .B(n87973), .Z(n84966) );
  IV U104726 ( .A(n84963), .Z(n84964) );
  NOR U104727 ( .A(n84965), .B(n84964), .Z(n87969) );
  XOR U104728 ( .A(n84966), .B(n87969), .Z(n84967) );
  NOR U104729 ( .A(n87972), .B(n84967), .Z(n84972) );
  IV U104730 ( .A(n87972), .Z(n87967) );
  NOR U104731 ( .A(n87970), .B(n84968), .Z(n84969) );
  IV U104732 ( .A(n84969), .Z(n84970) );
  NOR U104733 ( .A(n87967), .B(n84970), .Z(n84971) );
  NOR U104734 ( .A(n84972), .B(n84971), .Z(n87955) );
  XOR U104735 ( .A(n87956), .B(n87955), .Z(n87957) );
  IV U104736 ( .A(n84973), .Z(n84975) );
  NOR U104737 ( .A(n84975), .B(n84974), .Z(n84980) );
  IV U104738 ( .A(n84976), .Z(n84977) );
  NOR U104739 ( .A(n84978), .B(n84977), .Z(n84979) );
  NOR U104740 ( .A(n84980), .B(n84979), .Z(n87959) );
  XOR U104741 ( .A(n87957), .B(n87959), .Z(n90741) );
  XOR U104742 ( .A(n90738), .B(n90741), .Z(n84981) );
  NOR U104743 ( .A(n84982), .B(n84981), .Z(n90737) );
  IV U104744 ( .A(n84983), .Z(n84985) );
  NOR U104745 ( .A(n84985), .B(n84984), .Z(n90740) );
  NOR U104746 ( .A(n90738), .B(n90740), .Z(n84986) );
  XOR U104747 ( .A(n90741), .B(n84986), .Z(n84987) );
  NOR U104748 ( .A(n84988), .B(n84987), .Z(n84989) );
  NOR U104749 ( .A(n90737), .B(n84989), .Z(n84990) );
  IV U104750 ( .A(n84990), .Z(n90734) );
  XOR U104751 ( .A(n90733), .B(n90734), .Z(n90726) );
  XOR U104752 ( .A(n90725), .B(n90726), .Z(n90730) );
  IV U104753 ( .A(n84991), .Z(n84994) );
  IV U104754 ( .A(n84992), .Z(n84993) );
  NOR U104755 ( .A(n84994), .B(n84993), .Z(n90728) );
  XOR U104756 ( .A(n90730), .B(n90728), .Z(n87887) );
  XOR U104757 ( .A(n87889), .B(n87887), .Z(n87901) );
  IV U104758 ( .A(n84995), .Z(n84996) );
  NOR U104759 ( .A(n84997), .B(n84996), .Z(n87886) );
  IV U104760 ( .A(n84998), .Z(n84999) );
  NOR U104761 ( .A(n84999), .B(n85002), .Z(n87899) );
  NOR U104762 ( .A(n87886), .B(n87899), .Z(n85000) );
  XOR U104763 ( .A(n87901), .B(n85000), .Z(n87896) );
  IV U104764 ( .A(n85001), .Z(n85003) );
  NOR U104765 ( .A(n85003), .B(n85002), .Z(n85004) );
  IV U104766 ( .A(n85004), .Z(n87897) );
  XOR U104767 ( .A(n87896), .B(n87897), .Z(n87883) );
  IV U104768 ( .A(n85005), .Z(n85007) );
  NOR U104769 ( .A(n85007), .B(n85006), .Z(n85013) );
  IV U104770 ( .A(n85013), .Z(n85008) );
  NOR U104771 ( .A(n87883), .B(n85008), .Z(n87915) );
  NOR U104772 ( .A(n85010), .B(n85009), .Z(n85011) );
  IV U104773 ( .A(n85011), .Z(n87884) );
  XOR U104774 ( .A(n87884), .B(n87883), .Z(n85012) );
  NOR U104775 ( .A(n85013), .B(n85012), .Z(n85017) );
  NOR U104776 ( .A(n87915), .B(n85017), .Z(n85014) );
  NOR U104777 ( .A(n85015), .B(n85014), .Z(n85018) );
  IV U104778 ( .A(n85015), .Z(n85016) );
  NOR U104779 ( .A(n85017), .B(n85016), .Z(n87914) );
  NOR U104780 ( .A(n85018), .B(n87914), .Z(n87906) );
  XOR U104781 ( .A(n87908), .B(n87906), .Z(n87910) );
  XOR U104782 ( .A(n87909), .B(n87910), .Z(n87920) );
  NOR U104783 ( .A(n85019), .B(n85020), .Z(n85029) );
  IV U104784 ( .A(n85020), .Z(n85021) );
  NOR U104785 ( .A(n85022), .B(n85021), .Z(n85027) );
  NOR U104786 ( .A(n85024), .B(n85023), .Z(n85025) );
  IV U104787 ( .A(n85025), .Z(n85026) );
  NOR U104788 ( .A(n85027), .B(n85026), .Z(n85028) );
  NOR U104789 ( .A(n85029), .B(n85028), .Z(n87918) );
  XOR U104790 ( .A(n87920), .B(n87918), .Z(n87923) );
  IV U104791 ( .A(n85030), .Z(n85032) );
  NOR U104792 ( .A(n85032), .B(n85031), .Z(n87921) );
  XOR U104793 ( .A(n87923), .B(n87921), .Z(n90754) );
  XOR U104794 ( .A(n90753), .B(n90754), .Z(n90757) );
  XOR U104795 ( .A(n90756), .B(n90757), .Z(n85038) );
  NOR U104796 ( .A(n85042), .B(n85038), .Z(n85037) );
  NOR U104797 ( .A(n85034), .B(n85033), .Z(n85039) );
  IV U104798 ( .A(n85039), .Z(n85035) );
  NOR U104799 ( .A(n90757), .B(n85035), .Z(n85036) );
  NOR U104800 ( .A(n85037), .B(n85036), .Z(n90752) );
  IV U104801 ( .A(n90752), .Z(n85041) );
  IV U104802 ( .A(n85038), .Z(n85043) );
  NOR U104803 ( .A(n85039), .B(n85043), .Z(n85040) );
  NOR U104804 ( .A(n85041), .B(n85040), .Z(n85045) );
  NOR U104805 ( .A(n85043), .B(n85042), .Z(n85044) );
  NOR U104806 ( .A(n85045), .B(n85044), .Z(n90750) );
  IV U104807 ( .A(n85046), .Z(n85048) );
  NOR U104808 ( .A(n85048), .B(n85047), .Z(n85049) );
  NOR U104809 ( .A(n90748), .B(n85049), .Z(n85050) );
  XOR U104810 ( .A(n90750), .B(n85050), .Z(n87857) );
  IV U104811 ( .A(n85051), .Z(n85053) );
  NOR U104812 ( .A(n85053), .B(n85052), .Z(n87858) );
  IV U104813 ( .A(n85054), .Z(n90745) );
  IV U104814 ( .A(n85055), .Z(n85056) );
  NOR U104815 ( .A(n90745), .B(n85056), .Z(n85057) );
  NOR U104816 ( .A(n87858), .B(n85057), .Z(n85058) );
  XOR U104817 ( .A(n87857), .B(n85058), .Z(n87856) );
  XOR U104818 ( .A(n87854), .B(n87856), .Z(n87866) );
  XOR U104819 ( .A(n87865), .B(n87866), .Z(n87869) );
  IV U104820 ( .A(n85059), .Z(n85060) );
  NOR U104821 ( .A(n85061), .B(n85060), .Z(n87868) );
  IV U104822 ( .A(n85062), .Z(n85064) );
  NOR U104823 ( .A(n85064), .B(n85063), .Z(n87863) );
  NOR U104824 ( .A(n87868), .B(n87863), .Z(n85065) );
  XOR U104825 ( .A(n87869), .B(n85065), .Z(n85066) );
  NOR U104826 ( .A(n85067), .B(n85066), .Z(n85070) );
  IV U104827 ( .A(n85067), .Z(n85069) );
  XOR U104828 ( .A(n87863), .B(n87869), .Z(n85068) );
  NOR U104829 ( .A(n85069), .B(n85068), .Z(n87882) );
  NOR U104830 ( .A(n85070), .B(n87882), .Z(n87878) );
  NOR U104831 ( .A(n85072), .B(n85071), .Z(n85079) );
  NOR U104832 ( .A(n85074), .B(n85073), .Z(n85077) );
  IV U104833 ( .A(n85075), .Z(n85076) );
  NOR U104834 ( .A(n85077), .B(n85076), .Z(n85078) );
  NOR U104835 ( .A(n85079), .B(n85078), .Z(n87880) );
  XOR U104836 ( .A(n87878), .B(n87880), .Z(n87830) );
  XOR U104837 ( .A(n87829), .B(n87830), .Z(n87832) );
  IV U104838 ( .A(n85080), .Z(n85081) );
  NOR U104839 ( .A(n85082), .B(n85081), .Z(n85087) );
  IV U104840 ( .A(n85083), .Z(n85085) );
  NOR U104841 ( .A(n85085), .B(n85084), .Z(n85086) );
  NOR U104842 ( .A(n85087), .B(n85086), .Z(n87833) );
  XOR U104843 ( .A(n87832), .B(n87833), .Z(n85088) );
  IV U104844 ( .A(n85088), .Z(n87822) );
  XOR U104845 ( .A(n87821), .B(n87822), .Z(n87825) );
  XOR U104846 ( .A(n87824), .B(n87825), .Z(n87847) );
  XOR U104847 ( .A(n87846), .B(n87847), .Z(n87851) );
  XOR U104848 ( .A(n87849), .B(n87851), .Z(n90779) );
  XOR U104849 ( .A(n90778), .B(n90779), .Z(n90783) );
  XOR U104850 ( .A(n90781), .B(n90783), .Z(n90777) );
  XOR U104851 ( .A(n90775), .B(n90777), .Z(n87840) );
  XOR U104852 ( .A(n87838), .B(n87840), .Z(n87843) );
  XOR U104853 ( .A(n87841), .B(n87843), .Z(n87809) );
  XOR U104854 ( .A(n87808), .B(n87809), .Z(n87812) );
  XOR U104855 ( .A(n87811), .B(n87812), .Z(n87818) );
  XOR U104856 ( .A(n85089), .B(n87818), .Z(n87801) );
  XOR U104857 ( .A(n87803), .B(n87801), .Z(n87760) );
  XOR U104858 ( .A(n87758), .B(n87760), .Z(n87761) );
  XOR U104859 ( .A(n87762), .B(n87761), .Z(n87768) );
  IV U104860 ( .A(n87768), .Z(n87776) );
  NOR U104861 ( .A(n85090), .B(n87776), .Z(n87777) );
  IV U104862 ( .A(n85091), .Z(n85092) );
  NOR U104863 ( .A(n85093), .B(n85092), .Z(n87774) );
  XOR U104864 ( .A(n87768), .B(n87774), .Z(n85094) );
  NOR U104865 ( .A(n85095), .B(n85094), .Z(n87772) );
  NOR U104866 ( .A(n87777), .B(n87772), .Z(n85103) );
  IV U104867 ( .A(n85096), .Z(n85097) );
  NOR U104868 ( .A(n85098), .B(n85097), .Z(n87767) );
  IV U104869 ( .A(n85099), .Z(n85101) );
  NOR U104870 ( .A(n85101), .B(n85100), .Z(n87771) );
  NOR U104871 ( .A(n87767), .B(n87771), .Z(n85102) );
  XOR U104872 ( .A(n85103), .B(n85102), .Z(n87753) );
  IV U104873 ( .A(n85104), .Z(n85106) );
  NOR U104874 ( .A(n85106), .B(n85105), .Z(n87751) );
  XOR U104875 ( .A(n87753), .B(n87751), .Z(n87754) );
  XOR U104876 ( .A(n85107), .B(n87754), .Z(n87787) );
  XOR U104877 ( .A(n87788), .B(n87787), .Z(n85114) );
  NOR U104878 ( .A(n85113), .B(n85114), .Z(n85108) );
  IV U104879 ( .A(n85108), .Z(n85112) );
  IV U104880 ( .A(n85109), .Z(n85111) );
  NOR U104881 ( .A(n85111), .B(n85110), .Z(n85117) );
  NOR U104882 ( .A(n85112), .B(n85117), .Z(n85123) );
  IV U104883 ( .A(n85113), .Z(n85118) );
  XOR U104884 ( .A(n85117), .B(n85118), .Z(n85116) );
  IV U104885 ( .A(n85114), .Z(n85115) );
  NOR U104886 ( .A(n85116), .B(n85115), .Z(n85121) );
  IV U104887 ( .A(n85117), .Z(n85119) );
  NOR U104888 ( .A(n85119), .B(n85118), .Z(n85120) );
  NOR U104889 ( .A(n85121), .B(n85120), .Z(n85122) );
  IV U104890 ( .A(n85122), .Z(n87749) );
  NOR U104891 ( .A(n85123), .B(n87749), .Z(n85124) );
  IV U104892 ( .A(n85124), .Z(n87747) );
  XOR U104893 ( .A(n87746), .B(n87747), .Z(n87791) );
  XOR U104894 ( .A(n87789), .B(n87791), .Z(n87793) );
  XOR U104895 ( .A(n87792), .B(n87793), .Z(n87734) );
  XOR U104896 ( .A(n87732), .B(n87734), .Z(n87735) );
  XOR U104897 ( .A(n87736), .B(n87735), .Z(n85125) );
  IV U104898 ( .A(n85125), .Z(n90796) );
  XOR U104899 ( .A(n90797), .B(n90796), .Z(n85126) );
  IV U104900 ( .A(n85126), .Z(n90801) );
  NOR U104901 ( .A(n90804), .B(n90801), .Z(n85135) );
  NOR U104902 ( .A(n85127), .B(n85126), .Z(n85133) );
  IV U104903 ( .A(n85128), .Z(n85129) );
  NOR U104904 ( .A(n85129), .B(n85138), .Z(n85130) );
  IV U104905 ( .A(n85130), .Z(n85131) );
  NOR U104906 ( .A(n85132), .B(n85131), .Z(n90803) );
  XOR U104907 ( .A(n85133), .B(n90803), .Z(n85134) );
  NOR U104908 ( .A(n85135), .B(n85134), .Z(n85136) );
  IV U104909 ( .A(n85136), .Z(n90800) );
  IV U104910 ( .A(n85137), .Z(n85139) );
  NOR U104911 ( .A(n85139), .B(n85138), .Z(n90798) );
  XOR U104912 ( .A(n90800), .B(n90798), .Z(n90831) );
  XOR U104913 ( .A(n85140), .B(n90831), .Z(n85141) );
  IV U104914 ( .A(n85141), .Z(n87743) );
  IV U104915 ( .A(n85142), .Z(n85144) );
  NOR U104916 ( .A(n85144), .B(n85143), .Z(n87741) );
  XOR U104917 ( .A(n87743), .B(n87741), .Z(n90822) );
  XOR U104918 ( .A(n90821), .B(n90822), .Z(n90825) );
  IV U104919 ( .A(n85145), .Z(n85147) );
  NOR U104920 ( .A(n85147), .B(n85146), .Z(n90824) );
  IV U104921 ( .A(n85148), .Z(n85150) );
  NOR U104922 ( .A(n85150), .B(n85149), .Z(n87727) );
  NOR U104923 ( .A(n90824), .B(n87727), .Z(n85151) );
  XOR U104924 ( .A(n90825), .B(n85151), .Z(n87720) );
  IV U104925 ( .A(n85152), .Z(n85154) );
  NOR U104926 ( .A(n85154), .B(n85153), .Z(n87726) );
  IV U104927 ( .A(n85155), .Z(n85156) );
  NOR U104928 ( .A(n85157), .B(n85156), .Z(n87721) );
  NOR U104929 ( .A(n87726), .B(n87721), .Z(n85158) );
  XOR U104930 ( .A(n87720), .B(n85158), .Z(n87718) );
  XOR U104931 ( .A(n87717), .B(n87718), .Z(n90857) );
  IV U104932 ( .A(n85159), .Z(n85160) );
  NOR U104933 ( .A(n85161), .B(n85160), .Z(n87715) );
  IV U104934 ( .A(n85162), .Z(n85163) );
  NOR U104935 ( .A(n85164), .B(n85163), .Z(n90855) );
  NOR U104936 ( .A(n87715), .B(n90855), .Z(n85165) );
  XOR U104937 ( .A(n90857), .B(n85165), .Z(n90851) );
  XOR U104938 ( .A(n90852), .B(n90851), .Z(n90844) );
  XOR U104939 ( .A(n90846), .B(n90844), .Z(n87712) );
  IV U104940 ( .A(n85166), .Z(n85168) );
  NOR U104941 ( .A(n85168), .B(n85167), .Z(n87710) );
  NOR U104942 ( .A(n90848), .B(n87710), .Z(n85169) );
  XOR U104943 ( .A(n87712), .B(n85169), .Z(n87681) );
  XOR U104944 ( .A(n85170), .B(n87681), .Z(n87685) );
  XOR U104945 ( .A(n87684), .B(n87685), .Z(n87675) );
  XOR U104946 ( .A(n87673), .B(n87675), .Z(n87677) );
  XOR U104947 ( .A(n87676), .B(n87677), .Z(n87701) );
  XOR U104948 ( .A(n87699), .B(n87701), .Z(n87704) );
  XOR U104949 ( .A(n87702), .B(n87704), .Z(n87663) );
  XOR U104950 ( .A(n87661), .B(n87663), .Z(n87666) );
  XOR U104951 ( .A(n87664), .B(n87666), .Z(n87692) );
  XOR U104952 ( .A(n87691), .B(n87692), .Z(n87696) );
  XOR U104953 ( .A(n87694), .B(n87696), .Z(n87669) );
  XOR U104954 ( .A(n87670), .B(n87669), .Z(n90882) );
  XOR U104955 ( .A(n90884), .B(n90882), .Z(n90887) );
  IV U104956 ( .A(n85171), .Z(n85173) );
  NOR U104957 ( .A(n85173), .B(n85172), .Z(n90885) );
  XOR U104958 ( .A(n90887), .B(n90885), .Z(n90875) );
  XOR U104959 ( .A(n90874), .B(n90875), .Z(n90878) );
  XOR U104960 ( .A(n90877), .B(n90878), .Z(n87659) );
  IV U104961 ( .A(n87659), .Z(n85182) );
  XOR U104962 ( .A(n87656), .B(n85182), .Z(n85177) );
  IV U104963 ( .A(n90907), .Z(n85175) );
  NOR U104964 ( .A(n85175), .B(n85174), .Z(n90905) );
  IV U104965 ( .A(n90905), .Z(n85176) );
  NOR U104966 ( .A(n85177), .B(n85176), .Z(n85184) );
  IV U104967 ( .A(n85178), .Z(n85179) );
  NOR U104968 ( .A(n85180), .B(n85179), .Z(n87658) );
  NOR U104969 ( .A(n87656), .B(n87658), .Z(n85181) );
  XOR U104970 ( .A(n85182), .B(n85181), .Z(n90908) );
  NOR U104971 ( .A(n90905), .B(n90908), .Z(n85183) );
  NOR U104972 ( .A(n85184), .B(n85183), .Z(n90917) );
  XOR U104973 ( .A(n85194), .B(n90917), .Z(n85185) );
  NOR U104974 ( .A(n85186), .B(n85185), .Z(n90915) );
  IV U104975 ( .A(n85187), .Z(n85188) );
  NOR U104976 ( .A(n85189), .B(n85188), .Z(n85190) );
  IV U104977 ( .A(n85190), .Z(n90920) );
  IV U104978 ( .A(n85191), .Z(n85193) );
  NOR U104979 ( .A(n85193), .B(n85192), .Z(n90916) );
  NOR U104980 ( .A(n85194), .B(n90916), .Z(n85195) );
  IV U104981 ( .A(n85195), .Z(n85196) );
  XOR U104982 ( .A(n85196), .B(n90917), .Z(n90919) );
  XOR U104983 ( .A(n90920), .B(n90919), .Z(n85197) );
  NOR U104984 ( .A(n85198), .B(n85197), .Z(n85199) );
  NOR U104985 ( .A(n90915), .B(n85199), .Z(n90911) );
  IV U104986 ( .A(n85200), .Z(n85201) );
  NOR U104987 ( .A(n85201), .B(n85211), .Z(n85202) );
  IV U104988 ( .A(n85202), .Z(n90912) );
  XOR U104989 ( .A(n90911), .B(n90912), .Z(n87647) );
  IV U104990 ( .A(n85203), .Z(n85205) );
  NOR U104991 ( .A(n85205), .B(n85204), .Z(n87642) );
  IV U104992 ( .A(n85206), .Z(n85208) );
  NOR U104993 ( .A(n85208), .B(n85207), .Z(n85213) );
  IV U104994 ( .A(n85209), .Z(n85210) );
  NOR U104995 ( .A(n85211), .B(n85210), .Z(n85212) );
  NOR U104996 ( .A(n85213), .B(n85212), .Z(n87641) );
  IV U104997 ( .A(n87641), .Z(n87648) );
  XOR U104998 ( .A(n87642), .B(n87648), .Z(n85214) );
  XOR U104999 ( .A(n87647), .B(n85214), .Z(n87640) );
  XOR U105000 ( .A(n85215), .B(n87640), .Z(n87652) );
  XOR U105001 ( .A(n87653), .B(n87652), .Z(n87654) );
  IV U105002 ( .A(n85216), .Z(n85217) );
  NOR U105003 ( .A(n85218), .B(n85217), .Z(n85223) );
  IV U105004 ( .A(n85219), .Z(n85221) );
  NOR U105005 ( .A(n85221), .B(n85220), .Z(n85222) );
  NOR U105006 ( .A(n85223), .B(n85222), .Z(n87655) );
  XOR U105007 ( .A(n87654), .B(n87655), .Z(n85224) );
  IV U105008 ( .A(n85224), .Z(n90933) );
  XOR U105009 ( .A(n90932), .B(n90933), .Z(n90937) );
  XOR U105010 ( .A(n90935), .B(n90937), .Z(n87629) );
  XOR U105011 ( .A(n87628), .B(n87629), .Z(n85231) );
  IV U105012 ( .A(n85231), .Z(n90926) );
  XOR U105013 ( .A(n87631), .B(n90926), .Z(n85225) );
  NOR U105014 ( .A(n85226), .B(n85225), .Z(n87635) );
  IV U105015 ( .A(n85227), .Z(n90929) );
  IV U105016 ( .A(n85228), .Z(n85229) );
  NOR U105017 ( .A(n85230), .B(n85229), .Z(n90925) );
  NOR U105018 ( .A(n90925), .B(n87631), .Z(n85232) );
  XOR U105019 ( .A(n85232), .B(n85231), .Z(n90928) );
  XOR U105020 ( .A(n90929), .B(n90928), .Z(n85233) );
  NOR U105021 ( .A(n85234), .B(n85233), .Z(n85235) );
  NOR U105022 ( .A(n87635), .B(n85235), .Z(n85236) );
  IV U105023 ( .A(n85236), .Z(n90959) );
  XOR U105024 ( .A(n90958), .B(n90959), .Z(n90963) );
  XOR U105025 ( .A(n90961), .B(n90963), .Z(n90951) );
  XOR U105026 ( .A(n90950), .B(n90951), .Z(n90955) );
  XOR U105027 ( .A(n90953), .B(n90955), .Z(n87621) );
  XOR U105028 ( .A(n87620), .B(n87621), .Z(n87624) );
  XOR U105029 ( .A(n87623), .B(n87624), .Z(n90973) );
  XOR U105030 ( .A(n90972), .B(n90973), .Z(n90983) );
  XOR U105031 ( .A(n90975), .B(n90983), .Z(n85237) );
  NOR U105032 ( .A(n85238), .B(n85237), .Z(n90986) );
  IV U105033 ( .A(n85239), .Z(n85241) );
  NOR U105034 ( .A(n85241), .B(n85240), .Z(n90982) );
  NOR U105035 ( .A(n90975), .B(n90982), .Z(n85242) );
  XOR U105036 ( .A(n90983), .B(n85242), .Z(n85243) );
  NOR U105037 ( .A(n85244), .B(n85243), .Z(n85245) );
  NOR U105038 ( .A(n90986), .B(n85245), .Z(n90979) );
  IV U105039 ( .A(n85246), .Z(n85248) );
  NOR U105040 ( .A(n85248), .B(n85247), .Z(n85249) );
  IV U105041 ( .A(n85249), .Z(n90981) );
  XOR U105042 ( .A(n90979), .B(n90981), .Z(n87613) );
  XOR U105043 ( .A(n87612), .B(n87613), .Z(n87617) );
  XOR U105044 ( .A(n87615), .B(n87617), .Z(n87586) );
  XOR U105045 ( .A(n87585), .B(n87586), .Z(n87589) );
  XOR U105046 ( .A(n87588), .B(n87589), .Z(n87567) );
  XOR U105047 ( .A(n85250), .B(n87567), .Z(n87572) );
  XOR U105048 ( .A(n87570), .B(n87572), .Z(n87580) );
  IV U105049 ( .A(n85251), .Z(n85252) );
  NOR U105050 ( .A(n85253), .B(n85252), .Z(n87569) );
  IV U105051 ( .A(n85254), .Z(n85255) );
  NOR U105052 ( .A(n85256), .B(n85255), .Z(n87578) );
  NOR U105053 ( .A(n87569), .B(n87578), .Z(n85257) );
  XOR U105054 ( .A(n87580), .B(n85257), .Z(n87575) );
  XOR U105055 ( .A(n87577), .B(n87575), .Z(n87562) );
  IV U105056 ( .A(n85258), .Z(n85260) );
  NOR U105057 ( .A(n85260), .B(n85259), .Z(n87560) );
  XOR U105058 ( .A(n87562), .B(n87560), .Z(n87563) );
  XOR U105059 ( .A(n87564), .B(n87563), .Z(n85261) );
  NOR U105060 ( .A(n85262), .B(n85261), .Z(n87600) );
  IV U105061 ( .A(n85262), .Z(n85263) );
  NOR U105062 ( .A(n85263), .B(n87563), .Z(n87598) );
  NOR U105063 ( .A(n87600), .B(n87598), .Z(n85267) );
  IV U105064 ( .A(n85264), .Z(n85265) );
  NOR U105065 ( .A(n85265), .B(n87602), .Z(n85266) );
  XOR U105066 ( .A(n85267), .B(n85266), .Z(n85275) );
  IV U105067 ( .A(n85268), .Z(n85270) );
  NOR U105068 ( .A(n85270), .B(n85269), .Z(n87597) );
  IV U105069 ( .A(n85271), .Z(n85272) );
  NOR U105070 ( .A(n85272), .B(n87602), .Z(n85273) );
  NOR U105071 ( .A(n87597), .B(n85273), .Z(n85274) );
  XOR U105072 ( .A(n85275), .B(n85274), .Z(n87596) );
  IV U105073 ( .A(n87596), .Z(n87605) );
  XOR U105074 ( .A(n87605), .B(n87595), .Z(n87551) );
  XOR U105075 ( .A(n87550), .B(n87551), .Z(n87554) );
  XOR U105076 ( .A(n87553), .B(n87554), .Z(n87544) );
  XOR U105077 ( .A(n87543), .B(n87544), .Z(n87546) );
  XOR U105078 ( .A(n85279), .B(n87546), .Z(n87538) );
  XOR U105079 ( .A(n85280), .B(n87538), .Z(n91012) );
  XOR U105080 ( .A(n91011), .B(n91012), .Z(n91015) );
  XOR U105081 ( .A(n91014), .B(n91015), .Z(n91001) );
  XOR U105082 ( .A(n91000), .B(n91001), .Z(n91004) );
  XOR U105083 ( .A(n91003), .B(n91004), .Z(n91058) );
  XOR U105084 ( .A(n91056), .B(n91058), .Z(n91060) );
  XOR U105085 ( .A(n91059), .B(n91060), .Z(n85287) );
  IV U105086 ( .A(n85281), .Z(n85285) );
  NOR U105087 ( .A(n85283), .B(n85282), .Z(n85284) );
  IV U105088 ( .A(n85284), .Z(n85296) );
  NOR U105089 ( .A(n85285), .B(n85296), .Z(n85293) );
  IV U105090 ( .A(n85293), .Z(n85286) );
  NOR U105091 ( .A(n85287), .B(n85286), .Z(n91033) );
  IV U105092 ( .A(n85288), .Z(n85290) );
  NOR U105093 ( .A(n85290), .B(n85289), .Z(n91030) );
  NOR U105094 ( .A(n91059), .B(n91030), .Z(n85291) );
  XOR U105095 ( .A(n91060), .B(n85291), .Z(n85292) );
  NOR U105096 ( .A(n85293), .B(n85292), .Z(n85294) );
  NOR U105097 ( .A(n91033), .B(n85294), .Z(n91036) );
  IV U105098 ( .A(n85295), .Z(n85297) );
  NOR U105099 ( .A(n85297), .B(n85296), .Z(n85298) );
  IV U105100 ( .A(n85298), .Z(n91037) );
  XOR U105101 ( .A(n91036), .B(n91037), .Z(n91040) );
  XOR U105102 ( .A(n91039), .B(n91040), .Z(n91029) );
  IV U105103 ( .A(n85299), .Z(n85300) );
  NOR U105104 ( .A(n85301), .B(n85300), .Z(n85302) );
  IV U105105 ( .A(n85302), .Z(n91028) );
  XOR U105106 ( .A(n91029), .B(n91028), .Z(n85303) );
  NOR U105107 ( .A(n85313), .B(n85303), .Z(n85315) );
  IV U105108 ( .A(n85304), .Z(n85305) );
  NOR U105109 ( .A(n85306), .B(n85305), .Z(n85311) );
  IV U105110 ( .A(n85307), .Z(n85308) );
  NOR U105111 ( .A(n85309), .B(n85308), .Z(n85310) );
  NOR U105112 ( .A(n85311), .B(n85310), .Z(n85312) );
  NOR U105113 ( .A(n85315), .B(n85312), .Z(n91051) );
  IV U105114 ( .A(n85312), .Z(n85317) );
  IV U105115 ( .A(n85313), .Z(n85314) );
  NOR U105116 ( .A(n85314), .B(n91029), .Z(n91050) );
  NOR U105117 ( .A(n85315), .B(n91050), .Z(n85316) );
  NOR U105118 ( .A(n85317), .B(n85316), .Z(n85318) );
  NOR U105119 ( .A(n91051), .B(n85318), .Z(n85319) );
  IV U105120 ( .A(n85319), .Z(n91048) );
  XOR U105121 ( .A(n91049), .B(n91048), .Z(n87535) );
  XOR U105122 ( .A(n87531), .B(n87535), .Z(n85327) );
  IV U105123 ( .A(n85320), .Z(n85321) );
  NOR U105124 ( .A(n85322), .B(n85321), .Z(n87528) );
  IV U105125 ( .A(n85323), .Z(n85325) );
  NOR U105126 ( .A(n85325), .B(n85324), .Z(n87530) );
  NOR U105127 ( .A(n87528), .B(n87530), .Z(n85326) );
  XOR U105128 ( .A(n85327), .B(n85326), .Z(n91078) );
  XOR U105129 ( .A(n91076), .B(n91078), .Z(n91081) );
  IV U105130 ( .A(n85328), .Z(n85335) );
  NOR U105131 ( .A(n85330), .B(n85329), .Z(n85331) );
  IV U105132 ( .A(n85331), .Z(n85332) );
  NOR U105133 ( .A(n85333), .B(n85332), .Z(n85334) );
  IV U105134 ( .A(n85334), .Z(n85337) );
  NOR U105135 ( .A(n85335), .B(n85337), .Z(n91079) );
  XOR U105136 ( .A(n91081), .B(n91079), .Z(n91071) );
  IV U105137 ( .A(n91071), .Z(n91069) );
  IV U105138 ( .A(n85336), .Z(n85338) );
  NOR U105139 ( .A(n85338), .B(n85337), .Z(n91068) );
  IV U105140 ( .A(n91068), .Z(n91070) );
  XOR U105141 ( .A(n91069), .B(n91070), .Z(n91095) );
  IV U105142 ( .A(n91095), .Z(n85346) );
  IV U105143 ( .A(n85339), .Z(n85340) );
  NOR U105144 ( .A(n85341), .B(n85340), .Z(n91073) );
  IV U105145 ( .A(n85342), .Z(n85343) );
  NOR U105146 ( .A(n85344), .B(n85343), .Z(n91093) );
  NOR U105147 ( .A(n91073), .B(n91093), .Z(n85345) );
  XOR U105148 ( .A(n85346), .B(n85345), .Z(n91092) );
  XOR U105149 ( .A(n91090), .B(n91092), .Z(n87521) );
  XOR U105150 ( .A(n87522), .B(n87521), .Z(n85347) );
  IV U105151 ( .A(n85347), .Z(n87525) );
  IV U105152 ( .A(n85348), .Z(n85351) );
  IV U105153 ( .A(n85349), .Z(n85350) );
  NOR U105154 ( .A(n85351), .B(n85350), .Z(n87523) );
  XOR U105155 ( .A(n87525), .B(n87523), .Z(n91100) );
  XOR U105156 ( .A(n91101), .B(n91100), .Z(n91102) );
  IV U105157 ( .A(n85352), .Z(n85353) );
  NOR U105158 ( .A(n85354), .B(n85353), .Z(n85359) );
  IV U105159 ( .A(n85355), .Z(n85356) );
  NOR U105160 ( .A(n85357), .B(n85356), .Z(n85358) );
  NOR U105161 ( .A(n85359), .B(n85358), .Z(n91104) );
  XOR U105162 ( .A(n91102), .B(n91104), .Z(n91121) );
  XOR U105163 ( .A(n85360), .B(n91121), .Z(n91113) );
  NOR U105164 ( .A(n85362), .B(n85361), .Z(n85372) );
  IV U105165 ( .A(n85372), .Z(n91115) );
  NOR U105166 ( .A(n91113), .B(n91115), .Z(n85374) );
  IV U105167 ( .A(n85363), .Z(n85365) );
  NOR U105168 ( .A(n85365), .B(n85364), .Z(n85368) );
  IV U105169 ( .A(n85368), .Z(n85367) );
  XOR U105170 ( .A(n91120), .B(n91121), .Z(n85366) );
  NOR U105171 ( .A(n85367), .B(n85366), .Z(n91123) );
  NOR U105172 ( .A(n91113), .B(n85368), .Z(n85369) );
  NOR U105173 ( .A(n91123), .B(n85369), .Z(n85370) );
  IV U105174 ( .A(n85370), .Z(n85371) );
  NOR U105175 ( .A(n85372), .B(n85371), .Z(n85373) );
  NOR U105176 ( .A(n85374), .B(n85373), .Z(n91116) );
  XOR U105177 ( .A(n91117), .B(n91116), .Z(n87513) );
  XOR U105178 ( .A(n87515), .B(n87513), .Z(n87517) );
  XOR U105179 ( .A(n87516), .B(n87517), .Z(n91143) );
  XOR U105180 ( .A(n91144), .B(n91143), .Z(n85381) );
  IV U105181 ( .A(n85381), .Z(n85375) );
  NOR U105182 ( .A(n85376), .B(n85375), .Z(n91132) );
  IV U105183 ( .A(n85377), .Z(n85380) );
  IV U105184 ( .A(n85378), .Z(n85379) );
  NOR U105185 ( .A(n85380), .B(n85379), .Z(n85382) );
  NOR U105186 ( .A(n85382), .B(n85381), .Z(n85384) );
  IV U105187 ( .A(n85382), .Z(n85383) );
  NOR U105188 ( .A(n85383), .B(n87517), .Z(n91131) );
  NOR U105189 ( .A(n85384), .B(n91131), .Z(n91163) );
  NOR U105190 ( .A(n85385), .B(n91163), .Z(n85386) );
  NOR U105191 ( .A(n91132), .B(n85386), .Z(n91133) );
  XOR U105192 ( .A(n85387), .B(n91133), .Z(n91150) );
  XOR U105193 ( .A(n85388), .B(n91150), .Z(n91162) );
  XOR U105194 ( .A(n91160), .B(n91162), .Z(n91146) );
  XOR U105195 ( .A(n91145), .B(n91146), .Z(n91176) );
  XOR U105196 ( .A(n91175), .B(n91176), .Z(n91178) );
  XOR U105197 ( .A(n91179), .B(n91178), .Z(n91157) );
  XOR U105198 ( .A(n91159), .B(n91157), .Z(n91180) );
  XOR U105199 ( .A(n91181), .B(n91180), .Z(n85391) );
  IV U105200 ( .A(n85391), .Z(n85389) );
  NOR U105201 ( .A(n85390), .B(n85389), .Z(n87511) );
  NOR U105202 ( .A(n85392), .B(n85391), .Z(n87509) );
  IV U105203 ( .A(n85393), .Z(n85394) );
  NOR U105204 ( .A(n85395), .B(n85394), .Z(n87508) );
  XOR U105205 ( .A(n87509), .B(n87508), .Z(n85396) );
  NOR U105206 ( .A(n87511), .B(n85396), .Z(n91196) );
  IV U105207 ( .A(n85397), .Z(n85398) );
  NOR U105208 ( .A(n85399), .B(n85398), .Z(n85400) );
  IV U105209 ( .A(n85400), .Z(n91197) );
  XOR U105210 ( .A(n91196), .B(n91197), .Z(n91201) );
  XOR U105211 ( .A(n91199), .B(n91201), .Z(n91194) );
  XOR U105212 ( .A(n91193), .B(n91194), .Z(n91188) );
  XOR U105213 ( .A(n91186), .B(n91188), .Z(n91189) );
  XOR U105214 ( .A(n91190), .B(n91189), .Z(n85407) );
  NOR U105215 ( .A(n85406), .B(n85407), .Z(n85401) );
  IV U105216 ( .A(n85401), .Z(n85405) );
  IV U105217 ( .A(n85402), .Z(n85404) );
  NOR U105218 ( .A(n85404), .B(n85403), .Z(n85410) );
  NOR U105219 ( .A(n85405), .B(n85410), .Z(n85416) );
  IV U105220 ( .A(n85406), .Z(n85411) );
  XOR U105221 ( .A(n85410), .B(n85411), .Z(n85409) );
  IV U105222 ( .A(n85407), .Z(n85408) );
  NOR U105223 ( .A(n85409), .B(n85408), .Z(n85414) );
  IV U105224 ( .A(n85410), .Z(n85412) );
  NOR U105225 ( .A(n85412), .B(n85411), .Z(n85413) );
  NOR U105226 ( .A(n85414), .B(n85413), .Z(n85415) );
  IV U105227 ( .A(n85415), .Z(n87491) );
  NOR U105228 ( .A(n85416), .B(n87491), .Z(n85417) );
  IV U105229 ( .A(n85417), .Z(n87488) );
  XOR U105230 ( .A(n87487), .B(n87488), .Z(n87498) );
  IV U105231 ( .A(n85418), .Z(n85421) );
  IV U105232 ( .A(n85419), .Z(n85420) );
  NOR U105233 ( .A(n85421), .B(n85420), .Z(n85422) );
  NOR U105234 ( .A(n85423), .B(n85422), .Z(n87494) );
  IV U105235 ( .A(n87494), .Z(n87499) );
  XOR U105236 ( .A(n87498), .B(n87499), .Z(n85424) );
  XOR U105237 ( .A(n85425), .B(n85424), .Z(n91217) );
  XOR U105238 ( .A(n91218), .B(n91217), .Z(n91220) );
  IV U105239 ( .A(n85426), .Z(n85427) );
  NOR U105240 ( .A(n85428), .B(n85427), .Z(n85433) );
  IV U105241 ( .A(n85429), .Z(n85430) );
  NOR U105242 ( .A(n85431), .B(n85430), .Z(n85432) );
  NOR U105243 ( .A(n85433), .B(n85432), .Z(n91221) );
  XOR U105244 ( .A(n91220), .B(n91221), .Z(n85434) );
  IV U105245 ( .A(n85434), .Z(n91232) );
  XOR U105246 ( .A(n91231), .B(n91232), .Z(n85435) );
  XOR U105247 ( .A(n85436), .B(n85435), .Z(n85437) );
  XOR U105248 ( .A(n85438), .B(n85437), .Z(n85439) );
  IV U105249 ( .A(n85439), .Z(n91238) );
  XOR U105250 ( .A(n91239), .B(n91238), .Z(n91252) );
  XOR U105251 ( .A(n91250), .B(n91252), .Z(n91246) );
  IV U105252 ( .A(n85440), .Z(n85441) );
  NOR U105253 ( .A(n85441), .B(n85444), .Z(n85450) );
  IV U105254 ( .A(n85450), .Z(n85442) );
  NOR U105255 ( .A(n91246), .B(n85442), .Z(n87484) );
  IV U105256 ( .A(n85443), .Z(n85445) );
  NOR U105257 ( .A(n85445), .B(n85444), .Z(n91251) );
  IV U105258 ( .A(n85446), .Z(n85448) );
  NOR U105259 ( .A(n85448), .B(n85447), .Z(n91244) );
  NOR U105260 ( .A(n91251), .B(n91244), .Z(n85449) );
  XOR U105261 ( .A(n85449), .B(n91246), .Z(n91241) );
  NOR U105262 ( .A(n85450), .B(n91241), .Z(n85451) );
  NOR U105263 ( .A(n87484), .B(n85451), .Z(n87478) );
  IV U105264 ( .A(n87478), .Z(n87476) );
  XOR U105265 ( .A(n87477), .B(n87476), .Z(n87458) );
  IV U105266 ( .A(n85452), .Z(n85453) );
  NOR U105267 ( .A(n85454), .B(n85453), .Z(n87457) );
  IV U105268 ( .A(n85455), .Z(n85456) );
  NOR U105269 ( .A(n85457), .B(n85456), .Z(n87480) );
  NOR U105270 ( .A(n91240), .B(n87480), .Z(n85458) );
  IV U105271 ( .A(n85458), .Z(n85459) );
  NOR U105272 ( .A(n87457), .B(n85459), .Z(n85460) );
  XOR U105273 ( .A(n87458), .B(n85460), .Z(n87471) );
  XOR U105274 ( .A(n87469), .B(n87471), .Z(n87464) );
  XOR U105275 ( .A(n85461), .B(n87464), .Z(n85462) );
  IV U105276 ( .A(n85462), .Z(n87462) );
  XOR U105277 ( .A(n87461), .B(n87462), .Z(n85463) );
  NOR U105278 ( .A(n85464), .B(n85463), .Z(n85475) );
  IV U105279 ( .A(n85465), .Z(n85472) );
  NOR U105280 ( .A(n85467), .B(n85466), .Z(n85468) );
  IV U105281 ( .A(n85468), .Z(n85469) );
  NOR U105282 ( .A(n85470), .B(n85469), .Z(n85471) );
  IV U105283 ( .A(n85471), .Z(n85480) );
  NOR U105284 ( .A(n85472), .B(n85480), .Z(n85477) );
  IV U105285 ( .A(n85477), .Z(n85473) );
  NOR U105286 ( .A(n85475), .B(n85473), .Z(n91275) );
  NOR U105287 ( .A(n87462), .B(n85474), .Z(n91276) );
  NOR U105288 ( .A(n85475), .B(n91276), .Z(n85476) );
  NOR U105289 ( .A(n85477), .B(n85476), .Z(n85478) );
  NOR U105290 ( .A(n91275), .B(n85478), .Z(n91268) );
  IV U105291 ( .A(n85479), .Z(n85481) );
  NOR U105292 ( .A(n85481), .B(n85480), .Z(n85482) );
  IV U105293 ( .A(n85482), .Z(n91269) );
  XOR U105294 ( .A(n91268), .B(n91269), .Z(n91271) );
  XOR U105295 ( .A(n91272), .B(n91271), .Z(n87450) );
  XOR U105296 ( .A(n87452), .B(n87450), .Z(n87399) );
  XOR U105297 ( .A(n85483), .B(n87399), .Z(n87394) );
  XOR U105298 ( .A(n87395), .B(n87394), .Z(n87405) );
  IV U105299 ( .A(n85484), .Z(n85485) );
  NOR U105300 ( .A(n85486), .B(n85485), .Z(n87404) );
  IV U105301 ( .A(n85487), .Z(n85488) );
  NOR U105302 ( .A(n85489), .B(n85488), .Z(n87392) );
  NOR U105303 ( .A(n87404), .B(n87392), .Z(n85490) );
  XOR U105304 ( .A(n87405), .B(n85490), .Z(n87408) );
  XOR U105305 ( .A(n85491), .B(n87408), .Z(n87426) );
  XOR U105306 ( .A(n85492), .B(n87426), .Z(n87421) );
  XOR U105307 ( .A(n87422), .B(n87421), .Z(n85493) );
  IV U105308 ( .A(n85493), .Z(n87435) );
  NOR U105309 ( .A(n87438), .B(n87435), .Z(n85500) );
  NOR U105310 ( .A(n85494), .B(n85493), .Z(n85498) );
  IV U105311 ( .A(n85495), .Z(n85508) );
  IV U105312 ( .A(n85496), .Z(n85497) );
  NOR U105313 ( .A(n85508), .B(n85497), .Z(n87437) );
  XOR U105314 ( .A(n85498), .B(n87437), .Z(n85499) );
  NOR U105315 ( .A(n85500), .B(n85499), .Z(n87432) );
  IV U105316 ( .A(n85501), .Z(n85503) );
  NOR U105317 ( .A(n85503), .B(n85502), .Z(n91290) );
  NOR U105318 ( .A(n85505), .B(n85504), .Z(n85506) );
  IV U105319 ( .A(n85506), .Z(n85507) );
  NOR U105320 ( .A(n85508), .B(n85507), .Z(n87433) );
  NOR U105321 ( .A(n91290), .B(n87433), .Z(n85509) );
  XOR U105322 ( .A(n87432), .B(n85509), .Z(n91300) );
  XOR U105323 ( .A(n85510), .B(n91300), .Z(n85511) );
  IV U105324 ( .A(n85511), .Z(n91303) );
  IV U105325 ( .A(n85512), .Z(n85514) );
  NOR U105326 ( .A(n85514), .B(n85513), .Z(n85515) );
  IV U105327 ( .A(n85515), .Z(n91302) );
  XOR U105328 ( .A(n91303), .B(n91302), .Z(n85516) );
  NOR U105329 ( .A(n85517), .B(n85516), .Z(n85520) );
  IV U105330 ( .A(n85517), .Z(n85519) );
  XOR U105331 ( .A(n91293), .B(n91300), .Z(n85518) );
  NOR U105332 ( .A(n85519), .B(n85518), .Z(n91289) );
  NOR U105333 ( .A(n85520), .B(n91289), .Z(n91285) );
  NOR U105334 ( .A(n85522), .B(n85521), .Z(n85523) );
  IV U105335 ( .A(n85523), .Z(n91287) );
  XOR U105336 ( .A(n91285), .B(n91287), .Z(n87339) );
  XOR U105337 ( .A(n87338), .B(n87339), .Z(n87342) );
  XOR U105338 ( .A(n87341), .B(n87342), .Z(n87349) );
  XOR U105339 ( .A(n87348), .B(n87349), .Z(n87352) );
  XOR U105340 ( .A(n87351), .B(n87352), .Z(n87332) );
  XOR U105341 ( .A(n87331), .B(n87332), .Z(n87335) );
  XOR U105342 ( .A(n87334), .B(n87335), .Z(n87368) );
  XOR U105343 ( .A(n87366), .B(n87368), .Z(n87381) );
  XOR U105344 ( .A(n85524), .B(n87381), .Z(n87384) );
  XOR U105345 ( .A(n87386), .B(n87384), .Z(n87378) );
  IV U105346 ( .A(n85525), .Z(n85526) );
  NOR U105347 ( .A(n85527), .B(n85526), .Z(n85531) );
  NOR U105348 ( .A(n85529), .B(n85528), .Z(n85530) );
  NOR U105349 ( .A(n85531), .B(n85530), .Z(n87379) );
  XOR U105350 ( .A(n87378), .B(n87379), .Z(n85532) );
  IV U105351 ( .A(n85532), .Z(n87358) );
  NOR U105352 ( .A(n87361), .B(n87358), .Z(n85539) );
  NOR U105353 ( .A(n85533), .B(n85532), .Z(n85537) );
  IV U105354 ( .A(n85534), .Z(n85536) );
  NOR U105355 ( .A(n85536), .B(n85535), .Z(n87360) );
  XOR U105356 ( .A(n85537), .B(n87360), .Z(n85538) );
  NOR U105357 ( .A(n85539), .B(n85538), .Z(n91315) );
  XOR U105358 ( .A(n91317), .B(n91315), .Z(n91329) );
  XOR U105359 ( .A(n85540), .B(n91329), .Z(n91324) );
  XOR U105360 ( .A(n91326), .B(n91324), .Z(n91336) );
  XOR U105361 ( .A(n91334), .B(n91336), .Z(n91339) );
  XOR U105362 ( .A(n91337), .B(n91339), .Z(n91332) );
  XOR U105363 ( .A(n91333), .B(n91332), .Z(n91350) );
  XOR U105364 ( .A(n91352), .B(n91350), .Z(n91378) );
  XOR U105365 ( .A(n85541), .B(n91378), .Z(n91373) );
  XOR U105366 ( .A(n91374), .B(n91373), .Z(n91361) );
  XOR U105367 ( .A(n91360), .B(n91361), .Z(n91365) );
  XOR U105368 ( .A(n91363), .B(n91365), .Z(n91358) );
  XOR U105369 ( .A(n91357), .B(n91358), .Z(n87300) );
  XOR U105370 ( .A(n87299), .B(n87300), .Z(n87303) );
  XOR U105371 ( .A(n87302), .B(n87303), .Z(n87292) );
  XOR U105372 ( .A(n87291), .B(n87292), .Z(n87295) );
  XOR U105373 ( .A(n87294), .B(n87295), .Z(n87289) );
  XOR U105374 ( .A(n87288), .B(n87289), .Z(n91394) );
  XOR U105375 ( .A(n91395), .B(n91394), .Z(n85542) );
  IV U105376 ( .A(n85542), .Z(n91398) );
  IV U105377 ( .A(n85543), .Z(n85545) );
  NOR U105378 ( .A(n85545), .B(n85544), .Z(n85546) );
  IV U105379 ( .A(n85546), .Z(n85551) );
  NOR U105380 ( .A(n85548), .B(n85547), .Z(n85549) );
  IV U105381 ( .A(n85549), .Z(n85550) );
  NOR U105382 ( .A(n85551), .B(n85550), .Z(n91396) );
  XOR U105383 ( .A(n91398), .B(n91396), .Z(n87321) );
  IV U105384 ( .A(n85552), .Z(n85557) );
  IV U105385 ( .A(n85553), .Z(n85554) );
  NOR U105386 ( .A(n85554), .B(n85559), .Z(n85555) );
  IV U105387 ( .A(n85555), .Z(n85556) );
  NOR U105388 ( .A(n85557), .B(n85556), .Z(n87319) );
  XOR U105389 ( .A(n87321), .B(n87319), .Z(n87324) );
  IV U105390 ( .A(n85558), .Z(n85560) );
  NOR U105391 ( .A(n85560), .B(n85559), .Z(n87322) );
  XOR U105392 ( .A(n87324), .B(n87322), .Z(n87313) );
  IV U105393 ( .A(n85561), .Z(n85562) );
  NOR U105394 ( .A(n85563), .B(n85562), .Z(n87311) );
  XOR U105395 ( .A(n87313), .B(n87311), .Z(n87315) );
  XOR U105396 ( .A(n87314), .B(n87315), .Z(n91408) );
  IV U105397 ( .A(n91408), .Z(n91405) );
  NOR U105398 ( .A(n85565), .B(n85564), .Z(n91406) );
  XOR U105399 ( .A(n91405), .B(n91406), .Z(n85572) );
  IV U105400 ( .A(n85566), .Z(n85567) );
  NOR U105401 ( .A(n85568), .B(n85567), .Z(n91409) );
  NOR U105402 ( .A(n85570), .B(n85569), .Z(n91410) );
  NOR U105403 ( .A(n91409), .B(n91410), .Z(n85571) );
  XOR U105404 ( .A(n85572), .B(n85571), .Z(n91388) );
  IV U105405 ( .A(n85576), .Z(n85574) );
  NOR U105406 ( .A(n85574), .B(n85573), .Z(n85584) );
  NOR U105407 ( .A(n85576), .B(n85575), .Z(n85582) );
  IV U105408 ( .A(n85577), .Z(n85578) );
  NOR U105409 ( .A(n85579), .B(n85578), .Z(n85580) );
  IV U105410 ( .A(n85580), .Z(n85581) );
  NOR U105411 ( .A(n85582), .B(n85581), .Z(n85583) );
  NOR U105412 ( .A(n85584), .B(n85583), .Z(n91387) );
  XOR U105413 ( .A(n91388), .B(n91387), .Z(n91389) );
  XOR U105414 ( .A(n91391), .B(n91389), .Z(n91429) );
  IV U105415 ( .A(n85585), .Z(n85592) );
  NOR U105416 ( .A(n85587), .B(n85586), .Z(n85588) );
  IV U105417 ( .A(n85588), .Z(n85589) );
  NOR U105418 ( .A(n85590), .B(n85589), .Z(n85591) );
  IV U105419 ( .A(n85591), .Z(n85594) );
  NOR U105420 ( .A(n85592), .B(n85594), .Z(n91427) );
  XOR U105421 ( .A(n91429), .B(n91427), .Z(n91432) );
  IV U105422 ( .A(n85593), .Z(n85595) );
  NOR U105423 ( .A(n85595), .B(n85594), .Z(n91430) );
  XOR U105424 ( .A(n91432), .B(n91430), .Z(n91420) );
  XOR U105425 ( .A(n91421), .B(n91420), .Z(n91422) );
  XOR U105426 ( .A(n91424), .B(n91422), .Z(n91418) );
  XOR U105427 ( .A(n91417), .B(n91418), .Z(n87260) );
  IV U105428 ( .A(n85596), .Z(n85598) );
  NOR U105429 ( .A(n85598), .B(n85597), .Z(n87258) );
  XOR U105430 ( .A(n87260), .B(n87258), .Z(n87262) );
  XOR U105431 ( .A(n87261), .B(n87262), .Z(n87251) );
  IV U105432 ( .A(n85599), .Z(n85601) );
  NOR U105433 ( .A(n85601), .B(n85600), .Z(n85602) );
  IV U105434 ( .A(n85602), .Z(n87250) );
  XOR U105435 ( .A(n87251), .B(n87250), .Z(n85603) );
  NOR U105436 ( .A(n85604), .B(n85603), .Z(n87253) );
  IV U105437 ( .A(n85604), .Z(n85605) );
  NOR U105438 ( .A(n85605), .B(n87251), .Z(n87255) );
  NOR U105439 ( .A(n87253), .B(n87255), .Z(n85606) );
  XOR U105440 ( .A(n87252), .B(n85606), .Z(n87269) );
  IV U105441 ( .A(n87269), .Z(n87271) );
  IV U105442 ( .A(n85607), .Z(n85609) );
  NOR U105443 ( .A(n85609), .B(n85608), .Z(n85613) );
  NOR U105444 ( .A(n85611), .B(n85610), .Z(n85612) );
  NOR U105445 ( .A(n85613), .B(n85612), .Z(n87268) );
  IV U105446 ( .A(n87268), .Z(n87270) );
  XOR U105447 ( .A(n87271), .B(n87270), .Z(n85614) );
  XOR U105448 ( .A(n87272), .B(n85614), .Z(n87275) );
  IV U105449 ( .A(n85615), .Z(n85616) );
  NOR U105450 ( .A(n85617), .B(n85616), .Z(n87274) );
  XOR U105451 ( .A(n87275), .B(n87274), .Z(n87277) );
  XOR U105452 ( .A(n87276), .B(n87277), .Z(n85618) );
  NOR U105453 ( .A(n85619), .B(n85618), .Z(n87283) );
  IV U105454 ( .A(n85620), .Z(n85622) );
  NOR U105455 ( .A(n85622), .B(n85621), .Z(n87273) );
  NOR U105456 ( .A(n87276), .B(n87273), .Z(n85623) );
  XOR U105457 ( .A(n85623), .B(n87277), .Z(n87279) );
  NOR U105458 ( .A(n85624), .B(n87279), .Z(n85625) );
  NOR U105459 ( .A(n87283), .B(n85625), .Z(n87218) );
  IV U105460 ( .A(n85626), .Z(n85627) );
  NOR U105461 ( .A(n85633), .B(n85627), .Z(n87278) );
  IV U105462 ( .A(n85628), .Z(n85630) );
  NOR U105463 ( .A(n85630), .B(n85629), .Z(n87217) );
  NOR U105464 ( .A(n87278), .B(n87217), .Z(n85631) );
  XOR U105465 ( .A(n87218), .B(n85631), .Z(n87237) );
  IV U105466 ( .A(n85632), .Z(n85634) );
  NOR U105467 ( .A(n85634), .B(n85633), .Z(n87235) );
  XOR U105468 ( .A(n87237), .B(n87235), .Z(n87238) );
  XOR U105469 ( .A(n87239), .B(n87238), .Z(n85635) );
  IV U105470 ( .A(n85635), .Z(n87244) );
  NOR U105471 ( .A(n87247), .B(n87244), .Z(n85641) );
  NOR U105472 ( .A(n87243), .B(n85635), .Z(n85639) );
  IV U105473 ( .A(n85636), .Z(n85638) );
  NOR U105474 ( .A(n85638), .B(n85637), .Z(n87242) );
  XOR U105475 ( .A(n85639), .B(n87242), .Z(n85640) );
  NOR U105476 ( .A(n85641), .B(n85640), .Z(n87207) );
  IV U105477 ( .A(n85642), .Z(n85644) );
  NOR U105478 ( .A(n85644), .B(n85643), .Z(n85645) );
  IV U105479 ( .A(n85645), .Z(n87208) );
  XOR U105480 ( .A(n87207), .B(n87208), .Z(n87212) );
  XOR U105481 ( .A(n87210), .B(n87212), .Z(n87200) );
  XOR U105482 ( .A(n87199), .B(n87200), .Z(n87203) );
  XOR U105483 ( .A(n87202), .B(n87203), .Z(n87223) );
  XOR U105484 ( .A(n87221), .B(n87223), .Z(n87228) );
  XOR U105485 ( .A(n87229), .B(n87228), .Z(n87224) );
  XOR U105486 ( .A(n87226), .B(n87224), .Z(n91455) );
  XOR U105487 ( .A(n91453), .B(n91455), .Z(n91456) );
  XOR U105488 ( .A(n91457), .B(n91456), .Z(n91460) );
  IV U105489 ( .A(n85646), .Z(n85647) );
  NOR U105490 ( .A(n85648), .B(n85647), .Z(n85650) );
  NOR U105491 ( .A(n85650), .B(n85649), .Z(n91462) );
  XOR U105492 ( .A(n91460), .B(n91462), .Z(n91470) );
  XOR U105493 ( .A(n91471), .B(n91470), .Z(n91467) );
  XOR U105494 ( .A(n91469), .B(n91467), .Z(n87198) );
  XOR U105495 ( .A(n85651), .B(n87198), .Z(n87150) );
  IV U105496 ( .A(n87150), .Z(n87153) );
  XOR U105497 ( .A(n87152), .B(n87153), .Z(n85655) );
  NOR U105498 ( .A(n85653), .B(n85652), .Z(n87154) );
  NOR U105499 ( .A(n87154), .B(n87155), .Z(n85654) );
  XOR U105500 ( .A(n85655), .B(n85654), .Z(n87178) );
  IV U105501 ( .A(n85656), .Z(n85659) );
  IV U105502 ( .A(n85657), .Z(n85658) );
  NOR U105503 ( .A(n85659), .B(n85658), .Z(n87176) );
  XOR U105504 ( .A(n87178), .B(n87176), .Z(n87181) );
  XOR U105505 ( .A(n87179), .B(n87181), .Z(n87167) );
  XOR U105506 ( .A(n87168), .B(n87167), .Z(n87169) );
  NOR U105507 ( .A(n85661), .B(n85660), .Z(n85663) );
  NOR U105508 ( .A(n85663), .B(n85662), .Z(n85664) );
  IV U105509 ( .A(n85664), .Z(n87170) );
  XOR U105510 ( .A(n87169), .B(n87170), .Z(n87161) );
  XOR U105511 ( .A(n87160), .B(n87161), .Z(n87163) );
  IV U105512 ( .A(n85665), .Z(n85666) );
  NOR U105513 ( .A(n85667), .B(n85666), .Z(n85668) );
  NOR U105514 ( .A(n85669), .B(n85668), .Z(n87164) );
  XOR U105515 ( .A(n87163), .B(n87164), .Z(n91515) );
  XOR U105516 ( .A(n91516), .B(n91515), .Z(n87193) );
  XOR U105517 ( .A(n85670), .B(n87193), .Z(n87188) );
  XOR U105518 ( .A(n85671), .B(n87188), .Z(n91493) );
  XOR U105519 ( .A(n91492), .B(n91493), .Z(n91501) );
  XOR U105520 ( .A(n91499), .B(n91501), .Z(n91507) );
  XOR U105521 ( .A(n91506), .B(n91507), .Z(n91504) );
  XOR U105522 ( .A(n91502), .B(n91504), .Z(n91537) );
  XOR U105523 ( .A(n91536), .B(n91537), .Z(n91540) );
  XOR U105524 ( .A(n91539), .B(n91540), .Z(n91535) );
  XOR U105525 ( .A(n91534), .B(n91535), .Z(n91527) );
  XOR U105526 ( .A(n91529), .B(n91527), .Z(n87117) );
  XOR U105527 ( .A(n85672), .B(n87117), .Z(n87109) );
  XOR U105528 ( .A(n85673), .B(n87109), .Z(n87122) );
  XOR U105529 ( .A(n87123), .B(n87122), .Z(n87124) );
  IV U105530 ( .A(n85674), .Z(n85676) );
  NOR U105531 ( .A(n85676), .B(n85675), .Z(n85677) );
  IV U105532 ( .A(n85677), .Z(n87125) );
  XOR U105533 ( .A(n87124), .B(n87125), .Z(n87139) );
  XOR U105534 ( .A(n87138), .B(n87139), .Z(n87143) );
  NOR U105535 ( .A(n85679), .B(n85678), .Z(n85685) );
  IV U105536 ( .A(n85679), .Z(n85680) );
  NOR U105537 ( .A(n85681), .B(n85680), .Z(n85682) );
  NOR U105538 ( .A(n85683), .B(n85682), .Z(n85684) );
  NOR U105539 ( .A(n85685), .B(n85684), .Z(n87141) );
  XOR U105540 ( .A(n87143), .B(n87141), .Z(n87132) );
  XOR U105541 ( .A(n87131), .B(n87132), .Z(n87134) );
  IV U105542 ( .A(n85686), .Z(n85687) );
  NOR U105543 ( .A(n85688), .B(n85687), .Z(n85693) );
  IV U105544 ( .A(n85689), .Z(n85691) );
  NOR U105545 ( .A(n85691), .B(n85690), .Z(n85692) );
  NOR U105546 ( .A(n85693), .B(n85692), .Z(n87135) );
  XOR U105547 ( .A(n87134), .B(n87135), .Z(n87101) );
  XOR U105548 ( .A(n87103), .B(n87101), .Z(n87105) );
  XOR U105549 ( .A(n87085), .B(n87105), .Z(n85697) );
  IV U105550 ( .A(n85694), .Z(n85695) );
  NOR U105551 ( .A(n85696), .B(n85695), .Z(n87104) );
  XOR U105552 ( .A(n85697), .B(n87104), .Z(n85698) );
  NOR U105553 ( .A(n87082), .B(n85698), .Z(n85702) );
  IV U105554 ( .A(n87082), .Z(n87083) );
  IV U105555 ( .A(n87105), .Z(n87080) );
  NOR U105556 ( .A(n87085), .B(n87080), .Z(n85699) );
  IV U105557 ( .A(n85699), .Z(n85700) );
  NOR U105558 ( .A(n87083), .B(n85700), .Z(n85701) );
  NOR U105559 ( .A(n85702), .B(n85701), .Z(n87092) );
  XOR U105560 ( .A(n85703), .B(n87092), .Z(n87095) );
  XOR U105561 ( .A(n87094), .B(n87095), .Z(n87090) );
  XOR U105562 ( .A(n87089), .B(n87090), .Z(n87051) );
  IV U105563 ( .A(n85704), .Z(n85706) );
  NOR U105564 ( .A(n85706), .B(n85705), .Z(n87088) );
  IV U105565 ( .A(n85707), .Z(n85708) );
  NOR U105566 ( .A(n85712), .B(n85708), .Z(n87049) );
  NOR U105567 ( .A(n87088), .B(n87049), .Z(n85709) );
  XOR U105568 ( .A(n87051), .B(n85709), .Z(n85710) );
  IV U105569 ( .A(n85710), .Z(n87056) );
  IV U105570 ( .A(n85711), .Z(n85713) );
  NOR U105571 ( .A(n85713), .B(n85712), .Z(n87047) );
  IV U105572 ( .A(n85714), .Z(n85716) );
  NOR U105573 ( .A(n85716), .B(n85715), .Z(n87054) );
  NOR U105574 ( .A(n87047), .B(n87054), .Z(n85717) );
  XOR U105575 ( .A(n87056), .B(n85717), .Z(n87057) );
  IV U105576 ( .A(n85718), .Z(n85719) );
  NOR U105577 ( .A(n85720), .B(n85719), .Z(n85730) );
  IV U105578 ( .A(n85730), .Z(n87059) );
  NOR U105579 ( .A(n87057), .B(n87059), .Z(n85732) );
  IV U105580 ( .A(n85721), .Z(n85722) );
  NOR U105581 ( .A(n85723), .B(n85722), .Z(n85726) );
  IV U105582 ( .A(n85726), .Z(n85725) );
  XOR U105583 ( .A(n87047), .B(n87056), .Z(n85724) );
  NOR U105584 ( .A(n85725), .B(n85724), .Z(n87064) );
  NOR U105585 ( .A(n87057), .B(n85726), .Z(n85727) );
  NOR U105586 ( .A(n87064), .B(n85727), .Z(n85728) );
  IV U105587 ( .A(n85728), .Z(n85729) );
  NOR U105588 ( .A(n85730), .B(n85729), .Z(n85731) );
  NOR U105589 ( .A(n85732), .B(n85731), .Z(n87068) );
  XOR U105590 ( .A(n87067), .B(n87068), .Z(n87071) );
  XOR U105591 ( .A(n87070), .B(n87071), .Z(n91563) );
  XOR U105592 ( .A(n91564), .B(n91563), .Z(n91565) );
  IV U105593 ( .A(n85733), .Z(n85735) );
  NOR U105594 ( .A(n85735), .B(n85734), .Z(n85736) );
  IV U105595 ( .A(n85736), .Z(n91566) );
  XOR U105596 ( .A(n91565), .B(n91566), .Z(n91568) );
  IV U105597 ( .A(n85737), .Z(n85738) );
  NOR U105598 ( .A(n85739), .B(n85738), .Z(n85744) );
  IV U105599 ( .A(n85740), .Z(n85741) );
  NOR U105600 ( .A(n85742), .B(n85741), .Z(n85743) );
  NOR U105601 ( .A(n85744), .B(n85743), .Z(n91569) );
  XOR U105602 ( .A(n91568), .B(n91569), .Z(n85745) );
  IV U105603 ( .A(n85745), .Z(n87078) );
  XOR U105604 ( .A(n87077), .B(n87078), .Z(n91582) );
  XOR U105605 ( .A(n85746), .B(n91582), .Z(n85749) );
  XOR U105606 ( .A(n91578), .B(n85749), .Z(n85747) );
  NOR U105607 ( .A(n85748), .B(n85747), .Z(n91598) );
  IV U105608 ( .A(n85749), .Z(n91595) );
  IV U105609 ( .A(n85750), .Z(n85752) );
  NOR U105610 ( .A(n85752), .B(n85751), .Z(n91594) );
  NOR U105611 ( .A(n85753), .B(n91594), .Z(n85754) );
  XOR U105612 ( .A(n91595), .B(n85754), .Z(n85755) );
  NOR U105613 ( .A(n85756), .B(n85755), .Z(n85757) );
  NOR U105614 ( .A(n91598), .B(n85757), .Z(n91591) );
  IV U105615 ( .A(n85758), .Z(n85760) );
  NOR U105616 ( .A(n85760), .B(n85759), .Z(n85767) );
  IV U105617 ( .A(n85761), .Z(n85765) );
  NOR U105618 ( .A(n85763), .B(n85762), .Z(n85764) );
  IV U105619 ( .A(n85764), .Z(n85769) );
  NOR U105620 ( .A(n85765), .B(n85769), .Z(n85766) );
  NOR U105621 ( .A(n85767), .B(n85766), .Z(n91593) );
  XOR U105622 ( .A(n91591), .B(n91593), .Z(n87025) );
  IV U105623 ( .A(n85768), .Z(n85770) );
  NOR U105624 ( .A(n85770), .B(n85769), .Z(n87023) );
  XOR U105625 ( .A(n87025), .B(n87023), .Z(n87028) );
  NOR U105626 ( .A(n85772), .B(n85771), .Z(n87026) );
  XOR U105627 ( .A(n87028), .B(n87026), .Z(n87010) );
  IV U105628 ( .A(n87010), .Z(n87012) );
  XOR U105629 ( .A(n87011), .B(n87012), .Z(n85778) );
  IV U105630 ( .A(n85773), .Z(n85775) );
  NOR U105631 ( .A(n85775), .B(n85774), .Z(n85776) );
  NOR U105632 ( .A(n87016), .B(n85776), .Z(n85777) );
  XOR U105633 ( .A(n85778), .B(n85777), .Z(n87006) );
  IV U105634 ( .A(n85779), .Z(n85781) );
  IV U105635 ( .A(n85780), .Z(n87014) );
  NOR U105636 ( .A(n85781), .B(n87014), .Z(n87007) );
  IV U105637 ( .A(n85782), .Z(n85783) );
  NOR U105638 ( .A(n87014), .B(n85783), .Z(n85784) );
  NOR U105639 ( .A(n87007), .B(n85784), .Z(n85785) );
  XOR U105640 ( .A(n87006), .B(n85785), .Z(n87036) );
  XOR U105641 ( .A(n87037), .B(n87036), .Z(n87033) );
  IV U105642 ( .A(n85786), .Z(n85787) );
  NOR U105643 ( .A(n85788), .B(n85787), .Z(n85789) );
  NOR U105644 ( .A(n85790), .B(n85789), .Z(n87035) );
  XOR U105645 ( .A(n87033), .B(n87035), .Z(n87039) );
  XOR U105646 ( .A(n87038), .B(n87039), .Z(n91630) );
  XOR U105647 ( .A(n91629), .B(n91630), .Z(n91633) );
  XOR U105648 ( .A(n91632), .B(n91633), .Z(n91617) );
  XOR U105649 ( .A(n91616), .B(n91617), .Z(n91619) );
  XOR U105650 ( .A(n91620), .B(n91619), .Z(n85791) );
  IV U105651 ( .A(n85791), .Z(n91609) );
  XOR U105652 ( .A(n91608), .B(n91609), .Z(n91613) );
  IV U105653 ( .A(n85792), .Z(n85794) );
  NOR U105654 ( .A(n85794), .B(n85793), .Z(n91611) );
  XOR U105655 ( .A(n91613), .B(n91611), .Z(n91642) );
  IV U105656 ( .A(n91642), .Z(n91639) );
  IV U105657 ( .A(n85795), .Z(n85797) );
  NOR U105658 ( .A(n85797), .B(n85796), .Z(n91640) );
  XOR U105659 ( .A(n91639), .B(n91640), .Z(n85807) );
  IV U105660 ( .A(n85798), .Z(n85801) );
  NOR U105661 ( .A(n85809), .B(n85799), .Z(n85800) );
  IV U105662 ( .A(n85800), .Z(n85804) );
  NOR U105663 ( .A(n85801), .B(n85804), .Z(n91644) );
  NOR U105664 ( .A(n85803), .B(n85802), .Z(n85805) );
  NOR U105665 ( .A(n85805), .B(n85804), .Z(n91643) );
  NOR U105666 ( .A(n91644), .B(n91643), .Z(n85806) );
  XOR U105667 ( .A(n85807), .B(n85806), .Z(n87001) );
  NOR U105668 ( .A(n85809), .B(n85808), .Z(n86999) );
  XOR U105669 ( .A(n87001), .B(n86999), .Z(n87002) );
  XOR U105670 ( .A(n87003), .B(n87002), .Z(n86979) );
  IV U105671 ( .A(n86979), .Z(n86982) );
  XOR U105672 ( .A(n86980), .B(n86982), .Z(n85810) );
  XOR U105673 ( .A(n85811), .B(n85810), .Z(n86991) );
  XOR U105674 ( .A(n86989), .B(n86991), .Z(n86993) );
  XOR U105675 ( .A(n86992), .B(n86993), .Z(n91670) );
  XOR U105676 ( .A(n91671), .B(n91670), .Z(n85812) );
  IV U105677 ( .A(n85812), .Z(n91673) );
  XOR U105678 ( .A(n85813), .B(n91673), .Z(n91660) );
  IV U105679 ( .A(n85814), .Z(n85815) );
  NOR U105680 ( .A(n85815), .B(n85817), .Z(n85825) );
  IV U105681 ( .A(n85825), .Z(n91661) );
  NOR U105682 ( .A(n91660), .B(n91661), .Z(n85827) );
  XOR U105683 ( .A(n91672), .B(n91673), .Z(n85820) );
  IV U105684 ( .A(n85816), .Z(n85818) );
  NOR U105685 ( .A(n85818), .B(n85817), .Z(n85821) );
  IV U105686 ( .A(n85821), .Z(n85819) );
  NOR U105687 ( .A(n85820), .B(n85819), .Z(n91664) );
  NOR U105688 ( .A(n91660), .B(n85821), .Z(n85822) );
  NOR U105689 ( .A(n91664), .B(n85822), .Z(n85823) );
  IV U105690 ( .A(n85823), .Z(n85824) );
  NOR U105691 ( .A(n85825), .B(n85824), .Z(n85826) );
  NOR U105692 ( .A(n85827), .B(n85826), .Z(n91659) );
  XOR U105693 ( .A(n91657), .B(n91659), .Z(n86956) );
  XOR U105694 ( .A(n85828), .B(n86956), .Z(n86958) );
  IV U105695 ( .A(n85829), .Z(n85831) );
  NOR U105696 ( .A(n85831), .B(n85830), .Z(n86959) );
  XOR U105697 ( .A(n86958), .B(n86959), .Z(n86947) );
  IV U105698 ( .A(n85832), .Z(n85833) );
  NOR U105699 ( .A(n85834), .B(n85833), .Z(n85837) );
  NOR U105700 ( .A(n85835), .B(n85842), .Z(n85836) );
  NOR U105701 ( .A(n85837), .B(n85836), .Z(n86949) );
  XOR U105702 ( .A(n86947), .B(n86949), .Z(n86952) );
  XOR U105703 ( .A(n86950), .B(n86952), .Z(n91686) );
  XOR U105704 ( .A(n91685), .B(n91686), .Z(n91689) );
  IV U105705 ( .A(n85838), .Z(n85839) );
  NOR U105706 ( .A(n85840), .B(n85839), .Z(n91688) );
  IV U105707 ( .A(n85841), .Z(n85847) );
  XOR U105708 ( .A(n85843), .B(n85842), .Z(n85844) );
  XOR U105709 ( .A(n85845), .B(n85844), .Z(n85846) );
  NOR U105710 ( .A(n85847), .B(n85846), .Z(n91683) );
  NOR U105711 ( .A(n91688), .B(n91683), .Z(n85848) );
  XOR U105712 ( .A(n91689), .B(n85848), .Z(n85849) );
  NOR U105713 ( .A(n85852), .B(n85849), .Z(n85857) );
  IV U105714 ( .A(n85850), .Z(n85851) );
  NOR U105715 ( .A(n85866), .B(n85851), .Z(n85859) );
  XOR U105716 ( .A(n91683), .B(n91689), .Z(n85854) );
  IV U105717 ( .A(n85852), .Z(n85853) );
  NOR U105718 ( .A(n85854), .B(n85853), .Z(n85855) );
  NOR U105719 ( .A(n85859), .B(n85855), .Z(n85856) );
  NOR U105720 ( .A(n85857), .B(n85856), .Z(n86976) );
  IV U105721 ( .A(n85857), .Z(n85858) );
  NOR U105722 ( .A(n85859), .B(n85858), .Z(n85860) );
  NOR U105723 ( .A(n86976), .B(n85860), .Z(n86968) );
  IV U105724 ( .A(n85861), .Z(n85862) );
  NOR U105725 ( .A(n85863), .B(n85862), .Z(n85868) );
  IV U105726 ( .A(n85864), .Z(n85865) );
  NOR U105727 ( .A(n85866), .B(n85865), .Z(n85867) );
  NOR U105728 ( .A(n85868), .B(n85867), .Z(n86970) );
  XOR U105729 ( .A(n86968), .B(n86970), .Z(n86972) );
  XOR U105730 ( .A(n86971), .B(n86972), .Z(n85876) );
  IV U105731 ( .A(n85876), .Z(n85869) );
  NOR U105732 ( .A(n85870), .B(n85869), .Z(n85874) );
  IV U105733 ( .A(n85877), .Z(n85872) );
  NOR U105734 ( .A(n85872), .B(n85871), .Z(n85873) );
  NOR U105735 ( .A(n85874), .B(n85873), .Z(n85875) );
  IV U105736 ( .A(n85875), .Z(n86930) );
  NOR U105737 ( .A(n85877), .B(n85876), .Z(n85878) );
  IV U105738 ( .A(n85878), .Z(n85879) );
  NOR U105739 ( .A(n85880), .B(n85879), .Z(n86932) );
  NOR U105740 ( .A(n86930), .B(n86932), .Z(n85881) );
  XOR U105741 ( .A(n85882), .B(n85881), .Z(n85883) );
  XOR U105742 ( .A(n86920), .B(n85883), .Z(n86934) );
  IV U105743 ( .A(n85884), .Z(n85885) );
  NOR U105744 ( .A(n85886), .B(n85885), .Z(n85891) );
  IV U105745 ( .A(n85887), .Z(n85888) );
  NOR U105746 ( .A(n85889), .B(n85888), .Z(n85890) );
  NOR U105747 ( .A(n85891), .B(n85890), .Z(n86933) );
  XOR U105748 ( .A(n86934), .B(n86933), .Z(n86937) );
  NOR U105749 ( .A(n86936), .B(n86937), .Z(n85895) );
  NOR U105750 ( .A(n85895), .B(n85896), .Z(n86942) );
  IV U105751 ( .A(n85896), .Z(n85898) );
  XOR U105752 ( .A(n86937), .B(n86936), .Z(n85897) );
  NOR U105753 ( .A(n85898), .B(n85897), .Z(n85899) );
  NOR U105754 ( .A(n86942), .B(n85899), .Z(n91703) );
  XOR U105755 ( .A(n91703), .B(n91702), .Z(n85900) );
  IV U105756 ( .A(n85900), .Z(n91708) );
  NOR U105757 ( .A(n91711), .B(n91708), .Z(n85903) );
  NOR U105758 ( .A(n91707), .B(n85900), .Z(n85901) );
  XOR U105759 ( .A(n85901), .B(n91706), .Z(n85902) );
  NOR U105760 ( .A(n85903), .B(n85902), .Z(n86910) );
  IV U105761 ( .A(n85904), .Z(n85906) );
  NOR U105762 ( .A(n85906), .B(n85905), .Z(n85907) );
  IV U105763 ( .A(n85907), .Z(n86912) );
  XOR U105764 ( .A(n86910), .B(n86912), .Z(n86914) );
  XOR U105765 ( .A(n86913), .B(n86914), .Z(n86903) );
  XOR U105766 ( .A(n86902), .B(n86903), .Z(n86907) );
  XOR U105767 ( .A(n86905), .B(n86907), .Z(n86891) );
  XOR U105768 ( .A(n85908), .B(n86891), .Z(n86886) );
  NOR U105769 ( .A(n86886), .B(n86888), .Z(n85912) );
  IV U105770 ( .A(n86888), .Z(n85910) );
  XOR U105771 ( .A(n86889), .B(n86891), .Z(n85909) );
  NOR U105772 ( .A(n85910), .B(n85909), .Z(n85911) );
  NOR U105773 ( .A(n85912), .B(n85911), .Z(n86873) );
  XOR U105774 ( .A(n85913), .B(n86873), .Z(n86878) );
  XOR U105775 ( .A(n86876), .B(n86878), .Z(n86879) );
  XOR U105776 ( .A(n86880), .B(n86879), .Z(n86893) );
  XOR U105777 ( .A(n86894), .B(n86893), .Z(n86842) );
  XOR U105778 ( .A(n85914), .B(n86842), .Z(n86833) );
  XOR U105779 ( .A(n86838), .B(n86833), .Z(n86831) );
  IV U105780 ( .A(n85915), .Z(n85916) );
  NOR U105781 ( .A(n85923), .B(n85916), .Z(n86830) );
  IV U105782 ( .A(n85917), .Z(n85919) );
  NOR U105783 ( .A(n85919), .B(n85918), .Z(n86834) );
  NOR U105784 ( .A(n86830), .B(n86834), .Z(n85920) );
  XOR U105785 ( .A(n86831), .B(n85920), .Z(n86854) );
  IV U105786 ( .A(n85921), .Z(n85922) );
  NOR U105787 ( .A(n85923), .B(n85922), .Z(n85924) );
  IV U105788 ( .A(n85924), .Z(n86855) );
  XOR U105789 ( .A(n86854), .B(n86855), .Z(n86858) );
  XOR U105790 ( .A(n86857), .B(n86858), .Z(n86848) );
  XOR U105791 ( .A(n86847), .B(n86848), .Z(n86850) );
  XOR U105792 ( .A(n86851), .B(n86850), .Z(n85925) );
  IV U105793 ( .A(n85925), .Z(n86866) );
  IV U105794 ( .A(n85928), .Z(n85927) );
  NOR U105795 ( .A(n85927), .B(n85926), .Z(n85933) );
  NOR U105796 ( .A(n85929), .B(n85928), .Z(n85930) );
  NOR U105797 ( .A(n85931), .B(n85930), .Z(n85932) );
  NOR U105798 ( .A(n85933), .B(n85932), .Z(n86864) );
  XOR U105799 ( .A(n86866), .B(n86864), .Z(n86777) );
  IV U105800 ( .A(n86777), .Z(n85941) );
  IV U105801 ( .A(n85934), .Z(n85936) );
  NOR U105802 ( .A(n85936), .B(n85935), .Z(n86865) );
  IV U105803 ( .A(n85937), .Z(n85939) );
  NOR U105804 ( .A(n85939), .B(n85938), .Z(n86775) );
  NOR U105805 ( .A(n86865), .B(n86775), .Z(n85940) );
  XOR U105806 ( .A(n85941), .B(n85940), .Z(n86774) );
  XOR U105807 ( .A(n86773), .B(n86774), .Z(n86783) );
  XOR U105808 ( .A(n86784), .B(n86783), .Z(n86769) );
  XOR U105809 ( .A(n85942), .B(n86769), .Z(n86765) );
  XOR U105810 ( .A(n86766), .B(n86765), .Z(n86803) );
  XOR U105811 ( .A(n86802), .B(n86803), .Z(n86805) );
  XOR U105812 ( .A(n86806), .B(n86805), .Z(n86799) );
  XOR U105813 ( .A(n86801), .B(n86799), .Z(n86793) );
  NOR U105814 ( .A(n85943), .B(n86793), .Z(n86814) );
  IV U105815 ( .A(n85944), .Z(n85946) );
  NOR U105816 ( .A(n85946), .B(n85945), .Z(n85947) );
  IV U105817 ( .A(n85947), .Z(n86792) );
  XOR U105818 ( .A(n86793), .B(n86792), .Z(n85948) );
  NOR U105819 ( .A(n85949), .B(n85948), .Z(n86817) );
  NOR U105820 ( .A(n86814), .B(n86817), .Z(n85950) );
  IV U105821 ( .A(n85950), .Z(n86795) );
  IV U105822 ( .A(n85951), .Z(n85953) );
  NOR U105823 ( .A(n85953), .B(n85952), .Z(n86815) );
  IV U105824 ( .A(n85954), .Z(n85956) );
  NOR U105825 ( .A(n85956), .B(n85955), .Z(n86794) );
  NOR U105826 ( .A(n86815), .B(n86794), .Z(n85957) );
  XOR U105827 ( .A(n86795), .B(n85957), .Z(n85960) );
  IV U105828 ( .A(n85960), .Z(n85958) );
  NOR U105829 ( .A(n85959), .B(n85958), .Z(n86755) );
  NOR U105830 ( .A(n85961), .B(n85960), .Z(n86753) );
  XOR U105831 ( .A(n86753), .B(n86752), .Z(n85962) );
  NOR U105832 ( .A(n86755), .B(n85962), .Z(n86758) );
  XOR U105833 ( .A(n86760), .B(n86758), .Z(n86823) );
  XOR U105834 ( .A(n86822), .B(n86823), .Z(n86826) );
  IV U105835 ( .A(n85963), .Z(n85967) );
  NOR U105836 ( .A(n85965), .B(n85964), .Z(n85966) );
  IV U105837 ( .A(n85966), .Z(n85984) );
  NOR U105838 ( .A(n85967), .B(n85984), .Z(n85981) );
  IV U105839 ( .A(n85981), .Z(n85968) );
  NOR U105840 ( .A(n86826), .B(n85968), .Z(n86751) );
  IV U105841 ( .A(n85969), .Z(n85973) );
  IV U105842 ( .A(n85970), .Z(n85979) );
  NOR U105843 ( .A(n85979), .B(n85971), .Z(n85972) );
  IV U105844 ( .A(n85972), .Z(n85976) );
  NOR U105845 ( .A(n85973), .B(n85976), .Z(n85974) );
  IV U105846 ( .A(n85974), .Z(n86749) );
  IV U105847 ( .A(n85975), .Z(n85977) );
  NOR U105848 ( .A(n85977), .B(n85976), .Z(n86729) );
  NOR U105849 ( .A(n85979), .B(n85978), .Z(n86825) );
  XOR U105850 ( .A(n86825), .B(n86826), .Z(n86730) );
  XOR U105851 ( .A(n86729), .B(n86730), .Z(n86748) );
  XOR U105852 ( .A(n86749), .B(n86748), .Z(n85980) );
  NOR U105853 ( .A(n85981), .B(n85980), .Z(n85982) );
  NOR U105854 ( .A(n86751), .B(n85982), .Z(n86722) );
  IV U105855 ( .A(n85983), .Z(n85985) );
  NOR U105856 ( .A(n85985), .B(n85984), .Z(n85986) );
  IV U105857 ( .A(n85986), .Z(n86723) );
  XOR U105858 ( .A(n86722), .B(n86723), .Z(n86725) );
  XOR U105859 ( .A(n86726), .B(n86725), .Z(n86738) );
  XOR U105860 ( .A(n86739), .B(n86738), .Z(n86742) );
  XOR U105861 ( .A(n86741), .B(n86742), .Z(n86732) );
  XOR U105862 ( .A(n86733), .B(n86732), .Z(n91743) );
  XOR U105863 ( .A(n91745), .B(n91743), .Z(n91739) );
  XOR U105864 ( .A(n85987), .B(n91739), .Z(n91734) );
  XOR U105865 ( .A(n91735), .B(n91734), .Z(n91753) );
  XOR U105866 ( .A(n91752), .B(n91753), .Z(n91755) );
  XOR U105867 ( .A(n91756), .B(n91755), .Z(n85988) );
  IV U105868 ( .A(n85988), .Z(n86691) );
  NOR U105869 ( .A(n86694), .B(n86691), .Z(n85995) );
  NOR U105870 ( .A(n85989), .B(n85988), .Z(n85993) );
  IV U105871 ( .A(n85990), .Z(n85992) );
  NOR U105872 ( .A(n85992), .B(n85991), .Z(n86693) );
  XOR U105873 ( .A(n85993), .B(n86693), .Z(n85994) );
  NOR U105874 ( .A(n85995), .B(n85994), .Z(n86688) );
  XOR U105875 ( .A(n86687), .B(n86688), .Z(n86679) );
  XOR U105876 ( .A(n86677), .B(n86679), .Z(n86672) );
  XOR U105877 ( .A(n85996), .B(n86672), .Z(n86668) );
  XOR U105878 ( .A(n86669), .B(n86668), .Z(n86711) );
  XOR U105879 ( .A(n86712), .B(n86711), .Z(n85997) );
  IV U105880 ( .A(n85997), .Z(n86714) );
  XOR U105881 ( .A(n86713), .B(n86714), .Z(n91795) );
  XOR U105882 ( .A(n91796), .B(n91795), .Z(n85998) );
  IV U105883 ( .A(n85998), .Z(n91798) );
  XOR U105884 ( .A(n91797), .B(n91798), .Z(n86706) );
  IV U105885 ( .A(n86706), .Z(n86704) );
  IV U105886 ( .A(n85999), .Z(n86000) );
  NOR U105887 ( .A(n86001), .B(n86000), .Z(n86703) );
  IV U105888 ( .A(n86703), .Z(n86705) );
  XOR U105889 ( .A(n86704), .B(n86705), .Z(n91788) );
  XOR U105890 ( .A(n91787), .B(n91788), .Z(n91785) );
  IV U105891 ( .A(n91785), .Z(n91781) );
  XOR U105892 ( .A(n91784), .B(n91781), .Z(n86002) );
  XOR U105893 ( .A(n86003), .B(n86002), .Z(n91770) );
  IV U105894 ( .A(n86004), .Z(n86006) );
  NOR U105895 ( .A(n86006), .B(n86005), .Z(n91768) );
  XOR U105896 ( .A(n91770), .B(n91768), .Z(n91773) );
  XOR U105897 ( .A(n91771), .B(n91773), .Z(n91767) );
  IV U105898 ( .A(n86007), .Z(n86008) );
  NOR U105899 ( .A(n86009), .B(n86008), .Z(n91765) );
  IV U105900 ( .A(n86010), .Z(n86011) );
  NOR U105901 ( .A(n86012), .B(n86011), .Z(n91766) );
  NOR U105902 ( .A(n91765), .B(n91766), .Z(n86013) );
  XOR U105903 ( .A(n91767), .B(n86013), .Z(n86014) );
  NOR U105904 ( .A(n86024), .B(n86014), .Z(n86029) );
  IV U105905 ( .A(n86015), .Z(n86016) );
  NOR U105906 ( .A(n86017), .B(n86016), .Z(n86022) );
  IV U105907 ( .A(n86018), .Z(n86019) );
  NOR U105908 ( .A(n86020), .B(n86019), .Z(n86021) );
  NOR U105909 ( .A(n86022), .B(n86021), .Z(n86023) );
  IV U105910 ( .A(n86023), .Z(n86031) );
  IV U105911 ( .A(n86024), .Z(n86026) );
  XOR U105912 ( .A(n91765), .B(n91767), .Z(n86025) );
  NOR U105913 ( .A(n86026), .B(n86025), .Z(n86027) );
  NOR U105914 ( .A(n86031), .B(n86027), .Z(n86028) );
  NOR U105915 ( .A(n86029), .B(n86028), .Z(n91827) );
  IV U105916 ( .A(n86029), .Z(n86030) );
  NOR U105917 ( .A(n86031), .B(n86030), .Z(n86032) );
  NOR U105918 ( .A(n91827), .B(n86032), .Z(n86033) );
  IV U105919 ( .A(n86033), .Z(n91813) );
  XOR U105920 ( .A(n91812), .B(n91813), .Z(n91816) );
  XOR U105921 ( .A(n91815), .B(n91816), .Z(n91811) );
  IV U105922 ( .A(n86034), .Z(n86036) );
  NOR U105923 ( .A(n86036), .B(n86035), .Z(n91808) );
  XOR U105924 ( .A(n91811), .B(n91808), .Z(n91824) );
  IV U105925 ( .A(n86037), .Z(n86046) );
  IV U105926 ( .A(n86040), .Z(n86038) );
  NOR U105927 ( .A(n86046), .B(n86038), .Z(n91809) );
  IV U105928 ( .A(n86039), .Z(n86042) );
  XOR U105929 ( .A(n86046), .B(n86040), .Z(n86041) );
  NOR U105930 ( .A(n86042), .B(n86041), .Z(n91823) );
  NOR U105931 ( .A(n91809), .B(n91823), .Z(n86043) );
  XOR U105932 ( .A(n91824), .B(n86043), .Z(n86660) );
  IV U105933 ( .A(n86044), .Z(n86045) );
  NOR U105934 ( .A(n86046), .B(n86045), .Z(n86051) );
  IV U105935 ( .A(n86047), .Z(n86048) );
  NOR U105936 ( .A(n86049), .B(n86048), .Z(n86050) );
  NOR U105937 ( .A(n86051), .B(n86050), .Z(n86661) );
  XOR U105938 ( .A(n86660), .B(n86661), .Z(n86664) );
  XOR U105939 ( .A(n86663), .B(n86664), .Z(n86658) );
  IV U105940 ( .A(n86052), .Z(n86054) );
  NOR U105941 ( .A(n86054), .B(n86053), .Z(n86656) );
  IV U105942 ( .A(n86656), .Z(n86657) );
  XOR U105943 ( .A(n86658), .B(n86657), .Z(n86055) );
  XOR U105944 ( .A(n86659), .B(n86055), .Z(n91850) );
  XOR U105945 ( .A(n91848), .B(n91850), .Z(n91852) );
  XOR U105946 ( .A(n91851), .B(n91852), .Z(n91837) );
  XOR U105947 ( .A(n91835), .B(n91837), .Z(n91840) );
  XOR U105948 ( .A(n86056), .B(n91840), .Z(n86645) );
  XOR U105949 ( .A(n86647), .B(n86645), .Z(n86655) );
  IV U105950 ( .A(n86057), .Z(n86058) );
  NOR U105951 ( .A(n86059), .B(n86058), .Z(n86654) );
  IV U105952 ( .A(n86060), .Z(n86062) );
  NOR U105953 ( .A(n86062), .B(n86061), .Z(n86653) );
  NOR U105954 ( .A(n86654), .B(n86653), .Z(n86063) );
  XOR U105955 ( .A(n86655), .B(n86063), .Z(n86064) );
  NOR U105956 ( .A(n86065), .B(n86064), .Z(n86068) );
  IV U105957 ( .A(n86065), .Z(n86067) );
  XOR U105958 ( .A(n86654), .B(n86655), .Z(n86066) );
  NOR U105959 ( .A(n86067), .B(n86066), .Z(n86652) );
  NOR U105960 ( .A(n86068), .B(n86652), .Z(n86650) );
  NOR U105961 ( .A(n86070), .B(n86069), .Z(n86077) );
  NOR U105962 ( .A(n86072), .B(n86071), .Z(n86075) );
  IV U105963 ( .A(n86073), .Z(n86074) );
  NOR U105964 ( .A(n86075), .B(n86074), .Z(n86076) );
  NOR U105965 ( .A(n86077), .B(n86076), .Z(n86651) );
  XOR U105966 ( .A(n86650), .B(n86651), .Z(n86084) );
  IV U105967 ( .A(n86084), .Z(n86078) );
  NOR U105968 ( .A(n86083), .B(n86078), .Z(n86079) );
  IV U105969 ( .A(n86079), .Z(n86082) );
  IV U105970 ( .A(n86080), .Z(n86081) );
  NOR U105971 ( .A(n86095), .B(n86081), .Z(n86086) );
  NOR U105972 ( .A(n86082), .B(n86086), .Z(n86092) );
  IV U105973 ( .A(n86083), .Z(n86087) );
  XOR U105974 ( .A(n86086), .B(n86087), .Z(n86085) );
  NOR U105975 ( .A(n86085), .B(n86084), .Z(n86090) );
  IV U105976 ( .A(n86086), .Z(n86088) );
  NOR U105977 ( .A(n86088), .B(n86087), .Z(n86089) );
  NOR U105978 ( .A(n86090), .B(n86089), .Z(n91868) );
  IV U105979 ( .A(n91868), .Z(n86091) );
  NOR U105980 ( .A(n86092), .B(n86091), .Z(n91858) );
  XOR U105981 ( .A(n91860), .B(n91858), .Z(n91864) );
  IV U105982 ( .A(n86093), .Z(n86094) );
  NOR U105983 ( .A(n86095), .B(n86094), .Z(n91861) );
  XOR U105984 ( .A(n91864), .B(n91861), .Z(n86628) );
  IV U105985 ( .A(n86096), .Z(n86097) );
  NOR U105986 ( .A(n86098), .B(n86097), .Z(n91862) );
  NOR U105987 ( .A(n86100), .B(n86099), .Z(n86626) );
  NOR U105988 ( .A(n91862), .B(n86626), .Z(n86101) );
  XOR U105989 ( .A(n86628), .B(n86101), .Z(n86640) );
  XOR U105990 ( .A(n86642), .B(n86640), .Z(n86630) );
  XOR U105991 ( .A(n86629), .B(n86630), .Z(n86633) );
  XOR U105992 ( .A(n86632), .B(n86633), .Z(n91877) );
  IV U105993 ( .A(n86102), .Z(n86103) );
  NOR U105994 ( .A(n86104), .B(n86103), .Z(n91875) );
  XOR U105995 ( .A(n91877), .B(n91875), .Z(n91885) );
  XOR U105996 ( .A(n91884), .B(n91885), .Z(n91882) );
  XOR U105997 ( .A(n91881), .B(n91882), .Z(n91880) );
  IV U105998 ( .A(n86105), .Z(n86109) );
  IV U105999 ( .A(n86106), .Z(n86118) );
  NOR U106000 ( .A(n86107), .B(n86118), .Z(n86108) );
  IV U106001 ( .A(n86108), .Z(n86111) );
  NOR U106002 ( .A(n86109), .B(n86111), .Z(n91878) );
  XOR U106003 ( .A(n91880), .B(n91878), .Z(n86597) );
  IV U106004 ( .A(n86597), .Z(n86599) );
  IV U106005 ( .A(n86110), .Z(n86112) );
  NOR U106006 ( .A(n86112), .B(n86111), .Z(n86598) );
  IV U106007 ( .A(n86598), .Z(n86596) );
  XOR U106008 ( .A(n86599), .B(n86596), .Z(n86123) );
  IV U106009 ( .A(n86113), .Z(n86114) );
  NOR U106010 ( .A(n86114), .B(n86118), .Z(n86601) );
  NOR U106011 ( .A(n86116), .B(n86115), .Z(n86117) );
  IV U106012 ( .A(n86117), .Z(n86121) );
  XOR U106013 ( .A(n86119), .B(n86118), .Z(n86120) );
  NOR U106014 ( .A(n86121), .B(n86120), .Z(n86600) );
  NOR U106015 ( .A(n86601), .B(n86600), .Z(n86122) );
  XOR U106016 ( .A(n86123), .B(n86122), .Z(n86126) );
  IV U106017 ( .A(n86126), .Z(n86124) );
  NOR U106018 ( .A(n86125), .B(n86124), .Z(n86620) );
  NOR U106019 ( .A(n86127), .B(n86126), .Z(n86617) );
  IV U106020 ( .A(n86128), .Z(n86130) );
  NOR U106021 ( .A(n86130), .B(n86129), .Z(n86616) );
  XOR U106022 ( .A(n86617), .B(n86616), .Z(n86131) );
  NOR U106023 ( .A(n86620), .B(n86131), .Z(n86613) );
  XOR U106024 ( .A(n86615), .B(n86613), .Z(n86612) );
  IV U106025 ( .A(n86132), .Z(n86136) );
  NOR U106026 ( .A(n86133), .B(n86142), .Z(n86134) );
  IV U106027 ( .A(n86134), .Z(n86135) );
  NOR U106028 ( .A(n86136), .B(n86135), .Z(n86610) );
  XOR U106029 ( .A(n86612), .B(n86610), .Z(n86608) );
  IV U106030 ( .A(n86137), .Z(n86139) );
  NOR U106031 ( .A(n86139), .B(n86138), .Z(n86140) );
  IV U106032 ( .A(n86145), .Z(n86149) );
  NOR U106033 ( .A(n86140), .B(n86149), .Z(n86147) );
  IV U106034 ( .A(n86141), .Z(n86143) );
  NOR U106035 ( .A(n86143), .B(n86142), .Z(n86144) );
  NOR U106036 ( .A(n86145), .B(n86144), .Z(n86146) );
  NOR U106037 ( .A(n86147), .B(n86146), .Z(n86607) );
  XOR U106038 ( .A(n86608), .B(n86607), .Z(n91916) );
  IV U106039 ( .A(n86148), .Z(n86153) );
  NOR U106040 ( .A(n86150), .B(n86149), .Z(n86151) );
  IV U106041 ( .A(n86151), .Z(n86152) );
  NOR U106042 ( .A(n86153), .B(n86152), .Z(n91914) );
  XOR U106043 ( .A(n91916), .B(n91914), .Z(n91918) );
  XOR U106044 ( .A(n91917), .B(n91918), .Z(n91907) );
  XOR U106045 ( .A(n91908), .B(n91907), .Z(n86154) );
  IV U106046 ( .A(n86154), .Z(n91911) );
  XOR U106047 ( .A(n91909), .B(n91911), .Z(n86590) );
  XOR U106048 ( .A(n86588), .B(n86590), .Z(n86592) );
  XOR U106049 ( .A(n86591), .B(n86592), .Z(n86569) );
  XOR U106050 ( .A(n86570), .B(n86569), .Z(n86554) );
  IV U106051 ( .A(n86155), .Z(n86156) );
  NOR U106052 ( .A(n86157), .B(n86156), .Z(n86561) );
  IV U106053 ( .A(n86161), .Z(n86159) );
  NOR U106054 ( .A(n86159), .B(n86158), .Z(n86166) );
  NOR U106055 ( .A(n86161), .B(n86160), .Z(n86164) );
  IV U106056 ( .A(n86162), .Z(n86163) );
  NOR U106057 ( .A(n86164), .B(n86163), .Z(n86165) );
  NOR U106058 ( .A(n86166), .B(n86165), .Z(n86556) );
  XOR U106059 ( .A(n86561), .B(n86556), .Z(n86167) );
  XOR U106060 ( .A(n86554), .B(n86167), .Z(n86566) );
  XOR U106061 ( .A(n86168), .B(n86566), .Z(n86182) );
  XOR U106062 ( .A(n86181), .B(n86182), .Z(n86177) );
  IV U106063 ( .A(n86169), .Z(n86171) );
  NOR U106064 ( .A(n86171), .B(n86170), .Z(n86178) );
  IV U106065 ( .A(n86172), .Z(n86174) );
  NOR U106066 ( .A(n86174), .B(n86173), .Z(n86180) );
  NOR U106067 ( .A(n86178), .B(n86180), .Z(n86175) );
  IV U106068 ( .A(n86175), .Z(n86176) );
  NOR U106069 ( .A(n86177), .B(n86176), .Z(n86188) );
  IV U106070 ( .A(n86178), .Z(n86179) );
  IV U106071 ( .A(n86182), .Z(n86572) );
  NOR U106072 ( .A(n86179), .B(n86572), .Z(n86186) );
  IV U106073 ( .A(n86180), .Z(n86184) );
  IV U106074 ( .A(n86181), .Z(n86571) );
  XOR U106075 ( .A(n86182), .B(n86571), .Z(n86183) );
  NOR U106076 ( .A(n86184), .B(n86183), .Z(n86185) );
  NOR U106077 ( .A(n86186), .B(n86185), .Z(n86187) );
  IV U106078 ( .A(n86187), .Z(n86584) );
  NOR U106079 ( .A(n86188), .B(n86584), .Z(n86578) );
  IV U106080 ( .A(n86578), .Z(n86575) );
  XOR U106081 ( .A(n86576), .B(n86575), .Z(n86197) );
  IV U106082 ( .A(n86189), .Z(n86191) );
  NOR U106083 ( .A(n86191), .B(n86190), .Z(n86196) );
  IV U106084 ( .A(n86192), .Z(n86194) );
  IV U106085 ( .A(n86193), .Z(n86199) );
  NOR U106086 ( .A(n86194), .B(n86199), .Z(n86195) );
  NOR U106087 ( .A(n86196), .B(n86195), .Z(n86579) );
  XOR U106088 ( .A(n86197), .B(n86579), .Z(n86509) );
  IV U106089 ( .A(n86198), .Z(n86200) );
  NOR U106090 ( .A(n86200), .B(n86199), .Z(n86507) );
  XOR U106091 ( .A(n86509), .B(n86507), .Z(n86512) );
  XOR U106092 ( .A(n86510), .B(n86512), .Z(n86506) );
  XOR U106093 ( .A(n86505), .B(n86506), .Z(n86502) );
  XOR U106094 ( .A(n86501), .B(n86502), .Z(n86504) );
  XOR U106095 ( .A(n86503), .B(n86504), .Z(n86515) );
  XOR U106096 ( .A(n86514), .B(n86515), .Z(n86205) );
  IV U106097 ( .A(n86201), .Z(n86203) );
  NOR U106098 ( .A(n86203), .B(n86202), .Z(n86211) );
  IV U106099 ( .A(n86211), .Z(n86204) );
  NOR U106100 ( .A(n86205), .B(n86204), .Z(n86517) );
  IV U106101 ( .A(n86206), .Z(n86207) );
  NOR U106102 ( .A(n86208), .B(n86207), .Z(n86513) );
  NOR U106103 ( .A(n86513), .B(n86514), .Z(n86209) );
  XOR U106104 ( .A(n86515), .B(n86209), .Z(n86210) );
  NOR U106105 ( .A(n86211), .B(n86210), .Z(n86212) );
  NOR U106106 ( .A(n86517), .B(n86212), .Z(n86213) );
  IV U106107 ( .A(n86213), .Z(n86529) );
  XOR U106108 ( .A(n86528), .B(n86529), .Z(n86532) );
  XOR U106109 ( .A(n86531), .B(n86532), .Z(n86526) );
  XOR U106110 ( .A(n86525), .B(n86526), .Z(n86542) );
  XOR U106111 ( .A(n86541), .B(n86542), .Z(n86545) );
  XOR U106112 ( .A(n86544), .B(n86545), .Z(n86518) );
  XOR U106113 ( .A(n86519), .B(n86518), .Z(n86214) );
  IV U106114 ( .A(n86214), .Z(n86494) );
  XOR U106115 ( .A(n86493), .B(n86494), .Z(n86521) );
  XOR U106116 ( .A(n86491), .B(n86521), .Z(n91945) );
  IV U106117 ( .A(n86215), .Z(n86217) );
  IV U106118 ( .A(n86216), .Z(n86224) );
  NOR U106119 ( .A(n86217), .B(n86224), .Z(n86218) );
  NOR U106120 ( .A(n86218), .B(n91944), .Z(n86219) );
  XOR U106121 ( .A(n91945), .B(n86219), .Z(n86229) );
  IV U106122 ( .A(n86220), .Z(n86221) );
  NOR U106123 ( .A(n86222), .B(n86221), .Z(n86227) );
  IV U106124 ( .A(n86223), .Z(n86225) );
  NOR U106125 ( .A(n86225), .B(n86224), .Z(n86226) );
  NOR U106126 ( .A(n86227), .B(n86226), .Z(n86228) );
  XOR U106127 ( .A(n86229), .B(n86228), .Z(n91953) );
  XOR U106128 ( .A(n91952), .B(n91953), .Z(n91943) );
  IV U106129 ( .A(n86230), .Z(n86231) );
  NOR U106130 ( .A(n86232), .B(n86231), .Z(n91941) );
  XOR U106131 ( .A(n91943), .B(n91941), .Z(n91937) );
  IV U106132 ( .A(n91937), .Z(n86233) );
  NOR U106133 ( .A(n91936), .B(n86233), .Z(n86238) );
  IV U106134 ( .A(n86234), .Z(n86235) );
  NOR U106135 ( .A(n86236), .B(n86235), .Z(n86240) );
  IV U106136 ( .A(n86240), .Z(n86237) );
  NOR U106137 ( .A(n86238), .B(n86237), .Z(n91939) );
  XOR U106138 ( .A(n91936), .B(n91937), .Z(n86244) );
  IV U106139 ( .A(n86244), .Z(n86239) );
  NOR U106140 ( .A(n86240), .B(n86239), .Z(n86241) );
  NOR U106141 ( .A(n91939), .B(n86241), .Z(n86242) );
  NOR U106142 ( .A(n86243), .B(n86242), .Z(n86249) );
  IV U106143 ( .A(n86243), .Z(n86245) );
  NOR U106144 ( .A(n86245), .B(n86244), .Z(n91962) );
  NOR U106145 ( .A(n86249), .B(n91962), .Z(n86246) );
  NOR U106146 ( .A(n86247), .B(n86246), .Z(n86250) );
  IV U106147 ( .A(n86247), .Z(n86248) );
  NOR U106148 ( .A(n86249), .B(n86248), .Z(n91961) );
  NOR U106149 ( .A(n86250), .B(n91961), .Z(n86251) );
  IV U106150 ( .A(n86251), .Z(n91979) );
  XOR U106151 ( .A(n91978), .B(n91979), .Z(n91971) );
  XOR U106152 ( .A(n91972), .B(n91971), .Z(n91982) );
  IV U106153 ( .A(n91982), .Z(n91974) );
  XOR U106154 ( .A(n91981), .B(n91974), .Z(n91967) );
  IV U106155 ( .A(n86252), .Z(n86254) );
  NOR U106156 ( .A(n86254), .B(n86253), .Z(n91983) );
  IV U106157 ( .A(n86255), .Z(n86256) );
  NOR U106158 ( .A(n86257), .B(n86256), .Z(n91966) );
  NOR U106159 ( .A(n91983), .B(n91966), .Z(n86258) );
  XOR U106160 ( .A(n91967), .B(n86258), .Z(n86439) );
  XOR U106161 ( .A(n86259), .B(n86439), .Z(n86437) );
  XOR U106162 ( .A(n86438), .B(n86437), .Z(n86444) );
  IV U106163 ( .A(n86260), .Z(n86261) );
  NOR U106164 ( .A(n86265), .B(n86261), .Z(n86445) );
  NOR U106165 ( .A(n86444), .B(n86445), .Z(n86269) );
  IV U106166 ( .A(n86262), .Z(n86263) );
  NOR U106167 ( .A(n86263), .B(n86276), .Z(n86268) );
  IV U106168 ( .A(n86264), .Z(n86266) );
  NOR U106169 ( .A(n86266), .B(n86265), .Z(n86267) );
  NOR U106170 ( .A(n86268), .B(n86267), .Z(n86270) );
  NOR U106171 ( .A(n86269), .B(n86270), .Z(n86448) );
  IV U106172 ( .A(n86270), .Z(n86272) );
  XOR U106173 ( .A(n86445), .B(n86444), .Z(n86271) );
  NOR U106174 ( .A(n86272), .B(n86271), .Z(n86273) );
  NOR U106175 ( .A(n86448), .B(n86273), .Z(n86452) );
  IV U106176 ( .A(n86274), .Z(n86275) );
  NOR U106177 ( .A(n86276), .B(n86275), .Z(n86277) );
  IV U106178 ( .A(n86277), .Z(n86454) );
  XOR U106179 ( .A(n86452), .B(n86454), .Z(n86456) );
  XOR U106180 ( .A(n86455), .B(n86456), .Z(n92001) );
  XOR U106181 ( .A(n91999), .B(n92001), .Z(n92003) );
  XOR U106182 ( .A(n92002), .B(n92003), .Z(n86482) );
  XOR U106183 ( .A(n86278), .B(n86482), .Z(n86279) );
  NOR U106184 ( .A(n86280), .B(n86279), .Z(n86284) );
  IV U106185 ( .A(n86280), .Z(n86282) );
  XOR U106186 ( .A(n86469), .B(n86482), .Z(n86281) );
  NOR U106187 ( .A(n86282), .B(n86281), .Z(n86283) );
  NOR U106188 ( .A(n86284), .B(n86283), .Z(n86285) );
  XOR U106189 ( .A(n86286), .B(n86285), .Z(n86462) );
  XOR U106190 ( .A(n86464), .B(n86462), .Z(n86465) );
  XOR U106191 ( .A(n86466), .B(n86465), .Z(n92026) );
  XOR U106192 ( .A(n92028), .B(n92026), .Z(n92031) );
  IV U106193 ( .A(n86287), .Z(n86289) );
  NOR U106194 ( .A(n86289), .B(n86288), .Z(n92029) );
  XOR U106195 ( .A(n92031), .B(n92029), .Z(n92017) );
  XOR U106196 ( .A(n92016), .B(n92017), .Z(n92020) );
  XOR U106197 ( .A(n92019), .B(n92020), .Z(n92010) );
  XOR U106198 ( .A(n92009), .B(n92010), .Z(n92013) );
  IV U106199 ( .A(n86290), .Z(n86292) );
  NOR U106200 ( .A(n86292), .B(n86291), .Z(n86293) );
  IV U106201 ( .A(n86293), .Z(n92012) );
  XOR U106202 ( .A(n92013), .B(n92012), .Z(n86294) );
  NOR U106203 ( .A(n86298), .B(n86294), .Z(n86300) );
  NOR U106204 ( .A(n86296), .B(n86295), .Z(n86302) );
  IV U106205 ( .A(n86302), .Z(n86297) );
  NOR U106206 ( .A(n86300), .B(n86297), .Z(n86412) );
  IV U106207 ( .A(n86298), .Z(n86299) );
  NOR U106208 ( .A(n92013), .B(n86299), .Z(n86413) );
  NOR U106209 ( .A(n86413), .B(n86300), .Z(n86301) );
  NOR U106210 ( .A(n86302), .B(n86301), .Z(n86303) );
  NOR U106211 ( .A(n86412), .B(n86303), .Z(n86427) );
  IV U106212 ( .A(n86427), .Z(n86429) );
  XOR U106213 ( .A(n86429), .B(n86428), .Z(n86416) );
  XOR U106214 ( .A(n86304), .B(n86416), .Z(n86417) );
  XOR U106215 ( .A(n86418), .B(n86417), .Z(n92062) );
  IV U106216 ( .A(n92062), .Z(n92060) );
  XOR U106217 ( .A(n86305), .B(n92060), .Z(n86306) );
  XOR U106218 ( .A(n92061), .B(n86306), .Z(n92046) );
  IV U106219 ( .A(n86307), .Z(n86309) );
  NOR U106220 ( .A(n86309), .B(n86308), .Z(n86310) );
  IV U106221 ( .A(n86310), .Z(n92045) );
  XOR U106222 ( .A(n92046), .B(n92045), .Z(n86311) );
  IV U106223 ( .A(n86311), .Z(n92047) );
  NOR U106224 ( .A(n92050), .B(n92047), .Z(n86319) );
  NOR U106225 ( .A(n86312), .B(n86311), .Z(n86317) );
  IV U106226 ( .A(n86313), .Z(n86316) );
  IV U106227 ( .A(n86314), .Z(n86315) );
  NOR U106228 ( .A(n86316), .B(n86315), .Z(n92049) );
  XOR U106229 ( .A(n86317), .B(n92049), .Z(n86318) );
  NOR U106230 ( .A(n86319), .B(n86318), .Z(n86323) );
  NOR U106231 ( .A(n86326), .B(n86323), .Z(n86320) );
  IV U106232 ( .A(n86320), .Z(n86321) );
  NOR U106233 ( .A(n86321), .B(n86322), .Z(n86332) );
  IV U106234 ( .A(n86322), .Z(n86327) );
  XOR U106235 ( .A(n86326), .B(n86327), .Z(n86325) );
  IV U106236 ( .A(n86323), .Z(n86324) );
  NOR U106237 ( .A(n86325), .B(n86324), .Z(n86330) );
  IV U106238 ( .A(n86326), .Z(n86328) );
  NOR U106239 ( .A(n86328), .B(n86327), .Z(n86329) );
  NOR U106240 ( .A(n86330), .B(n86329), .Z(n86331) );
  IV U106241 ( .A(n86331), .Z(n92043) );
  NOR U106242 ( .A(n86332), .B(n92043), .Z(n92040) );
  NOR U106243 ( .A(n86334), .B(n86333), .Z(n86335) );
  IV U106244 ( .A(n86335), .Z(n86336) );
  NOR U106245 ( .A(n86337), .B(n86336), .Z(n86338) );
  IV U106246 ( .A(n86338), .Z(n92041) );
  XOR U106247 ( .A(n92040), .B(n92041), .Z(n92078) );
  XOR U106248 ( .A(n92077), .B(n92078), .Z(n92081) );
  XOR U106249 ( .A(n92080), .B(n92081), .Z(n92088) );
  XOR U106250 ( .A(n92087), .B(n92088), .Z(n92091) );
  XOR U106251 ( .A(n92090), .B(n92091), .Z(n86339) );
  NOR U106252 ( .A(n86340), .B(n86339), .Z(n92076) );
  NOR U106253 ( .A(n86342), .B(n86341), .Z(n92073) );
  NOR U106254 ( .A(n92090), .B(n92073), .Z(n86343) );
  XOR U106255 ( .A(n92091), .B(n86343), .Z(n86344) );
  NOR U106256 ( .A(n86345), .B(n86344), .Z(n86346) );
  NOR U106257 ( .A(n92076), .B(n86346), .Z(n86347) );
  IV U106258 ( .A(n86347), .Z(n92309) );
  IV U106259 ( .A(n86348), .Z(n86350) );
  NOR U106260 ( .A(n86350), .B(n86349), .Z(n92308) );
  XOR U106261 ( .A(n92309), .B(n92308), .Z(n92311) );
  XOR U106262 ( .A(n86351), .B(n92311), .Z(n92306) );
  XOR U106263 ( .A(n92307), .B(n92306), .Z(n92252) );
  IV U106264 ( .A(n92252), .Z(n86377) );
  NOR U106265 ( .A(n86353), .B(n86352), .Z(n86354) );
  XOR U106266 ( .A(n86355), .B(n86354), .Z(n86381) );
  XOR U106267 ( .A(n86357), .B(n86356), .Z(n86382) );
  NOR U106268 ( .A(n86359), .B(n86358), .Z(n86360) );
  XOR U106269 ( .A(n86361), .B(n86360), .Z(n92106) );
  IV U106270 ( .A(n92106), .Z(n86402) );
  XOR U106271 ( .A(n86363), .B(n86362), .Z(n86384) );
  IV U106272 ( .A(n86364), .Z(n86366) );
  NOR U106273 ( .A(n86366), .B(n86365), .Z(n92118) );
  IV U106274 ( .A(n92118), .Z(n86367) );
  NOR U106275 ( .A(n86368), .B(n86367), .Z(n92116) );
  IV U106276 ( .A(n92116), .Z(n86369) );
  NOR U106277 ( .A(n86370), .B(n86369), .Z(n86385) );
  IV U106278 ( .A(n86385), .Z(n86371) );
  NOR U106279 ( .A(n86384), .B(n86371), .Z(n92105) );
  IV U106280 ( .A(n92105), .Z(n86372) );
  NOR U106281 ( .A(n86402), .B(n86372), .Z(n86383) );
  IV U106282 ( .A(n86383), .Z(n86373) );
  NOR U106283 ( .A(n86382), .B(n86373), .Z(n92132) );
  IV U106284 ( .A(n92132), .Z(n86374) );
  NOR U106285 ( .A(n86374), .B(n86404), .Z(n86378) );
  IV U106286 ( .A(n86378), .Z(n86375) );
  NOR U106287 ( .A(n86381), .B(n86375), .Z(n92250) );
  IV U106288 ( .A(n92250), .Z(n86376) );
  NOR U106289 ( .A(n86377), .B(n86376), .Z(n86411) );
  NOR U106290 ( .A(n92252), .B(n92250), .Z(n86409) );
  NOR U106291 ( .A(n86379), .B(n86378), .Z(n86380) );
  XOR U106292 ( .A(n86381), .B(n86380), .Z(n92241) );
  IV U106293 ( .A(n92241), .Z(n92173) );
  XOR U106294 ( .A(n86383), .B(n86382), .Z(n92102) );
  XOR U106295 ( .A(n86385), .B(n86384), .Z(n92108) );
  NOR U106296 ( .A(n86387), .B(n86386), .Z(n86389) );
  NOR U106297 ( .A(n86389), .B(n86388), .Z(n86390) );
  XOR U106298 ( .A(n92112), .B(n86390), .Z(n92117) );
  IV U106299 ( .A(n92117), .Z(n92136) );
  XOR U106300 ( .A(n86391), .B(n92121), .Z(n86396) );
  IV U106301 ( .A(n86392), .Z(n86394) );
  NOR U106302 ( .A(n86394), .B(n86393), .Z(n92142) );
  IV U106303 ( .A(n92142), .Z(n86395) );
  NOR U106304 ( .A(n86396), .B(n86395), .Z(n92115) );
  IV U106305 ( .A(n92115), .Z(n86397) );
  NOR U106306 ( .A(n92136), .B(n86397), .Z(n86398) );
  IV U106307 ( .A(n86398), .Z(n86399) );
  NOR U106308 ( .A(n92113), .B(n86399), .Z(n92109) );
  IV U106309 ( .A(n92109), .Z(n86400) );
  NOR U106310 ( .A(n92108), .B(n86400), .Z(n92104) );
  IV U106311 ( .A(n92104), .Z(n86401) );
  NOR U106312 ( .A(n86402), .B(n86401), .Z(n92103) );
  IV U106313 ( .A(n92103), .Z(n86403) );
  NOR U106314 ( .A(n92102), .B(n86403), .Z(n92131) );
  IV U106315 ( .A(n92131), .Z(n86406) );
  XOR U106316 ( .A(n86405), .B(n86404), .Z(n92134) );
  NOR U106317 ( .A(n86406), .B(n92134), .Z(n92242) );
  IV U106318 ( .A(n92242), .Z(n86407) );
  NOR U106319 ( .A(n92173), .B(n86407), .Z(n92246) );
  IV U106320 ( .A(n92246), .Z(n86408) );
  NOR U106321 ( .A(n86409), .B(n86408), .Z(n86410) );
  NOR U106322 ( .A(n86411), .B(n86410), .Z(n92100) );
  NOR U106323 ( .A(n86413), .B(n86412), .Z(n92072) );
  IV U106324 ( .A(n86414), .Z(n86415) );
  NOR U106325 ( .A(n86416), .B(n86415), .Z(n86426) );
  IV U106326 ( .A(n86417), .Z(n86419) );
  NOR U106327 ( .A(n86419), .B(n86418), .Z(n86423) );
  IV U106328 ( .A(n86420), .Z(n86421) );
  NOR U106329 ( .A(n86421), .B(n92062), .Z(n86422) );
  NOR U106330 ( .A(n86423), .B(n86422), .Z(n86424) );
  IV U106331 ( .A(n86424), .Z(n86425) );
  NOR U106332 ( .A(n86426), .B(n86425), .Z(n86436) );
  NOR U106333 ( .A(n86428), .B(n86427), .Z(n86434) );
  IV U106334 ( .A(n86428), .Z(n86430) );
  NOR U106335 ( .A(n86430), .B(n86429), .Z(n86431) );
  NOR U106336 ( .A(n86432), .B(n86431), .Z(n86433) );
  NOR U106337 ( .A(n86434), .B(n86433), .Z(n86435) );
  XOR U106338 ( .A(n86436), .B(n86435), .Z(n92039) );
  NOR U106339 ( .A(n86438), .B(n86437), .Z(n86443) );
  IV U106340 ( .A(n86439), .Z(n91964) );
  IV U106341 ( .A(n86440), .Z(n86441) );
  NOR U106342 ( .A(n91964), .B(n86441), .Z(n86442) );
  NOR U106343 ( .A(n86443), .B(n86442), .Z(n86451) );
  IV U106344 ( .A(n86444), .Z(n86447) );
  IV U106345 ( .A(n86445), .Z(n86446) );
  NOR U106346 ( .A(n86447), .B(n86446), .Z(n86449) );
  NOR U106347 ( .A(n86449), .B(n86448), .Z(n86450) );
  XOR U106348 ( .A(n86451), .B(n86450), .Z(n86461) );
  IV U106349 ( .A(n86452), .Z(n86453) );
  NOR U106350 ( .A(n86454), .B(n86453), .Z(n86459) );
  IV U106351 ( .A(n86455), .Z(n86457) );
  NOR U106352 ( .A(n86457), .B(n86456), .Z(n86458) );
  NOR U106353 ( .A(n86459), .B(n86458), .Z(n86460) );
  XOR U106354 ( .A(n86461), .B(n86460), .Z(n86488) );
  IV U106355 ( .A(n86462), .Z(n86463) );
  NOR U106356 ( .A(n86464), .B(n86463), .Z(n86468) );
  NOR U106357 ( .A(n86466), .B(n86465), .Z(n86467) );
  NOR U106358 ( .A(n86468), .B(n86467), .Z(n86486) );
  IV U106359 ( .A(n86469), .Z(n86470) );
  NOR U106360 ( .A(n86482), .B(n86470), .Z(n86478) );
  XOR U106361 ( .A(n86482), .B(n86470), .Z(n86471) );
  NOR U106362 ( .A(n86480), .B(n86471), .Z(n86476) );
  NOR U106363 ( .A(n86473), .B(n86472), .Z(n86474) );
  IV U106364 ( .A(n86474), .Z(n86475) );
  NOR U106365 ( .A(n86476), .B(n86475), .Z(n86477) );
  NOR U106366 ( .A(n86478), .B(n86477), .Z(n86479) );
  IV U106367 ( .A(n86479), .Z(n86484) );
  IV U106368 ( .A(n86480), .Z(n86481) );
  NOR U106369 ( .A(n86482), .B(n86481), .Z(n86483) );
  NOR U106370 ( .A(n86484), .B(n86483), .Z(n86485) );
  XOR U106371 ( .A(n86486), .B(n86485), .Z(n86487) );
  XOR U106372 ( .A(n86488), .B(n86487), .Z(n91998) );
  IV U106373 ( .A(n86489), .Z(n86490) );
  NOR U106374 ( .A(n86490), .B(n91945), .Z(n86500) );
  IV U106375 ( .A(n86491), .Z(n86492) );
  NOR U106376 ( .A(n86492), .B(n86521), .Z(n86497) );
  IV U106377 ( .A(n86493), .Z(n86495) );
  NOR U106378 ( .A(n86495), .B(n86494), .Z(n86496) );
  NOR U106379 ( .A(n86497), .B(n86496), .Z(n86498) );
  IV U106380 ( .A(n86498), .Z(n86499) );
  NOR U106381 ( .A(n86500), .B(n86499), .Z(n91935) );
  IV U106382 ( .A(n86507), .Z(n86508) );
  IV U106383 ( .A(n86510), .Z(n86511) );
  IV U106384 ( .A(n86514), .Z(n86516) );
  NOR U106385 ( .A(n86519), .B(n86518), .Z(n86524) );
  IV U106386 ( .A(n86520), .Z(n86522) );
  NOR U106387 ( .A(n86522), .B(n86521), .Z(n86523) );
  NOR U106388 ( .A(n86524), .B(n86523), .Z(n86540) );
  IV U106389 ( .A(n86525), .Z(n86527) );
  NOR U106390 ( .A(n86527), .B(n86526), .Z(n86538) );
  IV U106391 ( .A(n86528), .Z(n86530) );
  NOR U106392 ( .A(n86530), .B(n86529), .Z(n86535) );
  IV U106393 ( .A(n86531), .Z(n86533) );
  NOR U106394 ( .A(n86533), .B(n86532), .Z(n86534) );
  NOR U106395 ( .A(n86535), .B(n86534), .Z(n86536) );
  IV U106396 ( .A(n86536), .Z(n86537) );
  NOR U106397 ( .A(n86538), .B(n86537), .Z(n86539) );
  XOR U106398 ( .A(n86540), .B(n86539), .Z(n86550) );
  IV U106399 ( .A(n86541), .Z(n86543) );
  NOR U106400 ( .A(n86543), .B(n86542), .Z(n86548) );
  IV U106401 ( .A(n86544), .Z(n86546) );
  NOR U106402 ( .A(n86546), .B(n86545), .Z(n86547) );
  NOR U106403 ( .A(n86548), .B(n86547), .Z(n86549) );
  XOR U106404 ( .A(n86550), .B(n86549), .Z(n86551) );
  XOR U106405 ( .A(n86552), .B(n86551), .Z(n91933) );
  IV U106406 ( .A(n86556), .Z(n86553) );
  NOR U106407 ( .A(n86554), .B(n86553), .Z(n86563) );
  IV U106408 ( .A(n86554), .Z(n86555) );
  NOR U106409 ( .A(n86556), .B(n86555), .Z(n86557) );
  NOR U106410 ( .A(n86558), .B(n86557), .Z(n86559) );
  IV U106411 ( .A(n86559), .Z(n86560) );
  NOR U106412 ( .A(n86561), .B(n86560), .Z(n86562) );
  NOR U106413 ( .A(n86563), .B(n86562), .Z(n86568) );
  IV U106414 ( .A(n86564), .Z(n86565) );
  NOR U106415 ( .A(n86566), .B(n86565), .Z(n86567) );
  NOR U106416 ( .A(n86568), .B(n86567), .Z(n91931) );
  NOR U106417 ( .A(n86570), .B(n86569), .Z(n86574) );
  NOR U106418 ( .A(n86572), .B(n86571), .Z(n86573) );
  NOR U106419 ( .A(n86574), .B(n86573), .Z(n86587) );
  NOR U106420 ( .A(n86576), .B(n86575), .Z(n86582) );
  IV U106421 ( .A(n86576), .Z(n86577) );
  NOR U106422 ( .A(n86578), .B(n86577), .Z(n86580) );
  NOR U106423 ( .A(n86580), .B(n86579), .Z(n86581) );
  NOR U106424 ( .A(n86582), .B(n86581), .Z(n86583) );
  IV U106425 ( .A(n86583), .Z(n86585) );
  NOR U106426 ( .A(n86585), .B(n86584), .Z(n86586) );
  XOR U106427 ( .A(n86587), .B(n86586), .Z(n91929) );
  IV U106428 ( .A(n86588), .Z(n86589) );
  NOR U106429 ( .A(n86590), .B(n86589), .Z(n86595) );
  IV U106430 ( .A(n86591), .Z(n86593) );
  NOR U106431 ( .A(n86593), .B(n86592), .Z(n86594) );
  NOR U106432 ( .A(n86595), .B(n86594), .Z(n91927) );
  NOR U106433 ( .A(n86597), .B(n86596), .Z(n86606) );
  NOR U106434 ( .A(n86599), .B(n86598), .Z(n86604) );
  XOR U106435 ( .A(n86601), .B(n86600), .Z(n86602) );
  IV U106436 ( .A(n86602), .Z(n86603) );
  NOR U106437 ( .A(n86604), .B(n86603), .Z(n86605) );
  NOR U106438 ( .A(n86606), .B(n86605), .Z(n91906) );
  IV U106439 ( .A(n86607), .Z(n86609) );
  NOR U106440 ( .A(n86609), .B(n86608), .Z(n91898) );
  IV U106441 ( .A(n86610), .Z(n86611) );
  NOR U106442 ( .A(n86612), .B(n86611), .Z(n86625) );
  IV U106443 ( .A(n86613), .Z(n86614) );
  NOR U106444 ( .A(n86615), .B(n86614), .Z(n86623) );
  IV U106445 ( .A(n86616), .Z(n86618) );
  NOR U106446 ( .A(n86618), .B(n86617), .Z(n86619) );
  NOR U106447 ( .A(n86620), .B(n86619), .Z(n86621) );
  IV U106448 ( .A(n86621), .Z(n86622) );
  NOR U106449 ( .A(n86623), .B(n86622), .Z(n86624) );
  IV U106450 ( .A(n86624), .Z(n91900) );
  NOR U106451 ( .A(n86625), .B(n91900), .Z(n91896) );
  IV U106452 ( .A(n86626), .Z(n86627) );
  NOR U106453 ( .A(n86628), .B(n86627), .Z(n86639) );
  IV U106454 ( .A(n86629), .Z(n86631) );
  NOR U106455 ( .A(n86631), .B(n86630), .Z(n86636) );
  IV U106456 ( .A(n86632), .Z(n86634) );
  NOR U106457 ( .A(n86634), .B(n86633), .Z(n86635) );
  NOR U106458 ( .A(n86636), .B(n86635), .Z(n86637) );
  IV U106459 ( .A(n86637), .Z(n86638) );
  NOR U106460 ( .A(n86639), .B(n86638), .Z(n91874) );
  IV U106461 ( .A(n86640), .Z(n86641) );
  NOR U106462 ( .A(n86642), .B(n86641), .Z(n91872) );
  IV U106463 ( .A(n86643), .Z(n86644) );
  NOR U106464 ( .A(n91840), .B(n86644), .Z(n86649) );
  IV U106465 ( .A(n86645), .Z(n86646) );
  NOR U106466 ( .A(n86647), .B(n86646), .Z(n86648) );
  NOR U106467 ( .A(n86649), .B(n86648), .Z(n91857) );
  IV U106468 ( .A(n86660), .Z(n86662) );
  NOR U106469 ( .A(n86662), .B(n86661), .Z(n86667) );
  IV U106470 ( .A(n86663), .Z(n86665) );
  NOR U106471 ( .A(n86665), .B(n86664), .Z(n86666) );
  NOR U106472 ( .A(n86667), .B(n86666), .Z(n91807) );
  IV U106473 ( .A(n86668), .Z(n86670) );
  NOR U106474 ( .A(n86670), .B(n86669), .Z(n86675) );
  IV U106475 ( .A(n86671), .Z(n86673) );
  NOR U106476 ( .A(n86673), .B(n86672), .Z(n86674) );
  NOR U106477 ( .A(n86675), .B(n86674), .Z(n86686) );
  IV U106478 ( .A(n86679), .Z(n86676) );
  NOR U106479 ( .A(n86677), .B(n86676), .Z(n86684) );
  IV U106480 ( .A(n86678), .Z(n86682) );
  NOR U106481 ( .A(n86680), .B(n86679), .Z(n86681) );
  NOR U106482 ( .A(n86682), .B(n86681), .Z(n86683) );
  NOR U106483 ( .A(n86684), .B(n86683), .Z(n86685) );
  XOR U106484 ( .A(n86686), .B(n86685), .Z(n86702) );
  IV U106485 ( .A(n86687), .Z(n86690) );
  IV U106486 ( .A(n86688), .Z(n86689) );
  NOR U106487 ( .A(n86690), .B(n86689), .Z(n86700) );
  XOR U106488 ( .A(n86693), .B(n86694), .Z(n86692) );
  NOR U106489 ( .A(n86692), .B(n86691), .Z(n86697) );
  IV U106490 ( .A(n86693), .Z(n86695) );
  NOR U106491 ( .A(n86695), .B(n86694), .Z(n86696) );
  NOR U106492 ( .A(n86697), .B(n86696), .Z(n86698) );
  IV U106493 ( .A(n86698), .Z(n86699) );
  NOR U106494 ( .A(n86700), .B(n86699), .Z(n86701) );
  XOR U106495 ( .A(n86702), .B(n86701), .Z(n86721) );
  NOR U106496 ( .A(n86704), .B(n86703), .Z(n86710) );
  NOR U106497 ( .A(n86706), .B(n86705), .Z(n86707) );
  NOR U106498 ( .A(n86708), .B(n86707), .Z(n86709) );
  NOR U106499 ( .A(n86710), .B(n86709), .Z(n86719) );
  NOR U106500 ( .A(n86712), .B(n86711), .Z(n86717) );
  IV U106501 ( .A(n86713), .Z(n86715) );
  NOR U106502 ( .A(n86715), .B(n86714), .Z(n86716) );
  NOR U106503 ( .A(n86717), .B(n86716), .Z(n86718) );
  XOR U106504 ( .A(n86719), .B(n86718), .Z(n86720) );
  XOR U106505 ( .A(n86721), .B(n86720), .Z(n91764) );
  IV U106506 ( .A(n86722), .Z(n86724) );
  NOR U106507 ( .A(n86724), .B(n86723), .Z(n86728) );
  NOR U106508 ( .A(n86726), .B(n86725), .Z(n86727) );
  NOR U106509 ( .A(n86728), .B(n86727), .Z(n86737) );
  IV U106510 ( .A(n86729), .Z(n86731) );
  NOR U106511 ( .A(n86731), .B(n86730), .Z(n86735) );
  NOR U106512 ( .A(n86733), .B(n86732), .Z(n86734) );
  NOR U106513 ( .A(n86735), .B(n86734), .Z(n86736) );
  XOR U106514 ( .A(n86737), .B(n86736), .Z(n86747) );
  IV U106515 ( .A(n86738), .Z(n86740) );
  NOR U106516 ( .A(n86740), .B(n86739), .Z(n86745) );
  IV U106517 ( .A(n86741), .Z(n86743) );
  NOR U106518 ( .A(n86743), .B(n86742), .Z(n86744) );
  NOR U106519 ( .A(n86745), .B(n86744), .Z(n86746) );
  XOR U106520 ( .A(n86747), .B(n86746), .Z(n91733) );
  NOR U106521 ( .A(n86749), .B(n86748), .Z(n86750) );
  NOR U106522 ( .A(n86751), .B(n86750), .Z(n86764) );
  IV U106523 ( .A(n86752), .Z(n86754) );
  NOR U106524 ( .A(n86754), .B(n86753), .Z(n86756) );
  NOR U106525 ( .A(n86756), .B(n86755), .Z(n86757) );
  IV U106526 ( .A(n86757), .Z(n86762) );
  IV U106527 ( .A(n86758), .Z(n86759) );
  NOR U106528 ( .A(n86760), .B(n86759), .Z(n86761) );
  NOR U106529 ( .A(n86762), .B(n86761), .Z(n86763) );
  XOR U106530 ( .A(n86764), .B(n86763), .Z(n91731) );
  IV U106531 ( .A(n86765), .Z(n86767) );
  NOR U106532 ( .A(n86767), .B(n86766), .Z(n86772) );
  IV U106533 ( .A(n86768), .Z(n86770) );
  NOR U106534 ( .A(n86770), .B(n86769), .Z(n86771) );
  NOR U106535 ( .A(n86772), .B(n86771), .Z(n86781) );
  NOR U106536 ( .A(n86774), .B(n86773), .Z(n86779) );
  IV U106537 ( .A(n86775), .Z(n86776) );
  NOR U106538 ( .A(n86777), .B(n86776), .Z(n86778) );
  NOR U106539 ( .A(n86779), .B(n86778), .Z(n86780) );
  XOR U106540 ( .A(n86781), .B(n86780), .Z(n86791) );
  NOR U106541 ( .A(n86783), .B(n86782), .Z(n86789) );
  IV U106542 ( .A(n86783), .Z(n86785) );
  NOR U106543 ( .A(n86785), .B(n86784), .Z(n86786) );
  NOR U106544 ( .A(n86787), .B(n86786), .Z(n86788) );
  NOR U106545 ( .A(n86789), .B(n86788), .Z(n86790) );
  XOR U106546 ( .A(n86791), .B(n86790), .Z(n86821) );
  NOR U106547 ( .A(n86793), .B(n86792), .Z(n86798) );
  IV U106548 ( .A(n86794), .Z(n86796) );
  NOR U106549 ( .A(n86796), .B(n86795), .Z(n86797) );
  NOR U106550 ( .A(n86798), .B(n86797), .Z(n86813) );
  IV U106551 ( .A(n86799), .Z(n86800) );
  NOR U106552 ( .A(n86801), .B(n86800), .Z(n86811) );
  IV U106553 ( .A(n86802), .Z(n86804) );
  NOR U106554 ( .A(n86804), .B(n86803), .Z(n86808) );
  NOR U106555 ( .A(n86806), .B(n86805), .Z(n86807) );
  NOR U106556 ( .A(n86808), .B(n86807), .Z(n86809) );
  IV U106557 ( .A(n86809), .Z(n86810) );
  NOR U106558 ( .A(n86811), .B(n86810), .Z(n86812) );
  XOR U106559 ( .A(n86813), .B(n86812), .Z(n86819) );
  NOR U106560 ( .A(n86815), .B(n86814), .Z(n86816) );
  NOR U106561 ( .A(n86817), .B(n86816), .Z(n86818) );
  XOR U106562 ( .A(n86819), .B(n86818), .Z(n86820) );
  XOR U106563 ( .A(n86821), .B(n86820), .Z(n91729) );
  IV U106564 ( .A(n86822), .Z(n86824) );
  NOR U106565 ( .A(n86824), .B(n86823), .Z(n86829) );
  IV U106566 ( .A(n86825), .Z(n86827) );
  NOR U106567 ( .A(n86827), .B(n86826), .Z(n86828) );
  NOR U106568 ( .A(n86829), .B(n86828), .Z(n91727) );
  IV U106569 ( .A(n86830), .Z(n86832) );
  NOR U106570 ( .A(n86832), .B(n86831), .Z(n86837) );
  IV U106571 ( .A(n86833), .Z(n86839) );
  IV U106572 ( .A(n86834), .Z(n86835) );
  NOR U106573 ( .A(n86839), .B(n86835), .Z(n86836) );
  XOR U106574 ( .A(n86837), .B(n86836), .Z(n86846) );
  NOR U106575 ( .A(n86839), .B(n86838), .Z(n86844) );
  IV U106576 ( .A(n86840), .Z(n86841) );
  NOR U106577 ( .A(n86842), .B(n86841), .Z(n86843) );
  NOR U106578 ( .A(n86844), .B(n86843), .Z(n86845) );
  XOR U106579 ( .A(n86846), .B(n86845), .Z(n86871) );
  IV U106580 ( .A(n86847), .Z(n86849) );
  NOR U106581 ( .A(n86849), .B(n86848), .Z(n86853) );
  NOR U106582 ( .A(n86851), .B(n86850), .Z(n86852) );
  NOR U106583 ( .A(n86853), .B(n86852), .Z(n86863) );
  IV U106584 ( .A(n86854), .Z(n86856) );
  NOR U106585 ( .A(n86856), .B(n86855), .Z(n86861) );
  IV U106586 ( .A(n86857), .Z(n86859) );
  NOR U106587 ( .A(n86859), .B(n86858), .Z(n86860) );
  NOR U106588 ( .A(n86861), .B(n86860), .Z(n86862) );
  XOR U106589 ( .A(n86863), .B(n86862), .Z(n86869) );
  NOR U106590 ( .A(n86865), .B(n86864), .Z(n86867) );
  NOR U106591 ( .A(n86867), .B(n86866), .Z(n86868) );
  XOR U106592 ( .A(n86869), .B(n86868), .Z(n86870) );
  XOR U106593 ( .A(n86871), .B(n86870), .Z(n91725) );
  IV U106594 ( .A(n86872), .Z(n86875) );
  IV U106595 ( .A(n86873), .Z(n86874) );
  NOR U106596 ( .A(n86875), .B(n86874), .Z(n86885) );
  IV U106597 ( .A(n86876), .Z(n86877) );
  NOR U106598 ( .A(n86878), .B(n86877), .Z(n86882) );
  NOR U106599 ( .A(n86880), .B(n86879), .Z(n86881) );
  NOR U106600 ( .A(n86882), .B(n86881), .Z(n86883) );
  IV U106601 ( .A(n86883), .Z(n86884) );
  NOR U106602 ( .A(n86885), .B(n86884), .Z(n91723) );
  NOR U106603 ( .A(n86893), .B(n86892), .Z(n86899) );
  IV U106604 ( .A(n86893), .Z(n86895) );
  NOR U106605 ( .A(n86895), .B(n86894), .Z(n86896) );
  NOR U106606 ( .A(n86897), .B(n86896), .Z(n86898) );
  NOR U106607 ( .A(n86899), .B(n86898), .Z(n86900) );
  XOR U106608 ( .A(n86901), .B(n86900), .Z(n91721) );
  IV U106609 ( .A(n86902), .Z(n86904) );
  NOR U106610 ( .A(n86904), .B(n86903), .Z(n86909) );
  IV U106611 ( .A(n86905), .Z(n86906) );
  NOR U106612 ( .A(n86907), .B(n86906), .Z(n86908) );
  NOR U106613 ( .A(n86909), .B(n86908), .Z(n86919) );
  IV U106614 ( .A(n86910), .Z(n86911) );
  NOR U106615 ( .A(n86912), .B(n86911), .Z(n86917) );
  IV U106616 ( .A(n86913), .Z(n86915) );
  NOR U106617 ( .A(n86915), .B(n86914), .Z(n86916) );
  NOR U106618 ( .A(n86917), .B(n86916), .Z(n86918) );
  XOR U106619 ( .A(n86919), .B(n86918), .Z(n91719) );
  NOR U106620 ( .A(n86921), .B(n86920), .Z(n86922) );
  NOR U106621 ( .A(n86922), .B(n86923), .Z(n86927) );
  IV U106622 ( .A(n86923), .Z(n86924) );
  NOR U106623 ( .A(n86925), .B(n86924), .Z(n86926) );
  NOR U106624 ( .A(n86927), .B(n86926), .Z(n86928) );
  IV U106625 ( .A(n86928), .Z(n86929) );
  NOR U106626 ( .A(n86930), .B(n86929), .Z(n86931) );
  NOR U106627 ( .A(n86932), .B(n86931), .Z(n91701) );
  NOR U106628 ( .A(n86934), .B(n86933), .Z(n86935) );
  XOR U106629 ( .A(n86935), .B(n86942), .Z(n86944) );
  IV U106630 ( .A(n86936), .Z(n86939) );
  IV U106631 ( .A(n86937), .Z(n86938) );
  NOR U106632 ( .A(n86939), .B(n86938), .Z(n86940) );
  IV U106633 ( .A(n86940), .Z(n86941) );
  NOR U106634 ( .A(n86942), .B(n86941), .Z(n86943) );
  NOR U106635 ( .A(n86944), .B(n86943), .Z(n91699) );
  IV U106636 ( .A(n86945), .Z(n86946) );
  NOR U106637 ( .A(n86946), .B(n86956), .Z(n86967) );
  IV U106638 ( .A(n86947), .Z(n86948) );
  NOR U106639 ( .A(n86949), .B(n86948), .Z(n86954) );
  IV U106640 ( .A(n86950), .Z(n86951) );
  NOR U106641 ( .A(n86952), .B(n86951), .Z(n86953) );
  NOR U106642 ( .A(n86954), .B(n86953), .Z(n86965) );
  IV U106643 ( .A(n86955), .Z(n86957) );
  NOR U106644 ( .A(n86957), .B(n86956), .Z(n86963) );
  IV U106645 ( .A(n86958), .Z(n86961) );
  IV U106646 ( .A(n86959), .Z(n86960) );
  NOR U106647 ( .A(n86961), .B(n86960), .Z(n86962) );
  NOR U106648 ( .A(n86963), .B(n86962), .Z(n86964) );
  XOR U106649 ( .A(n86965), .B(n86964), .Z(n86966) );
  XOR U106650 ( .A(n86967), .B(n86966), .Z(n86978) );
  IV U106651 ( .A(n86968), .Z(n86969) );
  NOR U106652 ( .A(n86970), .B(n86969), .Z(n86974) );
  NOR U106653 ( .A(n86972), .B(n86971), .Z(n86973) );
  NOR U106654 ( .A(n86974), .B(n86973), .Z(n86975) );
  XOR U106655 ( .A(n86976), .B(n86975), .Z(n86977) );
  XOR U106656 ( .A(n86978), .B(n86977), .Z(n91682) );
  NOR U106657 ( .A(n86979), .B(n86980), .Z(n86988) );
  IV U106658 ( .A(n86980), .Z(n86981) );
  NOR U106659 ( .A(n86982), .B(n86981), .Z(n86986) );
  XOR U106660 ( .A(n86984), .B(n86983), .Z(n86985) );
  NOR U106661 ( .A(n86986), .B(n86985), .Z(n86987) );
  NOR U106662 ( .A(n86988), .B(n86987), .Z(n86998) );
  IV U106663 ( .A(n86989), .Z(n86990) );
  NOR U106664 ( .A(n86991), .B(n86990), .Z(n86996) );
  IV U106665 ( .A(n86992), .Z(n86994) );
  NOR U106666 ( .A(n86994), .B(n86993), .Z(n86995) );
  NOR U106667 ( .A(n86996), .B(n86995), .Z(n86997) );
  XOR U106668 ( .A(n86998), .B(n86997), .Z(n91654) );
  IV U106669 ( .A(n86999), .Z(n87000) );
  NOR U106670 ( .A(n87001), .B(n87000), .Z(n87005) );
  NOR U106671 ( .A(n87003), .B(n87002), .Z(n87004) );
  NOR U106672 ( .A(n87005), .B(n87004), .Z(n91652) );
  IV U106673 ( .A(n87006), .Z(n87009) );
  IV U106674 ( .A(n87007), .Z(n87008) );
  NOR U106675 ( .A(n87009), .B(n87008), .Z(n91628) );
  NOR U106676 ( .A(n87011), .B(n87010), .Z(n87022) );
  NOR U106677 ( .A(n87013), .B(n87012), .Z(n87020) );
  NOR U106678 ( .A(n87015), .B(n87014), .Z(n87017) );
  XOR U106679 ( .A(n87017), .B(n87016), .Z(n87018) );
  IV U106680 ( .A(n87018), .Z(n87019) );
  NOR U106681 ( .A(n87020), .B(n87019), .Z(n87021) );
  NOR U106682 ( .A(n87022), .B(n87021), .Z(n87032) );
  IV U106683 ( .A(n87023), .Z(n87024) );
  NOR U106684 ( .A(n87025), .B(n87024), .Z(n87030) );
  IV U106685 ( .A(n87026), .Z(n87027) );
  NOR U106686 ( .A(n87028), .B(n87027), .Z(n87029) );
  NOR U106687 ( .A(n87030), .B(n87029), .Z(n87031) );
  XOR U106688 ( .A(n87032), .B(n87031), .Z(n87046) );
  IV U106689 ( .A(n87033), .Z(n87034) );
  NOR U106690 ( .A(n87035), .B(n87034), .Z(n87044) );
  NOR U106691 ( .A(n87037), .B(n87036), .Z(n87042) );
  IV U106692 ( .A(n87038), .Z(n87040) );
  NOR U106693 ( .A(n87040), .B(n87039), .Z(n87041) );
  NOR U106694 ( .A(n87042), .B(n87041), .Z(n87043) );
  XOR U106695 ( .A(n87044), .B(n87043), .Z(n87045) );
  XOR U106696 ( .A(n87046), .B(n87045), .Z(n91607) );
  IV U106697 ( .A(n87047), .Z(n87048) );
  NOR U106698 ( .A(n87056), .B(n87048), .Z(n87053) );
  IV U106699 ( .A(n87049), .Z(n87050) );
  NOR U106700 ( .A(n87051), .B(n87050), .Z(n87052) );
  NOR U106701 ( .A(n87053), .B(n87052), .Z(n87066) );
  IV U106702 ( .A(n87054), .Z(n87055) );
  NOR U106703 ( .A(n87056), .B(n87055), .Z(n87061) );
  IV U106704 ( .A(n87057), .Z(n87058) );
  NOR U106705 ( .A(n87059), .B(n87058), .Z(n87060) );
  NOR U106706 ( .A(n87061), .B(n87060), .Z(n87062) );
  IV U106707 ( .A(n87062), .Z(n87063) );
  NOR U106708 ( .A(n87064), .B(n87063), .Z(n87065) );
  XOR U106709 ( .A(n87066), .B(n87065), .Z(n87076) );
  IV U106710 ( .A(n87067), .Z(n87069) );
  NOR U106711 ( .A(n87069), .B(n87068), .Z(n87074) );
  IV U106712 ( .A(n87070), .Z(n87072) );
  NOR U106713 ( .A(n87072), .B(n87071), .Z(n87073) );
  NOR U106714 ( .A(n87074), .B(n87073), .Z(n87075) );
  XOR U106715 ( .A(n87076), .B(n87075), .Z(n91562) );
  IV U106716 ( .A(n87077), .Z(n87079) );
  NOR U106717 ( .A(n87079), .B(n87078), .Z(n91560) );
  XOR U106718 ( .A(n87104), .B(n87080), .Z(n87081) );
  NOR U106719 ( .A(n87082), .B(n87081), .Z(n87087) );
  NOR U106720 ( .A(n87105), .B(n87083), .Z(n87084) );
  NOR U106721 ( .A(n87085), .B(n87084), .Z(n87086) );
  NOR U106722 ( .A(n87087), .B(n87086), .Z(n91558) );
  NOR U106723 ( .A(n87089), .B(n87088), .Z(n87091) );
  NOR U106724 ( .A(n87091), .B(n87090), .Z(n87100) );
  NOR U106725 ( .A(n87093), .B(n87092), .Z(n87098) );
  IV U106726 ( .A(n87094), .Z(n87096) );
  NOR U106727 ( .A(n87096), .B(n87095), .Z(n87097) );
  NOR U106728 ( .A(n87098), .B(n87097), .Z(n87099) );
  XOR U106729 ( .A(n87100), .B(n87099), .Z(n91556) );
  IV U106730 ( .A(n87101), .Z(n87102) );
  NOR U106731 ( .A(n87103), .B(n87102), .Z(n87108) );
  IV U106732 ( .A(n87104), .Z(n87106) );
  NOR U106733 ( .A(n87106), .B(n87105), .Z(n87107) );
  NOR U106734 ( .A(n87108), .B(n87107), .Z(n91554) );
  IV U106735 ( .A(n87109), .Z(n87114) );
  IV U106736 ( .A(n87110), .Z(n87111) );
  NOR U106737 ( .A(n87114), .B(n87111), .Z(n87121) );
  IV U106738 ( .A(n87112), .Z(n87113) );
  NOR U106739 ( .A(n87114), .B(n87113), .Z(n87119) );
  IV U106740 ( .A(n87115), .Z(n87116) );
  NOR U106741 ( .A(n87117), .B(n87116), .Z(n87118) );
  NOR U106742 ( .A(n87119), .B(n87118), .Z(n87120) );
  XOR U106743 ( .A(n87121), .B(n87120), .Z(n87130) );
  NOR U106744 ( .A(n87123), .B(n87122), .Z(n87128) );
  IV U106745 ( .A(n87124), .Z(n87126) );
  NOR U106746 ( .A(n87126), .B(n87125), .Z(n87127) );
  NOR U106747 ( .A(n87128), .B(n87127), .Z(n87129) );
  XOR U106748 ( .A(n87130), .B(n87129), .Z(n87149) );
  IV U106749 ( .A(n87131), .Z(n87133) );
  NOR U106750 ( .A(n87133), .B(n87132), .Z(n87137) );
  NOR U106751 ( .A(n87135), .B(n87134), .Z(n87136) );
  NOR U106752 ( .A(n87137), .B(n87136), .Z(n87147) );
  IV U106753 ( .A(n87138), .Z(n87140) );
  NOR U106754 ( .A(n87140), .B(n87139), .Z(n87145) );
  IV U106755 ( .A(n87141), .Z(n87142) );
  NOR U106756 ( .A(n87143), .B(n87142), .Z(n87144) );
  NOR U106757 ( .A(n87145), .B(n87144), .Z(n87146) );
  XOR U106758 ( .A(n87147), .B(n87146), .Z(n87148) );
  XOR U106759 ( .A(n87149), .B(n87148), .Z(n91552) );
  NOR U106760 ( .A(n87151), .B(n87150), .Z(n87159) );
  NOR U106761 ( .A(n87153), .B(n87152), .Z(n87157) );
  XOR U106762 ( .A(n87155), .B(n87154), .Z(n87156) );
  NOR U106763 ( .A(n87157), .B(n87156), .Z(n87158) );
  NOR U106764 ( .A(n87159), .B(n87158), .Z(n87187) );
  IV U106765 ( .A(n87160), .Z(n87162) );
  NOR U106766 ( .A(n87162), .B(n87161), .Z(n87166) );
  NOR U106767 ( .A(n87164), .B(n87163), .Z(n87165) );
  NOR U106768 ( .A(n87166), .B(n87165), .Z(n87175) );
  NOR U106769 ( .A(n87168), .B(n87167), .Z(n87173) );
  IV U106770 ( .A(n87169), .Z(n87171) );
  NOR U106771 ( .A(n87171), .B(n87170), .Z(n87172) );
  NOR U106772 ( .A(n87173), .B(n87172), .Z(n87174) );
  XOR U106773 ( .A(n87175), .B(n87174), .Z(n87185) );
  IV U106774 ( .A(n87176), .Z(n87177) );
  NOR U106775 ( .A(n87178), .B(n87177), .Z(n87183) );
  IV U106776 ( .A(n87179), .Z(n87180) );
  NOR U106777 ( .A(n87181), .B(n87180), .Z(n87182) );
  NOR U106778 ( .A(n87183), .B(n87182), .Z(n87184) );
  XOR U106779 ( .A(n87185), .B(n87184), .Z(n87186) );
  XOR U106780 ( .A(n87187), .B(n87186), .Z(n91488) );
  IV U106781 ( .A(n87188), .Z(n91491) );
  IV U106782 ( .A(n87189), .Z(n87190) );
  NOR U106783 ( .A(n91491), .B(n87190), .Z(n87195) );
  IV U106784 ( .A(n87191), .Z(n87192) );
  NOR U106785 ( .A(n87193), .B(n87192), .Z(n87194) );
  NOR U106786 ( .A(n87195), .B(n87194), .Z(n91486) );
  IV U106787 ( .A(n87196), .Z(n87197) );
  NOR U106788 ( .A(n87198), .B(n87197), .Z(n91484) );
  IV U106789 ( .A(n87199), .Z(n87201) );
  NOR U106790 ( .A(n87201), .B(n87200), .Z(n87206) );
  IV U106791 ( .A(n87202), .Z(n87204) );
  NOR U106792 ( .A(n87204), .B(n87203), .Z(n87205) );
  NOR U106793 ( .A(n87206), .B(n87205), .Z(n87216) );
  IV U106794 ( .A(n87207), .Z(n87209) );
  NOR U106795 ( .A(n87209), .B(n87208), .Z(n87214) );
  IV U106796 ( .A(n87210), .Z(n87211) );
  NOR U106797 ( .A(n87212), .B(n87211), .Z(n87213) );
  NOR U106798 ( .A(n87214), .B(n87213), .Z(n87215) );
  XOR U106799 ( .A(n87216), .B(n87215), .Z(n91452) );
  IV U106800 ( .A(n87217), .Z(n87220) );
  IV U106801 ( .A(n87218), .Z(n87219) );
  NOR U106802 ( .A(n87220), .B(n87219), .Z(n91450) );
  IV U106803 ( .A(n87221), .Z(n87222) );
  NOR U106804 ( .A(n87223), .B(n87222), .Z(n87227) );
  IV U106805 ( .A(n87224), .Z(n87225) );
  NOR U106806 ( .A(n87226), .B(n87225), .Z(n87232) );
  XOR U106807 ( .A(n87227), .B(n87232), .Z(n87234) );
  NOR U106808 ( .A(n87229), .B(n87228), .Z(n87230) );
  IV U106809 ( .A(n87230), .Z(n87231) );
  NOR U106810 ( .A(n87232), .B(n87231), .Z(n87233) );
  NOR U106811 ( .A(n87234), .B(n87233), .Z(n91448) );
  IV U106812 ( .A(n87235), .Z(n87236) );
  NOR U106813 ( .A(n87237), .B(n87236), .Z(n87241) );
  NOR U106814 ( .A(n87239), .B(n87238), .Z(n87240) );
  NOR U106815 ( .A(n87241), .B(n87240), .Z(n91446) );
  IV U106816 ( .A(n87242), .Z(n87246) );
  XOR U106817 ( .A(n87243), .B(n87246), .Z(n87245) );
  NOR U106818 ( .A(n87245), .B(n87244), .Z(n87249) );
  NOR U106819 ( .A(n87247), .B(n87246), .Z(n87248) );
  NOR U106820 ( .A(n87249), .B(n87248), .Z(n91444) );
  NOR U106821 ( .A(n87251), .B(n87250), .Z(n87257) );
  NOR U106822 ( .A(n87253), .B(n87252), .Z(n87254) );
  NOR U106823 ( .A(n87255), .B(n87254), .Z(n87256) );
  XOR U106824 ( .A(n87257), .B(n87256), .Z(n87267) );
  IV U106825 ( .A(n87258), .Z(n87259) );
  NOR U106826 ( .A(n87260), .B(n87259), .Z(n87265) );
  IV U106827 ( .A(n87261), .Z(n87263) );
  NOR U106828 ( .A(n87263), .B(n87262), .Z(n87264) );
  NOR U106829 ( .A(n87265), .B(n87264), .Z(n87266) );
  XOR U106830 ( .A(n87267), .B(n87266), .Z(n87287) );
  IV U106831 ( .A(n87278), .Z(n87281) );
  IV U106832 ( .A(n87279), .Z(n87280) );
  NOR U106833 ( .A(n87281), .B(n87280), .Z(n87282) );
  NOR U106834 ( .A(n87283), .B(n87282), .Z(n87284) );
  XOR U106835 ( .A(n87285), .B(n87284), .Z(n87286) );
  XOR U106836 ( .A(n87287), .B(n87286), .Z(n91442) );
  IV U106837 ( .A(n87288), .Z(n87290) );
  NOR U106838 ( .A(n87290), .B(n87289), .Z(n87310) );
  IV U106839 ( .A(n87291), .Z(n87293) );
  NOR U106840 ( .A(n87293), .B(n87292), .Z(n87298) );
  IV U106841 ( .A(n87294), .Z(n87296) );
  NOR U106842 ( .A(n87296), .B(n87295), .Z(n87297) );
  NOR U106843 ( .A(n87298), .B(n87297), .Z(n87308) );
  IV U106844 ( .A(n87299), .Z(n87301) );
  NOR U106845 ( .A(n87301), .B(n87300), .Z(n87306) );
  IV U106846 ( .A(n87302), .Z(n87304) );
  NOR U106847 ( .A(n87304), .B(n87303), .Z(n87305) );
  NOR U106848 ( .A(n87306), .B(n87305), .Z(n87307) );
  XOR U106849 ( .A(n87308), .B(n87307), .Z(n87309) );
  XOR U106850 ( .A(n87310), .B(n87309), .Z(n87330) );
  IV U106851 ( .A(n87311), .Z(n87312) );
  NOR U106852 ( .A(n87313), .B(n87312), .Z(n87318) );
  IV U106853 ( .A(n87314), .Z(n87316) );
  NOR U106854 ( .A(n87316), .B(n87315), .Z(n87317) );
  NOR U106855 ( .A(n87318), .B(n87317), .Z(n87328) );
  IV U106856 ( .A(n87319), .Z(n87320) );
  NOR U106857 ( .A(n87321), .B(n87320), .Z(n87326) );
  IV U106858 ( .A(n87322), .Z(n87323) );
  NOR U106859 ( .A(n87324), .B(n87323), .Z(n87325) );
  NOR U106860 ( .A(n87326), .B(n87325), .Z(n87327) );
  XOR U106861 ( .A(n87328), .B(n87327), .Z(n87329) );
  XOR U106862 ( .A(n87330), .B(n87329), .Z(n91386) );
  IV U106863 ( .A(n87331), .Z(n87333) );
  NOR U106864 ( .A(n87333), .B(n87332), .Z(n87337) );
  NOR U106865 ( .A(n87335), .B(n87334), .Z(n87336) );
  NOR U106866 ( .A(n87337), .B(n87336), .Z(n87347) );
  IV U106867 ( .A(n87338), .Z(n87340) );
  NOR U106868 ( .A(n87340), .B(n87339), .Z(n87345) );
  IV U106869 ( .A(n87341), .Z(n87343) );
  NOR U106870 ( .A(n87343), .B(n87342), .Z(n87344) );
  NOR U106871 ( .A(n87345), .B(n87344), .Z(n87346) );
  XOR U106872 ( .A(n87347), .B(n87346), .Z(n87357) );
  IV U106873 ( .A(n87348), .Z(n87350) );
  NOR U106874 ( .A(n87350), .B(n87349), .Z(n87355) );
  IV U106875 ( .A(n87351), .Z(n87353) );
  NOR U106876 ( .A(n87353), .B(n87352), .Z(n87354) );
  NOR U106877 ( .A(n87355), .B(n87354), .Z(n87356) );
  XOR U106878 ( .A(n87357), .B(n87356), .Z(n87377) );
  XOR U106879 ( .A(n87360), .B(n87361), .Z(n87359) );
  NOR U106880 ( .A(n87359), .B(n87358), .Z(n87364) );
  IV U106881 ( .A(n87360), .Z(n87362) );
  NOR U106882 ( .A(n87362), .B(n87361), .Z(n87363) );
  NOR U106883 ( .A(n87364), .B(n87363), .Z(n87375) );
  IV U106884 ( .A(n87368), .Z(n87365) );
  NOR U106885 ( .A(n87366), .B(n87365), .Z(n87373) );
  IV U106886 ( .A(n87367), .Z(n87371) );
  NOR U106887 ( .A(n87369), .B(n87368), .Z(n87370) );
  NOR U106888 ( .A(n87371), .B(n87370), .Z(n87372) );
  NOR U106889 ( .A(n87373), .B(n87372), .Z(n87374) );
  XOR U106890 ( .A(n87375), .B(n87374), .Z(n87376) );
  XOR U106891 ( .A(n87377), .B(n87376), .Z(n91313) );
  NOR U106892 ( .A(n87379), .B(n87378), .Z(n87383) );
  IV U106893 ( .A(n87380), .Z(n87382) );
  NOR U106894 ( .A(n87382), .B(n87381), .Z(n87389) );
  XOR U106895 ( .A(n87383), .B(n87389), .Z(n87391) );
  IV U106896 ( .A(n87384), .Z(n87385) );
  NOR U106897 ( .A(n87386), .B(n87385), .Z(n87387) );
  IV U106898 ( .A(n87387), .Z(n87388) );
  NOR U106899 ( .A(n87389), .B(n87388), .Z(n87390) );
  NOR U106900 ( .A(n87391), .B(n87390), .Z(n91311) );
  IV U106901 ( .A(n87392), .Z(n87393) );
  NOR U106902 ( .A(n87405), .B(n87393), .Z(n87403) );
  IV U106903 ( .A(n87394), .Z(n87396) );
  NOR U106904 ( .A(n87396), .B(n87395), .Z(n87401) );
  IV U106905 ( .A(n87397), .Z(n87398) );
  NOR U106906 ( .A(n87399), .B(n87398), .Z(n87400) );
  NOR U106907 ( .A(n87401), .B(n87400), .Z(n87402) );
  XOR U106908 ( .A(n87403), .B(n87402), .Z(n87413) );
  IV U106909 ( .A(n87404), .Z(n87406) );
  NOR U106910 ( .A(n87406), .B(n87405), .Z(n87411) );
  IV U106911 ( .A(n87407), .Z(n87409) );
  IV U106912 ( .A(n87408), .Z(n87418) );
  NOR U106913 ( .A(n87409), .B(n87418), .Z(n87410) );
  NOR U106914 ( .A(n87411), .B(n87410), .Z(n87412) );
  XOR U106915 ( .A(n87413), .B(n87412), .Z(n87448) );
  IV U106916 ( .A(n87414), .Z(n87415) );
  NOR U106917 ( .A(n87415), .B(n87426), .Z(n87420) );
  IV U106918 ( .A(n87416), .Z(n87417) );
  NOR U106919 ( .A(n87418), .B(n87417), .Z(n87419) );
  NOR U106920 ( .A(n87420), .B(n87419), .Z(n87431) );
  IV U106921 ( .A(n87421), .Z(n87424) );
  IV U106922 ( .A(n87422), .Z(n87423) );
  NOR U106923 ( .A(n87424), .B(n87423), .Z(n87429) );
  IV U106924 ( .A(n87425), .Z(n87427) );
  NOR U106925 ( .A(n87427), .B(n87426), .Z(n87428) );
  NOR U106926 ( .A(n87429), .B(n87428), .Z(n87430) );
  XOR U106927 ( .A(n87431), .B(n87430), .Z(n87446) );
  IV U106928 ( .A(n87432), .Z(n91292) );
  IV U106929 ( .A(n87433), .Z(n87434) );
  NOR U106930 ( .A(n91292), .B(n87434), .Z(n87444) );
  XOR U106931 ( .A(n87437), .B(n87438), .Z(n87436) );
  NOR U106932 ( .A(n87436), .B(n87435), .Z(n87441) );
  IV U106933 ( .A(n87437), .Z(n87439) );
  NOR U106934 ( .A(n87439), .B(n87438), .Z(n87440) );
  NOR U106935 ( .A(n87441), .B(n87440), .Z(n87442) );
  IV U106936 ( .A(n87442), .Z(n87443) );
  NOR U106937 ( .A(n87444), .B(n87443), .Z(n87445) );
  XOR U106938 ( .A(n87446), .B(n87445), .Z(n87447) );
  XOR U106939 ( .A(n87448), .B(n87447), .Z(n91284) );
  NOR U106940 ( .A(n87449), .B(n87450), .Z(n87456) );
  IV U106941 ( .A(n87450), .Z(n87451) );
  NOR U106942 ( .A(n87452), .B(n87451), .Z(n87453) );
  NOR U106943 ( .A(n87454), .B(n87453), .Z(n87455) );
  NOR U106944 ( .A(n87456), .B(n87455), .Z(n91282) );
  IV U106945 ( .A(n87457), .Z(n87460) );
  IV U106946 ( .A(n87458), .Z(n87459) );
  NOR U106947 ( .A(n87460), .B(n87459), .Z(n87475) );
  NOR U106948 ( .A(n87462), .B(n87461), .Z(n87467) );
  IV U106949 ( .A(n87463), .Z(n87465) );
  NOR U106950 ( .A(n87465), .B(n87464), .Z(n87466) );
  NOR U106951 ( .A(n87467), .B(n87466), .Z(n87473) );
  NOR U106952 ( .A(n87469), .B(n87468), .Z(n87470) );
  NOR U106953 ( .A(n87471), .B(n87470), .Z(n87472) );
  XOR U106954 ( .A(n87473), .B(n87472), .Z(n87474) );
  XOR U106955 ( .A(n87475), .B(n87474), .Z(n91267) );
  NOR U106956 ( .A(n87477), .B(n87476), .Z(n87486) );
  NOR U106957 ( .A(n87479), .B(n87478), .Z(n87482) );
  IV U106958 ( .A(n87480), .Z(n87481) );
  NOR U106959 ( .A(n87482), .B(n87481), .Z(n87483) );
  XOR U106960 ( .A(n87484), .B(n87483), .Z(n87485) );
  NOR U106961 ( .A(n87486), .B(n87485), .Z(n91265) );
  IV U106962 ( .A(n87487), .Z(n87489) );
  NOR U106963 ( .A(n87489), .B(n87488), .Z(n87490) );
  NOR U106964 ( .A(n87491), .B(n87490), .Z(n87507) );
  IV U106965 ( .A(n87492), .Z(n87493) );
  NOR U106966 ( .A(n87493), .B(n87498), .Z(n87497) );
  NOR U106967 ( .A(n87494), .B(n87498), .Z(n87495) );
  NOR U106968 ( .A(n87496), .B(n87495), .Z(n87503) );
  XOR U106969 ( .A(n87497), .B(n87503), .Z(n87505) );
  IV U106970 ( .A(n87498), .Z(n87500) );
  NOR U106971 ( .A(n87500), .B(n87499), .Z(n87501) );
  IV U106972 ( .A(n87501), .Z(n87502) );
  NOR U106973 ( .A(n87503), .B(n87502), .Z(n87504) );
  NOR U106974 ( .A(n87505), .B(n87504), .Z(n87506) );
  XOR U106975 ( .A(n87507), .B(n87506), .Z(n91216) );
  IV U106976 ( .A(n87508), .Z(n87510) );
  NOR U106977 ( .A(n87510), .B(n87509), .Z(n87512) );
  NOR U106978 ( .A(n87512), .B(n87511), .Z(n91214) );
  IV U106979 ( .A(n87513), .Z(n87514) );
  NOR U106980 ( .A(n87515), .B(n87514), .Z(n87520) );
  IV U106981 ( .A(n87516), .Z(n87518) );
  NOR U106982 ( .A(n87518), .B(n87517), .Z(n87519) );
  NOR U106983 ( .A(n87520), .B(n87519), .Z(n91142) );
  NOR U106984 ( .A(n87522), .B(n87521), .Z(n87527) );
  IV U106985 ( .A(n87523), .Z(n87524) );
  NOR U106986 ( .A(n87525), .B(n87524), .Z(n87526) );
  NOR U106987 ( .A(n87527), .B(n87526), .Z(n91130) );
  XOR U106988 ( .A(n87530), .B(n87528), .Z(n87529) );
  NOR U106989 ( .A(n87531), .B(n87529), .Z(n87537) );
  IV U106990 ( .A(n87530), .Z(n87533) );
  IV U106991 ( .A(n87531), .Z(n87532) );
  NOR U106992 ( .A(n87533), .B(n87532), .Z(n87534) );
  NOR U106993 ( .A(n87535), .B(n87534), .Z(n87536) );
  NOR U106994 ( .A(n87537), .B(n87536), .Z(n91089) );
  NOR U106995 ( .A(n87539), .B(n87538), .Z(n87540) );
  IV U106996 ( .A(n87540), .Z(n91009) );
  IV U106997 ( .A(n87541), .Z(n87542) );
  NOR U106998 ( .A(n91009), .B(n87542), .Z(n91027) );
  IV U106999 ( .A(n87543), .Z(n87545) );
  NOR U107000 ( .A(n87545), .B(n87544), .Z(n87549) );
  NOR U107001 ( .A(n87547), .B(n87546), .Z(n87548) );
  NOR U107002 ( .A(n87549), .B(n87548), .Z(n87559) );
  IV U107003 ( .A(n87550), .Z(n87552) );
  NOR U107004 ( .A(n87552), .B(n87551), .Z(n87557) );
  IV U107005 ( .A(n87553), .Z(n87555) );
  NOR U107006 ( .A(n87555), .B(n87554), .Z(n87556) );
  NOR U107007 ( .A(n87557), .B(n87556), .Z(n87558) );
  XOR U107008 ( .A(n87559), .B(n87558), .Z(n90999) );
  IV U107009 ( .A(n87560), .Z(n87561) );
  NOR U107010 ( .A(n87562), .B(n87561), .Z(n87566) );
  NOR U107011 ( .A(n87564), .B(n87563), .Z(n87565) );
  NOR U107012 ( .A(n87566), .B(n87565), .Z(n90997) );
  NOR U107013 ( .A(n87568), .B(n87567), .Z(n87574) );
  NOR U107014 ( .A(n87570), .B(n87569), .Z(n87571) );
  NOR U107015 ( .A(n87572), .B(n87571), .Z(n87573) );
  NOR U107016 ( .A(n87574), .B(n87573), .Z(n87584) );
  IV U107017 ( .A(n87575), .Z(n87576) );
  NOR U107018 ( .A(n87577), .B(n87576), .Z(n87582) );
  IV U107019 ( .A(n87578), .Z(n87579) );
  NOR U107020 ( .A(n87580), .B(n87579), .Z(n87581) );
  NOR U107021 ( .A(n87582), .B(n87581), .Z(n87583) );
  XOR U107022 ( .A(n87584), .B(n87583), .Z(n87594) );
  IV U107023 ( .A(n87585), .Z(n87587) );
  NOR U107024 ( .A(n87587), .B(n87586), .Z(n87592) );
  IV U107025 ( .A(n87588), .Z(n87590) );
  NOR U107026 ( .A(n87590), .B(n87589), .Z(n87591) );
  NOR U107027 ( .A(n87592), .B(n87591), .Z(n87593) );
  XOR U107028 ( .A(n87594), .B(n87593), .Z(n87611) );
  NOR U107029 ( .A(n87596), .B(n87595), .Z(n87609) );
  NOR U107030 ( .A(n87598), .B(n87597), .Z(n87599) );
  NOR U107031 ( .A(n87600), .B(n87599), .Z(n87607) );
  NOR U107032 ( .A(n87602), .B(n87601), .Z(n87603) );
  IV U107033 ( .A(n87603), .Z(n87604) );
  NOR U107034 ( .A(n87605), .B(n87604), .Z(n87606) );
  NOR U107035 ( .A(n87607), .B(n87606), .Z(n87608) );
  XOR U107036 ( .A(n87609), .B(n87608), .Z(n87610) );
  XOR U107037 ( .A(n87611), .B(n87610), .Z(n90995) );
  IV U107038 ( .A(n87612), .Z(n87614) );
  NOR U107039 ( .A(n87614), .B(n87613), .Z(n87619) );
  IV U107040 ( .A(n87615), .Z(n87616) );
  NOR U107041 ( .A(n87617), .B(n87616), .Z(n87618) );
  NOR U107042 ( .A(n87619), .B(n87618), .Z(n90971) );
  IV U107043 ( .A(n87620), .Z(n87622) );
  NOR U107044 ( .A(n87622), .B(n87621), .Z(n87627) );
  IV U107045 ( .A(n87623), .Z(n87625) );
  NOR U107046 ( .A(n87625), .B(n87624), .Z(n87626) );
  NOR U107047 ( .A(n87627), .B(n87626), .Z(n90949) );
  NOR U107048 ( .A(n87629), .B(n87628), .Z(n87630) );
  XOR U107049 ( .A(n87630), .B(n87635), .Z(n87637) );
  IV U107050 ( .A(n87631), .Z(n87632) );
  NOR U107051 ( .A(n87632), .B(n90926), .Z(n87633) );
  IV U107052 ( .A(n87633), .Z(n87634) );
  NOR U107053 ( .A(n87635), .B(n87634), .Z(n87636) );
  NOR U107054 ( .A(n87637), .B(n87636), .Z(n90947) );
  IV U107055 ( .A(n87638), .Z(n87639) );
  NOR U107056 ( .A(n87640), .B(n87639), .Z(n90945) );
  NOR U107057 ( .A(n87641), .B(n87647), .Z(n87646) );
  NOR U107058 ( .A(n87643), .B(n87642), .Z(n87644) );
  IV U107059 ( .A(n87644), .Z(n87645) );
  NOR U107060 ( .A(n87646), .B(n87645), .Z(n87651) );
  IV U107061 ( .A(n87647), .Z(n87649) );
  NOR U107062 ( .A(n87649), .B(n87648), .Z(n87650) );
  NOR U107063 ( .A(n87651), .B(n87650), .Z(n90924) );
  IV U107064 ( .A(n87656), .Z(n87657) );
  IV U107065 ( .A(n87658), .Z(n87660) );
  IV U107066 ( .A(n87661), .Z(n87662) );
  NOR U107067 ( .A(n87663), .B(n87662), .Z(n87668) );
  IV U107068 ( .A(n87664), .Z(n87665) );
  NOR U107069 ( .A(n87666), .B(n87665), .Z(n87667) );
  NOR U107070 ( .A(n87668), .B(n87667), .Z(n87672) );
  NOR U107071 ( .A(n87670), .B(n87669), .Z(n87671) );
  IV U107072 ( .A(n87673), .Z(n87674) );
  NOR U107073 ( .A(n87675), .B(n87674), .Z(n87680) );
  IV U107074 ( .A(n87676), .Z(n87678) );
  NOR U107075 ( .A(n87678), .B(n87677), .Z(n87679) );
  NOR U107076 ( .A(n87680), .B(n87679), .Z(n87690) );
  IV U107077 ( .A(n87681), .Z(n87709) );
  IV U107078 ( .A(n87682), .Z(n87683) );
  NOR U107079 ( .A(n87709), .B(n87683), .Z(n87688) );
  IV U107080 ( .A(n87684), .Z(n87686) );
  NOR U107081 ( .A(n87686), .B(n87685), .Z(n87687) );
  NOR U107082 ( .A(n87688), .B(n87687), .Z(n87689) );
  XOR U107083 ( .A(n87690), .B(n87689), .Z(n90873) );
  IV U107084 ( .A(n87691), .Z(n87693) );
  NOR U107085 ( .A(n87693), .B(n87692), .Z(n87698) );
  IV U107086 ( .A(n87694), .Z(n87695) );
  NOR U107087 ( .A(n87696), .B(n87695), .Z(n87697) );
  NOR U107088 ( .A(n87698), .B(n87697), .Z(n90871) );
  IV U107089 ( .A(n87699), .Z(n87700) );
  NOR U107090 ( .A(n87701), .B(n87700), .Z(n87706) );
  IV U107091 ( .A(n87702), .Z(n87703) );
  NOR U107092 ( .A(n87704), .B(n87703), .Z(n87705) );
  NOR U107093 ( .A(n87706), .B(n87705), .Z(n90869) );
  IV U107094 ( .A(n87707), .Z(n87708) );
  NOR U107095 ( .A(n87709), .B(n87708), .Z(n87714) );
  IV U107096 ( .A(n87710), .Z(n87711) );
  NOR U107097 ( .A(n87712), .B(n87711), .Z(n87713) );
  NOR U107098 ( .A(n87714), .B(n87713), .Z(n90867) );
  IV U107099 ( .A(n87715), .Z(n87716) );
  NOR U107100 ( .A(n87718), .B(n87716), .Z(n90865) );
  IV U107101 ( .A(n87717), .Z(n87719) );
  NOR U107102 ( .A(n87719), .B(n87718), .Z(n87725) );
  IV U107103 ( .A(n87720), .Z(n87723) );
  IV U107104 ( .A(n87721), .Z(n87722) );
  NOR U107105 ( .A(n87723), .B(n87722), .Z(n87724) );
  NOR U107106 ( .A(n87725), .B(n87724), .Z(n87731) );
  NOR U107107 ( .A(n87727), .B(n87726), .Z(n87729) );
  XOR U107108 ( .A(n90824), .B(n90825), .Z(n87728) );
  NOR U107109 ( .A(n87729), .B(n87728), .Z(n87730) );
  XOR U107110 ( .A(n87731), .B(n87730), .Z(n90842) );
  IV U107111 ( .A(n87732), .Z(n87733) );
  NOR U107112 ( .A(n87734), .B(n87733), .Z(n87738) );
  NOR U107113 ( .A(n87736), .B(n87735), .Z(n87737) );
  NOR U107114 ( .A(n87738), .B(n87737), .Z(n90820) );
  IV U107115 ( .A(n87739), .Z(n87740) );
  NOR U107116 ( .A(n87740), .B(n90831), .Z(n87745) );
  IV U107117 ( .A(n87741), .Z(n87742) );
  NOR U107118 ( .A(n87743), .B(n87742), .Z(n87744) );
  NOR U107119 ( .A(n87745), .B(n87744), .Z(n90818) );
  IV U107120 ( .A(n87746), .Z(n87748) );
  NOR U107121 ( .A(n87748), .B(n87747), .Z(n87750) );
  NOR U107122 ( .A(n87750), .B(n87749), .Z(n90816) );
  IV U107123 ( .A(n87751), .Z(n87752) );
  NOR U107124 ( .A(n87753), .B(n87752), .Z(n87757) );
  NOR U107125 ( .A(n87755), .B(n87754), .Z(n87756) );
  NOR U107126 ( .A(n87757), .B(n87756), .Z(n87766) );
  IV U107127 ( .A(n87758), .Z(n87759) );
  NOR U107128 ( .A(n87760), .B(n87759), .Z(n87764) );
  NOR U107129 ( .A(n87762), .B(n87761), .Z(n87763) );
  NOR U107130 ( .A(n87764), .B(n87763), .Z(n87765) );
  XOR U107131 ( .A(n87766), .B(n87765), .Z(n87786) );
  IV U107132 ( .A(n87767), .Z(n87770) );
  NOR U107133 ( .A(n87768), .B(n87774), .Z(n87769) );
  NOR U107134 ( .A(n87770), .B(n87769), .Z(n87784) );
  IV U107135 ( .A(n87771), .Z(n87773) );
  NOR U107136 ( .A(n87773), .B(n87772), .Z(n87781) );
  IV U107137 ( .A(n87774), .Z(n87775) );
  NOR U107138 ( .A(n87776), .B(n87775), .Z(n87778) );
  NOR U107139 ( .A(n87778), .B(n87777), .Z(n87779) );
  IV U107140 ( .A(n87779), .Z(n87780) );
  NOR U107141 ( .A(n87781), .B(n87780), .Z(n87782) );
  IV U107142 ( .A(n87782), .Z(n87783) );
  NOR U107143 ( .A(n87784), .B(n87783), .Z(n87785) );
  XOR U107144 ( .A(n87786), .B(n87785), .Z(n87800) );
  NOR U107145 ( .A(n87788), .B(n87787), .Z(n87798) );
  IV U107146 ( .A(n87789), .Z(n87790) );
  NOR U107147 ( .A(n87791), .B(n87790), .Z(n87796) );
  IV U107148 ( .A(n87792), .Z(n87794) );
  NOR U107149 ( .A(n87794), .B(n87793), .Z(n87795) );
  NOR U107150 ( .A(n87796), .B(n87795), .Z(n87797) );
  XOR U107151 ( .A(n87798), .B(n87797), .Z(n87799) );
  XOR U107152 ( .A(n87800), .B(n87799), .Z(n90795) );
  IV U107153 ( .A(n87801), .Z(n87802) );
  NOR U107154 ( .A(n87803), .B(n87802), .Z(n87807) );
  IV U107155 ( .A(n87804), .Z(n87805) );
  NOR U107156 ( .A(n87818), .B(n87805), .Z(n87806) );
  NOR U107157 ( .A(n87807), .B(n87806), .Z(n90793) );
  IV U107158 ( .A(n87808), .Z(n87810) );
  NOR U107159 ( .A(n87810), .B(n87809), .Z(n87815) );
  IV U107160 ( .A(n87811), .Z(n87813) );
  NOR U107161 ( .A(n87813), .B(n87812), .Z(n87814) );
  NOR U107162 ( .A(n87815), .B(n87814), .Z(n87820) );
  IV U107163 ( .A(n87816), .Z(n87817) );
  NOR U107164 ( .A(n87818), .B(n87817), .Z(n87819) );
  XOR U107165 ( .A(n87820), .B(n87819), .Z(n90791) );
  IV U107166 ( .A(n87821), .Z(n87823) );
  NOR U107167 ( .A(n87823), .B(n87822), .Z(n87828) );
  IV U107168 ( .A(n87824), .Z(n87826) );
  NOR U107169 ( .A(n87826), .B(n87825), .Z(n87827) );
  NOR U107170 ( .A(n87828), .B(n87827), .Z(n87837) );
  IV U107171 ( .A(n87829), .Z(n87831) );
  NOR U107172 ( .A(n87831), .B(n87830), .Z(n87835) );
  NOR U107173 ( .A(n87833), .B(n87832), .Z(n87834) );
  NOR U107174 ( .A(n87835), .B(n87834), .Z(n87836) );
  XOR U107175 ( .A(n87837), .B(n87836), .Z(n90774) );
  IV U107176 ( .A(n87838), .Z(n87839) );
  NOR U107177 ( .A(n87840), .B(n87839), .Z(n87845) );
  IV U107178 ( .A(n87841), .Z(n87842) );
  NOR U107179 ( .A(n87843), .B(n87842), .Z(n87844) );
  NOR U107180 ( .A(n87845), .B(n87844), .Z(n90772) );
  IV U107181 ( .A(n87846), .Z(n87848) );
  NOR U107182 ( .A(n87848), .B(n87847), .Z(n87853) );
  IV U107183 ( .A(n87849), .Z(n87850) );
  NOR U107184 ( .A(n87851), .B(n87850), .Z(n87852) );
  NOR U107185 ( .A(n87853), .B(n87852), .Z(n90770) );
  IV U107186 ( .A(n87854), .Z(n87855) );
  NOR U107187 ( .A(n87856), .B(n87855), .Z(n87862) );
  IV U107188 ( .A(n87857), .Z(n87860) );
  IV U107189 ( .A(n87858), .Z(n87859) );
  NOR U107190 ( .A(n87860), .B(n87859), .Z(n87861) );
  NOR U107191 ( .A(n87862), .B(n87861), .Z(n87877) );
  IV U107192 ( .A(n87863), .Z(n87864) );
  NOR U107193 ( .A(n87869), .B(n87864), .Z(n87875) );
  IV U107194 ( .A(n87865), .Z(n87867) );
  NOR U107195 ( .A(n87867), .B(n87866), .Z(n87872) );
  IV U107196 ( .A(n87868), .Z(n87870) );
  NOR U107197 ( .A(n87870), .B(n87869), .Z(n87871) );
  NOR U107198 ( .A(n87872), .B(n87871), .Z(n87873) );
  IV U107199 ( .A(n87873), .Z(n87874) );
  NOR U107200 ( .A(n87875), .B(n87874), .Z(n87876) );
  XOR U107201 ( .A(n87877), .B(n87876), .Z(n90768) );
  IV U107202 ( .A(n87878), .Z(n87879) );
  NOR U107203 ( .A(n87880), .B(n87879), .Z(n87881) );
  NOR U107204 ( .A(n87882), .B(n87881), .Z(n90766) );
  NOR U107205 ( .A(n87884), .B(n87883), .Z(n87895) );
  IV U107206 ( .A(n87889), .Z(n87885) );
  NOR U107207 ( .A(n87885), .B(n87887), .Z(n87893) );
  IV U107208 ( .A(n87886), .Z(n87891) );
  IV U107209 ( .A(n87887), .Z(n87888) );
  NOR U107210 ( .A(n87889), .B(n87888), .Z(n87890) );
  NOR U107211 ( .A(n87891), .B(n87890), .Z(n87892) );
  NOR U107212 ( .A(n87893), .B(n87892), .Z(n87894) );
  XOR U107213 ( .A(n87895), .B(n87894), .Z(n87905) );
  IV U107214 ( .A(n87896), .Z(n87898) );
  NOR U107215 ( .A(n87898), .B(n87897), .Z(n87903) );
  IV U107216 ( .A(n87899), .Z(n87900) );
  NOR U107217 ( .A(n87901), .B(n87900), .Z(n87902) );
  NOR U107218 ( .A(n87903), .B(n87902), .Z(n87904) );
  XOR U107219 ( .A(n87905), .B(n87904), .Z(n87929) );
  IV U107220 ( .A(n87906), .Z(n87907) );
  NOR U107221 ( .A(n87908), .B(n87907), .Z(n87913) );
  IV U107222 ( .A(n87909), .Z(n87911) );
  NOR U107223 ( .A(n87911), .B(n87910), .Z(n87912) );
  NOR U107224 ( .A(n87913), .B(n87912), .Z(n87917) );
  NOR U107225 ( .A(n87915), .B(n87914), .Z(n87916) );
  XOR U107226 ( .A(n87917), .B(n87916), .Z(n87927) );
  IV U107227 ( .A(n87918), .Z(n87919) );
  NOR U107228 ( .A(n87920), .B(n87919), .Z(n87925) );
  IV U107229 ( .A(n87921), .Z(n87922) );
  NOR U107230 ( .A(n87923), .B(n87922), .Z(n87924) );
  NOR U107231 ( .A(n87925), .B(n87924), .Z(n87926) );
  XOR U107232 ( .A(n87927), .B(n87926), .Z(n87928) );
  XOR U107233 ( .A(n87929), .B(n87928), .Z(n90744) );
  IV U107234 ( .A(n87930), .Z(n87933) );
  IV U107235 ( .A(n87931), .Z(n87932) );
  NOR U107236 ( .A(n87933), .B(n87932), .Z(n87941) );
  NOR U107237 ( .A(n87935), .B(n87934), .Z(n87939) );
  NOR U107238 ( .A(n87937), .B(n87936), .Z(n87938) );
  NOR U107239 ( .A(n87939), .B(n87938), .Z(n87940) );
  IV U107240 ( .A(n87942), .Z(n87944) );
  NOR U107241 ( .A(n87944), .B(n87943), .Z(n87954) );
  XOR U107242 ( .A(n87947), .B(n87948), .Z(n87946) );
  NOR U107243 ( .A(n87946), .B(n87945), .Z(n87951) );
  IV U107244 ( .A(n87947), .Z(n87949) );
  NOR U107245 ( .A(n87949), .B(n87948), .Z(n87950) );
  NOR U107246 ( .A(n87951), .B(n87950), .Z(n87952) );
  IV U107247 ( .A(n87952), .Z(n87953) );
  NOR U107248 ( .A(n87956), .B(n87955), .Z(n87961) );
  IV U107249 ( .A(n87957), .Z(n87958) );
  NOR U107250 ( .A(n87959), .B(n87958), .Z(n87960) );
  NOR U107251 ( .A(n87961), .B(n87960), .Z(n87966) );
  IV U107252 ( .A(n87969), .Z(n87962) );
  IV U107253 ( .A(n87970), .Z(n87968) );
  NOR U107254 ( .A(n87962), .B(n87968), .Z(n87963) );
  NOR U107255 ( .A(n87964), .B(n87963), .Z(n87965) );
  NOR U107256 ( .A(n87968), .B(n87967), .Z(n87976) );
  XOR U107257 ( .A(n87970), .B(n87969), .Z(n87971) );
  NOR U107258 ( .A(n87972), .B(n87971), .Z(n87974) );
  NOR U107259 ( .A(n87974), .B(n87973), .Z(n87975) );
  IV U107260 ( .A(n87979), .Z(n87980) );
  NOR U107261 ( .A(n87981), .B(n87980), .Z(n87986) );
  IV U107262 ( .A(n87982), .Z(n87984) );
  NOR U107263 ( .A(n87984), .B(n87983), .Z(n87985) );
  NOR U107264 ( .A(n87986), .B(n87985), .Z(n87996) );
  IV U107265 ( .A(n87987), .Z(n87988) );
  NOR U107266 ( .A(n87989), .B(n87988), .Z(n87994) );
  IV U107267 ( .A(n87990), .Z(n87991) );
  NOR U107268 ( .A(n87992), .B(n87991), .Z(n87993) );
  NOR U107269 ( .A(n87994), .B(n87993), .Z(n87995) );
  XOR U107270 ( .A(n87996), .B(n87995), .Z(n88004) );
  NOR U107271 ( .A(n87998), .B(n87997), .Z(n88002) );
  NOR U107272 ( .A(n88000), .B(n87999), .Z(n88001) );
  NOR U107273 ( .A(n88002), .B(n88001), .Z(n88003) );
  XOR U107274 ( .A(n88004), .B(n88003), .Z(n88023) );
  IV U107275 ( .A(n88005), .Z(n88006) );
  NOR U107276 ( .A(n88007), .B(n88006), .Z(n88011) );
  NOR U107277 ( .A(n88009), .B(n88008), .Z(n88010) );
  NOR U107278 ( .A(n88011), .B(n88010), .Z(n88021) );
  IV U107279 ( .A(n88012), .Z(n88014) );
  NOR U107280 ( .A(n88014), .B(n88013), .Z(n88019) );
  IV U107281 ( .A(n88015), .Z(n88017) );
  NOR U107282 ( .A(n88017), .B(n88016), .Z(n88018) );
  NOR U107283 ( .A(n88019), .B(n88018), .Z(n88020) );
  XOR U107284 ( .A(n88021), .B(n88020), .Z(n88022) );
  XOR U107285 ( .A(n88023), .B(n88022), .Z(n90724) );
  IV U107286 ( .A(n88024), .Z(n88026) );
  NOR U107287 ( .A(n88026), .B(n88025), .Z(n88031) );
  IV U107288 ( .A(n88027), .Z(n88028) );
  NOR U107289 ( .A(n88029), .B(n88028), .Z(n88030) );
  NOR U107290 ( .A(n88031), .B(n88030), .Z(n90722) );
  IV U107291 ( .A(n88032), .Z(n88036) );
  XOR U107292 ( .A(n88033), .B(n88036), .Z(n88035) );
  NOR U107293 ( .A(n88035), .B(n88034), .Z(n88039) );
  NOR U107294 ( .A(n88037), .B(n88036), .Z(n88038) );
  NOR U107295 ( .A(n88039), .B(n88038), .Z(n88048) );
  NOR U107296 ( .A(n88041), .B(n88040), .Z(n88046) );
  IV U107297 ( .A(n88042), .Z(n88044) );
  NOR U107298 ( .A(n88044), .B(n88043), .Z(n88045) );
  NOR U107299 ( .A(n88046), .B(n88045), .Z(n88047) );
  XOR U107300 ( .A(n88048), .B(n88047), .Z(n88058) );
  NOR U107301 ( .A(n88049), .B(n88050), .Z(n88056) );
  IV U107302 ( .A(n88050), .Z(n88051) );
  NOR U107303 ( .A(n88052), .B(n88051), .Z(n88053) );
  NOR U107304 ( .A(n88054), .B(n88053), .Z(n88055) );
  NOR U107305 ( .A(n88056), .B(n88055), .Z(n88057) );
  XOR U107306 ( .A(n88058), .B(n88057), .Z(n88077) );
  IV U107307 ( .A(n88059), .Z(n88061) );
  NOR U107308 ( .A(n88061), .B(n88060), .Z(n88065) );
  NOR U107309 ( .A(n88063), .B(n88062), .Z(n88064) );
  NOR U107310 ( .A(n88065), .B(n88064), .Z(n88075) );
  NOR U107311 ( .A(n88067), .B(n88066), .Z(n88073) );
  IV U107312 ( .A(n88067), .Z(n88069) );
  NOR U107313 ( .A(n88069), .B(n88068), .Z(n88070) );
  NOR U107314 ( .A(n88071), .B(n88070), .Z(n88072) );
  NOR U107315 ( .A(n88073), .B(n88072), .Z(n88074) );
  XOR U107316 ( .A(n88075), .B(n88074), .Z(n88076) );
  XOR U107317 ( .A(n88077), .B(n88076), .Z(n90720) );
  IV U107318 ( .A(n88078), .Z(n88079) );
  NOR U107319 ( .A(n88080), .B(n88079), .Z(n88084) );
  NOR U107320 ( .A(n88082), .B(n88081), .Z(n88083) );
  NOR U107321 ( .A(n88084), .B(n88083), .Z(n90697) );
  IV U107322 ( .A(n88085), .Z(n88087) );
  NOR U107323 ( .A(n88087), .B(n88086), .Z(n88088) );
  XOR U107324 ( .A(n88088), .B(n88093), .Z(n88095) );
  IV U107325 ( .A(n88089), .Z(n88090) );
  NOR U107326 ( .A(n88097), .B(n88090), .Z(n88091) );
  IV U107327 ( .A(n88091), .Z(n88092) );
  NOR U107328 ( .A(n88093), .B(n88092), .Z(n88094) );
  NOR U107329 ( .A(n88095), .B(n88094), .Z(n90666) );
  IV U107330 ( .A(n88096), .Z(n88098) );
  NOR U107331 ( .A(n88098), .B(n88097), .Z(n88103) );
  IV U107332 ( .A(n88099), .Z(n88101) );
  NOR U107333 ( .A(n88101), .B(n88100), .Z(n88102) );
  XOR U107334 ( .A(n88103), .B(n88102), .Z(n90652) );
  IV U107335 ( .A(n88104), .Z(n88105) );
  NOR U107336 ( .A(n88106), .B(n88105), .Z(n88133) );
  IV U107337 ( .A(n88110), .Z(n88107) );
  NOR U107338 ( .A(n88108), .B(n88107), .Z(n88118) );
  NOR U107339 ( .A(n88110), .B(n88109), .Z(n88116) );
  IV U107340 ( .A(n88111), .Z(n88112) );
  NOR U107341 ( .A(n88113), .B(n88112), .Z(n88114) );
  IV U107342 ( .A(n88114), .Z(n88115) );
  NOR U107343 ( .A(n88116), .B(n88115), .Z(n88117) );
  NOR U107344 ( .A(n88118), .B(n88117), .Z(n88131) );
  NOR U107345 ( .A(n88119), .B(n88120), .Z(n88129) );
  IV U107346 ( .A(n88120), .Z(n88121) );
  NOR U107347 ( .A(n88122), .B(n88121), .Z(n88127) );
  NOR U107348 ( .A(n88124), .B(n88123), .Z(n88125) );
  IV U107349 ( .A(n88125), .Z(n88126) );
  NOR U107350 ( .A(n88127), .B(n88126), .Z(n88128) );
  NOR U107351 ( .A(n88129), .B(n88128), .Z(n88130) );
  XOR U107352 ( .A(n88131), .B(n88130), .Z(n88132) );
  XOR U107353 ( .A(n88133), .B(n88132), .Z(n88161) );
  IV U107354 ( .A(n88134), .Z(n88135) );
  NOR U107355 ( .A(n88135), .B(n90622), .Z(n88144) );
  IV U107356 ( .A(n88136), .Z(n88142) );
  IV U107357 ( .A(n88137), .Z(n88139) );
  NOR U107358 ( .A(n88139), .B(n88138), .Z(n88140) );
  IV U107359 ( .A(n88140), .Z(n88141) );
  NOR U107360 ( .A(n88142), .B(n88141), .Z(n88143) );
  NOR U107361 ( .A(n88144), .B(n88143), .Z(n88159) );
  IV U107362 ( .A(n88145), .Z(n88146) );
  NOR U107363 ( .A(n88147), .B(n88146), .Z(n88157) );
  IV U107364 ( .A(n88148), .Z(n88149) );
  NOR U107365 ( .A(n88150), .B(n88149), .Z(n88155) );
  IV U107366 ( .A(n88151), .Z(n88153) );
  NOR U107367 ( .A(n88153), .B(n88152), .Z(n88154) );
  XOR U107368 ( .A(n88155), .B(n88154), .Z(n88156) );
  NOR U107369 ( .A(n88157), .B(n88156), .Z(n88158) );
  XOR U107370 ( .A(n88159), .B(n88158), .Z(n88160) );
  XOR U107371 ( .A(n88161), .B(n88160), .Z(n90616) );
  IV U107372 ( .A(n88162), .Z(n88164) );
  NOR U107373 ( .A(n88164), .B(n88163), .Z(n88168) );
  NOR U107374 ( .A(n88166), .B(n88165), .Z(n88167) );
  NOR U107375 ( .A(n88168), .B(n88167), .Z(n90587) );
  NOR U107376 ( .A(n88170), .B(n88169), .Z(n88175) );
  IV U107377 ( .A(n88171), .Z(n88172) );
  NOR U107378 ( .A(n88173), .B(n88172), .Z(n88174) );
  NOR U107379 ( .A(n88175), .B(n88174), .Z(n88185) );
  IV U107380 ( .A(n88176), .Z(n88177) );
  NOR U107381 ( .A(n88178), .B(n88177), .Z(n88183) );
  IV U107382 ( .A(n88179), .Z(n88181) );
  NOR U107383 ( .A(n88181), .B(n88180), .Z(n88182) );
  NOR U107384 ( .A(n88183), .B(n88182), .Z(n88184) );
  XOR U107385 ( .A(n88185), .B(n88184), .Z(n90562) );
  IV U107386 ( .A(n88186), .Z(n88188) );
  NOR U107387 ( .A(n88188), .B(n88187), .Z(n88192) );
  IV U107388 ( .A(n88189), .Z(n88190) );
  NOR U107389 ( .A(n88190), .B(n88195), .Z(n88191) );
  NOR U107390 ( .A(n88192), .B(n88191), .Z(n90548) );
  IV U107391 ( .A(n88196), .Z(n88193) );
  NOR U107392 ( .A(n88193), .B(n88195), .Z(n88200) );
  IV U107393 ( .A(n88194), .Z(n88198) );
  XOR U107394 ( .A(n88196), .B(n88195), .Z(n88197) );
  NOR U107395 ( .A(n88198), .B(n88197), .Z(n88199) );
  NOR U107396 ( .A(n88200), .B(n88199), .Z(n90524) );
  NOR U107397 ( .A(n88202), .B(n88201), .Z(n90505) );
  IV U107398 ( .A(n88206), .Z(n88203) );
  NOR U107399 ( .A(n88203), .B(n88204), .Z(n88211) );
  IV U107400 ( .A(n88204), .Z(n88205) );
  NOR U107401 ( .A(n88206), .B(n88205), .Z(n88209) );
  IV U107402 ( .A(n88207), .Z(n88208) );
  NOR U107403 ( .A(n88209), .B(n88208), .Z(n88210) );
  NOR U107404 ( .A(n88211), .B(n88210), .Z(n90503) );
  IV U107405 ( .A(n88223), .Z(n88225) );
  XOR U107406 ( .A(n88233), .B(n88232), .Z(n90501) );
  IV U107407 ( .A(n88234), .Z(n88235) );
  NOR U107408 ( .A(n88236), .B(n88235), .Z(n90499) );
  IV U107409 ( .A(n88237), .Z(n88239) );
  NOR U107410 ( .A(n88239), .B(n88238), .Z(n90497) );
  IV U107411 ( .A(n88240), .Z(n88241) );
  NOR U107412 ( .A(n88242), .B(n88241), .Z(n90495) );
  NOR U107413 ( .A(n88244), .B(n88243), .Z(n88249) );
  IV U107414 ( .A(n88245), .Z(n88247) );
  NOR U107415 ( .A(n88247), .B(n88246), .Z(n88248) );
  NOR U107416 ( .A(n88249), .B(n88248), .Z(n90493) );
  IV U107417 ( .A(n88250), .Z(n90478) );
  IV U107418 ( .A(n88251), .Z(n88252) );
  NOR U107419 ( .A(n90478), .B(n88252), .Z(n90477) );
  IV U107420 ( .A(n88253), .Z(n88254) );
  NOR U107421 ( .A(n88255), .B(n88254), .Z(n90475) );
  IV U107422 ( .A(n88256), .Z(n88257) );
  NOR U107423 ( .A(n88258), .B(n88257), .Z(n88262) );
  NOR U107424 ( .A(n88260), .B(n88259), .Z(n88261) );
  NOR U107425 ( .A(n88262), .B(n88261), .Z(n88267) );
  IV U107426 ( .A(n88263), .Z(n88265) );
  NOR U107427 ( .A(n88265), .B(n88264), .Z(n88266) );
  XOR U107428 ( .A(n88267), .B(n88266), .Z(n90473) );
  NOR U107429 ( .A(n88269), .B(n88268), .Z(n88274) );
  IV U107430 ( .A(n88270), .Z(n88271) );
  NOR U107431 ( .A(n88272), .B(n88271), .Z(n88273) );
  NOR U107432 ( .A(n88274), .B(n88273), .Z(n90436) );
  NOR U107433 ( .A(n88276), .B(n88275), .Z(n90411) );
  NOR U107434 ( .A(n88278), .B(n88277), .Z(n88283) );
  IV U107435 ( .A(n88279), .Z(n88281) );
  NOR U107436 ( .A(n88281), .B(n88280), .Z(n88282) );
  NOR U107437 ( .A(n88283), .B(n88282), .Z(n88296) );
  NOR U107438 ( .A(n88285), .B(n88284), .Z(n88292) );
  XOR U107439 ( .A(n88286), .B(n88292), .Z(n88294) );
  IV U107440 ( .A(n88287), .Z(n88289) );
  NOR U107441 ( .A(n88289), .B(n88288), .Z(n88290) );
  IV U107442 ( .A(n88290), .Z(n88291) );
  NOR U107443 ( .A(n88292), .B(n88291), .Z(n88293) );
  NOR U107444 ( .A(n88294), .B(n88293), .Z(n88295) );
  XOR U107445 ( .A(n88296), .B(n88295), .Z(n90386) );
  NOR U107446 ( .A(n88298), .B(n88297), .Z(n88303) );
  IV U107447 ( .A(n88299), .Z(n88300) );
  NOR U107448 ( .A(n88301), .B(n88300), .Z(n88302) );
  NOR U107449 ( .A(n88303), .B(n88302), .Z(n90355) );
  NOR U107450 ( .A(n88304), .B(n88305), .Z(n88312) );
  IV U107451 ( .A(n88305), .Z(n88307) );
  NOR U107452 ( .A(n88307), .B(n88306), .Z(n88310) );
  IV U107453 ( .A(n88308), .Z(n88309) );
  NOR U107454 ( .A(n88310), .B(n88309), .Z(n88311) );
  NOR U107455 ( .A(n88312), .B(n88311), .Z(n90353) );
  IV U107456 ( .A(n88313), .Z(n88315) );
  NOR U107457 ( .A(n88315), .B(n88314), .Z(n88319) );
  NOR U107458 ( .A(n88317), .B(n88316), .Z(n88318) );
  NOR U107459 ( .A(n88319), .B(n88318), .Z(n88329) );
  IV U107460 ( .A(n88320), .Z(n88322) );
  NOR U107461 ( .A(n88322), .B(n88321), .Z(n88327) );
  IV U107462 ( .A(n88323), .Z(n88325) );
  NOR U107463 ( .A(n88325), .B(n88324), .Z(n88326) );
  NOR U107464 ( .A(n88327), .B(n88326), .Z(n88328) );
  XOR U107465 ( .A(n88329), .B(n88328), .Z(n88338) );
  NOR U107466 ( .A(n88331), .B(n88330), .Z(n88336) );
  NOR U107467 ( .A(n88336), .B(n88335), .Z(n88337) );
  XOR U107468 ( .A(n88338), .B(n88337), .Z(n88356) );
  IV U107469 ( .A(n88339), .Z(n88340) );
  NOR U107470 ( .A(n88341), .B(n88340), .Z(n88347) );
  IV U107471 ( .A(n88342), .Z(n88345) );
  IV U107472 ( .A(n88343), .Z(n88344) );
  NOR U107473 ( .A(n88345), .B(n88344), .Z(n88346) );
  NOR U107474 ( .A(n88347), .B(n88346), .Z(n88354) );
  IV U107475 ( .A(n88348), .Z(n88350) );
  NOR U107476 ( .A(n88350), .B(n88349), .Z(n88351) );
  NOR U107477 ( .A(n88352), .B(n88351), .Z(n88353) );
  XOR U107478 ( .A(n88354), .B(n88353), .Z(n88355) );
  XOR U107479 ( .A(n88356), .B(n88355), .Z(n90351) );
  IV U107480 ( .A(n88357), .Z(n88359) );
  NOR U107481 ( .A(n88359), .B(n88358), .Z(n88364) );
  IV U107482 ( .A(n88360), .Z(n88362) );
  NOR U107483 ( .A(n88362), .B(n88361), .Z(n88363) );
  NOR U107484 ( .A(n88364), .B(n88363), .Z(n90349) );
  IV U107485 ( .A(n88365), .Z(n88367) );
  NOR U107486 ( .A(n88367), .B(n88366), .Z(n88372) );
  IV U107487 ( .A(n88368), .Z(n88370) );
  NOR U107488 ( .A(n88370), .B(n88369), .Z(n88371) );
  NOR U107489 ( .A(n88372), .B(n88371), .Z(n88376) );
  NOR U107490 ( .A(n88374), .B(n88373), .Z(n88375) );
  XOR U107491 ( .A(n88376), .B(n88375), .Z(n90347) );
  IV U107492 ( .A(n88377), .Z(n88378) );
  NOR U107493 ( .A(n88379), .B(n88378), .Z(n88384) );
  IV U107494 ( .A(n88380), .Z(n88381) );
  NOR U107495 ( .A(n88382), .B(n88381), .Z(n88383) );
  XOR U107496 ( .A(n88384), .B(n88383), .Z(n90345) );
  IV U107497 ( .A(n88385), .Z(n88386) );
  NOR U107498 ( .A(n88387), .B(n88386), .Z(n88391) );
  NOR U107499 ( .A(n88389), .B(n88388), .Z(n88390) );
  NOR U107500 ( .A(n88391), .B(n88390), .Z(n90343) );
  NOR U107501 ( .A(n88393), .B(n88392), .Z(n88395) );
  NOR U107502 ( .A(n88395), .B(n88394), .Z(n90341) );
  IV U107503 ( .A(n88396), .Z(n88397) );
  NOR U107504 ( .A(n88398), .B(n88397), .Z(n88402) );
  IV U107505 ( .A(n88399), .Z(n88400) );
  NOR U107506 ( .A(n88400), .B(n90330), .Z(n88401) );
  NOR U107507 ( .A(n88402), .B(n88401), .Z(n90339) );
  IV U107508 ( .A(n88403), .Z(n88404) );
  NOR U107509 ( .A(n88405), .B(n88404), .Z(n88410) );
  IV U107510 ( .A(n88406), .Z(n88408) );
  NOR U107511 ( .A(n88408), .B(n88407), .Z(n88409) );
  NOR U107512 ( .A(n88410), .B(n88409), .Z(n90310) );
  IV U107513 ( .A(n88411), .Z(n88413) );
  NOR U107514 ( .A(n88413), .B(n88412), .Z(n88415) );
  NOR U107515 ( .A(n88415), .B(n88414), .Z(n90308) );
  IV U107516 ( .A(n88416), .Z(n88418) );
  NOR U107517 ( .A(n88418), .B(n88417), .Z(n88422) );
  NOR U107518 ( .A(n88420), .B(n88419), .Z(n88421) );
  NOR U107519 ( .A(n88422), .B(n88421), .Z(n90306) );
  NOR U107520 ( .A(n88424), .B(n88423), .Z(n90304) );
  IV U107521 ( .A(n88425), .Z(n88426) );
  NOR U107522 ( .A(n88427), .B(n88426), .Z(n88433) );
  IV U107523 ( .A(n88428), .Z(n88431) );
  IV U107524 ( .A(n88429), .Z(n88430) );
  NOR U107525 ( .A(n88431), .B(n88430), .Z(n88432) );
  NOR U107526 ( .A(n88433), .B(n88432), .Z(n90253) );
  NOR U107527 ( .A(n88435), .B(n88434), .Z(n90251) );
  IV U107528 ( .A(n88436), .Z(n88437) );
  NOR U107529 ( .A(n88438), .B(n88437), .Z(n88443) );
  IV U107530 ( .A(n88439), .Z(n88441) );
  NOR U107531 ( .A(n88441), .B(n88440), .Z(n88442) );
  NOR U107532 ( .A(n88443), .B(n88442), .Z(n88452) );
  IV U107533 ( .A(n88444), .Z(n88445) );
  NOR U107534 ( .A(n88446), .B(n88445), .Z(n88450) );
  NOR U107535 ( .A(n88448), .B(n88447), .Z(n88449) );
  NOR U107536 ( .A(n88450), .B(n88449), .Z(n88451) );
  XOR U107537 ( .A(n88452), .B(n88451), .Z(n88462) );
  IV U107538 ( .A(n88453), .Z(n88454) );
  NOR U107539 ( .A(n88455), .B(n88454), .Z(n88460) );
  IV U107540 ( .A(n88456), .Z(n88458) );
  NOR U107541 ( .A(n88458), .B(n88457), .Z(n88459) );
  NOR U107542 ( .A(n88460), .B(n88459), .Z(n88461) );
  XOR U107543 ( .A(n88462), .B(n88461), .Z(n90240) );
  NOR U107544 ( .A(n88464), .B(n88463), .Z(n90238) );
  IV U107545 ( .A(n88465), .Z(n88467) );
  IV U107546 ( .A(n88468), .Z(n88471) );
  NOR U107547 ( .A(n88469), .B(n88499), .Z(n88470) );
  IV U107548 ( .A(n88470), .Z(n88508) );
  IV U107549 ( .A(n88476), .Z(n88480) );
  IV U107550 ( .A(n88477), .Z(n88478) );
  IV U107551 ( .A(n88479), .Z(n88481) );
  IV U107552 ( .A(n88484), .Z(n88486) );
  IV U107553 ( .A(n88487), .Z(n88489) );
  NOR U107554 ( .A(n88489), .B(n88488), .Z(n88493) );
  NOR U107555 ( .A(n88491), .B(n88490), .Z(n88492) );
  IV U107556 ( .A(n88495), .Z(n88496) );
  NOR U107557 ( .A(n88497), .B(n88496), .Z(n88502) );
  IV U107558 ( .A(n88498), .Z(n88500) );
  NOR U107559 ( .A(n88500), .B(n88499), .Z(n88501) );
  NOR U107560 ( .A(n88502), .B(n88501), .Z(n90234) );
  IV U107561 ( .A(n88503), .Z(n88505) );
  NOR U107562 ( .A(n88505), .B(n88504), .Z(n88510) );
  IV U107563 ( .A(n88506), .Z(n88507) );
  NOR U107564 ( .A(n88508), .B(n88507), .Z(n88509) );
  XOR U107565 ( .A(n88510), .B(n88509), .Z(n90232) );
  IV U107566 ( .A(n88511), .Z(n88513) );
  NOR U107567 ( .A(n88513), .B(n88512), .Z(n88517) );
  NOR U107568 ( .A(n88515), .B(n88514), .Z(n88516) );
  NOR U107569 ( .A(n88517), .B(n88516), .Z(n88527) );
  IV U107570 ( .A(n88518), .Z(n88520) );
  NOR U107571 ( .A(n88520), .B(n88519), .Z(n88525) );
  IV U107572 ( .A(n88521), .Z(n88523) );
  NOR U107573 ( .A(n88523), .B(n88522), .Z(n88524) );
  NOR U107574 ( .A(n88525), .B(n88524), .Z(n88526) );
  XOR U107575 ( .A(n88527), .B(n88526), .Z(n90230) );
  IV U107576 ( .A(n88528), .Z(n88529) );
  NOR U107577 ( .A(n88529), .B(n90216), .Z(n90228) );
  IV U107578 ( .A(n88532), .Z(n88530) );
  NOR U107579 ( .A(n88531), .B(n88530), .Z(n88537) );
  NOR U107580 ( .A(n88533), .B(n88532), .Z(n88535) );
  NOR U107581 ( .A(n88535), .B(n88534), .Z(n88536) );
  NOR U107582 ( .A(n88537), .B(n88536), .Z(n90226) );
  NOR U107583 ( .A(n88539), .B(n88538), .Z(n88544) );
  IV U107584 ( .A(n88540), .Z(n88541) );
  NOR U107585 ( .A(n88542), .B(n88541), .Z(n88543) );
  NOR U107586 ( .A(n88544), .B(n88543), .Z(n90224) );
  IV U107587 ( .A(n88545), .Z(n88547) );
  NOR U107588 ( .A(n88547), .B(n88546), .Z(n88552) );
  IV U107589 ( .A(n88548), .Z(n88550) );
  NOR U107590 ( .A(n88550), .B(n88549), .Z(n88551) );
  NOR U107591 ( .A(n88552), .B(n88551), .Z(n90175) );
  NOR U107592 ( .A(n88554), .B(n88553), .Z(n88559) );
  IV U107593 ( .A(n88555), .Z(n88556) );
  NOR U107594 ( .A(n88557), .B(n88556), .Z(n88558) );
  NOR U107595 ( .A(n88559), .B(n88558), .Z(n88569) );
  IV U107596 ( .A(n88560), .Z(n88562) );
  NOR U107597 ( .A(n88562), .B(n88561), .Z(n88567) );
  IV U107598 ( .A(n88563), .Z(n88564) );
  NOR U107599 ( .A(n88565), .B(n88564), .Z(n88566) );
  NOR U107600 ( .A(n88567), .B(n88566), .Z(n88568) );
  XOR U107601 ( .A(n88569), .B(n88568), .Z(n90173) );
  IV U107602 ( .A(n88570), .Z(n88572) );
  NOR U107603 ( .A(n88572), .B(n88571), .Z(n88577) );
  IV U107604 ( .A(n88573), .Z(n88574) );
  NOR U107605 ( .A(n88575), .B(n88574), .Z(n88576) );
  NOR U107606 ( .A(n88577), .B(n88576), .Z(n88583) );
  NOR U107607 ( .A(n88579), .B(n88578), .Z(n88581) );
  NOR U107608 ( .A(n88581), .B(n88580), .Z(n88582) );
  XOR U107609 ( .A(n88583), .B(n88582), .Z(n88593) );
  IV U107610 ( .A(n88584), .Z(n88586) );
  NOR U107611 ( .A(n88586), .B(n88585), .Z(n88591) );
  IV U107612 ( .A(n88587), .Z(n88589) );
  NOR U107613 ( .A(n88589), .B(n88588), .Z(n88590) );
  NOR U107614 ( .A(n88591), .B(n88590), .Z(n88592) );
  XOR U107615 ( .A(n88593), .B(n88592), .Z(n90171) );
  IV U107616 ( .A(n88594), .Z(n88595) );
  NOR U107617 ( .A(n88596), .B(n88595), .Z(n90169) );
  IV U107618 ( .A(n88597), .Z(n88598) );
  NOR U107619 ( .A(n88599), .B(n88598), .Z(n88604) );
  IV U107620 ( .A(n88600), .Z(n88601) );
  NOR U107621 ( .A(n88602), .B(n88601), .Z(n88603) );
  NOR U107622 ( .A(n88604), .B(n88603), .Z(n90167) );
  IV U107623 ( .A(n88605), .Z(n88606) );
  NOR U107624 ( .A(n88607), .B(n88606), .Z(n88612) );
  IV U107625 ( .A(n88608), .Z(n88610) );
  NOR U107626 ( .A(n88610), .B(n88609), .Z(n88611) );
  NOR U107627 ( .A(n88612), .B(n88611), .Z(n90106) );
  IV U107628 ( .A(n88613), .Z(n88614) );
  NOR U107629 ( .A(n88614), .B(n90112), .Z(n88618) );
  IV U107630 ( .A(n88615), .Z(n88616) );
  NOR U107631 ( .A(n88617), .B(n88616), .Z(n88624) );
  XOR U107632 ( .A(n88618), .B(n88624), .Z(n88626) );
  IV U107633 ( .A(n88619), .Z(n88620) );
  NOR U107634 ( .A(n88621), .B(n88620), .Z(n88622) );
  IV U107635 ( .A(n88622), .Z(n88623) );
  NOR U107636 ( .A(n88624), .B(n88623), .Z(n88625) );
  NOR U107637 ( .A(n88626), .B(n88625), .Z(n90104) );
  IV U107638 ( .A(n88627), .Z(n88629) );
  NOR U107639 ( .A(n88629), .B(n88628), .Z(n88634) );
  IV U107640 ( .A(n88630), .Z(n88631) );
  NOR U107641 ( .A(n88632), .B(n88631), .Z(n88633) );
  NOR U107642 ( .A(n88634), .B(n88633), .Z(n90092) );
  NOR U107643 ( .A(n88636), .B(n88635), .Z(n90090) );
  IV U107644 ( .A(n88637), .Z(n88638) );
  NOR U107645 ( .A(n88638), .B(n88642), .Z(n88639) );
  NOR U107646 ( .A(n88640), .B(n88639), .Z(n90088) );
  IV U107647 ( .A(n88641), .Z(n88643) );
  NOR U107648 ( .A(n88643), .B(n88642), .Z(n88653) );
  XOR U107649 ( .A(n88646), .B(n88647), .Z(n88645) );
  NOR U107650 ( .A(n88645), .B(n88644), .Z(n88650) );
  IV U107651 ( .A(n88646), .Z(n88648) );
  NOR U107652 ( .A(n88648), .B(n88647), .Z(n88649) );
  NOR U107653 ( .A(n88650), .B(n88649), .Z(n88651) );
  IV U107654 ( .A(n88651), .Z(n88652) );
  NOR U107655 ( .A(n88653), .B(n88652), .Z(n90057) );
  NOR U107656 ( .A(n88655), .B(n88654), .Z(n88656) );
  NOR U107657 ( .A(n88656), .B(n88657), .Z(n88660) );
  IV U107658 ( .A(n88657), .Z(n90061) );
  NOR U107659 ( .A(n90061), .B(n88658), .Z(n88659) );
  NOR U107660 ( .A(n88660), .B(n88659), .Z(n90055) );
  IV U107661 ( .A(n88661), .Z(n88663) );
  NOR U107662 ( .A(n88663), .B(n88662), .Z(n88668) );
  IV U107663 ( .A(n88664), .Z(n88666) );
  NOR U107664 ( .A(n88666), .B(n88665), .Z(n88667) );
  NOR U107665 ( .A(n88668), .B(n88667), .Z(n90053) );
  IV U107666 ( .A(n88679), .Z(n88680) );
  NOR U107667 ( .A(n88681), .B(n88680), .Z(n88685) );
  NOR U107668 ( .A(n88683), .B(n88682), .Z(n88684) );
  NOR U107669 ( .A(n88685), .B(n88684), .Z(n88686) );
  XOR U107670 ( .A(n88687), .B(n88686), .Z(n88699) );
  NOR U107671 ( .A(n88689), .B(n88688), .Z(n88697) );
  IV U107672 ( .A(n88689), .Z(n88691) );
  NOR U107673 ( .A(n88691), .B(n88690), .Z(n88695) );
  XOR U107674 ( .A(n88693), .B(n88692), .Z(n88694) );
  NOR U107675 ( .A(n88695), .B(n88694), .Z(n88696) );
  NOR U107676 ( .A(n88697), .B(n88696), .Z(n88698) );
  XOR U107677 ( .A(n88699), .B(n88698), .Z(n90036) );
  IV U107678 ( .A(n88700), .Z(n88702) );
  NOR U107679 ( .A(n88702), .B(n88701), .Z(n88707) );
  IV U107680 ( .A(n88703), .Z(n88705) );
  NOR U107681 ( .A(n88705), .B(n88704), .Z(n88706) );
  NOR U107682 ( .A(n88707), .B(n88706), .Z(n89997) );
  IV U107683 ( .A(n88708), .Z(n88709) );
  NOR U107684 ( .A(n88709), .B(n89957), .Z(n88713) );
  NOR U107685 ( .A(n88711), .B(n88710), .Z(n88712) );
  NOR U107686 ( .A(n88713), .B(n88712), .Z(n88722) );
  IV U107687 ( .A(n88714), .Z(n88716) );
  NOR U107688 ( .A(n88716), .B(n88715), .Z(n88720) );
  NOR U107689 ( .A(n88718), .B(n88717), .Z(n88719) );
  NOR U107690 ( .A(n88720), .B(n88719), .Z(n88721) );
  XOR U107691 ( .A(n88722), .B(n88721), .Z(n88737) );
  IV U107692 ( .A(n88723), .Z(n88725) );
  NOR U107693 ( .A(n88725), .B(n88724), .Z(n88735) );
  IV U107694 ( .A(n88726), .Z(n88728) );
  NOR U107695 ( .A(n88728), .B(n88727), .Z(n88733) );
  IV U107696 ( .A(n88729), .Z(n88731) );
  NOR U107697 ( .A(n88731), .B(n88730), .Z(n88732) );
  NOR U107698 ( .A(n88733), .B(n88732), .Z(n88734) );
  XOR U107699 ( .A(n88735), .B(n88734), .Z(n88736) );
  XOR U107700 ( .A(n88737), .B(n88736), .Z(n89954) );
  IV U107701 ( .A(n88738), .Z(n88739) );
  NOR U107702 ( .A(n88740), .B(n88739), .Z(n89952) );
  IV U107703 ( .A(n88741), .Z(n88743) );
  NOR U107704 ( .A(n88743), .B(n88742), .Z(n88747) );
  NOR U107705 ( .A(n88745), .B(n88744), .Z(n88746) );
  NOR U107706 ( .A(n88747), .B(n88746), .Z(n89950) );
  IV U107707 ( .A(n88748), .Z(n88749) );
  NOR U107708 ( .A(n88750), .B(n88749), .Z(n88754) );
  NOR U107709 ( .A(n88752), .B(n88751), .Z(n88753) );
  NOR U107710 ( .A(n88754), .B(n88753), .Z(n89924) );
  NOR U107711 ( .A(n88756), .B(n88755), .Z(n89922) );
  IV U107712 ( .A(n88757), .Z(n88759) );
  NOR U107713 ( .A(n88759), .B(n88758), .Z(n88763) );
  NOR U107714 ( .A(n88761), .B(n88760), .Z(n88762) );
  NOR U107715 ( .A(n88763), .B(n88762), .Z(n89920) );
  IV U107716 ( .A(n88764), .Z(n88765) );
  NOR U107717 ( .A(n88765), .B(n89891), .Z(n88771) );
  IV U107718 ( .A(n88766), .Z(n88769) );
  IV U107719 ( .A(n88767), .Z(n88768) );
  NOR U107720 ( .A(n88769), .B(n88768), .Z(n88770) );
  NOR U107721 ( .A(n88771), .B(n88770), .Z(n89918) );
  IV U107722 ( .A(n88772), .Z(n88773) );
  NOR U107723 ( .A(n88774), .B(n88773), .Z(n88779) );
  IV U107724 ( .A(n88775), .Z(n88777) );
  NOR U107725 ( .A(n88777), .B(n88776), .Z(n88778) );
  NOR U107726 ( .A(n88779), .B(n88778), .Z(n89865) );
  IV U107727 ( .A(n88792), .Z(n88796) );
  XOR U107728 ( .A(n88795), .B(n88796), .Z(n88794) );
  NOR U107729 ( .A(n88794), .B(n88793), .Z(n88799) );
  IV U107730 ( .A(n88795), .Z(n88797) );
  NOR U107731 ( .A(n88797), .B(n88796), .Z(n88798) );
  NOR U107732 ( .A(n88799), .B(n88798), .Z(n89787) );
  IV U107733 ( .A(n88800), .Z(n88801) );
  NOR U107734 ( .A(n88802), .B(n88801), .Z(n88803) );
  NOR U107735 ( .A(n88804), .B(n88803), .Z(n89785) );
  IV U107736 ( .A(n88805), .Z(n88807) );
  NOR U107737 ( .A(n88807), .B(n88806), .Z(n88812) );
  IV U107738 ( .A(n88808), .Z(n88810) );
  NOR U107739 ( .A(n88810), .B(n88809), .Z(n88811) );
  NOR U107740 ( .A(n88812), .B(n88811), .Z(n88822) );
  IV U107741 ( .A(n88813), .Z(n88815) );
  NOR U107742 ( .A(n88815), .B(n88814), .Z(n88820) );
  IV U107743 ( .A(n88816), .Z(n88817) );
  NOR U107744 ( .A(n88818), .B(n88817), .Z(n88819) );
  NOR U107745 ( .A(n88820), .B(n88819), .Z(n88821) );
  XOR U107746 ( .A(n88822), .B(n88821), .Z(n89783) );
  NOR U107747 ( .A(n88824), .B(n88823), .Z(n88825) );
  NOR U107748 ( .A(n88826), .B(n88825), .Z(n88836) );
  IV U107749 ( .A(n88827), .Z(n88828) );
  NOR U107750 ( .A(n88829), .B(n88828), .Z(n88834) );
  IV U107751 ( .A(n88830), .Z(n88831) );
  NOR U107752 ( .A(n88832), .B(n88831), .Z(n88833) );
  NOR U107753 ( .A(n88834), .B(n88833), .Z(n88835) );
  XOR U107754 ( .A(n88836), .B(n88835), .Z(n88846) );
  NOR U107755 ( .A(n88838), .B(n88837), .Z(n88844) );
  IV U107756 ( .A(n88839), .Z(n88842) );
  IV U107757 ( .A(n88840), .Z(n88841) );
  NOR U107758 ( .A(n88842), .B(n88841), .Z(n88843) );
  NOR U107759 ( .A(n88844), .B(n88843), .Z(n88845) );
  XOR U107760 ( .A(n88846), .B(n88845), .Z(n89781) );
  IV U107761 ( .A(n88847), .Z(n88849) );
  NOR U107762 ( .A(n88849), .B(n88848), .Z(n88850) );
  NOR U107763 ( .A(n88851), .B(n88850), .Z(n89779) );
  IV U107764 ( .A(n88855), .Z(n88852) );
  NOR U107765 ( .A(n88852), .B(n88853), .Z(n88860) );
  IV U107766 ( .A(n88853), .Z(n88854) );
  NOR U107767 ( .A(n88855), .B(n88854), .Z(n88858) );
  IV U107768 ( .A(n88856), .Z(n88857) );
  NOR U107769 ( .A(n88858), .B(n88857), .Z(n88859) );
  NOR U107770 ( .A(n88860), .B(n88859), .Z(n88875) );
  IV U107771 ( .A(n88861), .Z(n88862) );
  NOR U107772 ( .A(n88862), .B(n88877), .Z(n88873) );
  IV U107773 ( .A(n88863), .Z(n88864) );
  NOR U107774 ( .A(n88865), .B(n88864), .Z(n88870) );
  IV U107775 ( .A(n88866), .Z(n88868) );
  NOR U107776 ( .A(n88868), .B(n88867), .Z(n88869) );
  NOR U107777 ( .A(n88870), .B(n88869), .Z(n88871) );
  IV U107778 ( .A(n88871), .Z(n88872) );
  NOR U107779 ( .A(n88873), .B(n88872), .Z(n88874) );
  XOR U107780 ( .A(n88875), .B(n88874), .Z(n88888) );
  IV U107781 ( .A(n88876), .Z(n88878) );
  NOR U107782 ( .A(n88878), .B(n88877), .Z(n88883) );
  IV U107783 ( .A(n88879), .Z(n88881) );
  NOR U107784 ( .A(n88881), .B(n88880), .Z(n88882) );
  NOR U107785 ( .A(n88883), .B(n88882), .Z(n88884) );
  IV U107786 ( .A(n88884), .Z(n88885) );
  NOR U107787 ( .A(n88886), .B(n88885), .Z(n88887) );
  XOR U107788 ( .A(n88888), .B(n88887), .Z(n89777) );
  IV U107789 ( .A(n88889), .Z(n88890) );
  NOR U107790 ( .A(n88891), .B(n88890), .Z(n89775) );
  NOR U107791 ( .A(n88893), .B(n88892), .Z(n88895) );
  NOR U107792 ( .A(n88895), .B(n88894), .Z(n88905) );
  IV U107793 ( .A(n88896), .Z(n88898) );
  NOR U107794 ( .A(n88898), .B(n88897), .Z(n88903) );
  IV U107795 ( .A(n88899), .Z(n88900) );
  NOR U107796 ( .A(n88901), .B(n88900), .Z(n88902) );
  NOR U107797 ( .A(n88903), .B(n88902), .Z(n88904) );
  XOR U107798 ( .A(n88905), .B(n88904), .Z(n88915) );
  IV U107799 ( .A(n88906), .Z(n88908) );
  NOR U107800 ( .A(n88908), .B(n88907), .Z(n88913) );
  IV U107801 ( .A(n88909), .Z(n88911) );
  NOR U107802 ( .A(n88911), .B(n88910), .Z(n88912) );
  NOR U107803 ( .A(n88913), .B(n88912), .Z(n88914) );
  XOR U107804 ( .A(n88915), .B(n88914), .Z(n88935) );
  IV U107805 ( .A(n88916), .Z(n88918) );
  NOR U107806 ( .A(n88918), .B(n88917), .Z(n88923) );
  IV U107807 ( .A(n88919), .Z(n88921) );
  NOR U107808 ( .A(n88921), .B(n88920), .Z(n88922) );
  NOR U107809 ( .A(n88923), .B(n88922), .Z(n88933) );
  IV U107810 ( .A(n88924), .Z(n88926) );
  NOR U107811 ( .A(n88926), .B(n88925), .Z(n88931) );
  IV U107812 ( .A(n88927), .Z(n88929) );
  NOR U107813 ( .A(n88929), .B(n88928), .Z(n88930) );
  NOR U107814 ( .A(n88931), .B(n88930), .Z(n88932) );
  XOR U107815 ( .A(n88933), .B(n88932), .Z(n88934) );
  XOR U107816 ( .A(n88935), .B(n88934), .Z(n89773) );
  IV U107817 ( .A(n88936), .Z(n88937) );
  NOR U107818 ( .A(n88938), .B(n88937), .Z(n88949) );
  IV U107819 ( .A(n88939), .Z(n88941) );
  NOR U107820 ( .A(n88941), .B(n88940), .Z(n88946) );
  IV U107821 ( .A(n88942), .Z(n88943) );
  NOR U107822 ( .A(n88944), .B(n88943), .Z(n88945) );
  NOR U107823 ( .A(n88946), .B(n88945), .Z(n88947) );
  IV U107824 ( .A(n88947), .Z(n88948) );
  NOR U107825 ( .A(n88949), .B(n88948), .Z(n89752) );
  IV U107826 ( .A(n88950), .Z(n88952) );
  NOR U107827 ( .A(n88952), .B(n88951), .Z(n89750) );
  IV U107828 ( .A(n88953), .Z(n88955) );
  IV U107829 ( .A(n88954), .Z(n89690) );
  NOR U107830 ( .A(n88955), .B(n89690), .Z(n88960) );
  IV U107831 ( .A(n88956), .Z(n88958) );
  NOR U107832 ( .A(n88958), .B(n88957), .Z(n88959) );
  NOR U107833 ( .A(n88960), .B(n88959), .Z(n89732) );
  NOR U107834 ( .A(n88961), .B(n89671), .Z(n88969) );
  XOR U107835 ( .A(n89670), .B(n88962), .Z(n88963) );
  NOR U107836 ( .A(n88964), .B(n88963), .Z(n88967) );
  IV U107837 ( .A(n88965), .Z(n88966) );
  NOR U107838 ( .A(n88967), .B(n88966), .Z(n88968) );
  NOR U107839 ( .A(n88969), .B(n88968), .Z(n89688) );
  IV U107840 ( .A(n88970), .Z(n88971) );
  NOR U107841 ( .A(n88972), .B(n88971), .Z(n88977) );
  IV U107842 ( .A(n88973), .Z(n88975) );
  NOR U107843 ( .A(n88975), .B(n88974), .Z(n88976) );
  NOR U107844 ( .A(n88977), .B(n88976), .Z(n89631) );
  NOR U107845 ( .A(n88979), .B(n88978), .Z(n88981) );
  NOR U107846 ( .A(n88981), .B(n88980), .Z(n89629) );
  IV U107847 ( .A(n88982), .Z(n88984) );
  NOR U107848 ( .A(n88984), .B(n88983), .Z(n88989) );
  IV U107849 ( .A(n88985), .Z(n88987) );
  NOR U107850 ( .A(n88987), .B(n88986), .Z(n88988) );
  NOR U107851 ( .A(n88989), .B(n88988), .Z(n88998) );
  NOR U107852 ( .A(n88991), .B(n88990), .Z(n88996) );
  IV U107853 ( .A(n88992), .Z(n88993) );
  NOR U107854 ( .A(n88994), .B(n88993), .Z(n88995) );
  NOR U107855 ( .A(n88996), .B(n88995), .Z(n88997) );
  XOR U107856 ( .A(n88998), .B(n88997), .Z(n89026) );
  IV U107857 ( .A(n88999), .Z(n89000) );
  NOR U107858 ( .A(n89001), .B(n89000), .Z(n89012) );
  IV U107859 ( .A(n89002), .Z(n89003) );
  NOR U107860 ( .A(n89004), .B(n89003), .Z(n89009) );
  IV U107861 ( .A(n89005), .Z(n89006) );
  NOR U107862 ( .A(n89007), .B(n89006), .Z(n89008) );
  NOR U107863 ( .A(n89009), .B(n89008), .Z(n89010) );
  IV U107864 ( .A(n89010), .Z(n89011) );
  NOR U107865 ( .A(n89012), .B(n89011), .Z(n89024) );
  IV U107866 ( .A(n89013), .Z(n89014) );
  NOR U107867 ( .A(n89015), .B(n89014), .Z(n89022) );
  NOR U107868 ( .A(n89016), .B(n89594), .Z(n89017) );
  IV U107869 ( .A(n89017), .Z(n89020) );
  IV U107870 ( .A(n89018), .Z(n89019) );
  NOR U107871 ( .A(n89020), .B(n89019), .Z(n89021) );
  NOR U107872 ( .A(n89022), .B(n89021), .Z(n89023) );
  XOR U107873 ( .A(n89024), .B(n89023), .Z(n89025) );
  XOR U107874 ( .A(n89026), .B(n89025), .Z(n89591) );
  NOR U107875 ( .A(n89028), .B(n89027), .Z(n89030) );
  NOR U107876 ( .A(n89030), .B(n89029), .Z(n89589) );
  NOR U107877 ( .A(n89032), .B(n89031), .Z(n89037) );
  IV U107878 ( .A(n89033), .Z(n89034) );
  NOR U107879 ( .A(n89035), .B(n89034), .Z(n89036) );
  NOR U107880 ( .A(n89037), .B(n89036), .Z(n89587) );
  IV U107881 ( .A(n89038), .Z(n89039) );
  NOR U107882 ( .A(n89040), .B(n89039), .Z(n89046) );
  NOR U107883 ( .A(n89042), .B(n89041), .Z(n89043) );
  NOR U107884 ( .A(n89044), .B(n89043), .Z(n89045) );
  NOR U107885 ( .A(n89046), .B(n89045), .Z(n89585) );
  IV U107886 ( .A(n89047), .Z(n89048) );
  NOR U107887 ( .A(n89049), .B(n89048), .Z(n89054) );
  IV U107888 ( .A(n89050), .Z(n89051) );
  NOR U107889 ( .A(n89052), .B(n89051), .Z(n89053) );
  NOR U107890 ( .A(n89054), .B(n89053), .Z(n89583) );
  IV U107891 ( .A(n89055), .Z(n89057) );
  NOR U107892 ( .A(n89057), .B(n89056), .Z(n89062) );
  IV U107893 ( .A(n89058), .Z(n89060) );
  NOR U107894 ( .A(n89060), .B(n89059), .Z(n89061) );
  NOR U107895 ( .A(n89062), .B(n89061), .Z(n89552) );
  IV U107896 ( .A(n89063), .Z(n89064) );
  NOR U107897 ( .A(n89065), .B(n89064), .Z(n89070) );
  IV U107898 ( .A(n89066), .Z(n89068) );
  NOR U107899 ( .A(n89068), .B(n89067), .Z(n89069) );
  NOR U107900 ( .A(n89070), .B(n89069), .Z(n89535) );
  XOR U107901 ( .A(n89073), .B(n89074), .Z(n89072) );
  NOR U107902 ( .A(n89072), .B(n89071), .Z(n89077) );
  IV U107903 ( .A(n89073), .Z(n89075) );
  NOR U107904 ( .A(n89075), .B(n89074), .Z(n89076) );
  NOR U107905 ( .A(n89077), .B(n89076), .Z(n89533) );
  IV U107906 ( .A(n89078), .Z(n89080) );
  NOR U107907 ( .A(n89080), .B(n89079), .Z(n89085) );
  IV U107908 ( .A(n89081), .Z(n89083) );
  NOR U107909 ( .A(n89083), .B(n89082), .Z(n89084) );
  NOR U107910 ( .A(n89085), .B(n89084), .Z(n89525) );
  NOR U107911 ( .A(n89087), .B(n89086), .Z(n89097) );
  IV U107912 ( .A(n89088), .Z(n89089) );
  NOR U107913 ( .A(n89090), .B(n89089), .Z(n89094) );
  NOR U107914 ( .A(n89092), .B(n89091), .Z(n89093) );
  NOR U107915 ( .A(n89094), .B(n89093), .Z(n89095) );
  IV U107916 ( .A(n89095), .Z(n89096) );
  NOR U107917 ( .A(n89097), .B(n89096), .Z(n89523) );
  IV U107918 ( .A(n89098), .Z(n89099) );
  NOR U107919 ( .A(n89100), .B(n89099), .Z(n89110) );
  IV U107920 ( .A(n89101), .Z(n89108) );
  NOR U107921 ( .A(n89103), .B(n89102), .Z(n89104) );
  IV U107922 ( .A(n89104), .Z(n89105) );
  NOR U107923 ( .A(n89106), .B(n89105), .Z(n89107) );
  IV U107924 ( .A(n89107), .Z(n89112) );
  NOR U107925 ( .A(n89108), .B(n89112), .Z(n89109) );
  NOR U107926 ( .A(n89110), .B(n89109), .Z(n89521) );
  IV U107927 ( .A(n89111), .Z(n89113) );
  NOR U107928 ( .A(n89113), .B(n89112), .Z(n89519) );
  XOR U107929 ( .A(n89116), .B(n89117), .Z(n89115) );
  NOR U107930 ( .A(n89115), .B(n89114), .Z(n89120) );
  IV U107931 ( .A(n89116), .Z(n89118) );
  NOR U107932 ( .A(n89118), .B(n89117), .Z(n89119) );
  NOR U107933 ( .A(n89120), .B(n89119), .Z(n89121) );
  IV U107934 ( .A(n89121), .Z(n89126) );
  IV U107935 ( .A(n89122), .Z(n89124) );
  NOR U107936 ( .A(n89124), .B(n89123), .Z(n89125) );
  NOR U107937 ( .A(n89126), .B(n89125), .Z(n89488) );
  IV U107938 ( .A(n89127), .Z(n89129) );
  NOR U107939 ( .A(n89129), .B(n89128), .Z(n89468) );
  IV U107940 ( .A(n89130), .Z(n89131) );
  NOR U107941 ( .A(n89132), .B(n89131), .Z(n89135) );
  NOR U107942 ( .A(n89134), .B(n89133), .Z(n89140) );
  XOR U107943 ( .A(n89135), .B(n89140), .Z(n89142) );
  NOR U107944 ( .A(n89137), .B(n89136), .Z(n89138) );
  IV U107945 ( .A(n89138), .Z(n89139) );
  NOR U107946 ( .A(n89140), .B(n89139), .Z(n89141) );
  NOR U107947 ( .A(n89142), .B(n89141), .Z(n89451) );
  IV U107948 ( .A(n89143), .Z(n89145) );
  NOR U107949 ( .A(n89145), .B(n89144), .Z(n89449) );
  IV U107950 ( .A(n89146), .Z(n89147) );
  NOR U107951 ( .A(n89148), .B(n89147), .Z(n89153) );
  IV U107952 ( .A(n89149), .Z(n89151) );
  NOR U107953 ( .A(n89151), .B(n89150), .Z(n89152) );
  NOR U107954 ( .A(n89153), .B(n89152), .Z(n89447) );
  IV U107955 ( .A(n89154), .Z(n89156) );
  NOR U107956 ( .A(n89156), .B(n89155), .Z(n89161) );
  IV U107957 ( .A(n89157), .Z(n89159) );
  NOR U107958 ( .A(n89159), .B(n89158), .Z(n89160) );
  NOR U107959 ( .A(n89161), .B(n89160), .Z(n89171) );
  IV U107960 ( .A(n89162), .Z(n89163) );
  NOR U107961 ( .A(n89164), .B(n89163), .Z(n89169) );
  IV U107962 ( .A(n89165), .Z(n89167) );
  NOR U107963 ( .A(n89167), .B(n89166), .Z(n89168) );
  NOR U107964 ( .A(n89169), .B(n89168), .Z(n89170) );
  XOR U107965 ( .A(n89171), .B(n89170), .Z(n89445) );
  IV U107966 ( .A(n89172), .Z(n89173) );
  NOR U107967 ( .A(n89174), .B(n89173), .Z(n89175) );
  NOR U107968 ( .A(n89176), .B(n89175), .Z(n89443) );
  IV U107969 ( .A(n89177), .Z(n89179) );
  NOR U107970 ( .A(n89179), .B(n89178), .Z(n89184) );
  IV U107971 ( .A(n89180), .Z(n89182) );
  NOR U107972 ( .A(n89182), .B(n89181), .Z(n89183) );
  NOR U107973 ( .A(n89184), .B(n89183), .Z(n89411) );
  IV U107974 ( .A(n89185), .Z(n89186) );
  NOR U107975 ( .A(n89187), .B(n89186), .Z(n89192) );
  IV U107976 ( .A(n89188), .Z(n89190) );
  NOR U107977 ( .A(n89190), .B(n89189), .Z(n89191) );
  NOR U107978 ( .A(n89192), .B(n89191), .Z(n89390) );
  IV U107979 ( .A(n89193), .Z(n89194) );
  NOR U107980 ( .A(n89195), .B(n89194), .Z(n89200) );
  IV U107981 ( .A(n89196), .Z(n89198) );
  NOR U107982 ( .A(n89198), .B(n89197), .Z(n89199) );
  NOR U107983 ( .A(n89200), .B(n89199), .Z(n89388) );
  IV U107984 ( .A(n89205), .Z(n89201) );
  NOR U107985 ( .A(n89202), .B(n89201), .Z(n89203) );
  NOR U107986 ( .A(n89204), .B(n89203), .Z(n89208) );
  NOR U107987 ( .A(n89206), .B(n89205), .Z(n89207) );
  NOR U107988 ( .A(n89208), .B(n89207), .Z(n89368) );
  IV U107989 ( .A(n89213), .Z(n89209) );
  NOR U107990 ( .A(n89210), .B(n89209), .Z(n89211) );
  NOR U107991 ( .A(n89212), .B(n89211), .Z(n89216) );
  NOR U107992 ( .A(n89214), .B(n89213), .Z(n89215) );
  NOR U107993 ( .A(n89216), .B(n89215), .Z(n89366) );
  NOR U107994 ( .A(n89218), .B(n89217), .Z(n89223) );
  IV U107995 ( .A(n89219), .Z(n89221) );
  NOR U107996 ( .A(n89221), .B(n89220), .Z(n89222) );
  NOR U107997 ( .A(n89223), .B(n89222), .Z(n89364) );
  IV U107998 ( .A(n89224), .Z(n89226) );
  NOR U107999 ( .A(n89226), .B(n89225), .Z(n89231) );
  IV U108000 ( .A(n89227), .Z(n89229) );
  NOR U108001 ( .A(n89229), .B(n89228), .Z(n89230) );
  NOR U108002 ( .A(n89231), .B(n89230), .Z(n89362) );
  IV U108003 ( .A(n89232), .Z(n89233) );
  NOR U108004 ( .A(n89234), .B(n89233), .Z(n89360) );
  IV U108005 ( .A(n89235), .Z(n89237) );
  NOR U108006 ( .A(n89237), .B(n89236), .Z(n89241) );
  NOR U108007 ( .A(n89239), .B(n89238), .Z(n89240) );
  NOR U108008 ( .A(n89241), .B(n89240), .Z(n89253) );
  IV U108009 ( .A(n89242), .Z(n89244) );
  NOR U108010 ( .A(n89244), .B(n89243), .Z(n89251) );
  IV U108011 ( .A(n89245), .Z(n89247) );
  NOR U108012 ( .A(n89247), .B(n89246), .Z(n89249) );
  NOR U108013 ( .A(n89249), .B(n89248), .Z(n89250) );
  XOR U108014 ( .A(n89251), .B(n89250), .Z(n89252) );
  XOR U108015 ( .A(n89253), .B(n89252), .Z(n89272) );
  IV U108016 ( .A(n89254), .Z(n89255) );
  NOR U108017 ( .A(n89256), .B(n89255), .Z(n89261) );
  IV U108018 ( .A(n89257), .Z(n89259) );
  NOR U108019 ( .A(n89259), .B(n89258), .Z(n89260) );
  NOR U108020 ( .A(n89261), .B(n89260), .Z(n89270) );
  NOR U108021 ( .A(n89263), .B(n89262), .Z(n89268) );
  IV U108022 ( .A(n89264), .Z(n89266) );
  NOR U108023 ( .A(n89266), .B(n89265), .Z(n89267) );
  NOR U108024 ( .A(n89268), .B(n89267), .Z(n89269) );
  XOR U108025 ( .A(n89270), .B(n89269), .Z(n89271) );
  XOR U108026 ( .A(n89272), .B(n89271), .Z(n89358) );
  XOR U108027 ( .A(n89275), .B(n89276), .Z(n89274) );
  NOR U108028 ( .A(n89274), .B(n89273), .Z(n89279) );
  IV U108029 ( .A(n89275), .Z(n89277) );
  NOR U108030 ( .A(n89277), .B(n89276), .Z(n89278) );
  NOR U108031 ( .A(n89279), .B(n89278), .Z(n89356) );
  IV U108032 ( .A(n89280), .Z(n89282) );
  NOR U108033 ( .A(n89282), .B(n89281), .Z(n89286) );
  NOR U108034 ( .A(n89284), .B(n89283), .Z(n89285) );
  NOR U108035 ( .A(n89286), .B(n89285), .Z(n89344) );
  NOR U108036 ( .A(n89288), .B(n89287), .Z(n89289) );
  IV U108037 ( .A(n89289), .Z(n89290) );
  NOR U108038 ( .A(n89291), .B(n89290), .Z(n89292) );
  NOR U108039 ( .A(n89293), .B(n89292), .Z(n89303) );
  IV U108040 ( .A(n89294), .Z(n89295) );
  NOR U108041 ( .A(n89296), .B(n89295), .Z(n89301) );
  IV U108042 ( .A(n89296), .Z(n89299) );
  IV U108043 ( .A(n89297), .Z(n89298) );
  NOR U108044 ( .A(n89299), .B(n89298), .Z(n89300) );
  NOR U108045 ( .A(n89301), .B(n89300), .Z(n89302) );
  XOR U108046 ( .A(n89303), .B(n89302), .Z(n89318) );
  IV U108047 ( .A(n89304), .Z(n89306) );
  NOR U108048 ( .A(n89306), .B(n89305), .Z(n89316) );
  IV U108049 ( .A(n89307), .Z(n89309) );
  NOR U108050 ( .A(n89309), .B(n89308), .Z(n89313) );
  NOR U108051 ( .A(n89311), .B(n89310), .Z(n89312) );
  NOR U108052 ( .A(n89313), .B(n89312), .Z(n89314) );
  IV U108053 ( .A(n89314), .Z(n89315) );
  NOR U108054 ( .A(n89316), .B(n89315), .Z(n89317) );
  XOR U108055 ( .A(n89318), .B(n89317), .Z(n89342) );
  IV U108056 ( .A(n89319), .Z(n89321) );
  NOR U108057 ( .A(n89321), .B(n89320), .Z(n89326) );
  IV U108058 ( .A(n89322), .Z(n89323) );
  NOR U108059 ( .A(n89324), .B(n89323), .Z(n89325) );
  NOR U108060 ( .A(n89326), .B(n89325), .Z(n89331) );
  IV U108061 ( .A(n89327), .Z(n89328) );
  NOR U108062 ( .A(n89329), .B(n89328), .Z(n89330) );
  XOR U108063 ( .A(n89331), .B(n89330), .Z(n89340) );
  NOR U108064 ( .A(n89333), .B(n89332), .Z(n89335) );
  NOR U108065 ( .A(n89335), .B(n89334), .Z(n89336) );
  IV U108066 ( .A(n89336), .Z(n89337) );
  NOR U108067 ( .A(n89338), .B(n89337), .Z(n89339) );
  XOR U108068 ( .A(n89340), .B(n89339), .Z(n89341) );
  XOR U108069 ( .A(n89342), .B(n89341), .Z(n89343) );
  XOR U108070 ( .A(n89344), .B(n89343), .Z(n89354) );
  IV U108071 ( .A(n89347), .Z(n89345) );
  NOR U108072 ( .A(n89346), .B(n89345), .Z(n89352) );
  IV U108073 ( .A(n89346), .Z(n89348) );
  NOR U108074 ( .A(n89348), .B(n89347), .Z(n89349) );
  NOR U108075 ( .A(n89350), .B(n89349), .Z(n89351) );
  NOR U108076 ( .A(n89352), .B(n89351), .Z(n89353) );
  XOR U108077 ( .A(n89354), .B(n89353), .Z(n89355) );
  XOR U108078 ( .A(n89356), .B(n89355), .Z(n89357) );
  XOR U108079 ( .A(n89358), .B(n89357), .Z(n89359) );
  XOR U108080 ( .A(n89360), .B(n89359), .Z(n89361) );
  XOR U108081 ( .A(n89362), .B(n89361), .Z(n89363) );
  XOR U108082 ( .A(n89364), .B(n89363), .Z(n89365) );
  XOR U108083 ( .A(n89366), .B(n89365), .Z(n89367) );
  XOR U108084 ( .A(n89368), .B(n89367), .Z(n89386) );
  IV U108085 ( .A(n89369), .Z(n89371) );
  NOR U108086 ( .A(n89371), .B(n89370), .Z(n89375) );
  NOR U108087 ( .A(n89373), .B(n89372), .Z(n89374) );
  NOR U108088 ( .A(n89375), .B(n89374), .Z(n89384) );
  IV U108089 ( .A(n89376), .Z(n89378) );
  NOR U108090 ( .A(n89378), .B(n89377), .Z(n89382) );
  NOR U108091 ( .A(n89380), .B(n89379), .Z(n89381) );
  NOR U108092 ( .A(n89382), .B(n89381), .Z(n89383) );
  XOR U108093 ( .A(n89384), .B(n89383), .Z(n89385) );
  XOR U108094 ( .A(n89386), .B(n89385), .Z(n89387) );
  XOR U108095 ( .A(n89388), .B(n89387), .Z(n89389) );
  XOR U108096 ( .A(n89390), .B(n89389), .Z(n89409) );
  IV U108097 ( .A(n89391), .Z(n89393) );
  IV U108098 ( .A(n89392), .Z(n89429) );
  NOR U108099 ( .A(n89393), .B(n89429), .Z(n89397) );
  IV U108100 ( .A(n89394), .Z(n89395) );
  NOR U108101 ( .A(n89395), .B(n89425), .Z(n89396) );
  NOR U108102 ( .A(n89397), .B(n89396), .Z(n89407) );
  NOR U108103 ( .A(n89398), .B(n89399), .Z(n89405) );
  IV U108104 ( .A(n89399), .Z(n89400) );
  NOR U108105 ( .A(n89401), .B(n89400), .Z(n89402) );
  NOR U108106 ( .A(n89403), .B(n89402), .Z(n89404) );
  NOR U108107 ( .A(n89405), .B(n89404), .Z(n89406) );
  XOR U108108 ( .A(n89407), .B(n89406), .Z(n89408) );
  XOR U108109 ( .A(n89409), .B(n89408), .Z(n89410) );
  XOR U108110 ( .A(n89411), .B(n89410), .Z(n89439) );
  IV U108111 ( .A(n89412), .Z(n89413) );
  NOR U108112 ( .A(n89414), .B(n89413), .Z(n89419) );
  IV U108113 ( .A(n89415), .Z(n89416) );
  NOR U108114 ( .A(n89417), .B(n89416), .Z(n89418) );
  NOR U108115 ( .A(n89419), .B(n89418), .Z(n89420) );
  XOR U108116 ( .A(n89421), .B(n89420), .Z(n89437) );
  NOR U108117 ( .A(n89423), .B(n89422), .Z(n89430) );
  IV U108118 ( .A(n89424), .Z(n89426) );
  NOR U108119 ( .A(n89426), .B(n89425), .Z(n89427) );
  XOR U108120 ( .A(n89430), .B(n89427), .Z(n89435) );
  IV U108121 ( .A(n89428), .Z(n89433) );
  NOR U108122 ( .A(n89430), .B(n89429), .Z(n89431) );
  IV U108123 ( .A(n89431), .Z(n89432) );
  NOR U108124 ( .A(n89433), .B(n89432), .Z(n89434) );
  NOR U108125 ( .A(n89435), .B(n89434), .Z(n89436) );
  XOR U108126 ( .A(n89437), .B(n89436), .Z(n89438) );
  XOR U108127 ( .A(n89439), .B(n89438), .Z(n89440) );
  XOR U108128 ( .A(n89441), .B(n89440), .Z(n89442) );
  XOR U108129 ( .A(n89443), .B(n89442), .Z(n89444) );
  XOR U108130 ( .A(n89445), .B(n89444), .Z(n89446) );
  XOR U108131 ( .A(n89447), .B(n89446), .Z(n89448) );
  XOR U108132 ( .A(n89449), .B(n89448), .Z(n89450) );
  XOR U108133 ( .A(n89451), .B(n89450), .Z(n89466) );
  NOR U108134 ( .A(n89452), .B(n89453), .Z(n89464) );
  IV U108135 ( .A(n89452), .Z(n89455) );
  IV U108136 ( .A(n89453), .Z(n89454) );
  NOR U108137 ( .A(n89455), .B(n89454), .Z(n89462) );
  NOR U108138 ( .A(n89457), .B(n89456), .Z(n89458) );
  XOR U108139 ( .A(n89459), .B(n89458), .Z(n89460) );
  IV U108140 ( .A(n89460), .Z(n89461) );
  NOR U108141 ( .A(n89462), .B(n89461), .Z(n89463) );
  NOR U108142 ( .A(n89464), .B(n89463), .Z(n89465) );
  XOR U108143 ( .A(n89466), .B(n89465), .Z(n89467) );
  XOR U108144 ( .A(n89468), .B(n89467), .Z(n89486) );
  IV U108145 ( .A(n89469), .Z(n89470) );
  NOR U108146 ( .A(n89471), .B(n89470), .Z(n89475) );
  NOR U108147 ( .A(n89473), .B(n89472), .Z(n89474) );
  NOR U108148 ( .A(n89475), .B(n89474), .Z(n89484) );
  IV U108149 ( .A(n89476), .Z(n89477) );
  NOR U108150 ( .A(n89478), .B(n89477), .Z(n89482) );
  NOR U108151 ( .A(n89480), .B(n89479), .Z(n89481) );
  NOR U108152 ( .A(n89482), .B(n89481), .Z(n89483) );
  XOR U108153 ( .A(n89484), .B(n89483), .Z(n89485) );
  XOR U108154 ( .A(n89486), .B(n89485), .Z(n89487) );
  XOR U108155 ( .A(n89488), .B(n89487), .Z(n89517) );
  NOR U108156 ( .A(n89490), .B(n89489), .Z(n89506) );
  IV U108157 ( .A(n89491), .Z(n89497) );
  IV U108158 ( .A(n89492), .Z(n89494) );
  NOR U108159 ( .A(n89494), .B(n89493), .Z(n89495) );
  IV U108160 ( .A(n89495), .Z(n89496) );
  NOR U108161 ( .A(n89497), .B(n89496), .Z(n89504) );
  NOR U108162 ( .A(n89499), .B(n89498), .Z(n89501) );
  NOR U108163 ( .A(n89501), .B(n89500), .Z(n89502) );
  IV U108164 ( .A(n89502), .Z(n89503) );
  NOR U108165 ( .A(n89504), .B(n89503), .Z(n89505) );
  NOR U108166 ( .A(n89506), .B(n89505), .Z(n89515) );
  IV U108167 ( .A(n89507), .Z(n89509) );
  NOR U108168 ( .A(n89509), .B(n89508), .Z(n89513) );
  NOR U108169 ( .A(n89511), .B(n89510), .Z(n89512) );
  NOR U108170 ( .A(n89513), .B(n89512), .Z(n89514) );
  XOR U108171 ( .A(n89515), .B(n89514), .Z(n89516) );
  XOR U108172 ( .A(n89517), .B(n89516), .Z(n89518) );
  XOR U108173 ( .A(n89519), .B(n89518), .Z(n89520) );
  XOR U108174 ( .A(n89521), .B(n89520), .Z(n89522) );
  XOR U108175 ( .A(n89523), .B(n89522), .Z(n89524) );
  XOR U108176 ( .A(n89525), .B(n89524), .Z(n89531) );
  NOR U108177 ( .A(n89527), .B(n89526), .Z(n89529) );
  NOR U108178 ( .A(n89529), .B(n89528), .Z(n89530) );
  XOR U108179 ( .A(n89531), .B(n89530), .Z(n89532) );
  XOR U108180 ( .A(n89533), .B(n89532), .Z(n89534) );
  XOR U108181 ( .A(n89535), .B(n89534), .Z(n89550) );
  IV U108182 ( .A(n89536), .Z(n89537) );
  NOR U108183 ( .A(n89538), .B(n89537), .Z(n89543) );
  IV U108184 ( .A(n89539), .Z(n89541) );
  NOR U108185 ( .A(n89541), .B(n89540), .Z(n89542) );
  NOR U108186 ( .A(n89543), .B(n89542), .Z(n89548) );
  IV U108187 ( .A(n89544), .Z(n89546) );
  NOR U108188 ( .A(n89546), .B(n89545), .Z(n89547) );
  XOR U108189 ( .A(n89548), .B(n89547), .Z(n89549) );
  XOR U108190 ( .A(n89550), .B(n89549), .Z(n89551) );
  XOR U108191 ( .A(n89552), .B(n89551), .Z(n89581) );
  IV U108192 ( .A(n89553), .Z(n89554) );
  NOR U108193 ( .A(n89555), .B(n89554), .Z(n89559) );
  NOR U108194 ( .A(n89557), .B(n89556), .Z(n89558) );
  NOR U108195 ( .A(n89559), .B(n89558), .Z(n89569) );
  IV U108196 ( .A(n89560), .Z(n89562) );
  NOR U108197 ( .A(n89562), .B(n89561), .Z(n89567) );
  IV U108198 ( .A(n89563), .Z(n89565) );
  NOR U108199 ( .A(n89565), .B(n89564), .Z(n89566) );
  NOR U108200 ( .A(n89567), .B(n89566), .Z(n89568) );
  XOR U108201 ( .A(n89569), .B(n89568), .Z(n89579) );
  IV U108202 ( .A(n89573), .Z(n89571) );
  IV U108203 ( .A(n89572), .Z(n89570) );
  NOR U108204 ( .A(n89571), .B(n89570), .Z(n89577) );
  NOR U108205 ( .A(n89573), .B(n89572), .Z(n89575) );
  NOR U108206 ( .A(n89575), .B(n89574), .Z(n89576) );
  NOR U108207 ( .A(n89577), .B(n89576), .Z(n89578) );
  XOR U108208 ( .A(n89579), .B(n89578), .Z(n89580) );
  XOR U108209 ( .A(n89581), .B(n89580), .Z(n89582) );
  XOR U108210 ( .A(n89583), .B(n89582), .Z(n89584) );
  XOR U108211 ( .A(n89585), .B(n89584), .Z(n89586) );
  XOR U108212 ( .A(n89587), .B(n89586), .Z(n89588) );
  XOR U108213 ( .A(n89589), .B(n89588), .Z(n89590) );
  XOR U108214 ( .A(n89591), .B(n89590), .Z(n89600) );
  NOR U108215 ( .A(n89593), .B(n89592), .Z(n89595) );
  NOR U108216 ( .A(n89595), .B(n89594), .Z(n89596) );
  IV U108217 ( .A(n89596), .Z(n89597) );
  NOR U108218 ( .A(n89598), .B(n89597), .Z(n89599) );
  XOR U108219 ( .A(n89600), .B(n89599), .Z(n89615) );
  IV U108220 ( .A(n89601), .Z(n89604) );
  IV U108221 ( .A(n89602), .Z(n89603) );
  NOR U108222 ( .A(n89604), .B(n89603), .Z(n89609) );
  IV U108223 ( .A(n89605), .Z(n89607) );
  NOR U108224 ( .A(n89607), .B(n89606), .Z(n89608) );
  NOR U108225 ( .A(n89609), .B(n89608), .Z(n89613) );
  NOR U108226 ( .A(n89611), .B(n89610), .Z(n89612) );
  XOR U108227 ( .A(n89613), .B(n89612), .Z(n89614) );
  XOR U108228 ( .A(n89615), .B(n89614), .Z(n89627) );
  IV U108229 ( .A(n89616), .Z(n89618) );
  NOR U108230 ( .A(n89618), .B(n89617), .Z(n89620) );
  NOR U108231 ( .A(n89620), .B(n89619), .Z(n89625) );
  IV U108232 ( .A(n89621), .Z(n89623) );
  NOR U108233 ( .A(n89623), .B(n89622), .Z(n89624) );
  XOR U108234 ( .A(n89625), .B(n89624), .Z(n89626) );
  XOR U108235 ( .A(n89627), .B(n89626), .Z(n89628) );
  XOR U108236 ( .A(n89629), .B(n89628), .Z(n89630) );
  XOR U108237 ( .A(n89631), .B(n89630), .Z(n89666) );
  IV U108238 ( .A(n89632), .Z(n89633) );
  NOR U108239 ( .A(n89634), .B(n89633), .Z(n89645) );
  IV U108240 ( .A(n89635), .Z(n89637) );
  NOR U108241 ( .A(n89637), .B(n89636), .Z(n89642) );
  IV U108242 ( .A(n89638), .Z(n89640) );
  NOR U108243 ( .A(n89640), .B(n89639), .Z(n89641) );
  NOR U108244 ( .A(n89642), .B(n89641), .Z(n89643) );
  IV U108245 ( .A(n89643), .Z(n89644) );
  NOR U108246 ( .A(n89645), .B(n89644), .Z(n89664) );
  IV U108247 ( .A(n89646), .Z(n89648) );
  NOR U108248 ( .A(n89648), .B(n89647), .Z(n89652) );
  NOR U108249 ( .A(n89650), .B(n89649), .Z(n89651) );
  NOR U108250 ( .A(n89652), .B(n89651), .Z(n89662) );
  IV U108251 ( .A(n89653), .Z(n89654) );
  NOR U108252 ( .A(n89655), .B(n89654), .Z(n89660) );
  IV U108253 ( .A(n89656), .Z(n89658) );
  NOR U108254 ( .A(n89658), .B(n89657), .Z(n89659) );
  NOR U108255 ( .A(n89660), .B(n89659), .Z(n89661) );
  XOR U108256 ( .A(n89662), .B(n89661), .Z(n89663) );
  XOR U108257 ( .A(n89664), .B(n89663), .Z(n89665) );
  XOR U108258 ( .A(n89666), .B(n89665), .Z(n89686) );
  IV U108259 ( .A(n89667), .Z(n89668) );
  NOR U108260 ( .A(n89669), .B(n89668), .Z(n89674) );
  IV U108261 ( .A(n89670), .Z(n89672) );
  NOR U108262 ( .A(n89672), .B(n89671), .Z(n89673) );
  NOR U108263 ( .A(n89674), .B(n89673), .Z(n89684) );
  IV U108264 ( .A(n89675), .Z(n89677) );
  NOR U108265 ( .A(n89677), .B(n89676), .Z(n89682) );
  IV U108266 ( .A(n89678), .Z(n89680) );
  NOR U108267 ( .A(n89680), .B(n89679), .Z(n89681) );
  NOR U108268 ( .A(n89682), .B(n89681), .Z(n89683) );
  XOR U108269 ( .A(n89684), .B(n89683), .Z(n89685) );
  XOR U108270 ( .A(n89686), .B(n89685), .Z(n89687) );
  XOR U108271 ( .A(n89688), .B(n89687), .Z(n89712) );
  IV U108272 ( .A(n89689), .Z(n89691) );
  NOR U108273 ( .A(n89691), .B(n89690), .Z(n89710) );
  IV U108274 ( .A(n89692), .Z(n89693) );
  NOR U108275 ( .A(n89694), .B(n89693), .Z(n89698) );
  NOR U108276 ( .A(n89696), .B(n89695), .Z(n89697) );
  NOR U108277 ( .A(n89698), .B(n89697), .Z(n89708) );
  IV U108278 ( .A(n89699), .Z(n89700) );
  NOR U108279 ( .A(n89701), .B(n89700), .Z(n89706) );
  IV U108280 ( .A(n89702), .Z(n89704) );
  NOR U108281 ( .A(n89704), .B(n89703), .Z(n89705) );
  NOR U108282 ( .A(n89706), .B(n89705), .Z(n89707) );
  XOR U108283 ( .A(n89708), .B(n89707), .Z(n89709) );
  XOR U108284 ( .A(n89710), .B(n89709), .Z(n89711) );
  XOR U108285 ( .A(n89712), .B(n89711), .Z(n89730) );
  IV U108286 ( .A(n89713), .Z(n89715) );
  NOR U108287 ( .A(n89715), .B(n89714), .Z(n89718) );
  IV U108288 ( .A(n89741), .Z(n89716) );
  NOR U108289 ( .A(n89716), .B(n89740), .Z(n89717) );
  NOR U108290 ( .A(n89718), .B(n89717), .Z(n89728) );
  IV U108291 ( .A(n89719), .Z(n89721) );
  NOR U108292 ( .A(n89721), .B(n89720), .Z(n89726) );
  IV U108293 ( .A(n89722), .Z(n89724) );
  NOR U108294 ( .A(n89724), .B(n89723), .Z(n89725) );
  NOR U108295 ( .A(n89726), .B(n89725), .Z(n89727) );
  XOR U108296 ( .A(n89728), .B(n89727), .Z(n89729) );
  XOR U108297 ( .A(n89730), .B(n89729), .Z(n89731) );
  XOR U108298 ( .A(n89732), .B(n89731), .Z(n89748) );
  IV U108299 ( .A(n89733), .Z(n89734) );
  NOR U108300 ( .A(n89734), .B(n89740), .Z(n89739) );
  IV U108301 ( .A(n89735), .Z(n89737) );
  NOR U108302 ( .A(n89737), .B(n89736), .Z(n89738) );
  NOR U108303 ( .A(n89739), .B(n89738), .Z(n89746) );
  XOR U108304 ( .A(n89741), .B(n89740), .Z(n89744) );
  IV U108305 ( .A(n89742), .Z(n89743) );
  NOR U108306 ( .A(n89744), .B(n89743), .Z(n89745) );
  XOR U108307 ( .A(n89746), .B(n89745), .Z(n89747) );
  XOR U108308 ( .A(n89748), .B(n89747), .Z(n89749) );
  XOR U108309 ( .A(n89750), .B(n89749), .Z(n89751) );
  XOR U108310 ( .A(n89752), .B(n89751), .Z(n89771) );
  IV U108311 ( .A(n89753), .Z(n89754) );
  NOR U108312 ( .A(n89755), .B(n89754), .Z(n89760) );
  IV U108313 ( .A(n89756), .Z(n89757) );
  NOR U108314 ( .A(n89758), .B(n89757), .Z(n89759) );
  NOR U108315 ( .A(n89760), .B(n89759), .Z(n89769) );
  NOR U108316 ( .A(n89762), .B(n89761), .Z(n89767) );
  IV U108317 ( .A(n89763), .Z(n89764) );
  NOR U108318 ( .A(n89765), .B(n89764), .Z(n89766) );
  NOR U108319 ( .A(n89767), .B(n89766), .Z(n89768) );
  XOR U108320 ( .A(n89769), .B(n89768), .Z(n89770) );
  XOR U108321 ( .A(n89771), .B(n89770), .Z(n89772) );
  XOR U108322 ( .A(n89773), .B(n89772), .Z(n89774) );
  XOR U108323 ( .A(n89775), .B(n89774), .Z(n89776) );
  XOR U108324 ( .A(n89777), .B(n89776), .Z(n89778) );
  XOR U108325 ( .A(n89779), .B(n89778), .Z(n89780) );
  XOR U108326 ( .A(n89781), .B(n89780), .Z(n89782) );
  XOR U108327 ( .A(n89783), .B(n89782), .Z(n89784) );
  XOR U108328 ( .A(n89785), .B(n89784), .Z(n89786) );
  XOR U108329 ( .A(n89787), .B(n89786), .Z(n89788) );
  XOR U108330 ( .A(n89789), .B(n89788), .Z(n89801) );
  IV U108331 ( .A(n89790), .Z(n89791) );
  NOR U108332 ( .A(n89791), .B(n89793), .Z(n89799) );
  IV U108333 ( .A(n89792), .Z(n89794) );
  NOR U108334 ( .A(n89794), .B(n89793), .Z(n89796) );
  NOR U108335 ( .A(n89796), .B(n89795), .Z(n89797) );
  IV U108336 ( .A(n89797), .Z(n89798) );
  NOR U108337 ( .A(n89799), .B(n89798), .Z(n89800) );
  XOR U108338 ( .A(n89801), .B(n89800), .Z(n89821) );
  IV U108339 ( .A(n89802), .Z(n89804) );
  NOR U108340 ( .A(n89804), .B(n89803), .Z(n89809) );
  IV U108341 ( .A(n89805), .Z(n89807) );
  NOR U108342 ( .A(n89807), .B(n89806), .Z(n89808) );
  NOR U108343 ( .A(n89809), .B(n89808), .Z(n89819) );
  IV U108344 ( .A(n89810), .Z(n89812) );
  NOR U108345 ( .A(n89812), .B(n89811), .Z(n89817) );
  IV U108346 ( .A(n89813), .Z(n89815) );
  NOR U108347 ( .A(n89815), .B(n89814), .Z(n89816) );
  NOR U108348 ( .A(n89817), .B(n89816), .Z(n89818) );
  XOR U108349 ( .A(n89819), .B(n89818), .Z(n89820) );
  XOR U108350 ( .A(n89821), .B(n89820), .Z(n89844) );
  IV U108351 ( .A(n89822), .Z(n89824) );
  NOR U108352 ( .A(n89824), .B(n89823), .Z(n89826) );
  NOR U108353 ( .A(n89826), .B(n89825), .Z(n89842) );
  IV U108354 ( .A(n89827), .Z(n89830) );
  IV U108355 ( .A(n89828), .Z(n89829) );
  NOR U108356 ( .A(n89830), .B(n89829), .Z(n89840) );
  IV U108357 ( .A(n89831), .Z(n89832) );
  NOR U108358 ( .A(n89833), .B(n89832), .Z(n89837) );
  NOR U108359 ( .A(n89835), .B(n89834), .Z(n89836) );
  NOR U108360 ( .A(n89837), .B(n89836), .Z(n89838) );
  IV U108361 ( .A(n89838), .Z(n89839) );
  NOR U108362 ( .A(n89840), .B(n89839), .Z(n89841) );
  XOR U108363 ( .A(n89842), .B(n89841), .Z(n89843) );
  XOR U108364 ( .A(n89844), .B(n89843), .Z(n89863) );
  IV U108365 ( .A(n89845), .Z(n89846) );
  NOR U108366 ( .A(n89847), .B(n89846), .Z(n89851) );
  NOR U108367 ( .A(n89849), .B(n89848), .Z(n89850) );
  NOR U108368 ( .A(n89851), .B(n89850), .Z(n89861) );
  IV U108369 ( .A(n89852), .Z(n89854) );
  NOR U108370 ( .A(n89854), .B(n89853), .Z(n89859) );
  IV U108371 ( .A(n89855), .Z(n89857) );
  NOR U108372 ( .A(n89857), .B(n89856), .Z(n89858) );
  NOR U108373 ( .A(n89859), .B(n89858), .Z(n89860) );
  XOR U108374 ( .A(n89861), .B(n89860), .Z(n89862) );
  XOR U108375 ( .A(n89863), .B(n89862), .Z(n89864) );
  XOR U108376 ( .A(n89865), .B(n89864), .Z(n89875) );
  IV U108377 ( .A(n89866), .Z(n89867) );
  NOR U108378 ( .A(n89868), .B(n89867), .Z(n89873) );
  IV U108379 ( .A(n89869), .Z(n89871) );
  NOR U108380 ( .A(n89871), .B(n89870), .Z(n89872) );
  NOR U108381 ( .A(n89873), .B(n89872), .Z(n89874) );
  XOR U108382 ( .A(n89875), .B(n89874), .Z(n89888) );
  IV U108383 ( .A(n89876), .Z(n89878) );
  NOR U108384 ( .A(n89878), .B(n89877), .Z(n89886) );
  IV U108385 ( .A(n89879), .Z(n89881) );
  NOR U108386 ( .A(n89881), .B(n89880), .Z(n89882) );
  NOR U108387 ( .A(n89883), .B(n89882), .Z(n89884) );
  IV U108388 ( .A(n89884), .Z(n89885) );
  NOR U108389 ( .A(n89886), .B(n89885), .Z(n89887) );
  XOR U108390 ( .A(n89888), .B(n89887), .Z(n89893) );
  IV U108391 ( .A(n89889), .Z(n89890) );
  NOR U108392 ( .A(n89891), .B(n89890), .Z(n89892) );
  XOR U108393 ( .A(n89893), .B(n89892), .Z(n89900) );
  IV U108394 ( .A(n89894), .Z(n89896) );
  NOR U108395 ( .A(n89896), .B(n89895), .Z(n89898) );
  NOR U108396 ( .A(n89898), .B(n89897), .Z(n89899) );
  XOR U108397 ( .A(n89900), .B(n89899), .Z(n89910) );
  NOR U108398 ( .A(n89902), .B(n89901), .Z(n89908) );
  IV U108399 ( .A(n89903), .Z(n89906) );
  IV U108400 ( .A(n89904), .Z(n89905) );
  NOR U108401 ( .A(n89906), .B(n89905), .Z(n89907) );
  NOR U108402 ( .A(n89908), .B(n89907), .Z(n89909) );
  XOR U108403 ( .A(n89910), .B(n89909), .Z(n89916) );
  NOR U108404 ( .A(n89912), .B(n89911), .Z(n89913) );
  NOR U108405 ( .A(n89914), .B(n89913), .Z(n89915) );
  XOR U108406 ( .A(n89916), .B(n89915), .Z(n89917) );
  XOR U108407 ( .A(n89918), .B(n89917), .Z(n89919) );
  XOR U108408 ( .A(n89920), .B(n89919), .Z(n89921) );
  XOR U108409 ( .A(n89922), .B(n89921), .Z(n89923) );
  XOR U108410 ( .A(n89924), .B(n89923), .Z(n89948) );
  IV U108411 ( .A(n89925), .Z(n89926) );
  NOR U108412 ( .A(n89927), .B(n89926), .Z(n89931) );
  NOR U108413 ( .A(n89929), .B(n89928), .Z(n89930) );
  NOR U108414 ( .A(n89931), .B(n89930), .Z(n89946) );
  XOR U108415 ( .A(n89934), .B(n89935), .Z(n89933) );
  NOR U108416 ( .A(n89933), .B(n89932), .Z(n89938) );
  IV U108417 ( .A(n89934), .Z(n89936) );
  NOR U108418 ( .A(n89936), .B(n89935), .Z(n89937) );
  NOR U108419 ( .A(n89938), .B(n89937), .Z(n89939) );
  IV U108420 ( .A(n89939), .Z(n89944) );
  IV U108421 ( .A(n89940), .Z(n89942) );
  NOR U108422 ( .A(n89942), .B(n89941), .Z(n89943) );
  NOR U108423 ( .A(n89944), .B(n89943), .Z(n89945) );
  XOR U108424 ( .A(n89946), .B(n89945), .Z(n89947) );
  XOR U108425 ( .A(n89948), .B(n89947), .Z(n89949) );
  XOR U108426 ( .A(n89950), .B(n89949), .Z(n89951) );
  XOR U108427 ( .A(n89952), .B(n89951), .Z(n89953) );
  XOR U108428 ( .A(n89954), .B(n89953), .Z(n89959) );
  IV U108429 ( .A(n89955), .Z(n89956) );
  NOR U108430 ( .A(n89957), .B(n89956), .Z(n89958) );
  XOR U108431 ( .A(n89959), .B(n89958), .Z(n89968) );
  NOR U108432 ( .A(n89960), .B(n89961), .Z(n89966) );
  IV U108433 ( .A(n89961), .Z(n89962) );
  NOR U108434 ( .A(n89963), .B(n89962), .Z(n89964) );
  NOR U108435 ( .A(n89990), .B(n89964), .Z(n89965) );
  NOR U108436 ( .A(n89966), .B(n89965), .Z(n89967) );
  XOR U108437 ( .A(n89968), .B(n89967), .Z(n89978) );
  NOR U108438 ( .A(n89970), .B(n89969), .Z(n89976) );
  IV U108439 ( .A(n89971), .Z(n89974) );
  IV U108440 ( .A(n89972), .Z(n89973) );
  NOR U108441 ( .A(n89974), .B(n89973), .Z(n89975) );
  NOR U108442 ( .A(n89976), .B(n89975), .Z(n89977) );
  XOR U108443 ( .A(n89978), .B(n89977), .Z(n89995) );
  IV U108444 ( .A(n89979), .Z(n89980) );
  NOR U108445 ( .A(n89981), .B(n89980), .Z(n89986) );
  IV U108446 ( .A(n89982), .Z(n89984) );
  NOR U108447 ( .A(n89984), .B(n89983), .Z(n89985) );
  NOR U108448 ( .A(n89986), .B(n89985), .Z(n89993) );
  NOR U108449 ( .A(n89988), .B(n89987), .Z(n89989) );
  IV U108450 ( .A(n89989), .Z(n89991) );
  NOR U108451 ( .A(n89991), .B(n89990), .Z(n89992) );
  XOR U108452 ( .A(n89993), .B(n89992), .Z(n89994) );
  XOR U108453 ( .A(n89995), .B(n89994), .Z(n89996) );
  XOR U108454 ( .A(n89997), .B(n89996), .Z(n90008) );
  NOR U108455 ( .A(n89998), .B(n90000), .Z(n90006) );
  IV U108456 ( .A(n89999), .Z(n90004) );
  IV U108457 ( .A(n90000), .Z(n90002) );
  NOR U108458 ( .A(n90002), .B(n90001), .Z(n90003) );
  NOR U108459 ( .A(n90004), .B(n90003), .Z(n90005) );
  NOR U108460 ( .A(n90006), .B(n90005), .Z(n90007) );
  XOR U108461 ( .A(n90008), .B(n90007), .Z(n90018) );
  IV U108462 ( .A(n90009), .Z(n90011) );
  NOR U108463 ( .A(n90011), .B(n90010), .Z(n90016) );
  IV U108464 ( .A(n90012), .Z(n90013) );
  NOR U108465 ( .A(n90014), .B(n90013), .Z(n90015) );
  NOR U108466 ( .A(n90016), .B(n90015), .Z(n90017) );
  XOR U108467 ( .A(n90018), .B(n90017), .Z(n90034) );
  IV U108468 ( .A(n90019), .Z(n90020) );
  NOR U108469 ( .A(n90027), .B(n90020), .Z(n90021) );
  NOR U108470 ( .A(n90022), .B(n90021), .Z(n90032) );
  IV U108471 ( .A(n90023), .Z(n90025) );
  NOR U108472 ( .A(n90025), .B(n90024), .Z(n90030) );
  IV U108473 ( .A(n90026), .Z(n90028) );
  NOR U108474 ( .A(n90028), .B(n90027), .Z(n90029) );
  NOR U108475 ( .A(n90030), .B(n90029), .Z(n90031) );
  XOR U108476 ( .A(n90032), .B(n90031), .Z(n90033) );
  XOR U108477 ( .A(n90034), .B(n90033), .Z(n90035) );
  XOR U108478 ( .A(n90036), .B(n90035), .Z(n90051) );
  IV U108479 ( .A(n90037), .Z(n90039) );
  NOR U108480 ( .A(n90039), .B(n90038), .Z(n90044) );
  IV U108481 ( .A(n90040), .Z(n90042) );
  NOR U108482 ( .A(n90042), .B(n90041), .Z(n90043) );
  NOR U108483 ( .A(n90044), .B(n90043), .Z(n90049) );
  IV U108484 ( .A(n90045), .Z(n90046) );
  NOR U108485 ( .A(n90047), .B(n90046), .Z(n90048) );
  XOR U108486 ( .A(n90049), .B(n90048), .Z(n90050) );
  XOR U108487 ( .A(n90051), .B(n90050), .Z(n90052) );
  XOR U108488 ( .A(n90053), .B(n90052), .Z(n90054) );
  XOR U108489 ( .A(n90055), .B(n90054), .Z(n90056) );
  XOR U108490 ( .A(n90057), .B(n90056), .Z(n90066) );
  NOR U108491 ( .A(n90059), .B(n90058), .Z(n90064) );
  IV U108492 ( .A(n90060), .Z(n90062) );
  NOR U108493 ( .A(n90062), .B(n90061), .Z(n90063) );
  NOR U108494 ( .A(n90064), .B(n90063), .Z(n90065) );
  XOR U108495 ( .A(n90066), .B(n90065), .Z(n90086) );
  IV U108496 ( .A(n90067), .Z(n90069) );
  NOR U108497 ( .A(n90069), .B(n90068), .Z(n90074) );
  IV U108498 ( .A(n90070), .Z(n90072) );
  NOR U108499 ( .A(n90072), .B(n90071), .Z(n90073) );
  NOR U108500 ( .A(n90074), .B(n90073), .Z(n90084) );
  IV U108501 ( .A(n90075), .Z(n90077) );
  NOR U108502 ( .A(n90077), .B(n90076), .Z(n90082) );
  IV U108503 ( .A(n90078), .Z(n90080) );
  NOR U108504 ( .A(n90080), .B(n90079), .Z(n90081) );
  NOR U108505 ( .A(n90082), .B(n90081), .Z(n90083) );
  XOR U108506 ( .A(n90084), .B(n90083), .Z(n90085) );
  XOR U108507 ( .A(n90086), .B(n90085), .Z(n90087) );
  XOR U108508 ( .A(n90088), .B(n90087), .Z(n90089) );
  XOR U108509 ( .A(n90090), .B(n90089), .Z(n90091) );
  XOR U108510 ( .A(n90092), .B(n90091), .Z(n90102) );
  IV U108511 ( .A(n90095), .Z(n90093) );
  NOR U108512 ( .A(n90094), .B(n90093), .Z(n90100) );
  NOR U108513 ( .A(n90096), .B(n90095), .Z(n90098) );
  NOR U108514 ( .A(n90098), .B(n90097), .Z(n90099) );
  NOR U108515 ( .A(n90100), .B(n90099), .Z(n90101) );
  XOR U108516 ( .A(n90102), .B(n90101), .Z(n90103) );
  XOR U108517 ( .A(n90104), .B(n90103), .Z(n90105) );
  XOR U108518 ( .A(n90106), .B(n90105), .Z(n90140) );
  IV U108519 ( .A(n90107), .Z(n90109) );
  NOR U108520 ( .A(n90109), .B(n90108), .Z(n90114) );
  IV U108521 ( .A(n90110), .Z(n90111) );
  NOR U108522 ( .A(n90112), .B(n90111), .Z(n90113) );
  NOR U108523 ( .A(n90114), .B(n90113), .Z(n90124) );
  IV U108524 ( .A(n90115), .Z(n90117) );
  NOR U108525 ( .A(n90117), .B(n90116), .Z(n90122) );
  IV U108526 ( .A(n90118), .Z(n90120) );
  NOR U108527 ( .A(n90120), .B(n90119), .Z(n90121) );
  NOR U108528 ( .A(n90122), .B(n90121), .Z(n90123) );
  XOR U108529 ( .A(n90124), .B(n90123), .Z(n90138) );
  NOR U108530 ( .A(n90126), .B(n90125), .Z(n90131) );
  IV U108531 ( .A(n90127), .Z(n90129) );
  NOR U108532 ( .A(n90129), .B(n90128), .Z(n90130) );
  NOR U108533 ( .A(n90131), .B(n90130), .Z(n90136) );
  IV U108534 ( .A(n90132), .Z(n90133) );
  NOR U108535 ( .A(n90134), .B(n90133), .Z(n90135) );
  XOR U108536 ( .A(n90136), .B(n90135), .Z(n90137) );
  XOR U108537 ( .A(n90138), .B(n90137), .Z(n90139) );
  XOR U108538 ( .A(n90140), .B(n90139), .Z(n90146) );
  NOR U108539 ( .A(n90142), .B(n90141), .Z(n90144) );
  NOR U108540 ( .A(n90144), .B(n90143), .Z(n90145) );
  XOR U108541 ( .A(n90146), .B(n90145), .Z(n90165) );
  IV U108542 ( .A(n90147), .Z(n90148) );
  NOR U108543 ( .A(n90149), .B(n90148), .Z(n90153) );
  NOR U108544 ( .A(n90151), .B(n90150), .Z(n90152) );
  NOR U108545 ( .A(n90153), .B(n90152), .Z(n90163) );
  IV U108546 ( .A(n90154), .Z(n90155) );
  NOR U108547 ( .A(n90156), .B(n90155), .Z(n90161) );
  IV U108548 ( .A(n90157), .Z(n90158) );
  NOR U108549 ( .A(n90159), .B(n90158), .Z(n90160) );
  NOR U108550 ( .A(n90161), .B(n90160), .Z(n90162) );
  XOR U108551 ( .A(n90163), .B(n90162), .Z(n90164) );
  XOR U108552 ( .A(n90165), .B(n90164), .Z(n90166) );
  XOR U108553 ( .A(n90167), .B(n90166), .Z(n90168) );
  XOR U108554 ( .A(n90169), .B(n90168), .Z(n90170) );
  XOR U108555 ( .A(n90171), .B(n90170), .Z(n90172) );
  XOR U108556 ( .A(n90173), .B(n90172), .Z(n90174) );
  XOR U108557 ( .A(n90175), .B(n90174), .Z(n90207) );
  IV U108558 ( .A(n90176), .Z(n90177) );
  NOR U108559 ( .A(n90178), .B(n90177), .Z(n90183) );
  IV U108560 ( .A(n90179), .Z(n90180) );
  NOR U108561 ( .A(n90181), .B(n90180), .Z(n90182) );
  NOR U108562 ( .A(n90183), .B(n90182), .Z(n90194) );
  IV U108563 ( .A(n90188), .Z(n90184) );
  NOR U108564 ( .A(n90185), .B(n90184), .Z(n90192) );
  IV U108565 ( .A(n90186), .Z(n90190) );
  NOR U108566 ( .A(n90188), .B(n90187), .Z(n90189) );
  NOR U108567 ( .A(n90190), .B(n90189), .Z(n90191) );
  NOR U108568 ( .A(n90192), .B(n90191), .Z(n90193) );
  XOR U108569 ( .A(n90194), .B(n90193), .Z(n90205) );
  IV U108570 ( .A(n90195), .Z(n90197) );
  NOR U108571 ( .A(n90197), .B(n90196), .Z(n90203) );
  NOR U108572 ( .A(n90199), .B(n90198), .Z(n90200) );
  NOR U108573 ( .A(n90201), .B(n90200), .Z(n90202) );
  XOR U108574 ( .A(n90203), .B(n90202), .Z(n90204) );
  XOR U108575 ( .A(n90205), .B(n90204), .Z(n90206) );
  XOR U108576 ( .A(n90207), .B(n90206), .Z(n90222) );
  IV U108577 ( .A(n90208), .Z(n90210) );
  NOR U108578 ( .A(n90210), .B(n90209), .Z(n90220) );
  IV U108579 ( .A(n90211), .Z(n90213) );
  NOR U108580 ( .A(n90213), .B(n90212), .Z(n90218) );
  IV U108581 ( .A(n90214), .Z(n90215) );
  NOR U108582 ( .A(n90216), .B(n90215), .Z(n90217) );
  NOR U108583 ( .A(n90218), .B(n90217), .Z(n90219) );
  XOR U108584 ( .A(n90220), .B(n90219), .Z(n90221) );
  XOR U108585 ( .A(n90222), .B(n90221), .Z(n90223) );
  XOR U108586 ( .A(n90224), .B(n90223), .Z(n90225) );
  XOR U108587 ( .A(n90226), .B(n90225), .Z(n90227) );
  XOR U108588 ( .A(n90228), .B(n90227), .Z(n90229) );
  XOR U108589 ( .A(n90230), .B(n90229), .Z(n90231) );
  XOR U108590 ( .A(n90232), .B(n90231), .Z(n90233) );
  XOR U108591 ( .A(n90234), .B(n90233), .Z(n90235) );
  XOR U108592 ( .A(n90236), .B(n90235), .Z(n90237) );
  XOR U108593 ( .A(n90238), .B(n90237), .Z(n90239) );
  XOR U108594 ( .A(n90240), .B(n90239), .Z(n90249) );
  IV U108595 ( .A(n90241), .Z(n90242) );
  NOR U108596 ( .A(n90243), .B(n90242), .Z(n90247) );
  NOR U108597 ( .A(n90245), .B(n90244), .Z(n90246) );
  NOR U108598 ( .A(n90247), .B(n90246), .Z(n90248) );
  XOR U108599 ( .A(n90249), .B(n90248), .Z(n90250) );
  XOR U108600 ( .A(n90251), .B(n90250), .Z(n90252) );
  XOR U108601 ( .A(n90253), .B(n90252), .Z(n90274) );
  IV U108602 ( .A(n90254), .Z(n90255) );
  NOR U108603 ( .A(n90256), .B(n90255), .Z(n90257) );
  IV U108604 ( .A(n90257), .Z(n90259) );
  NOR U108605 ( .A(n90259), .B(n90258), .Z(n90262) );
  NOR U108606 ( .A(n90260), .B(n90267), .Z(n90261) );
  NOR U108607 ( .A(n90262), .B(n90261), .Z(n90272) );
  IV U108608 ( .A(n90263), .Z(n90277) );
  IV U108609 ( .A(n90264), .Z(n90265) );
  NOR U108610 ( .A(n90277), .B(n90265), .Z(n90270) );
  IV U108611 ( .A(n90266), .Z(n90268) );
  NOR U108612 ( .A(n90268), .B(n90267), .Z(n90269) );
  NOR U108613 ( .A(n90270), .B(n90269), .Z(n90271) );
  XOR U108614 ( .A(n90272), .B(n90271), .Z(n90273) );
  XOR U108615 ( .A(n90274), .B(n90273), .Z(n90302) );
  IV U108616 ( .A(n90275), .Z(n90276) );
  NOR U108617 ( .A(n90277), .B(n90276), .Z(n90300) );
  IV U108618 ( .A(n90278), .Z(n90282) );
  IV U108619 ( .A(n90286), .Z(n90279) );
  NOR U108620 ( .A(n90280), .B(n90279), .Z(n90281) );
  NOR U108621 ( .A(n90282), .B(n90281), .Z(n90291) );
  NOR U108622 ( .A(n90284), .B(n90283), .Z(n90288) );
  NOR U108623 ( .A(n90286), .B(n90285), .Z(n90287) );
  NOR U108624 ( .A(n90288), .B(n90287), .Z(n90289) );
  IV U108625 ( .A(n90289), .Z(n90290) );
  NOR U108626 ( .A(n90291), .B(n90290), .Z(n90298) );
  IV U108627 ( .A(n90292), .Z(n90294) );
  NOR U108628 ( .A(n90294), .B(n90293), .Z(n90295) );
  NOR U108629 ( .A(n90296), .B(n90295), .Z(n90297) );
  XOR U108630 ( .A(n90298), .B(n90297), .Z(n90299) );
  XOR U108631 ( .A(n90300), .B(n90299), .Z(n90301) );
  XOR U108632 ( .A(n90302), .B(n90301), .Z(n90303) );
  XOR U108633 ( .A(n90304), .B(n90303), .Z(n90305) );
  XOR U108634 ( .A(n90306), .B(n90305), .Z(n90307) );
  XOR U108635 ( .A(n90308), .B(n90307), .Z(n90309) );
  XOR U108636 ( .A(n90310), .B(n90309), .Z(n90321) );
  NOR U108637 ( .A(n90313), .B(n90311), .Z(n90319) );
  IV U108638 ( .A(n90312), .Z(n90317) );
  IV U108639 ( .A(n90313), .Z(n90314) );
  NOR U108640 ( .A(n90315), .B(n90314), .Z(n90316) );
  NOR U108641 ( .A(n90317), .B(n90316), .Z(n90318) );
  NOR U108642 ( .A(n90319), .B(n90318), .Z(n90320) );
  XOR U108643 ( .A(n90321), .B(n90320), .Z(n90337) );
  IV U108644 ( .A(n90322), .Z(n90323) );
  NOR U108645 ( .A(n90324), .B(n90323), .Z(n90328) );
  NOR U108646 ( .A(n90326), .B(n90325), .Z(n90327) );
  NOR U108647 ( .A(n90328), .B(n90327), .Z(n90335) );
  IV U108648 ( .A(n90329), .Z(n90331) );
  NOR U108649 ( .A(n90331), .B(n90330), .Z(n90332) );
  NOR U108650 ( .A(n90333), .B(n90332), .Z(n90334) );
  XOR U108651 ( .A(n90335), .B(n90334), .Z(n90336) );
  XOR U108652 ( .A(n90337), .B(n90336), .Z(n90338) );
  XOR U108653 ( .A(n90339), .B(n90338), .Z(n90340) );
  XOR U108654 ( .A(n90341), .B(n90340), .Z(n90342) );
  XOR U108655 ( .A(n90343), .B(n90342), .Z(n90344) );
  XOR U108656 ( .A(n90345), .B(n90344), .Z(n90346) );
  XOR U108657 ( .A(n90347), .B(n90346), .Z(n90348) );
  XOR U108658 ( .A(n90349), .B(n90348), .Z(n90350) );
  XOR U108659 ( .A(n90351), .B(n90350), .Z(n90352) );
  XOR U108660 ( .A(n90353), .B(n90352), .Z(n90354) );
  XOR U108661 ( .A(n90355), .B(n90354), .Z(n90384) );
  NOR U108662 ( .A(n90357), .B(n90356), .Z(n90364) );
  NOR U108663 ( .A(n90359), .B(n90358), .Z(n90362) );
  IV U108664 ( .A(n90360), .Z(n90361) );
  NOR U108665 ( .A(n90362), .B(n90361), .Z(n90363) );
  NOR U108666 ( .A(n90364), .B(n90363), .Z(n90382) );
  NOR U108667 ( .A(n90365), .B(n90366), .Z(n90375) );
  IV U108668 ( .A(n90365), .Z(n90368) );
  IV U108669 ( .A(n90366), .Z(n90367) );
  NOR U108670 ( .A(n90368), .B(n90367), .Z(n90369) );
  NOR U108671 ( .A(n90370), .B(n90369), .Z(n90371) );
  IV U108672 ( .A(n90371), .Z(n90372) );
  NOR U108673 ( .A(n90373), .B(n90372), .Z(n90374) );
  NOR U108674 ( .A(n90375), .B(n90374), .Z(n90380) );
  IV U108675 ( .A(n90376), .Z(n90378) );
  NOR U108676 ( .A(n90378), .B(n90377), .Z(n90379) );
  NOR U108677 ( .A(n90380), .B(n90379), .Z(n90381) );
  XOR U108678 ( .A(n90382), .B(n90381), .Z(n90383) );
  XOR U108679 ( .A(n90384), .B(n90383), .Z(n90385) );
  XOR U108680 ( .A(n90386), .B(n90385), .Z(n90409) );
  IV U108681 ( .A(n90387), .Z(n90389) );
  NOR U108682 ( .A(n90389), .B(n90388), .Z(n90397) );
  IV U108683 ( .A(n90390), .Z(n90432) );
  IV U108684 ( .A(n90391), .Z(n90392) );
  NOR U108685 ( .A(n90393), .B(n90392), .Z(n90394) );
  IV U108686 ( .A(n90394), .Z(n90395) );
  NOR U108687 ( .A(n90432), .B(n90395), .Z(n90396) );
  NOR U108688 ( .A(n90397), .B(n90396), .Z(n90407) );
  NOR U108689 ( .A(n90399), .B(n90398), .Z(n90405) );
  IV U108690 ( .A(n90400), .Z(n90403) );
  IV U108691 ( .A(n90401), .Z(n90402) );
  NOR U108692 ( .A(n90403), .B(n90402), .Z(n90404) );
  NOR U108693 ( .A(n90405), .B(n90404), .Z(n90406) );
  XOR U108694 ( .A(n90407), .B(n90406), .Z(n90408) );
  XOR U108695 ( .A(n90409), .B(n90408), .Z(n90410) );
  XOR U108696 ( .A(n90411), .B(n90410), .Z(n90422) );
  IV U108697 ( .A(n90416), .Z(n90413) );
  NOR U108698 ( .A(n90413), .B(n90412), .Z(n90420) );
  IV U108699 ( .A(n90414), .Z(n90418) );
  NOR U108700 ( .A(n90416), .B(n90415), .Z(n90417) );
  NOR U108701 ( .A(n90418), .B(n90417), .Z(n90419) );
  NOR U108702 ( .A(n90420), .B(n90419), .Z(n90421) );
  XOR U108703 ( .A(n90422), .B(n90421), .Z(n90434) );
  NOR U108704 ( .A(n90424), .B(n90423), .Z(n90425) );
  IV U108705 ( .A(n90425), .Z(n90426) );
  NOR U108706 ( .A(n90427), .B(n90426), .Z(n90428) );
  XOR U108707 ( .A(n90429), .B(n90428), .Z(n90430) );
  IV U108708 ( .A(n90430), .Z(n90431) );
  NOR U108709 ( .A(n90432), .B(n90431), .Z(n90433) );
  XOR U108710 ( .A(n90434), .B(n90433), .Z(n90435) );
  XOR U108711 ( .A(n90436), .B(n90435), .Z(n90471) );
  IV U108712 ( .A(n90440), .Z(n90437) );
  NOR U108713 ( .A(n90437), .B(n90438), .Z(n90444) );
  IV U108714 ( .A(n90438), .Z(n90439) );
  NOR U108715 ( .A(n90440), .B(n90439), .Z(n90441) );
  NOR U108716 ( .A(n90442), .B(n90441), .Z(n90443) );
  NOR U108717 ( .A(n90444), .B(n90443), .Z(n90460) );
  IV U108718 ( .A(n90445), .Z(n90447) );
  NOR U108719 ( .A(n90447), .B(n90446), .Z(n90458) );
  IV U108720 ( .A(n90448), .Z(n90450) );
  NOR U108721 ( .A(n90450), .B(n90449), .Z(n90455) );
  IV U108722 ( .A(n90451), .Z(n90453) );
  NOR U108723 ( .A(n90453), .B(n90452), .Z(n90454) );
  NOR U108724 ( .A(n90455), .B(n90454), .Z(n90456) );
  IV U108725 ( .A(n90456), .Z(n90457) );
  NOR U108726 ( .A(n90458), .B(n90457), .Z(n90459) );
  XOR U108727 ( .A(n90460), .B(n90459), .Z(n90469) );
  IV U108728 ( .A(n90461), .Z(n90463) );
  NOR U108729 ( .A(n90463), .B(n90462), .Z(n90467) );
  NOR U108730 ( .A(n90465), .B(n90464), .Z(n90466) );
  NOR U108731 ( .A(n90467), .B(n90466), .Z(n90468) );
  XOR U108732 ( .A(n90469), .B(n90468), .Z(n90470) );
  XOR U108733 ( .A(n90471), .B(n90470), .Z(n90472) );
  XOR U108734 ( .A(n90473), .B(n90472), .Z(n90474) );
  XOR U108735 ( .A(n90475), .B(n90474), .Z(n90476) );
  XOR U108736 ( .A(n90477), .B(n90476), .Z(n90491) );
  NOR U108737 ( .A(n90479), .B(n90478), .Z(n90489) );
  XOR U108738 ( .A(n90482), .B(n90483), .Z(n90481) );
  NOR U108739 ( .A(n90481), .B(n90480), .Z(n90486) );
  IV U108740 ( .A(n90482), .Z(n90484) );
  NOR U108741 ( .A(n90484), .B(n90483), .Z(n90485) );
  NOR U108742 ( .A(n90486), .B(n90485), .Z(n90487) );
  IV U108743 ( .A(n90487), .Z(n90488) );
  NOR U108744 ( .A(n90489), .B(n90488), .Z(n90490) );
  XOR U108745 ( .A(n90491), .B(n90490), .Z(n90492) );
  XOR U108746 ( .A(n90493), .B(n90492), .Z(n90494) );
  XOR U108747 ( .A(n90495), .B(n90494), .Z(n90496) );
  XOR U108748 ( .A(n90497), .B(n90496), .Z(n90498) );
  XOR U108749 ( .A(n90499), .B(n90498), .Z(n90500) );
  XOR U108750 ( .A(n90501), .B(n90500), .Z(n90502) );
  XOR U108751 ( .A(n90503), .B(n90502), .Z(n90504) );
  XOR U108752 ( .A(n90505), .B(n90504), .Z(n90522) );
  IV U108753 ( .A(n90506), .Z(n90507) );
  NOR U108754 ( .A(n90508), .B(n90507), .Z(n90514) );
  IV U108755 ( .A(n90509), .Z(n90512) );
  IV U108756 ( .A(n90510), .Z(n90511) );
  NOR U108757 ( .A(n90512), .B(n90511), .Z(n90513) );
  NOR U108758 ( .A(n90514), .B(n90513), .Z(n90520) );
  IV U108759 ( .A(n90515), .Z(n90518) );
  IV U108760 ( .A(n90516), .Z(n90517) );
  NOR U108761 ( .A(n90518), .B(n90517), .Z(n90519) );
  XOR U108762 ( .A(n90520), .B(n90519), .Z(n90521) );
  XOR U108763 ( .A(n90522), .B(n90521), .Z(n90523) );
  XOR U108764 ( .A(n90524), .B(n90523), .Z(n90546) );
  IV U108765 ( .A(n90528), .Z(n90525) );
  NOR U108766 ( .A(n90526), .B(n90525), .Z(n90533) );
  IV U108767 ( .A(n90526), .Z(n90527) );
  NOR U108768 ( .A(n90528), .B(n90527), .Z(n90531) );
  IV U108769 ( .A(n90529), .Z(n90530) );
  NOR U108770 ( .A(n90531), .B(n90530), .Z(n90532) );
  NOR U108771 ( .A(n90533), .B(n90532), .Z(n90544) );
  IV U108772 ( .A(n90534), .Z(n90537) );
  IV U108773 ( .A(n90535), .Z(n90536) );
  NOR U108774 ( .A(n90537), .B(n90536), .Z(n90542) );
  IV U108775 ( .A(n90538), .Z(n90539) );
  NOR U108776 ( .A(n90540), .B(n90539), .Z(n90541) );
  NOR U108777 ( .A(n90542), .B(n90541), .Z(n90543) );
  XOR U108778 ( .A(n90544), .B(n90543), .Z(n90545) );
  XOR U108779 ( .A(n90546), .B(n90545), .Z(n90547) );
  XOR U108780 ( .A(n90548), .B(n90547), .Z(n90560) );
  IV U108781 ( .A(n90549), .Z(n90550) );
  NOR U108782 ( .A(n90551), .B(n90550), .Z(n90556) );
  IV U108783 ( .A(n90552), .Z(n90554) );
  NOR U108784 ( .A(n90554), .B(n90553), .Z(n90555) );
  NOR U108785 ( .A(n90556), .B(n90555), .Z(n90557) );
  XOR U108786 ( .A(n90558), .B(n90557), .Z(n90559) );
  XOR U108787 ( .A(n90560), .B(n90559), .Z(n90561) );
  XOR U108788 ( .A(n90562), .B(n90561), .Z(n90585) );
  IV U108789 ( .A(n90565), .Z(n90563) );
  NOR U108790 ( .A(n90564), .B(n90563), .Z(n90573) );
  NOR U108791 ( .A(n90566), .B(n90565), .Z(n90571) );
  XOR U108792 ( .A(n90568), .B(n90567), .Z(n90569) );
  IV U108793 ( .A(n90569), .Z(n90570) );
  NOR U108794 ( .A(n90571), .B(n90570), .Z(n90572) );
  NOR U108795 ( .A(n90573), .B(n90572), .Z(n90583) );
  IV U108796 ( .A(n90574), .Z(n90575) );
  NOR U108797 ( .A(n90576), .B(n90575), .Z(n90581) );
  IV U108798 ( .A(n90577), .Z(n90579) );
  NOR U108799 ( .A(n90579), .B(n90578), .Z(n90580) );
  NOR U108800 ( .A(n90581), .B(n90580), .Z(n90582) );
  XOR U108801 ( .A(n90583), .B(n90582), .Z(n90584) );
  XOR U108802 ( .A(n90585), .B(n90584), .Z(n90586) );
  XOR U108803 ( .A(n90587), .B(n90586), .Z(n90614) );
  IV U108804 ( .A(n90588), .Z(n90590) );
  NOR U108805 ( .A(n90590), .B(n90589), .Z(n90594) );
  NOR U108806 ( .A(n90592), .B(n90591), .Z(n90593) );
  NOR U108807 ( .A(n90594), .B(n90593), .Z(n90603) );
  IV U108808 ( .A(n90595), .Z(n90597) );
  NOR U108809 ( .A(n90597), .B(n90596), .Z(n90601) );
  NOR U108810 ( .A(n90599), .B(n90598), .Z(n90600) );
  NOR U108811 ( .A(n90601), .B(n90600), .Z(n90602) );
  XOR U108812 ( .A(n90603), .B(n90602), .Z(n90612) );
  NOR U108813 ( .A(n90605), .B(n90604), .Z(n90610) );
  IV U108814 ( .A(n90606), .Z(n90607) );
  NOR U108815 ( .A(n90608), .B(n90607), .Z(n90609) );
  NOR U108816 ( .A(n90610), .B(n90609), .Z(n90611) );
  XOR U108817 ( .A(n90612), .B(n90611), .Z(n90613) );
  XOR U108818 ( .A(n90614), .B(n90613), .Z(n90615) );
  XOR U108819 ( .A(n90616), .B(n90615), .Z(n90626) );
  IV U108820 ( .A(n90617), .Z(n90619) );
  NOR U108821 ( .A(n90619), .B(n90618), .Z(n90624) );
  IV U108822 ( .A(n90620), .Z(n90621) );
  NOR U108823 ( .A(n90622), .B(n90621), .Z(n90623) );
  NOR U108824 ( .A(n90624), .B(n90623), .Z(n90625) );
  XOR U108825 ( .A(n90626), .B(n90625), .Z(n90650) );
  IV U108826 ( .A(n90627), .Z(n90629) );
  NOR U108827 ( .A(n90629), .B(n90628), .Z(n90630) );
  NOR U108828 ( .A(n90631), .B(n90630), .Z(n90637) );
  NOR U108829 ( .A(n90633), .B(n90632), .Z(n90634) );
  NOR U108830 ( .A(n90635), .B(n90634), .Z(n90636) );
  XOR U108831 ( .A(n90637), .B(n90636), .Z(n90648) );
  IV U108832 ( .A(n90642), .Z(n90639) );
  NOR U108833 ( .A(n90639), .B(n90638), .Z(n90646) );
  IV U108834 ( .A(n90640), .Z(n90644) );
  NOR U108835 ( .A(n90642), .B(n90641), .Z(n90643) );
  NOR U108836 ( .A(n90644), .B(n90643), .Z(n90645) );
  NOR U108837 ( .A(n90646), .B(n90645), .Z(n90647) );
  XOR U108838 ( .A(n90648), .B(n90647), .Z(n90649) );
  XOR U108839 ( .A(n90650), .B(n90649), .Z(n90651) );
  XOR U108840 ( .A(n90652), .B(n90651), .Z(n90664) );
  IV U108841 ( .A(n90656), .Z(n90653) );
  NOR U108842 ( .A(n90654), .B(n90653), .Z(n90662) );
  IV U108843 ( .A(n90654), .Z(n90655) );
  NOR U108844 ( .A(n90656), .B(n90655), .Z(n90660) );
  XOR U108845 ( .A(n90658), .B(n90657), .Z(n90659) );
  NOR U108846 ( .A(n90660), .B(n90659), .Z(n90661) );
  NOR U108847 ( .A(n90662), .B(n90661), .Z(n90663) );
  XOR U108848 ( .A(n90664), .B(n90663), .Z(n90665) );
  XOR U108849 ( .A(n90666), .B(n90665), .Z(n90695) );
  IV U108850 ( .A(n90667), .Z(n90669) );
  NOR U108851 ( .A(n90669), .B(n90668), .Z(n90673) );
  NOR U108852 ( .A(n90671), .B(n90670), .Z(n90672) );
  NOR U108853 ( .A(n90673), .B(n90672), .Z(n90683) );
  IV U108854 ( .A(n90674), .Z(n90675) );
  NOR U108855 ( .A(n90676), .B(n90675), .Z(n90681) );
  IV U108856 ( .A(n90677), .Z(n90678) );
  NOR U108857 ( .A(n90679), .B(n90678), .Z(n90680) );
  NOR U108858 ( .A(n90681), .B(n90680), .Z(n90682) );
  XOR U108859 ( .A(n90683), .B(n90682), .Z(n90693) );
  IV U108860 ( .A(n90686), .Z(n90684) );
  NOR U108861 ( .A(n90685), .B(n90684), .Z(n90691) );
  IV U108862 ( .A(n90685), .Z(n90687) );
  NOR U108863 ( .A(n90687), .B(n90686), .Z(n90689) );
  NOR U108864 ( .A(n90689), .B(n90688), .Z(n90690) );
  NOR U108865 ( .A(n90691), .B(n90690), .Z(n90692) );
  XOR U108866 ( .A(n90693), .B(n90692), .Z(n90694) );
  XOR U108867 ( .A(n90695), .B(n90694), .Z(n90696) );
  XOR U108868 ( .A(n90697), .B(n90696), .Z(n90718) );
  IV U108869 ( .A(n90698), .Z(n90701) );
  IV U108870 ( .A(n90699), .Z(n90700) );
  NOR U108871 ( .A(n90701), .B(n90700), .Z(n90702) );
  NOR U108872 ( .A(n90703), .B(n90702), .Z(n90708) );
  XOR U108873 ( .A(n90708), .B(n90707), .Z(n90716) );
  IV U108874 ( .A(n90709), .Z(n90712) );
  IV U108875 ( .A(n90710), .Z(n90711) );
  NOR U108876 ( .A(n90712), .B(n90711), .Z(n90713) );
  NOR U108877 ( .A(n90714), .B(n90713), .Z(n90715) );
  XOR U108878 ( .A(n90716), .B(n90715), .Z(n90717) );
  XOR U108879 ( .A(n90718), .B(n90717), .Z(n90719) );
  XOR U108880 ( .A(n90720), .B(n90719), .Z(n90721) );
  XOR U108881 ( .A(n90722), .B(n90721), .Z(n90723) );
  IV U108882 ( .A(n90725), .Z(n90727) );
  NOR U108883 ( .A(n90727), .B(n90726), .Z(n90732) );
  IV U108884 ( .A(n90728), .Z(n90729) );
  NOR U108885 ( .A(n90730), .B(n90729), .Z(n90731) );
  IV U108886 ( .A(n90733), .Z(n90735) );
  NOR U108887 ( .A(n90735), .B(n90734), .Z(n90736) );
  IV U108888 ( .A(n90738), .Z(n90739) );
  IV U108889 ( .A(n90740), .Z(n90742) );
  XOR U108890 ( .A(n90744), .B(n90743), .Z(n90764) );
  NOR U108891 ( .A(n90746), .B(n90745), .Z(n90747) );
  NOR U108892 ( .A(n90748), .B(n90747), .Z(n90749) );
  NOR U108893 ( .A(n90750), .B(n90749), .Z(n90751) );
  XOR U108894 ( .A(n90752), .B(n90751), .Z(n90762) );
  IV U108895 ( .A(n90753), .Z(n90755) );
  NOR U108896 ( .A(n90755), .B(n90754), .Z(n90760) );
  IV U108897 ( .A(n90756), .Z(n90758) );
  NOR U108898 ( .A(n90758), .B(n90757), .Z(n90759) );
  NOR U108899 ( .A(n90760), .B(n90759), .Z(n90761) );
  XOR U108900 ( .A(n90762), .B(n90761), .Z(n90763) );
  XOR U108901 ( .A(n90764), .B(n90763), .Z(n90765) );
  XOR U108902 ( .A(n90766), .B(n90765), .Z(n90767) );
  XOR U108903 ( .A(n90768), .B(n90767), .Z(n90769) );
  XOR U108904 ( .A(n90770), .B(n90769), .Z(n90771) );
  XOR U108905 ( .A(n90772), .B(n90771), .Z(n90773) );
  XOR U108906 ( .A(n90774), .B(n90773), .Z(n90789) );
  IV U108907 ( .A(n90775), .Z(n90776) );
  NOR U108908 ( .A(n90777), .B(n90776), .Z(n90787) );
  IV U108909 ( .A(n90778), .Z(n90780) );
  NOR U108910 ( .A(n90780), .B(n90779), .Z(n90785) );
  IV U108911 ( .A(n90781), .Z(n90782) );
  NOR U108912 ( .A(n90783), .B(n90782), .Z(n90784) );
  NOR U108913 ( .A(n90785), .B(n90784), .Z(n90786) );
  XOR U108914 ( .A(n90787), .B(n90786), .Z(n90788) );
  XOR U108915 ( .A(n90789), .B(n90788), .Z(n90790) );
  XOR U108916 ( .A(n90791), .B(n90790), .Z(n90792) );
  XOR U108917 ( .A(n90793), .B(n90792), .Z(n90794) );
  XOR U108918 ( .A(n90795), .B(n90794), .Z(n90814) );
  NOR U108919 ( .A(n90797), .B(n90796), .Z(n90812) );
  IV U108920 ( .A(n90798), .Z(n90799) );
  NOR U108921 ( .A(n90800), .B(n90799), .Z(n90810) );
  XOR U108922 ( .A(n90803), .B(n90804), .Z(n90802) );
  NOR U108923 ( .A(n90802), .B(n90801), .Z(n90807) );
  IV U108924 ( .A(n90803), .Z(n90805) );
  NOR U108925 ( .A(n90805), .B(n90804), .Z(n90806) );
  NOR U108926 ( .A(n90807), .B(n90806), .Z(n90808) );
  IV U108927 ( .A(n90808), .Z(n90809) );
  NOR U108928 ( .A(n90810), .B(n90809), .Z(n90811) );
  XOR U108929 ( .A(n90812), .B(n90811), .Z(n90813) );
  XOR U108930 ( .A(n90814), .B(n90813), .Z(n90815) );
  XOR U108931 ( .A(n90816), .B(n90815), .Z(n90817) );
  XOR U108932 ( .A(n90818), .B(n90817), .Z(n90819) );
  XOR U108933 ( .A(n90820), .B(n90819), .Z(n90840) );
  IV U108934 ( .A(n90821), .Z(n90823) );
  NOR U108935 ( .A(n90823), .B(n90822), .Z(n90828) );
  IV U108936 ( .A(n90824), .Z(n90826) );
  NOR U108937 ( .A(n90826), .B(n90825), .Z(n90827) );
  NOR U108938 ( .A(n90828), .B(n90827), .Z(n90838) );
  IV U108939 ( .A(n90832), .Z(n90829) );
  NOR U108940 ( .A(n90831), .B(n90829), .Z(n90836) );
  IV U108941 ( .A(n90830), .Z(n90834) );
  XOR U108942 ( .A(n90832), .B(n90831), .Z(n90833) );
  NOR U108943 ( .A(n90834), .B(n90833), .Z(n90835) );
  NOR U108944 ( .A(n90836), .B(n90835), .Z(n90837) );
  XOR U108945 ( .A(n90838), .B(n90837), .Z(n90839) );
  XOR U108946 ( .A(n90840), .B(n90839), .Z(n90841) );
  XOR U108947 ( .A(n90842), .B(n90841), .Z(n90863) );
  NOR U108948 ( .A(n90843), .B(n90844), .Z(n90850) );
  IV U108949 ( .A(n90844), .Z(n90845) );
  NOR U108950 ( .A(n90846), .B(n90845), .Z(n90847) );
  NOR U108951 ( .A(n90848), .B(n90847), .Z(n90849) );
  NOR U108952 ( .A(n90850), .B(n90849), .Z(n90861) );
  IV U108953 ( .A(n90851), .Z(n90854) );
  IV U108954 ( .A(n90852), .Z(n90853) );
  NOR U108955 ( .A(n90854), .B(n90853), .Z(n90859) );
  IV U108956 ( .A(n90855), .Z(n90856) );
  NOR U108957 ( .A(n90857), .B(n90856), .Z(n90858) );
  NOR U108958 ( .A(n90859), .B(n90858), .Z(n90860) );
  XOR U108959 ( .A(n90861), .B(n90860), .Z(n90862) );
  XOR U108960 ( .A(n90863), .B(n90862), .Z(n90864) );
  XOR U108961 ( .A(n90865), .B(n90864), .Z(n90866) );
  XOR U108962 ( .A(n90867), .B(n90866), .Z(n90868) );
  XOR U108963 ( .A(n90869), .B(n90868), .Z(n90870) );
  XOR U108964 ( .A(n90871), .B(n90870), .Z(n90872) );
  XOR U108965 ( .A(n90873), .B(n90872), .Z(n90893) );
  IV U108966 ( .A(n90874), .Z(n90876) );
  NOR U108967 ( .A(n90876), .B(n90875), .Z(n90881) );
  IV U108968 ( .A(n90877), .Z(n90879) );
  NOR U108969 ( .A(n90879), .B(n90878), .Z(n90880) );
  NOR U108970 ( .A(n90881), .B(n90880), .Z(n90891) );
  IV U108971 ( .A(n90882), .Z(n90883) );
  NOR U108972 ( .A(n90884), .B(n90883), .Z(n90889) );
  IV U108973 ( .A(n90885), .Z(n90886) );
  NOR U108974 ( .A(n90887), .B(n90886), .Z(n90888) );
  NOR U108975 ( .A(n90889), .B(n90888), .Z(n90890) );
  XOR U108976 ( .A(n90891), .B(n90890), .Z(n90892) );
  NOR U108977 ( .A(n90895), .B(n90894), .Z(n90896) );
  IV U108978 ( .A(n90896), .Z(n90903) );
  XOR U108979 ( .A(n90898), .B(n90897), .Z(n90899) );
  NOR U108980 ( .A(n90900), .B(n90899), .Z(n90901) );
  IV U108981 ( .A(n90901), .Z(n90902) );
  NOR U108982 ( .A(n90903), .B(n90902), .Z(n90904) );
  NOR U108983 ( .A(n90907), .B(n90906), .Z(n90909) );
  NOR U108984 ( .A(n90909), .B(n90908), .Z(n90910) );
  IV U108985 ( .A(n90911), .Z(n90913) );
  NOR U108986 ( .A(n90913), .B(n90912), .Z(n90914) );
  IV U108987 ( .A(n90916), .Z(n90918) );
  NOR U108988 ( .A(n90918), .B(n90917), .Z(n90922) );
  NOR U108989 ( .A(n90920), .B(n90919), .Z(n90921) );
  XOR U108990 ( .A(n90924), .B(n90923), .Z(n90943) );
  IV U108991 ( .A(n90925), .Z(n90927) );
  NOR U108992 ( .A(n90927), .B(n90926), .Z(n90931) );
  NOR U108993 ( .A(n90929), .B(n90928), .Z(n90930) );
  NOR U108994 ( .A(n90931), .B(n90930), .Z(n90941) );
  IV U108995 ( .A(n90932), .Z(n90934) );
  NOR U108996 ( .A(n90934), .B(n90933), .Z(n90939) );
  IV U108997 ( .A(n90935), .Z(n90936) );
  NOR U108998 ( .A(n90937), .B(n90936), .Z(n90938) );
  NOR U108999 ( .A(n90939), .B(n90938), .Z(n90940) );
  XOR U109000 ( .A(n90941), .B(n90940), .Z(n90942) );
  XOR U109001 ( .A(n90943), .B(n90942), .Z(n90944) );
  XOR U109002 ( .A(n90945), .B(n90944), .Z(n90946) );
  XOR U109003 ( .A(n90947), .B(n90946), .Z(n90948) );
  XOR U109004 ( .A(n90949), .B(n90948), .Z(n90969) );
  IV U109005 ( .A(n90950), .Z(n90952) );
  NOR U109006 ( .A(n90952), .B(n90951), .Z(n90957) );
  IV U109007 ( .A(n90953), .Z(n90954) );
  NOR U109008 ( .A(n90955), .B(n90954), .Z(n90956) );
  NOR U109009 ( .A(n90957), .B(n90956), .Z(n90967) );
  IV U109010 ( .A(n90958), .Z(n90960) );
  NOR U109011 ( .A(n90960), .B(n90959), .Z(n90965) );
  IV U109012 ( .A(n90961), .Z(n90962) );
  NOR U109013 ( .A(n90963), .B(n90962), .Z(n90964) );
  NOR U109014 ( .A(n90965), .B(n90964), .Z(n90966) );
  XOR U109015 ( .A(n90967), .B(n90966), .Z(n90968) );
  XOR U109016 ( .A(n90969), .B(n90968), .Z(n90970) );
  XOR U109017 ( .A(n90971), .B(n90970), .Z(n90993) );
  IV U109018 ( .A(n90972), .Z(n90974) );
  NOR U109019 ( .A(n90974), .B(n90973), .Z(n90978) );
  IV U109020 ( .A(n90975), .Z(n90976) );
  NOR U109021 ( .A(n90976), .B(n90983), .Z(n90977) );
  NOR U109022 ( .A(n90978), .B(n90977), .Z(n90991) );
  IV U109023 ( .A(n90979), .Z(n90980) );
  NOR U109024 ( .A(n90981), .B(n90980), .Z(n90989) );
  IV U109025 ( .A(n90982), .Z(n90984) );
  NOR U109026 ( .A(n90984), .B(n90983), .Z(n90985) );
  NOR U109027 ( .A(n90986), .B(n90985), .Z(n90987) );
  IV U109028 ( .A(n90987), .Z(n90988) );
  NOR U109029 ( .A(n90989), .B(n90988), .Z(n90990) );
  XOR U109030 ( .A(n90991), .B(n90990), .Z(n90992) );
  XOR U109031 ( .A(n90993), .B(n90992), .Z(n90994) );
  XOR U109032 ( .A(n90995), .B(n90994), .Z(n90996) );
  XOR U109033 ( .A(n90997), .B(n90996), .Z(n90998) );
  XOR U109034 ( .A(n90999), .B(n90998), .Z(n91025) );
  IV U109035 ( .A(n91000), .Z(n91002) );
  NOR U109036 ( .A(n91002), .B(n91001), .Z(n91007) );
  IV U109037 ( .A(n91003), .Z(n91005) );
  NOR U109038 ( .A(n91005), .B(n91004), .Z(n91006) );
  NOR U109039 ( .A(n91007), .B(n91006), .Z(n91023) );
  IV U109040 ( .A(n91008), .Z(n91010) );
  NOR U109041 ( .A(n91010), .B(n91009), .Z(n91021) );
  IV U109042 ( .A(n91011), .Z(n91013) );
  NOR U109043 ( .A(n91013), .B(n91012), .Z(n91018) );
  IV U109044 ( .A(n91014), .Z(n91016) );
  NOR U109045 ( .A(n91016), .B(n91015), .Z(n91017) );
  NOR U109046 ( .A(n91018), .B(n91017), .Z(n91019) );
  IV U109047 ( .A(n91019), .Z(n91020) );
  NOR U109048 ( .A(n91021), .B(n91020), .Z(n91022) );
  XOR U109049 ( .A(n91023), .B(n91022), .Z(n91024) );
  XOR U109050 ( .A(n91025), .B(n91024), .Z(n91026) );
  XOR U109051 ( .A(n91027), .B(n91026), .Z(n91047) );
  NOR U109052 ( .A(n91029), .B(n91028), .Z(n91035) );
  IV U109053 ( .A(n91030), .Z(n91031) );
  NOR U109054 ( .A(n91031), .B(n91060), .Z(n91032) );
  NOR U109055 ( .A(n91033), .B(n91032), .Z(n91034) );
  XOR U109056 ( .A(n91035), .B(n91034), .Z(n91045) );
  IV U109057 ( .A(n91036), .Z(n91038) );
  NOR U109058 ( .A(n91038), .B(n91037), .Z(n91043) );
  IV U109059 ( .A(n91039), .Z(n91041) );
  NOR U109060 ( .A(n91041), .B(n91040), .Z(n91042) );
  NOR U109061 ( .A(n91043), .B(n91042), .Z(n91044) );
  XOR U109062 ( .A(n91045), .B(n91044), .Z(n91046) );
  XOR U109063 ( .A(n91047), .B(n91046), .Z(n91067) );
  NOR U109064 ( .A(n91049), .B(n91048), .Z(n91053) );
  XOR U109065 ( .A(n91050), .B(n91053), .Z(n91055) );
  IV U109066 ( .A(n91051), .Z(n91052) );
  NOR U109067 ( .A(n91053), .B(n91052), .Z(n91054) );
  NOR U109068 ( .A(n91055), .B(n91054), .Z(n91065) );
  IV U109069 ( .A(n91056), .Z(n91057) );
  NOR U109070 ( .A(n91058), .B(n91057), .Z(n91063) );
  IV U109071 ( .A(n91059), .Z(n91061) );
  NOR U109072 ( .A(n91061), .B(n91060), .Z(n91062) );
  NOR U109073 ( .A(n91063), .B(n91062), .Z(n91064) );
  XOR U109074 ( .A(n91065), .B(n91064), .Z(n91066) );
  XOR U109075 ( .A(n91067), .B(n91066), .Z(n91087) );
  NOR U109076 ( .A(n91069), .B(n91068), .Z(n91075) );
  NOR U109077 ( .A(n91071), .B(n91070), .Z(n91072) );
  NOR U109078 ( .A(n91073), .B(n91072), .Z(n91074) );
  NOR U109079 ( .A(n91075), .B(n91074), .Z(n91085) );
  IV U109080 ( .A(n91076), .Z(n91077) );
  NOR U109081 ( .A(n91078), .B(n91077), .Z(n91083) );
  IV U109082 ( .A(n91079), .Z(n91080) );
  NOR U109083 ( .A(n91081), .B(n91080), .Z(n91082) );
  NOR U109084 ( .A(n91083), .B(n91082), .Z(n91084) );
  XOR U109085 ( .A(n91085), .B(n91084), .Z(n91086) );
  XOR U109086 ( .A(n91087), .B(n91086), .Z(n91088) );
  XOR U109087 ( .A(n91089), .B(n91088), .Z(n91112) );
  IV U109088 ( .A(n91090), .Z(n91091) );
  NOR U109089 ( .A(n91092), .B(n91091), .Z(n91097) );
  IV U109090 ( .A(n91093), .Z(n91094) );
  NOR U109091 ( .A(n91095), .B(n91094), .Z(n91096) );
  NOR U109092 ( .A(n91097), .B(n91096), .Z(n91110) );
  IV U109093 ( .A(n91098), .Z(n91099) );
  NOR U109094 ( .A(n91099), .B(n91121), .Z(n91108) );
  NOR U109095 ( .A(n91101), .B(n91100), .Z(n91106) );
  IV U109096 ( .A(n91102), .Z(n91103) );
  NOR U109097 ( .A(n91104), .B(n91103), .Z(n91105) );
  NOR U109098 ( .A(n91106), .B(n91105), .Z(n91107) );
  XOR U109099 ( .A(n91108), .B(n91107), .Z(n91109) );
  XOR U109100 ( .A(n91110), .B(n91109), .Z(n91111) );
  XOR U109101 ( .A(n91112), .B(n91111), .Z(n91128) );
  IV U109102 ( .A(n91113), .Z(n91114) );
  NOR U109103 ( .A(n91115), .B(n91114), .Z(n91119) );
  NOR U109104 ( .A(n91117), .B(n91116), .Z(n91118) );
  NOR U109105 ( .A(n91119), .B(n91118), .Z(n91126) );
  IV U109106 ( .A(n91120), .Z(n91122) );
  NOR U109107 ( .A(n91122), .B(n91121), .Z(n91124) );
  NOR U109108 ( .A(n91124), .B(n91123), .Z(n91125) );
  XOR U109109 ( .A(n91126), .B(n91125), .Z(n91127) );
  XOR U109110 ( .A(n91128), .B(n91127), .Z(n91129) );
  XOR U109111 ( .A(n91130), .B(n91129), .Z(n91140) );
  NOR U109112 ( .A(n91132), .B(n91131), .Z(n91138) );
  IV U109113 ( .A(n91133), .Z(n91136) );
  IV U109114 ( .A(n91134), .Z(n91135) );
  NOR U109115 ( .A(n91136), .B(n91135), .Z(n91137) );
  XOR U109116 ( .A(n91138), .B(n91137), .Z(n91139) );
  XOR U109117 ( .A(n91140), .B(n91139), .Z(n91141) );
  XOR U109118 ( .A(n91142), .B(n91141), .Z(n91156) );
  NOR U109119 ( .A(n91144), .B(n91143), .Z(n91154) );
  IV U109120 ( .A(n91145), .Z(n91147) );
  NOR U109121 ( .A(n91147), .B(n91146), .Z(n91152) );
  IV U109122 ( .A(n91148), .Z(n91149) );
  NOR U109123 ( .A(n91150), .B(n91149), .Z(n91151) );
  NOR U109124 ( .A(n91152), .B(n91151), .Z(n91153) );
  XOR U109125 ( .A(n91154), .B(n91153), .Z(n91155) );
  XOR U109126 ( .A(n91156), .B(n91155), .Z(n91174) );
  IV U109127 ( .A(n91157), .Z(n91158) );
  NOR U109128 ( .A(n91159), .B(n91158), .Z(n91172) );
  IV U109129 ( .A(n91160), .Z(n91161) );
  NOR U109130 ( .A(n91162), .B(n91161), .Z(n91170) );
  IV U109131 ( .A(n91163), .Z(n91168) );
  NOR U109132 ( .A(n91165), .B(n91164), .Z(n91166) );
  IV U109133 ( .A(n91166), .Z(n91167) );
  NOR U109134 ( .A(n91168), .B(n91167), .Z(n91169) );
  XOR U109135 ( .A(n91170), .B(n91169), .Z(n91171) );
  XOR U109136 ( .A(n91172), .B(n91171), .Z(n91173) );
  XOR U109137 ( .A(n91174), .B(n91173), .Z(n91212) );
  IV U109138 ( .A(n91175), .Z(n91177) );
  NOR U109139 ( .A(n91177), .B(n91176), .Z(n91185) );
  NOR U109140 ( .A(n91179), .B(n91178), .Z(n91183) );
  NOR U109141 ( .A(n91181), .B(n91180), .Z(n91182) );
  NOR U109142 ( .A(n91183), .B(n91182), .Z(n91184) );
  XOR U109143 ( .A(n91185), .B(n91184), .Z(n91210) );
  IV U109144 ( .A(n91186), .Z(n91187) );
  NOR U109145 ( .A(n91188), .B(n91187), .Z(n91192) );
  NOR U109146 ( .A(n91190), .B(n91189), .Z(n91191) );
  NOR U109147 ( .A(n91192), .B(n91191), .Z(n91208) );
  IV U109148 ( .A(n91193), .Z(n91195) );
  NOR U109149 ( .A(n91195), .B(n91194), .Z(n91206) );
  IV U109150 ( .A(n91196), .Z(n91198) );
  NOR U109151 ( .A(n91198), .B(n91197), .Z(n91203) );
  IV U109152 ( .A(n91199), .Z(n91200) );
  NOR U109153 ( .A(n91201), .B(n91200), .Z(n91202) );
  NOR U109154 ( .A(n91203), .B(n91202), .Z(n91204) );
  IV U109155 ( .A(n91204), .Z(n91205) );
  NOR U109156 ( .A(n91206), .B(n91205), .Z(n91207) );
  XOR U109157 ( .A(n91208), .B(n91207), .Z(n91209) );
  XOR U109158 ( .A(n91210), .B(n91209), .Z(n91211) );
  XOR U109159 ( .A(n91212), .B(n91211), .Z(n91213) );
  XOR U109160 ( .A(n91214), .B(n91213), .Z(n91215) );
  XOR U109161 ( .A(n91216), .B(n91215), .Z(n91225) );
  IV U109162 ( .A(n91217), .Z(n91219) );
  NOR U109163 ( .A(n91219), .B(n91218), .Z(n91223) );
  NOR U109164 ( .A(n91221), .B(n91220), .Z(n91222) );
  NOR U109165 ( .A(n91223), .B(n91222), .Z(n91224) );
  XOR U109166 ( .A(n91225), .B(n91224), .Z(n91237) );
  IV U109167 ( .A(n91231), .Z(n91226) );
  NOR U109168 ( .A(n91227), .B(n91226), .Z(n91235) );
  XOR U109169 ( .A(n91229), .B(n91228), .Z(n91230) );
  NOR U109170 ( .A(n91231), .B(n91230), .Z(n91233) );
  NOR U109171 ( .A(n91233), .B(n91232), .Z(n91234) );
  NOR U109172 ( .A(n91235), .B(n91234), .Z(n91236) );
  XOR U109173 ( .A(n91237), .B(n91236), .Z(n91263) );
  NOR U109174 ( .A(n91239), .B(n91238), .Z(n91261) );
  IV U109175 ( .A(n91240), .Z(n91243) );
  IV U109176 ( .A(n91241), .Z(n91242) );
  NOR U109177 ( .A(n91243), .B(n91242), .Z(n91248) );
  IV U109178 ( .A(n91244), .Z(n91245) );
  NOR U109179 ( .A(n91246), .B(n91245), .Z(n91247) );
  NOR U109180 ( .A(n91248), .B(n91247), .Z(n91259) );
  IV U109181 ( .A(n91252), .Z(n91249) );
  NOR U109182 ( .A(n91250), .B(n91249), .Z(n91257) );
  IV U109183 ( .A(n91251), .Z(n91255) );
  NOR U109184 ( .A(n91253), .B(n91252), .Z(n91254) );
  NOR U109185 ( .A(n91255), .B(n91254), .Z(n91256) );
  NOR U109186 ( .A(n91257), .B(n91256), .Z(n91258) );
  XOR U109187 ( .A(n91259), .B(n91258), .Z(n91260) );
  XOR U109188 ( .A(n91261), .B(n91260), .Z(n91262) );
  XOR U109189 ( .A(n91263), .B(n91262), .Z(n91264) );
  XOR U109190 ( .A(n91265), .B(n91264), .Z(n91266) );
  XOR U109191 ( .A(n91267), .B(n91266), .Z(n91280) );
  IV U109192 ( .A(n91268), .Z(n91270) );
  NOR U109193 ( .A(n91270), .B(n91269), .Z(n91274) );
  NOR U109194 ( .A(n91272), .B(n91271), .Z(n91273) );
  NOR U109195 ( .A(n91274), .B(n91273), .Z(n91278) );
  NOR U109196 ( .A(n91276), .B(n91275), .Z(n91277) );
  XOR U109197 ( .A(n91278), .B(n91277), .Z(n91279) );
  XOR U109198 ( .A(n91280), .B(n91279), .Z(n91281) );
  XOR U109199 ( .A(n91282), .B(n91281), .Z(n91283) );
  XOR U109200 ( .A(n91284), .B(n91283), .Z(n91309) );
  IV U109201 ( .A(n91285), .Z(n91286) );
  NOR U109202 ( .A(n91287), .B(n91286), .Z(n91288) );
  NOR U109203 ( .A(n91289), .B(n91288), .Z(n91298) );
  IV U109204 ( .A(n91290), .Z(n91291) );
  NOR U109205 ( .A(n91292), .B(n91291), .Z(n91296) );
  IV U109206 ( .A(n91293), .Z(n91294) );
  NOR U109207 ( .A(n91294), .B(n91300), .Z(n91295) );
  NOR U109208 ( .A(n91296), .B(n91295), .Z(n91297) );
  XOR U109209 ( .A(n91298), .B(n91297), .Z(n91307) );
  IV U109210 ( .A(n91299), .Z(n91301) );
  NOR U109211 ( .A(n91301), .B(n91300), .Z(n91305) );
  NOR U109212 ( .A(n91303), .B(n91302), .Z(n91304) );
  NOR U109213 ( .A(n91305), .B(n91304), .Z(n91306) );
  XOR U109214 ( .A(n91307), .B(n91306), .Z(n91308) );
  XOR U109215 ( .A(n91309), .B(n91308), .Z(n91310) );
  XOR U109216 ( .A(n91311), .B(n91310), .Z(n91312) );
  XOR U109217 ( .A(n91313), .B(n91312), .Z(n91323) );
  NOR U109218 ( .A(n91314), .B(n91315), .Z(n91321) );
  IV U109219 ( .A(n91315), .Z(n91316) );
  NOR U109220 ( .A(n91317), .B(n91316), .Z(n91318) );
  NOR U109221 ( .A(n91319), .B(n91318), .Z(n91320) );
  NOR U109222 ( .A(n91321), .B(n91320), .Z(n91322) );
  XOR U109223 ( .A(n91323), .B(n91322), .Z(n91348) );
  IV U109224 ( .A(n91324), .Z(n91325) );
  NOR U109225 ( .A(n91326), .B(n91325), .Z(n91331) );
  IV U109226 ( .A(n91327), .Z(n91328) );
  NOR U109227 ( .A(n91329), .B(n91328), .Z(n91330) );
  NOR U109228 ( .A(n91331), .B(n91330), .Z(n91346) );
  NOR U109229 ( .A(n91333), .B(n91332), .Z(n91344) );
  IV U109230 ( .A(n91334), .Z(n91335) );
  NOR U109231 ( .A(n91336), .B(n91335), .Z(n91341) );
  IV U109232 ( .A(n91337), .Z(n91338) );
  NOR U109233 ( .A(n91339), .B(n91338), .Z(n91340) );
  NOR U109234 ( .A(n91341), .B(n91340), .Z(n91342) );
  IV U109235 ( .A(n91342), .Z(n91343) );
  NOR U109236 ( .A(n91344), .B(n91343), .Z(n91345) );
  XOR U109237 ( .A(n91346), .B(n91345), .Z(n91347) );
  XOR U109238 ( .A(n91348), .B(n91347), .Z(n91384) );
  NOR U109239 ( .A(n91349), .B(n91350), .Z(n91356) );
  IV U109240 ( .A(n91350), .Z(n91351) );
  NOR U109241 ( .A(n91352), .B(n91351), .Z(n91353) );
  NOR U109242 ( .A(n91354), .B(n91353), .Z(n91355) );
  NOR U109243 ( .A(n91356), .B(n91355), .Z(n91372) );
  IV U109244 ( .A(n91357), .Z(n91359) );
  NOR U109245 ( .A(n91359), .B(n91358), .Z(n91370) );
  IV U109246 ( .A(n91360), .Z(n91362) );
  NOR U109247 ( .A(n91362), .B(n91361), .Z(n91367) );
  IV U109248 ( .A(n91363), .Z(n91364) );
  NOR U109249 ( .A(n91365), .B(n91364), .Z(n91366) );
  NOR U109250 ( .A(n91367), .B(n91366), .Z(n91368) );
  IV U109251 ( .A(n91368), .Z(n91369) );
  NOR U109252 ( .A(n91370), .B(n91369), .Z(n91371) );
  XOR U109253 ( .A(n91372), .B(n91371), .Z(n91382) );
  IV U109254 ( .A(n91373), .Z(n91375) );
  NOR U109255 ( .A(n91375), .B(n91374), .Z(n91380) );
  IV U109256 ( .A(n91376), .Z(n91377) );
  NOR U109257 ( .A(n91378), .B(n91377), .Z(n91379) );
  NOR U109258 ( .A(n91380), .B(n91379), .Z(n91381) );
  XOR U109259 ( .A(n91382), .B(n91381), .Z(n91383) );
  XOR U109260 ( .A(n91384), .B(n91383), .Z(n91385) );
  XOR U109261 ( .A(n91386), .B(n91385), .Z(n91404) );
  NOR U109262 ( .A(n91388), .B(n91387), .Z(n91393) );
  IV U109263 ( .A(n91389), .Z(n91390) );
  NOR U109264 ( .A(n91391), .B(n91390), .Z(n91392) );
  NOR U109265 ( .A(n91393), .B(n91392), .Z(n91402) );
  NOR U109266 ( .A(n91395), .B(n91394), .Z(n91400) );
  IV U109267 ( .A(n91396), .Z(n91397) );
  NOR U109268 ( .A(n91398), .B(n91397), .Z(n91399) );
  NOR U109269 ( .A(n91400), .B(n91399), .Z(n91401) );
  XOR U109270 ( .A(n91402), .B(n91401), .Z(n91403) );
  XOR U109271 ( .A(n91404), .B(n91403), .Z(n91416) );
  NOR U109272 ( .A(n91405), .B(n91406), .Z(n91414) );
  IV U109273 ( .A(n91406), .Z(n91407) );
  NOR U109274 ( .A(n91408), .B(n91407), .Z(n91412) );
  XOR U109275 ( .A(n91410), .B(n91409), .Z(n91411) );
  NOR U109276 ( .A(n91412), .B(n91411), .Z(n91413) );
  NOR U109277 ( .A(n91414), .B(n91413), .Z(n91415) );
  XOR U109278 ( .A(n91416), .B(n91415), .Z(n91440) );
  IV U109279 ( .A(n91417), .Z(n91419) );
  NOR U109280 ( .A(n91419), .B(n91418), .Z(n91438) );
  NOR U109281 ( .A(n91421), .B(n91420), .Z(n91426) );
  IV U109282 ( .A(n91422), .Z(n91423) );
  NOR U109283 ( .A(n91424), .B(n91423), .Z(n91425) );
  NOR U109284 ( .A(n91426), .B(n91425), .Z(n91436) );
  IV U109285 ( .A(n91427), .Z(n91428) );
  NOR U109286 ( .A(n91429), .B(n91428), .Z(n91434) );
  IV U109287 ( .A(n91430), .Z(n91431) );
  NOR U109288 ( .A(n91432), .B(n91431), .Z(n91433) );
  NOR U109289 ( .A(n91434), .B(n91433), .Z(n91435) );
  XOR U109290 ( .A(n91436), .B(n91435), .Z(n91437) );
  XOR U109291 ( .A(n91438), .B(n91437), .Z(n91439) );
  XOR U109292 ( .A(n91440), .B(n91439), .Z(n91441) );
  XOR U109293 ( .A(n91442), .B(n91441), .Z(n91443) );
  XOR U109294 ( .A(n91444), .B(n91443), .Z(n91445) );
  XOR U109295 ( .A(n91446), .B(n91445), .Z(n91447) );
  XOR U109296 ( .A(n91448), .B(n91447), .Z(n91449) );
  XOR U109297 ( .A(n91450), .B(n91449), .Z(n91451) );
  XOR U109298 ( .A(n91452), .B(n91451), .Z(n91482) );
  IV U109299 ( .A(n91453), .Z(n91454) );
  NOR U109300 ( .A(n91455), .B(n91454), .Z(n91459) );
  NOR U109301 ( .A(n91457), .B(n91456), .Z(n91458) );
  NOR U109302 ( .A(n91459), .B(n91458), .Z(n91480) );
  IV U109303 ( .A(n91460), .Z(n91461) );
  NOR U109304 ( .A(n91462), .B(n91461), .Z(n91478) );
  IV U109305 ( .A(n91463), .Z(n91466) );
  NOR U109306 ( .A(n91464), .B(n91467), .Z(n91465) );
  NOR U109307 ( .A(n91466), .B(n91465), .Z(n91476) );
  IV U109308 ( .A(n91467), .Z(n91468) );
  NOR U109309 ( .A(n91469), .B(n91468), .Z(n91473) );
  NOR U109310 ( .A(n91471), .B(n91470), .Z(n91472) );
  NOR U109311 ( .A(n91473), .B(n91472), .Z(n91474) );
  IV U109312 ( .A(n91474), .Z(n91475) );
  NOR U109313 ( .A(n91476), .B(n91475), .Z(n91477) );
  XOR U109314 ( .A(n91478), .B(n91477), .Z(n91479) );
  XOR U109315 ( .A(n91480), .B(n91479), .Z(n91481) );
  XOR U109316 ( .A(n91482), .B(n91481), .Z(n91483) );
  XOR U109317 ( .A(n91484), .B(n91483), .Z(n91485) );
  XOR U109318 ( .A(n91486), .B(n91485), .Z(n91487) );
  XOR U109319 ( .A(n91488), .B(n91487), .Z(n91498) );
  IV U109320 ( .A(n91489), .Z(n91490) );
  NOR U109321 ( .A(n91491), .B(n91490), .Z(n91496) );
  IV U109322 ( .A(n91492), .Z(n91494) );
  NOR U109323 ( .A(n91494), .B(n91493), .Z(n91495) );
  NOR U109324 ( .A(n91496), .B(n91495), .Z(n91497) );
  XOR U109325 ( .A(n91498), .B(n91497), .Z(n91525) );
  IV U109326 ( .A(n91499), .Z(n91500) );
  NOR U109327 ( .A(n91501), .B(n91500), .Z(n91505) );
  IV U109328 ( .A(n91502), .Z(n91503) );
  NOR U109329 ( .A(n91504), .B(n91503), .Z(n91511) );
  XOR U109330 ( .A(n91505), .B(n91511), .Z(n91513) );
  IV U109331 ( .A(n91506), .Z(n91508) );
  NOR U109332 ( .A(n91508), .B(n91507), .Z(n91509) );
  IV U109333 ( .A(n91509), .Z(n91510) );
  NOR U109334 ( .A(n91511), .B(n91510), .Z(n91512) );
  NOR U109335 ( .A(n91513), .B(n91512), .Z(n91523) );
  NOR U109336 ( .A(n91515), .B(n91514), .Z(n91521) );
  IV U109337 ( .A(n91515), .Z(n91517) );
  NOR U109338 ( .A(n91517), .B(n91516), .Z(n91518) );
  NOR U109339 ( .A(n91519), .B(n91518), .Z(n91520) );
  NOR U109340 ( .A(n91521), .B(n91520), .Z(n91522) );
  XOR U109341 ( .A(n91523), .B(n91522), .Z(n91524) );
  XOR U109342 ( .A(n91525), .B(n91524), .Z(n91550) );
  NOR U109343 ( .A(n91526), .B(n91527), .Z(n91533) );
  IV U109344 ( .A(n91527), .Z(n91528) );
  NOR U109345 ( .A(n91529), .B(n91528), .Z(n91530) );
  NOR U109346 ( .A(n91531), .B(n91530), .Z(n91532) );
  NOR U109347 ( .A(n91533), .B(n91532), .Z(n91548) );
  NOR U109348 ( .A(n91535), .B(n91534), .Z(n91546) );
  IV U109349 ( .A(n91536), .Z(n91538) );
  NOR U109350 ( .A(n91538), .B(n91537), .Z(n91543) );
  IV U109351 ( .A(n91539), .Z(n91541) );
  NOR U109352 ( .A(n91541), .B(n91540), .Z(n91542) );
  NOR U109353 ( .A(n91543), .B(n91542), .Z(n91544) );
  IV U109354 ( .A(n91544), .Z(n91545) );
  NOR U109355 ( .A(n91546), .B(n91545), .Z(n91547) );
  XOR U109356 ( .A(n91548), .B(n91547), .Z(n91549) );
  XOR U109357 ( .A(n91550), .B(n91549), .Z(n91551) );
  XOR U109358 ( .A(n91552), .B(n91551), .Z(n91553) );
  XOR U109359 ( .A(n91554), .B(n91553), .Z(n91555) );
  XOR U109360 ( .A(n91556), .B(n91555), .Z(n91557) );
  XOR U109361 ( .A(n91558), .B(n91557), .Z(n91559) );
  XOR U109362 ( .A(n91560), .B(n91559), .Z(n91561) );
  XOR U109363 ( .A(n91562), .B(n91561), .Z(n91575) );
  NOR U109364 ( .A(n91564), .B(n91563), .Z(n91573) );
  IV U109365 ( .A(n91565), .Z(n91567) );
  NOR U109366 ( .A(n91567), .B(n91566), .Z(n91571) );
  NOR U109367 ( .A(n91569), .B(n91568), .Z(n91570) );
  NOR U109368 ( .A(n91571), .B(n91570), .Z(n91572) );
  XOR U109369 ( .A(n91573), .B(n91572), .Z(n91574) );
  XOR U109370 ( .A(n91575), .B(n91574), .Z(n91605) );
  IV U109371 ( .A(n91576), .Z(n91577) );
  NOR U109372 ( .A(n91577), .B(n91582), .Z(n91580) );
  NOR U109373 ( .A(n91578), .B(n91595), .Z(n91579) );
  NOR U109374 ( .A(n91580), .B(n91579), .Z(n91590) );
  IV U109375 ( .A(n91583), .Z(n91581) );
  NOR U109376 ( .A(n91581), .B(n91582), .Z(n91588) );
  XOR U109377 ( .A(n91583), .B(n91582), .Z(n91586) );
  IV U109378 ( .A(n91584), .Z(n91585) );
  NOR U109379 ( .A(n91586), .B(n91585), .Z(n91587) );
  NOR U109380 ( .A(n91588), .B(n91587), .Z(n91589) );
  XOR U109381 ( .A(n91590), .B(n91589), .Z(n91603) );
  IV U109382 ( .A(n91591), .Z(n91592) );
  NOR U109383 ( .A(n91593), .B(n91592), .Z(n91601) );
  IV U109384 ( .A(n91594), .Z(n91596) );
  NOR U109385 ( .A(n91596), .B(n91595), .Z(n91597) );
  NOR U109386 ( .A(n91598), .B(n91597), .Z(n91599) );
  IV U109387 ( .A(n91599), .Z(n91600) );
  NOR U109388 ( .A(n91601), .B(n91600), .Z(n91602) );
  XOR U109389 ( .A(n91603), .B(n91602), .Z(n91604) );
  XOR U109390 ( .A(n91605), .B(n91604), .Z(n91606) );
  XOR U109391 ( .A(n91607), .B(n91606), .Z(n91626) );
  IV U109392 ( .A(n91608), .Z(n91610) );
  NOR U109393 ( .A(n91610), .B(n91609), .Z(n91615) );
  IV U109394 ( .A(n91611), .Z(n91612) );
  NOR U109395 ( .A(n91613), .B(n91612), .Z(n91614) );
  NOR U109396 ( .A(n91615), .B(n91614), .Z(n91624) );
  IV U109397 ( .A(n91616), .Z(n91618) );
  NOR U109398 ( .A(n91618), .B(n91617), .Z(n91622) );
  NOR U109399 ( .A(n91620), .B(n91619), .Z(n91621) );
  NOR U109400 ( .A(n91622), .B(n91621), .Z(n91623) );
  XOR U109401 ( .A(n91624), .B(n91623), .Z(n91625) );
  XOR U109402 ( .A(n91626), .B(n91625), .Z(n91627) );
  XOR U109403 ( .A(n91628), .B(n91627), .Z(n91638) );
  IV U109404 ( .A(n91629), .Z(n91631) );
  NOR U109405 ( .A(n91631), .B(n91630), .Z(n91636) );
  IV U109406 ( .A(n91632), .Z(n91634) );
  NOR U109407 ( .A(n91634), .B(n91633), .Z(n91635) );
  NOR U109408 ( .A(n91636), .B(n91635), .Z(n91637) );
  XOR U109409 ( .A(n91638), .B(n91637), .Z(n91650) );
  NOR U109410 ( .A(n91639), .B(n91640), .Z(n91648) );
  IV U109411 ( .A(n91640), .Z(n91641) );
  NOR U109412 ( .A(n91642), .B(n91641), .Z(n91646) );
  XOR U109413 ( .A(n91644), .B(n91643), .Z(n91645) );
  NOR U109414 ( .A(n91646), .B(n91645), .Z(n91647) );
  NOR U109415 ( .A(n91648), .B(n91647), .Z(n91649) );
  XOR U109416 ( .A(n91650), .B(n91649), .Z(n91651) );
  XOR U109417 ( .A(n91652), .B(n91651), .Z(n91653) );
  XOR U109418 ( .A(n91654), .B(n91653), .Z(n91680) );
  IV U109419 ( .A(n91655), .Z(n91656) );
  NOR U109420 ( .A(n91656), .B(n91673), .Z(n91669) );
  IV U109421 ( .A(n91657), .Z(n91658) );
  NOR U109422 ( .A(n91659), .B(n91658), .Z(n91667) );
  IV U109423 ( .A(n91660), .Z(n91662) );
  NOR U109424 ( .A(n91662), .B(n91661), .Z(n91663) );
  NOR U109425 ( .A(n91664), .B(n91663), .Z(n91665) );
  IV U109426 ( .A(n91665), .Z(n91666) );
  NOR U109427 ( .A(n91667), .B(n91666), .Z(n91668) );
  XOR U109428 ( .A(n91669), .B(n91668), .Z(n91678) );
  NOR U109429 ( .A(n91671), .B(n91670), .Z(n91676) );
  IV U109430 ( .A(n91672), .Z(n91674) );
  NOR U109431 ( .A(n91674), .B(n91673), .Z(n91675) );
  NOR U109432 ( .A(n91676), .B(n91675), .Z(n91677) );
  XOR U109433 ( .A(n91678), .B(n91677), .Z(n91679) );
  XOR U109434 ( .A(n91680), .B(n91679), .Z(n91681) );
  XOR U109435 ( .A(n91682), .B(n91681), .Z(n91697) );
  IV U109436 ( .A(n91683), .Z(n91684) );
  NOR U109437 ( .A(n91689), .B(n91684), .Z(n91695) );
  IV U109438 ( .A(n91685), .Z(n91687) );
  NOR U109439 ( .A(n91687), .B(n91686), .Z(n91692) );
  IV U109440 ( .A(n91688), .Z(n91690) );
  NOR U109441 ( .A(n91690), .B(n91689), .Z(n91691) );
  NOR U109442 ( .A(n91692), .B(n91691), .Z(n91693) );
  IV U109443 ( .A(n91693), .Z(n91694) );
  NOR U109444 ( .A(n91695), .B(n91694), .Z(n91696) );
  XOR U109445 ( .A(n91697), .B(n91696), .Z(n91698) );
  XOR U109446 ( .A(n91699), .B(n91698), .Z(n91700) );
  XOR U109447 ( .A(n91701), .B(n91700), .Z(n91717) );
  IV U109448 ( .A(n91702), .Z(n91705) );
  IV U109449 ( .A(n91703), .Z(n91704) );
  NOR U109450 ( .A(n91705), .B(n91704), .Z(n91715) );
  IV U109451 ( .A(n91706), .Z(n91710) );
  XOR U109452 ( .A(n91707), .B(n91710), .Z(n91709) );
  NOR U109453 ( .A(n91709), .B(n91708), .Z(n91713) );
  NOR U109454 ( .A(n91711), .B(n91710), .Z(n91712) );
  NOR U109455 ( .A(n91713), .B(n91712), .Z(n91714) );
  XOR U109456 ( .A(n91715), .B(n91714), .Z(n91716) );
  XOR U109457 ( .A(n91717), .B(n91716), .Z(n91718) );
  XOR U109458 ( .A(n91719), .B(n91718), .Z(n91720) );
  XOR U109459 ( .A(n91721), .B(n91720), .Z(n91722) );
  XOR U109460 ( .A(n91723), .B(n91722), .Z(n91724) );
  XOR U109461 ( .A(n91725), .B(n91724), .Z(n91726) );
  XOR U109462 ( .A(n91727), .B(n91726), .Z(n91728) );
  XOR U109463 ( .A(n91729), .B(n91728), .Z(n91730) );
  XOR U109464 ( .A(n91731), .B(n91730), .Z(n91732) );
  XOR U109465 ( .A(n91733), .B(n91732), .Z(n91762) );
  IV U109466 ( .A(n91734), .Z(n91736) );
  NOR U109467 ( .A(n91736), .B(n91735), .Z(n91741) );
  IV U109468 ( .A(n91737), .Z(n91738) );
  NOR U109469 ( .A(n91739), .B(n91738), .Z(n91740) );
  NOR U109470 ( .A(n91741), .B(n91740), .Z(n91751) );
  NOR U109471 ( .A(n91742), .B(n91743), .Z(n91749) );
  IV U109472 ( .A(n91743), .Z(n91744) );
  NOR U109473 ( .A(n91745), .B(n91744), .Z(n91746) );
  NOR U109474 ( .A(n91747), .B(n91746), .Z(n91748) );
  NOR U109475 ( .A(n91749), .B(n91748), .Z(n91750) );
  XOR U109476 ( .A(n91751), .B(n91750), .Z(n91760) );
  IV U109477 ( .A(n91752), .Z(n91754) );
  NOR U109478 ( .A(n91754), .B(n91753), .Z(n91758) );
  NOR U109479 ( .A(n91756), .B(n91755), .Z(n91757) );
  NOR U109480 ( .A(n91758), .B(n91757), .Z(n91759) );
  XOR U109481 ( .A(n91760), .B(n91759), .Z(n91761) );
  XOR U109482 ( .A(n91762), .B(n91761), .Z(n91763) );
  XOR U109483 ( .A(n91764), .B(n91763), .Z(n91779) );
  IV U109484 ( .A(n91768), .Z(n91769) );
  NOR U109485 ( .A(n91770), .B(n91769), .Z(n91775) );
  IV U109486 ( .A(n91771), .Z(n91772) );
  NOR U109487 ( .A(n91773), .B(n91772), .Z(n91774) );
  NOR U109488 ( .A(n91775), .B(n91774), .Z(n91776) );
  XOR U109489 ( .A(n91777), .B(n91776), .Z(n91778) );
  XOR U109490 ( .A(n91779), .B(n91778), .Z(n91805) );
  IV U109491 ( .A(n91780), .Z(n91783) );
  NOR U109492 ( .A(n91784), .B(n91781), .Z(n91782) );
  NOR U109493 ( .A(n91783), .B(n91782), .Z(n91794) );
  IV U109494 ( .A(n91784), .Z(n91786) );
  NOR U109495 ( .A(n91786), .B(n91785), .Z(n91791) );
  IV U109496 ( .A(n91787), .Z(n91789) );
  NOR U109497 ( .A(n91789), .B(n91788), .Z(n91790) );
  NOR U109498 ( .A(n91791), .B(n91790), .Z(n91792) );
  IV U109499 ( .A(n91792), .Z(n91793) );
  NOR U109500 ( .A(n91794), .B(n91793), .Z(n91803) );
  NOR U109501 ( .A(n91796), .B(n91795), .Z(n91801) );
  IV U109502 ( .A(n91797), .Z(n91799) );
  NOR U109503 ( .A(n91799), .B(n91798), .Z(n91800) );
  NOR U109504 ( .A(n91801), .B(n91800), .Z(n91802) );
  XOR U109505 ( .A(n91803), .B(n91802), .Z(n91804) );
  XOR U109506 ( .A(n91805), .B(n91804), .Z(n91806) );
  XOR U109507 ( .A(n91807), .B(n91806), .Z(n91831) );
  NOR U109508 ( .A(n91809), .B(n91808), .Z(n91810) );
  NOR U109509 ( .A(n91811), .B(n91810), .Z(n91822) );
  IV U109510 ( .A(n91812), .Z(n91814) );
  NOR U109511 ( .A(n91814), .B(n91813), .Z(n91819) );
  IV U109512 ( .A(n91815), .Z(n91817) );
  NOR U109513 ( .A(n91817), .B(n91816), .Z(n91818) );
  NOR U109514 ( .A(n91819), .B(n91818), .Z(n91820) );
  IV U109515 ( .A(n91820), .Z(n91821) );
  NOR U109516 ( .A(n91822), .B(n91821), .Z(n91829) );
  IV U109517 ( .A(n91823), .Z(n91825) );
  NOR U109518 ( .A(n91825), .B(n91824), .Z(n91826) );
  NOR U109519 ( .A(n91827), .B(n91826), .Z(n91828) );
  XOR U109520 ( .A(n91829), .B(n91828), .Z(n91830) );
  XOR U109521 ( .A(n91831), .B(n91830), .Z(n91847) );
  IV U109522 ( .A(n91832), .Z(n91834) );
  XOR U109523 ( .A(n91838), .B(n91840), .Z(n91833) );
  NOR U109524 ( .A(n91834), .B(n91833), .Z(n91845) );
  IV U109525 ( .A(n91835), .Z(n91836) );
  NOR U109526 ( .A(n91837), .B(n91836), .Z(n91842) );
  IV U109527 ( .A(n91838), .Z(n91839) );
  NOR U109528 ( .A(n91840), .B(n91839), .Z(n91841) );
  NOR U109529 ( .A(n91842), .B(n91841), .Z(n91843) );
  IV U109530 ( .A(n91843), .Z(n91844) );
  NOR U109531 ( .A(n91845), .B(n91844), .Z(n91846) );
  IV U109532 ( .A(n91848), .Z(n91849) );
  NOR U109533 ( .A(n91850), .B(n91849), .Z(n91855) );
  IV U109534 ( .A(n91851), .Z(n91853) );
  NOR U109535 ( .A(n91853), .B(n91852), .Z(n91854) );
  XOR U109536 ( .A(n91857), .B(n91856), .Z(n91870) );
  IV U109537 ( .A(n91858), .Z(n91859) );
  NOR U109538 ( .A(n91860), .B(n91859), .Z(n91866) );
  NOR U109539 ( .A(n91862), .B(n91861), .Z(n91863) );
  NOR U109540 ( .A(n91864), .B(n91863), .Z(n91865) );
  NOR U109541 ( .A(n91866), .B(n91865), .Z(n91867) );
  XOR U109542 ( .A(n91868), .B(n91867), .Z(n91869) );
  XOR U109543 ( .A(n91870), .B(n91869), .Z(n91871) );
  XOR U109544 ( .A(n91872), .B(n91871), .Z(n91873) );
  XOR U109545 ( .A(n91874), .B(n91873), .Z(n91895) );
  IV U109546 ( .A(n91875), .Z(n91876) );
  NOR U109547 ( .A(n91877), .B(n91876), .Z(n91893) );
  IV U109548 ( .A(n91878), .Z(n91879) );
  NOR U109549 ( .A(n91880), .B(n91879), .Z(n91891) );
  IV U109550 ( .A(n91881), .Z(n91883) );
  NOR U109551 ( .A(n91883), .B(n91882), .Z(n91888) );
  IV U109552 ( .A(n91884), .Z(n91886) );
  NOR U109553 ( .A(n91886), .B(n91885), .Z(n91887) );
  NOR U109554 ( .A(n91888), .B(n91887), .Z(n91889) );
  IV U109555 ( .A(n91889), .Z(n91890) );
  NOR U109556 ( .A(n91891), .B(n91890), .Z(n91892) );
  XOR U109557 ( .A(n91893), .B(n91892), .Z(n91894) );
  XOR U109558 ( .A(n91895), .B(n91894), .Z(n91899) );
  XOR U109559 ( .A(n91896), .B(n91899), .Z(n91897) );
  NOR U109560 ( .A(n91898), .B(n91897), .Z(n91904) );
  IV U109561 ( .A(n91898), .Z(n91902) );
  XOR U109562 ( .A(n91900), .B(n91899), .Z(n91901) );
  NOR U109563 ( .A(n91902), .B(n91901), .Z(n91903) );
  NOR U109564 ( .A(n91904), .B(n91903), .Z(n91905) );
  XOR U109565 ( .A(n91906), .B(n91905), .Z(n91925) );
  NOR U109566 ( .A(n91908), .B(n91907), .Z(n91913) );
  IV U109567 ( .A(n91909), .Z(n91910) );
  NOR U109568 ( .A(n91911), .B(n91910), .Z(n91912) );
  NOR U109569 ( .A(n91913), .B(n91912), .Z(n91923) );
  IV U109570 ( .A(n91914), .Z(n91915) );
  NOR U109571 ( .A(n91916), .B(n91915), .Z(n91921) );
  IV U109572 ( .A(n91917), .Z(n91919) );
  NOR U109573 ( .A(n91919), .B(n91918), .Z(n91920) );
  NOR U109574 ( .A(n91921), .B(n91920), .Z(n91922) );
  XOR U109575 ( .A(n91923), .B(n91922), .Z(n91924) );
  XOR U109576 ( .A(n91925), .B(n91924), .Z(n91926) );
  XOR U109577 ( .A(n91927), .B(n91926), .Z(n91928) );
  XOR U109578 ( .A(n91929), .B(n91928), .Z(n91930) );
  XOR U109579 ( .A(n91931), .B(n91930), .Z(n91932) );
  XOR U109580 ( .A(n91933), .B(n91932), .Z(n91934) );
  XOR U109581 ( .A(n91935), .B(n91934), .Z(n91960) );
  IV U109582 ( .A(n91936), .Z(n91938) );
  NOR U109583 ( .A(n91938), .B(n91937), .Z(n91940) );
  NOR U109584 ( .A(n91940), .B(n91939), .Z(n91958) );
  IV U109585 ( .A(n91941), .Z(n91942) );
  NOR U109586 ( .A(n91943), .B(n91942), .Z(n91950) );
  IV U109587 ( .A(n91953), .Z(n91948) );
  NOR U109588 ( .A(n91945), .B(n91944), .Z(n91946) );
  IV U109589 ( .A(n91946), .Z(n91947) );
  NOR U109590 ( .A(n91948), .B(n91947), .Z(n91949) );
  NOR U109591 ( .A(n91950), .B(n91949), .Z(n91951) );
  IV U109592 ( .A(n91951), .Z(n91956) );
  IV U109593 ( .A(n91952), .Z(n91954) );
  NOR U109594 ( .A(n91954), .B(n91953), .Z(n91955) );
  NOR U109595 ( .A(n91956), .B(n91955), .Z(n91957) );
  XOR U109596 ( .A(n91958), .B(n91957), .Z(n91959) );
  XOR U109597 ( .A(n91960), .B(n91959), .Z(n91996) );
  NOR U109598 ( .A(n91962), .B(n91961), .Z(n91994) );
  IV U109599 ( .A(n91963), .Z(n91965) );
  NOR U109600 ( .A(n91965), .B(n91964), .Z(n91970) );
  IV U109601 ( .A(n91966), .Z(n91968) );
  NOR U109602 ( .A(n91968), .B(n91967), .Z(n91969) );
  NOR U109603 ( .A(n91970), .B(n91969), .Z(n91992) );
  NOR U109604 ( .A(n91972), .B(n91971), .Z(n91976) );
  IV U109605 ( .A(n91981), .Z(n91973) );
  NOR U109606 ( .A(n91974), .B(n91973), .Z(n91975) );
  NOR U109607 ( .A(n91976), .B(n91975), .Z(n91977) );
  IV U109608 ( .A(n91977), .Z(n91990) );
  IV U109609 ( .A(n91978), .Z(n91980) );
  NOR U109610 ( .A(n91980), .B(n91979), .Z(n91987) );
  NOR U109611 ( .A(n91982), .B(n91981), .Z(n91985) );
  IV U109612 ( .A(n91983), .Z(n91984) );
  NOR U109613 ( .A(n91985), .B(n91984), .Z(n91986) );
  NOR U109614 ( .A(n91987), .B(n91986), .Z(n91988) );
  IV U109615 ( .A(n91988), .Z(n91989) );
  NOR U109616 ( .A(n91990), .B(n91989), .Z(n91991) );
  XOR U109617 ( .A(n91992), .B(n91991), .Z(n91993) );
  XOR U109618 ( .A(n91994), .B(n91993), .Z(n91995) );
  XOR U109619 ( .A(n91996), .B(n91995), .Z(n91997) );
  XOR U109620 ( .A(n91998), .B(n91997), .Z(n92008) );
  IV U109621 ( .A(n91999), .Z(n92000) );
  NOR U109622 ( .A(n92001), .B(n92000), .Z(n92006) );
  IV U109623 ( .A(n92002), .Z(n92004) );
  NOR U109624 ( .A(n92004), .B(n92003), .Z(n92005) );
  NOR U109625 ( .A(n92006), .B(n92005), .Z(n92007) );
  XOR U109626 ( .A(n92008), .B(n92007), .Z(n92037) );
  IV U109627 ( .A(n92009), .Z(n92011) );
  NOR U109628 ( .A(n92011), .B(n92010), .Z(n92015) );
  NOR U109629 ( .A(n92013), .B(n92012), .Z(n92014) );
  NOR U109630 ( .A(n92015), .B(n92014), .Z(n92025) );
  IV U109631 ( .A(n92016), .Z(n92018) );
  NOR U109632 ( .A(n92018), .B(n92017), .Z(n92023) );
  IV U109633 ( .A(n92019), .Z(n92021) );
  NOR U109634 ( .A(n92021), .B(n92020), .Z(n92022) );
  NOR U109635 ( .A(n92023), .B(n92022), .Z(n92024) );
  XOR U109636 ( .A(n92025), .B(n92024), .Z(n92035) );
  IV U109637 ( .A(n92026), .Z(n92027) );
  NOR U109638 ( .A(n92028), .B(n92027), .Z(n92033) );
  IV U109639 ( .A(n92029), .Z(n92030) );
  NOR U109640 ( .A(n92031), .B(n92030), .Z(n92032) );
  NOR U109641 ( .A(n92033), .B(n92032), .Z(n92034) );
  XOR U109642 ( .A(n92035), .B(n92034), .Z(n92036) );
  XOR U109643 ( .A(n92037), .B(n92036), .Z(n92038) );
  XOR U109644 ( .A(n92039), .B(n92038), .Z(n92070) );
  IV U109645 ( .A(n92040), .Z(n92042) );
  NOR U109646 ( .A(n92042), .B(n92041), .Z(n92044) );
  NOR U109647 ( .A(n92044), .B(n92043), .Z(n92058) );
  NOR U109648 ( .A(n92046), .B(n92045), .Z(n92056) );
  XOR U109649 ( .A(n92049), .B(n92050), .Z(n92048) );
  NOR U109650 ( .A(n92048), .B(n92047), .Z(n92053) );
  IV U109651 ( .A(n92049), .Z(n92051) );
  NOR U109652 ( .A(n92051), .B(n92050), .Z(n92052) );
  NOR U109653 ( .A(n92053), .B(n92052), .Z(n92054) );
  IV U109654 ( .A(n92054), .Z(n92055) );
  NOR U109655 ( .A(n92056), .B(n92055), .Z(n92057) );
  XOR U109656 ( .A(n92058), .B(n92057), .Z(n92068) );
  NOR U109657 ( .A(n92060), .B(n92059), .Z(n92066) );
  NOR U109658 ( .A(n92062), .B(n92061), .Z(n92063) );
  NOR U109659 ( .A(n92064), .B(n92063), .Z(n92065) );
  NOR U109660 ( .A(n92066), .B(n92065), .Z(n92067) );
  XOR U109661 ( .A(n92068), .B(n92067), .Z(n92069) );
  XOR U109662 ( .A(n92070), .B(n92069), .Z(n92071) );
  XOR U109663 ( .A(n92072), .B(n92071), .Z(n92098) );
  IV U109664 ( .A(n92073), .Z(n92074) );
  NOR U109665 ( .A(n92074), .B(n92091), .Z(n92075) );
  NOR U109666 ( .A(n92076), .B(n92075), .Z(n92086) );
  IV U109667 ( .A(n92077), .Z(n92079) );
  NOR U109668 ( .A(n92079), .B(n92078), .Z(n92084) );
  IV U109669 ( .A(n92080), .Z(n92082) );
  NOR U109670 ( .A(n92082), .B(n92081), .Z(n92083) );
  NOR U109671 ( .A(n92084), .B(n92083), .Z(n92085) );
  XOR U109672 ( .A(n92086), .B(n92085), .Z(n92096) );
  IV U109673 ( .A(n92087), .Z(n92089) );
  NOR U109674 ( .A(n92089), .B(n92088), .Z(n92094) );
  IV U109675 ( .A(n92090), .Z(n92092) );
  NOR U109676 ( .A(n92092), .B(n92091), .Z(n92093) );
  NOR U109677 ( .A(n92094), .B(n92093), .Z(n92095) );
  XOR U109678 ( .A(n92096), .B(n92095), .Z(n92097) );
  XOR U109679 ( .A(n92098), .B(n92097), .Z(n92099) );
  XOR U109680 ( .A(n92100), .B(n92099), .Z(n92101) );
  IV U109681 ( .A(n92101), .Z(n92321) );
  XOR U109682 ( .A(n92103), .B(n92102), .Z(n92155) );
  NOR U109683 ( .A(n92105), .B(n92104), .Z(n92107) );
  XOR U109684 ( .A(n92107), .B(n92106), .Z(n92198) );
  XOR U109685 ( .A(n92109), .B(n92108), .Z(n92196) );
  NOR U109686 ( .A(n92198), .B(n92196), .Z(n92110) );
  IV U109687 ( .A(n92110), .Z(n92154) );
  NOR U109688 ( .A(n92112), .B(n92111), .Z(n92114) );
  XOR U109689 ( .A(n92114), .B(n92113), .Z(n92140) );
  NOR U109690 ( .A(n92116), .B(n92115), .Z(n92135) );
  XOR U109691 ( .A(n92135), .B(n92117), .Z(n92188) );
  NOR U109692 ( .A(n92119), .B(n92118), .Z(n92120) );
  XOR U109693 ( .A(n92121), .B(n92120), .Z(n92144) );
  IV U109694 ( .A(n92122), .Z(n92124) );
  NOR U109695 ( .A(n92124), .B(n92123), .Z(n92141) );
  IV U109696 ( .A(n92141), .Z(n92125) );
  NOR U109697 ( .A(n92144), .B(n92125), .Z(n92126) );
  IV U109698 ( .A(n92126), .Z(n92189) );
  NOR U109699 ( .A(n92188), .B(n92189), .Z(n92137) );
  IV U109700 ( .A(n92137), .Z(n92127) );
  NOR U109701 ( .A(n92140), .B(n92127), .Z(n92166) );
  IV U109702 ( .A(n92166), .Z(n92128) );
  NOR U109703 ( .A(n92154), .B(n92128), .Z(n92156) );
  IV U109704 ( .A(n92156), .Z(n92129) );
  NOR U109705 ( .A(n92155), .B(n92129), .Z(n92130) );
  IV U109706 ( .A(n92130), .Z(n92175) );
  NOR U109707 ( .A(n92132), .B(n92131), .Z(n92133) );
  XOR U109708 ( .A(n92134), .B(n92133), .Z(n92174) );
  XOR U109709 ( .A(n92175), .B(n92174), .Z(n92206) );
  NOR U109710 ( .A(n92136), .B(n92135), .Z(n92138) );
  NOR U109711 ( .A(n92138), .B(n92137), .Z(n92139) );
  XOR U109712 ( .A(n92140), .B(n92139), .Z(n92163) );
  IV U109713 ( .A(n92163), .Z(n92152) );
  NOR U109714 ( .A(n92142), .B(n92141), .Z(n92143) );
  XOR U109715 ( .A(n92144), .B(n92143), .Z(n92145) );
  IV U109716 ( .A(n92145), .Z(n92212) );
  NOR U109717 ( .A(n92212), .B(n92188), .Z(n92146) );
  IV U109718 ( .A(n92146), .Z(n92161) );
  IV U109719 ( .A(n92147), .Z(n92149) );
  NOR U109720 ( .A(n92149), .B(n92148), .Z(n92183) );
  IV U109721 ( .A(n92183), .Z(n92150) );
  NOR U109722 ( .A(n92161), .B(n92150), .Z(n92151) );
  IV U109723 ( .A(n92151), .Z(n92162) );
  NOR U109724 ( .A(n92152), .B(n92162), .Z(n92165) );
  IV U109725 ( .A(n92165), .Z(n92153) );
  NOR U109726 ( .A(n92154), .B(n92153), .Z(n92177) );
  XOR U109727 ( .A(n92156), .B(n92155), .Z(n92179) );
  XOR U109728 ( .A(n92177), .B(n92179), .Z(n92262) );
  IV U109729 ( .A(n92157), .Z(n92159) );
  NOR U109730 ( .A(n92159), .B(n92158), .Z(n92182) );
  IV U109731 ( .A(n92182), .Z(n92160) );
  NOR U109732 ( .A(n92161), .B(n92160), .Z(n92193) );
  IV U109733 ( .A(n92193), .Z(n92164) );
  XOR U109734 ( .A(n92163), .B(n92162), .Z(n92192) );
  NOR U109735 ( .A(n92164), .B(n92192), .Z(n92181) );
  IV U109736 ( .A(n92181), .Z(n92168) );
  IV U109737 ( .A(n92196), .Z(n92167) );
  NOR U109738 ( .A(n92166), .B(n92165), .Z(n92197) );
  XOR U109739 ( .A(n92167), .B(n92197), .Z(n92226) );
  NOR U109740 ( .A(n92168), .B(n92226), .Z(n92209) );
  IV U109741 ( .A(n92209), .Z(n92169) );
  NOR U109742 ( .A(n92262), .B(n92169), .Z(n92170) );
  IV U109743 ( .A(n92170), .Z(n92171) );
  NOR U109744 ( .A(n92198), .B(n92171), .Z(n92203) );
  IV U109745 ( .A(n92203), .Z(n92172) );
  NOR U109746 ( .A(n92206), .B(n92172), .Z(n92236) );
  XOR U109747 ( .A(n92242), .B(n92173), .Z(n92296) );
  IV U109748 ( .A(n92174), .Z(n92176) );
  NOR U109749 ( .A(n92176), .B(n92175), .Z(n92244) );
  IV U109750 ( .A(n92177), .Z(n92178) );
  NOR U109751 ( .A(n92179), .B(n92178), .Z(n92204) );
  IV U109752 ( .A(n92204), .Z(n92180) );
  NOR U109753 ( .A(n92206), .B(n92180), .Z(n92243) );
  NOR U109754 ( .A(n92244), .B(n92243), .Z(n92297) );
  XOR U109755 ( .A(n92296), .B(n92297), .Z(n92237) );
  XOR U109756 ( .A(n92236), .B(n92237), .Z(n92344) );
  IV U109757 ( .A(n92344), .Z(n92286) );
  XOR U109758 ( .A(n92181), .B(n92226), .Z(n92266) );
  NOR U109759 ( .A(n92183), .B(n92182), .Z(n92211) );
  XOR U109760 ( .A(n92211), .B(n92212), .Z(n92270) );
  IV U109761 ( .A(n92270), .Z(n92221) );
  IV U109762 ( .A(n92184), .Z(n92186) );
  NOR U109763 ( .A(n92186), .B(n92185), .Z(n92268) );
  IV U109764 ( .A(n92268), .Z(n92187) );
  NOR U109765 ( .A(n92221), .B(n92187), .Z(n92213) );
  IV U109766 ( .A(n92213), .Z(n92191) );
  XOR U109767 ( .A(n92189), .B(n92188), .Z(n92216) );
  IV U109768 ( .A(n92216), .Z(n92190) );
  NOR U109769 ( .A(n92191), .B(n92190), .Z(n92275) );
  IV U109770 ( .A(n92275), .Z(n92194) );
  XOR U109771 ( .A(n92193), .B(n92192), .Z(n92274) );
  NOR U109772 ( .A(n92194), .B(n92274), .Z(n92264) );
  IV U109773 ( .A(n92264), .Z(n92195) );
  NOR U109774 ( .A(n92266), .B(n92195), .Z(n92208) );
  IV U109775 ( .A(n92208), .Z(n92200) );
  NOR U109776 ( .A(n92197), .B(n92196), .Z(n92199) );
  XOR U109777 ( .A(n92199), .B(n92198), .Z(n92257) );
  NOR U109778 ( .A(n92200), .B(n92257), .Z(n92201) );
  IV U109779 ( .A(n92201), .Z(n92202) );
  NOR U109780 ( .A(n92262), .B(n92202), .Z(n92254) );
  IV U109781 ( .A(n92254), .Z(n92207) );
  NOR U109782 ( .A(n92204), .B(n92203), .Z(n92205) );
  XOR U109783 ( .A(n92206), .B(n92205), .Z(n92256) );
  IV U109784 ( .A(n92256), .Z(n92230) );
  NOR U109785 ( .A(n92207), .B(n92230), .Z(n92231) );
  IV U109786 ( .A(n92231), .Z(n92343) );
  NOR U109787 ( .A(n92286), .B(n92343), .Z(n92235) );
  NOR U109788 ( .A(n92209), .B(n92208), .Z(n92258) );
  XOR U109789 ( .A(n92257), .B(n92258), .Z(n92210) );
  IV U109790 ( .A(n92210), .Z(n92335) );
  NOR U109791 ( .A(n92212), .B(n92211), .Z(n92214) );
  NOR U109792 ( .A(n92214), .B(n92213), .Z(n92215) );
  XOR U109793 ( .A(n92216), .B(n92215), .Z(n92328) );
  IV U109794 ( .A(n92217), .Z(n92219) );
  NOR U109795 ( .A(n92219), .B(n92218), .Z(n92267) );
  IV U109796 ( .A(n92267), .Z(n92220) );
  NOR U109797 ( .A(n92221), .B(n92220), .Z(n92325) );
  IV U109798 ( .A(n92325), .Z(n92222) );
  NOR U109799 ( .A(n92328), .B(n92222), .Z(n92223) );
  IV U109800 ( .A(n92223), .Z(n92224) );
  NOR U109801 ( .A(n92274), .B(n92224), .Z(n92263) );
  IV U109802 ( .A(n92263), .Z(n92225) );
  NOR U109803 ( .A(n92226), .B(n92225), .Z(n92334) );
  IV U109804 ( .A(n92334), .Z(n92227) );
  NOR U109805 ( .A(n92335), .B(n92227), .Z(n92259) );
  IV U109806 ( .A(n92259), .Z(n92228) );
  NOR U109807 ( .A(n92262), .B(n92228), .Z(n92253) );
  IV U109808 ( .A(n92253), .Z(n92229) );
  NOR U109809 ( .A(n92230), .B(n92229), .Z(n92342) );
  IV U109810 ( .A(n92342), .Z(n92233) );
  NOR U109811 ( .A(n92344), .B(n92231), .Z(n92232) );
  NOR U109812 ( .A(n92233), .B(n92232), .Z(n92234) );
  NOR U109813 ( .A(n92235), .B(n92234), .Z(n92289) );
  IV U109814 ( .A(n92236), .Z(n92239) );
  IV U109815 ( .A(n92237), .Z(n92238) );
  NOR U109816 ( .A(n92239), .B(n92238), .Z(n92240) );
  IV U109817 ( .A(n92240), .Z(n92295) );
  NOR U109818 ( .A(n92242), .B(n92241), .Z(n92248) );
  XOR U109819 ( .A(n92244), .B(n92243), .Z(n92245) );
  NOR U109820 ( .A(n92246), .B(n92245), .Z(n92247) );
  NOR U109821 ( .A(n92248), .B(n92247), .Z(n92249) );
  XOR U109822 ( .A(n92250), .B(n92249), .Z(n92251) );
  XOR U109823 ( .A(n92252), .B(n92251), .Z(n92300) );
  XOR U109824 ( .A(n92295), .B(n92300), .Z(n92288) );
  NOR U109825 ( .A(n92289), .B(n92288), .Z(n92292) );
  NOR U109826 ( .A(n92254), .B(n92253), .Z(n92255) );
  XOR U109827 ( .A(n92256), .B(n92255), .Z(n92340) );
  NOR U109828 ( .A(n92258), .B(n92257), .Z(n92260) );
  NOR U109829 ( .A(n92260), .B(n92259), .Z(n92261) );
  XOR U109830 ( .A(n92262), .B(n92261), .Z(n92338) );
  IV U109831 ( .A(n92338), .Z(n92283) );
  NOR U109832 ( .A(n92264), .B(n92263), .Z(n92265) );
  XOR U109833 ( .A(n92266), .B(n92265), .Z(n92332) );
  IV U109834 ( .A(n92332), .Z(n92280) );
  NOR U109835 ( .A(n92268), .B(n92267), .Z(n92269) );
  XOR U109836 ( .A(n92270), .B(n92269), .Z(n92323) );
  NOR U109837 ( .A(n92272), .B(n92271), .Z(n92273) );
  IV U109838 ( .A(n92273), .Z(n92322) );
  NOR U109839 ( .A(n92323), .B(n92322), .Z(n92324) );
  IV U109840 ( .A(n92324), .Z(n92276) );
  XOR U109841 ( .A(n92275), .B(n92274), .Z(n92326) );
  NOR U109842 ( .A(n92276), .B(n92326), .Z(n92277) );
  IV U109843 ( .A(n92277), .Z(n92278) );
  NOR U109844 ( .A(n92328), .B(n92278), .Z(n92331) );
  IV U109845 ( .A(n92331), .Z(n92279) );
  NOR U109846 ( .A(n92280), .B(n92279), .Z(n92333) );
  IV U109847 ( .A(n92333), .Z(n92281) );
  NOR U109848 ( .A(n92335), .B(n92281), .Z(n92337) );
  IV U109849 ( .A(n92337), .Z(n92282) );
  NOR U109850 ( .A(n92283), .B(n92282), .Z(n92284) );
  IV U109851 ( .A(n92284), .Z(n92339) );
  NOR U109852 ( .A(n92340), .B(n92339), .Z(n92341) );
  IV U109853 ( .A(n92341), .Z(n92285) );
  NOR U109854 ( .A(n92286), .B(n92285), .Z(n92287) );
  IV U109855 ( .A(n92287), .Z(n92348) );
  XOR U109856 ( .A(n92289), .B(n92288), .Z(n92290) );
  IV U109857 ( .A(n92290), .Z(n92347) );
  NOR U109858 ( .A(n92348), .B(n92347), .Z(n92291) );
  NOR U109859 ( .A(n92292), .B(n92291), .Z(n92293) );
  IV U109860 ( .A(n92293), .Z(n92305) );
  IV U109861 ( .A(n92300), .Z(n92294) );
  NOR U109862 ( .A(n92295), .B(n92294), .Z(n92302) );
  NOR U109863 ( .A(n92297), .B(n92296), .Z(n92298) );
  IV U109864 ( .A(n92298), .Z(n92299) );
  NOR U109865 ( .A(n92300), .B(n92299), .Z(n92301) );
  NOR U109866 ( .A(n92302), .B(n92301), .Z(n92303) );
  IV U109867 ( .A(n92303), .Z(n92304) );
  NOR U109868 ( .A(n92305), .B(n92304), .Z(n92319) );
  NOR U109869 ( .A(n92307), .B(n92306), .Z(n92317) );
  IV U109870 ( .A(n92308), .Z(n92310) );
  NOR U109871 ( .A(n92310), .B(n92309), .Z(n92314) );
  NOR U109872 ( .A(n92312), .B(n92311), .Z(n92313) );
  NOR U109873 ( .A(n92314), .B(n92313), .Z(n92315) );
  IV U109874 ( .A(n92315), .Z(n92316) );
  NOR U109875 ( .A(n92317), .B(n92316), .Z(n92318) );
  XOR U109876 ( .A(n92319), .B(n92318), .Z(n92320) );
  XOR U109877 ( .A(n92321), .B(n92320), .Z(o[10]) );
  XOR U109878 ( .A(n92323), .B(n92322), .Z(o[1]) );
  NOR U109879 ( .A(n92325), .B(n92324), .Z(n92327) );
  XOR U109880 ( .A(n92328), .B(n92327), .Z(o[2]) );
  IV U109881 ( .A(n92326), .Z(n92330) );
  NOR U109882 ( .A(n92328), .B(n92327), .Z(n92329) );
  XOR U109883 ( .A(n92330), .B(n92329), .Z(o[3]) );
  XOR U109884 ( .A(n92332), .B(n92331), .Z(o[4]) );
  NOR U109885 ( .A(n92334), .B(n92333), .Z(n92336) );
  XOR U109886 ( .A(n92336), .B(n92335), .Z(o[5]) );
  XOR U109887 ( .A(n92338), .B(n92337), .Z(o[6]) );
  XOR U109888 ( .A(n92340), .B(n92339), .Z(o[7]) );
  NOR U109889 ( .A(n92342), .B(n92341), .Z(n92346) );
  XOR U109890 ( .A(n92344), .B(n92343), .Z(n92345) );
  XOR U109891 ( .A(n92346), .B(n92345), .Z(o[8]) );
  XOR U109892 ( .A(n92348), .B(n92347), .Z(o[9]) );
endmodule

