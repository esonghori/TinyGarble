
module hamming_N32_CC1 ( clk, rst, g_input, e_input, o );
  input [31:0] g_input;
  input [31:0] e_input;
  output [5:0] o;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146;

  MUX U33 ( .IN0(n100), .IN1(n98), .SEL(n99), .F(n94) );
  MUX U34 ( .IN0(n33), .IN1(n36), .SEL(n34), .F(n26) );
  XOR U35 ( .A(n57), .B(n56), .Z(n41) );
  MUX U36 ( .IN0(n97), .IN1(n95), .SEL(n96), .F(n1) );
  IV U37 ( .A(n1), .Z(n50) );
  MUX U38 ( .IN0(n108), .IN1(n106), .SEL(n107), .F(n2) );
  IV U39 ( .A(n2), .Z(n55) );
  MUX U40 ( .IN0(n78), .IN1(n76), .SEL(n77), .F(n70) );
  XNOR U41 ( .A(n43), .B(n44), .Z(n24) );
  XOR U42 ( .A(n30), .B(n29), .Z(n23) );
  MUX U43 ( .IN0(n112), .IN1(n110), .SEL(n111), .F(n3) );
  IV U44 ( .A(n3), .Z(n62) );
  MUX U45 ( .IN0(n120), .IN1(n118), .SEL(n119), .F(n4) );
  IV U46 ( .A(n4), .Z(n66) );
  MUX U47 ( .IN0(n88), .IN1(n86), .SEL(n87), .F(n51) );
  XOR U48 ( .A(n36), .B(n34), .Z(n47) );
  MUX U49 ( .IN0(n55), .IN1(n5), .SEL(n56), .F(n28) );
  IV U50 ( .A(n57), .Z(n5) );
  MUX U51 ( .IN0(n21), .IN1(n6), .SEL(n22), .F(n12) );
  IV U52 ( .A(n23), .Z(n6) );
  MUX U53 ( .IN0(n105), .IN1(n103), .SEL(n104), .F(n63) );
  MUX U54 ( .IN0(n7), .IN1(n79), .SEL(n80), .F(n36) );
  IV U55 ( .A(n81), .Z(n7) );
  MUX U56 ( .IN0(n8), .IN1(n84), .SEL(n83), .F(n37) );
  IV U57 ( .A(n82), .Z(n8) );
  MUX U58 ( .IN0(n48), .IN1(n51), .SEL(n49), .F(n42) );
  MUX U59 ( .IN0(n28), .IN1(n9), .SEL(n29), .F(n16) );
  IV U60 ( .A(n30), .Z(n9) );
  MUX U61 ( .IN0(n115), .IN1(n113), .SEL(n114), .F(n109) );
  MUX U62 ( .IN0(n64), .IN1(n67), .SEL(n65), .F(n30) );
  MUX U63 ( .IN0(n24), .IN1(n26), .SEL(n25), .F(n19) );
  NOR U64 ( .A(o[4]), .B(n10), .Z(o[5]) );
  XNOR U65 ( .A(n11), .B(n12), .Z(o[4]) );
  XOR U66 ( .A(n10), .B(n13), .Z(n11) );
  AND U67 ( .A(n14), .B(n15), .Z(n13) );
  XOR U68 ( .A(n16), .B(n12), .Z(n15) );
  OR U69 ( .A(n17), .B(o[3]), .Z(n10) );
  XNOR U70 ( .A(n18), .B(n14), .Z(o[3]) );
  XOR U71 ( .A(n19), .B(n20), .Z(n14) );
  IV U72 ( .A(n12), .Z(n20) );
  XOR U73 ( .A(n16), .B(n17), .Z(n18) );
  OR U74 ( .A(n27), .B(o[2]), .Z(n17) );
  XNOR U75 ( .A(n31), .B(n22), .Z(o[2]) );
  XOR U76 ( .A(n32), .B(n26), .Z(n22) );
  XNOR U77 ( .A(n25), .B(n21), .Z(n32) );
  XOR U78 ( .A(n37), .B(n38), .Z(n21) );
  AND U79 ( .A(n39), .B(n40), .Z(n38) );
  XNOR U80 ( .A(n41), .B(n37), .Z(n40) );
  XOR U81 ( .A(n42), .B(n24), .Z(n25) );
  AND U82 ( .A(n45), .B(n46), .Z(n44) );
  XNOR U83 ( .A(n43), .B(n47), .Z(n46) );
  XNOR U84 ( .A(n23), .B(n27), .Z(n31) );
  OR U85 ( .A(n52), .B(o[1]), .Z(n27) );
  XOR U86 ( .A(n53), .B(n54), .Z(n29) );
  IV U87 ( .A(n28), .Z(n54) );
  XOR U88 ( .A(n58), .B(n59), .Z(n53) );
  AND U89 ( .A(n60), .B(n61), .Z(n59) );
  XNOR U90 ( .A(n62), .B(n63), .Z(n61) );
  XNOR U91 ( .A(n68), .B(n39), .Z(o[1]) );
  XOR U92 ( .A(n69), .B(n47), .Z(n39) );
  XOR U93 ( .A(n70), .B(n33), .Z(n34) );
  IV U94 ( .A(n35), .Z(n33) );
  XNOR U95 ( .A(n71), .B(n72), .Z(n35) );
  ANDN U96 ( .A(n73), .B(n74), .Z(n72) );
  XOR U97 ( .A(n71), .B(n75), .Z(n73) );
  XNOR U98 ( .A(n45), .B(n37), .Z(n69) );
  XOR U99 ( .A(n85), .B(n51), .Z(n45) );
  XNOR U100 ( .A(n49), .B(n43), .Z(n85) );
  XNOR U101 ( .A(n89), .B(n90), .Z(n43) );
  ANDN U102 ( .A(n91), .B(n92), .Z(n90) );
  XOR U103 ( .A(n89), .B(n93), .Z(n91) );
  XOR U104 ( .A(n94), .B(n48), .Z(n49) );
  IV U105 ( .A(n50), .Z(n48) );
  XNOR U106 ( .A(n41), .B(n52), .Z(n68) );
  OR U107 ( .A(n101), .B(o[0]), .Z(n52) );
  XOR U108 ( .A(n102), .B(n63), .Z(n56) );
  XNOR U109 ( .A(n60), .B(n55), .Z(n102) );
  XOR U110 ( .A(n109), .B(n58), .Z(n60) );
  IV U111 ( .A(n62), .Z(n58) );
  XNOR U112 ( .A(n67), .B(n116), .Z(n57) );
  IV U113 ( .A(n65), .Z(n116) );
  XOR U114 ( .A(n117), .B(n64), .Z(n65) );
  IV U115 ( .A(n66), .Z(n64) );
  XOR U116 ( .A(n121), .B(n122), .Z(n117) );
  ANDN U117 ( .A(n123), .B(n124), .Z(n122) );
  XOR U118 ( .A(n121), .B(n125), .Z(n123) );
  XOR U119 ( .A(n126), .B(n127), .Z(n67) );
  ANDN U120 ( .A(n128), .B(n129), .Z(n127) );
  XNOR U121 ( .A(n126), .B(n130), .Z(n128) );
  XNOR U122 ( .A(n131), .B(n83), .Z(o[0]) );
  XOR U123 ( .A(n132), .B(n93), .Z(n83) );
  XNOR U124 ( .A(n75), .B(n74), .Z(n93) );
  XNOR U125 ( .A(n133), .B(n78), .Z(n74) );
  XNOR U126 ( .A(g_input[24]), .B(e_input[24]), .Z(n78) );
  XNOR U127 ( .A(n77), .B(n71), .Z(n133) );
  XNOR U128 ( .A(g_input[18]), .B(e_input[18]), .Z(n71) );
  XNOR U129 ( .A(n134), .B(n76), .Z(n77) );
  XNOR U130 ( .A(g_input[22]), .B(e_input[22]), .Z(n76) );
  XNOR U131 ( .A(g_input[23]), .B(e_input[23]), .Z(n134) );
  XOR U132 ( .A(n81), .B(n80), .Z(n75) );
  XNOR U133 ( .A(n135), .B(n79), .Z(n80) );
  XNOR U134 ( .A(g_input[19]), .B(e_input[19]), .Z(n79) );
  XNOR U135 ( .A(g_input[20]), .B(e_input[20]), .Z(n135) );
  XOR U136 ( .A(g_input[21]), .B(e_input[21]), .Z(n81) );
  XNOR U137 ( .A(n92), .B(n82), .Z(n132) );
  XNOR U138 ( .A(g_input[1]), .B(e_input[1]), .Z(n82) );
  XNOR U139 ( .A(n136), .B(n97), .Z(n92) );
  XNOR U140 ( .A(n88), .B(n87), .Z(n97) );
  XNOR U141 ( .A(n137), .B(n86), .Z(n87) );
  XNOR U142 ( .A(g_input[26]), .B(e_input[26]), .Z(n86) );
  XNOR U143 ( .A(g_input[27]), .B(e_input[27]), .Z(n137) );
  XNOR U144 ( .A(g_input[28]), .B(e_input[28]), .Z(n88) );
  XNOR U145 ( .A(n96), .B(n89), .Z(n136) );
  XNOR U146 ( .A(g_input[17]), .B(e_input[17]), .Z(n89) );
  XNOR U147 ( .A(n138), .B(n100), .Z(n96) );
  XNOR U148 ( .A(g_input[31]), .B(e_input[31]), .Z(n100) );
  XNOR U149 ( .A(n99), .B(n95), .Z(n138) );
  XNOR U150 ( .A(g_input[25]), .B(e_input[25]), .Z(n95) );
  XNOR U151 ( .A(n139), .B(n98), .Z(n99) );
  XNOR U152 ( .A(g_input[29]), .B(e_input[29]), .Z(n98) );
  XNOR U153 ( .A(g_input[30]), .B(e_input[30]), .Z(n139) );
  XOR U154 ( .A(n101), .B(n84), .Z(n131) );
  XOR U155 ( .A(n108), .B(n107), .Z(n84) );
  XNOR U156 ( .A(n140), .B(n112), .Z(n107) );
  XNOR U157 ( .A(n105), .B(n104), .Z(n112) );
  XNOR U158 ( .A(n141), .B(n103), .Z(n104) );
  XNOR U159 ( .A(g_input[11]), .B(e_input[11]), .Z(n103) );
  XNOR U160 ( .A(g_input[12]), .B(e_input[12]), .Z(n141) );
  XNOR U161 ( .A(g_input[13]), .B(e_input[13]), .Z(n105) );
  XNOR U162 ( .A(n111), .B(n106), .Z(n140) );
  XNOR U163 ( .A(g_input[2]), .B(e_input[2]), .Z(n106) );
  XNOR U164 ( .A(n142), .B(n115), .Z(n111) );
  XNOR U165 ( .A(g_input[16]), .B(e_input[16]), .Z(n115) );
  XNOR U166 ( .A(n114), .B(n110), .Z(n142) );
  XNOR U167 ( .A(g_input[10]), .B(e_input[10]), .Z(n110) );
  XNOR U168 ( .A(n143), .B(n113), .Z(n114) );
  XNOR U169 ( .A(g_input[14]), .B(e_input[14]), .Z(n113) );
  XNOR U170 ( .A(g_input[15]), .B(e_input[15]), .Z(n143) );
  XNOR U171 ( .A(n120), .B(n119), .Z(n108) );
  XNOR U172 ( .A(n144), .B(n125), .Z(n119) );
  XNOR U173 ( .A(g_input[9]), .B(e_input[9]), .Z(n125) );
  XNOR U174 ( .A(n124), .B(n118), .Z(n144) );
  XNOR U175 ( .A(g_input[3]), .B(e_input[3]), .Z(n118) );
  XNOR U176 ( .A(n145), .B(n121), .Z(n124) );
  XNOR U177 ( .A(g_input[7]), .B(e_input[7]), .Z(n121) );
  XNOR U178 ( .A(g_input[8]), .B(e_input[8]), .Z(n145) );
  XOR U179 ( .A(n130), .B(n129), .Z(n120) );
  XNOR U180 ( .A(n146), .B(n126), .Z(n129) );
  XNOR U181 ( .A(g_input[4]), .B(e_input[4]), .Z(n126) );
  XNOR U182 ( .A(g_input[5]), .B(e_input[5]), .Z(n146) );
  XOR U183 ( .A(g_input[6]), .B(e_input[6]), .Z(n130) );
  XNOR U184 ( .A(g_input[0]), .B(e_input[0]), .Z(n101) );
endmodule

