
module mult_N256_CC8 ( clk, rst, a, b, c );
  input [255:0] a;
  input [31:0] b;
  output [511:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
         n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
         n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
         n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
         n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345,
         n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
         n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
         n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369,
         n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377,
         n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
         n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
         n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401,
         n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409,
         n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417,
         n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425,
         n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
         n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441,
         n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
         n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
         n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465,
         n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473,
         n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
         n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489,
         n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
         n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
         n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
         n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521,
         n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
         n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537,
         n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545,
         n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553,
         n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561,
         n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569,
         n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
         n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585,
         n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593,
         n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601,
         n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609,
         n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617,
         n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625,
         n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633,
         n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
         n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
         n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657,
         n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665,
         n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673,
         n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681,
         n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689,
         n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697,
         n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705,
         n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713,
         n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721,
         n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729,
         n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737,
         n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745,
         n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753,
         n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761,
         n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769,
         n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777,
         n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785,
         n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793,
         n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801,
         n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809,
         n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817,
         n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825,
         n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833,
         n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841,
         n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849,
         n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857,
         n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865,
         n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873,
         n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881,
         n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889,
         n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897,
         n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905,
         n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913,
         n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921,
         n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929,
         n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937,
         n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945,
         n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953,
         n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961,
         n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969,
         n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977,
         n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985,
         n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993,
         n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001,
         n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009,
         n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017,
         n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025,
         n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033,
         n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041,
         n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049,
         n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057,
         n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065,
         n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073,
         n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081,
         n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089,
         n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097,
         n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
         n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113,
         n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121,
         n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129,
         n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137,
         n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145,
         n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153,
         n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161,
         n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169,
         n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177,
         n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185,
         n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193,
         n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201,
         n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209,
         n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217,
         n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225,
         n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233,
         n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241,
         n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249,
         n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257,
         n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265,
         n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273,
         n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281,
         n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289,
         n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297,
         n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305,
         n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313,
         n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321,
         n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329,
         n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337,
         n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345,
         n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353,
         n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361,
         n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369,
         n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377,
         n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385,
         n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393,
         n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401,
         n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409,
         n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417,
         n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425,
         n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433,
         n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441,
         n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449,
         n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457,
         n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465,
         n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473,
         n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481,
         n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489,
         n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497,
         n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505,
         n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513,
         n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521,
         n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529,
         n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537,
         n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545,
         n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553,
         n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561,
         n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569,
         n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577,
         n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585,
         n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593,
         n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601,
         n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609,
         n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617,
         n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625,
         n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633,
         n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641,
         n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649,
         n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657,
         n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665,
         n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673,
         n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681,
         n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689,
         n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697,
         n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705,
         n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713,
         n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721,
         n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729,
         n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737,
         n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745,
         n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753,
         n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761,
         n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769,
         n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777,
         n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785,
         n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793,
         n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801,
         n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809,
         n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817,
         n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825,
         n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833,
         n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841,
         n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849,
         n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857,
         n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865,
         n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873,
         n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881,
         n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889,
         n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897,
         n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905,
         n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913,
         n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921,
         n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929,
         n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937,
         n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945,
         n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953,
         n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961,
         n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969,
         n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977,
         n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985,
         n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993,
         n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001,
         n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009,
         n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017,
         n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025,
         n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033,
         n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041,
         n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049,
         n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057,
         n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065,
         n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073,
         n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081,
         n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089,
         n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097,
         n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105,
         n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113,
         n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121,
         n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129,
         n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137,
         n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145,
         n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153,
         n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161,
         n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169,
         n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177,
         n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185,
         n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193,
         n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201,
         n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209,
         n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217,
         n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225,
         n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233,
         n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241,
         n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249,
         n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257,
         n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265,
         n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273,
         n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281,
         n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289,
         n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297,
         n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305,
         n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313,
         n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321,
         n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329,
         n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337,
         n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345,
         n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353,
         n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361,
         n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369,
         n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377,
         n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385,
         n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393,
         n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401,
         n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409,
         n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417,
         n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425,
         n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433,
         n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441,
         n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449,
         n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457,
         n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465,
         n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473,
         n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481,
         n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489,
         n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497,
         n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505,
         n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513,
         n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521,
         n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529,
         n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537,
         n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545,
         n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553,
         n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561,
         n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569,
         n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577,
         n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585,
         n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593,
         n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601,
         n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609,
         n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617,
         n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625,
         n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633,
         n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641,
         n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649,
         n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657,
         n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665,
         n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673,
         n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681,
         n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689,
         n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697,
         n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705,
         n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713,
         n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721,
         n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729,
         n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737,
         n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745,
         n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753,
         n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761,
         n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769,
         n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777,
         n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785,
         n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793,
         n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801,
         n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809,
         n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817,
         n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825,
         n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833,
         n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841,
         n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849,
         n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857,
         n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865,
         n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873,
         n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881,
         n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889,
         n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897,
         n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905,
         n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913,
         n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921,
         n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929,
         n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937,
         n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945,
         n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953,
         n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961,
         n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969,
         n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977,
         n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985,
         n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993,
         n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001,
         n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009,
         n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017,
         n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025,
         n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033,
         n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041,
         n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049,
         n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057,
         n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065,
         n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073,
         n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081,
         n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089,
         n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097,
         n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105,
         n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113,
         n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121,
         n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129,
         n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137,
         n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145,
         n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153,
         n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161,
         n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169,
         n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177,
         n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185,
         n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193,
         n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201,
         n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209,
         n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217,
         n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225,
         n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233,
         n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241,
         n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249,
         n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257,
         n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265,
         n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273,
         n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281,
         n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289,
         n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297,
         n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305,
         n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313,
         n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321,
         n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329,
         n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337,
         n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345,
         n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353,
         n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361,
         n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369,
         n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377,
         n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385,
         n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393,
         n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401,
         n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409,
         n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417,
         n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425,
         n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433,
         n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441,
         n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449,
         n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457,
         n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465,
         n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473,
         n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481,
         n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489,
         n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497,
         n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505,
         n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513,
         n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521,
         n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529,
         n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537,
         n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545,
         n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553,
         n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561,
         n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569,
         n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577,
         n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585,
         n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593,
         n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601,
         n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609,
         n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617,
         n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625,
         n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633,
         n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641,
         n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649,
         n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657,
         n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665,
         n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673,
         n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681,
         n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689,
         n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697,
         n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705,
         n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713,
         n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721,
         n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729,
         n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737,
         n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745,
         n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753,
         n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761,
         n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769,
         n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777,
         n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785,
         n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793,
         n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801,
         n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809,
         n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817,
         n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825,
         n24826, n24827, n24828, n24829, n24830, n24831, n24832, n24833,
         n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841,
         n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849,
         n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857,
         n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865,
         n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873,
         n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881,
         n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889,
         n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897,
         n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905,
         n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913,
         n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921,
         n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929,
         n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937,
         n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945,
         n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953,
         n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961,
         n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969,
         n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977,
         n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985,
         n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993,
         n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001,
         n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009,
         n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017,
         n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025,
         n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033,
         n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041,
         n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049,
         n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057,
         n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065,
         n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073,
         n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081,
         n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089,
         n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097,
         n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105,
         n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113,
         n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121,
         n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129,
         n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137,
         n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145,
         n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153,
         n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161,
         n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169,
         n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177,
         n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185,
         n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193,
         n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201,
         n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209,
         n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217,
         n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225,
         n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233,
         n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241,
         n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249,
         n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257,
         n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265,
         n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273,
         n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281,
         n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289,
         n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297,
         n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305,
         n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313,
         n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321,
         n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329,
         n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337,
         n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345,
         n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353,
         n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361,
         n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369,
         n25370, n25371, n25372, n25373, n25374, n25375, n25376, n25377,
         n25378, n25379, n25380, n25381, n25382, n25383, n25384, n25385,
         n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393,
         n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401,
         n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409,
         n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417,
         n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425,
         n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433,
         n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441,
         n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449,
         n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457,
         n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465,
         n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473,
         n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481,
         n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489,
         n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497,
         n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505,
         n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513,
         n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521,
         n25522, n25523, n25524, n25525, n25526, n25527, n25528, n25529,
         n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537,
         n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545,
         n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553,
         n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561,
         n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569,
         n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577,
         n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585,
         n25586, n25587, n25588, n25589, n25590, n25591, n25592, n25593,
         n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601,
         n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609,
         n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617,
         n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625,
         n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25633,
         n25634, n25635, n25636, n25637, n25638, n25639, n25640, n25641,
         n25642, n25643, n25644, n25645, n25646, n25647, n25648, n25649,
         n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657,
         n25658, n25659, n25660, n25661, n25662, n25663, n25664, n25665,
         n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673,
         n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681,
         n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689,
         n25690, n25691, n25692, n25693, n25694, n25695, n25696, n25697,
         n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25705,
         n25706, n25707, n25708, n25709, n25710, n25711, n25712, n25713,
         n25714, n25715, n25716, n25717, n25718, n25719, n25720, n25721,
         n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729,
         n25730, n25731, n25732, n25733, n25734, n25735, n25736, n25737,
         n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745,
         n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753,
         n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761,
         n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769,
         n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777,
         n25778, n25779, n25780, n25781, n25782, n25783, n25784, n25785,
         n25786, n25787, n25788, n25789, n25790, n25791, n25792, n25793,
         n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801,
         n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809,
         n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817,
         n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825,
         n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833,
         n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841,
         n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849,
         n25850, n25851, n25852, n25853, n25854, n25855, n25856, n25857,
         n25858, n25859, n25860, n25861, n25862, n25863, n25864, n25865,
         n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873,
         n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881,
         n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25889,
         n25890, n25891, n25892, n25893, n25894, n25895, n25896, n25897,
         n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905,
         n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913,
         n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921,
         n25922, n25923, n25924, n25925, n25926, n25927, n25928, n25929,
         n25930, n25931, n25932, n25933, n25934, n25935, n25936, n25937,
         n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25945,
         n25946, n25947, n25948, n25949, n25950, n25951, n25952, n25953,
         n25954, n25955, n25956, n25957, n25958, n25959, n25960, n25961,
         n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969,
         n25970, n25971, n25972, n25973, n25974, n25975, n25976, n25977,
         n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25985,
         n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993,
         n25994, n25995, n25996, n25997, n25998, n25999, n26000, n26001,
         n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26009,
         n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017,
         n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025,
         n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26033,
         n26034, n26035, n26036, n26037, n26038, n26039, n26040, n26041,
         n26042, n26043, n26044, n26045, n26046, n26047, n26048, n26049,
         n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057,
         n26058, n26059, n26060, n26061, n26062, n26063, n26064, n26065,
         n26066, n26067, n26068, n26069, n26070, n26071, n26072, n26073,
         n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081,
         n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089,
         n26090, n26091, n26092, n26093, n26094, n26095, n26096, n26097,
         n26098, n26099, n26100, n26101, n26102, n26103, n26104, n26105,
         n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113,
         n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121,
         n26122, n26123, n26124, n26125, n26126, n26127, n26128, n26129,
         n26130, n26131, n26132, n26133, n26134, n26135, n26136, n26137,
         n26138, n26139, n26140, n26141, n26142, n26143, n26144, n26145,
         n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153,
         n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161,
         n26162, n26163, n26164, n26165, n26166, n26167, n26168, n26169,
         n26170, n26171, n26172, n26173, n26174, n26175, n26176, n26177,
         n26178, n26179, n26180, n26181, n26182, n26183, n26184, n26185,
         n26186, n26187, n26188, n26189, n26190, n26191, n26192, n26193,
         n26194, n26195, n26196, n26197, n26198, n26199, n26200, n26201,
         n26202, n26203, n26204, n26205, n26206, n26207, n26208, n26209,
         n26210, n26211, n26212, n26213, n26214, n26215, n26216, n26217,
         n26218, n26219, n26220, n26221, n26222, n26223, n26224, n26225,
         n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233,
         n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241,
         n26242, n26243, n26244, n26245, n26246, n26247, n26248, n26249,
         n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257,
         n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265,
         n26266, n26267, n26268, n26269, n26270, n26271, n26272, n26273,
         n26274, n26275, n26276, n26277, n26278, n26279, n26280, n26281,
         n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289,
         n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297,
         n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305,
         n26306, n26307, n26308, n26309, n26310, n26311, n26312, n26313,
         n26314, n26315, n26316, n26317, n26318, n26319, n26320, n26321,
         n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329,
         n26330, n26331, n26332, n26333, n26334, n26335, n26336, n26337,
         n26338, n26339, n26340, n26341, n26342, n26343, n26344, n26345,
         n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26353,
         n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361,
         n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369,
         n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377,
         n26378, n26379, n26380, n26381, n26382, n26383, n26384, n26385,
         n26386, n26387, n26388, n26389, n26390, n26391, n26392, n26393,
         n26394, n26395, n26396, n26397, n26398, n26399, n26400, n26401,
         n26402, n26403, n26404, n26405, n26406, n26407, n26408, n26409,
         n26410, n26411, n26412, n26413, n26414, n26415, n26416, n26417,
         n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425,
         n26426, n26427, n26428, n26429, n26430, n26431, n26432, n26433,
         n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441,
         n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449,
         n26450, n26451, n26452, n26453, n26454, n26455, n26456, n26457,
         n26458, n26459, n26460, n26461, n26462, n26463, n26464, n26465,
         n26466, n26467, n26468, n26469, n26470, n26471, n26472, n26473,
         n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481,
         n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489,
         n26490, n26491, n26492, n26493, n26494, n26495, n26496, n26497,
         n26498, n26499, n26500, n26501, n26502, n26503, n26504, n26505,
         n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513,
         n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521,
         n26522, n26523, n26524, n26525, n26526, n26527, n26528, n26529,
         n26530, n26531, n26532, n26533, n26534, n26535, n26536, n26537,
         n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545,
         n26546, n26547, n26548, n26549, n26550, n26551, n26552, n26553,
         n26554, n26555, n26556, n26557, n26558, n26559, n26560, n26561,
         n26562, n26563, n26564, n26565, n26566, n26567, n26568, n26569,
         n26570, n26571, n26572, n26573, n26574, n26575, n26576, n26577,
         n26578, n26579, n26580, n26581, n26582, n26583, n26584, n26585,
         n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593,
         n26594, n26595, n26596, n26597, n26598, n26599, n26600, n26601,
         n26602, n26603, n26604, n26605, n26606, n26607, n26608, n26609,
         n26610, n26611, n26612, n26613, n26614, n26615, n26616, n26617,
         n26618, n26619, n26620, n26621, n26622, n26623, n26624, n26625,
         n26626, n26627, n26628, n26629, n26630, n26631, n26632, n26633,
         n26634, n26635, n26636, n26637, n26638, n26639, n26640, n26641,
         n26642, n26643, n26644, n26645, n26646, n26647, n26648, n26649,
         n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657,
         n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665,
         n26666, n26667, n26668, n26669, n26670, n26671, n26672, n26673,
         n26674, n26675, n26676, n26677, n26678, n26679, n26680, n26681,
         n26682, n26683, n26684, n26685, n26686, n26687, n26688, n26689,
         n26690, n26691, n26692, n26693, n26694, n26695, n26696, n26697,
         n26698, n26699, n26700, n26701, n26702, n26703, n26704, n26705,
         n26706, n26707, n26708, n26709, n26710, n26711, n26712, n26713,
         n26714, n26715, n26716, n26717, n26718, n26719, n26720, n26721,
         n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729,
         n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737,
         n26738, n26739, n26740, n26741, n26742, n26743, n26744, n26745,
         n26746, n26747, n26748, n26749, n26750, n26751, n26752, n26753,
         n26754, n26755, n26756, n26757, n26758, n26759, n26760, n26761,
         n26762, n26763, n26764, n26765, n26766, n26767, n26768, n26769,
         n26770, n26771, n26772, n26773, n26774, n26775, n26776, n26777,
         n26778, n26779, n26780, n26781, n26782, n26783, n26784, n26785,
         n26786, n26787, n26788, n26789, n26790, n26791, n26792, n26793,
         n26794, n26795, n26796, n26797, n26798, n26799, n26800, n26801,
         n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809,
         n26810, n26811, n26812, n26813, n26814, n26815, n26816, n26817,
         n26818, n26819, n26820, n26821, n26822, n26823, n26824, n26825,
         n26826, n26827, n26828, n26829, n26830, n26831, n26832, n26833,
         n26834, n26835, n26836, n26837, n26838, n26839, n26840, n26841,
         n26842, n26843, n26844, n26845, n26846, n26847, n26848, n26849,
         n26850, n26851, n26852, n26853, n26854, n26855, n26856, n26857,
         n26858, n26859, n26860, n26861, n26862, n26863, n26864, n26865,
         n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873,
         n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881,
         n26882, n26883, n26884, n26885, n26886, n26887, n26888, n26889,
         n26890, n26891, n26892, n26893, n26894, n26895, n26896, n26897,
         n26898, n26899, n26900, n26901, n26902, n26903, n26904, n26905,
         n26906, n26907, n26908, n26909, n26910, n26911, n26912, n26913,
         n26914, n26915, n26916, n26917, n26918, n26919, n26920, n26921,
         n26922, n26923, n26924, n26925, n26926, n26927, n26928, n26929,
         n26930, n26931, n26932, n26933, n26934, n26935, n26936, n26937,
         n26938, n26939, n26940, n26941, n26942, n26943, n26944, n26945,
         n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953,
         n26954, n26955, n26956, n26957, n26958, n26959, n26960, n26961,
         n26962, n26963, n26964, n26965, n26966, n26967, n26968, n26969,
         n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977,
         n26978, n26979, n26980, n26981, n26982, n26983, n26984, n26985,
         n26986, n26987, n26988, n26989, n26990, n26991, n26992, n26993,
         n26994, n26995, n26996, n26997, n26998, n26999, n27000, n27001,
         n27002, n27003, n27004, n27005, n27006, n27007, n27008, n27009,
         n27010, n27011, n27012, n27013, n27014, n27015, n27016, n27017,
         n27018, n27019, n27020, n27021, n27022, n27023, n27024, n27025,
         n27026, n27027, n27028, n27029, n27030, n27031, n27032, n27033,
         n27034, n27035, n27036, n27037, n27038, n27039, n27040, n27041,
         n27042, n27043, n27044, n27045, n27046, n27047, n27048, n27049,
         n27050, n27051, n27052, n27053, n27054, n27055, n27056, n27057,
         n27058, n27059, n27060, n27061, n27062, n27063, n27064, n27065,
         n27066, n27067, n27068, n27069, n27070, n27071, n27072, n27073,
         n27074, n27075, n27076, n27077, n27078, n27079, n27080, n27081,
         n27082, n27083, n27084, n27085, n27086, n27087, n27088, n27089,
         n27090, n27091, n27092, n27093, n27094, n27095, n27096, n27097,
         n27098, n27099, n27100, n27101, n27102, n27103, n27104, n27105,
         n27106, n27107, n27108, n27109, n27110, n27111, n27112, n27113,
         n27114, n27115, n27116, n27117, n27118, n27119, n27120, n27121,
         n27122, n27123, n27124, n27125, n27126, n27127, n27128, n27129,
         n27130, n27131, n27132, n27133, n27134, n27135, n27136, n27137,
         n27138, n27139, n27140, n27141, n27142, n27143, n27144, n27145,
         n27146, n27147, n27148, n27149, n27150, n27151, n27152, n27153,
         n27154, n27155, n27156, n27157, n27158, n27159, n27160, n27161,
         n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169,
         n27170, n27171, n27172, n27173, n27174, n27175, n27176, n27177,
         n27178, n27179, n27180, n27181, n27182, n27183, n27184, n27185,
         n27186, n27187, n27188, n27189, n27190, n27191, n27192, n27193,
         n27194, n27195, n27196, n27197, n27198, n27199, n27200, n27201,
         n27202, n27203, n27204, n27205, n27206, n27207, n27208, n27209,
         n27210, n27211, n27212, n27213, n27214, n27215, n27216, n27217,
         n27218, n27219, n27220, n27221, n27222, n27223, n27224, n27225,
         n27226, n27227, n27228, n27229, n27230, n27231, n27232, n27233,
         n27234, n27235, n27236, n27237, n27238, n27239, n27240, n27241,
         n27242, n27243, n27244, n27245, n27246, n27247, n27248, n27249,
         n27250, n27251, n27252, n27253, n27254, n27255, n27256, n27257,
         n27258, n27259, n27260, n27261, n27262, n27263, n27264, n27265,
         n27266, n27267, n27268, n27269, n27270, n27271, n27272, n27273,
         n27274, n27275, n27276, n27277, n27278, n27279, n27280, n27281,
         n27282, n27283, n27284, n27285, n27286, n27287, n27288, n27289,
         n27290, n27291, n27292, n27293, n27294, n27295, n27296, n27297,
         n27298, n27299, n27300, n27301, n27302, n27303, n27304, n27305,
         n27306, n27307, n27308, n27309, n27310, n27311, n27312, n27313,
         n27314, n27315, n27316, n27317, n27318, n27319, n27320, n27321,
         n27322, n27323, n27324, n27325, n27326, n27327, n27328, n27329,
         n27330, n27331, n27332, n27333, n27334, n27335, n27336, n27337,
         n27338, n27339, n27340, n27341, n27342, n27343, n27344, n27345,
         n27346, n27347, n27348, n27349, n27350, n27351, n27352, n27353,
         n27354, n27355, n27356, n27357, n27358, n27359, n27360, n27361,
         n27362, n27363, n27364, n27365, n27366, n27367, n27368, n27369,
         n27370, n27371, n27372, n27373, n27374, n27375, n27376, n27377,
         n27378, n27379, n27380, n27381, n27382, n27383, n27384, n27385,
         n27386, n27387, n27388, n27389, n27390, n27391, n27392, n27393,
         n27394, n27395, n27396, n27397, n27398, n27399, n27400, n27401,
         n27402, n27403, n27404, n27405, n27406, n27407, n27408, n27409,
         n27410, n27411, n27412, n27413, n27414, n27415, n27416, n27417,
         n27418, n27419, n27420, n27421, n27422, n27423, n27424, n27425,
         n27426, n27427, n27428, n27429, n27430, n27431, n27432, n27433,
         n27434, n27435, n27436, n27437, n27438, n27439, n27440, n27441,
         n27442, n27443, n27444, n27445, n27446, n27447, n27448, n27449,
         n27450, n27451, n27452, n27453, n27454, n27455, n27456, n27457,
         n27458, n27459, n27460, n27461, n27462, n27463, n27464, n27465,
         n27466, n27467, n27468, n27469, n27470, n27471, n27472, n27473,
         n27474, n27475, n27476, n27477, n27478, n27479, n27480, n27481,
         n27482, n27483, n27484, n27485, n27486, n27487, n27488, n27489,
         n27490, n27491, n27492, n27493, n27494, n27495, n27496, n27497,
         n27498, n27499, n27500, n27501, n27502, n27503, n27504, n27505,
         n27506, n27507, n27508, n27509, n27510, n27511, n27512, n27513,
         n27514, n27515, n27516, n27517, n27518, n27519, n27520, n27521,
         n27522, n27523, n27524, n27525, n27526, n27527, n27528, n27529,
         n27530, n27531, n27532, n27533, n27534, n27535, n27536, n27537,
         n27538, n27539, n27540, n27541, n27542, n27543, n27544, n27545,
         n27546, n27547, n27548, n27549, n27550, n27551, n27552, n27553,
         n27554, n27555, n27556, n27557, n27558, n27559, n27560, n27561,
         n27562, n27563, n27564, n27565, n27566, n27567, n27568, n27569,
         n27570, n27571, n27572, n27573, n27574, n27575, n27576, n27577,
         n27578, n27579, n27580, n27581, n27582, n27583, n27584, n27585,
         n27586, n27587, n27588, n27589, n27590, n27591, n27592, n27593,
         n27594, n27595, n27596, n27597, n27598, n27599, n27600, n27601,
         n27602, n27603, n27604, n27605, n27606, n27607, n27608, n27609,
         n27610, n27611, n27612, n27613, n27614, n27615, n27616, n27617,
         n27618, n27619, n27620, n27621, n27622, n27623, n27624, n27625,
         n27626, n27627, n27628, n27629, n27630, n27631, n27632, n27633,
         n27634, n27635, n27636, n27637, n27638, n27639, n27640, n27641,
         n27642, n27643, n27644, n27645, n27646, n27647, n27648, n27649,
         n27650, n27651, n27652, n27653, n27654, n27655, n27656, n27657,
         n27658, n27659, n27660, n27661, n27662, n27663, n27664, n27665,
         n27666, n27667, n27668, n27669, n27670, n27671, n27672, n27673,
         n27674, n27675, n27676, n27677, n27678, n27679, n27680, n27681,
         n27682, n27683, n27684, n27685, n27686, n27687, n27688, n27689,
         n27690, n27691, n27692, n27693, n27694, n27695, n27696, n27697,
         n27698, n27699, n27700, n27701, n27702, n27703, n27704, n27705,
         n27706, n27707, n27708, n27709, n27710, n27711, n27712, n27713,
         n27714, n27715, n27716, n27717, n27718, n27719, n27720, n27721,
         n27722, n27723, n27724, n27725, n27726, n27727, n27728, n27729,
         n27730, n27731, n27732, n27733, n27734, n27735, n27736, n27737,
         n27738, n27739, n27740, n27741, n27742, n27743, n27744, n27745,
         n27746, n27747, n27748, n27749, n27750, n27751, n27752, n27753,
         n27754, n27755, n27756, n27757, n27758, n27759, n27760, n27761,
         n27762, n27763, n27764, n27765, n27766, n27767, n27768, n27769,
         n27770, n27771, n27772, n27773, n27774, n27775, n27776, n27777,
         n27778, n27779, n27780, n27781, n27782, n27783, n27784, n27785,
         n27786, n27787, n27788, n27789, n27790, n27791, n27792, n27793,
         n27794, n27795, n27796, n27797, n27798, n27799, n27800, n27801,
         n27802, n27803, n27804, n27805, n27806, n27807, n27808, n27809,
         n27810, n27811, n27812, n27813, n27814, n27815, n27816, n27817,
         n27818, n27819, n27820, n27821, n27822, n27823, n27824, n27825,
         n27826, n27827, n27828, n27829, n27830, n27831, n27832, n27833,
         n27834, n27835, n27836, n27837, n27838, n27839, n27840, n27841,
         n27842, n27843, n27844, n27845, n27846, n27847, n27848, n27849,
         n27850, n27851, n27852, n27853, n27854, n27855, n27856, n27857,
         n27858, n27859, n27860, n27861, n27862, n27863, n27864, n27865,
         n27866, n27867, n27868, n27869, n27870, n27871, n27872, n27873,
         n27874, n27875, n27876, n27877, n27878, n27879, n27880, n27881,
         n27882, n27883, n27884, n27885, n27886, n27887, n27888, n27889,
         n27890, n27891, n27892, n27893, n27894, n27895, n27896, n27897,
         n27898, n27899, n27900, n27901, n27902, n27903, n27904, n27905,
         n27906, n27907, n27908, n27909, n27910, n27911, n27912, n27913,
         n27914, n27915, n27916, n27917, n27918, n27919, n27920, n27921,
         n27922, n27923, n27924, n27925, n27926, n27927, n27928, n27929,
         n27930, n27931, n27932, n27933, n27934, n27935, n27936, n27937,
         n27938, n27939, n27940, n27941, n27942, n27943, n27944, n27945,
         n27946, n27947, n27948, n27949, n27950, n27951, n27952, n27953,
         n27954, n27955, n27956, n27957, n27958, n27959, n27960, n27961,
         n27962, n27963, n27964, n27965, n27966, n27967, n27968, n27969,
         n27970, n27971, n27972, n27973, n27974, n27975, n27976, n27977,
         n27978, n27979, n27980, n27981, n27982, n27983, n27984, n27985,
         n27986, n27987, n27988, n27989, n27990, n27991, n27992, n27993,
         n27994, n27995, n27996, n27997, n27998, n27999, n28000, n28001,
         n28002, n28003, n28004, n28005, n28006, n28007, n28008, n28009,
         n28010, n28011, n28012, n28013, n28014, n28015, n28016, n28017,
         n28018, n28019, n28020, n28021, n28022, n28023, n28024, n28025,
         n28026, n28027, n28028, n28029, n28030, n28031, n28032, n28033,
         n28034, n28035, n28036, n28037, n28038, n28039, n28040, n28041,
         n28042, n28043, n28044, n28045, n28046, n28047, n28048, n28049,
         n28050, n28051, n28052, n28053, n28054, n28055, n28056, n28057,
         n28058, n28059, n28060, n28061, n28062, n28063, n28064, n28065,
         n28066, n28067, n28068, n28069, n28070, n28071, n28072, n28073,
         n28074, n28075, n28076, n28077, n28078, n28079, n28080, n28081,
         n28082, n28083, n28084, n28085, n28086, n28087, n28088, n28089,
         n28090, n28091, n28092, n28093, n28094, n28095, n28096, n28097,
         n28098, n28099, n28100, n28101, n28102, n28103, n28104, n28105,
         n28106, n28107, n28108, n28109, n28110, n28111, n28112, n28113,
         n28114, n28115, n28116, n28117, n28118, n28119, n28120, n28121,
         n28122, n28123, n28124, n28125, n28126, n28127, n28128, n28129,
         n28130, n28131, n28132, n28133, n28134, n28135, n28136, n28137,
         n28138, n28139, n28140, n28141, n28142, n28143, n28144, n28145,
         n28146, n28147, n28148, n28149, n28150, n28151, n28152, n28153,
         n28154, n28155, n28156, n28157, n28158, n28159, n28160, n28161,
         n28162, n28163, n28164, n28165, n28166, n28167, n28168, n28169,
         n28170, n28171, n28172, n28173, n28174, n28175, n28176, n28177,
         n28178, n28179, n28180, n28181, n28182, n28183, n28184, n28185,
         n28186, n28187, n28188, n28189, n28190, n28191, n28192, n28193,
         n28194, n28195, n28196, n28197, n28198, n28199, n28200, n28201,
         n28202, n28203, n28204, n28205, n28206, n28207, n28208, n28209,
         n28210, n28211, n28212, n28213, n28214, n28215, n28216, n28217,
         n28218, n28219, n28220, n28221, n28222, n28223, n28224, n28225,
         n28226, n28227, n28228, n28229, n28230, n28231, n28232, n28233,
         n28234, n28235, n28236, n28237, n28238, n28239, n28240, n28241,
         n28242, n28243, n28244, n28245, n28246, n28247, n28248, n28249,
         n28250, n28251, n28252, n28253, n28254, n28255, n28256, n28257,
         n28258, n28259, n28260, n28261, n28262, n28263, n28264, n28265,
         n28266, n28267, n28268, n28269, n28270, n28271, n28272, n28273,
         n28274, n28275, n28276, n28277, n28278, n28279, n28280, n28281,
         n28282, n28283, n28284, n28285, n28286, n28287, n28288, n28289,
         n28290, n28291, n28292, n28293, n28294, n28295, n28296, n28297,
         n28298, n28299, n28300, n28301, n28302, n28303, n28304, n28305,
         n28306, n28307, n28308, n28309, n28310, n28311, n28312, n28313,
         n28314, n28315, n28316, n28317, n28318, n28319, n28320, n28321,
         n28322, n28323, n28324, n28325, n28326, n28327, n28328, n28329,
         n28330, n28331, n28332, n28333, n28334, n28335, n28336, n28337,
         n28338, n28339, n28340, n28341, n28342, n28343, n28344, n28345,
         n28346, n28347, n28348, n28349, n28350, n28351, n28352, n28353,
         n28354, n28355, n28356, n28357, n28358, n28359, n28360, n28361,
         n28362, n28363, n28364, n28365, n28366, n28367, n28368, n28369,
         n28370, n28371, n28372, n28373, n28374, n28375, n28376, n28377,
         n28378, n28379, n28380, n28381, n28382, n28383, n28384, n28385,
         n28386, n28387, n28388, n28389, n28390, n28391, n28392, n28393,
         n28394, n28395, n28396, n28397, n28398, n28399, n28400, n28401,
         n28402, n28403, n28404, n28405, n28406, n28407, n28408, n28409,
         n28410, n28411, n28412, n28413, n28414, n28415, n28416, n28417,
         n28418, n28419, n28420, n28421, n28422, n28423, n28424, n28425,
         n28426, n28427, n28428, n28429, n28430, n28431, n28432, n28433,
         n28434, n28435, n28436, n28437, n28438, n28439, n28440, n28441,
         n28442, n28443, n28444, n28445, n28446, n28447, n28448, n28449,
         n28450, n28451, n28452, n28453, n28454, n28455, n28456, n28457,
         n28458, n28459, n28460, n28461, n28462, n28463, n28464, n28465,
         n28466, n28467, n28468, n28469, n28470, n28471, n28472, n28473,
         n28474, n28475, n28476, n28477, n28478, n28479, n28480, n28481,
         n28482, n28483, n28484, n28485, n28486, n28487, n28488, n28489,
         n28490, n28491, n28492, n28493, n28494, n28495, n28496, n28497,
         n28498, n28499, n28500, n28501, n28502, n28503, n28504, n28505,
         n28506, n28507, n28508, n28509, n28510, n28511, n28512, n28513,
         n28514, n28515, n28516, n28517, n28518, n28519, n28520, n28521,
         n28522, n28523, n28524, n28525, n28526, n28527, n28528, n28529,
         n28530, n28531, n28532, n28533, n28534, n28535, n28536, n28537,
         n28538, n28539, n28540, n28541, n28542, n28543, n28544, n28545,
         n28546, n28547, n28548, n28549, n28550, n28551, n28552, n28553,
         n28554, n28555, n28556, n28557, n28558, n28559, n28560, n28561,
         n28562, n28563, n28564, n28565, n28566, n28567, n28568, n28569,
         n28570, n28571, n28572, n28573, n28574, n28575, n28576, n28577,
         n28578, n28579, n28580, n28581, n28582, n28583, n28584, n28585,
         n28586, n28587, n28588, n28589, n28590, n28591, n28592, n28593,
         n28594, n28595, n28596, n28597, n28598, n28599, n28600, n28601,
         n28602, n28603, n28604, n28605, n28606, n28607, n28608, n28609,
         n28610, n28611, n28612, n28613, n28614, n28615, n28616, n28617,
         n28618, n28619, n28620, n28621, n28622, n28623, n28624, n28625,
         n28626, n28627, n28628, n28629, n28630, n28631, n28632, n28633,
         n28634, n28635, n28636, n28637, n28638, n28639, n28640, n28641,
         n28642, n28643, n28644, n28645, n28646, n28647, n28648, n28649,
         n28650, n28651, n28652, n28653, n28654, n28655, n28656, n28657,
         n28658, n28659, n28660, n28661, n28662, n28663, n28664, n28665,
         n28666, n28667, n28668, n28669, n28670, n28671, n28672, n28673,
         n28674, n28675, n28676, n28677, n28678, n28679, n28680, n28681,
         n28682, n28683, n28684, n28685, n28686, n28687, n28688, n28689,
         n28690, n28691, n28692, n28693, n28694, n28695, n28696, n28697,
         n28698, n28699, n28700, n28701, n28702, n28703, n28704, n28705,
         n28706, n28707, n28708, n28709, n28710, n28711, n28712, n28713,
         n28714, n28715, n28716, n28717, n28718, n28719, n28720, n28721,
         n28722, n28723, n28724, n28725, n28726, n28727, n28728, n28729,
         n28730, n28731, n28732, n28733, n28734, n28735, n28736, n28737,
         n28738, n28739, n28740, n28741, n28742, n28743, n28744, n28745,
         n28746, n28747, n28748, n28749, n28750, n28751, n28752, n28753,
         n28754, n28755, n28756, n28757, n28758, n28759, n28760, n28761,
         n28762, n28763, n28764, n28765, n28766, n28767, n28768, n28769,
         n28770, n28771, n28772, n28773, n28774, n28775, n28776, n28777,
         n28778, n28779, n28780, n28781, n28782, n28783, n28784, n28785,
         n28786, n28787, n28788, n28789, n28790, n28791, n28792, n28793,
         n28794, n28795, n28796, n28797, n28798, n28799, n28800, n28801,
         n28802, n28803, n28804, n28805, n28806, n28807, n28808, n28809,
         n28810, n28811, n28812, n28813, n28814, n28815, n28816, n28817,
         n28818, n28819, n28820, n28821, n28822, n28823, n28824, n28825,
         n28826, n28827, n28828, n28829, n28830, n28831, n28832, n28833,
         n28834, n28835, n28836, n28837, n28838, n28839, n28840, n28841,
         n28842, n28843, n28844, n28845, n28846, n28847, n28848, n28849,
         n28850, n28851, n28852, n28853, n28854, n28855, n28856, n28857,
         n28858, n28859, n28860, n28861, n28862, n28863, n28864, n28865,
         n28866, n28867, n28868, n28869, n28870, n28871, n28872, n28873,
         n28874, n28875, n28876, n28877, n28878, n28879, n28880, n28881,
         n28882, n28883, n28884, n28885, n28886, n28887, n28888, n28889,
         n28890, n28891, n28892, n28893, n28894, n28895, n28896, n28897,
         n28898, n28899, n28900, n28901, n28902, n28903, n28904, n28905,
         n28906, n28907, n28908, n28909, n28910, n28911, n28912, n28913,
         n28914, n28915, n28916, n28917, n28918, n28919, n28920, n28921,
         n28922, n28923, n28924, n28925, n28926, n28927, n28928, n28929,
         n28930, n28931, n28932, n28933, n28934, n28935, n28936, n28937,
         n28938, n28939, n28940, n28941, n28942, n28943, n28944, n28945,
         n28946, n28947, n28948, n28949, n28950, n28951, n28952, n28953,
         n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961,
         n28962, n28963, n28964, n28965, n28966, n28967, n28968, n28969,
         n28970, n28971, n28972, n28973, n28974, n28975, n28976, n28977,
         n28978, n28979, n28980, n28981, n28982, n28983, n28984, n28985,
         n28986, n28987, n28988, n28989, n28990, n28991, n28992, n28993,
         n28994, n28995, n28996, n28997, n28998, n28999, n29000, n29001,
         n29002, n29003, n29004, n29005, n29006, n29007, n29008, n29009,
         n29010, n29011, n29012, n29013, n29014, n29015, n29016, n29017,
         n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025,
         n29026, n29027, n29028, n29029, n29030, n29031, n29032, n29033,
         n29034, n29035, n29036, n29037, n29038, n29039, n29040, n29041,
         n29042, n29043, n29044, n29045, n29046, n29047, n29048, n29049,
         n29050, n29051, n29052, n29053, n29054, n29055, n29056, n29057,
         n29058, n29059, n29060, n29061, n29062, n29063, n29064, n29065,
         n29066, n29067, n29068, n29069, n29070, n29071, n29072, n29073,
         n29074, n29075, n29076, n29077, n29078, n29079, n29080, n29081,
         n29082, n29083, n29084, n29085, n29086, n29087, n29088, n29089,
         n29090, n29091, n29092, n29093, n29094, n29095, n29096, n29097,
         n29098, n29099, n29100, n29101, n29102, n29103, n29104, n29105,
         n29106, n29107, n29108, n29109, n29110, n29111, n29112, n29113,
         n29114, n29115, n29116, n29117, n29118, n29119, n29120, n29121,
         n29122, n29123, n29124, n29125, n29126, n29127, n29128, n29129,
         n29130, n29131, n29132, n29133, n29134, n29135, n29136, n29137,
         n29138, n29139, n29140, n29141, n29142, n29143, n29144, n29145,
         n29146, n29147, n29148, n29149, n29150, n29151, n29152, n29153,
         n29154, n29155, n29156, n29157, n29158, n29159, n29160, n29161,
         n29162, n29163, n29164, n29165, n29166, n29167, n29168, n29169,
         n29170, n29171, n29172, n29173, n29174, n29175, n29176, n29177,
         n29178, n29179, n29180, n29181, n29182, n29183, n29184, n29185,
         n29186, n29187, n29188, n29189, n29190, n29191, n29192, n29193,
         n29194, n29195, n29196, n29197, n29198, n29199, n29200, n29201,
         n29202, n29203, n29204, n29205, n29206, n29207, n29208, n29209,
         n29210, n29211, n29212, n29213, n29214, n29215, n29216, n29217,
         n29218, n29219, n29220, n29221, n29222, n29223, n29224, n29225,
         n29226, n29227, n29228, n29229, n29230, n29231, n29232, n29233,
         n29234, n29235, n29236, n29237, n29238, n29239, n29240, n29241,
         n29242, n29243, n29244, n29245, n29246, n29247, n29248, n29249,
         n29250, n29251, n29252, n29253, n29254, n29255, n29256, n29257,
         n29258, n29259, n29260, n29261, n29262, n29263, n29264, n29265,
         n29266, n29267, n29268, n29269, n29270, n29271, n29272, n29273,
         n29274, n29275, n29276, n29277, n29278, n29279, n29280, n29281,
         n29282, n29283, n29284, n29285, n29286, n29287, n29288, n29289,
         n29290, n29291, n29292, n29293, n29294, n29295, n29296, n29297,
         n29298, n29299, n29300, n29301, n29302, n29303, n29304, n29305,
         n29306, n29307, n29308, n29309, n29310, n29311, n29312, n29313,
         n29314, n29315, n29316, n29317, n29318, n29319, n29320, n29321,
         n29322, n29323, n29324, n29325, n29326, n29327, n29328, n29329,
         n29330, n29331, n29332, n29333, n29334, n29335, n29336, n29337,
         n29338, n29339, n29340, n29341, n29342, n29343, n29344, n29345,
         n29346, n29347, n29348, n29349, n29350, n29351, n29352, n29353,
         n29354, n29355, n29356, n29357, n29358, n29359, n29360, n29361,
         n29362, n29363, n29364, n29365, n29366, n29367, n29368, n29369,
         n29370, n29371, n29372, n29373, n29374, n29375, n29376, n29377,
         n29378, n29379, n29380, n29381, n29382, n29383, n29384, n29385,
         n29386, n29387, n29388, n29389, n29390, n29391, n29392, n29393,
         n29394, n29395, n29396, n29397, n29398, n29399, n29400, n29401,
         n29402, n29403, n29404, n29405, n29406, n29407, n29408, n29409,
         n29410, n29411, n29412, n29413, n29414, n29415, n29416, n29417,
         n29418, n29419, n29420, n29421, n29422, n29423, n29424, n29425,
         n29426, n29427, n29428, n29429, n29430, n29431, n29432, n29433,
         n29434, n29435, n29436, n29437, n29438, n29439, n29440, n29441,
         n29442, n29443, n29444, n29445, n29446, n29447, n29448, n29449,
         n29450, n29451, n29452, n29453, n29454, n29455, n29456, n29457,
         n29458, n29459, n29460, n29461, n29462, n29463, n29464, n29465,
         n29466, n29467, n29468, n29469, n29470, n29471, n29472, n29473,
         n29474, n29475, n29476, n29477, n29478, n29479, n29480, n29481,
         n29482, n29483, n29484, n29485, n29486, n29487, n29488, n29489,
         n29490, n29491, n29492, n29493, n29494, n29495, n29496, n29497,
         n29498, n29499, n29500, n29501, n29502, n29503, n29504, n29505,
         n29506, n29507, n29508, n29509, n29510, n29511, n29512, n29513,
         n29514, n29515, n29516, n29517, n29518, n29519, n29520, n29521,
         n29522, n29523, n29524, n29525, n29526, n29527, n29528, n29529,
         n29530, n29531, n29532, n29533, n29534, n29535, n29536, n29537,
         n29538, n29539, n29540, n29541, n29542, n29543, n29544, n29545,
         n29546, n29547, n29548, n29549, n29550, n29551, n29552, n29553,
         n29554, n29555, n29556, n29557, n29558, n29559, n29560, n29561,
         n29562, n29563, n29564, n29565, n29566, n29567, n29568, n29569,
         n29570, n29571, n29572, n29573, n29574, n29575, n29576, n29577,
         n29578, n29579, n29580, n29581, n29582, n29583, n29584, n29585,
         n29586, n29587, n29588, n29589, n29590, n29591, n29592, n29593,
         n29594, n29595, n29596, n29597, n29598, n29599, n29600, n29601,
         n29602, n29603, n29604, n29605, n29606, n29607, n29608, n29609,
         n29610, n29611, n29612, n29613, n29614, n29615, n29616, n29617,
         n29618, n29619, n29620, n29621, n29622, n29623, n29624, n29625,
         n29626, n29627, n29628, n29629, n29630, n29631, n29632, n29633,
         n29634, n29635, n29636, n29637, n29638, n29639, n29640, n29641,
         n29642, n29643, n29644, n29645, n29646, n29647, n29648, n29649,
         n29650, n29651, n29652, n29653, n29654, n29655, n29656, n29657,
         n29658, n29659, n29660, n29661, n29662, n29663, n29664, n29665,
         n29666, n29667, n29668, n29669, n29670, n29671, n29672, n29673,
         n29674, n29675, n29676, n29677, n29678, n29679, n29680, n29681,
         n29682, n29683, n29684, n29685, n29686, n29687, n29688, n29689,
         n29690, n29691, n29692, n29693, n29694, n29695, n29696, n29697,
         n29698, n29699, n29700, n29701, n29702, n29703, n29704, n29705,
         n29706, n29707, n29708, n29709, n29710, n29711, n29712, n29713,
         n29714, n29715, n29716, n29717, n29718, n29719, n29720, n29721,
         n29722, n29723, n29724, n29725, n29726, n29727, n29728, n29729,
         n29730, n29731, n29732, n29733, n29734, n29735, n29736, n29737,
         n29738, n29739, n29740, n29741, n29742, n29743, n29744, n29745,
         n29746, n29747, n29748, n29749, n29750, n29751, n29752, n29753,
         n29754, n29755, n29756, n29757, n29758, n29759, n29760, n29761,
         n29762, n29763, n29764, n29765, n29766, n29767, n29768, n29769,
         n29770, n29771, n29772, n29773, n29774, n29775, n29776, n29777,
         n29778, n29779, n29780, n29781, n29782, n29783, n29784, n29785,
         n29786, n29787, n29788, n29789, n29790, n29791, n29792, n29793,
         n29794, n29795, n29796, n29797, n29798, n29799, n29800, n29801,
         n29802, n29803, n29804, n29805, n29806, n29807, n29808, n29809,
         n29810, n29811, n29812, n29813, n29814, n29815, n29816, n29817,
         n29818, n29819, n29820, n29821, n29822, n29823, n29824, n29825,
         n29826, n29827, n29828, n29829, n29830, n29831, n29832, n29833,
         n29834, n29835, n29836, n29837, n29838, n29839, n29840, n29841,
         n29842, n29843, n29844, n29845, n29846, n29847, n29848, n29849,
         n29850, n29851, n29852, n29853, n29854, n29855, n29856, n29857,
         n29858, n29859, n29860, n29861, n29862, n29863, n29864, n29865,
         n29866, n29867, n29868, n29869, n29870, n29871, n29872, n29873,
         n29874, n29875, n29876, n29877, n29878, n29879, n29880, n29881,
         n29882, n29883, n29884, n29885, n29886, n29887, n29888, n29889,
         n29890, n29891, n29892, n29893, n29894, n29895, n29896, n29897,
         n29898, n29899, n29900, n29901, n29902, n29903, n29904, n29905,
         n29906, n29907, n29908, n29909, n29910, n29911, n29912, n29913,
         n29914, n29915, n29916, n29917, n29918, n29919, n29920, n29921,
         n29922, n29923, n29924, n29925, n29926, n29927, n29928, n29929,
         n29930, n29931, n29932, n29933, n29934, n29935, n29936, n29937,
         n29938, n29939, n29940, n29941, n29942, n29943, n29944, n29945,
         n29946, n29947, n29948, n29949, n29950, n29951, n29952, n29953,
         n29954, n29955, n29956, n29957, n29958, n29959, n29960, n29961,
         n29962, n29963, n29964, n29965, n29966, n29967, n29968, n29969,
         n29970, n29971, n29972, n29973, n29974, n29975, n29976, n29977,
         n29978, n29979, n29980, n29981, n29982, n29983, n29984, n29985,
         n29986, n29987, n29988, n29989, n29990, n29991, n29992, n29993,
         n29994, n29995, n29996, n29997, n29998, n29999, n30000, n30001,
         n30002, n30003, n30004, n30005, n30006, n30007, n30008, n30009,
         n30010, n30011, n30012, n30013, n30014, n30015, n30016, n30017,
         n30018, n30019, n30020, n30021, n30022, n30023, n30024, n30025,
         n30026, n30027, n30028, n30029, n30030, n30031, n30032, n30033,
         n30034, n30035, n30036, n30037, n30038, n30039, n30040, n30041,
         n30042, n30043, n30044, n30045, n30046, n30047, n30048, n30049,
         n30050, n30051, n30052, n30053, n30054, n30055, n30056, n30057,
         n30058, n30059, n30060, n30061, n30062, n30063, n30064, n30065,
         n30066, n30067, n30068, n30069, n30070, n30071, n30072, n30073,
         n30074, n30075, n30076, n30077, n30078, n30079, n30080, n30081,
         n30082, n30083, n30084, n30085, n30086, n30087, n30088, n30089,
         n30090, n30091, n30092, n30093, n30094, n30095, n30096, n30097,
         n30098, n30099, n30100, n30101, n30102, n30103, n30104, n30105,
         n30106, n30107, n30108, n30109, n30110, n30111, n30112, n30113,
         n30114, n30115, n30116, n30117, n30118, n30119, n30120, n30121,
         n30122, n30123, n30124, n30125, n30126, n30127, n30128, n30129,
         n30130, n30131, n30132, n30133, n30134, n30135, n30136, n30137,
         n30138, n30139, n30140, n30141, n30142, n30143, n30144, n30145,
         n30146, n30147, n30148, n30149, n30150, n30151, n30152, n30153,
         n30154, n30155, n30156, n30157, n30158, n30159, n30160, n30161,
         n30162, n30163, n30164, n30165, n30166, n30167, n30168, n30169,
         n30170, n30171, n30172, n30173, n30174, n30175, n30176, n30177,
         n30178, n30179, n30180, n30181, n30182, n30183, n30184, n30185,
         n30186, n30187, n30188, n30189, n30190, n30191, n30192, n30193,
         n30194, n30195, n30196, n30197, n30198, n30199, n30200, n30201,
         n30202, n30203, n30204, n30205, n30206, n30207, n30208, n30209,
         n30210, n30211, n30212, n30213, n30214, n30215, n30216, n30217,
         n30218, n30219, n30220, n30221, n30222, n30223, n30224, n30225,
         n30226, n30227, n30228, n30229, n30230, n30231, n30232, n30233,
         n30234, n30235, n30236, n30237, n30238, n30239, n30240, n30241,
         n30242, n30243, n30244, n30245, n30246, n30247, n30248, n30249,
         n30250, n30251, n30252, n30253, n30254, n30255, n30256, n30257,
         n30258, n30259, n30260, n30261, n30262, n30263, n30264, n30265,
         n30266, n30267, n30268, n30269, n30270, n30271, n30272, n30273,
         n30274, n30275, n30276, n30277, n30278, n30279, n30280, n30281,
         n30282, n30283, n30284, n30285, n30286, n30287, n30288, n30289,
         n30290, n30291, n30292, n30293, n30294, n30295, n30296, n30297,
         n30298, n30299, n30300, n30301, n30302, n30303, n30304, n30305,
         n30306, n30307, n30308, n30309, n30310, n30311, n30312, n30313,
         n30314, n30315, n30316, n30317, n30318, n30319, n30320, n30321,
         n30322, n30323, n30324, n30325, n30326, n30327, n30328, n30329,
         n30330, n30331, n30332, n30333, n30334, n30335, n30336, n30337,
         n30338, n30339, n30340, n30341, n30342, n30343, n30344, n30345,
         n30346, n30347, n30348, n30349, n30350, n30351, n30352, n30353,
         n30354, n30355, n30356, n30357, n30358, n30359, n30360, n30361,
         n30362, n30363, n30364, n30365, n30366, n30367, n30368, n30369,
         n30370, n30371, n30372, n30373, n30374, n30375, n30376, n30377,
         n30378, n30379, n30380, n30381, n30382, n30383, n30384, n30385,
         n30386, n30387, n30388, n30389, n30390, n30391, n30392, n30393,
         n30394, n30395, n30396, n30397, n30398, n30399, n30400, n30401,
         n30402, n30403, n30404, n30405, n30406, n30407, n30408, n30409,
         n30410, n30411, n30412, n30413, n30414, n30415, n30416, n30417,
         n30418, n30419, n30420, n30421, n30422, n30423, n30424, n30425,
         n30426, n30427, n30428, n30429, n30430, n30431, n30432, n30433,
         n30434, n30435, n30436, n30437, n30438, n30439, n30440, n30441,
         n30442, n30443, n30444, n30445, n30446, n30447, n30448, n30449,
         n30450, n30451, n30452, n30453, n30454, n30455, n30456, n30457,
         n30458, n30459, n30460, n30461, n30462, n30463, n30464, n30465,
         n30466, n30467, n30468, n30469, n30470, n30471, n30472, n30473,
         n30474, n30475, n30476, n30477, n30478, n30479, n30480, n30481,
         n30482, n30483, n30484, n30485, n30486, n30487, n30488, n30489,
         n30490, n30491, n30492, n30493, n30494, n30495, n30496, n30497,
         n30498, n30499, n30500, n30501, n30502, n30503, n30504, n30505,
         n30506, n30507, n30508, n30509, n30510, n30511, n30512, n30513,
         n30514, n30515, n30516, n30517, n30518, n30519, n30520, n30521,
         n30522, n30523, n30524, n30525, n30526, n30527, n30528, n30529,
         n30530, n30531, n30532, n30533, n30534, n30535, n30536, n30537,
         n30538, n30539, n30540, n30541, n30542, n30543, n30544, n30545,
         n30546, n30547, n30548, n30549, n30550, n30551, n30552, n30553,
         n30554, n30555, n30556, n30557, n30558, n30559, n30560, n30561,
         n30562, n30563, n30564, n30565, n30566, n30567, n30568, n30569,
         n30570, n30571, n30572, n30573, n30574, n30575, n30576, n30577,
         n30578, n30579, n30580, n30581, n30582, n30583, n30584, n30585,
         n30586, n30587, n30588, n30589, n30590, n30591, n30592, n30593,
         n30594, n30595, n30596, n30597, n30598, n30599, n30600, n30601,
         n30602, n30603, n30604, n30605, n30606, n30607, n30608, n30609,
         n30610, n30611, n30612, n30613, n30614, n30615, n30616, n30617,
         n30618, n30619, n30620, n30621, n30622, n30623, n30624, n30625,
         n30626, n30627, n30628, n30629, n30630, n30631, n30632, n30633,
         n30634, n30635, n30636, n30637, n30638, n30639, n30640, n30641,
         n30642, n30643, n30644, n30645, n30646, n30647, n30648, n30649,
         n30650, n30651, n30652, n30653, n30654, n30655, n30656, n30657,
         n30658, n30659, n30660, n30661, n30662, n30663, n30664, n30665,
         n30666, n30667, n30668, n30669, n30670, n30671, n30672, n30673,
         n30674, n30675, n30676, n30677, n30678, n30679, n30680, n30681,
         n30682, n30683, n30684, n30685, n30686, n30687, n30688, n30689,
         n30690, n30691, n30692, n30693, n30694, n30695, n30696, n30697,
         n30698, n30699, n30700, n30701, n30702, n30703, n30704, n30705,
         n30706, n30707, n30708, n30709, n30710, n30711, n30712, n30713,
         n30714, n30715, n30716, n30717, n30718, n30719, n30720, n30721,
         n30722, n30723, n30724, n30725, n30726, n30727, n30728, n30729,
         n30730, n30731, n30732, n30733, n30734, n30735, n30736, n30737,
         n30738, n30739, n30740, n30741, n30742, n30743, n30744, n30745,
         n30746, n30747, n30748, n30749, n30750, n30751, n30752, n30753,
         n30754, n30755, n30756, n30757, n30758, n30759, n30760, n30761,
         n30762, n30763, n30764, n30765, n30766, n30767, n30768, n30769,
         n30770, n30771, n30772, n30773, n30774, n30775, n30776, n30777,
         n30778, n30779, n30780, n30781, n30782, n30783, n30784, n30785,
         n30786, n30787, n30788, n30789, n30790, n30791, n30792, n30793,
         n30794, n30795, n30796, n30797, n30798, n30799, n30800, n30801,
         n30802, n30803, n30804, n30805, n30806, n30807, n30808, n30809,
         n30810, n30811, n30812, n30813, n30814, n30815, n30816, n30817,
         n30818, n30819, n30820, n30821, n30822, n30823, n30824, n30825,
         n30826, n30827, n30828, n30829, n30830, n30831, n30832, n30833,
         n30834, n30835, n30836, n30837, n30838, n30839, n30840, n30841,
         n30842, n30843, n30844, n30845, n30846, n30847, n30848, n30849,
         n30850, n30851, n30852, n30853, n30854, n30855, n30856, n30857,
         n30858, n30859, n30860, n30861, n30862, n30863, n30864, n30865,
         n30866, n30867, n30868, n30869, n30870, n30871, n30872, n30873,
         n30874, n30875, n30876, n30877, n30878, n30879, n30880, n30881,
         n30882, n30883, n30884, n30885, n30886, n30887, n30888, n30889,
         n30890, n30891, n30892, n30893, n30894, n30895, n30896, n30897,
         n30898, n30899, n30900, n30901, n30902, n30903, n30904, n30905,
         n30906, n30907, n30908, n30909, n30910, n30911, n30912, n30913,
         n30914, n30915, n30916, n30917, n30918, n30919, n30920, n30921,
         n30922, n30923, n30924, n30925, n30926, n30927, n30928, n30929,
         n30930, n30931, n30932, n30933, n30934, n30935, n30936, n30937,
         n30938, n30939, n30940, n30941, n30942, n30943, n30944, n30945,
         n30946, n30947, n30948, n30949, n30950, n30951, n30952, n30953,
         n30954, n30955, n30956, n30957, n30958, n30959, n30960, n30961,
         n30962, n30963, n30964, n30965, n30966, n30967, n30968, n30969,
         n30970, n30971, n30972, n30973, n30974, n30975, n30976, n30977,
         n30978, n30979, n30980, n30981, n30982, n30983, n30984, n30985,
         n30986, n30987, n30988, n30989, n30990, n30991, n30992, n30993,
         n30994, n30995, n30996, n30997, n30998, n30999, n31000, n31001,
         n31002, n31003, n31004, n31005, n31006, n31007, n31008, n31009,
         n31010, n31011, n31012, n31013, n31014, n31015, n31016, n31017,
         n31018, n31019, n31020, n31021, n31022, n31023, n31024, n31025,
         n31026, n31027, n31028, n31029, n31030, n31031, n31032, n31033,
         n31034, n31035, n31036, n31037, n31038, n31039, n31040, n31041,
         n31042, n31043, n31044, n31045, n31046, n31047, n31048, n31049,
         n31050, n31051, n31052, n31053, n31054, n31055, n31056, n31057,
         n31058, n31059, n31060, n31061, n31062, n31063, n31064, n31065,
         n31066, n31067, n31068, n31069, n31070, n31071, n31072, n31073,
         n31074, n31075, n31076, n31077, n31078, n31079, n31080, n31081,
         n31082, n31083, n31084, n31085, n31086, n31087, n31088, n31089,
         n31090, n31091, n31092, n31093, n31094, n31095, n31096, n31097,
         n31098, n31099, n31100, n31101, n31102, n31103, n31104, n31105,
         n31106, n31107, n31108, n31109, n31110, n31111, n31112, n31113,
         n31114, n31115, n31116, n31117, n31118, n31119, n31120, n31121,
         n31122, n31123, n31124, n31125, n31126, n31127, n31128, n31129,
         n31130, n31131, n31132, n31133, n31134, n31135, n31136, n31137,
         n31138, n31139, n31140, n31141, n31142, n31143, n31144, n31145,
         n31146, n31147, n31148, n31149, n31150, n31151, n31152, n31153,
         n31154, n31155, n31156, n31157, n31158, n31159, n31160, n31161,
         n31162, n31163, n31164, n31165, n31166, n31167, n31168, n31169,
         n31170, n31171, n31172, n31173, n31174, n31175, n31176, n31177,
         n31178, n31179, n31180, n31181, n31182, n31183, n31184, n31185,
         n31186, n31187, n31188, n31189, n31190, n31191, n31192, n31193,
         n31194, n31195, n31196, n31197, n31198, n31199, n31200, n31201,
         n31202, n31203, n31204, n31205, n31206, n31207, n31208, n31209,
         n31210, n31211, n31212, n31213, n31214, n31215, n31216, n31217,
         n31218, n31219, n31220, n31221, n31222, n31223, n31224, n31225,
         n31226, n31227, n31228, n31229, n31230, n31231, n31232, n31233,
         n31234, n31235, n31236, n31237, n31238, n31239, n31240, n31241,
         n31242, n31243, n31244, n31245, n31246, n31247, n31248, n31249,
         n31250, n31251, n31252, n31253, n31254, n31255, n31256, n31257,
         n31258, n31259, n31260, n31261, n31262, n31263, n31264, n31265,
         n31266, n31267, n31268, n31269, n31270, n31271, n31272, n31273,
         n31274, n31275, n31276, n31277, n31278, n31279, n31280, n31281,
         n31282, n31283, n31284, n31285, n31286, n31287, n31288, n31289,
         n31290, n31291, n31292, n31293, n31294, n31295, n31296, n31297,
         n31298, n31299, n31300, n31301, n31302, n31303, n31304, n31305,
         n31306, n31307, n31308, n31309, n31310, n31311, n31312, n31313,
         n31314, n31315, n31316, n31317, n31318, n31319, n31320, n31321,
         n31322, n31323, n31324, n31325, n31326, n31327, n31328, n31329,
         n31330, n31331, n31332, n31333, n31334, n31335, n31336, n31337,
         n31338, n31339, n31340, n31341, n31342, n31343, n31344, n31345,
         n31346, n31347, n31348, n31349, n31350, n31351, n31352, n31353,
         n31354, n31355, n31356, n31357, n31358, n31359, n31360, n31361,
         n31362, n31363, n31364, n31365, n31366, n31367, n31368, n31369,
         n31370, n31371, n31372, n31373, n31374, n31375, n31376, n31377,
         n31378, n31379, n31380, n31381, n31382, n31383, n31384, n31385,
         n31386, n31387, n31388, n31389, n31390, n31391, n31392, n31393,
         n31394, n31395, n31396, n31397, n31398, n31399, n31400, n31401,
         n31402, n31403, n31404, n31405, n31406, n31407, n31408, n31409,
         n31410, n31411, n31412, n31413, n31414, n31415, n31416, n31417,
         n31418, n31419, n31420, n31421, n31422, n31423, n31424, n31425,
         n31426, n31427, n31428, n31429, n31430, n31431, n31432, n31433,
         n31434, n31435, n31436, n31437, n31438, n31439, n31440, n31441,
         n31442, n31443, n31444, n31445, n31446, n31447, n31448, n31449,
         n31450, n31451, n31452, n31453, n31454, n31455, n31456, n31457,
         n31458, n31459, n31460, n31461, n31462, n31463, n31464, n31465,
         n31466, n31467, n31468, n31469, n31470, n31471, n31472, n31473,
         n31474, n31475, n31476, n31477, n31478, n31479, n31480, n31481,
         n31482, n31483, n31484, n31485, n31486, n31487, n31488, n31489,
         n31490, n31491, n31492, n31493, n31494, n31495, n31496, n31497,
         n31498, n31499, n31500, n31501, n31502, n31503, n31504, n31505,
         n31506, n31507, n31508, n31509, n31510, n31511, n31512, n31513,
         n31514, n31515, n31516, n31517, n31518, n31519, n31520, n31521,
         n31522, n31523, n31524, n31525, n31526, n31527, n31528, n31529,
         n31530, n31531, n31532, n31533, n31534, n31535, n31536, n31537,
         n31538, n31539, n31540, n31541, n31542, n31543, n31544, n31545,
         n31546, n31547, n31548, n31549, n31550, n31551, n31552, n31553,
         n31554, n31555, n31556, n31557, n31558, n31559, n31560, n31561,
         n31562, n31563, n31564, n31565, n31566, n31567, n31568, n31569,
         n31570, n31571, n31572, n31573, n31574, n31575, n31576, n31577,
         n31578, n31579, n31580, n31581, n31582, n31583, n31584, n31585,
         n31586, n31587, n31588, n31589, n31590, n31591, n31592, n31593,
         n31594, n31595, n31596, n31597, n31598, n31599, n31600, n31601,
         n31602, n31603, n31604, n31605, n31606, n31607, n31608, n31609,
         n31610, n31611, n31612, n31613, n31614, n31615, n31616, n31617,
         n31618, n31619, n31620, n31621, n31622, n31623, n31624, n31625,
         n31626, n31627, n31628, n31629, n31630, n31631, n31632, n31633,
         n31634, n31635, n31636, n31637, n31638, n31639, n31640, n31641,
         n31642, n31643, n31644, n31645, n31646, n31647, n31648, n31649,
         n31650, n31651, n31652, n31653, n31654, n31655, n31656, n31657,
         n31658, n31659, n31660, n31661, n31662, n31663, n31664, n31665,
         n31666, n31667, n31668, n31669, n31670, n31671, n31672, n31673,
         n31674, n31675, n31676, n31677, n31678, n31679, n31680, n31681,
         n31682, n31683, n31684, n31685, n31686, n31687, n31688, n31689,
         n31690, n31691, n31692, n31693, n31694, n31695, n31696, n31697,
         n31698, n31699, n31700, n31701, n31702, n31703, n31704, n31705,
         n31706, n31707, n31708, n31709, n31710, n31711, n31712, n31713,
         n31714, n31715, n31716, n31717, n31718, n31719, n31720, n31721,
         n31722, n31723, n31724, n31725, n31726, n31727, n31728, n31729,
         n31730, n31731, n31732, n31733, n31734, n31735, n31736, n31737,
         n31738, n31739, n31740, n31741, n31742, n31743, n31744, n31745,
         n31746, n31747, n31748, n31749, n31750, n31751, n31752, n31753,
         n31754, n31755, n31756, n31757, n31758, n31759, n31760, n31761,
         n31762, n31763, n31764, n31765, n31766, n31767, n31768, n31769,
         n31770, n31771, n31772, n31773, n31774, n31775, n31776, n31777,
         n31778, n31779, n31780, n31781, n31782, n31783, n31784, n31785,
         n31786, n31787, n31788, n31789, n31790, n31791, n31792, n31793,
         n31794, n31795, n31796, n31797, n31798, n31799, n31800, n31801,
         n31802, n31803, n31804, n31805, n31806, n31807, n31808, n31809,
         n31810, n31811, n31812, n31813, n31814, n31815, n31816, n31817,
         n31818, n31819, n31820, n31821, n31822, n31823, n31824, n31825,
         n31826, n31827, n31828, n31829, n31830, n31831, n31832, n31833,
         n31834, n31835, n31836, n31837, n31838, n31839, n31840, n31841,
         n31842, n31843, n31844, n31845, n31846, n31847, n31848, n31849,
         n31850, n31851, n31852, n31853, n31854, n31855, n31856, n31857,
         n31858, n31859, n31860, n31861, n31862, n31863, n31864, n31865,
         n31866, n31867, n31868, n31869, n31870, n31871, n31872, n31873,
         n31874, n31875, n31876, n31877, n31878, n31879, n31880, n31881,
         n31882, n31883, n31884, n31885, n31886, n31887, n31888, n31889,
         n31890, n31891, n31892, n31893, n31894, n31895, n31896, n31897,
         n31898, n31899, n31900, n31901, n31902, n31903, n31904, n31905,
         n31906, n31907, n31908, n31909, n31910, n31911, n31912, n31913,
         n31914, n31915, n31916, n31917, n31918, n31919, n31920, n31921,
         n31922, n31923, n31924, n31925, n31926, n31927, n31928, n31929,
         n31930, n31931, n31932, n31933, n31934, n31935, n31936, n31937,
         n31938, n31939, n31940, n31941, n31942, n31943, n31944, n31945,
         n31946, n31947, n31948, n31949, n31950, n31951, n31952, n31953,
         n31954, n31955, n31956, n31957, n31958, n31959, n31960, n31961,
         n31962, n31963, n31964, n31965, n31966, n31967, n31968, n31969,
         n31970, n31971, n31972, n31973, n31974, n31975, n31976, n31977,
         n31978, n31979, n31980, n31981, n31982, n31983, n31984, n31985,
         n31986, n31987, n31988, n31989, n31990, n31991, n31992, n31993,
         n31994, n31995, n31996, n31997, n31998, n31999, n32000, n32001,
         n32002, n32003, n32004, n32005, n32006, n32007, n32008, n32009,
         n32010, n32011, n32012, n32013, n32014, n32015, n32016, n32017,
         n32018, n32019, n32020, n32021, n32022, n32023, n32024, n32025,
         n32026, n32027, n32028, n32029, n32030, n32031, n32032, n32033,
         n32034, n32035, n32036, n32037, n32038, n32039, n32040, n32041,
         n32042, n32043, n32044, n32045, n32046, n32047, n32048, n32049,
         n32050, n32051, n32052, n32053, n32054, n32055, n32056, n32057,
         n32058, n32059, n32060, n32061, n32062, n32063, n32064, n32065,
         n32066, n32067, n32068, n32069, n32070, n32071, n32072, n32073,
         n32074, n32075, n32076, n32077, n32078, n32079, n32080, n32081,
         n32082, n32083, n32084, n32085, n32086, n32087, n32088, n32089,
         n32090, n32091, n32092, n32093, n32094, n32095, n32096, n32097,
         n32098, n32099, n32100, n32101, n32102, n32103, n32104, n32105,
         n32106, n32107, n32108, n32109, n32110, n32111, n32112, n32113,
         n32114, n32115, n32116, n32117, n32118, n32119, n32120, n32121,
         n32122, n32123, n32124, n32125, n32126, n32127, n32128, n32129,
         n32130, n32131, n32132, n32133, n32134, n32135, n32136, n32137,
         n32138, n32139, n32140, n32141, n32142, n32143, n32144, n32145,
         n32146, n32147, n32148, n32149, n32150, n32151, n32152, n32153,
         n32154, n32155, n32156, n32157, n32158, n32159, n32160, n32161,
         n32162, n32163, n32164, n32165, n32166, n32167, n32168, n32169,
         n32170, n32171, n32172, n32173, n32174, n32175, n32176, n32177,
         n32178, n32179, n32180, n32181, n32182, n32183, n32184, n32185,
         n32186, n32187, n32188, n32189, n32190, n32191, n32192, n32193,
         n32194, n32195, n32196, n32197, n32198, n32199, n32200, n32201,
         n32202, n32203, n32204, n32205, n32206, n32207, n32208, n32209,
         n32210, n32211, n32212, n32213, n32214, n32215, n32216, n32217,
         n32218, n32219, n32220, n32221, n32222, n32223, n32224, n32225,
         n32226, n32227, n32228, n32229, n32230, n32231, n32232, n32233,
         n32234, n32235, n32236, n32237, n32238, n32239, n32240, n32241,
         n32242, n32243, n32244, n32245, n32246, n32247, n32248, n32249,
         n32250, n32251, n32252, n32253, n32254, n32255, n32256, n32257,
         n32258, n32259, n32260, n32261, n32262, n32263, n32264, n32265,
         n32266, n32267, n32268, n32269, n32270, n32271, n32272, n32273,
         n32274, n32275, n32276, n32277, n32278, n32279, n32280, n32281,
         n32282, n32283, n32284, n32285, n32286, n32287, n32288, n32289,
         n32290, n32291, n32292, n32293, n32294, n32295, n32296, n32297,
         n32298, n32299, n32300, n32301, n32302, n32303, n32304, n32305,
         n32306, n32307, n32308, n32309, n32310, n32311, n32312, n32313,
         n32314, n32315, n32316, n32317, n32318, n32319, n32320, n32321,
         n32322, n32323, n32324, n32325, n32326, n32327, n32328, n32329,
         n32330, n32331, n32332, n32333, n32334, n32335, n32336, n32337,
         n32338, n32339, n32340, n32341, n32342, n32343, n32344, n32345,
         n32346, n32347, n32348, n32349, n32350, n32351, n32352, n32353,
         n32354, n32355, n32356, n32357, n32358, n32359, n32360, n32361,
         n32362, n32363, n32364, n32365, n32366, n32367, n32368, n32369,
         n32370, n32371, n32372, n32373, n32374, n32375, n32376, n32377,
         n32378, n32379, n32380, n32381, n32382, n32383, n32384, n32385,
         n32386, n32387, n32388, n32389, n32390, n32391, n32392, n32393,
         n32394, n32395, n32396, n32397, n32398, n32399, n32400, n32401,
         n32402, n32403, n32404, n32405, n32406, n32407, n32408, n32409,
         n32410, n32411, n32412, n32413, n32414, n32415, n32416, n32417,
         n32418, n32419, n32420, n32421, n32422, n32423, n32424, n32425,
         n32426, n32427, n32428, n32429, n32430, n32431, n32432, n32433,
         n32434, n32435, n32436, n32437, n32438, n32439, n32440, n32441,
         n32442, n32443, n32444, n32445, n32446, n32447, n32448, n32449,
         n32450, n32451, n32452, n32453, n32454, n32455, n32456, n32457,
         n32458, n32459, n32460, n32461, n32462, n32463, n32464, n32465,
         n32466, n32467, n32468, n32469, n32470, n32471, n32472, n32473,
         n32474, n32475, n32476, n32477, n32478, n32479, n32480, n32481,
         n32482, n32483, n32484, n32485, n32486, n32487, n32488, n32489,
         n32490, n32491, n32492, n32493, n32494, n32495, n32496, n32497,
         n32498, n32499, n32500, n32501, n32502, n32503, n32504, n32505,
         n32506, n32507, n32508, n32509, n32510, n32511, n32512, n32513,
         n32514, n32515, n32516, n32517, n32518, n32519, n32520, n32521,
         n32522, n32523, n32524, n32525, n32526, n32527, n32528, n32529,
         n32530, n32531, n32532, n32533, n32534, n32535, n32536, n32537,
         n32538, n32539, n32540, n32541, n32542, n32543, n32544, n32545,
         n32546, n32547, n32548, n32549, n32550, n32551, n32552, n32553,
         n32554, n32555, n32556, n32557, n32558, n32559, n32560, n32561,
         n32562, n32563, n32564, n32565, n32566, n32567, n32568, n32569,
         n32570, n32571, n32572, n32573, n32574, n32575, n32576, n32577,
         n32578, n32579, n32580, n32581, n32582, n32583, n32584, n32585,
         n32586, n32587, n32588, n32589, n32590, n32591, n32592, n32593,
         n32594, n32595, n32596, n32597, n32598, n32599, n32600, n32601,
         n32602, n32603, n32604, n32605, n32606, n32607, n32608, n32609,
         n32610, n32611, n32612, n32613, n32614, n32615, n32616, n32617,
         n32618, n32619, n32620, n32621, n32622, n32623, n32624, n32625,
         n32626, n32627, n32628, n32629, n32630, n32631, n32632, n32633,
         n32634, n32635, n32636, n32637, n32638, n32639, n32640, n32641,
         n32642, n32643, n32644, n32645, n32646, n32647, n32648, n32649,
         n32650, n32651, n32652, n32653, n32654, n32655, n32656, n32657,
         n32658, n32659, n32660, n32661, n32662, n32663, n32664, n32665,
         n32666, n32667, n32668, n32669, n32670, n32671, n32672, n32673,
         n32674, n32675, n32676, n32677, n32678, n32679, n32680, n32681,
         n32682, n32683, n32684, n32685, n32686, n32687, n32688, n32689,
         n32690, n32691, n32692, n32693, n32694, n32695, n32696, n32697,
         n32698, n32699, n32700, n32701, n32702, n32703, n32704, n32705,
         n32706, n32707, n32708, n32709, n32710, n32711, n32712, n32713,
         n32714, n32715, n32716, n32717, n32718, n32719, n32720, n32721,
         n32722, n32723, n32724, n32725, n32726, n32727, n32728, n32729,
         n32730, n32731, n32732, n32733, n32734, n32735, n32736, n32737,
         n32738, n32739, n32740, n32741, n32742, n32743, n32744, n32745,
         n32746, n32747, n32748, n32749, n32750, n32751, n32752, n32753,
         n32754, n32755, n32756, n32757, n32758, n32759, n32760, n32761,
         n32762, n32763, n32764, n32765, n32766, n32767, n32768, n32769,
         n32770, n32771, n32772, n32773, n32774, n32775, n32776, n32777,
         n32778, n32779, n32780, n32781, n32782, n32783, n32784, n32785,
         n32786, n32787, n32788, n32789, n32790, n32791, n32792, n32793,
         n32794, n32795, n32796, n32797, n32798, n32799, n32800, n32801,
         n32802, n32803, n32804, n32805, n32806, n32807, n32808, n32809,
         n32810, n32811, n32812, n32813, n32814, n32815, n32816, n32817,
         n32818, n32819, n32820, n32821, n32822, n32823, n32824, n32825,
         n32826, n32827, n32828, n32829, n32830, n32831, n32832, n32833,
         n32834, n32835, n32836, n32837, n32838, n32839, n32840, n32841,
         n32842, n32843, n32844, n32845, n32846, n32847, n32848, n32849,
         n32850, n32851, n32852, n32853, n32854, n32855, n32856, n32857,
         n32858, n32859, n32860, n32861, n32862, n32863, n32864, n32865,
         n32866, n32867, n32868, n32869, n32870, n32871, n32872, n32873,
         n32874, n32875, n32876, n32877, n32878, n32879, n32880, n32881,
         n32882, n32883, n32884, n32885, n32886, n32887, n32888, n32889,
         n32890, n32891, n32892, n32893, n32894, n32895, n32896, n32897,
         n32898, n32899, n32900, n32901, n32902, n32903, n32904, n32905,
         n32906, n32907, n32908, n32909, n32910, n32911, n32912, n32913,
         n32914, n32915, n32916, n32917, n32918, n32919, n32920, n32921,
         n32922, n32923, n32924, n32925, n32926, n32927, n32928, n32929,
         n32930, n32931, n32932, n32933, n32934, n32935, n32936, n32937,
         n32938, n32939, n32940, n32941, n32942, n32943, n32944, n32945,
         n32946, n32947, n32948, n32949, n32950, n32951, n32952, n32953,
         n32954, n32955, n32956, n32957, n32958, n32959, n32960, n32961,
         n32962, n32963, n32964, n32965, n32966, n32967, n32968, n32969,
         n32970, n32971, n32972, n32973, n32974, n32975, n32976, n32977,
         n32978, n32979, n32980, n32981, n32982, n32983, n32984, n32985,
         n32986, n32987, n32988, n32989, n32990, n32991, n32992, n32993,
         n32994, n32995, n32996, n32997, n32998, n32999, n33000, n33001,
         n33002, n33003, n33004, n33005, n33006, n33007, n33008, n33009,
         n33010, n33011, n33012, n33013, n33014, n33015, n33016, n33017,
         n33018, n33019, n33020, n33021, n33022, n33023, n33024, n33025,
         n33026, n33027, n33028, n33029, n33030, n33031, n33032, n33033,
         n33034, n33035, n33036, n33037, n33038, n33039, n33040, n33041,
         n33042, n33043, n33044, n33045, n33046, n33047, n33048, n33049,
         n33050, n33051, n33052, n33053, n33054, n33055, n33056, n33057,
         n33058, n33059, n33060, n33061, n33062, n33063, n33064, n33065,
         n33066, n33067, n33068, n33069, n33070, n33071, n33072, n33073,
         n33074, n33075, n33076, n33077, n33078, n33079, n33080, n33081,
         n33082, n33083, n33084, n33085, n33086, n33087, n33088, n33089,
         n33090, n33091, n33092, n33093, n33094, n33095, n33096, n33097,
         n33098, n33099, n33100, n33101, n33102, n33103, n33104, n33105,
         n33106, n33107, n33108, n33109, n33110, n33111, n33112, n33113,
         n33114, n33115, n33116, n33117, n33118, n33119, n33120, n33121,
         n33122, n33123, n33124, n33125, n33126, n33127, n33128, n33129,
         n33130, n33131, n33132, n33133, n33134, n33135, n33136, n33137,
         n33138, n33139, n33140, n33141, n33142, n33143, n33144, n33145,
         n33146, n33147, n33148, n33149, n33150, n33151, n33152, n33153,
         n33154, n33155, n33156, n33157, n33158, n33159, n33160, n33161,
         n33162, n33163, n33164, n33165, n33166, n33167, n33168, n33169,
         n33170, n33171, n33172, n33173, n33174, n33175, n33176, n33177,
         n33178, n33179, n33180, n33181, n33182, n33183, n33184, n33185,
         n33186, n33187, n33188, n33189, n33190, n33191, n33192, n33193,
         n33194, n33195, n33196, n33197, n33198, n33199, n33200, n33201,
         n33202, n33203, n33204, n33205, n33206, n33207, n33208, n33209,
         n33210, n33211, n33212, n33213, n33214, n33215, n33216, n33217,
         n33218, n33219, n33220, n33221, n33222, n33223, n33224, n33225,
         n33226, n33227, n33228, n33229, n33230, n33231, n33232, n33233,
         n33234, n33235, n33236, n33237, n33238, n33239, n33240, n33241,
         n33242, n33243, n33244, n33245, n33246, n33247, n33248, n33249,
         n33250, n33251, n33252, n33253, n33254, n33255, n33256, n33257,
         n33258, n33259, n33260, n33261, n33262, n33263, n33264, n33265,
         n33266, n33267, n33268, n33269, n33270, n33271, n33272, n33273,
         n33274, n33275, n33276, n33277, n33278, n33279, n33280, n33281,
         n33282, n33283, n33284, n33285, n33286, n33287, n33288, n33289,
         n33290, n33291, n33292, n33293, n33294, n33295, n33296, n33297,
         n33298, n33299, n33300, n33301, n33302, n33303, n33304, n33305,
         n33306, n33307, n33308, n33309, n33310, n33311, n33312, n33313,
         n33314, n33315, n33316, n33317, n33318, n33319, n33320, n33321,
         n33322, n33323, n33324, n33325, n33326, n33327, n33328, n33329,
         n33330, n33331, n33332, n33333, n33334, n33335, n33336, n33337,
         n33338, n33339, n33340, n33341, n33342, n33343, n33344, n33345,
         n33346, n33347, n33348, n33349, n33350, n33351, n33352, n33353,
         n33354, n33355, n33356, n33357, n33358, n33359, n33360, n33361,
         n33362, n33363, n33364, n33365, n33366, n33367, n33368, n33369,
         n33370, n33371, n33372, n33373, n33374, n33375, n33376, n33377,
         n33378, n33379, n33380, n33381, n33382, n33383, n33384, n33385,
         n33386, n33387, n33388, n33389, n33390, n33391, n33392, n33393,
         n33394, n33395, n33396, n33397, n33398, n33399, n33400, n33401,
         n33402, n33403, n33404, n33405, n33406, n33407, n33408, n33409,
         n33410, n33411, n33412, n33413, n33414, n33415, n33416, n33417,
         n33418, n33419, n33420, n33421, n33422, n33423, n33424, n33425,
         n33426, n33427, n33428, n33429, n33430, n33431, n33432, n33433,
         n33434, n33435, n33436, n33437, n33438, n33439, n33440, n33441,
         n33442, n33443, n33444, n33445, n33446, n33447, n33448, n33449,
         n33450, n33451, n33452, n33453, n33454, n33455, n33456, n33457,
         n33458, n33459, n33460, n33461, n33462, n33463, n33464, n33465,
         n33466, n33467, n33468, n33469, n33470, n33471, n33472, n33473,
         n33474, n33475, n33476, n33477, n33478, n33479, n33480, n33481,
         n33482, n33483, n33484, n33485, n33486, n33487, n33488, n33489,
         n33490, n33491, n33492, n33493, n33494, n33495, n33496, n33497,
         n33498, n33499, n33500, n33501, n33502, n33503, n33504, n33505,
         n33506, n33507, n33508, n33509, n33510, n33511, n33512, n33513,
         n33514, n33515, n33516, n33517, n33518, n33519, n33520, n33521,
         n33522, n33523, n33524, n33525, n33526, n33527, n33528, n33529,
         n33530, n33531, n33532, n33533, n33534, n33535, n33536, n33537,
         n33538, n33539, n33540, n33541, n33542, n33543, n33544, n33545,
         n33546, n33547, n33548, n33549, n33550, n33551, n33552, n33553,
         n33554, n33555, n33556, n33557, n33558, n33559, n33560, n33561,
         n33562, n33563, n33564, n33565, n33566, n33567, n33568, n33569,
         n33570, n33571, n33572, n33573, n33574, n33575, n33576, n33577,
         n33578, n33579, n33580, n33581, n33582, n33583, n33584, n33585,
         n33586, n33587, n33588, n33589, n33590, n33591, n33592, n33593,
         n33594, n33595, n33596, n33597, n33598, n33599, n33600, n33601,
         n33602, n33603, n33604, n33605, n33606, n33607, n33608, n33609,
         n33610, n33611, n33612, n33613, n33614, n33615, n33616, n33617,
         n33618, n33619, n33620, n33621, n33622, n33623, n33624, n33625,
         n33626, n33627, n33628, n33629, n33630, n33631, n33632, n33633,
         n33634, n33635, n33636, n33637, n33638, n33639, n33640, n33641,
         n33642, n33643, n33644, n33645, n33646, n33647, n33648, n33649,
         n33650, n33651, n33652, n33653, n33654, n33655, n33656, n33657,
         n33658, n33659, n33660, n33661, n33662, n33663, n33664, n33665,
         n33666, n33667, n33668, n33669, n33670, n33671, n33672, n33673,
         n33674, n33675, n33676, n33677, n33678, n33679, n33680, n33681,
         n33682, n33683, n33684, n33685, n33686, n33687, n33688, n33689,
         n33690, n33691, n33692, n33693, n33694, n33695, n33696, n33697,
         n33698, n33699, n33700, n33701, n33702, n33703, n33704, n33705,
         n33706, n33707, n33708, n33709, n33710, n33711, n33712, n33713,
         n33714, n33715, n33716, n33717, n33718, n33719, n33720, n33721,
         n33722, n33723, n33724, n33725, n33726, n33727, n33728, n33729,
         n33730, n33731, n33732, n33733, n33734, n33735, n33736, n33737,
         n33738, n33739, n33740, n33741, n33742, n33743, n33744, n33745,
         n33746, n33747, n33748, n33749, n33750, n33751, n33752, n33753,
         n33754, n33755, n33756, n33757, n33758, n33759, n33760, n33761,
         n33762, n33763, n33764, n33765, n33766, n33767, n33768, n33769,
         n33770, n33771, n33772, n33773, n33774, n33775, n33776, n33777,
         n33778, n33779, n33780, n33781, n33782, n33783, n33784, n33785,
         n33786, n33787, n33788, n33789, n33790, n33791, n33792, n33793,
         n33794, n33795, n33796, n33797, n33798, n33799, n33800, n33801,
         n33802, n33803, n33804, n33805, n33806, n33807, n33808, n33809,
         n33810, n33811, n33812, n33813, n33814, n33815, n33816, n33817,
         n33818, n33819, n33820, n33821, n33822, n33823, n33824, n33825,
         n33826, n33827, n33828, n33829, n33830, n33831, n33832, n33833,
         n33834, n33835, n33836, n33837, n33838, n33839, n33840, n33841,
         n33842, n33843, n33844, n33845, n33846, n33847, n33848, n33849,
         n33850, n33851, n33852, n33853, n33854, n33855, n33856, n33857,
         n33858, n33859, n33860, n33861, n33862, n33863, n33864, n33865,
         n33866, n33867, n33868, n33869, n33870, n33871, n33872, n33873,
         n33874, n33875, n33876, n33877, n33878, n33879, n33880, n33881,
         n33882, n33883, n33884, n33885, n33886, n33887, n33888, n33889,
         n33890, n33891, n33892, n33893, n33894, n33895, n33896, n33897,
         n33898, n33899, n33900, n33901, n33902, n33903, n33904, n33905,
         n33906, n33907, n33908, n33909, n33910, n33911, n33912, n33913,
         n33914, n33915, n33916, n33917, n33918, n33919, n33920, n33921,
         n33922, n33923, n33924, n33925, n33926, n33927, n33928, n33929,
         n33930, n33931, n33932, n33933, n33934, n33935, n33936, n33937,
         n33938, n33939, n33940, n33941, n33942, n33943, n33944, n33945,
         n33946, n33947, n33948, n33949, n33950, n33951, n33952, n33953,
         n33954, n33955, n33956, n33957, n33958, n33959, n33960, n33961,
         n33962, n33963, n33964, n33965, n33966, n33967, n33968, n33969,
         n33970, n33971, n33972, n33973, n33974, n33975, n33976, n33977,
         n33978, n33979, n33980, n33981, n33982, n33983, n33984, n33985,
         n33986, n33987, n33988, n33989, n33990, n33991, n33992, n33993,
         n33994, n33995, n33996, n33997, n33998, n33999, n34000, n34001,
         n34002, n34003, n34004, n34005, n34006, n34007, n34008, n34009,
         n34010, n34011, n34012, n34013, n34014, n34015, n34016, n34017,
         n34018, n34019, n34020, n34021, n34022, n34023, n34024, n34025,
         n34026, n34027, n34028, n34029, n34030, n34031, n34032, n34033,
         n34034, n34035, n34036, n34037, n34038, n34039, n34040, n34041,
         n34042, n34043, n34044, n34045, n34046, n34047, n34048, n34049,
         n34050, n34051, n34052, n34053, n34054, n34055, n34056, n34057,
         n34058, n34059, n34060, n34061, n34062, n34063, n34064, n34065,
         n34066, n34067, n34068, n34069, n34070, n34071, n34072, n34073,
         n34074, n34075, n34076, n34077, n34078, n34079, n34080, n34081,
         n34082, n34083, n34084, n34085, n34086, n34087, n34088, n34089,
         n34090, n34091, n34092, n34093, n34094, n34095, n34096, n34097,
         n34098, n34099, n34100, n34101, n34102, n34103, n34104, n34105,
         n34106, n34107, n34108, n34109, n34110, n34111, n34112, n34113,
         n34114, n34115, n34116, n34117, n34118, n34119, n34120, n34121,
         n34122, n34123, n34124, n34125, n34126, n34127, n34128, n34129,
         n34130, n34131, n34132, n34133, n34134, n34135, n34136, n34137,
         n34138, n34139, n34140, n34141, n34142, n34143, n34144, n34145,
         n34146, n34147, n34148, n34149, n34150, n34151, n34152, n34153,
         n34154, n34155, n34156, n34157, n34158, n34159, n34160, n34161,
         n34162, n34163, n34164, n34165, n34166, n34167, n34168, n34169,
         n34170, n34171, n34172, n34173, n34174, n34175, n34176, n34177,
         n34178, n34179, n34180, n34181, n34182, n34183, n34184, n34185,
         n34186, n34187, n34188, n34189, n34190, n34191, n34192, n34193,
         n34194, n34195, n34196, n34197, n34198, n34199, n34200, n34201,
         n34202, n34203, n34204, n34205, n34206, n34207, n34208, n34209,
         n34210, n34211, n34212, n34213, n34214, n34215, n34216, n34217,
         n34218, n34219, n34220, n34221, n34222, n34223, n34224, n34225,
         n34226, n34227, n34228, n34229, n34230, n34231, n34232, n34233,
         n34234, n34235, n34236, n34237, n34238, n34239, n34240, n34241,
         n34242, n34243, n34244, n34245, n34246, n34247, n34248, n34249,
         n34250, n34251, n34252, n34253, n34254, n34255, n34256, n34257,
         n34258, n34259, n34260, n34261, n34262, n34263, n34264, n34265,
         n34266, n34267, n34268, n34269, n34270, n34271, n34272, n34273,
         n34274, n34275, n34276, n34277, n34278, n34279, n34280, n34281,
         n34282, n34283, n34284, n34285, n34286, n34287, n34288, n34289,
         n34290, n34291, n34292, n34293, n34294, n34295, n34296, n34297,
         n34298, n34299, n34300, n34301, n34302, n34303, n34304, n34305,
         n34306, n34307, n34308, n34309, n34310, n34311, n34312, n34313,
         n34314, n34315, n34316, n34317, n34318, n34319, n34320, n34321,
         n34322, n34323, n34324, n34325, n34326, n34327, n34328, n34329,
         n34330, n34331, n34332, n34333, n34334, n34335, n34336, n34337,
         n34338, n34339, n34340, n34341, n34342, n34343, n34344, n34345,
         n34346, n34347, n34348, n34349, n34350, n34351, n34352, n34353,
         n34354, n34355, n34356, n34357, n34358, n34359, n34360, n34361,
         n34362, n34363, n34364, n34365, n34366, n34367, n34368, n34369,
         n34370, n34371, n34372, n34373, n34374, n34375, n34376, n34377,
         n34378, n34379, n34380, n34381, n34382, n34383, n34384, n34385,
         n34386, n34387, n34388, n34389, n34390, n34391, n34392, n34393,
         n34394, n34395, n34396, n34397, n34398, n34399, n34400, n34401,
         n34402, n34403, n34404, n34405, n34406, n34407, n34408, n34409,
         n34410, n34411, n34412, n34413, n34414, n34415, n34416, n34417,
         n34418, n34419, n34420, n34421, n34422, n34423, n34424, n34425,
         n34426, n34427, n34428, n34429, n34430, n34431, n34432, n34433,
         n34434, n34435, n34436, n34437, n34438, n34439, n34440, n34441,
         n34442, n34443, n34444, n34445, n34446, n34447, n34448, n34449,
         n34450, n34451, n34452, n34453, n34454, n34455, n34456, n34457,
         n34458, n34459, n34460, n34461, n34462, n34463, n34464, n34465,
         n34466, n34467, n34468, n34469, n34470, n34471, n34472, n34473,
         n34474, n34475, n34476, n34477, n34478, n34479, n34480, n34481,
         n34482, n34483, n34484, n34485, n34486, n34487, n34488, n34489,
         n34490, n34491, n34492, n34493, n34494, n34495, n34496, n34497,
         n34498, n34499, n34500, n34501, n34502, n34503, n34504, n34505,
         n34506, n34507, n34508, n34509, n34510, n34511, n34512, n34513,
         n34514, n34515, n34516, n34517, n34518, n34519, n34520, n34521,
         n34522, n34523, n34524, n34525, n34526, n34527, n34528, n34529,
         n34530, n34531, n34532, n34533, n34534, n34535, n34536, n34537,
         n34538, n34539, n34540, n34541, n34542, n34543, n34544, n34545,
         n34546, n34547, n34548, n34549, n34550, n34551, n34552, n34553,
         n34554, n34555, n34556, n34557, n34558, n34559, n34560, n34561,
         n34562, n34563, n34564, n34565, n34566, n34567, n34568, n34569,
         n34570, n34571, n34572, n34573, n34574, n34575, n34576, n34577,
         n34578, n34579, n34580, n34581, n34582, n34583, n34584, n34585,
         n34586, n34587, n34588, n34589, n34590, n34591, n34592, n34593,
         n34594, n34595, n34596, n34597, n34598, n34599, n34600, n34601,
         n34602, n34603, n34604, n34605, n34606, n34607, n34608, n34609,
         n34610, n34611, n34612, n34613, n34614, n34615, n34616, n34617,
         n34618, n34619, n34620, n34621, n34622, n34623, n34624, n34625,
         n34626, n34627, n34628, n34629, n34630, n34631, n34632, n34633,
         n34634, n34635, n34636, n34637, n34638, n34639, n34640, n34641,
         n34642, n34643, n34644, n34645, n34646, n34647, n34648, n34649,
         n34650, n34651, n34652, n34653, n34654, n34655, n34656, n34657,
         n34658, n34659, n34660, n34661, n34662, n34663, n34664, n34665,
         n34666, n34667, n34668, n34669, n34670, n34671, n34672, n34673,
         n34674, n34675, n34676, n34677, n34678, n34679, n34680, n34681,
         n34682, n34683, n34684, n34685, n34686, n34687, n34688, n34689,
         n34690, n34691, n34692, n34693, n34694, n34695, n34696, n34697,
         n34698, n34699, n34700, n34701, n34702, n34703, n34704, n34705,
         n34706, n34707, n34708, n34709, n34710, n34711, n34712, n34713,
         n34714, n34715, n34716, n34717, n34718, n34719, n34720, n34721,
         n34722, n34723, n34724, n34725, n34726, n34727, n34728, n34729,
         n34730, n34731, n34732, n34733, n34734, n34735, n34736, n34737,
         n34738, n34739, n34740, n34741, n34742, n34743, n34744, n34745,
         n34746, n34747, n34748, n34749, n34750, n34751, n34752, n34753,
         n34754, n34755, n34756, n34757, n34758, n34759, n34760, n34761,
         n34762, n34763, n34764, n34765, n34766, n34767, n34768, n34769,
         n34770, n34771, n34772, n34773, n34774, n34775, n34776, n34777,
         n34778, n34779, n34780, n34781, n34782, n34783, n34784, n34785,
         n34786, n34787, n34788, n34789, n34790, n34791, n34792, n34793,
         n34794, n34795, n34796, n34797, n34798, n34799, n34800, n34801,
         n34802, n34803, n34804, n34805, n34806, n34807, n34808, n34809,
         n34810, n34811, n34812, n34813, n34814, n34815, n34816, n34817,
         n34818, n34819, n34820, n34821, n34822, n34823, n34824, n34825,
         n34826, n34827, n34828, n34829, n34830, n34831, n34832, n34833,
         n34834, n34835, n34836, n34837, n34838, n34839, n34840, n34841,
         n34842, n34843, n34844, n34845, n34846, n34847, n34848, n34849,
         n34850, n34851, n34852, n34853, n34854, n34855, n34856, n34857,
         n34858, n34859, n34860, n34861, n34862, n34863, n34864, n34865,
         n34866, n34867, n34868, n34869, n34870, n34871, n34872, n34873,
         n34874, n34875, n34876, n34877, n34878, n34879, n34880, n34881,
         n34882, n34883, n34884, n34885, n34886, n34887, n34888, n34889,
         n34890, n34891, n34892, n34893, n34894, n34895, n34896, n34897,
         n34898, n34899, n34900, n34901, n34902, n34903, n34904, n34905,
         n34906, n34907, n34908, n34909, n34910, n34911, n34912, n34913,
         n34914, n34915, n34916, n34917, n34918, n34919, n34920, n34921,
         n34922, n34923, n34924, n34925, n34926, n34927, n34928, n34929,
         n34930, n34931, n34932, n34933, n34934, n34935, n34936, n34937,
         n34938, n34939, n34940, n34941, n34942, n34943, n34944, n34945,
         n34946, n34947, n34948, n34949, n34950, n34951, n34952, n34953,
         n34954, n34955, n34956, n34957, n34958, n34959, n34960, n34961,
         n34962, n34963, n34964, n34965, n34966, n34967, n34968, n34969,
         n34970, n34971, n34972, n34973, n34974, n34975, n34976, n34977,
         n34978, n34979, n34980, n34981, n34982, n34983, n34984, n34985,
         n34986, n34987, n34988, n34989, n34990, n34991, n34992, n34993,
         n34994, n34995, n34996, n34997, n34998, n34999, n35000, n35001,
         n35002, n35003, n35004, n35005, n35006, n35007, n35008, n35009,
         n35010, n35011, n35012, n35013, n35014, n35015, n35016, n35017,
         n35018, n35019, n35020, n35021, n35022, n35023, n35024, n35025,
         n35026, n35027, n35028, n35029, n35030, n35031, n35032, n35033,
         n35034, n35035, n35036, n35037, n35038, n35039, n35040, n35041,
         n35042, n35043, n35044, n35045, n35046, n35047, n35048, n35049,
         n35050, n35051, n35052, n35053, n35054, n35055, n35056, n35057,
         n35058, n35059, n35060, n35061, n35062, n35063, n35064, n35065,
         n35066, n35067, n35068, n35069, n35070, n35071, n35072, n35073,
         n35074, n35075, n35076, n35077, n35078, n35079, n35080, n35081,
         n35082, n35083, n35084, n35085, n35086, n35087, n35088, n35089,
         n35090, n35091, n35092, n35093, n35094, n35095, n35096, n35097,
         n35098, n35099, n35100, n35101, n35102, n35103, n35104, n35105,
         n35106, n35107, n35108, n35109, n35110, n35111, n35112, n35113,
         n35114, n35115, n35116, n35117, n35118, n35119, n35120, n35121,
         n35122, n35123, n35124, n35125, n35126, n35127, n35128, n35129,
         n35130, n35131, n35132, n35133, n35134, n35135, n35136, n35137,
         n35138, n35139, n35140, n35141, n35142, n35143, n35144, n35145,
         n35146, n35147, n35148, n35149, n35150, n35151, n35152, n35153,
         n35154, n35155, n35156, n35157, n35158, n35159, n35160, n35161,
         n35162, n35163, n35164, n35165, n35166, n35167, n35168, n35169,
         n35170, n35171, n35172, n35173, n35174, n35175, n35176, n35177,
         n35178, n35179, n35180, n35181, n35182, n35183, n35184, n35185,
         n35186, n35187, n35188, n35189, n35190, n35191, n35192, n35193,
         n35194, n35195, n35196, n35197, n35198, n35199, n35200, n35201,
         n35202, n35203, n35204, n35205, n35206, n35207, n35208, n35209,
         n35210, n35211, n35212, n35213, n35214, n35215, n35216, n35217,
         n35218, n35219, n35220, n35221, n35222, n35223, n35224, n35225,
         n35226, n35227, n35228, n35229, n35230, n35231, n35232, n35233,
         n35234, n35235, n35236, n35237, n35238, n35239, n35240, n35241,
         n35242, n35243, n35244, n35245, n35246, n35247, n35248, n35249,
         n35250, n35251, n35252, n35253, n35254, n35255, n35256, n35257,
         n35258, n35259, n35260, n35261, n35262, n35263, n35264, n35265,
         n35266, n35267, n35268, n35269, n35270, n35271, n35272, n35273,
         n35274, n35275, n35276, n35277, n35278, n35279, n35280, n35281,
         n35282, n35283, n35284, n35285, n35286, n35287, n35288, n35289,
         n35290, n35291, n35292, n35293, n35294, n35295, n35296, n35297,
         n35298, n35299, n35300, n35301, n35302, n35303, n35304, n35305,
         n35306, n35307, n35308, n35309, n35310, n35311, n35312, n35313,
         n35314, n35315, n35316, n35317, n35318, n35319, n35320, n35321,
         n35322, n35323, n35324, n35325, n35326, n35327, n35328, n35329,
         n35330, n35331, n35332, n35333, n35334, n35335, n35336, n35337,
         n35338, n35339, n35340, n35341, n35342, n35343, n35344, n35345,
         n35346, n35347, n35348, n35349, n35350, n35351, n35352, n35353,
         n35354, n35355, n35356, n35357, n35358, n35359, n35360, n35361,
         n35362, n35363, n35364, n35365, n35366, n35367, n35368, n35369,
         n35370, n35371, n35372, n35373, n35374, n35375, n35376, n35377,
         n35378, n35379, n35380, n35381, n35382, n35383, n35384, n35385,
         n35386, n35387, n35388, n35389, n35390, n35391, n35392, n35393,
         n35394, n35395, n35396, n35397, n35398, n35399, n35400, n35401,
         n35402, n35403, n35404, n35405, n35406, n35407, n35408, n35409,
         n35410, n35411, n35412, n35413, n35414, n35415, n35416, n35417,
         n35418, n35419, n35420, n35421, n35422, n35423, n35424, n35425,
         n35426, n35427, n35428, n35429, n35430, n35431, n35432, n35433,
         n35434, n35435, n35436, n35437, n35438, n35439, n35440, n35441,
         n35442, n35443, n35444, n35445, n35446, n35447, n35448, n35449,
         n35450, n35451, n35452, n35453, n35454, n35455, n35456, n35457,
         n35458, n35459, n35460, n35461, n35462, n35463, n35464, n35465,
         n35466, n35467, n35468, n35469, n35470, n35471, n35472, n35473,
         n35474, n35475, n35476, n35477, n35478, n35479, n35480, n35481,
         n35482, n35483, n35484, n35485, n35486, n35487, n35488, n35489,
         n35490, n35491, n35492, n35493, n35494, n35495, n35496, n35497,
         n35498, n35499, n35500, n35501, n35502, n35503, n35504, n35505,
         n35506, n35507, n35508, n35509, n35510, n35511, n35512, n35513,
         n35514, n35515, n35516, n35517, n35518, n35519, n35520, n35521,
         n35522, n35523, n35524, n35525, n35526, n35527, n35528, n35529,
         n35530, n35531, n35532, n35533, n35534, n35535, n35536, n35537,
         n35538, n35539, n35540, n35541, n35542, n35543, n35544, n35545,
         n35546, n35547, n35548, n35549, n35550, n35551, n35552, n35553,
         n35554, n35555, n35556, n35557, n35558, n35559, n35560, n35561,
         n35562, n35563, n35564, n35565, n35566, n35567, n35568, n35569,
         n35570, n35571, n35572, n35573, n35574, n35575, n35576, n35577,
         n35578, n35579, n35580, n35581, n35582, n35583, n35584, n35585,
         n35586, n35587, n35588, n35589, n35590, n35591, n35592, n35593,
         n35594, n35595, n35596, n35597, n35598, n35599, n35600, n35601,
         n35602, n35603, n35604, n35605, n35606, n35607, n35608, n35609,
         n35610, n35611, n35612, n35613, n35614, n35615, n35616, n35617,
         n35618, n35619, n35620, n35621, n35622, n35623, n35624, n35625,
         n35626, n35627, n35628, n35629, n35630, n35631, n35632, n35633,
         n35634, n35635, n35636, n35637, n35638, n35639, n35640, n35641,
         n35642, n35643, n35644, n35645, n35646, n35647, n35648, n35649,
         n35650, n35651, n35652, n35653, n35654, n35655, n35656, n35657,
         n35658, n35659, n35660, n35661, n35662, n35663, n35664, n35665,
         n35666, n35667, n35668, n35669, n35670, n35671, n35672, n35673,
         n35674, n35675, n35676, n35677, n35678, n35679, n35680, n35681,
         n35682, n35683, n35684, n35685, n35686, n35687, n35688, n35689,
         n35690, n35691, n35692, n35693, n35694, n35695, n35696, n35697,
         n35698, n35699, n35700, n35701, n35702, n35703, n35704, n35705,
         n35706, n35707, n35708, n35709, n35710, n35711, n35712, n35713,
         n35714, n35715, n35716, n35717, n35718, n35719, n35720, n35721,
         n35722, n35723, n35724, n35725, n35726, n35727, n35728, n35729,
         n35730, n35731, n35732, n35733, n35734, n35735, n35736, n35737,
         n35738, n35739, n35740, n35741, n35742, n35743, n35744, n35745,
         n35746, n35747, n35748, n35749, n35750, n35751, n35752, n35753,
         n35754, n35755, n35756, n35757, n35758, n35759, n35760, n35761,
         n35762, n35763, n35764, n35765, n35766, n35767, n35768, n35769,
         n35770, n35771, n35772, n35773, n35774, n35775, n35776, n35777,
         n35778, n35779, n35780, n35781, n35782, n35783, n35784, n35785,
         n35786, n35787, n35788, n35789, n35790, n35791, n35792, n35793,
         n35794, n35795, n35796, n35797, n35798, n35799, n35800, n35801,
         n35802, n35803, n35804, n35805, n35806, n35807, n35808, n35809,
         n35810, n35811, n35812, n35813, n35814, n35815, n35816, n35817,
         n35818, n35819, n35820, n35821, n35822, n35823, n35824, n35825,
         n35826, n35827, n35828, n35829, n35830, n35831, n35832, n35833,
         n35834, n35835, n35836, n35837, n35838, n35839, n35840, n35841,
         n35842, n35843, n35844, n35845, n35846, n35847, n35848, n35849,
         n35850, n35851, n35852, n35853, n35854, n35855, n35856, n35857,
         n35858, n35859, n35860, n35861, n35862, n35863, n35864, n35865,
         n35866, n35867, n35868, n35869, n35870, n35871, n35872, n35873,
         n35874, n35875, n35876, n35877, n35878, n35879, n35880, n35881,
         n35882, n35883, n35884, n35885, n35886, n35887, n35888, n35889,
         n35890, n35891, n35892, n35893, n35894, n35895, n35896, n35897,
         n35898, n35899, n35900, n35901, n35902, n35903, n35904, n35905,
         n35906, n35907, n35908, n35909, n35910, n35911, n35912, n35913,
         n35914, n35915, n35916, n35917, n35918, n35919, n35920, n35921,
         n35922, n35923, n35924, n35925, n35926, n35927, n35928, n35929,
         n35930, n35931, n35932, n35933, n35934, n35935, n35936, n35937,
         n35938, n35939, n35940, n35941, n35942, n35943, n35944, n35945,
         n35946, n35947, n35948, n35949, n35950, n35951, n35952, n35953,
         n35954, n35955, n35956, n35957, n35958, n35959, n35960, n35961,
         n35962, n35963, n35964, n35965, n35966, n35967, n35968, n35969,
         n35970, n35971, n35972, n35973, n35974, n35975, n35976, n35977,
         n35978, n35979, n35980, n35981, n35982, n35983, n35984, n35985,
         n35986, n35987, n35988, n35989, n35990, n35991, n35992, n35993,
         n35994, n35995, n35996, n35997, n35998, n35999, n36000, n36001,
         n36002, n36003, n36004, n36005, n36006, n36007, n36008, n36009,
         n36010, n36011, n36012, n36013, n36014, n36015, n36016, n36017,
         n36018, n36019, n36020, n36021, n36022, n36023, n36024, n36025,
         n36026, n36027, n36028, n36029, n36030, n36031, n36032, n36033,
         n36034, n36035, n36036, n36037, n36038, n36039, n36040, n36041,
         n36042, n36043, n36044, n36045, n36046, n36047, n36048, n36049,
         n36050, n36051, n36052, n36053, n36054, n36055, n36056, n36057,
         n36058, n36059, n36060, n36061, n36062, n36063, n36064, n36065,
         n36066, n36067, n36068, n36069, n36070, n36071, n36072, n36073,
         n36074, n36075, n36076, n36077, n36078, n36079, n36080, n36081,
         n36082, n36083, n36084, n36085, n36086, n36087, n36088, n36089,
         n36090, n36091, n36092, n36093, n36094, n36095, n36096, n36097,
         n36098, n36099, n36100, n36101, n36102, n36103, n36104, n36105,
         n36106, n36107, n36108, n36109, n36110, n36111, n36112, n36113,
         n36114, n36115, n36116, n36117, n36118, n36119, n36120, n36121,
         n36122, n36123, n36124, n36125, n36126, n36127, n36128, n36129,
         n36130, n36131, n36132, n36133, n36134, n36135, n36136, n36137,
         n36138, n36139, n36140, n36141, n36142, n36143, n36144, n36145,
         n36146, n36147, n36148, n36149, n36150, n36151, n36152, n36153,
         n36154, n36155, n36156, n36157, n36158, n36159, n36160, n36161,
         n36162, n36163, n36164, n36165, n36166, n36167, n36168, n36169,
         n36170, n36171, n36172, n36173, n36174, n36175, n36176, n36177,
         n36178, n36179, n36180, n36181, n36182, n36183, n36184, n36185,
         n36186, n36187, n36188, n36189, n36190, n36191, n36192, n36193,
         n36194, n36195, n36196, n36197, n36198, n36199, n36200, n36201,
         n36202, n36203, n36204, n36205, n36206, n36207, n36208, n36209,
         n36210, n36211, n36212, n36213, n36214, n36215, n36216, n36217,
         n36218, n36219, n36220, n36221, n36222, n36223, n36224, n36225,
         n36226, n36227, n36228, n36229, n36230, n36231, n36232, n36233,
         n36234, n36235, n36236, n36237, n36238, n36239, n36240, n36241,
         n36242, n36243, n36244, n36245, n36246, n36247, n36248, n36249,
         n36250, n36251, n36252, n36253, n36254, n36255, n36256, n36257,
         n36258, n36259, n36260, n36261, n36262, n36263, n36264, n36265,
         n36266, n36267, n36268, n36269, n36270, n36271, n36272, n36273,
         n36274, n36275, n36276, n36277, n36278, n36279, n36280, n36281,
         n36282, n36283, n36284, n36285, n36286, n36287, n36288, n36289,
         n36290, n36291, n36292, n36293, n36294, n36295, n36296, n36297,
         n36298, n36299, n36300, n36301, n36302, n36303, n36304, n36305,
         n36306, n36307, n36308, n36309, n36310, n36311, n36312, n36313,
         n36314, n36315, n36316, n36317, n36318, n36319, n36320, n36321,
         n36322, n36323, n36324, n36325, n36326, n36327, n36328, n36329,
         n36330, n36331, n36332, n36333, n36334, n36335, n36336, n36337,
         n36338, n36339, n36340, n36341, n36342, n36343, n36344, n36345,
         n36346, n36347, n36348, n36349, n36350, n36351, n36352, n36353,
         n36354, n36355, n36356, n36357, n36358, n36359, n36360, n36361,
         n36362, n36363, n36364, n36365, n36366, n36367, n36368, n36369,
         n36370, n36371, n36372, n36373, n36374, n36375, n36376, n36377,
         n36378, n36379, n36380, n36381, n36382, n36383, n36384, n36385,
         n36386, n36387, n36388, n36389, n36390, n36391, n36392, n36393,
         n36394, n36395, n36396, n36397, n36398, n36399, n36400, n36401,
         n36402, n36403, n36404, n36405, n36406, n36407, n36408, n36409,
         n36410, n36411, n36412, n36413, n36414, n36415, n36416, n36417,
         n36418, n36419, n36420, n36421, n36422, n36423, n36424, n36425,
         n36426, n36427, n36428, n36429, n36430, n36431, n36432, n36433,
         n36434, n36435, n36436, n36437, n36438, n36439, n36440, n36441,
         n36442, n36443, n36444, n36445, n36446, n36447, n36448, n36449,
         n36450, n36451, n36452, n36453, n36454, n36455, n36456, n36457,
         n36458, n36459, n36460, n36461, n36462, n36463, n36464, n36465,
         n36466, n36467, n36468, n36469, n36470, n36471, n36472, n36473,
         n36474, n36475, n36476, n36477, n36478, n36479, n36480, n36481,
         n36482, n36483, n36484, n36485, n36486, n36487, n36488, n36489,
         n36490, n36491, n36492, n36493, n36494, n36495, n36496, n36497,
         n36498, n36499, n36500, n36501, n36502, n36503, n36504, n36505,
         n36506, n36507, n36508, n36509, n36510, n36511, n36512, n36513,
         n36514, n36515, n36516, n36517, n36518, n36519, n36520, n36521,
         n36522, n36523, n36524, n36525, n36526, n36527, n36528, n36529,
         n36530, n36531, n36532, n36533, n36534, n36535, n36536, n36537,
         n36538, n36539, n36540, n36541, n36542, n36543, n36544, n36545,
         n36546, n36547, n36548, n36549, n36550, n36551, n36552, n36553,
         n36554, n36555, n36556, n36557, n36558, n36559, n36560, n36561,
         n36562, n36563, n36564, n36565, n36566, n36567, n36568, n36569,
         n36570, n36571, n36572, n36573, n36574, n36575, n36576, n36577,
         n36578, n36579, n36580, n36581, n36582, n36583, n36584, n36585,
         n36586, n36587, n36588, n36589, n36590, n36591, n36592, n36593,
         n36594, n36595, n36596, n36597, n36598, n36599, n36600, n36601,
         n36602, n36603, n36604, n36605, n36606, n36607, n36608, n36609,
         n36610, n36611, n36612, n36613, n36614, n36615, n36616, n36617,
         n36618, n36619, n36620, n36621, n36622, n36623, n36624, n36625,
         n36626, n36627, n36628, n36629, n36630, n36631, n36632, n36633,
         n36634, n36635, n36636, n36637, n36638, n36639, n36640, n36641,
         n36642, n36643, n36644, n36645, n36646, n36647, n36648, n36649,
         n36650, n36651, n36652, n36653, n36654, n36655, n36656, n36657,
         n36658, n36659, n36660, n36661, n36662, n36663, n36664, n36665,
         n36666, n36667, n36668, n36669, n36670, n36671, n36672, n36673,
         n36674, n36675, n36676, n36677, n36678, n36679, n36680, n36681,
         n36682, n36683, n36684, n36685, n36686, n36687, n36688, n36689,
         n36690, n36691, n36692, n36693, n36694, n36695, n36696, n36697,
         n36698, n36699, n36700, n36701, n36702, n36703, n36704, n36705,
         n36706, n36707, n36708, n36709, n36710, n36711, n36712, n36713,
         n36714, n36715, n36716, n36717, n36718, n36719, n36720, n36721,
         n36722, n36723, n36724, n36725, n36726, n36727, n36728, n36729,
         n36730, n36731, n36732, n36733, n36734, n36735, n36736, n36737,
         n36738, n36739, n36740, n36741, n36742, n36743, n36744, n36745,
         n36746, n36747, n36748, n36749, n36750, n36751, n36752, n36753,
         n36754, n36755, n36756, n36757, n36758, n36759, n36760, n36761,
         n36762, n36763, n36764, n36765, n36766, n36767, n36768, n36769,
         n36770, n36771, n36772, n36773, n36774, n36775, n36776, n36777,
         n36778, n36779, n36780, n36781, n36782, n36783, n36784, n36785,
         n36786, n36787, n36788, n36789, n36790, n36791, n36792, n36793,
         n36794, n36795, n36796, n36797, n36798, n36799, n36800, n36801,
         n36802, n36803, n36804, n36805, n36806, n36807, n36808, n36809,
         n36810, n36811, n36812, n36813, n36814, n36815, n36816, n36817,
         n36818, n36819, n36820, n36821, n36822, n36823, n36824, n36825,
         n36826, n36827, n36828, n36829, n36830, n36831, n36832, n36833,
         n36834, n36835, n36836, n36837, n36838, n36839, n36840, n36841,
         n36842, n36843, n36844, n36845, n36846, n36847, n36848, n36849,
         n36850, n36851, n36852, n36853, n36854, n36855, n36856, n36857,
         n36858, n36859, n36860, n36861, n36862, n36863, n36864, n36865,
         n36866, n36867, n36868, n36869, n36870, n36871, n36872, n36873,
         n36874, n36875, n36876, n36877, n36878, n36879, n36880, n36881,
         n36882, n36883, n36884, n36885, n36886, n36887, n36888, n36889,
         n36890, n36891, n36892, n36893, n36894, n36895, n36896, n36897,
         n36898, n36899, n36900, n36901, n36902, n36903, n36904, n36905,
         n36906, n36907, n36908, n36909, n36910, n36911, n36912, n36913,
         n36914, n36915, n36916, n36917, n36918, n36919, n36920, n36921,
         n36922, n36923, n36924, n36925, n36926, n36927, n36928, n36929,
         n36930, n36931, n36932, n36933, n36934, n36935, n36936, n36937,
         n36938, n36939, n36940, n36941, n36942, n36943, n36944, n36945,
         n36946, n36947, n36948, n36949, n36950, n36951, n36952, n36953,
         n36954, n36955, n36956, n36957, n36958, n36959, n36960, n36961,
         n36962, n36963, n36964, n36965, n36966, n36967, n36968, n36969,
         n36970, n36971, n36972, n36973, n36974, n36975, n36976, n36977,
         n36978, n36979, n36980, n36981, n36982, n36983, n36984, n36985,
         n36986, n36987, n36988, n36989, n36990, n36991, n36992, n36993,
         n36994, n36995, n36996, n36997, n36998, n36999, n37000, n37001,
         n37002, n37003, n37004, n37005, n37006, n37007, n37008, n37009,
         n37010, n37011, n37012, n37013, n37014, n37015, n37016, n37017,
         n37018, n37019, n37020, n37021, n37022, n37023, n37024, n37025,
         n37026, n37027, n37028, n37029, n37030, n37031, n37032, n37033,
         n37034, n37035, n37036, n37037, n37038, n37039, n37040, n37041,
         n37042, n37043, n37044, n37045, n37046, n37047, n37048, n37049,
         n37050, n37051, n37052, n37053, n37054, n37055, n37056, n37057,
         n37058, n37059, n37060, n37061, n37062, n37063, n37064, n37065,
         n37066, n37067, n37068, n37069, n37070, n37071, n37072, n37073,
         n37074, n37075, n37076, n37077, n37078, n37079, n37080, n37081,
         n37082, n37083, n37084, n37085, n37086, n37087, n37088, n37089,
         n37090, n37091, n37092, n37093, n37094, n37095, n37096, n37097,
         n37098, n37099, n37100, n37101, n37102, n37103, n37104, n37105,
         n37106, n37107, n37108, n37109, n37110, n37111, n37112, n37113,
         n37114, n37115, n37116, n37117, n37118, n37119, n37120, n37121,
         n37122, n37123, n37124, n37125, n37126, n37127, n37128, n37129,
         n37130, n37131, n37132, n37133, n37134, n37135, n37136, n37137,
         n37138, n37139, n37140, n37141, n37142, n37143, n37144, n37145,
         n37146, n37147, n37148, n37149, n37150, n37151, n37152, n37153,
         n37154, n37155, n37156, n37157, n37158, n37159, n37160, n37161,
         n37162, n37163, n37164, n37165, n37166, n37167, n37168, n37169,
         n37170, n37171, n37172, n37173, n37174, n37175, n37176, n37177,
         n37178, n37179, n37180, n37181, n37182, n37183, n37184, n37185,
         n37186, n37187, n37188, n37189, n37190, n37191, n37192, n37193,
         n37194, n37195, n37196, n37197, n37198, n37199, n37200, n37201,
         n37202, n37203, n37204, n37205, n37206, n37207, n37208, n37209,
         n37210, n37211, n37212, n37213, n37214, n37215, n37216, n37217,
         n37218, n37219, n37220, n37221, n37222, n37223, n37224, n37225,
         n37226, n37227, n37228, n37229, n37230, n37231, n37232, n37233,
         n37234, n37235, n37236, n37237, n37238, n37239, n37240, n37241,
         n37242, n37243, n37244, n37245, n37246, n37247, n37248, n37249,
         n37250, n37251, n37252, n37253, n37254, n37255, n37256, n37257,
         n37258, n37259, n37260, n37261, n37262, n37263, n37264, n37265,
         n37266, n37267, n37268, n37269, n37270, n37271, n37272, n37273,
         n37274, n37275, n37276, n37277, n37278, n37279, n37280, n37281,
         n37282, n37283, n37284, n37285, n37286, n37287, n37288, n37289,
         n37290, n37291, n37292, n37293, n37294, n37295, n37296, n37297,
         n37298, n37299, n37300, n37301, n37302, n37303, n37304, n37305,
         n37306, n37307, n37308, n37309, n37310, n37311, n37312, n37313,
         n37314, n37315, n37316, n37317, n37318, n37319, n37320, n37321,
         n37322, n37323, n37324, n37325, n37326, n37327, n37328, n37329,
         n37330, n37331, n37332, n37333, n37334, n37335, n37336, n37337,
         n37338, n37339, n37340, n37341, n37342, n37343, n37344, n37345,
         n37346, n37347, n37348, n37349, n37350, n37351, n37352, n37353,
         n37354, n37355, n37356, n37357, n37358, n37359, n37360, n37361,
         n37362, n37363, n37364, n37365, n37366, n37367, n37368, n37369,
         n37370, n37371, n37372, n37373, n37374, n37375, n37376, n37377,
         n37378, n37379, n37380, n37381, n37382, n37383, n37384, n37385,
         n37386, n37387, n37388, n37389, n37390, n37391, n37392, n37393,
         n37394, n37395, n37396, n37397, n37398, n37399, n37400, n37401,
         n37402, n37403, n37404, n37405, n37406, n37407, n37408, n37409,
         n37410, n37411, n37412, n37413, n37414, n37415, n37416, n37417,
         n37418, n37419, n37420, n37421, n37422, n37423, n37424, n37425,
         n37426, n37427, n37428, n37429, n37430, n37431, n37432, n37433,
         n37434, n37435, n37436, n37437, n37438, n37439, n37440, n37441,
         n37442, n37443, n37444, n37445, n37446, n37447, n37448, n37449,
         n37450, n37451, n37452, n37453, n37454, n37455, n37456, n37457,
         n37458, n37459, n37460, n37461, n37462, n37463, n37464, n37465,
         n37466, n37467, n37468, n37469, n37470, n37471, n37472, n37473,
         n37474, n37475, n37476, n37477, n37478, n37479, n37480, n37481,
         n37482, n37483, n37484, n37485, n37486, n37487, n37488, n37489,
         n37490, n37491, n37492, n37493, n37494, n37495, n37496, n37497,
         n37498, n37499, n37500, n37501, n37502, n37503, n37504, n37505,
         n37506, n37507, n37508, n37509, n37510, n37511, n37512, n37513,
         n37514, n37515, n37516, n37517, n37518, n37519, n37520, n37521,
         n37522, n37523, n37524, n37525, n37526, n37527, n37528, n37529,
         n37530, n37531, n37532, n37533, n37534, n37535, n37536, n37537,
         n37538, n37539, n37540, n37541, n37542, n37543, n37544, n37545,
         n37546, n37547, n37548, n37549, n37550, n37551, n37552, n37553,
         n37554, n37555, n37556, n37557, n37558, n37559, n37560, n37561,
         n37562, n37563, n37564, n37565, n37566, n37567, n37568, n37569,
         n37570, n37571, n37572, n37573, n37574, n37575, n37576, n37577,
         n37578, n37579, n37580, n37581, n37582, n37583, n37584, n37585,
         n37586, n37587, n37588, n37589, n37590, n37591, n37592, n37593,
         n37594, n37595, n37596, n37597, n37598, n37599, n37600, n37601,
         n37602, n37603, n37604, n37605, n37606, n37607, n37608, n37609,
         n37610, n37611, n37612, n37613, n37614, n37615, n37616, n37617,
         n37618, n37619, n37620, n37621, n37622, n37623, n37624, n37625,
         n37626, n37627, n37628, n37629, n37630, n37631, n37632, n37633,
         n37634, n37635, n37636, n37637, n37638, n37639, n37640, n37641,
         n37642, n37643, n37644, n37645, n37646, n37647, n37648, n37649,
         n37650, n37651, n37652, n37653, n37654, n37655, n37656, n37657,
         n37658, n37659, n37660, n37661, n37662, n37663, n37664, n37665,
         n37666, n37667, n37668, n37669, n37670, n37671, n37672, n37673,
         n37674, n37675, n37676, n37677, n37678, n37679, n37680, n37681,
         n37682, n37683, n37684, n37685, n37686, n37687, n37688, n37689,
         n37690, n37691, n37692, n37693, n37694, n37695, n37696, n37697,
         n37698, n37699, n37700, n37701, n37702, n37703, n37704, n37705,
         n37706, n37707, n37708, n37709, n37710, n37711, n37712, n37713,
         n37714, n37715, n37716, n37717, n37718, n37719, n37720, n37721,
         n37722, n37723, n37724, n37725, n37726, n37727, n37728, n37729,
         n37730, n37731, n37732, n37733, n37734, n37735, n37736, n37737,
         n37738, n37739, n37740, n37741, n37742, n37743, n37744, n37745,
         n37746, n37747, n37748, n37749, n37750, n37751, n37752, n37753,
         n37754, n37755, n37756, n37757, n37758, n37759, n37760, n37761,
         n37762, n37763, n37764, n37765, n37766, n37767, n37768, n37769,
         n37770, n37771, n37772, n37773, n37774, n37775, n37776, n37777,
         n37778, n37779, n37780, n37781, n37782, n37783, n37784, n37785,
         n37786, n37787, n37788, n37789, n37790, n37791, n37792, n37793,
         n37794, n37795, n37796, n37797, n37798, n37799, n37800, n37801,
         n37802, n37803, n37804, n37805, n37806, n37807, n37808, n37809,
         n37810, n37811, n37812, n37813, n37814, n37815, n37816, n37817,
         n37818, n37819, n37820, n37821, n37822, n37823, n37824, n37825,
         n37826, n37827, n37828, n37829, n37830, n37831, n37832, n37833,
         n37834, n37835, n37836, n37837, n37838, n37839, n37840, n37841,
         n37842, n37843, n37844, n37845, n37846, n37847, n37848, n37849,
         n37850, n37851, n37852, n37853, n37854, n37855, n37856, n37857,
         n37858, n37859, n37860, n37861, n37862, n37863, n37864, n37865,
         n37866, n37867, n37868, n37869, n37870, n37871, n37872, n37873,
         n37874, n37875, n37876, n37877, n37878, n37879, n37880, n37881,
         n37882, n37883, n37884, n37885, n37886, n37887, n37888, n37889,
         n37890, n37891, n37892, n37893, n37894, n37895, n37896, n37897,
         n37898, n37899, n37900, n37901, n37902, n37903, n37904, n37905,
         n37906, n37907, n37908, n37909, n37910, n37911, n37912, n37913,
         n37914, n37915, n37916, n37917, n37918, n37919, n37920, n37921,
         n37922, n37923, n37924, n37925, n37926, n37927, n37928, n37929,
         n37930, n37931, n37932, n37933, n37934, n37935, n37936, n37937,
         n37938, n37939, n37940, n37941, n37942, n37943, n37944, n37945,
         n37946, n37947, n37948, n37949, n37950, n37951, n37952, n37953,
         n37954, n37955, n37956, n37957, n37958, n37959, n37960, n37961,
         n37962, n37963, n37964, n37965, n37966, n37967, n37968, n37969,
         n37970, n37971, n37972, n37973, n37974, n37975, n37976, n37977,
         n37978, n37979, n37980, n37981, n37982, n37983, n37984, n37985,
         n37986, n37987, n37988, n37989, n37990, n37991, n37992, n37993,
         n37994, n37995, n37996, n37997, n37998, n37999, n38000, n38001,
         n38002, n38003, n38004, n38005, n38006, n38007, n38008, n38009,
         n38010, n38011, n38012, n38013, n38014, n38015, n38016, n38017,
         n38018, n38019, n38020, n38021, n38022, n38023, n38024, n38025,
         n38026, n38027, n38028, n38029, n38030, n38031, n38032, n38033,
         n38034, n38035, n38036, n38037, n38038, n38039, n38040, n38041,
         n38042, n38043, n38044, n38045, n38046, n38047, n38048, n38049,
         n38050, n38051, n38052, n38053, n38054, n38055, n38056, n38057,
         n38058, n38059, n38060, n38061, n38062, n38063, n38064, n38065,
         n38066, n38067, n38068, n38069, n38070, n38071, n38072, n38073,
         n38074, n38075, n38076, n38077, n38078, n38079, n38080, n38081,
         n38082, n38083, n38084, n38085, n38086, n38087, n38088, n38089,
         n38090, n38091, n38092, n38093, n38094, n38095, n38096, n38097,
         n38098, n38099, n38100, n38101, n38102, n38103, n38104, n38105,
         n38106, n38107, n38108, n38109, n38110, n38111, n38112, n38113,
         n38114, n38115, n38116, n38117, n38118, n38119, n38120, n38121,
         n38122, n38123, n38124, n38125, n38126, n38127, n38128, n38129,
         n38130, n38131, n38132, n38133, n38134, n38135, n38136, n38137,
         n38138, n38139, n38140, n38141, n38142, n38143, n38144, n38145,
         n38146, n38147, n38148, n38149, n38150, n38151, n38152, n38153,
         n38154, n38155, n38156, n38157, n38158, n38159, n38160, n38161,
         n38162, n38163, n38164, n38165, n38166, n38167, n38168, n38169,
         n38170, n38171, n38172, n38173, n38174, n38175, n38176, n38177,
         n38178, n38179, n38180, n38181, n38182, n38183, n38184, n38185,
         n38186, n38187, n38188, n38189, n38190, n38191, n38192, n38193,
         n38194, n38195, n38196, n38197, n38198, n38199, n38200, n38201,
         n38202, n38203, n38204, n38205, n38206, n38207, n38208, n38209,
         n38210, n38211, n38212, n38213, n38214, n38215, n38216, n38217,
         n38218, n38219, n38220, n38221, n38222, n38223, n38224, n38225,
         n38226, n38227, n38228, n38229, n38230, n38231, n38232, n38233,
         n38234, n38235, n38236, n38237, n38238, n38239, n38240, n38241,
         n38242, n38243, n38244, n38245, n38246, n38247, n38248, n38249,
         n38250, n38251, n38252, n38253, n38254, n38255, n38256, n38257,
         n38258, n38259, n38260, n38261, n38262, n38263, n38264, n38265,
         n38266, n38267, n38268, n38269, n38270, n38271, n38272, n38273,
         n38274, n38275, n38276, n38277, n38278, n38279, n38280, n38281,
         n38282, n38283, n38284, n38285, n38286, n38287, n38288, n38289,
         n38290, n38291, n38292, n38293, n38294, n38295, n38296, n38297,
         n38298, n38299, n38300, n38301, n38302, n38303, n38304, n38305,
         n38306, n38307, n38308, n38309, n38310, n38311, n38312, n38313,
         n38314, n38315, n38316, n38317, n38318, n38319, n38320, n38321,
         n38322, n38323, n38324, n38325, n38326, n38327, n38328, n38329,
         n38330, n38331, n38332, n38333, n38334, n38335, n38336, n38337,
         n38338, n38339, n38340, n38341, n38342, n38343, n38344, n38345,
         n38346, n38347, n38348, n38349, n38350, n38351, n38352, n38353,
         n38354, n38355, n38356, n38357, n38358, n38359, n38360, n38361,
         n38362, n38363, n38364, n38365, n38366, n38367, n38368, n38369,
         n38370, n38371, n38372, n38373, n38374, n38375, n38376, n38377,
         n38378, n38379, n38380, n38381, n38382, n38383, n38384, n38385,
         n38386, n38387, n38388, n38389, n38390, n38391, n38392, n38393,
         n38394, n38395, n38396, n38397, n38398, n38399, n38400, n38401,
         n38402, n38403, n38404, n38405, n38406, n38407, n38408, n38409,
         n38410, n38411, n38412, n38413, n38414, n38415, n38416, n38417,
         n38418, n38419, n38420, n38421, n38422, n38423, n38424, n38425,
         n38426, n38427, n38428, n38429, n38430, n38431, n38432, n38433,
         n38434, n38435, n38436, n38437, n38438, n38439, n38440, n38441,
         n38442, n38443, n38444, n38445, n38446, n38447, n38448, n38449,
         n38450, n38451, n38452, n38453, n38454, n38455, n38456, n38457,
         n38458, n38459, n38460, n38461, n38462, n38463, n38464, n38465,
         n38466, n38467, n38468, n38469, n38470, n38471, n38472, n38473,
         n38474, n38475, n38476, n38477, n38478, n38479, n38480, n38481,
         n38482, n38483, n38484, n38485, n38486, n38487, n38488, n38489,
         n38490, n38491, n38492, n38493, n38494, n38495, n38496, n38497,
         n38498, n38499, n38500, n38501, n38502, n38503, n38504, n38505,
         n38506, n38507, n38508, n38509, n38510, n38511, n38512, n38513,
         n38514, n38515, n38516, n38517, n38518, n38519, n38520, n38521,
         n38522, n38523, n38524, n38525, n38526, n38527, n38528, n38529,
         n38530;
  wire   [511:0] sreg;

  DFF \sreg_reg[479]  ( .D(c[511]), .CLK(clk), .RST(rst), .Q(sreg[479]) );
  DFF \sreg_reg[478]  ( .D(c[510]), .CLK(clk), .RST(rst), .Q(sreg[478]) );
  DFF \sreg_reg[477]  ( .D(c[509]), .CLK(clk), .RST(rst), .Q(sreg[477]) );
  DFF \sreg_reg[476]  ( .D(c[508]), .CLK(clk), .RST(rst), .Q(sreg[476]) );
  DFF \sreg_reg[475]  ( .D(c[507]), .CLK(clk), .RST(rst), .Q(sreg[475]) );
  DFF \sreg_reg[474]  ( .D(c[506]), .CLK(clk), .RST(rst), .Q(sreg[474]) );
  DFF \sreg_reg[473]  ( .D(c[505]), .CLK(clk), .RST(rst), .Q(sreg[473]) );
  DFF \sreg_reg[472]  ( .D(c[504]), .CLK(clk), .RST(rst), .Q(sreg[472]) );
  DFF \sreg_reg[471]  ( .D(c[503]), .CLK(clk), .RST(rst), .Q(sreg[471]) );
  DFF \sreg_reg[470]  ( .D(c[502]), .CLK(clk), .RST(rst), .Q(sreg[470]) );
  DFF \sreg_reg[469]  ( .D(c[501]), .CLK(clk), .RST(rst), .Q(sreg[469]) );
  DFF \sreg_reg[468]  ( .D(c[500]), .CLK(clk), .RST(rst), .Q(sreg[468]) );
  DFF \sreg_reg[467]  ( .D(c[499]), .CLK(clk), .RST(rst), .Q(sreg[467]) );
  DFF \sreg_reg[466]  ( .D(c[498]), .CLK(clk), .RST(rst), .Q(sreg[466]) );
  DFF \sreg_reg[465]  ( .D(c[497]), .CLK(clk), .RST(rst), .Q(sreg[465]) );
  DFF \sreg_reg[464]  ( .D(c[496]), .CLK(clk), .RST(rst), .Q(sreg[464]) );
  DFF \sreg_reg[463]  ( .D(c[495]), .CLK(clk), .RST(rst), .Q(sreg[463]) );
  DFF \sreg_reg[462]  ( .D(c[494]), .CLK(clk), .RST(rst), .Q(sreg[462]) );
  DFF \sreg_reg[461]  ( .D(c[493]), .CLK(clk), .RST(rst), .Q(sreg[461]) );
  DFF \sreg_reg[460]  ( .D(c[492]), .CLK(clk), .RST(rst), .Q(sreg[460]) );
  DFF \sreg_reg[459]  ( .D(c[491]), .CLK(clk), .RST(rst), .Q(sreg[459]) );
  DFF \sreg_reg[458]  ( .D(c[490]), .CLK(clk), .RST(rst), .Q(sreg[458]) );
  DFF \sreg_reg[457]  ( .D(c[489]), .CLK(clk), .RST(rst), .Q(sreg[457]) );
  DFF \sreg_reg[456]  ( .D(c[488]), .CLK(clk), .RST(rst), .Q(sreg[456]) );
  DFF \sreg_reg[455]  ( .D(c[487]), .CLK(clk), .RST(rst), .Q(sreg[455]) );
  DFF \sreg_reg[454]  ( .D(c[486]), .CLK(clk), .RST(rst), .Q(sreg[454]) );
  DFF \sreg_reg[453]  ( .D(c[485]), .CLK(clk), .RST(rst), .Q(sreg[453]) );
  DFF \sreg_reg[452]  ( .D(c[484]), .CLK(clk), .RST(rst), .Q(sreg[452]) );
  DFF \sreg_reg[451]  ( .D(c[483]), .CLK(clk), .RST(rst), .Q(sreg[451]) );
  DFF \sreg_reg[450]  ( .D(c[482]), .CLK(clk), .RST(rst), .Q(sreg[450]) );
  DFF \sreg_reg[449]  ( .D(c[481]), .CLK(clk), .RST(rst), .Q(sreg[449]) );
  DFF \sreg_reg[448]  ( .D(c[480]), .CLK(clk), .RST(rst), .Q(sreg[448]) );
  DFF \sreg_reg[447]  ( .D(c[479]), .CLK(clk), .RST(rst), .Q(sreg[447]) );
  DFF \sreg_reg[446]  ( .D(c[478]), .CLK(clk), .RST(rst), .Q(sreg[446]) );
  DFF \sreg_reg[445]  ( .D(c[477]), .CLK(clk), .RST(rst), .Q(sreg[445]) );
  DFF \sreg_reg[444]  ( .D(c[476]), .CLK(clk), .RST(rst), .Q(sreg[444]) );
  DFF \sreg_reg[443]  ( .D(c[475]), .CLK(clk), .RST(rst), .Q(sreg[443]) );
  DFF \sreg_reg[442]  ( .D(c[474]), .CLK(clk), .RST(rst), .Q(sreg[442]) );
  DFF \sreg_reg[441]  ( .D(c[473]), .CLK(clk), .RST(rst), .Q(sreg[441]) );
  DFF \sreg_reg[440]  ( .D(c[472]), .CLK(clk), .RST(rst), .Q(sreg[440]) );
  DFF \sreg_reg[439]  ( .D(c[471]), .CLK(clk), .RST(rst), .Q(sreg[439]) );
  DFF \sreg_reg[438]  ( .D(c[470]), .CLK(clk), .RST(rst), .Q(sreg[438]) );
  DFF \sreg_reg[437]  ( .D(c[469]), .CLK(clk), .RST(rst), .Q(sreg[437]) );
  DFF \sreg_reg[436]  ( .D(c[468]), .CLK(clk), .RST(rst), .Q(sreg[436]) );
  DFF \sreg_reg[435]  ( .D(c[467]), .CLK(clk), .RST(rst), .Q(sreg[435]) );
  DFF \sreg_reg[434]  ( .D(c[466]), .CLK(clk), .RST(rst), .Q(sreg[434]) );
  DFF \sreg_reg[433]  ( .D(c[465]), .CLK(clk), .RST(rst), .Q(sreg[433]) );
  DFF \sreg_reg[432]  ( .D(c[464]), .CLK(clk), .RST(rst), .Q(sreg[432]) );
  DFF \sreg_reg[431]  ( .D(c[463]), .CLK(clk), .RST(rst), .Q(sreg[431]) );
  DFF \sreg_reg[430]  ( .D(c[462]), .CLK(clk), .RST(rst), .Q(sreg[430]) );
  DFF \sreg_reg[429]  ( .D(c[461]), .CLK(clk), .RST(rst), .Q(sreg[429]) );
  DFF \sreg_reg[428]  ( .D(c[460]), .CLK(clk), .RST(rst), .Q(sreg[428]) );
  DFF \sreg_reg[427]  ( .D(c[459]), .CLK(clk), .RST(rst), .Q(sreg[427]) );
  DFF \sreg_reg[426]  ( .D(c[458]), .CLK(clk), .RST(rst), .Q(sreg[426]) );
  DFF \sreg_reg[425]  ( .D(c[457]), .CLK(clk), .RST(rst), .Q(sreg[425]) );
  DFF \sreg_reg[424]  ( .D(c[456]), .CLK(clk), .RST(rst), .Q(sreg[424]) );
  DFF \sreg_reg[423]  ( .D(c[455]), .CLK(clk), .RST(rst), .Q(sreg[423]) );
  DFF \sreg_reg[422]  ( .D(c[454]), .CLK(clk), .RST(rst), .Q(sreg[422]) );
  DFF \sreg_reg[421]  ( .D(c[453]), .CLK(clk), .RST(rst), .Q(sreg[421]) );
  DFF \sreg_reg[420]  ( .D(c[452]), .CLK(clk), .RST(rst), .Q(sreg[420]) );
  DFF \sreg_reg[419]  ( .D(c[451]), .CLK(clk), .RST(rst), .Q(sreg[419]) );
  DFF \sreg_reg[418]  ( .D(c[450]), .CLK(clk), .RST(rst), .Q(sreg[418]) );
  DFF \sreg_reg[417]  ( .D(c[449]), .CLK(clk), .RST(rst), .Q(sreg[417]) );
  DFF \sreg_reg[416]  ( .D(c[448]), .CLK(clk), .RST(rst), .Q(sreg[416]) );
  DFF \sreg_reg[415]  ( .D(c[447]), .CLK(clk), .RST(rst), .Q(sreg[415]) );
  DFF \sreg_reg[414]  ( .D(c[446]), .CLK(clk), .RST(rst), .Q(sreg[414]) );
  DFF \sreg_reg[413]  ( .D(c[445]), .CLK(clk), .RST(rst), .Q(sreg[413]) );
  DFF \sreg_reg[412]  ( .D(c[444]), .CLK(clk), .RST(rst), .Q(sreg[412]) );
  DFF \sreg_reg[411]  ( .D(c[443]), .CLK(clk), .RST(rst), .Q(sreg[411]) );
  DFF \sreg_reg[410]  ( .D(c[442]), .CLK(clk), .RST(rst), .Q(sreg[410]) );
  DFF \sreg_reg[409]  ( .D(c[441]), .CLK(clk), .RST(rst), .Q(sreg[409]) );
  DFF \sreg_reg[408]  ( .D(c[440]), .CLK(clk), .RST(rst), .Q(sreg[408]) );
  DFF \sreg_reg[407]  ( .D(c[439]), .CLK(clk), .RST(rst), .Q(sreg[407]) );
  DFF \sreg_reg[406]  ( .D(c[438]), .CLK(clk), .RST(rst), .Q(sreg[406]) );
  DFF \sreg_reg[405]  ( .D(c[437]), .CLK(clk), .RST(rst), .Q(sreg[405]) );
  DFF \sreg_reg[404]  ( .D(c[436]), .CLK(clk), .RST(rst), .Q(sreg[404]) );
  DFF \sreg_reg[403]  ( .D(c[435]), .CLK(clk), .RST(rst), .Q(sreg[403]) );
  DFF \sreg_reg[402]  ( .D(c[434]), .CLK(clk), .RST(rst), .Q(sreg[402]) );
  DFF \sreg_reg[401]  ( .D(c[433]), .CLK(clk), .RST(rst), .Q(sreg[401]) );
  DFF \sreg_reg[400]  ( .D(c[432]), .CLK(clk), .RST(rst), .Q(sreg[400]) );
  DFF \sreg_reg[399]  ( .D(c[431]), .CLK(clk), .RST(rst), .Q(sreg[399]) );
  DFF \sreg_reg[398]  ( .D(c[430]), .CLK(clk), .RST(rst), .Q(sreg[398]) );
  DFF \sreg_reg[397]  ( .D(c[429]), .CLK(clk), .RST(rst), .Q(sreg[397]) );
  DFF \sreg_reg[396]  ( .D(c[428]), .CLK(clk), .RST(rst), .Q(sreg[396]) );
  DFF \sreg_reg[395]  ( .D(c[427]), .CLK(clk), .RST(rst), .Q(sreg[395]) );
  DFF \sreg_reg[394]  ( .D(c[426]), .CLK(clk), .RST(rst), .Q(sreg[394]) );
  DFF \sreg_reg[393]  ( .D(c[425]), .CLK(clk), .RST(rst), .Q(sreg[393]) );
  DFF \sreg_reg[392]  ( .D(c[424]), .CLK(clk), .RST(rst), .Q(sreg[392]) );
  DFF \sreg_reg[391]  ( .D(c[423]), .CLK(clk), .RST(rst), .Q(sreg[391]) );
  DFF \sreg_reg[390]  ( .D(c[422]), .CLK(clk), .RST(rst), .Q(sreg[390]) );
  DFF \sreg_reg[389]  ( .D(c[421]), .CLK(clk), .RST(rst), .Q(sreg[389]) );
  DFF \sreg_reg[388]  ( .D(c[420]), .CLK(clk), .RST(rst), .Q(sreg[388]) );
  DFF \sreg_reg[387]  ( .D(c[419]), .CLK(clk), .RST(rst), .Q(sreg[387]) );
  DFF \sreg_reg[386]  ( .D(c[418]), .CLK(clk), .RST(rst), .Q(sreg[386]) );
  DFF \sreg_reg[385]  ( .D(c[417]), .CLK(clk), .RST(rst), .Q(sreg[385]) );
  DFF \sreg_reg[384]  ( .D(c[416]), .CLK(clk), .RST(rst), .Q(sreg[384]) );
  DFF \sreg_reg[383]  ( .D(c[415]), .CLK(clk), .RST(rst), .Q(sreg[383]) );
  DFF \sreg_reg[382]  ( .D(c[414]), .CLK(clk), .RST(rst), .Q(sreg[382]) );
  DFF \sreg_reg[381]  ( .D(c[413]), .CLK(clk), .RST(rst), .Q(sreg[381]) );
  DFF \sreg_reg[380]  ( .D(c[412]), .CLK(clk), .RST(rst), .Q(sreg[380]) );
  DFF \sreg_reg[379]  ( .D(c[411]), .CLK(clk), .RST(rst), .Q(sreg[379]) );
  DFF \sreg_reg[378]  ( .D(c[410]), .CLK(clk), .RST(rst), .Q(sreg[378]) );
  DFF \sreg_reg[377]  ( .D(c[409]), .CLK(clk), .RST(rst), .Q(sreg[377]) );
  DFF \sreg_reg[376]  ( .D(c[408]), .CLK(clk), .RST(rst), .Q(sreg[376]) );
  DFF \sreg_reg[375]  ( .D(c[407]), .CLK(clk), .RST(rst), .Q(sreg[375]) );
  DFF \sreg_reg[374]  ( .D(c[406]), .CLK(clk), .RST(rst), .Q(sreg[374]) );
  DFF \sreg_reg[373]  ( .D(c[405]), .CLK(clk), .RST(rst), .Q(sreg[373]) );
  DFF \sreg_reg[372]  ( .D(c[404]), .CLK(clk), .RST(rst), .Q(sreg[372]) );
  DFF \sreg_reg[371]  ( .D(c[403]), .CLK(clk), .RST(rst), .Q(sreg[371]) );
  DFF \sreg_reg[370]  ( .D(c[402]), .CLK(clk), .RST(rst), .Q(sreg[370]) );
  DFF \sreg_reg[369]  ( .D(c[401]), .CLK(clk), .RST(rst), .Q(sreg[369]) );
  DFF \sreg_reg[368]  ( .D(c[400]), .CLK(clk), .RST(rst), .Q(sreg[368]) );
  DFF \sreg_reg[367]  ( .D(c[399]), .CLK(clk), .RST(rst), .Q(sreg[367]) );
  DFF \sreg_reg[366]  ( .D(c[398]), .CLK(clk), .RST(rst), .Q(sreg[366]) );
  DFF \sreg_reg[365]  ( .D(c[397]), .CLK(clk), .RST(rst), .Q(sreg[365]) );
  DFF \sreg_reg[364]  ( .D(c[396]), .CLK(clk), .RST(rst), .Q(sreg[364]) );
  DFF \sreg_reg[363]  ( .D(c[395]), .CLK(clk), .RST(rst), .Q(sreg[363]) );
  DFF \sreg_reg[362]  ( .D(c[394]), .CLK(clk), .RST(rst), .Q(sreg[362]) );
  DFF \sreg_reg[361]  ( .D(c[393]), .CLK(clk), .RST(rst), .Q(sreg[361]) );
  DFF \sreg_reg[360]  ( .D(c[392]), .CLK(clk), .RST(rst), .Q(sreg[360]) );
  DFF \sreg_reg[359]  ( .D(c[391]), .CLK(clk), .RST(rst), .Q(sreg[359]) );
  DFF \sreg_reg[358]  ( .D(c[390]), .CLK(clk), .RST(rst), .Q(sreg[358]) );
  DFF \sreg_reg[357]  ( .D(c[389]), .CLK(clk), .RST(rst), .Q(sreg[357]) );
  DFF \sreg_reg[356]  ( .D(c[388]), .CLK(clk), .RST(rst), .Q(sreg[356]) );
  DFF \sreg_reg[355]  ( .D(c[387]), .CLK(clk), .RST(rst), .Q(sreg[355]) );
  DFF \sreg_reg[354]  ( .D(c[386]), .CLK(clk), .RST(rst), .Q(sreg[354]) );
  DFF \sreg_reg[353]  ( .D(c[385]), .CLK(clk), .RST(rst), .Q(sreg[353]) );
  DFF \sreg_reg[352]  ( .D(c[384]), .CLK(clk), .RST(rst), .Q(sreg[352]) );
  DFF \sreg_reg[351]  ( .D(c[383]), .CLK(clk), .RST(rst), .Q(sreg[351]) );
  DFF \sreg_reg[350]  ( .D(c[382]), .CLK(clk), .RST(rst), .Q(sreg[350]) );
  DFF \sreg_reg[349]  ( .D(c[381]), .CLK(clk), .RST(rst), .Q(sreg[349]) );
  DFF \sreg_reg[348]  ( .D(c[380]), .CLK(clk), .RST(rst), .Q(sreg[348]) );
  DFF \sreg_reg[347]  ( .D(c[379]), .CLK(clk), .RST(rst), .Q(sreg[347]) );
  DFF \sreg_reg[346]  ( .D(c[378]), .CLK(clk), .RST(rst), .Q(sreg[346]) );
  DFF \sreg_reg[345]  ( .D(c[377]), .CLK(clk), .RST(rst), .Q(sreg[345]) );
  DFF \sreg_reg[344]  ( .D(c[376]), .CLK(clk), .RST(rst), .Q(sreg[344]) );
  DFF \sreg_reg[343]  ( .D(c[375]), .CLK(clk), .RST(rst), .Q(sreg[343]) );
  DFF \sreg_reg[342]  ( .D(c[374]), .CLK(clk), .RST(rst), .Q(sreg[342]) );
  DFF \sreg_reg[341]  ( .D(c[373]), .CLK(clk), .RST(rst), .Q(sreg[341]) );
  DFF \sreg_reg[340]  ( .D(c[372]), .CLK(clk), .RST(rst), .Q(sreg[340]) );
  DFF \sreg_reg[339]  ( .D(c[371]), .CLK(clk), .RST(rst), .Q(sreg[339]) );
  DFF \sreg_reg[338]  ( .D(c[370]), .CLK(clk), .RST(rst), .Q(sreg[338]) );
  DFF \sreg_reg[337]  ( .D(c[369]), .CLK(clk), .RST(rst), .Q(sreg[337]) );
  DFF \sreg_reg[336]  ( .D(c[368]), .CLK(clk), .RST(rst), .Q(sreg[336]) );
  DFF \sreg_reg[335]  ( .D(c[367]), .CLK(clk), .RST(rst), .Q(sreg[335]) );
  DFF \sreg_reg[334]  ( .D(c[366]), .CLK(clk), .RST(rst), .Q(sreg[334]) );
  DFF \sreg_reg[333]  ( .D(c[365]), .CLK(clk), .RST(rst), .Q(sreg[333]) );
  DFF \sreg_reg[332]  ( .D(c[364]), .CLK(clk), .RST(rst), .Q(sreg[332]) );
  DFF \sreg_reg[331]  ( .D(c[363]), .CLK(clk), .RST(rst), .Q(sreg[331]) );
  DFF \sreg_reg[330]  ( .D(c[362]), .CLK(clk), .RST(rst), .Q(sreg[330]) );
  DFF \sreg_reg[329]  ( .D(c[361]), .CLK(clk), .RST(rst), .Q(sreg[329]) );
  DFF \sreg_reg[328]  ( .D(c[360]), .CLK(clk), .RST(rst), .Q(sreg[328]) );
  DFF \sreg_reg[327]  ( .D(c[359]), .CLK(clk), .RST(rst), .Q(sreg[327]) );
  DFF \sreg_reg[326]  ( .D(c[358]), .CLK(clk), .RST(rst), .Q(sreg[326]) );
  DFF \sreg_reg[325]  ( .D(c[357]), .CLK(clk), .RST(rst), .Q(sreg[325]) );
  DFF \sreg_reg[324]  ( .D(c[356]), .CLK(clk), .RST(rst), .Q(sreg[324]) );
  DFF \sreg_reg[323]  ( .D(c[355]), .CLK(clk), .RST(rst), .Q(sreg[323]) );
  DFF \sreg_reg[322]  ( .D(c[354]), .CLK(clk), .RST(rst), .Q(sreg[322]) );
  DFF \sreg_reg[321]  ( .D(c[353]), .CLK(clk), .RST(rst), .Q(sreg[321]) );
  DFF \sreg_reg[320]  ( .D(c[352]), .CLK(clk), .RST(rst), .Q(sreg[320]) );
  DFF \sreg_reg[319]  ( .D(c[351]), .CLK(clk), .RST(rst), .Q(sreg[319]) );
  DFF \sreg_reg[318]  ( .D(c[350]), .CLK(clk), .RST(rst), .Q(sreg[318]) );
  DFF \sreg_reg[317]  ( .D(c[349]), .CLK(clk), .RST(rst), .Q(sreg[317]) );
  DFF \sreg_reg[316]  ( .D(c[348]), .CLK(clk), .RST(rst), .Q(sreg[316]) );
  DFF \sreg_reg[315]  ( .D(c[347]), .CLK(clk), .RST(rst), .Q(sreg[315]) );
  DFF \sreg_reg[314]  ( .D(c[346]), .CLK(clk), .RST(rst), .Q(sreg[314]) );
  DFF \sreg_reg[313]  ( .D(c[345]), .CLK(clk), .RST(rst), .Q(sreg[313]) );
  DFF \sreg_reg[312]  ( .D(c[344]), .CLK(clk), .RST(rst), .Q(sreg[312]) );
  DFF \sreg_reg[311]  ( .D(c[343]), .CLK(clk), .RST(rst), .Q(sreg[311]) );
  DFF \sreg_reg[310]  ( .D(c[342]), .CLK(clk), .RST(rst), .Q(sreg[310]) );
  DFF \sreg_reg[309]  ( .D(c[341]), .CLK(clk), .RST(rst), .Q(sreg[309]) );
  DFF \sreg_reg[308]  ( .D(c[340]), .CLK(clk), .RST(rst), .Q(sreg[308]) );
  DFF \sreg_reg[307]  ( .D(c[339]), .CLK(clk), .RST(rst), .Q(sreg[307]) );
  DFF \sreg_reg[306]  ( .D(c[338]), .CLK(clk), .RST(rst), .Q(sreg[306]) );
  DFF \sreg_reg[305]  ( .D(c[337]), .CLK(clk), .RST(rst), .Q(sreg[305]) );
  DFF \sreg_reg[304]  ( .D(c[336]), .CLK(clk), .RST(rst), .Q(sreg[304]) );
  DFF \sreg_reg[303]  ( .D(c[335]), .CLK(clk), .RST(rst), .Q(sreg[303]) );
  DFF \sreg_reg[302]  ( .D(c[334]), .CLK(clk), .RST(rst), .Q(sreg[302]) );
  DFF \sreg_reg[301]  ( .D(c[333]), .CLK(clk), .RST(rst), .Q(sreg[301]) );
  DFF \sreg_reg[300]  ( .D(c[332]), .CLK(clk), .RST(rst), .Q(sreg[300]) );
  DFF \sreg_reg[299]  ( .D(c[331]), .CLK(clk), .RST(rst), .Q(sreg[299]) );
  DFF \sreg_reg[298]  ( .D(c[330]), .CLK(clk), .RST(rst), .Q(sreg[298]) );
  DFF \sreg_reg[297]  ( .D(c[329]), .CLK(clk), .RST(rst), .Q(sreg[297]) );
  DFF \sreg_reg[296]  ( .D(c[328]), .CLK(clk), .RST(rst), .Q(sreg[296]) );
  DFF \sreg_reg[295]  ( .D(c[327]), .CLK(clk), .RST(rst), .Q(sreg[295]) );
  DFF \sreg_reg[294]  ( .D(c[326]), .CLK(clk), .RST(rst), .Q(sreg[294]) );
  DFF \sreg_reg[293]  ( .D(c[325]), .CLK(clk), .RST(rst), .Q(sreg[293]) );
  DFF \sreg_reg[292]  ( .D(c[324]), .CLK(clk), .RST(rst), .Q(sreg[292]) );
  DFF \sreg_reg[291]  ( .D(c[323]), .CLK(clk), .RST(rst), .Q(sreg[291]) );
  DFF \sreg_reg[290]  ( .D(c[322]), .CLK(clk), .RST(rst), .Q(sreg[290]) );
  DFF \sreg_reg[289]  ( .D(c[321]), .CLK(clk), .RST(rst), .Q(sreg[289]) );
  DFF \sreg_reg[288]  ( .D(c[320]), .CLK(clk), .RST(rst), .Q(sreg[288]) );
  DFF \sreg_reg[287]  ( .D(c[319]), .CLK(clk), .RST(rst), .Q(sreg[287]) );
  DFF \sreg_reg[286]  ( .D(c[318]), .CLK(clk), .RST(rst), .Q(sreg[286]) );
  DFF \sreg_reg[285]  ( .D(c[317]), .CLK(clk), .RST(rst), .Q(sreg[285]) );
  DFF \sreg_reg[284]  ( .D(c[316]), .CLK(clk), .RST(rst), .Q(sreg[284]) );
  DFF \sreg_reg[283]  ( .D(c[315]), .CLK(clk), .RST(rst), .Q(sreg[283]) );
  DFF \sreg_reg[282]  ( .D(c[314]), .CLK(clk), .RST(rst), .Q(sreg[282]) );
  DFF \sreg_reg[281]  ( .D(c[313]), .CLK(clk), .RST(rst), .Q(sreg[281]) );
  DFF \sreg_reg[280]  ( .D(c[312]), .CLK(clk), .RST(rst), .Q(sreg[280]) );
  DFF \sreg_reg[279]  ( .D(c[311]), .CLK(clk), .RST(rst), .Q(sreg[279]) );
  DFF \sreg_reg[278]  ( .D(c[310]), .CLK(clk), .RST(rst), .Q(sreg[278]) );
  DFF \sreg_reg[277]  ( .D(c[309]), .CLK(clk), .RST(rst), .Q(sreg[277]) );
  DFF \sreg_reg[276]  ( .D(c[308]), .CLK(clk), .RST(rst), .Q(sreg[276]) );
  DFF \sreg_reg[275]  ( .D(c[307]), .CLK(clk), .RST(rst), .Q(sreg[275]) );
  DFF \sreg_reg[274]  ( .D(c[306]), .CLK(clk), .RST(rst), .Q(sreg[274]) );
  DFF \sreg_reg[273]  ( .D(c[305]), .CLK(clk), .RST(rst), .Q(sreg[273]) );
  DFF \sreg_reg[272]  ( .D(c[304]), .CLK(clk), .RST(rst), .Q(sreg[272]) );
  DFF \sreg_reg[271]  ( .D(c[303]), .CLK(clk), .RST(rst), .Q(sreg[271]) );
  DFF \sreg_reg[270]  ( .D(c[302]), .CLK(clk), .RST(rst), .Q(sreg[270]) );
  DFF \sreg_reg[269]  ( .D(c[301]), .CLK(clk), .RST(rst), .Q(sreg[269]) );
  DFF \sreg_reg[268]  ( .D(c[300]), .CLK(clk), .RST(rst), .Q(sreg[268]) );
  DFF \sreg_reg[267]  ( .D(c[299]), .CLK(clk), .RST(rst), .Q(sreg[267]) );
  DFF \sreg_reg[266]  ( .D(c[298]), .CLK(clk), .RST(rst), .Q(sreg[266]) );
  DFF \sreg_reg[265]  ( .D(c[297]), .CLK(clk), .RST(rst), .Q(sreg[265]) );
  DFF \sreg_reg[264]  ( .D(c[296]), .CLK(clk), .RST(rst), .Q(sreg[264]) );
  DFF \sreg_reg[263]  ( .D(c[295]), .CLK(clk), .RST(rst), .Q(sreg[263]) );
  DFF \sreg_reg[262]  ( .D(c[294]), .CLK(clk), .RST(rst), .Q(sreg[262]) );
  DFF \sreg_reg[261]  ( .D(c[293]), .CLK(clk), .RST(rst), .Q(sreg[261]) );
  DFF \sreg_reg[260]  ( .D(c[292]), .CLK(clk), .RST(rst), .Q(sreg[260]) );
  DFF \sreg_reg[259]  ( .D(c[291]), .CLK(clk), .RST(rst), .Q(sreg[259]) );
  DFF \sreg_reg[258]  ( .D(c[290]), .CLK(clk), .RST(rst), .Q(sreg[258]) );
  DFF \sreg_reg[257]  ( .D(c[289]), .CLK(clk), .RST(rst), .Q(sreg[257]) );
  DFF \sreg_reg[256]  ( .D(c[288]), .CLK(clk), .RST(rst), .Q(sreg[256]) );
  DFF \sreg_reg[255]  ( .D(c[287]), .CLK(clk), .RST(rst), .Q(sreg[255]) );
  DFF \sreg_reg[254]  ( .D(c[286]), .CLK(clk), .RST(rst), .Q(sreg[254]) );
  DFF \sreg_reg[253]  ( .D(c[285]), .CLK(clk), .RST(rst), .Q(sreg[253]) );
  DFF \sreg_reg[252]  ( .D(c[284]), .CLK(clk), .RST(rst), .Q(sreg[252]) );
  DFF \sreg_reg[251]  ( .D(c[283]), .CLK(clk), .RST(rst), .Q(sreg[251]) );
  DFF \sreg_reg[250]  ( .D(c[282]), .CLK(clk), .RST(rst), .Q(sreg[250]) );
  DFF \sreg_reg[249]  ( .D(c[281]), .CLK(clk), .RST(rst), .Q(sreg[249]) );
  DFF \sreg_reg[248]  ( .D(c[280]), .CLK(clk), .RST(rst), .Q(sreg[248]) );
  DFF \sreg_reg[247]  ( .D(c[279]), .CLK(clk), .RST(rst), .Q(sreg[247]) );
  DFF \sreg_reg[246]  ( .D(c[278]), .CLK(clk), .RST(rst), .Q(sreg[246]) );
  DFF \sreg_reg[245]  ( .D(c[277]), .CLK(clk), .RST(rst), .Q(sreg[245]) );
  DFF \sreg_reg[244]  ( .D(c[276]), .CLK(clk), .RST(rst), .Q(sreg[244]) );
  DFF \sreg_reg[243]  ( .D(c[275]), .CLK(clk), .RST(rst), .Q(sreg[243]) );
  DFF \sreg_reg[242]  ( .D(c[274]), .CLK(clk), .RST(rst), .Q(sreg[242]) );
  DFF \sreg_reg[241]  ( .D(c[273]), .CLK(clk), .RST(rst), .Q(sreg[241]) );
  DFF \sreg_reg[240]  ( .D(c[272]), .CLK(clk), .RST(rst), .Q(sreg[240]) );
  DFF \sreg_reg[239]  ( .D(c[271]), .CLK(clk), .RST(rst), .Q(sreg[239]) );
  DFF \sreg_reg[238]  ( .D(c[270]), .CLK(clk), .RST(rst), .Q(sreg[238]) );
  DFF \sreg_reg[237]  ( .D(c[269]), .CLK(clk), .RST(rst), .Q(sreg[237]) );
  DFF \sreg_reg[236]  ( .D(c[268]), .CLK(clk), .RST(rst), .Q(sreg[236]) );
  DFF \sreg_reg[235]  ( .D(c[267]), .CLK(clk), .RST(rst), .Q(sreg[235]) );
  DFF \sreg_reg[234]  ( .D(c[266]), .CLK(clk), .RST(rst), .Q(sreg[234]) );
  DFF \sreg_reg[233]  ( .D(c[265]), .CLK(clk), .RST(rst), .Q(sreg[233]) );
  DFF \sreg_reg[232]  ( .D(c[264]), .CLK(clk), .RST(rst), .Q(sreg[232]) );
  DFF \sreg_reg[231]  ( .D(c[263]), .CLK(clk), .RST(rst), .Q(sreg[231]) );
  DFF \sreg_reg[230]  ( .D(c[262]), .CLK(clk), .RST(rst), .Q(sreg[230]) );
  DFF \sreg_reg[229]  ( .D(c[261]), .CLK(clk), .RST(rst), .Q(sreg[229]) );
  DFF \sreg_reg[228]  ( .D(c[260]), .CLK(clk), .RST(rst), .Q(sreg[228]) );
  DFF \sreg_reg[227]  ( .D(c[259]), .CLK(clk), .RST(rst), .Q(sreg[227]) );
  DFF \sreg_reg[226]  ( .D(c[258]), .CLK(clk), .RST(rst), .Q(sreg[226]) );
  DFF \sreg_reg[225]  ( .D(c[257]), .CLK(clk), .RST(rst), .Q(sreg[225]) );
  DFF \sreg_reg[224]  ( .D(c[256]), .CLK(clk), .RST(rst), .Q(sreg[224]) );
  DFF \sreg_reg[223]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(c[223]) );
  DFF \sreg_reg[222]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(c[222]) );
  DFF \sreg_reg[221]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(c[221]) );
  DFF \sreg_reg[220]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(c[220]) );
  DFF \sreg_reg[219]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(c[219]) );
  DFF \sreg_reg[218]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(c[218]) );
  DFF \sreg_reg[217]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(c[217]) );
  DFF \sreg_reg[216]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(c[216]) );
  DFF \sreg_reg[215]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(c[215]) );
  DFF \sreg_reg[214]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(c[214]) );
  DFF \sreg_reg[213]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(c[213]) );
  DFF \sreg_reg[212]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(c[212]) );
  DFF \sreg_reg[211]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(c[211]) );
  DFF \sreg_reg[210]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(c[210]) );
  DFF \sreg_reg[209]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(c[209]) );
  DFF \sreg_reg[208]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(c[208]) );
  DFF \sreg_reg[207]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(c[207]) );
  DFF \sreg_reg[206]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(c[206]) );
  DFF \sreg_reg[205]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(c[205]) );
  DFF \sreg_reg[204]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(c[204]) );
  DFF \sreg_reg[203]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(c[203]) );
  DFF \sreg_reg[202]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(c[202]) );
  DFF \sreg_reg[201]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(c[201]) );
  DFF \sreg_reg[200]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(c[200]) );
  DFF \sreg_reg[199]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(c[199]) );
  DFF \sreg_reg[198]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(c[198]) );
  DFF \sreg_reg[197]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(c[197]) );
  DFF \sreg_reg[196]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(c[196]) );
  DFF \sreg_reg[195]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(c[195]) );
  DFF \sreg_reg[194]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(c[194]) );
  DFF \sreg_reg[193]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(c[193]) );
  DFF \sreg_reg[192]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(c[192]) );
  DFF \sreg_reg[191]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(c[191]) );
  DFF \sreg_reg[190]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(c[190]) );
  DFF \sreg_reg[189]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(c[189]) );
  DFF \sreg_reg[188]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(c[188]) );
  DFF \sreg_reg[187]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(c[187]) );
  DFF \sreg_reg[186]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(c[186]) );
  DFF \sreg_reg[185]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(c[185]) );
  DFF \sreg_reg[184]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(c[184]) );
  DFF \sreg_reg[183]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(c[183]) );
  DFF \sreg_reg[182]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(c[182]) );
  DFF \sreg_reg[181]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(c[181]) );
  DFF \sreg_reg[180]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(c[180]) );
  DFF \sreg_reg[179]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(c[179]) );
  DFF \sreg_reg[178]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(c[178]) );
  DFF \sreg_reg[177]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(c[177]) );
  DFF \sreg_reg[176]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(c[176]) );
  DFF \sreg_reg[175]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(c[175]) );
  DFF \sreg_reg[174]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(c[174]) );
  DFF \sreg_reg[173]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(c[173]) );
  DFF \sreg_reg[172]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(c[172]) );
  DFF \sreg_reg[171]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(c[171]) );
  DFF \sreg_reg[170]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(c[170]) );
  DFF \sreg_reg[169]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(c[169]) );
  DFF \sreg_reg[168]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(c[168]) );
  DFF \sreg_reg[167]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(c[167]) );
  DFF \sreg_reg[166]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(c[166]) );
  DFF \sreg_reg[165]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(c[165]) );
  DFF \sreg_reg[164]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(c[164]) );
  DFF \sreg_reg[163]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(c[163]) );
  DFF \sreg_reg[162]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(c[162]) );
  DFF \sreg_reg[161]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(c[161]) );
  DFF \sreg_reg[160]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(c[160]) );
  DFF \sreg_reg[159]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(c[159]) );
  DFF \sreg_reg[158]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(c[158]) );
  DFF \sreg_reg[157]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(c[157]) );
  DFF \sreg_reg[156]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(c[156]) );
  DFF \sreg_reg[155]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(c[155]) );
  DFF \sreg_reg[154]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(c[154]) );
  DFF \sreg_reg[153]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(c[153]) );
  DFF \sreg_reg[152]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(c[152]) );
  DFF \sreg_reg[151]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(c[151]) );
  DFF \sreg_reg[150]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(c[150]) );
  DFF \sreg_reg[149]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(c[149]) );
  DFF \sreg_reg[148]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(c[148]) );
  DFF \sreg_reg[147]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(c[147]) );
  DFF \sreg_reg[146]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(c[146]) );
  DFF \sreg_reg[145]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(c[145]) );
  DFF \sreg_reg[144]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(c[144]) );
  DFF \sreg_reg[143]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(c[143]) );
  DFF \sreg_reg[142]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(c[142]) );
  DFF \sreg_reg[141]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(c[141]) );
  DFF \sreg_reg[140]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(c[140]) );
  DFF \sreg_reg[139]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(c[139]) );
  DFF \sreg_reg[138]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(c[138]) );
  DFF \sreg_reg[137]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(c[137]) );
  DFF \sreg_reg[136]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(c[136]) );
  DFF \sreg_reg[135]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(c[135]) );
  DFF \sreg_reg[134]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(c[134]) );
  DFF \sreg_reg[133]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(c[133]) );
  DFF \sreg_reg[132]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(c[132]) );
  DFF \sreg_reg[131]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(c[131]) );
  DFF \sreg_reg[130]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(c[130]) );
  DFF \sreg_reg[129]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(c[129]) );
  DFF \sreg_reg[128]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(c[128]) );
  DFF \sreg_reg[127]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(c[127]) );
  DFF \sreg_reg[126]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(c[126]) );
  DFF \sreg_reg[125]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(c[125]) );
  DFF \sreg_reg[124]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(c[124]) );
  DFF \sreg_reg[123]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(c[123]) );
  DFF \sreg_reg[122]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(c[122]) );
  DFF \sreg_reg[121]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(c[121]) );
  DFF \sreg_reg[120]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(c[120]) );
  DFF \sreg_reg[119]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[118]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[117]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[116]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[115]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[114]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[113]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[112]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[111]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[110]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[109]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[108]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[107]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[106]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[105]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[104]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[103]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[102]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[101]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[100]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[99]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[98]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[97]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[96]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[95]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[94]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[93]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[92]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[91]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[90]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[89]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[88]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[87]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[86]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[85]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[84]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[83]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[82]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[81]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[80]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[79]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[78]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[77]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[76]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[75]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[74]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[73]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[72]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[71]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[70]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[69]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[68]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[67]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[66]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[65]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[64]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[63]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[62]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[0]) );
  XOR U35 ( .A(n35961), .B(n35960), .Z(n35962) );
  XOR U36 ( .A(n35527), .B(n35526), .Z(n35528) );
  XOR U37 ( .A(n35535), .B(n35534), .Z(n35550) );
  XOR U38 ( .A(n37059), .B(n37058), .Z(n37045) );
  XOR U39 ( .A(n36986), .B(n36985), .Z(n36973) );
  XNOR U40 ( .A(n37492), .B(n37491), .Z(n37519) );
  XOR U41 ( .A(n37678), .B(n37677), .Z(n37695) );
  XOR U42 ( .A(n37913), .B(n37912), .Z(n37951) );
  XOR U43 ( .A(n37979), .B(n37978), .Z(n38005) );
  XOR U44 ( .A(n38000), .B(n37999), .Z(n38001) );
  XOR U45 ( .A(n37857), .B(n37856), .Z(n37874) );
  NANDN U46 ( .A(n38239), .B(n38238), .Z(n1) );
  NANDN U47 ( .A(n38295), .B(n38237), .Z(n2) );
  NAND U48 ( .A(n1), .B(n2), .Z(n38275) );
  NAND U49 ( .A(n38341), .B(n38340), .Z(n3) );
  NANDN U50 ( .A(n38376), .B(n38339), .Z(n4) );
  NAND U51 ( .A(n3), .B(n4), .Z(n38364) );
  XOR U52 ( .A(n35742), .B(n35741), .Z(n35743) );
  XOR U53 ( .A(n35963), .B(n35962), .Z(n35972) );
  XOR U54 ( .A(n36183), .B(n36182), .Z(n36184) );
  XOR U55 ( .A(n36701), .B(n36700), .Z(n36702) );
  XOR U56 ( .A(n36796), .B(n36795), .Z(n36797) );
  XOR U57 ( .A(n35396), .B(n35395), .Z(n35397) );
  XOR U58 ( .A(n35666), .B(n35665), .Z(n35705) );
  XOR U59 ( .A(n35893), .B(n35892), .Z(n35894) );
  XOR U60 ( .A(n35887), .B(n35886), .Z(n35888) );
  XOR U61 ( .A(n36478), .B(n36477), .Z(n36479) );
  XOR U62 ( .A(n36614), .B(n36613), .Z(n36615) );
  XOR U63 ( .A(n36721), .B(n36720), .Z(n36657) );
  XOR U64 ( .A(n36742), .B(n36741), .Z(n36651) );
  XOR U65 ( .A(n36823), .B(n36822), .Z(n36859) );
  XNOR U66 ( .A(n36792), .B(n36791), .Z(n36866) );
  XOR U67 ( .A(n37046), .B(n37045), .Z(n37047) );
  XOR U68 ( .A(n35756), .B(n35755), .Z(n35766) );
  XOR U69 ( .A(n36530), .B(n36529), .Z(n36539) );
  XOR U70 ( .A(n37190), .B(n37189), .Z(n37219) );
  XOR U71 ( .A(n37196), .B(n37195), .Z(n37135) );
  XOR U72 ( .A(n37290), .B(n37289), .Z(n37250) );
  XOR U73 ( .A(n37246), .B(n37245), .Z(n37308) );
  XOR U74 ( .A(n37409), .B(n37408), .Z(n37401) );
  XNOR U75 ( .A(n37498), .B(n37497), .Z(n37521) );
  NAND U76 ( .A(n37487), .B(n38064), .Z(n5) );
  NANDN U77 ( .A(n37488), .B(n37579), .Z(n6) );
  AND U78 ( .A(n5), .B(n6), .Z(n37546) );
  XOR U79 ( .A(n37567), .B(n37566), .Z(n37604) );
  XOR U80 ( .A(n37952), .B(n37951), .Z(n37953) );
  XOR U81 ( .A(n38056), .B(n38055), .Z(n38057) );
  XOR U82 ( .A(n35762), .B(n35761), .Z(n35645) );
  XOR U83 ( .A(n36197), .B(n36196), .Z(n36200) );
  XOR U84 ( .A(n36900), .B(n36899), .Z(n36995) );
  XOR U85 ( .A(n37016), .B(n37015), .Z(n37018) );
  XOR U86 ( .A(n37238), .B(n37237), .Z(n37239) );
  XOR U87 ( .A(n37728), .B(n37727), .Z(n37730) );
  XOR U88 ( .A(n37901), .B(n37900), .Z(n37894) );
  XOR U89 ( .A(n38002), .B(n38001), .Z(n38011) );
  NAND U90 ( .A(n37979), .B(n37978), .Z(n7) );
  NANDN U91 ( .A(n38044), .B(n37977), .Z(n8) );
  NAND U92 ( .A(n7), .B(n8), .Z(n38087) );
  XOR U93 ( .A(n38310), .B(n38309), .Z(n38274) );
  XOR U94 ( .A(n38336), .B(n38335), .Z(n38329) );
  XOR U95 ( .A(n38362), .B(n38361), .Z(n38363) );
  XOR U96 ( .A(n38423), .B(n38422), .Z(n38412) );
  XOR U97 ( .A(n37817), .B(n37816), .Z(n37808) );
  XNOR U98 ( .A(n38229), .B(n38230), .Z(n9) );
  XNOR U99 ( .A(n38228), .B(n9), .Z(n38222) );
  NAND U100 ( .A(n194), .B(n38419), .Z(n10) );
  NANDN U101 ( .A(n38457), .B(n38456), .Z(n11) );
  NAND U102 ( .A(n10), .B(n11), .Z(n38440) );
  XOR U103 ( .A(n38475), .B(n38474), .Z(n38478) );
  XOR U104 ( .A(n35748), .B(n35747), .Z(n35749) );
  XOR U105 ( .A(n36042), .B(n36041), .Z(n36043) );
  NANDN U106 ( .A(b[0]), .B(a[255]), .Z(n12) );
  AND U107 ( .A(b[1]), .B(n12), .Z(n35981) );
  XOR U108 ( .A(n36260), .B(n36259), .Z(n36261) );
  XOR U109 ( .A(n36466), .B(n36465), .Z(n36467) );
  XOR U110 ( .A(n35392), .B(n35391), .Z(n35426) );
  XOR U111 ( .A(n35533), .B(n35532), .Z(n35534) );
  XOR U112 ( .A(n35529), .B(n35528), .Z(n35538) );
  XOR U113 ( .A(n35589), .B(n35588), .Z(n35551) );
  XOR U114 ( .A(n35545), .B(n35544), .Z(n35547) );
  XNOR U115 ( .A(n35595), .B(n35594), .Z(n35497) );
  XOR U116 ( .A(n35664), .B(n35663), .Z(n35665) );
  XOR U117 ( .A(n35660), .B(n35659), .Z(n35669) );
  XNOR U118 ( .A(n35652), .B(n35651), .Z(n35654) );
  XOR U119 ( .A(n35889), .B(n35888), .Z(n35898) );
  XNOR U120 ( .A(n35895), .B(n35894), .Z(n35812) );
  XOR U121 ( .A(n35969), .B(n35968), .Z(n35999) );
  XNOR U122 ( .A(n35975), .B(n35974), .Z(n35956) );
  XOR U123 ( .A(n36094), .B(n36093), .Z(n36121) );
  XOR U124 ( .A(n36189), .B(n36188), .Z(n36190) );
  XNOR U125 ( .A(n36157), .B(n36156), .Z(n36159) );
  XNOR U126 ( .A(n36268), .B(n36267), .Z(n36278) );
  XNOR U127 ( .A(n36333), .B(n36332), .Z(n36238) );
  XOR U128 ( .A(n36486), .B(n36485), .Z(n36381) );
  XOR U129 ( .A(n36558), .B(n36557), .Z(n36559) );
  XNOR U130 ( .A(n36616), .B(n36615), .Z(n36522) );
  XOR U131 ( .A(n36516), .B(n36515), .Z(n36518) );
  XOR U132 ( .A(n36715), .B(n36714), .Z(n36653) );
  XOR U133 ( .A(n36860), .B(n36859), .Z(n36861) );
  XNOR U134 ( .A(n36850), .B(n36849), .Z(n36867) );
  XOR U135 ( .A(n36854), .B(n36853), .Z(n36856) );
  XOR U136 ( .A(n37063), .B(n37062), .Z(n37064) );
  XNOR U137 ( .A(n36968), .B(n36967), .Z(n36977) );
  XOR U138 ( .A(n36928), .B(n36927), .Z(n36983) );
  XOR U139 ( .A(n37358), .B(n37357), .Z(n37359) );
  XOR U140 ( .A(n37502), .B(n37501), .Z(n37503) );
  XOR U141 ( .A(n37599), .B(n37598), .Z(n37600) );
  XOR U142 ( .A(n37756), .B(n37755), .Z(n37757) );
  XOR U143 ( .A(n37843), .B(n37842), .Z(n37844) );
  XOR U144 ( .A(n37933), .B(n37932), .Z(n37935) );
  XOR U145 ( .A(n35601), .B(n35600), .Z(n35605) );
  XOR U146 ( .A(n36542), .B(n36541), .Z(n36509) );
  XOR U147 ( .A(n36660), .B(n36659), .Z(n36708) );
  XNOR U148 ( .A(n37106), .B(n37105), .Z(n37039) );
  XOR U149 ( .A(n37314), .B(n37313), .Z(n37315) );
  XNOR U150 ( .A(n37252), .B(n37251), .Z(n37307) );
  XNOR U151 ( .A(n37397), .B(n37396), .Z(n37400) );
  XNOR U152 ( .A(n37518), .B(n37517), .Z(n37463) );
  XNOR U153 ( .A(n37595), .B(n37594), .Z(n37545) );
  XOR U154 ( .A(n37696), .B(n37695), .Z(n37697) );
  XOR U155 ( .A(n37764), .B(n37763), .Z(n37788) );
  XNOR U156 ( .A(n37863), .B(n37862), .Z(n37849) );
  XOR U157 ( .A(n38058), .B(n38057), .Z(n38081) );
  XOR U158 ( .A(n38126), .B(n38125), .Z(n38127) );
  XOR U159 ( .A(n38191), .B(n38190), .Z(n38192) );
  XOR U160 ( .A(n38197), .B(n38196), .Z(n38199) );
  XOR U161 ( .A(n35646), .B(n35645), .Z(n35648) );
  XNOR U162 ( .A(n35907), .B(n35906), .Z(n35917) );
  XOR U163 ( .A(n35794), .B(n35793), .Z(n35796) );
  XOR U164 ( .A(n35945), .B(n35944), .Z(n36061) );
  XOR U165 ( .A(n35937), .B(n35936), .Z(n35938) );
  XOR U166 ( .A(n36201), .B(n36200), .Z(n36203) );
  XOR U167 ( .A(n36080), .B(n36079), .Z(n36082) );
  XOR U168 ( .A(n36369), .B(n36368), .Z(n36371) );
  XOR U169 ( .A(n36620), .B(n36619), .Z(n36621) );
  XOR U170 ( .A(n36772), .B(n36771), .Z(n36773) );
  XOR U171 ( .A(n36998), .B(n36997), .Z(n36894) );
  XNOR U172 ( .A(n37024), .B(n37023), .Z(n37017) );
  XOR U173 ( .A(n37130), .B(n37129), .Z(n37131) );
  XOR U174 ( .A(n37320), .B(n37319), .Z(n37321) );
  XOR U175 ( .A(n37526), .B(n37525), .Z(n37527) );
  XOR U176 ( .A(n37619), .B(n37618), .Z(n37541) );
  XOR U177 ( .A(n37643), .B(n37642), .Z(n37644) );
  XNOR U178 ( .A(n37797), .B(n37796), .Z(n37729) );
  XOR U179 ( .A(n38018), .B(n38017), .Z(n38019) );
  XOR U180 ( .A(n38088), .B(n38087), .Z(n38090) );
  XOR U181 ( .A(n38038), .B(n38037), .Z(n38039) );
  XOR U182 ( .A(n38328), .B(n38327), .Z(n38330) );
  XOR U183 ( .A(n38411), .B(n38410), .Z(n38413) );
  XOR U184 ( .A(n36345), .B(n36344), .Z(n36220) );
  XOR U185 ( .A(n36363), .B(n36362), .Z(n36364) );
  XOR U186 ( .A(n37809), .B(n37808), .Z(n37810) );
  XOR U187 ( .A(n37887), .B(n37886), .Z(n37888) );
  XOR U188 ( .A(n38170), .B(n38169), .Z(n38161) );
  XOR U189 ( .A(n38223), .B(n38222), .Z(n38224) );
  XNOR U190 ( .A(n38277), .B(n38276), .Z(n38269) );
  XOR U191 ( .A(n38364), .B(n38363), .Z(n38390) );
  XOR U192 ( .A(n38441), .B(n38440), .Z(n38443) );
  XOR U193 ( .A(n38497), .B(n38496), .Z(n38498) );
  XOR U194 ( .A(n35462), .B(n35461), .Z(n35463) );
  XOR U195 ( .A(n35468), .B(n35467), .Z(n35469) );
  XOR U196 ( .A(n35503), .B(n35502), .Z(n35504) );
  XOR U197 ( .A(n35694), .B(n35693), .Z(n35695) );
  XOR U198 ( .A(n35863), .B(n35862), .Z(n35864) );
  XOR U199 ( .A(n35851), .B(n35850), .Z(n35852) );
  XOR U200 ( .A(n35845), .B(n35844), .Z(n35846) );
  XOR U201 ( .A(n35967), .B(n35966), .Z(n35968) );
  XOR U202 ( .A(n36290), .B(n36289), .Z(n36291) );
  XOR U203 ( .A(n36393), .B(n36392), .Z(n36395) );
  XOR U204 ( .A(n36719), .B(n36718), .Z(n36720) );
  XOR U205 ( .A(n35390), .B(n35389), .Z(n35391) );
  XOR U206 ( .A(n35398), .B(n35397), .Z(n35403) );
  XOR U207 ( .A(n35539), .B(n35538), .Z(n35540) );
  XOR U208 ( .A(n35670), .B(n35669), .Z(n35671) );
  XOR U209 ( .A(n35750), .B(n35749), .Z(n35706) );
  XOR U210 ( .A(n35700), .B(n35699), .Z(n35702) );
  XOR U211 ( .A(n35806), .B(n35805), .Z(n35808) );
  XNOR U212 ( .A(n35901), .B(n35900), .Z(n35858) );
  XOR U213 ( .A(n36044), .B(n36043), .Z(n36000) );
  XNOR U214 ( .A(n35981), .B(n35980), .Z(n35955) );
  XOR U215 ( .A(n36122), .B(n36121), .Z(n36123) );
  XOR U216 ( .A(n36163), .B(n36162), .Z(n36165) );
  XNOR U217 ( .A(n36135), .B(n36134), .Z(n36128) );
  XOR U218 ( .A(n36414), .B(n36413), .Z(n36415) );
  XNOR U219 ( .A(n36446), .B(n36445), .Z(n36484) );
  XOR U220 ( .A(n36468), .B(n36467), .Z(n36489) );
  XOR U221 ( .A(n36552), .B(n36551), .Z(n36553) );
  XNOR U222 ( .A(n36560), .B(n36559), .Z(n36528) );
  XOR U223 ( .A(n36713), .B(n36712), .Z(n36714) );
  XOR U224 ( .A(n36652), .B(n36651), .Z(n36654) );
  XOR U225 ( .A(n36821), .B(n36820), .Z(n36822) );
  XOR U226 ( .A(n36798), .B(n36797), .Z(n36847) );
  XOR U227 ( .A(n36960), .B(n36959), .Z(n36962) );
  XOR U228 ( .A(n36966), .B(n36965), .Z(n36967) );
  XOR U229 ( .A(n36926), .B(n36925), .Z(n36927) );
  XNOR U230 ( .A(n36934), .B(n36933), .Z(n36979) );
  NANDN U231 ( .A(n36803), .B(n36802), .Z(n13) );
  NANDN U232 ( .A(n36937), .B(n36801), .Z(n14) );
  NAND U233 ( .A(n13), .B(n14), .Z(n36986) );
  XOR U234 ( .A(n37184), .B(n37183), .Z(n37187) );
  XOR U235 ( .A(n37268), .B(n37267), .Z(n37269) );
  XOR U236 ( .A(n37395), .B(n37394), .Z(n37396) );
  XOR U237 ( .A(n37490), .B(n37489), .Z(n37491) );
  XOR U238 ( .A(n37496), .B(n37495), .Z(n37497) );
  XOR U239 ( .A(n37593), .B(n37592), .Z(n37594) );
  XOR U240 ( .A(n37659), .B(n37658), .Z(n37660) );
  XOR U241 ( .A(n37762), .B(n37761), .Z(n37763) );
  XNOR U242 ( .A(n35553), .B(n35552), .Z(n35604) );
  XOR U243 ( .A(n35611), .B(n35610), .Z(n35612) );
  XOR U244 ( .A(n35800), .B(n35799), .Z(n35802) );
  XOR U245 ( .A(n35949), .B(n35948), .Z(n35950) );
  XOR U246 ( .A(n36056), .B(n36055), .Z(n35943) );
  XOR U247 ( .A(n36191), .B(n36190), .Z(n36086) );
  XOR U248 ( .A(n36337), .B(n36336), .Z(n36339) );
  XOR U249 ( .A(n36227), .B(n36226), .Z(n36228) );
  XOR U250 ( .A(n36233), .B(n36232), .Z(n36234) );
  XNOR U251 ( .A(n36480), .B(n36479), .Z(n36472) );
  XOR U252 ( .A(n36524), .B(n36523), .Z(n36540) );
  XOR U253 ( .A(n36972), .B(n36971), .Z(n36974) );
  XOR U254 ( .A(n36872), .B(n36871), .Z(n36873) );
  XOR U255 ( .A(n36990), .B(n36989), .Z(n36991) );
  XNOR U256 ( .A(n37065), .B(n37064), .Z(n37033) );
  XNOR U257 ( .A(n37054), .B(n37053), .Z(n37041) );
  XOR U258 ( .A(n37048), .B(n37047), .Z(n37027) );
  XNOR U259 ( .A(n37202), .B(n37201), .Z(n37194) );
  XOR U260 ( .A(n37218), .B(n37217), .Z(n37220) );
  XNOR U261 ( .A(n37258), .B(n37257), .Z(n37244) );
  XOR U262 ( .A(n37264), .B(n37263), .Z(n37249) );
  NAND U263 ( .A(n37290), .B(n37289), .Z(n15) );
  NANDN U264 ( .A(n37389), .B(n37288), .Z(n16) );
  AND U265 ( .A(n15), .B(n16), .Z(n37403) );
  XNOR U266 ( .A(n37360), .B(n37359), .Z(n37432) );
  XNOR U267 ( .A(n37601), .B(n37600), .Z(n37547) );
  XNOR U268 ( .A(n37667), .B(n37666), .Z(n37670) );
  XOR U269 ( .A(n37734), .B(n37733), .Z(n37736) );
  XNOR U270 ( .A(n37758), .B(n37757), .Z(n37782) );
  NAND U271 ( .A(n37678), .B(n37677), .Z(n17) );
  NANDN U272 ( .A(n37767), .B(n37676), .Z(n18) );
  NAND U273 ( .A(n17), .B(n18), .Z(n37791) );
  XOR U274 ( .A(n37861), .B(n37860), .Z(n37862) );
  XOR U275 ( .A(n37845), .B(n37844), .Z(n37854) );
  XOR U276 ( .A(n37911), .B(n37910), .Z(n37912) );
  XOR U277 ( .A(n38050), .B(n38049), .Z(n38052) );
  XNOR U278 ( .A(n38128), .B(n38127), .Z(n38119) );
  XOR U279 ( .A(n38232), .B(n38231), .Z(n38233) );
  XOR U280 ( .A(n38281), .B(n38280), .Z(n38283) );
  XNOR U281 ( .A(n35768), .B(n35767), .Z(n35647) );
  XNOR U282 ( .A(n35919), .B(n35918), .Z(n35795) );
  XNOR U283 ( .A(n36383), .B(n36382), .Z(n36374) );
  XOR U284 ( .A(n36512), .B(n36511), .Z(n36622) );
  XOR U285 ( .A(n36746), .B(n36745), .Z(n36747) );
  XOR U286 ( .A(n36634), .B(n36633), .Z(n36635) );
  XOR U287 ( .A(n37466), .B(n37465), .Z(n37451) );
  XOR U288 ( .A(n37617), .B(n37616), .Z(n37618) );
  XOR U289 ( .A(n37540), .B(n37539), .Z(n37542) );
  XOR U290 ( .A(n37893), .B(n37892), .Z(n37895) );
  XOR U291 ( .A(n38008), .B(n38007), .Z(n38013) );
  XOR U292 ( .A(n38193), .B(n38192), .Z(n38208) );
  XOR U293 ( .A(n38275), .B(n38274), .Z(n38276) );
  XOR U294 ( .A(n35774), .B(n35773), .Z(n35633) );
  XOR U295 ( .A(n36066), .B(n36065), .Z(n36067) );
  XOR U296 ( .A(n36207), .B(n36206), .Z(n36208) );
  XOR U297 ( .A(n36221), .B(n36220), .Z(n36222) );
  XNOR U298 ( .A(n36774), .B(n36773), .Z(n36766) );
  XOR U299 ( .A(n36886), .B(n36885), .Z(n36887) );
  XOR U300 ( .A(n37124), .B(n37123), .Z(n37125) );
  XNOR U301 ( .A(n37322), .B(n37321), .Z(n37325) );
  XOR U302 ( .A(n37348), .B(n37347), .Z(n37339) );
  XOR U303 ( .A(n37446), .B(n37445), .Z(n37447) );
  XNOR U304 ( .A(n37645), .B(n37644), .Z(n37637) );
  XOR U305 ( .A(n37722), .B(n37721), .Z(n37723) );
  XOR U306 ( .A(n38020), .B(n38019), .Z(n37965) );
  XNOR U307 ( .A(n38040), .B(n38039), .Z(n38032) );
  XNOR U308 ( .A(n38110), .B(n38109), .Z(n38101) );
  XOR U309 ( .A(n38162), .B(n38161), .Z(n38163) );
  NAND U310 ( .A(n38229), .B(n38230), .Z(n19) );
  XOR U311 ( .A(n38229), .B(n38230), .Z(n20) );
  NANDN U312 ( .A(n38228), .B(n20), .Z(n21) );
  NAND U313 ( .A(n19), .B(n21), .Z(n38271) );
  XOR U314 ( .A(n38322), .B(n38321), .Z(n38323) );
  XOR U315 ( .A(n38391), .B(n38390), .Z(n38392) );
  XOR U316 ( .A(n38405), .B(n38404), .Z(n38406) );
  XOR U317 ( .A(n38435), .B(n38434), .Z(n38436) );
  NANDN U318 ( .A(n247), .B(n246), .Z(n22) );
  NANDN U319 ( .A(n244), .B(n245), .Z(n23) );
  AND U320 ( .A(n22), .B(n23), .Z(n280) );
  XOR U321 ( .A(n35788), .B(n35787), .Z(n35789) );
  XOR U322 ( .A(n36365), .B(n36364), .Z(n36356) );
  XOR U323 ( .A(n37012), .B(n37011), .Z(n37003) );
  XOR U324 ( .A(n37811), .B(n37810), .Z(n37802) );
  XOR U325 ( .A(n37889), .B(n37888), .Z(n37880) );
  XOR U326 ( .A(n38225), .B(n38224), .Z(n38216) );
  XOR U327 ( .A(n38479), .B(n38478), .Z(n38480) );
  XOR U328 ( .A(n38510), .B(n38511), .Z(n38513) );
  NAND U329 ( .A(b[0]), .B(a[233]), .Z(n24) );
  XNOR U330 ( .A(b[1]), .B(n24), .Z(n25) );
  NANDN U331 ( .A(b[0]), .B(a[232]), .Z(n26) );
  AND U332 ( .A(n25), .B(n26), .Z(n32540) );
  XOR U333 ( .A(n35366), .B(n35365), .Z(n35367) );
  XOR U334 ( .A(n35587), .B(n35586), .Z(n35588) );
  XOR U335 ( .A(n35593), .B(n35592), .Z(n35594) );
  XOR U336 ( .A(n35973), .B(n35972), .Z(n35974) );
  XOR U337 ( .A(n36036), .B(n36035), .Z(n36037) );
  XOR U338 ( .A(n35979), .B(n35978), .Z(n35980) );
  XOR U339 ( .A(n36092), .B(n36091), .Z(n36093) );
  XOR U340 ( .A(n36253), .B(n36254), .Z(n36255) );
  XOR U341 ( .A(n36331), .B(n36330), .Z(n36332) );
  XOR U342 ( .A(n36266), .B(n36265), .Z(n36267) );
  XOR U343 ( .A(n36272), .B(n36271), .Z(n36273) );
  XOR U344 ( .A(n36444), .B(n36443), .Z(n36445) );
  XOR U345 ( .A(n36387), .B(n36386), .Z(n36388) );
  XOR U346 ( .A(n36583), .B(n36582), .Z(n36584) );
  XOR U347 ( .A(n36695), .B(n36694), .Z(n36697) );
  XOR U348 ( .A(n36790), .B(n36789), .Z(n36791) );
  XOR U349 ( .A(n36932), .B(n36931), .Z(n36933) );
  NANDN U350 ( .A(n2293), .B(n2294), .Z(n27) );
  NANDN U351 ( .A(n2292), .B(n2291), .Z(n28) );
  NAND U352 ( .A(n27), .B(n28), .Z(n2483) );
  NANDN U353 ( .A(n3357), .B(n3356), .Z(n29) );
  NANDN U354 ( .A(n3358), .B(n3359), .Z(n30) );
  AND U355 ( .A(n29), .B(n30), .Z(n3552) );
  NANDN U356 ( .A(n3492), .B(n3491), .Z(n31) );
  NANDN U357 ( .A(n3493), .B(n3494), .Z(n32) );
  AND U358 ( .A(n31), .B(n32), .Z(n3705) );
  NANDN U359 ( .A(n3645), .B(n3644), .Z(n33) );
  NANDN U360 ( .A(n3646), .B(n3647), .Z(n34) );
  AND U361 ( .A(n33), .B(n34), .Z(n3854) );
  NANDN U362 ( .A(n4102), .B(n4101), .Z(n35) );
  NANDN U363 ( .A(n4103), .B(n4104), .Z(n36) );
  AND U364 ( .A(n35), .B(n36), .Z(n4299) );
  NANDN U365 ( .A(n4994), .B(n4993), .Z(n37) );
  NANDN U366 ( .A(n4995), .B(n4996), .Z(n38) );
  AND U367 ( .A(n37), .B(n38), .Z(n5183) );
  NANDN U368 ( .A(n5123), .B(n5122), .Z(n39) );
  NANDN U369 ( .A(n5124), .B(n5125), .Z(n40) );
  AND U370 ( .A(n39), .B(n40), .Z(n5338) );
  NANDN U371 ( .A(n5586), .B(n5585), .Z(n41) );
  NANDN U372 ( .A(n5587), .B(n5588), .Z(n42) );
  AND U373 ( .A(n41), .B(n42), .Z(n5777) );
  NANDN U374 ( .A(n6180), .B(n6179), .Z(n43) );
  NANDN U375 ( .A(n6181), .B(n6182), .Z(n44) );
  AND U376 ( .A(n43), .B(n44), .Z(n6377) );
  NANDN U377 ( .A(n6917), .B(n6916), .Z(n45) );
  NANDN U378 ( .A(n6918), .B(n6919), .Z(n46) );
  AND U379 ( .A(n45), .B(n46), .Z(n7114) );
  NANDN U380 ( .A(n7964), .B(n7963), .Z(n47) );
  NANDN U381 ( .A(n7965), .B(n7966), .Z(n48) );
  AND U382 ( .A(n47), .B(n48), .Z(n8155) );
  NANDN U383 ( .A(n9303), .B(n9302), .Z(n49) );
  NANDN U384 ( .A(n9304), .B(n9305), .Z(n50) );
  AND U385 ( .A(n49), .B(n50), .Z(n9492) );
  NANDN U386 ( .A(n9432), .B(n9431), .Z(n51) );
  NANDN U387 ( .A(n9433), .B(n9434), .Z(n52) );
  AND U388 ( .A(n51), .B(n52), .Z(n9645) );
  NANDN U389 ( .A(n9585), .B(n9584), .Z(n53) );
  NANDN U390 ( .A(n9586), .B(n9587), .Z(n54) );
  AND U391 ( .A(n53), .B(n54), .Z(n9792) );
  NANDN U392 ( .A(n9732), .B(n9731), .Z(n55) );
  NANDN U393 ( .A(n9733), .B(n9734), .Z(n56) );
  AND U394 ( .A(n55), .B(n56), .Z(n9941) );
  NANDN U395 ( .A(n10040), .B(n10039), .Z(n57) );
  NANDN U396 ( .A(n10041), .B(n10042), .Z(n58) );
  AND U397 ( .A(n57), .B(n58), .Z(n10229) );
  NANDN U398 ( .A(n10169), .B(n10168), .Z(n59) );
  NANDN U399 ( .A(n10170), .B(n10171), .Z(n60) );
  AND U400 ( .A(n59), .B(n60), .Z(n10382) );
  NANDN U401 ( .A(n10322), .B(n10321), .Z(n61) );
  NANDN U402 ( .A(n10323), .B(n10324), .Z(n62) );
  AND U403 ( .A(n61), .B(n62), .Z(n10529) );
  NANDN U404 ( .A(n10469), .B(n10468), .Z(n63) );
  NANDN U405 ( .A(n10470), .B(n10471), .Z(n64) );
  AND U406 ( .A(n63), .B(n64), .Z(n10678) );
  NANDN U407 ( .A(n10777), .B(n10776), .Z(n65) );
  NANDN U408 ( .A(n10778), .B(n10779), .Z(n66) );
  AND U409 ( .A(n65), .B(n66), .Z(n10966) );
  NANDN U410 ( .A(n10906), .B(n10905), .Z(n67) );
  NANDN U411 ( .A(n10907), .B(n10908), .Z(n68) );
  AND U412 ( .A(n67), .B(n68), .Z(n11121) );
  NANDN U413 ( .A(n11369), .B(n11368), .Z(n69) );
  NANDN U414 ( .A(n11370), .B(n11371), .Z(n70) );
  AND U415 ( .A(n69), .B(n70), .Z(n11558) );
  NANDN U416 ( .A(n11498), .B(n11497), .Z(n71) );
  NANDN U417 ( .A(n11499), .B(n11500), .Z(n72) );
  AND U418 ( .A(n71), .B(n72), .Z(n11711) );
  NANDN U419 ( .A(n11651), .B(n11650), .Z(n73) );
  NANDN U420 ( .A(n11652), .B(n11653), .Z(n74) );
  AND U421 ( .A(n73), .B(n74), .Z(n11860) );
  NANDN U422 ( .A(n11959), .B(n11958), .Z(n75) );
  NANDN U423 ( .A(n11960), .B(n11961), .Z(n76) );
  AND U424 ( .A(n75), .B(n76), .Z(n12150) );
  NANDN U425 ( .A(n12702), .B(n12701), .Z(n77) );
  NANDN U426 ( .A(n12703), .B(n12704), .Z(n78) );
  AND U427 ( .A(n77), .B(n78), .Z(n12893) );
  NANDN U428 ( .A(n15829), .B(n15828), .Z(n79) );
  NANDN U429 ( .A(n15830), .B(n15831), .Z(n80) );
  AND U430 ( .A(n79), .B(n80), .Z(n16020) );
  NANDN U431 ( .A(n16125), .B(n16124), .Z(n81) );
  NANDN U432 ( .A(n16126), .B(n16127), .Z(n82) );
  AND U433 ( .A(n81), .B(n82), .Z(n16316) );
  NANDN U434 ( .A(n17160), .B(n17159), .Z(n83) );
  NANDN U435 ( .A(n17161), .B(n17162), .Z(n84) );
  AND U436 ( .A(n83), .B(n84), .Z(n17357) );
  NANDN U437 ( .A(n17611), .B(n17610), .Z(n85) );
  NANDN U438 ( .A(n17612), .B(n17613), .Z(n86) );
  AND U439 ( .A(n85), .B(n86), .Z(n17800) );
  NANDN U440 ( .A(n17740), .B(n17739), .Z(n87) );
  NANDN U441 ( .A(n17741), .B(n17742), .Z(n88) );
  AND U442 ( .A(n87), .B(n88), .Z(n17955) );
  NANDN U443 ( .A(n18197), .B(n18196), .Z(n89) );
  NANDN U444 ( .A(n18198), .B(n18199), .Z(n90) );
  AND U445 ( .A(n89), .B(n90), .Z(n18400) );
  NANDN U446 ( .A(n19095), .B(n19094), .Z(n91) );
  NANDN U447 ( .A(n19096), .B(n19097), .Z(n92) );
  AND U448 ( .A(n91), .B(n92), .Z(n19292) );
  NANDN U449 ( .A(n19391), .B(n19390), .Z(n93) );
  NANDN U450 ( .A(n19392), .B(n19393), .Z(n94) );
  AND U451 ( .A(n93), .B(n94), .Z(n19588) );
  NANDN U452 ( .A(n19985), .B(n19984), .Z(n95) );
  NANDN U453 ( .A(n19986), .B(n19987), .Z(n96) );
  AND U454 ( .A(n95), .B(n96), .Z(n20182) );
  NANDN U455 ( .A(n20579), .B(n20578), .Z(n97) );
  NANDN U456 ( .A(n20580), .B(n20581), .Z(n98) );
  AND U457 ( .A(n97), .B(n98), .Z(n20768) );
  NANDN U458 ( .A(n20708), .B(n20707), .Z(n99) );
  NANDN U459 ( .A(n20709), .B(n20710), .Z(n100) );
  AND U460 ( .A(n99), .B(n100), .Z(n20923) );
  NANDN U461 ( .A(n21022), .B(n21021), .Z(n101) );
  NANDN U462 ( .A(n21023), .B(n21024), .Z(n102) );
  AND U463 ( .A(n101), .B(n102), .Z(n21213) );
  NANDN U464 ( .A(n21765), .B(n21764), .Z(n103) );
  NANDN U465 ( .A(n21766), .B(n21767), .Z(n104) );
  AND U466 ( .A(n103), .B(n104), .Z(n21962) );
  NANDN U467 ( .A(n22210), .B(n22209), .Z(n105) );
  NANDN U468 ( .A(n22211), .B(n22212), .Z(n106) );
  AND U469 ( .A(n105), .B(n106), .Z(n22401) );
  NANDN U470 ( .A(n23394), .B(n23393), .Z(n107) );
  NANDN U471 ( .A(n23395), .B(n23396), .Z(n108) );
  AND U472 ( .A(n107), .B(n108), .Z(n23589) );
  NANDN U473 ( .A(n23529), .B(n23528), .Z(n109) );
  NANDN U474 ( .A(n23530), .B(n23531), .Z(n110) );
  AND U475 ( .A(n109), .B(n110), .Z(n23744) );
  NANDN U476 ( .A(n23843), .B(n23842), .Z(n111) );
  NANDN U477 ( .A(n23844), .B(n23845), .Z(n112) );
  AND U478 ( .A(n111), .B(n112), .Z(n24040) );
  NANDN U479 ( .A(n24139), .B(n24138), .Z(n113) );
  NANDN U480 ( .A(n24140), .B(n24141), .Z(n114) );
  AND U481 ( .A(n113), .B(n114), .Z(n24328) );
  NANDN U482 ( .A(n24268), .B(n24267), .Z(n115) );
  NANDN U483 ( .A(n24269), .B(n24270), .Z(n116) );
  AND U484 ( .A(n115), .B(n116), .Z(n24481) );
  NANDN U485 ( .A(n24421), .B(n24420), .Z(n117) );
  NANDN U486 ( .A(n24422), .B(n24423), .Z(n118) );
  AND U487 ( .A(n117), .B(n118), .Z(n24630) );
  NANDN U488 ( .A(n24878), .B(n24877), .Z(n119) );
  NANDN U489 ( .A(n24879), .B(n24880), .Z(n120) );
  AND U490 ( .A(n119), .B(n120), .Z(n25069) );
  NANDN U491 ( .A(n25919), .B(n25918), .Z(n121) );
  NANDN U492 ( .A(n25920), .B(n25921), .Z(n122) );
  AND U493 ( .A(n121), .B(n122), .Z(n26108) );
  NANDN U494 ( .A(n26048), .B(n26047), .Z(n123) );
  NANDN U495 ( .A(n26049), .B(n26050), .Z(n124) );
  AND U496 ( .A(n123), .B(n124), .Z(n26263) );
  NANDN U497 ( .A(n26958), .B(n26957), .Z(n125) );
  NANDN U498 ( .A(n26959), .B(n26960), .Z(n126) );
  AND U499 ( .A(n125), .B(n126), .Z(n27155) );
  NANDN U500 ( .A(n28595), .B(n28594), .Z(n127) );
  NANDN U501 ( .A(n28596), .B(n28597), .Z(n128) );
  AND U502 ( .A(n127), .B(n128), .Z(n28790) );
  NANDN U503 ( .A(n28730), .B(n28729), .Z(n129) );
  NANDN U504 ( .A(n28731), .B(n28732), .Z(n130) );
  AND U505 ( .A(n129), .B(n130), .Z(n28939) );
  NANDN U506 ( .A(n29187), .B(n29186), .Z(n131) );
  NANDN U507 ( .A(n29188), .B(n29189), .Z(n132) );
  AND U508 ( .A(n131), .B(n132), .Z(n29382) );
  NANDN U509 ( .A(n29322), .B(n29321), .Z(n133) );
  NANDN U510 ( .A(n29323), .B(n29324), .Z(n134) );
  AND U511 ( .A(n133), .B(n134), .Z(n29529) );
  NANDN U512 ( .A(n29469), .B(n29468), .Z(n135) );
  NANDN U513 ( .A(n29470), .B(n29471), .Z(n136) );
  AND U514 ( .A(n135), .B(n136), .Z(n29678) );
  NANDN U515 ( .A(n29777), .B(n29776), .Z(n137) );
  NANDN U516 ( .A(n29778), .B(n29779), .Z(n138) );
  AND U517 ( .A(n137), .B(n138), .Z(n29974) );
  NANDN U518 ( .A(n30669), .B(n30668), .Z(n139) );
  NANDN U519 ( .A(n30670), .B(n30671), .Z(n140) );
  AND U520 ( .A(n139), .B(n140), .Z(n30864) );
  NANDN U521 ( .A(n30804), .B(n30803), .Z(n141) );
  NANDN U522 ( .A(n30805), .B(n30806), .Z(n142) );
  AND U523 ( .A(n141), .B(n142), .Z(n31011) );
  NANDN U524 ( .A(n30951), .B(n30950), .Z(n143) );
  NANDN U525 ( .A(n30952), .B(n30953), .Z(n144) );
  AND U526 ( .A(n143), .B(n144), .Z(n31158) );
  NANDN U527 ( .A(n31098), .B(n31097), .Z(n145) );
  NANDN U528 ( .A(n31099), .B(n31100), .Z(n146) );
  AND U529 ( .A(n145), .B(n146), .Z(n31307) );
  NANDN U530 ( .A(n31852), .B(n31851), .Z(n147) );
  NANDN U531 ( .A(n31853), .B(n31854), .Z(n148) );
  AND U532 ( .A(n147), .B(n148), .Z(n32044) );
  NANDN U533 ( .A(n32593), .B(n32592), .Z(n149) );
  NANDN U534 ( .A(n32594), .B(n32595), .Z(n150) );
  AND U535 ( .A(n149), .B(n150), .Z(n32784) );
  NANDN U536 ( .A(n33932), .B(n33931), .Z(n151) );
  NANDN U537 ( .A(n33933), .B(n33934), .Z(n152) );
  AND U538 ( .A(n151), .B(n152), .Z(n34129) );
  XOR U539 ( .A(n35402), .B(n35401), .Z(n35404) );
  XNOR U540 ( .A(n35464), .B(n35463), .Z(n35408) );
  XOR U541 ( .A(n35470), .B(n35469), .Z(n35425) );
  XNOR U542 ( .A(n35541), .B(n35540), .Z(n35498) );
  XOR U543 ( .A(n35658), .B(n35657), .Z(n35659) );
  XNOR U544 ( .A(n35744), .B(n35743), .Z(n35652) );
  XOR U545 ( .A(n35899), .B(n35898), .Z(n35900) );
  XNOR U546 ( .A(n35853), .B(n35852), .Z(n35857) );
  XOR U547 ( .A(n36048), .B(n36047), .Z(n36049) );
  XOR U548 ( .A(n36116), .B(n36115), .Z(n36117) );
  XNOR U549 ( .A(n36262), .B(n36261), .Z(n36284) );
  XNOR U550 ( .A(n36185), .B(n36184), .Z(n36157) );
  XNOR U551 ( .A(n36416), .B(n36415), .Z(n36419) );
  XNOR U552 ( .A(n36492), .B(n36491), .Z(n36380) );
  XOR U553 ( .A(n36740), .B(n36739), .Z(n36741) );
  XOR U554 ( .A(n36703), .B(n36702), .Z(n36712) );
  NANDN U555 ( .A(n36565), .B(n36564), .Z(n153) );
  NANDN U556 ( .A(n36724), .B(n36563), .Z(n154) );
  NAND U557 ( .A(n153), .B(n154), .Z(n36660) );
  XOR U558 ( .A(n36848), .B(n36847), .Z(n36849) );
  XOR U559 ( .A(n37104), .B(n37103), .Z(n37105) );
  XOR U560 ( .A(n37052), .B(n37051), .Z(n37053) );
  XOR U561 ( .A(n37182), .B(n37181), .Z(n37183) );
  XOR U562 ( .A(n37142), .B(n37141), .Z(n37144) );
  XOR U563 ( .A(n37212), .B(n37211), .Z(n37213) );
  XOR U564 ( .A(n37200), .B(n37199), .Z(n37201) );
  XOR U565 ( .A(n37262), .B(n37261), .Z(n37263) );
  XOR U566 ( .A(n37256), .B(n37255), .Z(n37257) );
  NAND U567 ( .A(n37305), .B(n38185), .Z(n155) );
  NANDN U568 ( .A(n37306), .B(n37375), .Z(n156) );
  AND U569 ( .A(n155), .B(n156), .Z(n37409) );
  XOR U570 ( .A(n37504), .B(n37503), .Z(n37495) );
  XOR U571 ( .A(n37665), .B(n37664), .Z(n37666) );
  NANDN U572 ( .A(n2089), .B(n2088), .Z(n157) );
  NANDN U573 ( .A(n2090), .B(n2091), .Z(n158) );
  AND U574 ( .A(n157), .B(n158), .Z(n2210) );
  XOR U575 ( .A(n35599), .B(n35598), .Z(n35600) );
  XOR U576 ( .A(n35754), .B(n35753), .Z(n35755) );
  XOR U577 ( .A(n35760), .B(n35759), .Z(n35761) );
  XNOR U578 ( .A(n35708), .B(n35707), .Z(n35765) );
  XOR U579 ( .A(n35911), .B(n35910), .Z(n35912) );
  XOR U580 ( .A(n35905), .B(n35904), .Z(n35906) );
  XOR U581 ( .A(n36054), .B(n36053), .Z(n36055) );
  XNOR U582 ( .A(n36002), .B(n36001), .Z(n35942) );
  XOR U583 ( .A(n36195), .B(n36194), .Z(n36196) );
  XOR U584 ( .A(n36554), .B(n36553), .Z(n36546) );
  XOR U585 ( .A(n36534), .B(n36533), .Z(n36535) );
  XOR U586 ( .A(n36510), .B(n36509), .Z(n36511) );
  XOR U587 ( .A(n36707), .B(n36706), .Z(n36709) );
  XOR U588 ( .A(n36646), .B(n36645), .Z(n36647) );
  XOR U589 ( .A(n36640), .B(n36639), .Z(n36641) );
  XNOR U590 ( .A(n36862), .B(n36861), .Z(n36783) );
  XOR U591 ( .A(n37028), .B(n37027), .Z(n37030) );
  XOR U592 ( .A(n37110), .B(n37109), .Z(n37111) );
  XOR U593 ( .A(n37136), .B(n37135), .Z(n37137) );
  XOR U594 ( .A(n37432), .B(n37431), .Z(n37434) );
  XOR U595 ( .A(n37458), .B(n37457), .Z(n37459) );
  NAND U596 ( .A(n37518), .B(n37517), .Z(n159) );
  NANDN U597 ( .A(n37551), .B(n37516), .Z(n160) );
  AND U598 ( .A(n159), .B(n160), .Z(n37606) );
  XOR U599 ( .A(n37611), .B(n37610), .Z(n37613) );
  XNOR U600 ( .A(n37661), .B(n37660), .Z(n37672) );
  XOR U601 ( .A(n37702), .B(n37701), .Z(n37704) );
  XOR U602 ( .A(n37855), .B(n37854), .Z(n37856) );
  XOR U603 ( .A(n37905), .B(n37904), .Z(n37907) );
  XOR U604 ( .A(n37972), .B(n37971), .Z(n37973) );
  XOR U605 ( .A(n38006), .B(n38005), .Z(n38007) );
  XOR U606 ( .A(n38082), .B(n38081), .Z(n38084) );
  XNOR U607 ( .A(n38150), .B(n38149), .Z(n38121) );
  NANDN U608 ( .A(n772), .B(n773), .Z(n161) );
  NANDN U609 ( .A(n771), .B(n770), .Z(n162) );
  NAND U610 ( .A(n161), .B(n162), .Z(n796) );
  NANDN U611 ( .A(n1892), .B(n1891), .Z(n163) );
  NANDN U612 ( .A(n1893), .B(n1894), .Z(n164) );
  AND U613 ( .A(n163), .B(n164), .Z(n2116) );
  XOR U614 ( .A(n35613), .B(n35612), .Z(n35491) );
  XOR U615 ( .A(n35640), .B(n35639), .Z(n35642) );
  XOR U616 ( .A(n36060), .B(n36059), .Z(n36062) );
  XNOR U617 ( .A(n36088), .B(n36087), .Z(n36202) );
  XNOR U618 ( .A(n36229), .B(n36228), .Z(n36342) );
  XOR U619 ( .A(n36349), .B(n36348), .Z(n36350) );
  XNOR U620 ( .A(n36474), .B(n36473), .Z(n36376) );
  XNOR U621 ( .A(n36874), .B(n36873), .Z(n36779) );
  XOR U622 ( .A(n36996), .B(n36995), .Z(n36997) );
  XNOR U623 ( .A(n36992), .B(n36991), .Z(n36891) );
  XOR U624 ( .A(n37036), .B(n37035), .Z(n37022) );
  XOR U625 ( .A(n37224), .B(n37223), .Z(n37225) );
  XOR U626 ( .A(n37310), .B(n37309), .Z(n37240) );
  XOR U627 ( .A(n37352), .B(n37351), .Z(n37354) );
  XOR U628 ( .A(n37346), .B(n37345), .Z(n37347) );
  XOR U629 ( .A(n37452), .B(n37451), .Z(n37453) );
  XOR U630 ( .A(n37698), .B(n37697), .Z(n37707) );
  XOR U631 ( .A(n37791), .B(n37790), .Z(n37794) );
  XOR U632 ( .A(n37873), .B(n37872), .Z(n37875) );
  XOR U633 ( .A(n37815), .B(n37814), .Z(n37816) );
  XOR U634 ( .A(n37899), .B(n37898), .Z(n37900) );
  XOR U635 ( .A(n38012), .B(n38011), .Z(n38014) );
  XOR U636 ( .A(n38114), .B(n38113), .Z(n38116) );
  XNOR U637 ( .A(n38211), .B(n38210), .Z(n38167) );
  XNOR U638 ( .A(n38234), .B(n38233), .Z(n38255) );
  XOR U639 ( .A(n38308), .B(n38307), .Z(n38309) );
  XOR U640 ( .A(n38334), .B(n38333), .Z(n38335) );
  XOR U641 ( .A(n38368), .B(n38367), .Z(n38370) );
  NAND U642 ( .A(n1325), .B(n1324), .Z(n165) );
  NANDN U643 ( .A(n1322), .B(n1323), .Z(n166) );
  AND U644 ( .A(n165), .B(n166), .Z(n1509) );
  XOR U645 ( .A(n35923), .B(n35922), .Z(n35924) );
  XNOR U646 ( .A(n36068), .B(n36067), .Z(n35930) );
  XNOR U647 ( .A(n36768), .B(n36767), .Z(n36759) );
  XOR U648 ( .A(n36888), .B(n36887), .Z(n36879) );
  XNOR U649 ( .A(n37639), .B(n37638), .Z(n37630) );
  XOR U650 ( .A(n37724), .B(n37723), .Z(n37715) );
  XOR U651 ( .A(n38104), .B(n38103), .Z(n38095) );
  XNOR U652 ( .A(n38407), .B(n38406), .Z(n38398) );
  XOR U653 ( .A(n234), .B(n232), .Z(n167) );
  NANDN U654 ( .A(n233), .B(n167), .Z(n168) );
  NAND U655 ( .A(n234), .B(n232), .Z(n169) );
  AND U656 ( .A(n168), .B(n169), .Z(n247) );
  XOR U657 ( .A(n35790), .B(n35789), .Z(n35782) );
  XOR U658 ( .A(n36074), .B(n36073), .Z(n36075) );
  XOR U659 ( .A(n36215), .B(n36214), .Z(n36216) );
  XOR U660 ( .A(n36357), .B(n36356), .Z(n36358) );
  XOR U661 ( .A(n36498), .B(n36497), .Z(n36499) );
  XOR U662 ( .A(n36628), .B(n36627), .Z(n36629) );
  XOR U663 ( .A(n37004), .B(n37003), .Z(n37005) );
  XOR U664 ( .A(n37118), .B(n37117), .Z(n37119) );
  XOR U665 ( .A(n37232), .B(n37231), .Z(n37233) );
  XOR U666 ( .A(n37334), .B(n37333), .Z(n37335) );
  XOR U667 ( .A(n37534), .B(n37533), .Z(n37535) );
  XOR U668 ( .A(n37803), .B(n37802), .Z(n37804) );
  XOR U669 ( .A(n37881), .B(n37880), .Z(n37882) );
  XOR U670 ( .A(n37960), .B(n37959), .Z(n37961) );
  XOR U671 ( .A(n38026), .B(n38025), .Z(n38027) );
  XOR U672 ( .A(n38156), .B(n38155), .Z(n38157) );
  XOR U673 ( .A(n38217), .B(n38216), .Z(n38218) );
  XOR U674 ( .A(n38263), .B(n38262), .Z(n38264) );
  XOR U675 ( .A(n38316), .B(n38315), .Z(n38317) );
  XOR U676 ( .A(n38356), .B(n38355), .Z(n38357) );
  XOR U677 ( .A(n38463), .B(n38462), .Z(n38464) );
  XOR U678 ( .A(n38503), .B(n38502), .Z(n38505) );
  XNOR U679 ( .A(n38523), .B(n38524), .Z(n38512) );
  NAND U680 ( .A(n983), .B(n36922), .Z(n170) );
  NAND U681 ( .A(n698), .B(n1681), .Z(n171) );
  XNOR U682 ( .A(b[1]), .B(b[2]), .Z(n172) );
  NAND U683 ( .A(n283), .B(n622), .Z(n173) );
  NAND U684 ( .A(n1178), .B(n37589), .Z(n174) );
  NAND U685 ( .A(n361), .B(n572), .Z(n175) );
  NAND U686 ( .A(n559), .B(n2434), .Z(n176) );
  NAND U687 ( .A(n2336), .B(n193), .Z(n177) );
  NAND U688 ( .A(n840), .B(n37509), .Z(n178) );
  NAND U689 ( .A(n454), .B(n2052), .Z(n179) );
  NAND U690 ( .A(n235), .B(n172), .Z(n180) );
  IV U691 ( .A(n180), .Z(n181) );
  IV U692 ( .A(n172), .Z(n182) );
  IV U693 ( .A(n173), .Z(n183) );
  IV U694 ( .A(n175), .Z(n184) );
  IV U695 ( .A(n179), .Z(n185) );
  IV U696 ( .A(n176), .Z(n186) );
  IV U697 ( .A(n171), .Z(n187) );
  IV U698 ( .A(n178), .Z(n188) );
  IV U699 ( .A(n170), .Z(n189) );
  IV U700 ( .A(n174), .Z(n190) );
  IV U701 ( .A(n38289), .Z(n191) );
  IV U702 ( .A(n38385), .Z(n192) );
  IV U703 ( .A(n38456), .Z(n193) );
  IV U704 ( .A(n177), .Z(n194) );
  IV U705 ( .A(n38470), .Z(n195) );
  AND U706 ( .A(b[0]), .B(a[0]), .Z(n197) );
  XOR U707 ( .A(n197), .B(sreg[224]), .Z(c[224]) );
  AND U708 ( .A(b[0]), .B(a[1]), .Z(n207) );
  NAND U709 ( .A(a[0]), .B(b[1]), .Z(n196) );
  XOR U710 ( .A(n207), .B(n196), .Z(n198) );
  XNOR U711 ( .A(sreg[225]), .B(n198), .Z(n200) );
  AND U712 ( .A(n197), .B(sreg[224]), .Z(n199) );
  XOR U713 ( .A(n200), .B(n199), .Z(c[225]) );
  NANDN U714 ( .A(n198), .B(sreg[225]), .Z(n202) );
  NAND U715 ( .A(n200), .B(n199), .Z(n201) );
  AND U716 ( .A(n202), .B(n201), .Z(n222) );
  XNOR U717 ( .A(n222), .B(sreg[226]), .Z(n224) );
  NAND U718 ( .A(b[0]), .B(a[2]), .Z(n203) );
  XNOR U719 ( .A(b[1]), .B(n203), .Z(n205) );
  NANDN U720 ( .A(b[0]), .B(a[1]), .Z(n204) );
  NAND U721 ( .A(n205), .B(n204), .Z(n211) );
  NAND U722 ( .A(a[0]), .B(b[2]), .Z(n206) );
  XNOR U723 ( .A(b[1]), .B(n206), .Z(n209) );
  NANDN U724 ( .A(a[0]), .B(n207), .Z(n208) );
  NAND U725 ( .A(n209), .B(n208), .Z(n210) );
  XOR U726 ( .A(n211), .B(n210), .Z(n223) );
  XOR U727 ( .A(n224), .B(n223), .Z(c[226]) );
  NOR U728 ( .A(n211), .B(n210), .Z(n234) );
  NAND U729 ( .A(b[0]), .B(a[3]), .Z(n212) );
  XNOR U730 ( .A(b[1]), .B(n212), .Z(n214) );
  NANDN U731 ( .A(b[0]), .B(a[2]), .Z(n213) );
  NAND U732 ( .A(n214), .B(n213), .Z(n242) );
  XOR U733 ( .A(b[3]), .B(b[2]), .Z(n235) );
  XOR U734 ( .A(b[3]), .B(a[0]), .Z(n215) );
  NAND U735 ( .A(n235), .B(n215), .Z(n216) );
  NANDN U736 ( .A(n216), .B(n172), .Z(n218) );
  XOR U737 ( .A(b[3]), .B(a[1]), .Z(n236) );
  NANDN U738 ( .A(n172), .B(n236), .Z(n217) );
  AND U739 ( .A(n218), .B(n217), .Z(n243) );
  XNOR U740 ( .A(n242), .B(n243), .Z(n233) );
  NAND U741 ( .A(n182), .B(a[0]), .Z(n220) );
  NAND U742 ( .A(b[1]), .B(b[2]), .Z(n219) );
  NAND U743 ( .A(b[3]), .B(n219), .Z(n36408) );
  IV U744 ( .A(n36408), .Z(n36302) );
  AND U745 ( .A(n220), .B(n36302), .Z(n232) );
  XOR U746 ( .A(n233), .B(n232), .Z(n221) );
  XOR U747 ( .A(n234), .B(n221), .Z(n227) );
  XNOR U748 ( .A(sreg[227]), .B(n227), .Z(n229) );
  NANDN U749 ( .A(n222), .B(sreg[226]), .Z(n226) );
  NAND U750 ( .A(n224), .B(n223), .Z(n225) );
  NAND U751 ( .A(n226), .B(n225), .Z(n228) );
  XOR U752 ( .A(n229), .B(n228), .Z(c[227]) );
  NANDN U753 ( .A(n227), .B(sreg[227]), .Z(n231) );
  NAND U754 ( .A(n229), .B(n228), .Z(n230) );
  AND U755 ( .A(n231), .B(n230), .Z(n267) );
  XNOR U756 ( .A(n267), .B(sreg[228]), .Z(n269) );
  NAND U757 ( .A(n181), .B(n236), .Z(n238) );
  XOR U758 ( .A(b[3]), .B(a[2]), .Z(n248) );
  NAND U759 ( .A(n182), .B(n248), .Z(n237) );
  AND U760 ( .A(n238), .B(n237), .Z(n264) );
  XNOR U761 ( .A(b[3]), .B(b[4]), .Z(n622) );
  IV U762 ( .A(n622), .Z(n36296) );
  AND U763 ( .A(a[0]), .B(n36296), .Z(n261) );
  NAND U764 ( .A(b[0]), .B(a[4]), .Z(n239) );
  XNOR U765 ( .A(b[1]), .B(n239), .Z(n241) );
  NANDN U766 ( .A(b[0]), .B(a[3]), .Z(n240) );
  NAND U767 ( .A(n241), .B(n240), .Z(n262) );
  XNOR U768 ( .A(n261), .B(n262), .Z(n263) );
  XNOR U769 ( .A(n264), .B(n263), .Z(n245) );
  OR U770 ( .A(n243), .B(n242), .Z(n244) );
  XNOR U771 ( .A(n245), .B(n244), .Z(n246) );
  XNOR U772 ( .A(n247), .B(n246), .Z(n268) );
  XOR U773 ( .A(n269), .B(n268), .Z(c[228]) );
  NAND U774 ( .A(n181), .B(n248), .Z(n250) );
  XOR U775 ( .A(b[3]), .B(a[3]), .Z(n289) );
  NAND U776 ( .A(n182), .B(n289), .Z(n249) );
  AND U777 ( .A(n250), .B(n249), .Z(n296) );
  NAND U778 ( .A(b[3]), .B(b[4]), .Z(n251) );
  AND U779 ( .A(b[5]), .B(n251), .Z(n36572) );
  IV U780 ( .A(n36572), .Z(n36727) );
  NOR U781 ( .A(n36727), .B(n261), .Z(n295) );
  XNOR U782 ( .A(n296), .B(n295), .Z(n298) );
  NAND U783 ( .A(b[0]), .B(a[5]), .Z(n252) );
  XNOR U784 ( .A(b[1]), .B(n252), .Z(n254) );
  NANDN U785 ( .A(b[0]), .B(a[4]), .Z(n253) );
  NAND U786 ( .A(n254), .B(n253), .Z(n287) );
  XOR U787 ( .A(b[5]), .B(a[1]), .Z(n284) );
  NAND U788 ( .A(n36296), .B(n284), .Z(n260) );
  ANDN U789 ( .B(b[4]), .A(b[5]), .Z(n255) );
  NAND U790 ( .A(n255), .B(a[0]), .Z(n257) );
  NANDN U791 ( .A(a[0]), .B(n36572), .Z(n256) );
  NAND U792 ( .A(n257), .B(n256), .Z(n258) );
  NANDN U793 ( .A(n36296), .B(n258), .Z(n259) );
  NAND U794 ( .A(n260), .B(n259), .Z(n288) );
  XNOR U795 ( .A(n287), .B(n288), .Z(n297) );
  XOR U796 ( .A(n298), .B(n297), .Z(n278) );
  NANDN U797 ( .A(n262), .B(n261), .Z(n266) );
  NANDN U798 ( .A(n264), .B(n263), .Z(n265) );
  AND U799 ( .A(n266), .B(n265), .Z(n277) );
  XNOR U800 ( .A(n278), .B(n277), .Z(n279) );
  XOR U801 ( .A(n280), .B(n279), .Z(n272) );
  XNOR U802 ( .A(n272), .B(sreg[229]), .Z(n274) );
  NANDN U803 ( .A(n267), .B(sreg[228]), .Z(n271) );
  NAND U804 ( .A(n269), .B(n268), .Z(n270) );
  NAND U805 ( .A(n271), .B(n270), .Z(n273) );
  XOR U806 ( .A(n274), .B(n273), .Z(c[229]) );
  NANDN U807 ( .A(n272), .B(sreg[229]), .Z(n276) );
  NAND U808 ( .A(n274), .B(n273), .Z(n275) );
  AND U809 ( .A(n276), .B(n275), .Z(n333) );
  XNOR U810 ( .A(n333), .B(sreg[230]), .Z(n335) );
  NANDN U811 ( .A(n278), .B(n277), .Z(n282) );
  NAND U812 ( .A(n280), .B(n279), .Z(n281) );
  AND U813 ( .A(n282), .B(n281), .Z(n303) );
  XOR U814 ( .A(b[4]), .B(b[5]), .Z(n283) );
  NAND U815 ( .A(n183), .B(n284), .Z(n286) );
  XOR U816 ( .A(b[5]), .B(a[2]), .Z(n311) );
  NAND U817 ( .A(n36296), .B(n311), .Z(n285) );
  AND U818 ( .A(n286), .B(n285), .Z(n328) );
  ANDN U819 ( .B(n288), .A(n287), .Z(n327) );
  XNOR U820 ( .A(n328), .B(n327), .Z(n330) );
  NAND U821 ( .A(n181), .B(n289), .Z(n291) );
  XOR U822 ( .A(b[3]), .B(a[4]), .Z(n318) );
  NAND U823 ( .A(n182), .B(n318), .Z(n290) );
  AND U824 ( .A(n291), .B(n290), .Z(n324) );
  XNOR U825 ( .A(b[5]), .B(b[6]), .Z(n572) );
  IV U826 ( .A(n572), .Z(n36592) );
  AND U827 ( .A(a[0]), .B(n36592), .Z(n321) );
  NAND U828 ( .A(b[0]), .B(a[6]), .Z(n292) );
  XNOR U829 ( .A(b[1]), .B(n292), .Z(n294) );
  NANDN U830 ( .A(b[0]), .B(a[5]), .Z(n293) );
  NAND U831 ( .A(n294), .B(n293), .Z(n322) );
  XNOR U832 ( .A(n321), .B(n322), .Z(n323) );
  XNOR U833 ( .A(n324), .B(n323), .Z(n329) );
  XOR U834 ( .A(n330), .B(n329), .Z(n302) );
  NANDN U835 ( .A(n296), .B(n295), .Z(n300) );
  NAND U836 ( .A(n298), .B(n297), .Z(n299) );
  AND U837 ( .A(n300), .B(n299), .Z(n301) );
  XOR U838 ( .A(n302), .B(n301), .Z(n304) );
  XNOR U839 ( .A(n303), .B(n304), .Z(n334) );
  XOR U840 ( .A(n335), .B(n334), .Z(c[230]) );
  NANDN U841 ( .A(n302), .B(n301), .Z(n306) );
  OR U842 ( .A(n304), .B(n303), .Z(n305) );
  AND U843 ( .A(n306), .B(n305), .Z(n345) );
  XOR U844 ( .A(b[7]), .B(b[6]), .Z(n361) );
  XOR U845 ( .A(b[7]), .B(a[0]), .Z(n307) );
  NAND U846 ( .A(n361), .B(n307), .Z(n308) );
  NANDN U847 ( .A(n308), .B(n572), .Z(n310) );
  XOR U848 ( .A(b[7]), .B(a[1]), .Z(n362) );
  NANDN U849 ( .A(n572), .B(n362), .Z(n309) );
  AND U850 ( .A(n310), .B(n309), .Z(n369) );
  NAND U851 ( .A(n183), .B(n311), .Z(n313) );
  XOR U852 ( .A(b[5]), .B(a[3]), .Z(n373) );
  NAND U853 ( .A(n36296), .B(n373), .Z(n312) );
  AND U854 ( .A(n313), .B(n312), .Z(n368) );
  XOR U855 ( .A(n369), .B(n368), .Z(n358) );
  NAND U856 ( .A(b[5]), .B(b[6]), .Z(n314) );
  NAND U857 ( .A(b[7]), .B(n314), .Z(n36939) );
  NOR U858 ( .A(n36939), .B(n321), .Z(n356) );
  NAND U859 ( .A(b[0]), .B(a[7]), .Z(n315) );
  XNOR U860 ( .A(b[1]), .B(n315), .Z(n317) );
  NANDN U861 ( .A(b[0]), .B(a[6]), .Z(n316) );
  NAND U862 ( .A(n317), .B(n316), .Z(n355) );
  XNOR U863 ( .A(n356), .B(n355), .Z(n357) );
  XNOR U864 ( .A(n358), .B(n357), .Z(n349) );
  NANDN U865 ( .A(n180), .B(n318), .Z(n320) );
  XNOR U866 ( .A(b[3]), .B(a[5]), .Z(n365) );
  OR U867 ( .A(n365), .B(n172), .Z(n319) );
  NAND U868 ( .A(n320), .B(n319), .Z(n350) );
  XNOR U869 ( .A(n349), .B(n350), .Z(n351) );
  NANDN U870 ( .A(n322), .B(n321), .Z(n326) );
  NANDN U871 ( .A(n324), .B(n323), .Z(n325) );
  NAND U872 ( .A(n326), .B(n325), .Z(n352) );
  XNOR U873 ( .A(n351), .B(n352), .Z(n343) );
  NANDN U874 ( .A(n328), .B(n327), .Z(n332) );
  NAND U875 ( .A(n330), .B(n329), .Z(n331) );
  NAND U876 ( .A(n332), .B(n331), .Z(n344) );
  XOR U877 ( .A(n343), .B(n344), .Z(n346) );
  XOR U878 ( .A(n345), .B(n346), .Z(n338) );
  XNOR U879 ( .A(n338), .B(sreg[231]), .Z(n340) );
  NANDN U880 ( .A(n333), .B(sreg[230]), .Z(n337) );
  NAND U881 ( .A(n335), .B(n334), .Z(n336) );
  NAND U882 ( .A(n337), .B(n336), .Z(n339) );
  XOR U883 ( .A(n340), .B(n339), .Z(c[231]) );
  NANDN U884 ( .A(n338), .B(sreg[231]), .Z(n342) );
  NAND U885 ( .A(n340), .B(n339), .Z(n341) );
  AND U886 ( .A(n342), .B(n341), .Z(n417) );
  XNOR U887 ( .A(n417), .B(sreg[232]), .Z(n419) );
  NANDN U888 ( .A(n344), .B(n343), .Z(n348) );
  OR U889 ( .A(n346), .B(n345), .Z(n347) );
  AND U890 ( .A(n348), .B(n347), .Z(n413) );
  NANDN U891 ( .A(n350), .B(n349), .Z(n354) );
  NANDN U892 ( .A(n352), .B(n351), .Z(n353) );
  AND U893 ( .A(n354), .B(n353), .Z(n412) );
  NANDN U894 ( .A(n356), .B(n355), .Z(n360) );
  NANDN U895 ( .A(n358), .B(n357), .Z(n359) );
  AND U896 ( .A(n360), .B(n359), .Z(n379) );
  NAND U897 ( .A(n184), .B(n362), .Z(n364) );
  XOR U898 ( .A(b[7]), .B(a[2]), .Z(n393) );
  NAND U899 ( .A(n36592), .B(n393), .Z(n363) );
  AND U900 ( .A(n364), .B(n363), .Z(n383) );
  OR U901 ( .A(n365), .B(n180), .Z(n367) );
  XOR U902 ( .A(b[3]), .B(a[6]), .Z(n408) );
  NAND U903 ( .A(n182), .B(n408), .Z(n366) );
  NAND U904 ( .A(n367), .B(n366), .Z(n382) );
  XNOR U905 ( .A(n383), .B(n382), .Z(n385) );
  NOR U906 ( .A(n369), .B(n368), .Z(n384) );
  XOR U907 ( .A(n385), .B(n384), .Z(n377) );
  NAND U908 ( .A(b[0]), .B(a[8]), .Z(n370) );
  XNOR U909 ( .A(b[1]), .B(n370), .Z(n372) );
  NANDN U910 ( .A(b[0]), .B(a[7]), .Z(n371) );
  NAND U911 ( .A(n372), .B(n371), .Z(n390) );
  XNOR U912 ( .A(b[7]), .B(b[8]), .Z(n2052) );
  IV U913 ( .A(n2052), .Z(n36805) );
  AND U914 ( .A(a[0]), .B(n36805), .Z(n401) );
  NAND U915 ( .A(n183), .B(n373), .Z(n375) );
  XOR U916 ( .A(b[5]), .B(a[4]), .Z(n402) );
  NAND U917 ( .A(n36296), .B(n402), .Z(n374) );
  AND U918 ( .A(n375), .B(n374), .Z(n388) );
  XOR U919 ( .A(n401), .B(n388), .Z(n389) );
  XNOR U920 ( .A(n390), .B(n389), .Z(n376) );
  XNOR U921 ( .A(n377), .B(n376), .Z(n378) );
  XNOR U922 ( .A(n379), .B(n378), .Z(n411) );
  XOR U923 ( .A(n412), .B(n411), .Z(n414) );
  XNOR U924 ( .A(n413), .B(n414), .Z(n418) );
  XOR U925 ( .A(n419), .B(n418), .Z(c[232]) );
  NANDN U926 ( .A(n377), .B(n376), .Z(n381) );
  NANDN U927 ( .A(n379), .B(n378), .Z(n380) );
  AND U928 ( .A(n381), .B(n380), .Z(n427) );
  NANDN U929 ( .A(n383), .B(n382), .Z(n387) );
  NAND U930 ( .A(n385), .B(n384), .Z(n386) );
  AND U931 ( .A(n387), .B(n386), .Z(n466) );
  NANDN U932 ( .A(n388), .B(n401), .Z(n392) );
  OR U933 ( .A(n390), .B(n389), .Z(n391) );
  AND U934 ( .A(n392), .B(n391), .Z(n464) );
  NAND U935 ( .A(n184), .B(n393), .Z(n395) );
  XOR U936 ( .A(b[7]), .B(a[3]), .Z(n448) );
  NAND U937 ( .A(n36592), .B(n448), .Z(n394) );
  AND U938 ( .A(n395), .B(n394), .Z(n458) );
  XOR U939 ( .A(b[9]), .B(b[8]), .Z(n454) );
  XOR U940 ( .A(b[9]), .B(a[0]), .Z(n396) );
  NAND U941 ( .A(n454), .B(n396), .Z(n397) );
  NANDN U942 ( .A(n397), .B(n2052), .Z(n399) );
  XOR U943 ( .A(b[9]), .B(a[1]), .Z(n455) );
  NANDN U944 ( .A(n2052), .B(n455), .Z(n398) );
  NAND U945 ( .A(n399), .B(n398), .Z(n459) );
  XOR U946 ( .A(n458), .B(n459), .Z(n435) );
  NAND U947 ( .A(b[7]), .B(b[8]), .Z(n400) );
  NAND U948 ( .A(b[9]), .B(n400), .Z(n37205) );
  NOR U949 ( .A(n37205), .B(n401), .Z(n434) );
  NAND U950 ( .A(n183), .B(n402), .Z(n404) );
  XOR U951 ( .A(b[5]), .B(a[5]), .Z(n451) );
  NAND U952 ( .A(n36296), .B(n451), .Z(n403) );
  AND U953 ( .A(n404), .B(n403), .Z(n433) );
  XOR U954 ( .A(n434), .B(n433), .Z(n436) );
  XOR U955 ( .A(n435), .B(n436), .Z(n442) );
  NAND U956 ( .A(b[0]), .B(a[9]), .Z(n405) );
  XNOR U957 ( .A(b[1]), .B(n405), .Z(n407) );
  NANDN U958 ( .A(b[0]), .B(a[8]), .Z(n406) );
  NAND U959 ( .A(n407), .B(n406), .Z(n440) );
  NAND U960 ( .A(n181), .B(n408), .Z(n410) );
  XOR U961 ( .A(b[3]), .B(a[7]), .Z(n460) );
  NAND U962 ( .A(n182), .B(n460), .Z(n409) );
  NAND U963 ( .A(n410), .B(n409), .Z(n439) );
  XNOR U964 ( .A(n440), .B(n439), .Z(n441) );
  XOR U965 ( .A(n442), .B(n441), .Z(n463) );
  XNOR U966 ( .A(n464), .B(n463), .Z(n465) );
  XOR U967 ( .A(n466), .B(n465), .Z(n428) );
  XNOR U968 ( .A(n427), .B(n428), .Z(n429) );
  NANDN U969 ( .A(n412), .B(n411), .Z(n416) );
  OR U970 ( .A(n414), .B(n413), .Z(n415) );
  NAND U971 ( .A(n416), .B(n415), .Z(n430) );
  XOR U972 ( .A(n429), .B(n430), .Z(n422) );
  XNOR U973 ( .A(sreg[233]), .B(n422), .Z(n424) );
  NANDN U974 ( .A(n417), .B(sreg[232]), .Z(n421) );
  NAND U975 ( .A(n419), .B(n418), .Z(n420) );
  NAND U976 ( .A(n421), .B(n420), .Z(n423) );
  XOR U977 ( .A(n424), .B(n423), .Z(c[233]) );
  NANDN U978 ( .A(n422), .B(sreg[233]), .Z(n426) );
  NAND U979 ( .A(n424), .B(n423), .Z(n425) );
  AND U980 ( .A(n426), .B(n425), .Z(n469) );
  XNOR U981 ( .A(n469), .B(sreg[234]), .Z(n471) );
  NANDN U982 ( .A(n428), .B(n427), .Z(n432) );
  NANDN U983 ( .A(n430), .B(n429), .Z(n431) );
  AND U984 ( .A(n432), .B(n431), .Z(n477) );
  NANDN U985 ( .A(n434), .B(n433), .Z(n438) );
  NANDN U986 ( .A(n436), .B(n435), .Z(n437) );
  AND U987 ( .A(n438), .B(n437), .Z(n519) );
  NANDN U988 ( .A(n440), .B(n439), .Z(n444) );
  NAND U989 ( .A(n442), .B(n441), .Z(n443) );
  AND U990 ( .A(n444), .B(n443), .Z(n518) );
  XNOR U991 ( .A(n519), .B(n518), .Z(n520) );
  NAND U992 ( .A(b[0]), .B(a[10]), .Z(n445) );
  XNOR U993 ( .A(b[1]), .B(n445), .Z(n447) );
  NANDN U994 ( .A(b[0]), .B(a[9]), .Z(n446) );
  NAND U995 ( .A(n447), .B(n446), .Z(n488) );
  XNOR U996 ( .A(b[9]), .B(b[10]), .Z(n2434) );
  IV U997 ( .A(n2434), .Z(n37097) );
  AND U998 ( .A(a[0]), .B(n37097), .Z(n511) );
  NAND U999 ( .A(n184), .B(n448), .Z(n450) );
  XOR U1000 ( .A(b[7]), .B(a[4]), .Z(n512) );
  NAND U1001 ( .A(n36592), .B(n512), .Z(n449) );
  AND U1002 ( .A(n450), .B(n449), .Z(n486) );
  XOR U1003 ( .A(n511), .B(n486), .Z(n487) );
  XOR U1004 ( .A(n488), .B(n487), .Z(n483) );
  NAND U1005 ( .A(n183), .B(n451), .Z(n453) );
  XOR U1006 ( .A(b[5]), .B(a[6]), .Z(n507) );
  NAND U1007 ( .A(n36296), .B(n507), .Z(n452) );
  AND U1008 ( .A(n453), .B(n452), .Z(n492) );
  NAND U1009 ( .A(n185), .B(n455), .Z(n457) );
  XOR U1010 ( .A(b[9]), .B(a[2]), .Z(n501) );
  NAND U1011 ( .A(n36805), .B(n501), .Z(n456) );
  NAND U1012 ( .A(n457), .B(n456), .Z(n491) );
  XNOR U1013 ( .A(n492), .B(n491), .Z(n494) );
  ANDN U1014 ( .B(n459), .A(n458), .Z(n493) );
  XOR U1015 ( .A(n494), .B(n493), .Z(n481) );
  NANDN U1016 ( .A(n180), .B(n460), .Z(n462) );
  XNOR U1017 ( .A(b[3]), .B(a[8]), .Z(n515) );
  OR U1018 ( .A(n515), .B(n172), .Z(n461) );
  AND U1019 ( .A(n462), .B(n461), .Z(n480) );
  XNOR U1020 ( .A(n481), .B(n480), .Z(n482) );
  XOR U1021 ( .A(n483), .B(n482), .Z(n521) );
  XNOR U1022 ( .A(n520), .B(n521), .Z(n474) );
  NANDN U1023 ( .A(n464), .B(n463), .Z(n468) );
  NANDN U1024 ( .A(n466), .B(n465), .Z(n467) );
  NAND U1025 ( .A(n468), .B(n467), .Z(n475) );
  XNOR U1026 ( .A(n474), .B(n475), .Z(n476) );
  XNOR U1027 ( .A(n477), .B(n476), .Z(n470) );
  XOR U1028 ( .A(n471), .B(n470), .Z(c[234]) );
  NANDN U1029 ( .A(n469), .B(sreg[234]), .Z(n473) );
  NAND U1030 ( .A(n471), .B(n470), .Z(n472) );
  AND U1031 ( .A(n473), .B(n472), .Z(n526) );
  NANDN U1032 ( .A(n475), .B(n474), .Z(n479) );
  NAND U1033 ( .A(n477), .B(n476), .Z(n478) );
  AND U1034 ( .A(n479), .B(n478), .Z(n532) );
  NANDN U1035 ( .A(n481), .B(n480), .Z(n485) );
  NANDN U1036 ( .A(n483), .B(n482), .Z(n484) );
  AND U1037 ( .A(n485), .B(n484), .Z(n578) );
  NANDN U1038 ( .A(n486), .B(n511), .Z(n490) );
  OR U1039 ( .A(n488), .B(n487), .Z(n489) );
  AND U1040 ( .A(n490), .B(n489), .Z(n576) );
  NANDN U1041 ( .A(n492), .B(n491), .Z(n496) );
  NAND U1042 ( .A(n494), .B(n493), .Z(n495) );
  AND U1043 ( .A(n496), .B(n495), .Z(n538) );
  XOR U1044 ( .A(b[11]), .B(b[10]), .Z(n559) );
  XOR U1045 ( .A(b[11]), .B(a[0]), .Z(n497) );
  NAND U1046 ( .A(n559), .B(n497), .Z(n498) );
  NANDN U1047 ( .A(n498), .B(n2434), .Z(n500) );
  XOR U1048 ( .A(b[11]), .B(a[1]), .Z(n560) );
  NANDN U1049 ( .A(n2434), .B(n560), .Z(n499) );
  AND U1050 ( .A(n500), .B(n499), .Z(n567) );
  NAND U1051 ( .A(n185), .B(n501), .Z(n503) );
  XOR U1052 ( .A(b[9]), .B(a[3]), .Z(n550) );
  NAND U1053 ( .A(n36805), .B(n550), .Z(n502) );
  AND U1054 ( .A(n503), .B(n502), .Z(n566) );
  XOR U1055 ( .A(n567), .B(n566), .Z(n555) );
  NAND U1056 ( .A(b[0]), .B(a[11]), .Z(n504) );
  XNOR U1057 ( .A(b[1]), .B(n504), .Z(n506) );
  NANDN U1058 ( .A(b[0]), .B(a[10]), .Z(n505) );
  NAND U1059 ( .A(n506), .B(n505), .Z(n553) );
  NANDN U1060 ( .A(n173), .B(n507), .Z(n509) );
  XNOR U1061 ( .A(b[5]), .B(a[7]), .Z(n563) );
  OR U1062 ( .A(n563), .B(n622), .Z(n508) );
  NAND U1063 ( .A(n509), .B(n508), .Z(n554) );
  XOR U1064 ( .A(n553), .B(n554), .Z(n556) );
  XOR U1065 ( .A(n555), .B(n556), .Z(n536) );
  NAND U1066 ( .A(b[9]), .B(b[10]), .Z(n510) );
  AND U1067 ( .A(b[11]), .B(n510), .Z(n37301) );
  IV U1068 ( .A(n37301), .Z(n37390) );
  NOR U1069 ( .A(n37390), .B(n511), .Z(n542) );
  NANDN U1070 ( .A(n175), .B(n512), .Z(n514) );
  XNOR U1071 ( .A(b[7]), .B(a[5]), .Z(n571) );
  OR U1072 ( .A(n571), .B(n572), .Z(n513) );
  NAND U1073 ( .A(n514), .B(n513), .Z(n541) );
  XOR U1074 ( .A(n542), .B(n541), .Z(n544) );
  OR U1075 ( .A(n515), .B(n180), .Z(n517) );
  XNOR U1076 ( .A(b[3]), .B(a[9]), .Z(n568) );
  OR U1077 ( .A(n568), .B(n172), .Z(n516) );
  NAND U1078 ( .A(n517), .B(n516), .Z(n543) );
  XOR U1079 ( .A(n544), .B(n543), .Z(n535) );
  XNOR U1080 ( .A(n536), .B(n535), .Z(n537) );
  XNOR U1081 ( .A(n538), .B(n537), .Z(n575) );
  XNOR U1082 ( .A(n576), .B(n575), .Z(n577) );
  XOR U1083 ( .A(n578), .B(n577), .Z(n530) );
  NANDN U1084 ( .A(n519), .B(n518), .Z(n523) );
  NANDN U1085 ( .A(n521), .B(n520), .Z(n522) );
  NAND U1086 ( .A(n523), .B(n522), .Z(n529) );
  XNOR U1087 ( .A(n530), .B(n529), .Z(n531) );
  XNOR U1088 ( .A(n532), .B(n531), .Z(n524) );
  XNOR U1089 ( .A(sreg[235]), .B(n524), .Z(n525) );
  XNOR U1090 ( .A(n526), .B(n525), .Z(c[235]) );
  NANDN U1091 ( .A(sreg[235]), .B(n524), .Z(n528) );
  NAND U1092 ( .A(n526), .B(n525), .Z(n527) );
  NAND U1093 ( .A(n528), .B(n527), .Z(n643) );
  XNOR U1094 ( .A(sreg[236]), .B(n643), .Z(n645) );
  NANDN U1095 ( .A(n530), .B(n529), .Z(n534) );
  NANDN U1096 ( .A(n532), .B(n531), .Z(n533) );
  AND U1097 ( .A(n534), .B(n533), .Z(n583) );
  NANDN U1098 ( .A(n536), .B(n535), .Z(n540) );
  NANDN U1099 ( .A(n538), .B(n537), .Z(n539) );
  AND U1100 ( .A(n540), .B(n539), .Z(n638) );
  NAND U1101 ( .A(n542), .B(n541), .Z(n546) );
  NAND U1102 ( .A(n544), .B(n543), .Z(n545) );
  NAND U1103 ( .A(n546), .B(n545), .Z(n637) );
  XNOR U1104 ( .A(n638), .B(n637), .Z(n640) );
  AND U1105 ( .A(b[0]), .B(a[12]), .Z(n547) );
  XOR U1106 ( .A(b[1]), .B(n547), .Z(n549) );
  NANDN U1107 ( .A(b[0]), .B(a[11]), .Z(n548) );
  AND U1108 ( .A(n549), .B(n548), .Z(n627) );
  XNOR U1109 ( .A(b[11]), .B(b[12]), .Z(n1681) );
  IV U1110 ( .A(n1681), .Z(n37295) );
  AND U1111 ( .A(a[0]), .B(n37295), .Z(n625) );
  NAND U1112 ( .A(n185), .B(n550), .Z(n552) );
  XOR U1113 ( .A(b[9]), .B(a[4]), .Z(n618) );
  NAND U1114 ( .A(n36805), .B(n618), .Z(n551) );
  AND U1115 ( .A(n552), .B(n551), .Z(n626) );
  XOR U1116 ( .A(n625), .B(n626), .Z(n628) );
  XNOR U1117 ( .A(n627), .B(n628), .Z(n587) );
  NANDN U1118 ( .A(n554), .B(n553), .Z(n558) );
  OR U1119 ( .A(n556), .B(n555), .Z(n557) );
  NAND U1120 ( .A(n558), .B(n557), .Z(n588) );
  XNOR U1121 ( .A(n587), .B(n588), .Z(n589) );
  NAND U1122 ( .A(n186), .B(n560), .Z(n562) );
  XOR U1123 ( .A(b[11]), .B(a[2]), .Z(n605) );
  NAND U1124 ( .A(n37097), .B(n605), .Z(n561) );
  AND U1125 ( .A(n562), .B(n561), .Z(n596) );
  OR U1126 ( .A(n563), .B(n173), .Z(n565) );
  XOR U1127 ( .A(b[5]), .B(a[8]), .Z(n621) );
  NAND U1128 ( .A(n36296), .B(n621), .Z(n564) );
  AND U1129 ( .A(n565), .B(n564), .Z(n594) );
  NOR U1130 ( .A(n567), .B(n566), .Z(n633) );
  OR U1131 ( .A(n568), .B(n180), .Z(n570) );
  XNOR U1132 ( .A(b[3]), .B(a[10]), .Z(n615) );
  OR U1133 ( .A(n615), .B(n172), .Z(n569) );
  AND U1134 ( .A(n570), .B(n569), .Z(n631) );
  OR U1135 ( .A(n571), .B(n175), .Z(n574) );
  XNOR U1136 ( .A(b[7]), .B(a[6]), .Z(n602) );
  OR U1137 ( .A(n602), .B(n572), .Z(n573) );
  NAND U1138 ( .A(n574), .B(n573), .Z(n632) );
  XOR U1139 ( .A(n631), .B(n632), .Z(n634) );
  XNOR U1140 ( .A(n633), .B(n634), .Z(n593) );
  XNOR U1141 ( .A(n594), .B(n593), .Z(n595) );
  XOR U1142 ( .A(n596), .B(n595), .Z(n590) );
  XNOR U1143 ( .A(n589), .B(n590), .Z(n639) );
  XOR U1144 ( .A(n640), .B(n639), .Z(n582) );
  NANDN U1145 ( .A(n576), .B(n575), .Z(n580) );
  NAND U1146 ( .A(n578), .B(n577), .Z(n579) );
  AND U1147 ( .A(n580), .B(n579), .Z(n581) );
  XOR U1148 ( .A(n582), .B(n581), .Z(n584) );
  XNOR U1149 ( .A(n583), .B(n584), .Z(n644) );
  XOR U1150 ( .A(n645), .B(n644), .Z(c[236]) );
  NANDN U1151 ( .A(n582), .B(n581), .Z(n586) );
  OR U1152 ( .A(n584), .B(n583), .Z(n585) );
  AND U1153 ( .A(n586), .B(n585), .Z(n655) );
  NANDN U1154 ( .A(n588), .B(n587), .Z(n592) );
  NANDN U1155 ( .A(n590), .B(n589), .Z(n591) );
  AND U1156 ( .A(n592), .B(n591), .Z(n709) );
  NANDN U1157 ( .A(n594), .B(n593), .Z(n598) );
  NANDN U1158 ( .A(n596), .B(n595), .Z(n597) );
  AND U1159 ( .A(n598), .B(n597), .Z(n708) );
  NAND U1160 ( .A(b[0]), .B(a[13]), .Z(n599) );
  XNOR U1161 ( .A(b[1]), .B(n599), .Z(n601) );
  NANDN U1162 ( .A(b[0]), .B(a[12]), .Z(n600) );
  NAND U1163 ( .A(n601), .B(n600), .Z(n693) );
  OR U1164 ( .A(n602), .B(n175), .Z(n604) );
  XOR U1165 ( .A(b[7]), .B(a[7]), .Z(n686) );
  NAND U1166 ( .A(n36592), .B(n686), .Z(n603) );
  NAND U1167 ( .A(n604), .B(n603), .Z(n692) );
  XNOR U1168 ( .A(n693), .B(n692), .Z(n695) );
  NAND U1169 ( .A(n186), .B(n605), .Z(n607) );
  XOR U1170 ( .A(b[11]), .B(a[3]), .Z(n680) );
  NAND U1171 ( .A(n37097), .B(n680), .Z(n606) );
  AND U1172 ( .A(n607), .B(n606), .Z(n706) );
  XOR U1173 ( .A(b[13]), .B(a[1]), .Z(n699) );
  NAND U1174 ( .A(n37295), .B(n699), .Z(n614) );
  ANDN U1175 ( .B(b[12]), .A(b[13]), .Z(n608) );
  NAND U1176 ( .A(n608), .B(a[0]), .Z(n611) );
  NAND U1177 ( .A(b[11]), .B(b[12]), .Z(n609) );
  AND U1178 ( .A(b[13]), .B(n609), .Z(n37507) );
  NANDN U1179 ( .A(a[0]), .B(n37507), .Z(n610) );
  NAND U1180 ( .A(n611), .B(n610), .Z(n612) );
  NANDN U1181 ( .A(n37295), .B(n612), .Z(n613) );
  NAND U1182 ( .A(n614), .B(n613), .Z(n705) );
  XNOR U1183 ( .A(n706), .B(n705), .Z(n694) );
  XOR U1184 ( .A(n695), .B(n694), .Z(n667) );
  OR U1185 ( .A(n615), .B(n180), .Z(n617) );
  XOR U1186 ( .A(b[3]), .B(a[11]), .Z(n689) );
  NAND U1187 ( .A(n182), .B(n689), .Z(n616) );
  AND U1188 ( .A(n617), .B(n616), .Z(n672) );
  NAND U1189 ( .A(n185), .B(n618), .Z(n620) );
  XOR U1190 ( .A(b[9]), .B(a[5]), .Z(n702) );
  NAND U1191 ( .A(n36805), .B(n702), .Z(n619) );
  NAND U1192 ( .A(n620), .B(n619), .Z(n671) );
  XNOR U1193 ( .A(n672), .B(n671), .Z(n674) );
  IV U1194 ( .A(n37507), .Z(n37554) );
  NOR U1195 ( .A(n37554), .B(n625), .Z(n673) );
  XOR U1196 ( .A(n674), .B(n673), .Z(n666) );
  NANDN U1197 ( .A(n173), .B(n621), .Z(n624) );
  XNOR U1198 ( .A(b[5]), .B(a[9]), .Z(n683) );
  OR U1199 ( .A(n683), .B(n622), .Z(n623) );
  AND U1200 ( .A(n624), .B(n623), .Z(n665) );
  XOR U1201 ( .A(n666), .B(n665), .Z(n668) );
  XOR U1202 ( .A(n667), .B(n668), .Z(n662) );
  NANDN U1203 ( .A(n626), .B(n625), .Z(n630) );
  NANDN U1204 ( .A(n628), .B(n627), .Z(n629) );
  AND U1205 ( .A(n630), .B(n629), .Z(n660) );
  NANDN U1206 ( .A(n632), .B(n631), .Z(n636) );
  OR U1207 ( .A(n634), .B(n633), .Z(n635) );
  AND U1208 ( .A(n636), .B(n635), .Z(n659) );
  XNOR U1209 ( .A(n660), .B(n659), .Z(n661) );
  XNOR U1210 ( .A(n662), .B(n661), .Z(n707) );
  XOR U1211 ( .A(n708), .B(n707), .Z(n710) );
  XOR U1212 ( .A(n709), .B(n710), .Z(n654) );
  NANDN U1213 ( .A(n638), .B(n637), .Z(n642) );
  NAND U1214 ( .A(n640), .B(n639), .Z(n641) );
  AND U1215 ( .A(n642), .B(n641), .Z(n653) );
  XOR U1216 ( .A(n654), .B(n653), .Z(n656) );
  XOR U1217 ( .A(n655), .B(n656), .Z(n648) );
  XNOR U1218 ( .A(n648), .B(sreg[237]), .Z(n650) );
  NANDN U1219 ( .A(n643), .B(sreg[236]), .Z(n647) );
  NAND U1220 ( .A(n645), .B(n644), .Z(n646) );
  NAND U1221 ( .A(n647), .B(n646), .Z(n649) );
  XOR U1222 ( .A(n650), .B(n649), .Z(c[237]) );
  NANDN U1223 ( .A(n648), .B(sreg[237]), .Z(n652) );
  NAND U1224 ( .A(n650), .B(n649), .Z(n651) );
  AND U1225 ( .A(n652), .B(n651), .Z(n780) );
  XNOR U1226 ( .A(sreg[238]), .B(n780), .Z(n782) );
  NANDN U1227 ( .A(n654), .B(n653), .Z(n658) );
  OR U1228 ( .A(n656), .B(n655), .Z(n657) );
  AND U1229 ( .A(n658), .B(n657), .Z(n716) );
  NANDN U1230 ( .A(n660), .B(n659), .Z(n664) );
  NANDN U1231 ( .A(n662), .B(n661), .Z(n663) );
  AND U1232 ( .A(n664), .B(n663), .Z(n776) );
  NANDN U1233 ( .A(n666), .B(n665), .Z(n670) );
  OR U1234 ( .A(n668), .B(n667), .Z(n669) );
  AND U1235 ( .A(n670), .B(n669), .Z(n774) );
  NANDN U1236 ( .A(n672), .B(n671), .Z(n676) );
  NAND U1237 ( .A(n674), .B(n673), .Z(n675) );
  AND U1238 ( .A(n676), .B(n675), .Z(n761) );
  NAND U1239 ( .A(b[0]), .B(a[14]), .Z(n677) );
  XNOR U1240 ( .A(b[1]), .B(n677), .Z(n679) );
  NANDN U1241 ( .A(b[0]), .B(a[13]), .Z(n678) );
  NAND U1242 ( .A(n679), .B(n678), .Z(n767) );
  XNOR U1243 ( .A(b[13]), .B(b[14]), .Z(n37509) );
  IV U1244 ( .A(n37509), .Z(n37382) );
  AND U1245 ( .A(a[0]), .B(n37382), .Z(n764) );
  NAND U1246 ( .A(n186), .B(n680), .Z(n682) );
  XOR U1247 ( .A(b[11]), .B(a[4]), .Z(n734) );
  NAND U1248 ( .A(n37097), .B(n734), .Z(n681) );
  AND U1249 ( .A(n682), .B(n681), .Z(n765) );
  XNOR U1250 ( .A(n764), .B(n765), .Z(n766) );
  XNOR U1251 ( .A(n767), .B(n766), .Z(n758) );
  OR U1252 ( .A(n683), .B(n173), .Z(n685) );
  XOR U1253 ( .A(b[5]), .B(a[10]), .Z(n728) );
  NAND U1254 ( .A(n36296), .B(n728), .Z(n684) );
  AND U1255 ( .A(n685), .B(n684), .Z(n755) );
  NAND U1256 ( .A(n184), .B(n686), .Z(n688) );
  XOR U1257 ( .A(b[7]), .B(a[8]), .Z(n725) );
  NAND U1258 ( .A(n36592), .B(n725), .Z(n687) );
  AND U1259 ( .A(n688), .B(n687), .Z(n753) );
  NAND U1260 ( .A(n181), .B(n689), .Z(n691) );
  XOR U1261 ( .A(b[3]), .B(a[12]), .Z(n731) );
  NAND U1262 ( .A(n182), .B(n731), .Z(n690) );
  NAND U1263 ( .A(n691), .B(n690), .Z(n752) );
  XNOR U1264 ( .A(n753), .B(n752), .Z(n754) );
  XOR U1265 ( .A(n755), .B(n754), .Z(n759) );
  XNOR U1266 ( .A(n758), .B(n759), .Z(n760) );
  XNOR U1267 ( .A(n761), .B(n760), .Z(n721) );
  NANDN U1268 ( .A(n693), .B(n692), .Z(n697) );
  NAND U1269 ( .A(n695), .B(n694), .Z(n696) );
  AND U1270 ( .A(n697), .B(n696), .Z(n720) );
  XOR U1271 ( .A(b[12]), .B(b[13]), .Z(n698) );
  NAND U1272 ( .A(n187), .B(n699), .Z(n701) );
  XOR U1273 ( .A(b[13]), .B(a[2]), .Z(n749) );
  NAND U1274 ( .A(n37295), .B(n749), .Z(n700) );
  AND U1275 ( .A(n701), .B(n700), .Z(n771) );
  NAND U1276 ( .A(n185), .B(n702), .Z(n704) );
  XOR U1277 ( .A(b[9]), .B(a[6]), .Z(n741) );
  NAND U1278 ( .A(n36805), .B(n741), .Z(n703) );
  NAND U1279 ( .A(n704), .B(n703), .Z(n770) );
  XNOR U1280 ( .A(n771), .B(n770), .Z(n773) );
  NANDN U1281 ( .A(n706), .B(n705), .Z(n772) );
  XNOR U1282 ( .A(n773), .B(n772), .Z(n719) );
  XOR U1283 ( .A(n720), .B(n719), .Z(n722) );
  XOR U1284 ( .A(n721), .B(n722), .Z(n775) );
  XOR U1285 ( .A(n774), .B(n775), .Z(n777) );
  XOR U1286 ( .A(n776), .B(n777), .Z(n714) );
  NANDN U1287 ( .A(n708), .B(n707), .Z(n712) );
  OR U1288 ( .A(n710), .B(n709), .Z(n711) );
  AND U1289 ( .A(n712), .B(n711), .Z(n713) );
  XNOR U1290 ( .A(n714), .B(n713), .Z(n715) );
  XNOR U1291 ( .A(n716), .B(n715), .Z(n781) );
  XNOR U1292 ( .A(n782), .B(n781), .Z(c[238]) );
  NANDN U1293 ( .A(n714), .B(n713), .Z(n718) );
  NANDN U1294 ( .A(n716), .B(n715), .Z(n717) );
  AND U1295 ( .A(n718), .B(n717), .Z(n792) );
  NANDN U1296 ( .A(n720), .B(n719), .Z(n724) );
  NANDN U1297 ( .A(n722), .B(n721), .Z(n723) );
  AND U1298 ( .A(n724), .B(n723), .Z(n854) );
  NAND U1299 ( .A(n184), .B(n725), .Z(n727) );
  XOR U1300 ( .A(b[7]), .B(a[9]), .Z(n834) );
  NAND U1301 ( .A(n36592), .B(n834), .Z(n726) );
  AND U1302 ( .A(n727), .B(n726), .Z(n821) );
  NAND U1303 ( .A(n183), .B(n728), .Z(n730) );
  XOR U1304 ( .A(b[5]), .B(a[11]), .Z(n844) );
  NAND U1305 ( .A(n36296), .B(n844), .Z(n729) );
  AND U1306 ( .A(n730), .B(n729), .Z(n805) );
  NAND U1307 ( .A(n181), .B(n731), .Z(n733) );
  XOR U1308 ( .A(b[3]), .B(a[13]), .Z(n828) );
  NAND U1309 ( .A(n182), .B(n828), .Z(n732) );
  AND U1310 ( .A(n733), .B(n732), .Z(n803) );
  NAND U1311 ( .A(n186), .B(n734), .Z(n736) );
  XOR U1312 ( .A(b[11]), .B(a[5]), .Z(n837) );
  NAND U1313 ( .A(n37097), .B(n837), .Z(n735) );
  NAND U1314 ( .A(n736), .B(n735), .Z(n802) );
  XNOR U1315 ( .A(n803), .B(n802), .Z(n804) );
  XNOR U1316 ( .A(n805), .B(n804), .Z(n820) );
  XNOR U1317 ( .A(n821), .B(n820), .Z(n823) );
  NAND U1318 ( .A(b[13]), .B(b[14]), .Z(n737) );
  AND U1319 ( .A(b[15]), .B(n737), .Z(n37685) );
  IV U1320 ( .A(n37685), .Z(n37770) );
  NOR U1321 ( .A(n37770), .B(n764), .Z(n822) );
  XOR U1322 ( .A(n823), .B(n822), .Z(n849) );
  NAND U1323 ( .A(b[0]), .B(a[15]), .Z(n738) );
  XNOR U1324 ( .A(b[1]), .B(n738), .Z(n740) );
  NANDN U1325 ( .A(b[0]), .B(a[14]), .Z(n739) );
  NAND U1326 ( .A(n740), .B(n739), .Z(n815) );
  NAND U1327 ( .A(n185), .B(n741), .Z(n743) );
  XOR U1328 ( .A(b[9]), .B(a[7]), .Z(n831) );
  NAND U1329 ( .A(n36805), .B(n831), .Z(n742) );
  NAND U1330 ( .A(n743), .B(n742), .Z(n814) );
  XNOR U1331 ( .A(n815), .B(n814), .Z(n817) );
  XOR U1332 ( .A(b[15]), .B(a[0]), .Z(n746) );
  XOR U1333 ( .A(b[15]), .B(b[13]), .Z(n744) );
  XOR U1334 ( .A(b[15]), .B(b[14]), .Z(n840) );
  AND U1335 ( .A(n744), .B(n840), .Z(n745) );
  NAND U1336 ( .A(n746), .B(n745), .Z(n748) );
  XOR U1337 ( .A(b[15]), .B(a[1]), .Z(n841) );
  NANDN U1338 ( .A(n37509), .B(n841), .Z(n747) );
  AND U1339 ( .A(n748), .B(n747), .Z(n826) );
  NAND U1340 ( .A(n187), .B(n749), .Z(n751) );
  XOR U1341 ( .A(b[13]), .B(a[3]), .Z(n811) );
  NAND U1342 ( .A(n37295), .B(n811), .Z(n750) );
  NAND U1343 ( .A(n751), .B(n750), .Z(n827) );
  XNOR U1344 ( .A(n826), .B(n827), .Z(n816) );
  XOR U1345 ( .A(n817), .B(n816), .Z(n848) );
  NANDN U1346 ( .A(n753), .B(n752), .Z(n757) );
  NANDN U1347 ( .A(n755), .B(n754), .Z(n756) );
  AND U1348 ( .A(n757), .B(n756), .Z(n847) );
  XOR U1349 ( .A(n848), .B(n847), .Z(n850) );
  XNOR U1350 ( .A(n849), .B(n850), .Z(n853) );
  XNOR U1351 ( .A(n854), .B(n853), .Z(n856) );
  NANDN U1352 ( .A(n759), .B(n758), .Z(n763) );
  NANDN U1353 ( .A(n761), .B(n760), .Z(n762) );
  AND U1354 ( .A(n763), .B(n762), .Z(n799) );
  NANDN U1355 ( .A(n765), .B(n764), .Z(n769) );
  NANDN U1356 ( .A(n767), .B(n766), .Z(n768) );
  AND U1357 ( .A(n769), .B(n768), .Z(n797) );
  XNOR U1358 ( .A(n797), .B(n796), .Z(n798) );
  XNOR U1359 ( .A(n799), .B(n798), .Z(n855) );
  XOR U1360 ( .A(n856), .B(n855), .Z(n791) );
  NANDN U1361 ( .A(n775), .B(n774), .Z(n779) );
  OR U1362 ( .A(n777), .B(n776), .Z(n778) );
  AND U1363 ( .A(n779), .B(n778), .Z(n790) );
  XOR U1364 ( .A(n791), .B(n790), .Z(n793) );
  XOR U1365 ( .A(n792), .B(n793), .Z(n785) );
  XNOR U1366 ( .A(n785), .B(sreg[239]), .Z(n787) );
  NANDN U1367 ( .A(sreg[238]), .B(n780), .Z(n784) );
  NAND U1368 ( .A(n782), .B(n781), .Z(n783) );
  AND U1369 ( .A(n784), .B(n783), .Z(n786) );
  XOR U1370 ( .A(n787), .B(n786), .Z(c[239]) );
  NANDN U1371 ( .A(n785), .B(sreg[239]), .Z(n789) );
  NAND U1372 ( .A(n787), .B(n786), .Z(n788) );
  AND U1373 ( .A(n789), .B(n788), .Z(n859) );
  XNOR U1374 ( .A(n859), .B(sreg[240]), .Z(n861) );
  NANDN U1375 ( .A(n791), .B(n790), .Z(n795) );
  OR U1376 ( .A(n793), .B(n792), .Z(n794) );
  AND U1377 ( .A(n795), .B(n794), .Z(n866) );
  NANDN U1378 ( .A(n797), .B(n796), .Z(n801) );
  NANDN U1379 ( .A(n799), .B(n798), .Z(n800) );
  AND U1380 ( .A(n801), .B(n800), .Z(n939) );
  NANDN U1381 ( .A(n803), .B(n802), .Z(n807) );
  NANDN U1382 ( .A(n805), .B(n804), .Z(n806) );
  AND U1383 ( .A(n807), .B(n806), .Z(n934) );
  NAND U1384 ( .A(b[0]), .B(a[16]), .Z(n808) );
  XNOR U1385 ( .A(b[1]), .B(n808), .Z(n810) );
  NANDN U1386 ( .A(b[0]), .B(a[15]), .Z(n809) );
  NAND U1387 ( .A(n810), .B(n809), .Z(n872) );
  XNOR U1388 ( .A(b[15]), .B(b[16]), .Z(n36922) );
  IV U1389 ( .A(n36922), .Z(n37652) );
  AND U1390 ( .A(a[0]), .B(n37652), .Z(n885) );
  NAND U1391 ( .A(n187), .B(n811), .Z(n813) );
  XOR U1392 ( .A(b[13]), .B(a[4]), .Z(n913) );
  NAND U1393 ( .A(n37295), .B(n913), .Z(n812) );
  AND U1394 ( .A(n813), .B(n812), .Z(n870) );
  XOR U1395 ( .A(n885), .B(n870), .Z(n871) );
  XOR U1396 ( .A(n872), .B(n871), .Z(n932) );
  NANDN U1397 ( .A(n815), .B(n814), .Z(n819) );
  NAND U1398 ( .A(n817), .B(n816), .Z(n818) );
  AND U1399 ( .A(n819), .B(n818), .Z(n931) );
  XNOR U1400 ( .A(n932), .B(n931), .Z(n933) );
  XOR U1401 ( .A(n934), .B(n933), .Z(n928) );
  NANDN U1402 ( .A(n821), .B(n820), .Z(n825) );
  NAND U1403 ( .A(n823), .B(n822), .Z(n824) );
  AND U1404 ( .A(n825), .B(n824), .Z(n926) );
  ANDN U1405 ( .B(n827), .A(n826), .Z(n906) );
  NANDN U1406 ( .A(n180), .B(n828), .Z(n830) );
  XNOR U1407 ( .A(b[3]), .B(a[14]), .Z(n895) );
  OR U1408 ( .A(n895), .B(n172), .Z(n829) );
  AND U1409 ( .A(n830), .B(n829), .Z(n904) );
  NANDN U1410 ( .A(n179), .B(n831), .Z(n833) );
  XNOR U1411 ( .A(b[9]), .B(a[8]), .Z(n886) );
  OR U1412 ( .A(n886), .B(n2052), .Z(n832) );
  NAND U1413 ( .A(n833), .B(n832), .Z(n905) );
  XOR U1414 ( .A(n904), .B(n905), .Z(n907) );
  XOR U1415 ( .A(n906), .B(n907), .Z(n901) );
  NAND U1416 ( .A(n184), .B(n834), .Z(n836) );
  XOR U1417 ( .A(b[7]), .B(a[10]), .Z(n916) );
  NAND U1418 ( .A(n36592), .B(n916), .Z(n835) );
  AND U1419 ( .A(n836), .B(n835), .Z(n899) );
  NAND U1420 ( .A(n186), .B(n837), .Z(n839) );
  XOR U1421 ( .A(b[11]), .B(a[6]), .Z(n910) );
  NAND U1422 ( .A(n37097), .B(n910), .Z(n838) );
  AND U1423 ( .A(n839), .B(n838), .Z(n922) );
  NAND U1424 ( .A(n188), .B(n841), .Z(n843) );
  XOR U1425 ( .A(b[15]), .B(a[2]), .Z(n875) );
  NAND U1426 ( .A(n37382), .B(n875), .Z(n842) );
  AND U1427 ( .A(n843), .B(n842), .Z(n920) );
  NAND U1428 ( .A(n183), .B(n844), .Z(n846) );
  XOR U1429 ( .A(b[5]), .B(a[12]), .Z(n892) );
  NAND U1430 ( .A(n36296), .B(n892), .Z(n845) );
  NAND U1431 ( .A(n846), .B(n845), .Z(n919) );
  XNOR U1432 ( .A(n920), .B(n919), .Z(n921) );
  XNOR U1433 ( .A(n922), .B(n921), .Z(n898) );
  XNOR U1434 ( .A(n899), .B(n898), .Z(n900) );
  XNOR U1435 ( .A(n901), .B(n900), .Z(n925) );
  XNOR U1436 ( .A(n926), .B(n925), .Z(n927) );
  XNOR U1437 ( .A(n928), .B(n927), .Z(n937) );
  NANDN U1438 ( .A(n848), .B(n847), .Z(n852) );
  OR U1439 ( .A(n850), .B(n849), .Z(n851) );
  NAND U1440 ( .A(n852), .B(n851), .Z(n938) );
  XOR U1441 ( .A(n937), .B(n938), .Z(n940) );
  XOR U1442 ( .A(n939), .B(n940), .Z(n865) );
  NANDN U1443 ( .A(n854), .B(n853), .Z(n858) );
  NAND U1444 ( .A(n856), .B(n855), .Z(n857) );
  AND U1445 ( .A(n858), .B(n857), .Z(n864) );
  XOR U1446 ( .A(n865), .B(n864), .Z(n867) );
  XNOR U1447 ( .A(n866), .B(n867), .Z(n860) );
  XOR U1448 ( .A(n861), .B(n860), .Z(c[240]) );
  NANDN U1449 ( .A(n859), .B(sreg[240]), .Z(n863) );
  NAND U1450 ( .A(n861), .B(n860), .Z(n862) );
  AND U1451 ( .A(n863), .B(n862), .Z(n945) );
  NANDN U1452 ( .A(n865), .B(n864), .Z(n869) );
  OR U1453 ( .A(n867), .B(n866), .Z(n868) );
  AND U1454 ( .A(n869), .B(n868), .Z(n951) );
  NANDN U1455 ( .A(n870), .B(n885), .Z(n874) );
  OR U1456 ( .A(n872), .B(n871), .Z(n873) );
  AND U1457 ( .A(n874), .B(n873), .Z(n968) );
  NAND U1458 ( .A(n188), .B(n875), .Z(n877) );
  XOR U1459 ( .A(b[15]), .B(a[3]), .Z(n990) );
  NAND U1460 ( .A(n37382), .B(n990), .Z(n876) );
  AND U1461 ( .A(n877), .B(n876), .Z(n978) );
  XOR U1462 ( .A(b[17]), .B(a[1]), .Z(n984) );
  NAND U1463 ( .A(n37652), .B(n984), .Z(n884) );
  ANDN U1464 ( .B(b[16]), .A(b[17]), .Z(n878) );
  NAND U1465 ( .A(n878), .B(a[0]), .Z(n881) );
  NAND U1466 ( .A(b[15]), .B(b[16]), .Z(n879) );
  NAND U1467 ( .A(b[17]), .B(n879), .Z(n37940) );
  OR U1468 ( .A(a[0]), .B(n37940), .Z(n880) );
  NAND U1469 ( .A(n881), .B(n880), .Z(n882) );
  NANDN U1470 ( .A(n37652), .B(n882), .Z(n883) );
  AND U1471 ( .A(n884), .B(n883), .Z(n979) );
  XOR U1472 ( .A(n978), .B(n979), .Z(n995) );
  NOR U1473 ( .A(n37940), .B(n885), .Z(n994) );
  OR U1474 ( .A(n886), .B(n179), .Z(n888) );
  XNOR U1475 ( .A(b[9]), .B(a[9]), .Z(n1011) );
  OR U1476 ( .A(n1011), .B(n2052), .Z(n887) );
  AND U1477 ( .A(n888), .B(n887), .Z(n993) );
  XOR U1478 ( .A(n994), .B(n993), .Z(n996) );
  XOR U1479 ( .A(n995), .B(n996), .Z(n967) );
  NAND U1480 ( .A(b[0]), .B(a[17]), .Z(n889) );
  XNOR U1481 ( .A(b[1]), .B(n889), .Z(n891) );
  NANDN U1482 ( .A(b[0]), .B(a[16]), .Z(n890) );
  NAND U1483 ( .A(n891), .B(n890), .Z(n973) );
  NAND U1484 ( .A(n183), .B(n892), .Z(n894) );
  XOR U1485 ( .A(b[5]), .B(a[13]), .Z(n1005) );
  NAND U1486 ( .A(n36296), .B(n1005), .Z(n893) );
  NAND U1487 ( .A(n894), .B(n893), .Z(n972) );
  XNOR U1488 ( .A(n973), .B(n972), .Z(n975) );
  OR U1489 ( .A(n895), .B(n180), .Z(n897) );
  XNOR U1490 ( .A(b[3]), .B(a[15]), .Z(n1017) );
  OR U1491 ( .A(n1017), .B(n172), .Z(n896) );
  NAND U1492 ( .A(n897), .B(n896), .Z(n974) );
  XOR U1493 ( .A(n975), .B(n974), .Z(n966) );
  XOR U1494 ( .A(n967), .B(n966), .Z(n969) );
  XOR U1495 ( .A(n968), .B(n969), .Z(n955) );
  NANDN U1496 ( .A(n899), .B(n898), .Z(n903) );
  NANDN U1497 ( .A(n901), .B(n900), .Z(n902) );
  AND U1498 ( .A(n903), .B(n902), .Z(n954) );
  XNOR U1499 ( .A(n955), .B(n954), .Z(n957) );
  NANDN U1500 ( .A(n905), .B(n904), .Z(n909) );
  OR U1501 ( .A(n907), .B(n906), .Z(n908) );
  AND U1502 ( .A(n909), .B(n908), .Z(n961) );
  NAND U1503 ( .A(n186), .B(n910), .Z(n912) );
  XOR U1504 ( .A(b[11]), .B(a[7]), .Z(n980) );
  NAND U1505 ( .A(n37097), .B(n980), .Z(n911) );
  AND U1506 ( .A(n912), .B(n911), .Z(n1001) );
  NAND U1507 ( .A(n187), .B(n913), .Z(n915) );
  XOR U1508 ( .A(b[13]), .B(a[5]), .Z(n1014) );
  NAND U1509 ( .A(n37295), .B(n1014), .Z(n914) );
  AND U1510 ( .A(n915), .B(n914), .Z(n1000) );
  NAND U1511 ( .A(n184), .B(n916), .Z(n918) );
  XOR U1512 ( .A(b[7]), .B(a[11]), .Z(n1008) );
  NAND U1513 ( .A(n36592), .B(n1008), .Z(n917) );
  NAND U1514 ( .A(n918), .B(n917), .Z(n999) );
  XOR U1515 ( .A(n1000), .B(n999), .Z(n1002) );
  XNOR U1516 ( .A(n1001), .B(n1002), .Z(n960) );
  XNOR U1517 ( .A(n961), .B(n960), .Z(n962) );
  NANDN U1518 ( .A(n920), .B(n919), .Z(n924) );
  NANDN U1519 ( .A(n922), .B(n921), .Z(n923) );
  NAND U1520 ( .A(n924), .B(n923), .Z(n963) );
  XNOR U1521 ( .A(n962), .B(n963), .Z(n956) );
  XOR U1522 ( .A(n957), .B(n956), .Z(n1022) );
  NANDN U1523 ( .A(n926), .B(n925), .Z(n930) );
  NANDN U1524 ( .A(n928), .B(n927), .Z(n929) );
  AND U1525 ( .A(n930), .B(n929), .Z(n1021) );
  NANDN U1526 ( .A(n932), .B(n931), .Z(n936) );
  NAND U1527 ( .A(n934), .B(n933), .Z(n935) );
  AND U1528 ( .A(n936), .B(n935), .Z(n1020) );
  XOR U1529 ( .A(n1021), .B(n1020), .Z(n1023) );
  XOR U1530 ( .A(n1022), .B(n1023), .Z(n949) );
  NANDN U1531 ( .A(n938), .B(n937), .Z(n942) );
  OR U1532 ( .A(n940), .B(n939), .Z(n941) );
  AND U1533 ( .A(n942), .B(n941), .Z(n948) );
  XNOR U1534 ( .A(n949), .B(n948), .Z(n950) );
  XNOR U1535 ( .A(n951), .B(n950), .Z(n943) );
  XNOR U1536 ( .A(sreg[241]), .B(n943), .Z(n944) );
  XNOR U1537 ( .A(n945), .B(n944), .Z(c[241]) );
  NANDN U1538 ( .A(sreg[241]), .B(n943), .Z(n947) );
  NAND U1539 ( .A(n945), .B(n944), .Z(n946) );
  NAND U1540 ( .A(n947), .B(n946), .Z(n1112) );
  XNOR U1541 ( .A(sreg[242]), .B(n1112), .Z(n1114) );
  NANDN U1542 ( .A(n949), .B(n948), .Z(n953) );
  NANDN U1543 ( .A(n951), .B(n950), .Z(n952) );
  AND U1544 ( .A(n953), .B(n952), .Z(n1029) );
  NANDN U1545 ( .A(n955), .B(n954), .Z(n959) );
  NAND U1546 ( .A(n957), .B(n956), .Z(n958) );
  AND U1547 ( .A(n959), .B(n958), .Z(n1109) );
  NANDN U1548 ( .A(n961), .B(n960), .Z(n965) );
  NANDN U1549 ( .A(n963), .B(n962), .Z(n964) );
  AND U1550 ( .A(n965), .B(n964), .Z(n1106) );
  NANDN U1551 ( .A(n967), .B(n966), .Z(n971) );
  OR U1552 ( .A(n969), .B(n968), .Z(n970) );
  AND U1553 ( .A(n971), .B(n970), .Z(n1101) );
  NANDN U1554 ( .A(n973), .B(n972), .Z(n977) );
  NAND U1555 ( .A(n975), .B(n974), .Z(n976) );
  NAND U1556 ( .A(n977), .B(n976), .Z(n1100) );
  XNOR U1557 ( .A(n1101), .B(n1100), .Z(n1102) );
  NOR U1558 ( .A(n979), .B(n978), .Z(n1057) );
  NANDN U1559 ( .A(n176), .B(n980), .Z(n982) );
  XNOR U1560 ( .A(b[11]), .B(a[8]), .Z(n1091) );
  OR U1561 ( .A(n1091), .B(n2434), .Z(n981) );
  AND U1562 ( .A(n982), .B(n981), .Z(n1055) );
  XOR U1563 ( .A(b[16]), .B(b[17]), .Z(n983) );
  NANDN U1564 ( .A(n170), .B(n984), .Z(n986) );
  XNOR U1565 ( .A(b[17]), .B(a[2]), .Z(n1042) );
  OR U1566 ( .A(n1042), .B(n36922), .Z(n985) );
  NAND U1567 ( .A(n986), .B(n985), .Z(n1056) );
  XOR U1568 ( .A(n1055), .B(n1056), .Z(n1058) );
  XOR U1569 ( .A(n1057), .B(n1058), .Z(n1033) );
  NAND U1570 ( .A(b[0]), .B(a[18]), .Z(n987) );
  XNOR U1571 ( .A(b[1]), .B(n987), .Z(n989) );
  NANDN U1572 ( .A(b[0]), .B(a[17]), .Z(n988) );
  NAND U1573 ( .A(n989), .B(n988), .Z(n1070) );
  XNOR U1574 ( .A(b[17]), .B(b[18]), .Z(n37589) );
  IV U1575 ( .A(n37589), .Z(n37821) );
  AND U1576 ( .A(a[0]), .B(n37821), .Z(n1067) );
  NAND U1577 ( .A(n188), .B(n990), .Z(n992) );
  XOR U1578 ( .A(b[15]), .B(a[4]), .Z(n1079) );
  NAND U1579 ( .A(n37382), .B(n1079), .Z(n991) );
  AND U1580 ( .A(n992), .B(n991), .Z(n1068) );
  XNOR U1581 ( .A(n1067), .B(n1068), .Z(n1069) );
  XNOR U1582 ( .A(n1070), .B(n1069), .Z(n1032) );
  XNOR U1583 ( .A(n1033), .B(n1032), .Z(n1034) );
  NANDN U1584 ( .A(n994), .B(n993), .Z(n998) );
  OR U1585 ( .A(n996), .B(n995), .Z(n997) );
  NAND U1586 ( .A(n998), .B(n997), .Z(n1035) );
  XNOR U1587 ( .A(n1034), .B(n1035), .Z(n1096) );
  NANDN U1588 ( .A(n1000), .B(n999), .Z(n1004) );
  OR U1589 ( .A(n1002), .B(n1001), .Z(n1003) );
  AND U1590 ( .A(n1004), .B(n1003), .Z(n1095) );
  NAND U1591 ( .A(n183), .B(n1005), .Z(n1007) );
  XOR U1592 ( .A(b[5]), .B(a[14]), .Z(n1082) );
  NAND U1593 ( .A(n36296), .B(n1082), .Z(n1006) );
  AND U1594 ( .A(n1007), .B(n1006), .Z(n1062) );
  NAND U1595 ( .A(n184), .B(n1008), .Z(n1010) );
  XOR U1596 ( .A(b[7]), .B(a[12]), .Z(n1073) );
  NAND U1597 ( .A(n36592), .B(n1073), .Z(n1009) );
  NAND U1598 ( .A(n1010), .B(n1009), .Z(n1061) );
  XNOR U1599 ( .A(n1062), .B(n1061), .Z(n1063) );
  OR U1600 ( .A(n1011), .B(n179), .Z(n1013) );
  XOR U1601 ( .A(b[9]), .B(a[10]), .Z(n1046) );
  NAND U1602 ( .A(n36805), .B(n1046), .Z(n1012) );
  AND U1603 ( .A(n1013), .B(n1012), .Z(n1052) );
  NAND U1604 ( .A(n187), .B(n1014), .Z(n1016) );
  XOR U1605 ( .A(b[13]), .B(a[6]), .Z(n1076) );
  NAND U1606 ( .A(n37295), .B(n1076), .Z(n1015) );
  AND U1607 ( .A(n1016), .B(n1015), .Z(n1050) );
  OR U1608 ( .A(n1017), .B(n180), .Z(n1019) );
  XOR U1609 ( .A(b[3]), .B(a[16]), .Z(n1085) );
  NAND U1610 ( .A(n182), .B(n1085), .Z(n1018) );
  NAND U1611 ( .A(n1019), .B(n1018), .Z(n1049) );
  XNOR U1612 ( .A(n1050), .B(n1049), .Z(n1051) );
  XOR U1613 ( .A(n1052), .B(n1051), .Z(n1064) );
  XNOR U1614 ( .A(n1063), .B(n1064), .Z(n1094) );
  XOR U1615 ( .A(n1095), .B(n1094), .Z(n1097) );
  XOR U1616 ( .A(n1096), .B(n1097), .Z(n1103) );
  XOR U1617 ( .A(n1102), .B(n1103), .Z(n1107) );
  XNOR U1618 ( .A(n1106), .B(n1107), .Z(n1108) );
  XOR U1619 ( .A(n1109), .B(n1108), .Z(n1027) );
  NANDN U1620 ( .A(n1021), .B(n1020), .Z(n1025) );
  OR U1621 ( .A(n1023), .B(n1022), .Z(n1024) );
  AND U1622 ( .A(n1025), .B(n1024), .Z(n1026) );
  XNOR U1623 ( .A(n1027), .B(n1026), .Z(n1028) );
  XNOR U1624 ( .A(n1029), .B(n1028), .Z(n1113) );
  XNOR U1625 ( .A(n1114), .B(n1113), .Z(c[242]) );
  NANDN U1626 ( .A(n1027), .B(n1026), .Z(n1031) );
  NANDN U1627 ( .A(n1029), .B(n1028), .Z(n1030) );
  AND U1628 ( .A(n1031), .B(n1030), .Z(n1124) );
  NANDN U1629 ( .A(n1033), .B(n1032), .Z(n1037) );
  NANDN U1630 ( .A(n1035), .B(n1034), .Z(n1036) );
  AND U1631 ( .A(n1037), .B(n1036), .Z(n1135) );
  XOR U1632 ( .A(b[19]), .B(b[18]), .Z(n1178) );
  XOR U1633 ( .A(b[19]), .B(a[0]), .Z(n1038) );
  NAND U1634 ( .A(n1178), .B(n1038), .Z(n1039) );
  NANDN U1635 ( .A(n1039), .B(n37589), .Z(n1041) );
  XOR U1636 ( .A(b[19]), .B(a[1]), .Z(n1179) );
  NANDN U1637 ( .A(n37589), .B(n1179), .Z(n1040) );
  AND U1638 ( .A(n1041), .B(n1040), .Z(n1174) );
  OR U1639 ( .A(n1042), .B(n170), .Z(n1044) );
  XOR U1640 ( .A(b[17]), .B(a[3]), .Z(n1149) );
  NAND U1641 ( .A(n37652), .B(n1149), .Z(n1043) );
  AND U1642 ( .A(n1044), .B(n1043), .Z(n1173) );
  XOR U1643 ( .A(n1174), .B(n1173), .Z(n1163) );
  NAND U1644 ( .A(b[17]), .B(b[18]), .Z(n1045) );
  NAND U1645 ( .A(b[19]), .B(n1045), .Z(n38045) );
  NOR U1646 ( .A(n38045), .B(n1067), .Z(n1162) );
  NANDN U1647 ( .A(n179), .B(n1046), .Z(n1048) );
  XNOR U1648 ( .A(b[9]), .B(a[11]), .Z(n1182) );
  OR U1649 ( .A(n1182), .B(n2052), .Z(n1047) );
  AND U1650 ( .A(n1048), .B(n1047), .Z(n1161) );
  XOR U1651 ( .A(n1162), .B(n1161), .Z(n1164) );
  XOR U1652 ( .A(n1163), .B(n1164), .Z(n1192) );
  NANDN U1653 ( .A(n1050), .B(n1049), .Z(n1054) );
  NANDN U1654 ( .A(n1052), .B(n1051), .Z(n1053) );
  NAND U1655 ( .A(n1054), .B(n1053), .Z(n1191) );
  XNOR U1656 ( .A(n1192), .B(n1191), .Z(n1193) );
  NANDN U1657 ( .A(n1056), .B(n1055), .Z(n1060) );
  OR U1658 ( .A(n1058), .B(n1057), .Z(n1059) );
  NAND U1659 ( .A(n1060), .B(n1059), .Z(n1194) );
  XNOR U1660 ( .A(n1193), .B(n1194), .Z(n1134) );
  XNOR U1661 ( .A(n1135), .B(n1134), .Z(n1137) );
  NANDN U1662 ( .A(n1062), .B(n1061), .Z(n1066) );
  NANDN U1663 ( .A(n1064), .B(n1063), .Z(n1065) );
  AND U1664 ( .A(n1066), .B(n1065), .Z(n1129) );
  NANDN U1665 ( .A(n1068), .B(n1067), .Z(n1072) );
  NANDN U1666 ( .A(n1070), .B(n1069), .Z(n1071) );
  NAND U1667 ( .A(n1072), .B(n1071), .Z(n1128) );
  XNOR U1668 ( .A(n1129), .B(n1128), .Z(n1130) );
  NAND U1669 ( .A(n184), .B(n1073), .Z(n1075) );
  XOR U1670 ( .A(b[7]), .B(a[13]), .Z(n1155) );
  NAND U1671 ( .A(n36592), .B(n1155), .Z(n1074) );
  AND U1672 ( .A(n1075), .B(n1074), .Z(n1198) );
  NAND U1673 ( .A(n187), .B(n1076), .Z(n1078) );
  XOR U1674 ( .A(b[13]), .B(a[7]), .Z(n1188) );
  NAND U1675 ( .A(n37295), .B(n1188), .Z(n1077) );
  AND U1676 ( .A(n1078), .B(n1077), .Z(n1143) );
  NAND U1677 ( .A(n188), .B(n1079), .Z(n1081) );
  XOR U1678 ( .A(b[15]), .B(a[5]), .Z(n1185) );
  NAND U1679 ( .A(n37382), .B(n1185), .Z(n1080) );
  AND U1680 ( .A(n1081), .B(n1080), .Z(n1141) );
  NAND U1681 ( .A(n183), .B(n1082), .Z(n1084) );
  XOR U1682 ( .A(b[5]), .B(a[15]), .Z(n1152) );
  NAND U1683 ( .A(n36296), .B(n1152), .Z(n1083) );
  NAND U1684 ( .A(n1084), .B(n1083), .Z(n1140) );
  XNOR U1685 ( .A(n1141), .B(n1140), .Z(n1142) );
  XNOR U1686 ( .A(n1143), .B(n1142), .Z(n1197) );
  XNOR U1687 ( .A(n1198), .B(n1197), .Z(n1199) );
  NAND U1688 ( .A(n181), .B(n1085), .Z(n1087) );
  XOR U1689 ( .A(b[3]), .B(a[17]), .Z(n1158) );
  NAND U1690 ( .A(n182), .B(n1158), .Z(n1086) );
  AND U1691 ( .A(n1087), .B(n1086), .Z(n1170) );
  NAND U1692 ( .A(b[0]), .B(a[19]), .Z(n1088) );
  XNOR U1693 ( .A(b[1]), .B(n1088), .Z(n1090) );
  NANDN U1694 ( .A(b[0]), .B(a[18]), .Z(n1089) );
  NAND U1695 ( .A(n1090), .B(n1089), .Z(n1168) );
  OR U1696 ( .A(n1091), .B(n176), .Z(n1093) );
  XOR U1697 ( .A(b[11]), .B(a[9]), .Z(n1175) );
  NAND U1698 ( .A(n37097), .B(n1175), .Z(n1092) );
  NAND U1699 ( .A(n1093), .B(n1092), .Z(n1167) );
  XNOR U1700 ( .A(n1168), .B(n1167), .Z(n1169) );
  XOR U1701 ( .A(n1170), .B(n1169), .Z(n1200) );
  XOR U1702 ( .A(n1199), .B(n1200), .Z(n1131) );
  XNOR U1703 ( .A(n1130), .B(n1131), .Z(n1136) );
  XOR U1704 ( .A(n1137), .B(n1136), .Z(n1204) );
  NANDN U1705 ( .A(n1095), .B(n1094), .Z(n1099) );
  NANDN U1706 ( .A(n1097), .B(n1096), .Z(n1098) );
  AND U1707 ( .A(n1099), .B(n1098), .Z(n1203) );
  XNOR U1708 ( .A(n1204), .B(n1203), .Z(n1205) );
  NANDN U1709 ( .A(n1101), .B(n1100), .Z(n1105) );
  NANDN U1710 ( .A(n1103), .B(n1102), .Z(n1104) );
  NAND U1711 ( .A(n1105), .B(n1104), .Z(n1206) );
  XNOR U1712 ( .A(n1205), .B(n1206), .Z(n1122) );
  NANDN U1713 ( .A(n1107), .B(n1106), .Z(n1111) );
  NAND U1714 ( .A(n1109), .B(n1108), .Z(n1110) );
  NAND U1715 ( .A(n1111), .B(n1110), .Z(n1123) );
  XOR U1716 ( .A(n1122), .B(n1123), .Z(n1125) );
  XOR U1717 ( .A(n1124), .B(n1125), .Z(n1117) );
  XNOR U1718 ( .A(n1117), .B(sreg[243]), .Z(n1119) );
  NANDN U1719 ( .A(sreg[242]), .B(n1112), .Z(n1116) );
  NAND U1720 ( .A(n1114), .B(n1113), .Z(n1115) );
  AND U1721 ( .A(n1116), .B(n1115), .Z(n1118) );
  XOR U1722 ( .A(n1119), .B(n1118), .Z(c[243]) );
  NANDN U1723 ( .A(n1117), .B(sreg[243]), .Z(n1121) );
  NAND U1724 ( .A(n1119), .B(n1118), .Z(n1120) );
  AND U1725 ( .A(n1121), .B(n1120), .Z(n1306) );
  XNOR U1726 ( .A(sreg[244]), .B(n1306), .Z(n1308) );
  NANDN U1727 ( .A(n1123), .B(n1122), .Z(n1127) );
  OR U1728 ( .A(n1125), .B(n1124), .Z(n1126) );
  AND U1729 ( .A(n1127), .B(n1126), .Z(n1212) );
  NANDN U1730 ( .A(n1129), .B(n1128), .Z(n1133) );
  NANDN U1731 ( .A(n1131), .B(n1130), .Z(n1132) );
  AND U1732 ( .A(n1133), .B(n1132), .Z(n1301) );
  NANDN U1733 ( .A(n1135), .B(n1134), .Z(n1139) );
  NAND U1734 ( .A(n1137), .B(n1136), .Z(n1138) );
  NAND U1735 ( .A(n1139), .B(n1138), .Z(n1300) );
  XNOR U1736 ( .A(n1301), .B(n1300), .Z(n1303) );
  NANDN U1737 ( .A(n1141), .B(n1140), .Z(n1145) );
  NANDN U1738 ( .A(n1143), .B(n1142), .Z(n1144) );
  AND U1739 ( .A(n1145), .B(n1144), .Z(n1284) );
  NAND U1740 ( .A(b[0]), .B(a[20]), .Z(n1146) );
  XNOR U1741 ( .A(b[1]), .B(n1146), .Z(n1148) );
  NANDN U1742 ( .A(b[0]), .B(a[19]), .Z(n1147) );
  NAND U1743 ( .A(n1148), .B(n1147), .Z(n1217) );
  XNOR U1744 ( .A(b[19]), .B(b[20]), .Z(n37488) );
  IV U1745 ( .A(n37488), .Z(n37993) );
  AND U1746 ( .A(a[0]), .B(n37993), .Z(n1230) );
  NAND U1747 ( .A(n189), .B(n1149), .Z(n1151) );
  XOR U1748 ( .A(b[17]), .B(a[4]), .Z(n1258) );
  NAND U1749 ( .A(n37652), .B(n1258), .Z(n1150) );
  AND U1750 ( .A(n1151), .B(n1150), .Z(n1215) );
  XNOR U1751 ( .A(n1230), .B(n1215), .Z(n1216) );
  XNOR U1752 ( .A(n1217), .B(n1216), .Z(n1282) );
  NAND U1753 ( .A(n183), .B(n1152), .Z(n1154) );
  XOR U1754 ( .A(b[5]), .B(a[16]), .Z(n1252) );
  NAND U1755 ( .A(n36296), .B(n1252), .Z(n1153) );
  AND U1756 ( .A(n1154), .B(n1153), .Z(n1279) );
  NAND U1757 ( .A(n184), .B(n1155), .Z(n1157) );
  XOR U1758 ( .A(b[7]), .B(a[14]), .Z(n1249) );
  NAND U1759 ( .A(n36592), .B(n1249), .Z(n1156) );
  AND U1760 ( .A(n1157), .B(n1156), .Z(n1277) );
  NAND U1761 ( .A(n181), .B(n1158), .Z(n1160) );
  XOR U1762 ( .A(b[3]), .B(a[18]), .Z(n1234) );
  NAND U1763 ( .A(n182), .B(n1234), .Z(n1159) );
  NAND U1764 ( .A(n1160), .B(n1159), .Z(n1276) );
  XNOR U1765 ( .A(n1277), .B(n1276), .Z(n1278) );
  XOR U1766 ( .A(n1279), .B(n1278), .Z(n1283) );
  XOR U1767 ( .A(n1282), .B(n1283), .Z(n1285) );
  XOR U1768 ( .A(n1284), .B(n1285), .Z(n1290) );
  NANDN U1769 ( .A(n1162), .B(n1161), .Z(n1166) );
  OR U1770 ( .A(n1164), .B(n1163), .Z(n1165) );
  AND U1771 ( .A(n1166), .B(n1165), .Z(n1289) );
  NANDN U1772 ( .A(n1168), .B(n1167), .Z(n1172) );
  NANDN U1773 ( .A(n1170), .B(n1169), .Z(n1171) );
  AND U1774 ( .A(n1172), .B(n1171), .Z(n1266) );
  NOR U1775 ( .A(n1174), .B(n1173), .Z(n1245) );
  NANDN U1776 ( .A(n176), .B(n1175), .Z(n1177) );
  XNOR U1777 ( .A(b[11]), .B(a[10]), .Z(n1231) );
  OR U1778 ( .A(n1231), .B(n2434), .Z(n1176) );
  AND U1779 ( .A(n1177), .B(n1176), .Z(n1243) );
  NANDN U1780 ( .A(n174), .B(n1179), .Z(n1181) );
  XNOR U1781 ( .A(b[19]), .B(a[2]), .Z(n1220) );
  OR U1782 ( .A(n1220), .B(n37589), .Z(n1180) );
  NAND U1783 ( .A(n1181), .B(n1180), .Z(n1244) );
  XOR U1784 ( .A(n1243), .B(n1244), .Z(n1246) );
  XOR U1785 ( .A(n1245), .B(n1246), .Z(n1265) );
  OR U1786 ( .A(n1182), .B(n179), .Z(n1184) );
  XNOR U1787 ( .A(b[9]), .B(a[12]), .Z(n1240) );
  OR U1788 ( .A(n1240), .B(n2052), .Z(n1183) );
  NAND U1789 ( .A(n1184), .B(n1183), .Z(n1271) );
  NAND U1790 ( .A(n188), .B(n1185), .Z(n1187) );
  XOR U1791 ( .A(b[15]), .B(a[6]), .Z(n1261) );
  NAND U1792 ( .A(n37382), .B(n1261), .Z(n1186) );
  NAND U1793 ( .A(n1187), .B(n1186), .Z(n1270) );
  XOR U1794 ( .A(n1271), .B(n1270), .Z(n1273) );
  NANDN U1795 ( .A(n171), .B(n1188), .Z(n1190) );
  XNOR U1796 ( .A(b[13]), .B(a[8]), .Z(n1255) );
  OR U1797 ( .A(n1255), .B(n1681), .Z(n1189) );
  NAND U1798 ( .A(n1190), .B(n1189), .Z(n1272) );
  XOR U1799 ( .A(n1273), .B(n1272), .Z(n1264) );
  XOR U1800 ( .A(n1265), .B(n1264), .Z(n1267) );
  XNOR U1801 ( .A(n1266), .B(n1267), .Z(n1288) );
  XOR U1802 ( .A(n1289), .B(n1288), .Z(n1291) );
  XOR U1803 ( .A(n1290), .B(n1291), .Z(n1297) );
  NANDN U1804 ( .A(n1192), .B(n1191), .Z(n1196) );
  NANDN U1805 ( .A(n1194), .B(n1193), .Z(n1195) );
  AND U1806 ( .A(n1196), .B(n1195), .Z(n1295) );
  NANDN U1807 ( .A(n1198), .B(n1197), .Z(n1202) );
  NANDN U1808 ( .A(n1200), .B(n1199), .Z(n1201) );
  NAND U1809 ( .A(n1202), .B(n1201), .Z(n1294) );
  XNOR U1810 ( .A(n1295), .B(n1294), .Z(n1296) );
  XNOR U1811 ( .A(n1297), .B(n1296), .Z(n1302) );
  XOR U1812 ( .A(n1303), .B(n1302), .Z(n1210) );
  NANDN U1813 ( .A(n1204), .B(n1203), .Z(n1208) );
  NANDN U1814 ( .A(n1206), .B(n1205), .Z(n1207) );
  NAND U1815 ( .A(n1208), .B(n1207), .Z(n1209) );
  XNOR U1816 ( .A(n1210), .B(n1209), .Z(n1211) );
  XNOR U1817 ( .A(n1212), .B(n1211), .Z(n1307) );
  XNOR U1818 ( .A(n1308), .B(n1307), .Z(c[244]) );
  NANDN U1819 ( .A(n1210), .B(n1209), .Z(n1214) );
  NANDN U1820 ( .A(n1212), .B(n1211), .Z(n1213) );
  AND U1821 ( .A(n1214), .B(n1213), .Z(n1319) );
  NANDN U1822 ( .A(n1215), .B(n1230), .Z(n1219) );
  NANDN U1823 ( .A(n1217), .B(n1216), .Z(n1218) );
  NAND U1824 ( .A(n1219), .B(n1218), .Z(n1334) );
  OR U1825 ( .A(n1220), .B(n174), .Z(n1222) );
  XOR U1826 ( .A(b[19]), .B(a[3]), .Z(n1367) );
  NAND U1827 ( .A(n37821), .B(n1367), .Z(n1221) );
  AND U1828 ( .A(n1222), .B(n1221), .Z(n1362) );
  XOR U1829 ( .A(b[21]), .B(a[1]), .Z(n1383) );
  NAND U1830 ( .A(n37993), .B(n1383), .Z(n1229) );
  ANDN U1831 ( .B(b[20]), .A(b[21]), .Z(n1223) );
  NAND U1832 ( .A(n1223), .B(a[0]), .Z(n1226) );
  NAND U1833 ( .A(b[19]), .B(b[20]), .Z(n1224) );
  NAND U1834 ( .A(b[21]), .B(n1224), .Z(n38202) );
  OR U1835 ( .A(a[0]), .B(n38202), .Z(n1225) );
  NAND U1836 ( .A(n1226), .B(n1225), .Z(n1227) );
  NANDN U1837 ( .A(n37993), .B(n1227), .Z(n1228) );
  AND U1838 ( .A(n1229), .B(n1228), .Z(n1363) );
  XOR U1839 ( .A(n1362), .B(n1363), .Z(n1353) );
  NOR U1840 ( .A(n38202), .B(n1230), .Z(n1351) );
  OR U1841 ( .A(n1231), .B(n176), .Z(n1233) );
  XNOR U1842 ( .A(b[11]), .B(a[11]), .Z(n1389) );
  OR U1843 ( .A(n1389), .B(n2434), .Z(n1232) );
  AND U1844 ( .A(n1233), .B(n1232), .Z(n1350) );
  XNOR U1845 ( .A(n1351), .B(n1350), .Z(n1352) );
  XOR U1846 ( .A(n1353), .B(n1352), .Z(n1332) );
  NAND U1847 ( .A(n181), .B(n1234), .Z(n1236) );
  XOR U1848 ( .A(b[3]), .B(a[19]), .Z(n1356) );
  NAND U1849 ( .A(n182), .B(n1356), .Z(n1235) );
  AND U1850 ( .A(n1236), .B(n1235), .Z(n1400) );
  NAND U1851 ( .A(b[0]), .B(a[21]), .Z(n1237) );
  XNOR U1852 ( .A(b[1]), .B(n1237), .Z(n1239) );
  NANDN U1853 ( .A(b[0]), .B(a[20]), .Z(n1238) );
  NAND U1854 ( .A(n1239), .B(n1238), .Z(n1399) );
  OR U1855 ( .A(n1240), .B(n179), .Z(n1242) );
  XOR U1856 ( .A(b[9]), .B(a[13]), .Z(n1386) );
  NAND U1857 ( .A(n36805), .B(n1386), .Z(n1241) );
  NAND U1858 ( .A(n1242), .B(n1241), .Z(n1398) );
  XOR U1859 ( .A(n1399), .B(n1398), .Z(n1401) );
  XOR U1860 ( .A(n1400), .B(n1401), .Z(n1333) );
  XNOR U1861 ( .A(n1332), .B(n1333), .Z(n1335) );
  XOR U1862 ( .A(n1334), .B(n1335), .Z(n1340) );
  NANDN U1863 ( .A(n1244), .B(n1243), .Z(n1248) );
  OR U1864 ( .A(n1246), .B(n1245), .Z(n1247) );
  AND U1865 ( .A(n1248), .B(n1247), .Z(n1339) );
  NAND U1866 ( .A(n184), .B(n1249), .Z(n1251) );
  XOR U1867 ( .A(b[7]), .B(a[15]), .Z(n1370) );
  NAND U1868 ( .A(n36592), .B(n1370), .Z(n1250) );
  AND U1869 ( .A(n1251), .B(n1250), .Z(n1345) );
  NAND U1870 ( .A(n183), .B(n1252), .Z(n1254) );
  XOR U1871 ( .A(b[5]), .B(a[17]), .Z(n1373) );
  NAND U1872 ( .A(n36296), .B(n1373), .Z(n1253) );
  NAND U1873 ( .A(n1254), .B(n1253), .Z(n1344) );
  XNOR U1874 ( .A(n1345), .B(n1344), .Z(n1347) );
  OR U1875 ( .A(n1255), .B(n171), .Z(n1257) );
  XOR U1876 ( .A(b[13]), .B(a[9]), .Z(n1359) );
  NAND U1877 ( .A(n37295), .B(n1359), .Z(n1256) );
  AND U1878 ( .A(n1257), .B(n1256), .Z(n1395) );
  NAND U1879 ( .A(n189), .B(n1258), .Z(n1260) );
  XOR U1880 ( .A(b[17]), .B(a[5]), .Z(n1379) );
  NAND U1881 ( .A(n37652), .B(n1379), .Z(n1259) );
  AND U1882 ( .A(n1260), .B(n1259), .Z(n1393) );
  NAND U1883 ( .A(n188), .B(n1261), .Z(n1263) );
  XOR U1884 ( .A(b[15]), .B(a[7]), .Z(n1376) );
  NAND U1885 ( .A(n37382), .B(n1376), .Z(n1262) );
  NAND U1886 ( .A(n1263), .B(n1262), .Z(n1392) );
  XNOR U1887 ( .A(n1393), .B(n1392), .Z(n1394) );
  XNOR U1888 ( .A(n1395), .B(n1394), .Z(n1346) );
  XNOR U1889 ( .A(n1347), .B(n1346), .Z(n1338) );
  XOR U1890 ( .A(n1339), .B(n1338), .Z(n1341) );
  XNOR U1891 ( .A(n1340), .B(n1341), .Z(n1322) );
  NANDN U1892 ( .A(n1265), .B(n1264), .Z(n1269) );
  OR U1893 ( .A(n1267), .B(n1266), .Z(n1268) );
  NAND U1894 ( .A(n1269), .B(n1268), .Z(n1323) );
  XNOR U1895 ( .A(n1322), .B(n1323), .Z(n1325) );
  NAND U1896 ( .A(n1271), .B(n1270), .Z(n1275) );
  NAND U1897 ( .A(n1273), .B(n1272), .Z(n1274) );
  NAND U1898 ( .A(n1275), .B(n1274), .Z(n1327) );
  NANDN U1899 ( .A(n1277), .B(n1276), .Z(n1281) );
  NANDN U1900 ( .A(n1279), .B(n1278), .Z(n1280) );
  NAND U1901 ( .A(n1281), .B(n1280), .Z(n1326) );
  XOR U1902 ( .A(n1327), .B(n1326), .Z(n1329) );
  NANDN U1903 ( .A(n1283), .B(n1282), .Z(n1287) );
  OR U1904 ( .A(n1285), .B(n1284), .Z(n1286) );
  NAND U1905 ( .A(n1287), .B(n1286), .Z(n1328) );
  XOR U1906 ( .A(n1329), .B(n1328), .Z(n1324) );
  XOR U1907 ( .A(n1325), .B(n1324), .Z(n1405) );
  NANDN U1908 ( .A(n1289), .B(n1288), .Z(n1293) );
  OR U1909 ( .A(n1291), .B(n1290), .Z(n1292) );
  NAND U1910 ( .A(n1293), .B(n1292), .Z(n1404) );
  XNOR U1911 ( .A(n1405), .B(n1404), .Z(n1406) );
  NANDN U1912 ( .A(n1295), .B(n1294), .Z(n1299) );
  NANDN U1913 ( .A(n1297), .B(n1296), .Z(n1298) );
  NAND U1914 ( .A(n1299), .B(n1298), .Z(n1407) );
  XNOR U1915 ( .A(n1406), .B(n1407), .Z(n1316) );
  NANDN U1916 ( .A(n1301), .B(n1300), .Z(n1305) );
  NAND U1917 ( .A(n1303), .B(n1302), .Z(n1304) );
  NAND U1918 ( .A(n1305), .B(n1304), .Z(n1317) );
  XNOR U1919 ( .A(n1316), .B(n1317), .Z(n1318) );
  XNOR U1920 ( .A(n1319), .B(n1318), .Z(n1311) );
  XNOR U1921 ( .A(sreg[245]), .B(n1311), .Z(n1313) );
  NANDN U1922 ( .A(sreg[244]), .B(n1306), .Z(n1310) );
  NAND U1923 ( .A(n1308), .B(n1307), .Z(n1309) );
  NAND U1924 ( .A(n1310), .B(n1309), .Z(n1312) );
  XNOR U1925 ( .A(n1313), .B(n1312), .Z(c[245]) );
  NANDN U1926 ( .A(sreg[245]), .B(n1311), .Z(n1315) );
  NAND U1927 ( .A(n1313), .B(n1312), .Z(n1314) );
  NAND U1928 ( .A(n1315), .B(n1314), .Z(n1514) );
  XNOR U1929 ( .A(sreg[246]), .B(n1514), .Z(n1516) );
  NANDN U1930 ( .A(n1317), .B(n1316), .Z(n1321) );
  NANDN U1931 ( .A(n1319), .B(n1318), .Z(n1320) );
  AND U1932 ( .A(n1321), .B(n1320), .Z(n1413) );
  NAND U1933 ( .A(n1327), .B(n1326), .Z(n1331) );
  NAND U1934 ( .A(n1329), .B(n1328), .Z(n1330) );
  NAND U1935 ( .A(n1331), .B(n1330), .Z(n1508) );
  XNOR U1936 ( .A(n1509), .B(n1508), .Z(n1511) );
  NAND U1937 ( .A(n1333), .B(n1332), .Z(n1337) );
  NANDN U1938 ( .A(n1335), .B(n1334), .Z(n1336) );
  AND U1939 ( .A(n1337), .B(n1336), .Z(n1417) );
  NANDN U1940 ( .A(n1339), .B(n1338), .Z(n1343) );
  NANDN U1941 ( .A(n1341), .B(n1340), .Z(n1342) );
  AND U1942 ( .A(n1343), .B(n1342), .Z(n1416) );
  XNOR U1943 ( .A(n1417), .B(n1416), .Z(n1418) );
  NANDN U1944 ( .A(n1345), .B(n1344), .Z(n1349) );
  NAND U1945 ( .A(n1347), .B(n1346), .Z(n1348) );
  AND U1946 ( .A(n1349), .B(n1348), .Z(n1423) );
  NANDN U1947 ( .A(n1351), .B(n1350), .Z(n1355) );
  NANDN U1948 ( .A(n1353), .B(n1352), .Z(n1354) );
  AND U1949 ( .A(n1355), .B(n1354), .Z(n1430) );
  NAND U1950 ( .A(n181), .B(n1356), .Z(n1358) );
  XOR U1951 ( .A(b[3]), .B(a[20]), .Z(n1451) );
  NAND U1952 ( .A(n182), .B(n1451), .Z(n1357) );
  AND U1953 ( .A(n1358), .B(n1357), .Z(n1491) );
  NAND U1954 ( .A(n187), .B(n1359), .Z(n1361) );
  XOR U1955 ( .A(b[13]), .B(a[10]), .Z(n1465) );
  NAND U1956 ( .A(n37295), .B(n1465), .Z(n1360) );
  NAND U1957 ( .A(n1361), .B(n1360), .Z(n1490) );
  XNOR U1958 ( .A(n1491), .B(n1490), .Z(n1493) );
  NOR U1959 ( .A(n1363), .B(n1362), .Z(n1492) );
  XOR U1960 ( .A(n1493), .B(n1492), .Z(n1429) );
  NAND U1961 ( .A(b[0]), .B(a[22]), .Z(n1364) );
  XNOR U1962 ( .A(b[1]), .B(n1364), .Z(n1366) );
  NANDN U1963 ( .A(b[0]), .B(a[21]), .Z(n1365) );
  NAND U1964 ( .A(n1366), .B(n1365), .Z(n1448) );
  XNOR U1965 ( .A(b[21]), .B(b[22]), .Z(n37306) );
  IV U1966 ( .A(n37306), .Z(n38132) );
  AND U1967 ( .A(a[0]), .B(n38132), .Z(n1458) );
  NAND U1968 ( .A(n190), .B(n1367), .Z(n1369) );
  XOR U1969 ( .A(b[19]), .B(a[4]), .Z(n1462) );
  NAND U1970 ( .A(n37821), .B(n1462), .Z(n1368) );
  AND U1971 ( .A(n1369), .B(n1368), .Z(n1446) );
  XOR U1972 ( .A(n1458), .B(n1446), .Z(n1447) );
  XNOR U1973 ( .A(n1448), .B(n1447), .Z(n1428) );
  XOR U1974 ( .A(n1429), .B(n1428), .Z(n1431) );
  XNOR U1975 ( .A(n1430), .B(n1431), .Z(n1422) );
  XNOR U1976 ( .A(n1423), .B(n1422), .Z(n1424) );
  NAND U1977 ( .A(n184), .B(n1370), .Z(n1372) );
  XOR U1978 ( .A(b[7]), .B(a[16]), .Z(n1481) );
  NAND U1979 ( .A(n36592), .B(n1481), .Z(n1371) );
  AND U1980 ( .A(n1372), .B(n1371), .Z(n1504) );
  NAND U1981 ( .A(n183), .B(n1373), .Z(n1375) );
  XOR U1982 ( .A(b[5]), .B(a[18]), .Z(n1487) );
  NAND U1983 ( .A(n36296), .B(n1487), .Z(n1374) );
  AND U1984 ( .A(n1375), .B(n1374), .Z(n1503) );
  NAND U1985 ( .A(n188), .B(n1376), .Z(n1378) );
  XOR U1986 ( .A(b[15]), .B(a[8]), .Z(n1454) );
  NAND U1987 ( .A(n37382), .B(n1454), .Z(n1377) );
  NAND U1988 ( .A(n1378), .B(n1377), .Z(n1502) );
  XOR U1989 ( .A(n1503), .B(n1502), .Z(n1505) );
  XOR U1990 ( .A(n1504), .B(n1505), .Z(n1442) );
  NAND U1991 ( .A(n189), .B(n1379), .Z(n1381) );
  XOR U1992 ( .A(b[17]), .B(a[6]), .Z(n1459) );
  NAND U1993 ( .A(n37652), .B(n1459), .Z(n1380) );
  AND U1994 ( .A(n1381), .B(n1380), .Z(n1498) );
  XOR U1995 ( .A(b[20]), .B(b[21]), .Z(n1382) );
  AND U1996 ( .A(n1382), .B(n37488), .Z(n38064) );
  NAND U1997 ( .A(n38064), .B(n1383), .Z(n1385) );
  XOR U1998 ( .A(b[21]), .B(a[2]), .Z(n1474) );
  NAND U1999 ( .A(n37993), .B(n1474), .Z(n1384) );
  AND U2000 ( .A(n1385), .B(n1384), .Z(n1497) );
  NAND U2001 ( .A(n185), .B(n1386), .Z(n1388) );
  XOR U2002 ( .A(b[9]), .B(a[14]), .Z(n1484) );
  NAND U2003 ( .A(n36805), .B(n1484), .Z(n1387) );
  NAND U2004 ( .A(n1388), .B(n1387), .Z(n1496) );
  XOR U2005 ( .A(n1497), .B(n1496), .Z(n1499) );
  XOR U2006 ( .A(n1498), .B(n1499), .Z(n1441) );
  OR U2007 ( .A(n1389), .B(n176), .Z(n1391) );
  XNOR U2008 ( .A(b[11]), .B(a[12]), .Z(n1468) );
  OR U2009 ( .A(n1468), .B(n2434), .Z(n1390) );
  AND U2010 ( .A(n1391), .B(n1390), .Z(n1440) );
  XOR U2011 ( .A(n1441), .B(n1440), .Z(n1443) );
  XOR U2012 ( .A(n1442), .B(n1443), .Z(n1437) );
  NANDN U2013 ( .A(n1393), .B(n1392), .Z(n1397) );
  NANDN U2014 ( .A(n1395), .B(n1394), .Z(n1396) );
  AND U2015 ( .A(n1397), .B(n1396), .Z(n1435) );
  NANDN U2016 ( .A(n1399), .B(n1398), .Z(n1403) );
  OR U2017 ( .A(n1401), .B(n1400), .Z(n1402) );
  NAND U2018 ( .A(n1403), .B(n1402), .Z(n1434) );
  XNOR U2019 ( .A(n1435), .B(n1434), .Z(n1436) );
  XOR U2020 ( .A(n1437), .B(n1436), .Z(n1425) );
  XOR U2021 ( .A(n1424), .B(n1425), .Z(n1419) );
  XNOR U2022 ( .A(n1418), .B(n1419), .Z(n1510) );
  XOR U2023 ( .A(n1511), .B(n1510), .Z(n1411) );
  NANDN U2024 ( .A(n1405), .B(n1404), .Z(n1409) );
  NANDN U2025 ( .A(n1407), .B(n1406), .Z(n1408) );
  NAND U2026 ( .A(n1409), .B(n1408), .Z(n1410) );
  XNOR U2027 ( .A(n1411), .B(n1410), .Z(n1412) );
  XNOR U2028 ( .A(n1413), .B(n1412), .Z(n1515) );
  XNOR U2029 ( .A(n1516), .B(n1515), .Z(c[246]) );
  NANDN U2030 ( .A(n1411), .B(n1410), .Z(n1415) );
  NANDN U2031 ( .A(n1413), .B(n1412), .Z(n1414) );
  AND U2032 ( .A(n1415), .B(n1414), .Z(n1527) );
  NANDN U2033 ( .A(n1417), .B(n1416), .Z(n1421) );
  NANDN U2034 ( .A(n1419), .B(n1418), .Z(n1420) );
  AND U2035 ( .A(n1421), .B(n1420), .Z(n1625) );
  NANDN U2036 ( .A(n1423), .B(n1422), .Z(n1427) );
  NANDN U2037 ( .A(n1425), .B(n1424), .Z(n1426) );
  AND U2038 ( .A(n1427), .B(n1426), .Z(n1533) );
  NANDN U2039 ( .A(n1429), .B(n1428), .Z(n1433) );
  OR U2040 ( .A(n1431), .B(n1430), .Z(n1432) );
  AND U2041 ( .A(n1433), .B(n1432), .Z(n1531) );
  NANDN U2042 ( .A(n1435), .B(n1434), .Z(n1439) );
  NANDN U2043 ( .A(n1437), .B(n1436), .Z(n1438) );
  AND U2044 ( .A(n1439), .B(n1438), .Z(n1530) );
  XNOR U2045 ( .A(n1531), .B(n1530), .Z(n1532) );
  XOR U2046 ( .A(n1533), .B(n1532), .Z(n1624) );
  NANDN U2047 ( .A(n1441), .B(n1440), .Z(n1445) );
  OR U2048 ( .A(n1443), .B(n1442), .Z(n1444) );
  AND U2049 ( .A(n1445), .B(n1444), .Z(n1617) );
  NANDN U2050 ( .A(n1446), .B(n1458), .Z(n1450) );
  OR U2051 ( .A(n1448), .B(n1447), .Z(n1449) );
  AND U2052 ( .A(n1450), .B(n1449), .Z(n1614) );
  NAND U2053 ( .A(n181), .B(n1451), .Z(n1453) );
  XOR U2054 ( .A(b[3]), .B(a[21]), .Z(n1553) );
  NAND U2055 ( .A(n182), .B(n1553), .Z(n1452) );
  AND U2056 ( .A(n1453), .B(n1452), .Z(n1565) );
  NAND U2057 ( .A(n188), .B(n1454), .Z(n1456) );
  XOR U2058 ( .A(b[15]), .B(a[9]), .Z(n1589) );
  NAND U2059 ( .A(n37382), .B(n1589), .Z(n1455) );
  AND U2060 ( .A(n1456), .B(n1455), .Z(n1563) );
  NAND U2061 ( .A(b[21]), .B(b[22]), .Z(n1457) );
  AND U2062 ( .A(b[23]), .B(n1457), .Z(n38253) );
  IV U2063 ( .A(n38253), .Z(n38298) );
  NOR U2064 ( .A(n38298), .B(n1458), .Z(n1562) );
  XNOR U2065 ( .A(n1563), .B(n1562), .Z(n1564) );
  XNOR U2066 ( .A(n1565), .B(n1564), .Z(n1611) );
  NAND U2067 ( .A(n189), .B(n1459), .Z(n1461) );
  XOR U2068 ( .A(b[17]), .B(a[7]), .Z(n1586) );
  NAND U2069 ( .A(n37652), .B(n1586), .Z(n1460) );
  AND U2070 ( .A(n1461), .B(n1460), .Z(n1545) );
  NAND U2071 ( .A(n190), .B(n1462), .Z(n1464) );
  XOR U2072 ( .A(b[19]), .B(a[5]), .Z(n1595) );
  NAND U2073 ( .A(n37821), .B(n1595), .Z(n1463) );
  AND U2074 ( .A(n1464), .B(n1463), .Z(n1543) );
  NAND U2075 ( .A(n187), .B(n1465), .Z(n1467) );
  XOR U2076 ( .A(b[13]), .B(a[11]), .Z(n1550) );
  NAND U2077 ( .A(n37295), .B(n1550), .Z(n1466) );
  NAND U2078 ( .A(n1467), .B(n1466), .Z(n1542) );
  XNOR U2079 ( .A(n1543), .B(n1542), .Z(n1544) );
  XOR U2080 ( .A(n1545), .B(n1544), .Z(n1612) );
  XNOR U2081 ( .A(n1611), .B(n1612), .Z(n1613) );
  XOR U2082 ( .A(n1614), .B(n1613), .Z(n1618) );
  XNOR U2083 ( .A(n1617), .B(n1618), .Z(n1619) );
  OR U2084 ( .A(n1468), .B(n176), .Z(n1470) );
  XOR U2085 ( .A(b[11]), .B(a[13]), .Z(n1592) );
  NAND U2086 ( .A(n37097), .B(n1592), .Z(n1469) );
  NAND U2087 ( .A(n1470), .B(n1469), .Z(n1556) );
  NAND U2088 ( .A(b[0]), .B(a[23]), .Z(n1471) );
  XNOR U2089 ( .A(b[1]), .B(n1471), .Z(n1473) );
  NANDN U2090 ( .A(b[0]), .B(a[22]), .Z(n1472) );
  NAND U2091 ( .A(n1473), .B(n1472), .Z(n1557) );
  XNOR U2092 ( .A(n1556), .B(n1557), .Z(n1558) );
  NAND U2093 ( .A(n38064), .B(n1474), .Z(n1476) );
  XOR U2094 ( .A(b[21]), .B(a[3]), .Z(n1577) );
  NAND U2095 ( .A(n37993), .B(n1577), .Z(n1475) );
  AND U2096 ( .A(n1476), .B(n1475), .Z(n1548) );
  XOR U2097 ( .A(b[23]), .B(b[22]), .Z(n1598) );
  XOR U2098 ( .A(b[23]), .B(a[0]), .Z(n1477) );
  NAND U2099 ( .A(n1598), .B(n1477), .Z(n1478) );
  NANDN U2100 ( .A(n1478), .B(n37306), .Z(n1480) );
  XOR U2101 ( .A(b[23]), .B(a[1]), .Z(n1599) );
  NANDN U2102 ( .A(n37306), .B(n1599), .Z(n1479) );
  NAND U2103 ( .A(n1480), .B(n1479), .Z(n1549) );
  XOR U2104 ( .A(n1548), .B(n1549), .Z(n1559) );
  XNOR U2105 ( .A(n1558), .B(n1559), .Z(n1606) );
  NAND U2106 ( .A(n184), .B(n1481), .Z(n1483) );
  XOR U2107 ( .A(b[7]), .B(a[17]), .Z(n1580) );
  NAND U2108 ( .A(n36592), .B(n1580), .Z(n1482) );
  AND U2109 ( .A(n1483), .B(n1482), .Z(n1570) );
  NAND U2110 ( .A(n185), .B(n1484), .Z(n1486) );
  XOR U2111 ( .A(b[9]), .B(a[15]), .Z(n1602) );
  NAND U2112 ( .A(n36805), .B(n1602), .Z(n1485) );
  AND U2113 ( .A(n1486), .B(n1485), .Z(n1569) );
  NAND U2114 ( .A(n183), .B(n1487), .Z(n1489) );
  XOR U2115 ( .A(b[5]), .B(a[19]), .Z(n1583) );
  NAND U2116 ( .A(n36296), .B(n1583), .Z(n1488) );
  NAND U2117 ( .A(n1489), .B(n1488), .Z(n1568) );
  XOR U2118 ( .A(n1569), .B(n1568), .Z(n1571) );
  XOR U2119 ( .A(n1570), .B(n1571), .Z(n1605) );
  XOR U2120 ( .A(n1606), .B(n1605), .Z(n1608) );
  NANDN U2121 ( .A(n1491), .B(n1490), .Z(n1495) );
  NAND U2122 ( .A(n1493), .B(n1492), .Z(n1494) );
  NAND U2123 ( .A(n1495), .B(n1494), .Z(n1607) );
  XOR U2124 ( .A(n1608), .B(n1607), .Z(n1538) );
  NANDN U2125 ( .A(n1497), .B(n1496), .Z(n1501) );
  OR U2126 ( .A(n1499), .B(n1498), .Z(n1500) );
  AND U2127 ( .A(n1501), .B(n1500), .Z(n1537) );
  NANDN U2128 ( .A(n1503), .B(n1502), .Z(n1507) );
  OR U2129 ( .A(n1505), .B(n1504), .Z(n1506) );
  NAND U2130 ( .A(n1507), .B(n1506), .Z(n1536) );
  XOR U2131 ( .A(n1537), .B(n1536), .Z(n1539) );
  XOR U2132 ( .A(n1538), .B(n1539), .Z(n1620) );
  XNOR U2133 ( .A(n1619), .B(n1620), .Z(n1623) );
  XOR U2134 ( .A(n1624), .B(n1623), .Z(n1626) );
  XOR U2135 ( .A(n1625), .B(n1626), .Z(n1525) );
  NANDN U2136 ( .A(n1509), .B(n1508), .Z(n1513) );
  NAND U2137 ( .A(n1511), .B(n1510), .Z(n1512) );
  AND U2138 ( .A(n1513), .B(n1512), .Z(n1524) );
  XNOR U2139 ( .A(n1525), .B(n1524), .Z(n1526) );
  XNOR U2140 ( .A(n1527), .B(n1526), .Z(n1519) );
  XNOR U2141 ( .A(sreg[247]), .B(n1519), .Z(n1521) );
  NANDN U2142 ( .A(sreg[246]), .B(n1514), .Z(n1518) );
  NAND U2143 ( .A(n1516), .B(n1515), .Z(n1517) );
  NAND U2144 ( .A(n1518), .B(n1517), .Z(n1520) );
  XNOR U2145 ( .A(n1521), .B(n1520), .Z(c[247]) );
  NANDN U2146 ( .A(sreg[247]), .B(n1519), .Z(n1523) );
  NAND U2147 ( .A(n1521), .B(n1520), .Z(n1522) );
  NAND U2148 ( .A(n1523), .B(n1522), .Z(n1743) );
  XNOR U2149 ( .A(sreg[248]), .B(n1743), .Z(n1745) );
  NANDN U2150 ( .A(n1525), .B(n1524), .Z(n1529) );
  NANDN U2151 ( .A(n1527), .B(n1526), .Z(n1528) );
  AND U2152 ( .A(n1529), .B(n1528), .Z(n1632) );
  NANDN U2153 ( .A(n1531), .B(n1530), .Z(n1535) );
  NAND U2154 ( .A(n1533), .B(n1532), .Z(n1534) );
  AND U2155 ( .A(n1535), .B(n1534), .Z(n1638) );
  NANDN U2156 ( .A(n1537), .B(n1536), .Z(n1541) );
  NANDN U2157 ( .A(n1539), .B(n1538), .Z(n1540) );
  AND U2158 ( .A(n1541), .B(n1540), .Z(n1739) );
  NANDN U2159 ( .A(n1543), .B(n1542), .Z(n1547) );
  NANDN U2160 ( .A(n1545), .B(n1544), .Z(n1546) );
  AND U2161 ( .A(n1547), .B(n1546), .Z(n1653) );
  ANDN U2162 ( .B(n1549), .A(n1548), .Z(n1695) );
  NANDN U2163 ( .A(n171), .B(n1550), .Z(n1552) );
  XNOR U2164 ( .A(b[13]), .B(a[12]), .Z(n1680) );
  OR U2165 ( .A(n1680), .B(n1681), .Z(n1551) );
  AND U2166 ( .A(n1552), .B(n1551), .Z(n1692) );
  NANDN U2167 ( .A(n180), .B(n1553), .Z(n1555) );
  XNOR U2168 ( .A(b[3]), .B(a[22]), .Z(n1684) );
  OR U2169 ( .A(n1684), .B(n172), .Z(n1554) );
  NAND U2170 ( .A(n1555), .B(n1554), .Z(n1693) );
  XNOR U2171 ( .A(n1692), .B(n1693), .Z(n1694) );
  XOR U2172 ( .A(n1695), .B(n1694), .Z(n1654) );
  XNOR U2173 ( .A(n1653), .B(n1654), .Z(n1656) );
  NANDN U2174 ( .A(n1557), .B(n1556), .Z(n1561) );
  NANDN U2175 ( .A(n1559), .B(n1558), .Z(n1560) );
  AND U2176 ( .A(n1561), .B(n1560), .Z(n1655) );
  XOR U2177 ( .A(n1656), .B(n1655), .Z(n1738) );
  NANDN U2178 ( .A(n1563), .B(n1562), .Z(n1567) );
  NANDN U2179 ( .A(n1565), .B(n1564), .Z(n1566) );
  AND U2180 ( .A(n1567), .B(n1566), .Z(n1648) );
  NANDN U2181 ( .A(n1569), .B(n1568), .Z(n1573) );
  OR U2182 ( .A(n1571), .B(n1570), .Z(n1572) );
  NAND U2183 ( .A(n1573), .B(n1572), .Z(n1647) );
  XNOR U2184 ( .A(n1648), .B(n1647), .Z(n1649) );
  NAND U2185 ( .A(b[0]), .B(a[24]), .Z(n1574) );
  XNOR U2186 ( .A(b[1]), .B(n1574), .Z(n1576) );
  NANDN U2187 ( .A(b[0]), .B(a[23]), .Z(n1575) );
  NAND U2188 ( .A(n1576), .B(n1575), .Z(n1667) );
  XNOR U2189 ( .A(b[23]), .B(b[24]), .Z(n37513) );
  IV U2190 ( .A(n37513), .Z(n38247) );
  AND U2191 ( .A(a[0]), .B(n38247), .Z(n1691) );
  NAND U2192 ( .A(n38064), .B(n1577), .Z(n1579) );
  XOR U2193 ( .A(b[21]), .B(a[4]), .Z(n1728) );
  NAND U2194 ( .A(n37993), .B(n1728), .Z(n1578) );
  AND U2195 ( .A(n1579), .B(n1578), .Z(n1665) );
  XNOR U2196 ( .A(n1691), .B(n1665), .Z(n1666) );
  XNOR U2197 ( .A(n1667), .B(n1666), .Z(n1659) );
  NAND U2198 ( .A(n184), .B(n1580), .Z(n1582) );
  XOR U2199 ( .A(b[7]), .B(a[18]), .Z(n1716) );
  NAND U2200 ( .A(n36592), .B(n1716), .Z(n1581) );
  AND U2201 ( .A(n1582), .B(n1581), .Z(n1713) );
  NAND U2202 ( .A(n183), .B(n1583), .Z(n1585) );
  XOR U2203 ( .A(b[5]), .B(a[20]), .Z(n1719) );
  NAND U2204 ( .A(n36296), .B(n1719), .Z(n1584) );
  AND U2205 ( .A(n1585), .B(n1584), .Z(n1711) );
  NAND U2206 ( .A(n189), .B(n1586), .Z(n1588) );
  XOR U2207 ( .A(b[17]), .B(a[8]), .Z(n1722) );
  NAND U2208 ( .A(n37652), .B(n1722), .Z(n1587) );
  NAND U2209 ( .A(n1588), .B(n1587), .Z(n1710) );
  XNOR U2210 ( .A(n1711), .B(n1710), .Z(n1712) );
  XOR U2211 ( .A(n1713), .B(n1712), .Z(n1660) );
  XNOR U2212 ( .A(n1659), .B(n1660), .Z(n1661) );
  NAND U2213 ( .A(n188), .B(n1589), .Z(n1591) );
  XOR U2214 ( .A(b[15]), .B(a[10]), .Z(n1687) );
  NAND U2215 ( .A(n37382), .B(n1687), .Z(n1590) );
  AND U2216 ( .A(n1591), .B(n1590), .Z(n1705) );
  NAND U2217 ( .A(n186), .B(n1592), .Z(n1594) );
  XOR U2218 ( .A(b[11]), .B(a[14]), .Z(n1734) );
  NAND U2219 ( .A(n37097), .B(n1734), .Z(n1593) );
  NAND U2220 ( .A(n1594), .B(n1593), .Z(n1704) );
  XNOR U2221 ( .A(n1705), .B(n1704), .Z(n1706) );
  NAND U2222 ( .A(n190), .B(n1595), .Z(n1597) );
  XOR U2223 ( .A(b[19]), .B(a[6]), .Z(n1725) );
  NAND U2224 ( .A(n37821), .B(n1725), .Z(n1596) );
  AND U2225 ( .A(n1597), .B(n1596), .Z(n1701) );
  AND U2226 ( .A(n1598), .B(n37306), .Z(n38185) );
  NAND U2227 ( .A(n38185), .B(n1599), .Z(n1601) );
  XOR U2228 ( .A(b[23]), .B(a[2]), .Z(n1670) );
  NAND U2229 ( .A(n38132), .B(n1670), .Z(n1600) );
  AND U2230 ( .A(n1601), .B(n1600), .Z(n1699) );
  NAND U2231 ( .A(n185), .B(n1602), .Z(n1604) );
  XOR U2232 ( .A(b[9]), .B(a[16]), .Z(n1731) );
  NAND U2233 ( .A(n36805), .B(n1731), .Z(n1603) );
  NAND U2234 ( .A(n1604), .B(n1603), .Z(n1698) );
  XNOR U2235 ( .A(n1699), .B(n1698), .Z(n1700) );
  XOR U2236 ( .A(n1701), .B(n1700), .Z(n1707) );
  XOR U2237 ( .A(n1706), .B(n1707), .Z(n1662) );
  XOR U2238 ( .A(n1661), .B(n1662), .Z(n1650) );
  XNOR U2239 ( .A(n1649), .B(n1650), .Z(n1737) );
  XOR U2240 ( .A(n1738), .B(n1737), .Z(n1740) );
  XOR U2241 ( .A(n1739), .B(n1740), .Z(n1644) );
  NAND U2242 ( .A(n1606), .B(n1605), .Z(n1610) );
  NAND U2243 ( .A(n1608), .B(n1607), .Z(n1609) );
  AND U2244 ( .A(n1610), .B(n1609), .Z(n1641) );
  NANDN U2245 ( .A(n1612), .B(n1611), .Z(n1616) );
  NANDN U2246 ( .A(n1614), .B(n1613), .Z(n1615) );
  NAND U2247 ( .A(n1616), .B(n1615), .Z(n1642) );
  XNOR U2248 ( .A(n1641), .B(n1642), .Z(n1643) );
  XNOR U2249 ( .A(n1644), .B(n1643), .Z(n1635) );
  NANDN U2250 ( .A(n1618), .B(n1617), .Z(n1622) );
  NANDN U2251 ( .A(n1620), .B(n1619), .Z(n1621) );
  NAND U2252 ( .A(n1622), .B(n1621), .Z(n1636) );
  XNOR U2253 ( .A(n1635), .B(n1636), .Z(n1637) );
  XNOR U2254 ( .A(n1638), .B(n1637), .Z(n1629) );
  NANDN U2255 ( .A(n1624), .B(n1623), .Z(n1628) );
  OR U2256 ( .A(n1626), .B(n1625), .Z(n1627) );
  NAND U2257 ( .A(n1628), .B(n1627), .Z(n1630) );
  XNOR U2258 ( .A(n1629), .B(n1630), .Z(n1631) );
  XNOR U2259 ( .A(n1632), .B(n1631), .Z(n1744) );
  XNOR U2260 ( .A(n1745), .B(n1744), .Z(c[248]) );
  NANDN U2261 ( .A(n1630), .B(n1629), .Z(n1634) );
  NANDN U2262 ( .A(n1632), .B(n1631), .Z(n1633) );
  AND U2263 ( .A(n1634), .B(n1633), .Z(n1756) );
  NANDN U2264 ( .A(n1636), .B(n1635), .Z(n1640) );
  NANDN U2265 ( .A(n1638), .B(n1637), .Z(n1639) );
  AND U2266 ( .A(n1640), .B(n1639), .Z(n1754) );
  NANDN U2267 ( .A(n1642), .B(n1641), .Z(n1646) );
  NANDN U2268 ( .A(n1644), .B(n1643), .Z(n1645) );
  AND U2269 ( .A(n1646), .B(n1645), .Z(n1762) );
  NANDN U2270 ( .A(n1648), .B(n1647), .Z(n1652) );
  NANDN U2271 ( .A(n1650), .B(n1649), .Z(n1651) );
  AND U2272 ( .A(n1652), .B(n1651), .Z(n1862) );
  NANDN U2273 ( .A(n1654), .B(n1653), .Z(n1658) );
  NAND U2274 ( .A(n1656), .B(n1655), .Z(n1657) );
  AND U2275 ( .A(n1658), .B(n1657), .Z(n1861) );
  XNOR U2276 ( .A(n1862), .B(n1861), .Z(n1864) );
  NANDN U2277 ( .A(n1660), .B(n1659), .Z(n1664) );
  NANDN U2278 ( .A(n1662), .B(n1661), .Z(n1663) );
  AND U2279 ( .A(n1664), .B(n1663), .Z(n1856) );
  NANDN U2280 ( .A(n1665), .B(n1691), .Z(n1669) );
  NANDN U2281 ( .A(n1667), .B(n1666), .Z(n1668) );
  AND U2282 ( .A(n1669), .B(n1668), .Z(n1779) );
  NAND U2283 ( .A(n38185), .B(n1670), .Z(n1672) );
  XOR U2284 ( .A(b[23]), .B(a[3]), .Z(n1817) );
  NAND U2285 ( .A(n38132), .B(n1817), .Z(n1671) );
  AND U2286 ( .A(n1672), .B(n1671), .Z(n1832) );
  XOR U2287 ( .A(b[25]), .B(b[24]), .Z(n1792) );
  XOR U2288 ( .A(b[25]), .B(a[0]), .Z(n1673) );
  NAND U2289 ( .A(n1792), .B(n1673), .Z(n1674) );
  NANDN U2290 ( .A(n1674), .B(n37513), .Z(n1676) );
  XOR U2291 ( .A(b[25]), .B(a[1]), .Z(n1793) );
  NANDN U2292 ( .A(n37513), .B(n1793), .Z(n1675) );
  AND U2293 ( .A(n1676), .B(n1675), .Z(n1833) );
  XOR U2294 ( .A(n1832), .B(n1833), .Z(n1785) );
  NAND U2295 ( .A(b[0]), .B(a[25]), .Z(n1677) );
  XNOR U2296 ( .A(b[1]), .B(n1677), .Z(n1679) );
  NANDN U2297 ( .A(b[0]), .B(a[24]), .Z(n1678) );
  NAND U2298 ( .A(n1679), .B(n1678), .Z(n1783) );
  OR U2299 ( .A(n1680), .B(n171), .Z(n1683) );
  XNOR U2300 ( .A(b[13]), .B(a[13]), .Z(n1840) );
  OR U2301 ( .A(n1840), .B(n1681), .Z(n1682) );
  NAND U2302 ( .A(n1683), .B(n1682), .Z(n1784) );
  XOR U2303 ( .A(n1783), .B(n1784), .Z(n1786) );
  XOR U2304 ( .A(n1785), .B(n1786), .Z(n1778) );
  OR U2305 ( .A(n1684), .B(n180), .Z(n1686) );
  XOR U2306 ( .A(b[3]), .B(a[23]), .Z(n1837) );
  NAND U2307 ( .A(n182), .B(n1837), .Z(n1685) );
  AND U2308 ( .A(n1686), .B(n1685), .Z(n1802) );
  NAND U2309 ( .A(n188), .B(n1687), .Z(n1689) );
  XOR U2310 ( .A(b[15]), .B(a[11]), .Z(n1834) );
  NAND U2311 ( .A(n37382), .B(n1834), .Z(n1688) );
  AND U2312 ( .A(n1689), .B(n1688), .Z(n1800) );
  NAND U2313 ( .A(b[23]), .B(b[24]), .Z(n1690) );
  AND U2314 ( .A(b[25]), .B(n1690), .Z(n38352) );
  IV U2315 ( .A(n38352), .Z(n38379) );
  NOR U2316 ( .A(n38379), .B(n1691), .Z(n1799) );
  XNOR U2317 ( .A(n1800), .B(n1799), .Z(n1801) );
  XNOR U2318 ( .A(n1802), .B(n1801), .Z(n1777) );
  XOR U2319 ( .A(n1778), .B(n1777), .Z(n1780) );
  XOR U2320 ( .A(n1779), .B(n1780), .Z(n1773) );
  NANDN U2321 ( .A(n1693), .B(n1692), .Z(n1697) );
  NANDN U2322 ( .A(n1695), .B(n1694), .Z(n1696) );
  AND U2323 ( .A(n1697), .B(n1696), .Z(n1772) );
  NANDN U2324 ( .A(n1699), .B(n1698), .Z(n1703) );
  NANDN U2325 ( .A(n1701), .B(n1700), .Z(n1702) );
  AND U2326 ( .A(n1703), .B(n1702), .Z(n1771) );
  XOR U2327 ( .A(n1772), .B(n1771), .Z(n1774) );
  XNOR U2328 ( .A(n1773), .B(n1774), .Z(n1855) );
  XNOR U2329 ( .A(n1856), .B(n1855), .Z(n1857) );
  NANDN U2330 ( .A(n1705), .B(n1704), .Z(n1709) );
  NANDN U2331 ( .A(n1707), .B(n1706), .Z(n1708) );
  AND U2332 ( .A(n1709), .B(n1708), .Z(n1768) );
  NANDN U2333 ( .A(n1711), .B(n1710), .Z(n1715) );
  NANDN U2334 ( .A(n1713), .B(n1712), .Z(n1714) );
  AND U2335 ( .A(n1715), .B(n1714), .Z(n1766) );
  NAND U2336 ( .A(n184), .B(n1716), .Z(n1718) );
  XOR U2337 ( .A(b[7]), .B(a[19]), .Z(n1811) );
  NAND U2338 ( .A(n36592), .B(n1811), .Z(n1717) );
  AND U2339 ( .A(n1718), .B(n1717), .Z(n1828) );
  NAND U2340 ( .A(n183), .B(n1719), .Z(n1721) );
  XOR U2341 ( .A(b[5]), .B(a[21]), .Z(n1846) );
  NAND U2342 ( .A(n36296), .B(n1846), .Z(n1720) );
  AND U2343 ( .A(n1721), .B(n1720), .Z(n1827) );
  NAND U2344 ( .A(n189), .B(n1722), .Z(n1724) );
  XOR U2345 ( .A(b[17]), .B(a[9]), .Z(n1796) );
  NAND U2346 ( .A(n37652), .B(n1796), .Z(n1723) );
  NAND U2347 ( .A(n1724), .B(n1723), .Z(n1826) );
  XOR U2348 ( .A(n1827), .B(n1826), .Z(n1829) );
  XOR U2349 ( .A(n1828), .B(n1829), .Z(n1851) );
  NAND U2350 ( .A(n190), .B(n1725), .Z(n1727) );
  XOR U2351 ( .A(b[19]), .B(a[7]), .Z(n1843) );
  NAND U2352 ( .A(n37821), .B(n1843), .Z(n1726) );
  AND U2353 ( .A(n1727), .B(n1726), .Z(n1822) );
  NAND U2354 ( .A(n38064), .B(n1728), .Z(n1730) );
  XOR U2355 ( .A(b[21]), .B(a[5]), .Z(n1789) );
  NAND U2356 ( .A(n37993), .B(n1789), .Z(n1729) );
  AND U2357 ( .A(n1730), .B(n1729), .Z(n1821) );
  NAND U2358 ( .A(n185), .B(n1731), .Z(n1733) );
  XOR U2359 ( .A(b[9]), .B(a[17]), .Z(n1805) );
  NAND U2360 ( .A(n36805), .B(n1805), .Z(n1732) );
  NAND U2361 ( .A(n1733), .B(n1732), .Z(n1820) );
  XOR U2362 ( .A(n1821), .B(n1820), .Z(n1823) );
  XOR U2363 ( .A(n1822), .B(n1823), .Z(n1850) );
  NANDN U2364 ( .A(n176), .B(n1734), .Z(n1736) );
  XNOR U2365 ( .A(b[11]), .B(a[15]), .Z(n1808) );
  OR U2366 ( .A(n1808), .B(n2434), .Z(n1735) );
  AND U2367 ( .A(n1736), .B(n1735), .Z(n1849) );
  XOR U2368 ( .A(n1850), .B(n1849), .Z(n1852) );
  XNOR U2369 ( .A(n1851), .B(n1852), .Z(n1765) );
  XNOR U2370 ( .A(n1766), .B(n1765), .Z(n1767) );
  XOR U2371 ( .A(n1768), .B(n1767), .Z(n1858) );
  XNOR U2372 ( .A(n1857), .B(n1858), .Z(n1863) );
  XOR U2373 ( .A(n1864), .B(n1863), .Z(n1760) );
  NANDN U2374 ( .A(n1738), .B(n1737), .Z(n1742) );
  OR U2375 ( .A(n1740), .B(n1739), .Z(n1741) );
  AND U2376 ( .A(n1742), .B(n1741), .Z(n1759) );
  XNOR U2377 ( .A(n1760), .B(n1759), .Z(n1761) );
  XNOR U2378 ( .A(n1762), .B(n1761), .Z(n1753) );
  XNOR U2379 ( .A(n1754), .B(n1753), .Z(n1755) );
  XNOR U2380 ( .A(n1756), .B(n1755), .Z(n1748) );
  XNOR U2381 ( .A(sreg[249]), .B(n1748), .Z(n1750) );
  NANDN U2382 ( .A(sreg[248]), .B(n1743), .Z(n1747) );
  NAND U2383 ( .A(n1745), .B(n1744), .Z(n1746) );
  NAND U2384 ( .A(n1747), .B(n1746), .Z(n1749) );
  XNOR U2385 ( .A(n1750), .B(n1749), .Z(c[249]) );
  NANDN U2386 ( .A(sreg[249]), .B(n1748), .Z(n1752) );
  NAND U2387 ( .A(n1750), .B(n1749), .Z(n1751) );
  NAND U2388 ( .A(n1752), .B(n1751), .Z(n1987) );
  XNOR U2389 ( .A(sreg[250]), .B(n1987), .Z(n1989) );
  NANDN U2390 ( .A(n1754), .B(n1753), .Z(n1758) );
  NANDN U2391 ( .A(n1756), .B(n1755), .Z(n1757) );
  AND U2392 ( .A(n1758), .B(n1757), .Z(n1870) );
  NANDN U2393 ( .A(n1760), .B(n1759), .Z(n1764) );
  NANDN U2394 ( .A(n1762), .B(n1761), .Z(n1763) );
  AND U2395 ( .A(n1764), .B(n1763), .Z(n1868) );
  NANDN U2396 ( .A(n1766), .B(n1765), .Z(n1770) );
  NANDN U2397 ( .A(n1768), .B(n1767), .Z(n1769) );
  AND U2398 ( .A(n1770), .B(n1769), .Z(n1880) );
  NANDN U2399 ( .A(n1772), .B(n1771), .Z(n1776) );
  OR U2400 ( .A(n1774), .B(n1773), .Z(n1775) );
  AND U2401 ( .A(n1776), .B(n1775), .Z(n1879) );
  XNOR U2402 ( .A(n1880), .B(n1879), .Z(n1882) );
  NANDN U2403 ( .A(n1778), .B(n1777), .Z(n1782) );
  OR U2404 ( .A(n1780), .B(n1779), .Z(n1781) );
  AND U2405 ( .A(n1782), .B(n1781), .Z(n1892) );
  NANDN U2406 ( .A(n1784), .B(n1783), .Z(n1788) );
  OR U2407 ( .A(n1786), .B(n1785), .Z(n1787) );
  AND U2408 ( .A(n1788), .B(n1787), .Z(n1970) );
  NAND U2409 ( .A(n38064), .B(n1789), .Z(n1791) );
  XOR U2410 ( .A(b[21]), .B(a[6]), .Z(n1954) );
  NAND U2411 ( .A(n37993), .B(n1954), .Z(n1790) );
  AND U2412 ( .A(n1791), .B(n1790), .Z(n1925) );
  AND U2413 ( .A(n1792), .B(n37513), .Z(n38289) );
  NAND U2414 ( .A(n38289), .B(n1793), .Z(n1795) );
  XOR U2415 ( .A(b[25]), .B(a[2]), .Z(n1905) );
  NAND U2416 ( .A(n38247), .B(n1905), .Z(n1794) );
  AND U2417 ( .A(n1795), .B(n1794), .Z(n1924) );
  NAND U2418 ( .A(n189), .B(n1796), .Z(n1798) );
  XOR U2419 ( .A(b[17]), .B(a[10]), .Z(n1951) );
  NAND U2420 ( .A(n37652), .B(n1951), .Z(n1797) );
  NAND U2421 ( .A(n1798), .B(n1797), .Z(n1923) );
  XOR U2422 ( .A(n1924), .B(n1923), .Z(n1926) );
  XNOR U2423 ( .A(n1925), .B(n1926), .Z(n1969) );
  XNOR U2424 ( .A(n1970), .B(n1969), .Z(n1972) );
  NANDN U2425 ( .A(n1800), .B(n1799), .Z(n1804) );
  NANDN U2426 ( .A(n1802), .B(n1801), .Z(n1803) );
  AND U2427 ( .A(n1804), .B(n1803), .Z(n1971) );
  XNOR U2428 ( .A(n1972), .B(n1971), .Z(n1891) );
  XNOR U2429 ( .A(n1892), .B(n1891), .Z(n1894) );
  NAND U2430 ( .A(n185), .B(n1805), .Z(n1807) );
  XOR U2431 ( .A(b[9]), .B(a[18]), .Z(n1960) );
  NAND U2432 ( .A(n36805), .B(n1960), .Z(n1806) );
  AND U2433 ( .A(n1807), .B(n1806), .Z(n1931) );
  OR U2434 ( .A(n1808), .B(n176), .Z(n1810) );
  XOR U2435 ( .A(b[11]), .B(a[16]), .Z(n1948) );
  NAND U2436 ( .A(n37097), .B(n1948), .Z(n1809) );
  AND U2437 ( .A(n1810), .B(n1809), .Z(n1930) );
  NAND U2438 ( .A(n184), .B(n1811), .Z(n1813) );
  XOR U2439 ( .A(b[7]), .B(a[20]), .Z(n1908) );
  NAND U2440 ( .A(n36592), .B(n1908), .Z(n1812) );
  NAND U2441 ( .A(n1813), .B(n1812), .Z(n1929) );
  XOR U2442 ( .A(n1930), .B(n1929), .Z(n1932) );
  XOR U2443 ( .A(n1931), .B(n1932), .Z(n1976) );
  NAND U2444 ( .A(b[0]), .B(a[26]), .Z(n1814) );
  XNOR U2445 ( .A(b[1]), .B(n1814), .Z(n1816) );
  NANDN U2446 ( .A(b[0]), .B(a[25]), .Z(n1815) );
  NAND U2447 ( .A(n1816), .B(n1815), .Z(n1937) );
  XNOR U2448 ( .A(b[25]), .B(b[26]), .Z(n2105) );
  IV U2449 ( .A(n2105), .Z(n38343) );
  AND U2450 ( .A(a[0]), .B(n38343), .Z(n1947) );
  NAND U2451 ( .A(n38185), .B(n1817), .Z(n1819) );
  XOR U2452 ( .A(b[23]), .B(a[4]), .Z(n1957) );
  NAND U2453 ( .A(n38132), .B(n1957), .Z(n1818) );
  AND U2454 ( .A(n1819), .B(n1818), .Z(n1935) );
  XOR U2455 ( .A(n1947), .B(n1935), .Z(n1936) );
  XNOR U2456 ( .A(n1937), .B(n1936), .Z(n1975) );
  XNOR U2457 ( .A(n1976), .B(n1975), .Z(n1977) );
  NANDN U2458 ( .A(n1821), .B(n1820), .Z(n1825) );
  OR U2459 ( .A(n1823), .B(n1822), .Z(n1824) );
  NAND U2460 ( .A(n1825), .B(n1824), .Z(n1978) );
  XOR U2461 ( .A(n1977), .B(n1978), .Z(n1885) );
  NANDN U2462 ( .A(n1827), .B(n1826), .Z(n1831) );
  OR U2463 ( .A(n1829), .B(n1828), .Z(n1830) );
  AND U2464 ( .A(n1831), .B(n1830), .Z(n1984) );
  NOR U2465 ( .A(n1833), .B(n1832), .Z(n1919) );
  NANDN U2466 ( .A(n178), .B(n1834), .Z(n1836) );
  XNOR U2467 ( .A(b[15]), .B(a[12]), .Z(n1943) );
  OR U2468 ( .A(n1943), .B(n37509), .Z(n1835) );
  AND U2469 ( .A(n1836), .B(n1835), .Z(n1917) );
  NANDN U2470 ( .A(n180), .B(n1837), .Z(n1839) );
  XNOR U2471 ( .A(b[3]), .B(a[24]), .Z(n1940) );
  OR U2472 ( .A(n1940), .B(n172), .Z(n1838) );
  NAND U2473 ( .A(n1839), .B(n1838), .Z(n1918) );
  XOR U2474 ( .A(n1917), .B(n1918), .Z(n1920) );
  XOR U2475 ( .A(n1919), .B(n1920), .Z(n1982) );
  OR U2476 ( .A(n1840), .B(n171), .Z(n1842) );
  XOR U2477 ( .A(b[13]), .B(a[14]), .Z(n1898) );
  NAND U2478 ( .A(n37295), .B(n1898), .Z(n1841) );
  AND U2479 ( .A(n1842), .B(n1841), .Z(n1966) );
  NAND U2480 ( .A(n190), .B(n1843), .Z(n1845) );
  XOR U2481 ( .A(b[19]), .B(a[8]), .Z(n1914) );
  NAND U2482 ( .A(n37821), .B(n1914), .Z(n1844) );
  AND U2483 ( .A(n1845), .B(n1844), .Z(n1964) );
  NAND U2484 ( .A(n183), .B(n1846), .Z(n1848) );
  XOR U2485 ( .A(b[5]), .B(a[22]), .Z(n1911) );
  NAND U2486 ( .A(n36296), .B(n1911), .Z(n1847) );
  NAND U2487 ( .A(n1848), .B(n1847), .Z(n1963) );
  XNOR U2488 ( .A(n1964), .B(n1963), .Z(n1965) );
  XNOR U2489 ( .A(n1966), .B(n1965), .Z(n1981) );
  XNOR U2490 ( .A(n1982), .B(n1981), .Z(n1983) );
  XNOR U2491 ( .A(n1984), .B(n1983), .Z(n1886) );
  XOR U2492 ( .A(n1885), .B(n1886), .Z(n1888) );
  NANDN U2493 ( .A(n1850), .B(n1849), .Z(n1854) );
  OR U2494 ( .A(n1852), .B(n1851), .Z(n1853) );
  AND U2495 ( .A(n1854), .B(n1853), .Z(n1887) );
  XNOR U2496 ( .A(n1888), .B(n1887), .Z(n1893) );
  XNOR U2497 ( .A(n1894), .B(n1893), .Z(n1881) );
  XOR U2498 ( .A(n1882), .B(n1881), .Z(n1876) );
  NANDN U2499 ( .A(n1856), .B(n1855), .Z(n1860) );
  NANDN U2500 ( .A(n1858), .B(n1857), .Z(n1859) );
  AND U2501 ( .A(n1860), .B(n1859), .Z(n1873) );
  NANDN U2502 ( .A(n1862), .B(n1861), .Z(n1866) );
  NAND U2503 ( .A(n1864), .B(n1863), .Z(n1865) );
  NAND U2504 ( .A(n1866), .B(n1865), .Z(n1874) );
  XNOR U2505 ( .A(n1873), .B(n1874), .Z(n1875) );
  XNOR U2506 ( .A(n1876), .B(n1875), .Z(n1867) );
  XNOR U2507 ( .A(n1868), .B(n1867), .Z(n1869) );
  XNOR U2508 ( .A(n1870), .B(n1869), .Z(n1988) );
  XNOR U2509 ( .A(n1989), .B(n1988), .Z(c[250]) );
  NANDN U2510 ( .A(n1868), .B(n1867), .Z(n1872) );
  NANDN U2511 ( .A(n1870), .B(n1869), .Z(n1871) );
  AND U2512 ( .A(n1872), .B(n1871), .Z(n2000) );
  NANDN U2513 ( .A(n1874), .B(n1873), .Z(n1878) );
  NANDN U2514 ( .A(n1876), .B(n1875), .Z(n1877) );
  AND U2515 ( .A(n1878), .B(n1877), .Z(n1998) );
  NANDN U2516 ( .A(n1880), .B(n1879), .Z(n1884) );
  NAND U2517 ( .A(n1882), .B(n1881), .Z(n1883) );
  AND U2518 ( .A(n1884), .B(n1883), .Z(n2005) );
  NAND U2519 ( .A(n1886), .B(n1885), .Z(n1890) );
  NAND U2520 ( .A(n1888), .B(n1887), .Z(n1889) );
  AND U2521 ( .A(n1890), .B(n1889), .Z(n2003) );
  NAND U2522 ( .A(b[0]), .B(a[27]), .Z(n1895) );
  XNOR U2523 ( .A(b[1]), .B(n1895), .Z(n1897) );
  NANDN U2524 ( .A(b[0]), .B(a[26]), .Z(n1896) );
  NAND U2525 ( .A(n1897), .B(n1896), .Z(n2065) );
  NAND U2526 ( .A(n187), .B(n1898), .Z(n1900) );
  XOR U2527 ( .A(b[13]), .B(a[15]), .Z(n2061) );
  NAND U2528 ( .A(n37295), .B(n2061), .Z(n1899) );
  NAND U2529 ( .A(n1900), .B(n1899), .Z(n2064) );
  XNOR U2530 ( .A(n2065), .B(n2064), .Z(n2066) );
  XOR U2531 ( .A(b[27]), .B(b[26]), .Z(n2103) );
  XOR U2532 ( .A(b[27]), .B(a[0]), .Z(n1901) );
  NAND U2533 ( .A(n2103), .B(n1901), .Z(n1902) );
  NANDN U2534 ( .A(n1902), .B(n2105), .Z(n1904) );
  XOR U2535 ( .A(b[27]), .B(a[1]), .Z(n2104) );
  NANDN U2536 ( .A(n2105), .B(n2104), .Z(n1903) );
  AND U2537 ( .A(n1904), .B(n1903), .Z(n2098) );
  NAND U2538 ( .A(n38289), .B(n1905), .Z(n1907) );
  XOR U2539 ( .A(b[25]), .B(a[3]), .Z(n2095) );
  NAND U2540 ( .A(n38247), .B(n2095), .Z(n1906) );
  NAND U2541 ( .A(n1907), .B(n1906), .Z(n2099) );
  XOR U2542 ( .A(n2098), .B(n2099), .Z(n2067) );
  XNOR U2543 ( .A(n2066), .B(n2067), .Z(n2027) );
  NAND U2544 ( .A(n184), .B(n1908), .Z(n1910) );
  XOR U2545 ( .A(b[7]), .B(a[21]), .Z(n2048) );
  NAND U2546 ( .A(n36592), .B(n2048), .Z(n1909) );
  AND U2547 ( .A(n1910), .B(n1909), .Z(n2111) );
  NAND U2548 ( .A(n183), .B(n1911), .Z(n1913) );
  XOR U2549 ( .A(b[5]), .B(a[23]), .Z(n2039) );
  NAND U2550 ( .A(n36296), .B(n2039), .Z(n1912) );
  AND U2551 ( .A(n1913), .B(n1912), .Z(n2109) );
  NAND U2552 ( .A(n190), .B(n1914), .Z(n1916) );
  XOR U2553 ( .A(b[19]), .B(a[9]), .Z(n2033) );
  NAND U2554 ( .A(n37821), .B(n2033), .Z(n1915) );
  NAND U2555 ( .A(n1916), .B(n1915), .Z(n2108) );
  XNOR U2556 ( .A(n2109), .B(n2108), .Z(n2110) );
  XOR U2557 ( .A(n2111), .B(n2110), .Z(n2028) );
  XNOR U2558 ( .A(n2027), .B(n2028), .Z(n2029) );
  NANDN U2559 ( .A(n1918), .B(n1917), .Z(n1922) );
  OR U2560 ( .A(n1920), .B(n1919), .Z(n1921) );
  NAND U2561 ( .A(n1922), .B(n1921), .Z(n2030) );
  XNOR U2562 ( .A(n2029), .B(n2030), .Z(n2018) );
  NANDN U2563 ( .A(n1924), .B(n1923), .Z(n1928) );
  OR U2564 ( .A(n1926), .B(n1925), .Z(n1927) );
  NAND U2565 ( .A(n1928), .B(n1927), .Z(n2016) );
  NANDN U2566 ( .A(n1930), .B(n1929), .Z(n1934) );
  OR U2567 ( .A(n1932), .B(n1931), .Z(n1933) );
  NAND U2568 ( .A(n1934), .B(n1933), .Z(n2015) );
  XOR U2569 ( .A(n2016), .B(n2015), .Z(n2017) );
  XOR U2570 ( .A(n2018), .B(n2017), .Z(n2024) );
  NANDN U2571 ( .A(n1935), .B(n1947), .Z(n1939) );
  OR U2572 ( .A(n1937), .B(n1936), .Z(n1938) );
  AND U2573 ( .A(n1939), .B(n1938), .Z(n2077) );
  OR U2574 ( .A(n1940), .B(n180), .Z(n1942) );
  XOR U2575 ( .A(b[3]), .B(a[25]), .Z(n2055) );
  NAND U2576 ( .A(n182), .B(n2055), .Z(n1941) );
  AND U2577 ( .A(n1942), .B(n1941), .Z(n2089) );
  OR U2578 ( .A(n1943), .B(n178), .Z(n1945) );
  XOR U2579 ( .A(b[15]), .B(a[13]), .Z(n2100) );
  NAND U2580 ( .A(n37382), .B(n2100), .Z(n1944) );
  NAND U2581 ( .A(n1945), .B(n1944), .Z(n2088) );
  XNOR U2582 ( .A(n2089), .B(n2088), .Z(n2091) );
  NAND U2583 ( .A(b[25]), .B(b[26]), .Z(n1946) );
  NAND U2584 ( .A(b[27]), .B(n1946), .Z(n38448) );
  OR U2585 ( .A(n38448), .B(n1947), .Z(n2090) );
  XNOR U2586 ( .A(n2091), .B(n2090), .Z(n2076) );
  XNOR U2587 ( .A(n2077), .B(n2076), .Z(n2079) );
  NAND U2588 ( .A(n186), .B(n1948), .Z(n1950) );
  XOR U2589 ( .A(b[11]), .B(a[17]), .Z(n2042) );
  NAND U2590 ( .A(n37097), .B(n2042), .Z(n1949) );
  AND U2591 ( .A(n1950), .B(n1949), .Z(n2083) );
  NAND U2592 ( .A(n189), .B(n1951), .Z(n1953) );
  XOR U2593 ( .A(b[17]), .B(a[11]), .Z(n2045) );
  NAND U2594 ( .A(n37652), .B(n2045), .Z(n1952) );
  NAND U2595 ( .A(n1953), .B(n1952), .Z(n2082) );
  XNOR U2596 ( .A(n2083), .B(n2082), .Z(n2084) );
  NAND U2597 ( .A(n38064), .B(n1954), .Z(n1956) );
  XOR U2598 ( .A(b[21]), .B(a[7]), .Z(n2036) );
  NAND U2599 ( .A(n37993), .B(n2036), .Z(n1955) );
  AND U2600 ( .A(n1956), .B(n1955), .Z(n2073) );
  NAND U2601 ( .A(n38185), .B(n1957), .Z(n1959) );
  XOR U2602 ( .A(b[23]), .B(a[5]), .Z(n2058) );
  NAND U2603 ( .A(n38132), .B(n2058), .Z(n1958) );
  AND U2604 ( .A(n1959), .B(n1958), .Z(n2071) );
  NAND U2605 ( .A(n185), .B(n1960), .Z(n1962) );
  XOR U2606 ( .A(b[9]), .B(a[19]), .Z(n2051) );
  NAND U2607 ( .A(n36805), .B(n2051), .Z(n1961) );
  NAND U2608 ( .A(n1962), .B(n1961), .Z(n2070) );
  XNOR U2609 ( .A(n2071), .B(n2070), .Z(n2072) );
  XOR U2610 ( .A(n2073), .B(n2072), .Z(n2085) );
  XNOR U2611 ( .A(n2084), .B(n2085), .Z(n2078) );
  XOR U2612 ( .A(n2079), .B(n2078), .Z(n2022) );
  NANDN U2613 ( .A(n1964), .B(n1963), .Z(n1968) );
  NANDN U2614 ( .A(n1966), .B(n1965), .Z(n1967) );
  AND U2615 ( .A(n1968), .B(n1967), .Z(n2021) );
  XNOR U2616 ( .A(n2022), .B(n2021), .Z(n2023) );
  XNOR U2617 ( .A(n2024), .B(n2023), .Z(n2114) );
  NANDN U2618 ( .A(n1970), .B(n1969), .Z(n1974) );
  NAND U2619 ( .A(n1972), .B(n1971), .Z(n1973) );
  AND U2620 ( .A(n1974), .B(n1973), .Z(n2012) );
  NANDN U2621 ( .A(n1976), .B(n1975), .Z(n1980) );
  NANDN U2622 ( .A(n1978), .B(n1977), .Z(n1979) );
  AND U2623 ( .A(n1980), .B(n1979), .Z(n2010) );
  NANDN U2624 ( .A(n1982), .B(n1981), .Z(n1986) );
  NANDN U2625 ( .A(n1984), .B(n1983), .Z(n1985) );
  AND U2626 ( .A(n1986), .B(n1985), .Z(n2009) );
  XNOR U2627 ( .A(n2010), .B(n2009), .Z(n2011) );
  XOR U2628 ( .A(n2012), .B(n2011), .Z(n2115) );
  XOR U2629 ( .A(n2114), .B(n2115), .Z(n2117) );
  XOR U2630 ( .A(n2116), .B(n2117), .Z(n2004) );
  XOR U2631 ( .A(n2003), .B(n2004), .Z(n2006) );
  XNOR U2632 ( .A(n2005), .B(n2006), .Z(n1997) );
  XNOR U2633 ( .A(n1998), .B(n1997), .Z(n1999) );
  XNOR U2634 ( .A(n2000), .B(n1999), .Z(n1992) );
  XNOR U2635 ( .A(sreg[251]), .B(n1992), .Z(n1994) );
  NANDN U2636 ( .A(sreg[250]), .B(n1987), .Z(n1991) );
  NAND U2637 ( .A(n1989), .B(n1988), .Z(n1990) );
  NAND U2638 ( .A(n1991), .B(n1990), .Z(n1993) );
  XNOR U2639 ( .A(n1994), .B(n1993), .Z(c[251]) );
  NANDN U2640 ( .A(sreg[251]), .B(n1992), .Z(n1996) );
  NAND U2641 ( .A(n1994), .B(n1993), .Z(n1995) );
  NAND U2642 ( .A(n1996), .B(n1995), .Z(n2251) );
  XNOR U2643 ( .A(sreg[252]), .B(n2251), .Z(n2253) );
  NANDN U2644 ( .A(n1998), .B(n1997), .Z(n2002) );
  NANDN U2645 ( .A(n2000), .B(n1999), .Z(n2001) );
  AND U2646 ( .A(n2002), .B(n2001), .Z(n2123) );
  NANDN U2647 ( .A(n2004), .B(n2003), .Z(n2008) );
  NANDN U2648 ( .A(n2006), .B(n2005), .Z(n2007) );
  AND U2649 ( .A(n2008), .B(n2007), .Z(n2121) );
  NANDN U2650 ( .A(n2010), .B(n2009), .Z(n2014) );
  NANDN U2651 ( .A(n2012), .B(n2011), .Z(n2013) );
  AND U2652 ( .A(n2014), .B(n2013), .Z(n2129) );
  NAND U2653 ( .A(n2016), .B(n2015), .Z(n2020) );
  NAND U2654 ( .A(n2018), .B(n2017), .Z(n2019) );
  AND U2655 ( .A(n2020), .B(n2019), .Z(n2127) );
  NANDN U2656 ( .A(n2022), .B(n2021), .Z(n2026) );
  NANDN U2657 ( .A(n2024), .B(n2023), .Z(n2025) );
  AND U2658 ( .A(n2026), .B(n2025), .Z(n2126) );
  XNOR U2659 ( .A(n2127), .B(n2126), .Z(n2128) );
  XOR U2660 ( .A(n2129), .B(n2128), .Z(n2248) );
  NANDN U2661 ( .A(n2028), .B(n2027), .Z(n2032) );
  NANDN U2662 ( .A(n2030), .B(n2029), .Z(n2031) );
  AND U2663 ( .A(n2032), .B(n2031), .Z(n2218) );
  NAND U2664 ( .A(n190), .B(n2033), .Z(n2035) );
  XOR U2665 ( .A(b[19]), .B(a[10]), .Z(n2148) );
  NAND U2666 ( .A(n37821), .B(n2148), .Z(n2034) );
  AND U2667 ( .A(n2035), .B(n2034), .Z(n2168) );
  NAND U2668 ( .A(n38064), .B(n2036), .Z(n2038) );
  XOR U2669 ( .A(b[21]), .B(a[8]), .Z(n2175) );
  NAND U2670 ( .A(n37993), .B(n2175), .Z(n2037) );
  AND U2671 ( .A(n2038), .B(n2037), .Z(n2167) );
  NAND U2672 ( .A(n183), .B(n2039), .Z(n2041) );
  XOR U2673 ( .A(b[5]), .B(a[24]), .Z(n2179) );
  NAND U2674 ( .A(n36296), .B(n2179), .Z(n2040) );
  NAND U2675 ( .A(n2041), .B(n2040), .Z(n2166) );
  XOR U2676 ( .A(n2167), .B(n2166), .Z(n2169) );
  XOR U2677 ( .A(n2168), .B(n2169), .Z(n2236) );
  NAND U2678 ( .A(n186), .B(n2042), .Z(n2044) );
  XOR U2679 ( .A(b[11]), .B(a[18]), .Z(n2151) );
  NAND U2680 ( .A(n37097), .B(n2151), .Z(n2043) );
  AND U2681 ( .A(n2044), .B(n2043), .Z(n2205) );
  NAND U2682 ( .A(n189), .B(n2045), .Z(n2047) );
  XOR U2683 ( .A(b[17]), .B(a[12]), .Z(n2185) );
  NAND U2684 ( .A(n37652), .B(n2185), .Z(n2046) );
  AND U2685 ( .A(n2047), .B(n2046), .Z(n2204) );
  NAND U2686 ( .A(n184), .B(n2048), .Z(n2050) );
  XOR U2687 ( .A(b[7]), .B(a[22]), .Z(n2172) );
  NAND U2688 ( .A(n36592), .B(n2172), .Z(n2049) );
  NAND U2689 ( .A(n2050), .B(n2049), .Z(n2203) );
  XOR U2690 ( .A(n2204), .B(n2203), .Z(n2206) );
  XOR U2691 ( .A(n2205), .B(n2206), .Z(n2234) );
  NANDN U2692 ( .A(n179), .B(n2051), .Z(n2054) );
  XNOR U2693 ( .A(b[9]), .B(a[20]), .Z(n2194) );
  OR U2694 ( .A(n2194), .B(n2052), .Z(n2053) );
  AND U2695 ( .A(n2054), .B(n2053), .Z(n2233) );
  XNOR U2696 ( .A(n2234), .B(n2233), .Z(n2235) );
  XNOR U2697 ( .A(n2236), .B(n2235), .Z(n2215) );
  NAND U2698 ( .A(n181), .B(n2055), .Z(n2057) );
  XOR U2699 ( .A(b[3]), .B(a[26]), .Z(n2182) );
  NAND U2700 ( .A(n182), .B(n2182), .Z(n2056) );
  AND U2701 ( .A(n2057), .B(n2056), .Z(n2162) );
  NAND U2702 ( .A(n38185), .B(n2058), .Z(n2060) );
  XOR U2703 ( .A(b[23]), .B(a[6]), .Z(n2188) );
  NAND U2704 ( .A(n38132), .B(n2188), .Z(n2059) );
  AND U2705 ( .A(n2060), .B(n2059), .Z(n2161) );
  NAND U2706 ( .A(n187), .B(n2061), .Z(n2063) );
  XOR U2707 ( .A(b[13]), .B(a[16]), .Z(n2145) );
  NAND U2708 ( .A(n37295), .B(n2145), .Z(n2062) );
  NAND U2709 ( .A(n2063), .B(n2062), .Z(n2160) );
  XOR U2710 ( .A(n2161), .B(n2160), .Z(n2163) );
  XOR U2711 ( .A(n2162), .B(n2163), .Z(n2222) );
  NANDN U2712 ( .A(n2065), .B(n2064), .Z(n2069) );
  NANDN U2713 ( .A(n2067), .B(n2066), .Z(n2068) );
  AND U2714 ( .A(n2069), .B(n2068), .Z(n2221) );
  XNOR U2715 ( .A(n2222), .B(n2221), .Z(n2223) );
  NANDN U2716 ( .A(n2071), .B(n2070), .Z(n2075) );
  NANDN U2717 ( .A(n2073), .B(n2072), .Z(n2074) );
  NAND U2718 ( .A(n2075), .B(n2074), .Z(n2224) );
  XOR U2719 ( .A(n2223), .B(n2224), .Z(n2216) );
  XNOR U2720 ( .A(n2215), .B(n2216), .Z(n2217) );
  XOR U2721 ( .A(n2218), .B(n2217), .Z(n2241) );
  NANDN U2722 ( .A(n2077), .B(n2076), .Z(n2081) );
  NAND U2723 ( .A(n2079), .B(n2078), .Z(n2080) );
  AND U2724 ( .A(n2081), .B(n2080), .Z(n2240) );
  NANDN U2725 ( .A(n2083), .B(n2082), .Z(n2087) );
  NANDN U2726 ( .A(n2085), .B(n2084), .Z(n2086) );
  AND U2727 ( .A(n2087), .B(n2086), .Z(n2212) );
  NAND U2728 ( .A(b[0]), .B(a[28]), .Z(n2092) );
  XNOR U2729 ( .A(b[1]), .B(n2092), .Z(n2094) );
  NANDN U2730 ( .A(b[0]), .B(a[27]), .Z(n2093) );
  NAND U2731 ( .A(n2094), .B(n2093), .Z(n2200) );
  XOR U2732 ( .A(b[27]), .B(b[28]), .Z(n38456) );
  AND U2733 ( .A(a[0]), .B(n38456), .Z(n2197) );
  NAND U2734 ( .A(n38289), .B(n2095), .Z(n2097) );
  XOR U2735 ( .A(b[25]), .B(a[4]), .Z(n2191) );
  NAND U2736 ( .A(n38247), .B(n2191), .Z(n2096) );
  AND U2737 ( .A(n2097), .B(n2096), .Z(n2198) );
  XOR U2738 ( .A(n2197), .B(n2198), .Z(n2199) );
  XOR U2739 ( .A(n2200), .B(n2199), .Z(n2228) );
  ANDN U2740 ( .B(n2099), .A(n2098), .Z(n2157) );
  NANDN U2741 ( .A(n178), .B(n2100), .Z(n2102) );
  XNOR U2742 ( .A(b[15]), .B(a[14]), .Z(n2142) );
  OR U2743 ( .A(n2142), .B(n37509), .Z(n2101) );
  AND U2744 ( .A(n2102), .B(n2101), .Z(n2154) );
  AND U2745 ( .A(n2103), .B(n2105), .Z(n38385) );
  NANDN U2746 ( .A(n192), .B(n2104), .Z(n2107) );
  XNOR U2747 ( .A(b[27]), .B(a[2]), .Z(n2136) );
  OR U2748 ( .A(n2136), .B(n2105), .Z(n2106) );
  NAND U2749 ( .A(n2107), .B(n2106), .Z(n2155) );
  XNOR U2750 ( .A(n2154), .B(n2155), .Z(n2156) );
  XNOR U2751 ( .A(n2157), .B(n2156), .Z(n2227) );
  XNOR U2752 ( .A(n2228), .B(n2227), .Z(n2230) );
  NANDN U2753 ( .A(n2109), .B(n2108), .Z(n2113) );
  NANDN U2754 ( .A(n2111), .B(n2110), .Z(n2112) );
  AND U2755 ( .A(n2113), .B(n2112), .Z(n2229) );
  XNOR U2756 ( .A(n2230), .B(n2229), .Z(n2209) );
  XNOR U2757 ( .A(n2210), .B(n2209), .Z(n2211) );
  XNOR U2758 ( .A(n2212), .B(n2211), .Z(n2239) );
  XOR U2759 ( .A(n2240), .B(n2239), .Z(n2242) );
  XOR U2760 ( .A(n2241), .B(n2242), .Z(n2246) );
  NANDN U2761 ( .A(n2115), .B(n2114), .Z(n2119) );
  NANDN U2762 ( .A(n2117), .B(n2116), .Z(n2118) );
  NAND U2763 ( .A(n2119), .B(n2118), .Z(n2245) );
  XNOR U2764 ( .A(n2246), .B(n2245), .Z(n2247) );
  XNOR U2765 ( .A(n2248), .B(n2247), .Z(n2120) );
  XNOR U2766 ( .A(n2121), .B(n2120), .Z(n2122) );
  XNOR U2767 ( .A(n2123), .B(n2122), .Z(n2252) );
  XNOR U2768 ( .A(n2253), .B(n2252), .Z(c[252]) );
  NANDN U2769 ( .A(n2121), .B(n2120), .Z(n2125) );
  NANDN U2770 ( .A(n2123), .B(n2122), .Z(n2124) );
  AND U2771 ( .A(n2125), .B(n2124), .Z(n2264) );
  NANDN U2772 ( .A(n2127), .B(n2126), .Z(n2131) );
  NAND U2773 ( .A(n2129), .B(n2128), .Z(n2130) );
  AND U2774 ( .A(n2131), .B(n2130), .Z(n2387) );
  XOR U2775 ( .A(b[29]), .B(b[28]), .Z(n2336) );
  XOR U2776 ( .A(b[29]), .B(a[0]), .Z(n2132) );
  NAND U2777 ( .A(n2336), .B(n2132), .Z(n2133) );
  NANDN U2778 ( .A(n2133), .B(n193), .Z(n2135) );
  XOR U2779 ( .A(b[29]), .B(a[1]), .Z(n2337) );
  NANDN U2780 ( .A(n193), .B(n2337), .Z(n2134) );
  AND U2781 ( .A(n2135), .B(n2134), .Z(n2335) );
  OR U2782 ( .A(n2136), .B(n192), .Z(n2138) );
  XOR U2783 ( .A(b[27]), .B(a[3]), .Z(n2301) );
  NAND U2784 ( .A(n38343), .B(n2301), .Z(n2137) );
  AND U2785 ( .A(n2138), .B(n2137), .Z(n2334) );
  XOR U2786 ( .A(n2335), .B(n2334), .Z(n2369) );
  NAND U2787 ( .A(b[0]), .B(a[29]), .Z(n2139) );
  XNOR U2788 ( .A(b[1]), .B(n2139), .Z(n2141) );
  NANDN U2789 ( .A(b[0]), .B(a[28]), .Z(n2140) );
  NAND U2790 ( .A(n2141), .B(n2140), .Z(n2367) );
  OR U2791 ( .A(n2142), .B(n178), .Z(n2144) );
  XNOR U2792 ( .A(b[15]), .B(a[15]), .Z(n2349) );
  OR U2793 ( .A(n2349), .B(n37509), .Z(n2143) );
  NAND U2794 ( .A(n2144), .B(n2143), .Z(n2368) );
  XOR U2795 ( .A(n2367), .B(n2368), .Z(n2370) );
  XOR U2796 ( .A(n2369), .B(n2370), .Z(n2329) );
  NAND U2797 ( .A(n187), .B(n2145), .Z(n2147) );
  XOR U2798 ( .A(b[13]), .B(a[17]), .Z(n2358) );
  NAND U2799 ( .A(n37295), .B(n2358), .Z(n2146) );
  AND U2800 ( .A(n2147), .B(n2146), .Z(n2376) );
  NAND U2801 ( .A(n190), .B(n2148), .Z(n2150) );
  XOR U2802 ( .A(b[19]), .B(a[11]), .Z(n2361) );
  NAND U2803 ( .A(n37821), .B(n2361), .Z(n2149) );
  AND U2804 ( .A(n2150), .B(n2149), .Z(n2374) );
  NAND U2805 ( .A(n186), .B(n2151), .Z(n2153) );
  XOR U2806 ( .A(b[11]), .B(a[19]), .Z(n2352) );
  NAND U2807 ( .A(n37097), .B(n2352), .Z(n2152) );
  NAND U2808 ( .A(n2153), .B(n2152), .Z(n2373) );
  XNOR U2809 ( .A(n2374), .B(n2373), .Z(n2375) );
  XNOR U2810 ( .A(n2376), .B(n2375), .Z(n2328) );
  XNOR U2811 ( .A(n2329), .B(n2328), .Z(n2330) );
  NANDN U2812 ( .A(n2155), .B(n2154), .Z(n2159) );
  NANDN U2813 ( .A(n2157), .B(n2156), .Z(n2158) );
  NAND U2814 ( .A(n2159), .B(n2158), .Z(n2331) );
  XNOR U2815 ( .A(n2330), .B(n2331), .Z(n2276) );
  NANDN U2816 ( .A(n2161), .B(n2160), .Z(n2165) );
  OR U2817 ( .A(n2163), .B(n2162), .Z(n2164) );
  AND U2818 ( .A(n2165), .B(n2164), .Z(n2274) );
  NANDN U2819 ( .A(n2167), .B(n2166), .Z(n2171) );
  OR U2820 ( .A(n2169), .B(n2168), .Z(n2170) );
  AND U2821 ( .A(n2171), .B(n2170), .Z(n2282) );
  NAND U2822 ( .A(n184), .B(n2172), .Z(n2174) );
  XOR U2823 ( .A(b[7]), .B(a[23]), .Z(n2364) );
  NAND U2824 ( .A(n36592), .B(n2364), .Z(n2173) );
  AND U2825 ( .A(n2174), .B(n2173), .Z(n2292) );
  NAND U2826 ( .A(n38064), .B(n2175), .Z(n2177) );
  XOR U2827 ( .A(b[21]), .B(a[9]), .Z(n2313) );
  NAND U2828 ( .A(n37993), .B(n2313), .Z(n2176) );
  NAND U2829 ( .A(n2177), .B(n2176), .Z(n2291) );
  XNOR U2830 ( .A(n2292), .B(n2291), .Z(n2294) );
  NAND U2831 ( .A(b[27]), .B(b[28]), .Z(n2178) );
  NAND U2832 ( .A(b[29]), .B(n2178), .Z(n38486) );
  OR U2833 ( .A(n38486), .B(n2197), .Z(n2293) );
  XNOR U2834 ( .A(n2294), .B(n2293), .Z(n2279) );
  NAND U2835 ( .A(n183), .B(n2179), .Z(n2181) );
  XOR U2836 ( .A(b[5]), .B(a[25]), .Z(n2343) );
  NAND U2837 ( .A(n36296), .B(n2343), .Z(n2180) );
  AND U2838 ( .A(n2181), .B(n2180), .Z(n2298) );
  NAND U2839 ( .A(n181), .B(n2182), .Z(n2184) );
  XOR U2840 ( .A(b[3]), .B(a[27]), .Z(n2346) );
  NAND U2841 ( .A(n182), .B(n2346), .Z(n2183) );
  AND U2842 ( .A(n2184), .B(n2183), .Z(n2296) );
  NAND U2843 ( .A(n189), .B(n2185), .Z(n2187) );
  XOR U2844 ( .A(b[17]), .B(a[13]), .Z(n2340) );
  NAND U2845 ( .A(n37652), .B(n2340), .Z(n2186) );
  NAND U2846 ( .A(n2187), .B(n2186), .Z(n2295) );
  XNOR U2847 ( .A(n2296), .B(n2295), .Z(n2297) );
  XOR U2848 ( .A(n2298), .B(n2297), .Z(n2280) );
  XNOR U2849 ( .A(n2279), .B(n2280), .Z(n2281) );
  XNOR U2850 ( .A(n2282), .B(n2281), .Z(n2273) );
  XNOR U2851 ( .A(n2274), .B(n2273), .Z(n2275) );
  XOR U2852 ( .A(n2276), .B(n2275), .Z(n2380) );
  NAND U2853 ( .A(n38185), .B(n2188), .Z(n2190) );
  XOR U2854 ( .A(b[23]), .B(a[7]), .Z(n2307) );
  NAND U2855 ( .A(n38132), .B(n2307), .Z(n2189) );
  AND U2856 ( .A(n2190), .B(n2189), .Z(n2287) );
  NAND U2857 ( .A(n38289), .B(n2191), .Z(n2193) );
  XOR U2858 ( .A(b[25]), .B(a[5]), .Z(n2310) );
  NAND U2859 ( .A(n38247), .B(n2310), .Z(n2192) );
  AND U2860 ( .A(n2193), .B(n2192), .Z(n2286) );
  OR U2861 ( .A(n2194), .B(n179), .Z(n2196) );
  XOR U2862 ( .A(b[9]), .B(a[21]), .Z(n2355) );
  NAND U2863 ( .A(n36805), .B(n2355), .Z(n2195) );
  NAND U2864 ( .A(n2196), .B(n2195), .Z(n2285) );
  XOR U2865 ( .A(n2286), .B(n2285), .Z(n2288) );
  XOR U2866 ( .A(n2287), .B(n2288), .Z(n2323) );
  NANDN U2867 ( .A(n2198), .B(n2197), .Z(n2202) );
  OR U2868 ( .A(n2200), .B(n2199), .Z(n2201) );
  AND U2869 ( .A(n2202), .B(n2201), .Z(n2322) );
  XNOR U2870 ( .A(n2323), .B(n2322), .Z(n2324) );
  NANDN U2871 ( .A(n2204), .B(n2203), .Z(n2208) );
  OR U2872 ( .A(n2206), .B(n2205), .Z(n2207) );
  NAND U2873 ( .A(n2208), .B(n2207), .Z(n2325) );
  XNOR U2874 ( .A(n2324), .B(n2325), .Z(n2379) );
  XNOR U2875 ( .A(n2380), .B(n2379), .Z(n2381) );
  NANDN U2876 ( .A(n2210), .B(n2209), .Z(n2214) );
  NANDN U2877 ( .A(n2212), .B(n2211), .Z(n2213) );
  NAND U2878 ( .A(n2214), .B(n2213), .Z(n2382) );
  XNOR U2879 ( .A(n2381), .B(n2382), .Z(n2270) );
  NANDN U2880 ( .A(n2216), .B(n2215), .Z(n2220) );
  NAND U2881 ( .A(n2218), .B(n2217), .Z(n2219) );
  AND U2882 ( .A(n2220), .B(n2219), .Z(n2268) );
  NANDN U2883 ( .A(n2222), .B(n2221), .Z(n2226) );
  NANDN U2884 ( .A(n2224), .B(n2223), .Z(n2225) );
  AND U2885 ( .A(n2226), .B(n2225), .Z(n2319) );
  NANDN U2886 ( .A(n2228), .B(n2227), .Z(n2232) );
  NAND U2887 ( .A(n2230), .B(n2229), .Z(n2231) );
  AND U2888 ( .A(n2232), .B(n2231), .Z(n2317) );
  NANDN U2889 ( .A(n2234), .B(n2233), .Z(n2238) );
  NANDN U2890 ( .A(n2236), .B(n2235), .Z(n2237) );
  NAND U2891 ( .A(n2238), .B(n2237), .Z(n2316) );
  XNOR U2892 ( .A(n2317), .B(n2316), .Z(n2318) );
  XNOR U2893 ( .A(n2319), .B(n2318), .Z(n2267) );
  XNOR U2894 ( .A(n2268), .B(n2267), .Z(n2269) );
  XOR U2895 ( .A(n2270), .B(n2269), .Z(n2386) );
  NANDN U2896 ( .A(n2240), .B(n2239), .Z(n2244) );
  OR U2897 ( .A(n2242), .B(n2241), .Z(n2243) );
  NAND U2898 ( .A(n2244), .B(n2243), .Z(n2385) );
  XOR U2899 ( .A(n2386), .B(n2385), .Z(n2388) );
  XOR U2900 ( .A(n2387), .B(n2388), .Z(n2262) );
  NANDN U2901 ( .A(n2246), .B(n2245), .Z(n2250) );
  NANDN U2902 ( .A(n2248), .B(n2247), .Z(n2249) );
  NAND U2903 ( .A(n2250), .B(n2249), .Z(n2261) );
  XNOR U2904 ( .A(n2262), .B(n2261), .Z(n2263) );
  XNOR U2905 ( .A(n2264), .B(n2263), .Z(n2256) );
  XNOR U2906 ( .A(sreg[253]), .B(n2256), .Z(n2258) );
  NANDN U2907 ( .A(sreg[252]), .B(n2251), .Z(n2255) );
  NAND U2908 ( .A(n2253), .B(n2252), .Z(n2254) );
  NAND U2909 ( .A(n2255), .B(n2254), .Z(n2257) );
  XNOR U2910 ( .A(n2258), .B(n2257), .Z(c[253]) );
  NANDN U2911 ( .A(sreg[253]), .B(n2256), .Z(n2260) );
  NAND U2912 ( .A(n2258), .B(n2257), .Z(n2259) );
  NAND U2913 ( .A(n2260), .B(n2259), .Z(n2532) );
  XNOR U2914 ( .A(sreg[254]), .B(n2532), .Z(n2534) );
  NANDN U2915 ( .A(n2262), .B(n2261), .Z(n2266) );
  NANDN U2916 ( .A(n2264), .B(n2263), .Z(n2265) );
  AND U2917 ( .A(n2266), .B(n2265), .Z(n2394) );
  NANDN U2918 ( .A(n2268), .B(n2267), .Z(n2272) );
  NAND U2919 ( .A(n2270), .B(n2269), .Z(n2271) );
  AND U2920 ( .A(n2272), .B(n2271), .Z(n2529) );
  NANDN U2921 ( .A(n2274), .B(n2273), .Z(n2278) );
  NAND U2922 ( .A(n2276), .B(n2275), .Z(n2277) );
  AND U2923 ( .A(n2278), .B(n2277), .Z(n2522) );
  NANDN U2924 ( .A(n2280), .B(n2279), .Z(n2284) );
  NANDN U2925 ( .A(n2282), .B(n2281), .Z(n2283) );
  AND U2926 ( .A(n2284), .B(n2283), .Z(n2521) );
  NANDN U2927 ( .A(n2286), .B(n2285), .Z(n2290) );
  OR U2928 ( .A(n2288), .B(n2287), .Z(n2289) );
  AND U2929 ( .A(n2290), .B(n2289), .Z(n2484) );
  XNOR U2930 ( .A(n2484), .B(n2483), .Z(n2485) );
  NANDN U2931 ( .A(n2296), .B(n2295), .Z(n2300) );
  NANDN U2932 ( .A(n2298), .B(n2297), .Z(n2299) );
  AND U2933 ( .A(n2300), .B(n2299), .Z(n2406) );
  XNOR U2934 ( .A(b[29]), .B(b[30]), .Z(n38493) );
  IV U2935 ( .A(n38493), .Z(n38453) );
  AND U2936 ( .A(a[0]), .B(n38453), .Z(n2514) );
  NAND U2937 ( .A(n38385), .B(n2301), .Z(n2303) );
  XOR U2938 ( .A(b[27]), .B(a[4]), .Z(n2421) );
  NAND U2939 ( .A(n38343), .B(n2421), .Z(n2302) );
  AND U2940 ( .A(n2303), .B(n2302), .Z(n2515) );
  XNOR U2941 ( .A(n2514), .B(n2515), .Z(n2516) );
  NAND U2942 ( .A(b[0]), .B(a[30]), .Z(n2304) );
  XNOR U2943 ( .A(b[1]), .B(n2304), .Z(n2306) );
  NANDN U2944 ( .A(b[0]), .B(a[29]), .Z(n2305) );
  NAND U2945 ( .A(n2306), .B(n2305), .Z(n2517) );
  XNOR U2946 ( .A(n2516), .B(n2517), .Z(n2403) );
  NAND U2947 ( .A(n38185), .B(n2307), .Z(n2309) );
  XOR U2948 ( .A(b[23]), .B(a[8]), .Z(n2415) );
  NAND U2949 ( .A(n38132), .B(n2415), .Z(n2308) );
  AND U2950 ( .A(n2309), .B(n2308), .Z(n2468) );
  NAND U2951 ( .A(n38289), .B(n2310), .Z(n2312) );
  XOR U2952 ( .A(b[25]), .B(a[6]), .Z(n2418) );
  NAND U2953 ( .A(n38247), .B(n2418), .Z(n2311) );
  AND U2954 ( .A(n2312), .B(n2311), .Z(n2466) );
  NAND U2955 ( .A(n38064), .B(n2313), .Z(n2315) );
  XOR U2956 ( .A(b[21]), .B(a[10]), .Z(n2427) );
  NAND U2957 ( .A(n37993), .B(n2427), .Z(n2314) );
  NAND U2958 ( .A(n2315), .B(n2314), .Z(n2465) );
  XNOR U2959 ( .A(n2466), .B(n2465), .Z(n2467) );
  XOR U2960 ( .A(n2468), .B(n2467), .Z(n2404) );
  XNOR U2961 ( .A(n2403), .B(n2404), .Z(n2405) );
  XOR U2962 ( .A(n2406), .B(n2405), .Z(n2486) );
  XNOR U2963 ( .A(n2485), .B(n2486), .Z(n2520) );
  XOR U2964 ( .A(n2521), .B(n2520), .Z(n2523) );
  XOR U2965 ( .A(n2522), .B(n2523), .Z(n2399) );
  NANDN U2966 ( .A(n2317), .B(n2316), .Z(n2321) );
  NANDN U2967 ( .A(n2319), .B(n2318), .Z(n2320) );
  AND U2968 ( .A(n2321), .B(n2320), .Z(n2398) );
  NANDN U2969 ( .A(n2323), .B(n2322), .Z(n2327) );
  NANDN U2970 ( .A(n2325), .B(n2324), .Z(n2326) );
  AND U2971 ( .A(n2327), .B(n2326), .Z(n2480) );
  NANDN U2972 ( .A(n2329), .B(n2328), .Z(n2333) );
  NANDN U2973 ( .A(n2331), .B(n2330), .Z(n2332) );
  AND U2974 ( .A(n2333), .B(n2332), .Z(n2477) );
  NOR U2975 ( .A(n2335), .B(n2334), .Z(n2455) );
  NANDN U2976 ( .A(n177), .B(n2337), .Z(n2339) );
  XNOR U2977 ( .A(b[29]), .B(a[2]), .Z(n2501) );
  OR U2978 ( .A(n2501), .B(n193), .Z(n2338) );
  AND U2979 ( .A(n2339), .B(n2338), .Z(n2453) );
  NANDN U2980 ( .A(n170), .B(n2340), .Z(n2342) );
  XNOR U2981 ( .A(b[17]), .B(a[14]), .Z(n2449) );
  OR U2982 ( .A(n2449), .B(n36922), .Z(n2341) );
  NAND U2983 ( .A(n2342), .B(n2341), .Z(n2454) );
  XOR U2984 ( .A(n2453), .B(n2454), .Z(n2456) );
  XOR U2985 ( .A(n2455), .B(n2456), .Z(n2410) );
  NAND U2986 ( .A(n183), .B(n2343), .Z(n2345) );
  XOR U2987 ( .A(b[5]), .B(a[26]), .Z(n2440) );
  NAND U2988 ( .A(n36296), .B(n2440), .Z(n2344) );
  AND U2989 ( .A(n2345), .B(n2344), .Z(n2474) );
  NAND U2990 ( .A(n181), .B(n2346), .Z(n2348) );
  XOR U2991 ( .A(b[3]), .B(a[28]), .Z(n2446) );
  NAND U2992 ( .A(n182), .B(n2446), .Z(n2347) );
  AND U2993 ( .A(n2348), .B(n2347), .Z(n2472) );
  OR U2994 ( .A(n2349), .B(n178), .Z(n2351) );
  XOR U2995 ( .A(b[15]), .B(a[16]), .Z(n2511) );
  NAND U2996 ( .A(n37382), .B(n2511), .Z(n2350) );
  NAND U2997 ( .A(n2351), .B(n2350), .Z(n2471) );
  XNOR U2998 ( .A(n2472), .B(n2471), .Z(n2473) );
  XNOR U2999 ( .A(n2474), .B(n2473), .Z(n2409) );
  XNOR U3000 ( .A(n2410), .B(n2409), .Z(n2412) );
  NAND U3001 ( .A(n186), .B(n2352), .Z(n2354) );
  XOR U3002 ( .A(b[11]), .B(a[20]), .Z(n2433) );
  NAND U3003 ( .A(n37097), .B(n2433), .Z(n2353) );
  AND U3004 ( .A(n2354), .B(n2353), .Z(n2460) );
  NAND U3005 ( .A(n185), .B(n2355), .Z(n2357) );
  XOR U3006 ( .A(b[9]), .B(a[22]), .Z(n2430) );
  NAND U3007 ( .A(n36805), .B(n2430), .Z(n2356) );
  NAND U3008 ( .A(n2357), .B(n2356), .Z(n2459) );
  XNOR U3009 ( .A(n2460), .B(n2459), .Z(n2461) );
  NAND U3010 ( .A(n187), .B(n2358), .Z(n2360) );
  XOR U3011 ( .A(b[13]), .B(a[18]), .Z(n2424) );
  NAND U3012 ( .A(n37295), .B(n2424), .Z(n2359) );
  AND U3013 ( .A(n2360), .B(n2359), .Z(n2498) );
  NAND U3014 ( .A(n190), .B(n2361), .Z(n2363) );
  XOR U3015 ( .A(b[19]), .B(a[12]), .Z(n2443) );
  NAND U3016 ( .A(n37821), .B(n2443), .Z(n2362) );
  AND U3017 ( .A(n2363), .B(n2362), .Z(n2496) );
  NAND U3018 ( .A(n184), .B(n2364), .Z(n2366) );
  XOR U3019 ( .A(b[7]), .B(a[24]), .Z(n2437) );
  NAND U3020 ( .A(n36592), .B(n2437), .Z(n2365) );
  NAND U3021 ( .A(n2366), .B(n2365), .Z(n2495) );
  XNOR U3022 ( .A(n2496), .B(n2495), .Z(n2497) );
  XOR U3023 ( .A(n2498), .B(n2497), .Z(n2462) );
  XNOR U3024 ( .A(n2461), .B(n2462), .Z(n2411) );
  XOR U3025 ( .A(n2412), .B(n2411), .Z(n2492) );
  NANDN U3026 ( .A(n2368), .B(n2367), .Z(n2372) );
  OR U3027 ( .A(n2370), .B(n2369), .Z(n2371) );
  AND U3028 ( .A(n2372), .B(n2371), .Z(n2490) );
  NANDN U3029 ( .A(n2374), .B(n2373), .Z(n2378) );
  NANDN U3030 ( .A(n2376), .B(n2375), .Z(n2377) );
  AND U3031 ( .A(n2378), .B(n2377), .Z(n2489) );
  XNOR U3032 ( .A(n2490), .B(n2489), .Z(n2491) );
  XOR U3033 ( .A(n2492), .B(n2491), .Z(n2478) );
  XNOR U3034 ( .A(n2477), .B(n2478), .Z(n2479) );
  XNOR U3035 ( .A(n2480), .B(n2479), .Z(n2397) );
  XOR U3036 ( .A(n2398), .B(n2397), .Z(n2400) );
  XOR U3037 ( .A(n2399), .B(n2400), .Z(n2527) );
  NANDN U3038 ( .A(n2380), .B(n2379), .Z(n2384) );
  NANDN U3039 ( .A(n2382), .B(n2381), .Z(n2383) );
  AND U3040 ( .A(n2384), .B(n2383), .Z(n2526) );
  XNOR U3041 ( .A(n2527), .B(n2526), .Z(n2528) );
  XOR U3042 ( .A(n2529), .B(n2528), .Z(n2392) );
  NANDN U3043 ( .A(n2386), .B(n2385), .Z(n2390) );
  OR U3044 ( .A(n2388), .B(n2387), .Z(n2389) );
  AND U3045 ( .A(n2390), .B(n2389), .Z(n2391) );
  XNOR U3046 ( .A(n2392), .B(n2391), .Z(n2393) );
  XNOR U3047 ( .A(n2394), .B(n2393), .Z(n2533) );
  XNOR U3048 ( .A(n2534), .B(n2533), .Z(c[254]) );
  NANDN U3049 ( .A(n2392), .B(n2391), .Z(n2396) );
  NANDN U3050 ( .A(n2394), .B(n2393), .Z(n2395) );
  AND U3051 ( .A(n2396), .B(n2395), .Z(n2545) );
  NANDN U3052 ( .A(n2398), .B(n2397), .Z(n2402) );
  OR U3053 ( .A(n2400), .B(n2399), .Z(n2401) );
  AND U3054 ( .A(n2402), .B(n2401), .Z(n2679) );
  NANDN U3055 ( .A(n2404), .B(n2403), .Z(n2408) );
  NANDN U3056 ( .A(n2406), .B(n2405), .Z(n2407) );
  AND U3057 ( .A(n2408), .B(n2407), .Z(n2671) );
  NANDN U3058 ( .A(n2410), .B(n2409), .Z(n2414) );
  NAND U3059 ( .A(n2412), .B(n2411), .Z(n2413) );
  NAND U3060 ( .A(n2414), .B(n2413), .Z(n2670) );
  XNOR U3061 ( .A(n2671), .B(n2670), .Z(n2672) );
  NAND U3062 ( .A(n38185), .B(n2415), .Z(n2417) );
  XOR U3063 ( .A(b[23]), .B(a[9]), .Z(n2610) );
  NAND U3064 ( .A(n38132), .B(n2610), .Z(n2416) );
  AND U3065 ( .A(n2417), .B(n2416), .Z(n2586) );
  NAND U3066 ( .A(n38289), .B(n2418), .Z(n2420) );
  XOR U3067 ( .A(b[25]), .B(a[7]), .Z(n2566) );
  NAND U3068 ( .A(n38247), .B(n2566), .Z(n2419) );
  AND U3069 ( .A(n2420), .B(n2419), .Z(n2585) );
  NAND U3070 ( .A(n38385), .B(n2421), .Z(n2423) );
  XOR U3071 ( .A(b[27]), .B(a[5]), .Z(n2569) );
  NAND U3072 ( .A(n38343), .B(n2569), .Z(n2422) );
  NAND U3073 ( .A(n2423), .B(n2422), .Z(n2584) );
  XOR U3074 ( .A(n2585), .B(n2584), .Z(n2587) );
  XOR U3075 ( .A(n2586), .B(n2587), .Z(n2562) );
  NAND U3076 ( .A(n187), .B(n2424), .Z(n2426) );
  XOR U3077 ( .A(b[13]), .B(a[19]), .Z(n2637) );
  NAND U3078 ( .A(n37295), .B(n2637), .Z(n2425) );
  AND U3079 ( .A(n2426), .B(n2425), .Z(n2648) );
  NAND U3080 ( .A(n38064), .B(n2427), .Z(n2429) );
  XOR U3081 ( .A(b[21]), .B(a[11]), .Z(n2631) );
  NAND U3082 ( .A(n37993), .B(n2631), .Z(n2428) );
  AND U3083 ( .A(n2429), .B(n2428), .Z(n2647) );
  NAND U3084 ( .A(n185), .B(n2430), .Z(n2432) );
  XOR U3085 ( .A(b[9]), .B(a[23]), .Z(n2604) );
  NAND U3086 ( .A(n36805), .B(n2604), .Z(n2431) );
  NAND U3087 ( .A(n2432), .B(n2431), .Z(n2646) );
  XOR U3088 ( .A(n2647), .B(n2646), .Z(n2649) );
  XOR U3089 ( .A(n2648), .B(n2649), .Z(n2561) );
  NANDN U3090 ( .A(n176), .B(n2433), .Z(n2436) );
  XNOR U3091 ( .A(b[11]), .B(a[21]), .Z(n2572) );
  OR U3092 ( .A(n2572), .B(n2434), .Z(n2435) );
  AND U3093 ( .A(n2436), .B(n2435), .Z(n2560) );
  XOR U3094 ( .A(n2561), .B(n2560), .Z(n2563) );
  XOR U3095 ( .A(n2562), .B(n2563), .Z(n2665) );
  NAND U3096 ( .A(n184), .B(n2437), .Z(n2439) );
  XOR U3097 ( .A(b[7]), .B(a[25]), .Z(n2575) );
  NAND U3098 ( .A(n36592), .B(n2575), .Z(n2438) );
  AND U3099 ( .A(n2439), .B(n2438), .Z(n2593) );
  NAND U3100 ( .A(n183), .B(n2440), .Z(n2442) );
  XOR U3101 ( .A(b[5]), .B(a[27]), .Z(n2578) );
  NAND U3102 ( .A(n36296), .B(n2578), .Z(n2441) );
  AND U3103 ( .A(n2442), .B(n2441), .Z(n2591) );
  NAND U3104 ( .A(n190), .B(n2443), .Z(n2445) );
  XOR U3105 ( .A(b[19]), .B(a[13]), .Z(n2581) );
  NAND U3106 ( .A(n37821), .B(n2581), .Z(n2444) );
  NAND U3107 ( .A(n2445), .B(n2444), .Z(n2590) );
  XNOR U3108 ( .A(n2591), .B(n2590), .Z(n2592) );
  XNOR U3109 ( .A(n2593), .B(n2592), .Z(n2652) );
  NAND U3110 ( .A(n181), .B(n2446), .Z(n2448) );
  XOR U3111 ( .A(b[3]), .B(a[29]), .Z(n2598) );
  NAND U3112 ( .A(n182), .B(n2598), .Z(n2447) );
  AND U3113 ( .A(n2448), .B(n2447), .Z(n2622) );
  OR U3114 ( .A(n2449), .B(n170), .Z(n2451) );
  XOR U3115 ( .A(b[17]), .B(a[15]), .Z(n2601) );
  NAND U3116 ( .A(n37652), .B(n2601), .Z(n2450) );
  AND U3117 ( .A(n2451), .B(n2450), .Z(n2620) );
  AND U3118 ( .A(b[29]), .B(b[30]), .Z(n38519) );
  NOR U3119 ( .A(n38519), .B(n2514), .Z(n2452) );
  AND U3120 ( .A(b[31]), .B(n2452), .Z(n2619) );
  XNOR U3121 ( .A(n2620), .B(n2619), .Z(n2621) );
  XOR U3122 ( .A(n2622), .B(n2621), .Z(n2653) );
  XNOR U3123 ( .A(n2652), .B(n2653), .Z(n2654) );
  NANDN U3124 ( .A(n2454), .B(n2453), .Z(n2458) );
  OR U3125 ( .A(n2456), .B(n2455), .Z(n2457) );
  NAND U3126 ( .A(n2458), .B(n2457), .Z(n2655) );
  XNOR U3127 ( .A(n2654), .B(n2655), .Z(n2664) );
  XNOR U3128 ( .A(n2665), .B(n2664), .Z(n2666) );
  NANDN U3129 ( .A(n2460), .B(n2459), .Z(n2464) );
  NANDN U3130 ( .A(n2462), .B(n2461), .Z(n2463) );
  AND U3131 ( .A(n2464), .B(n2463), .Z(n2616) );
  NANDN U3132 ( .A(n2466), .B(n2465), .Z(n2470) );
  NANDN U3133 ( .A(n2468), .B(n2467), .Z(n2469) );
  AND U3134 ( .A(n2470), .B(n2469), .Z(n2614) );
  NANDN U3135 ( .A(n2472), .B(n2471), .Z(n2476) );
  NANDN U3136 ( .A(n2474), .B(n2473), .Z(n2475) );
  NAND U3137 ( .A(n2476), .B(n2475), .Z(n2613) );
  XNOR U3138 ( .A(n2614), .B(n2613), .Z(n2615) );
  XOR U3139 ( .A(n2616), .B(n2615), .Z(n2667) );
  XOR U3140 ( .A(n2666), .B(n2667), .Z(n2673) );
  XNOR U3141 ( .A(n2672), .B(n2673), .Z(n2548) );
  NANDN U3142 ( .A(n2478), .B(n2477), .Z(n2482) );
  NANDN U3143 ( .A(n2480), .B(n2479), .Z(n2481) );
  NAND U3144 ( .A(n2482), .B(n2481), .Z(n2549) );
  XNOR U3145 ( .A(n2548), .B(n2549), .Z(n2551) );
  NANDN U3146 ( .A(n2484), .B(n2483), .Z(n2488) );
  NANDN U3147 ( .A(n2486), .B(n2485), .Z(n2487) );
  AND U3148 ( .A(n2488), .B(n2487), .Z(n2557) );
  NANDN U3149 ( .A(n2490), .B(n2489), .Z(n2494) );
  NANDN U3150 ( .A(n2492), .B(n2491), .Z(n2493) );
  AND U3151 ( .A(n2494), .B(n2493), .Z(n2554) );
  NANDN U3152 ( .A(n2496), .B(n2495), .Z(n2500) );
  NANDN U3153 ( .A(n2498), .B(n2497), .Z(n2499) );
  AND U3154 ( .A(n2500), .B(n2499), .Z(n2661) );
  OR U3155 ( .A(n2501), .B(n177), .Z(n2503) );
  XOR U3156 ( .A(b[29]), .B(a[3]), .Z(n2643) );
  NAND U3157 ( .A(n38456), .B(n2643), .Z(n2502) );
  AND U3158 ( .A(n2503), .B(n2502), .Z(n2597) );
  XOR U3159 ( .A(b[30]), .B(b[31]), .Z(n2504) );
  AND U3160 ( .A(n2504), .B(n38493), .Z(n38470) );
  XOR U3161 ( .A(a[0]), .B(b[31]), .Z(n2505) );
  NAND U3162 ( .A(n38470), .B(n2505), .Z(n2507) );
  XOR U3163 ( .A(b[31]), .B(a[1]), .Z(n2607) );
  AND U3164 ( .A(n2607), .B(n38453), .Z(n2506) );
  ANDN U3165 ( .B(n2507), .A(n2506), .Z(n2596) );
  XOR U3166 ( .A(n2597), .B(n2596), .Z(n2627) );
  NAND U3167 ( .A(b[0]), .B(a[31]), .Z(n2508) );
  XNOR U3168 ( .A(b[1]), .B(n2508), .Z(n2510) );
  NANDN U3169 ( .A(b[0]), .B(a[30]), .Z(n2509) );
  NAND U3170 ( .A(n2510), .B(n2509), .Z(n2625) );
  NANDN U3171 ( .A(n178), .B(n2511), .Z(n2513) );
  XNOR U3172 ( .A(b[15]), .B(a[17]), .Z(n2634) );
  OR U3173 ( .A(n2634), .B(n37509), .Z(n2512) );
  NAND U3174 ( .A(n2513), .B(n2512), .Z(n2626) );
  XOR U3175 ( .A(n2625), .B(n2626), .Z(n2628) );
  XOR U3176 ( .A(n2627), .B(n2628), .Z(n2659) );
  NANDN U3177 ( .A(n2515), .B(n2514), .Z(n2519) );
  NANDN U3178 ( .A(n2517), .B(n2516), .Z(n2518) );
  NAND U3179 ( .A(n2519), .B(n2518), .Z(n2658) );
  XNOR U3180 ( .A(n2659), .B(n2658), .Z(n2660) );
  XOR U3181 ( .A(n2661), .B(n2660), .Z(n2555) );
  XNOR U3182 ( .A(n2554), .B(n2555), .Z(n2556) );
  XNOR U3183 ( .A(n2557), .B(n2556), .Z(n2550) );
  XOR U3184 ( .A(n2551), .B(n2550), .Z(n2677) );
  NANDN U3185 ( .A(n2521), .B(n2520), .Z(n2525) );
  OR U3186 ( .A(n2523), .B(n2522), .Z(n2524) );
  AND U3187 ( .A(n2525), .B(n2524), .Z(n2676) );
  XNOR U3188 ( .A(n2677), .B(n2676), .Z(n2678) );
  XNOR U3189 ( .A(n2679), .B(n2678), .Z(n2542) );
  NANDN U3190 ( .A(n2527), .B(n2526), .Z(n2531) );
  NAND U3191 ( .A(n2529), .B(n2528), .Z(n2530) );
  NAND U3192 ( .A(n2531), .B(n2530), .Z(n2543) );
  XNOR U3193 ( .A(n2542), .B(n2543), .Z(n2544) );
  XNOR U3194 ( .A(n2545), .B(n2544), .Z(n2537) );
  XNOR U3195 ( .A(sreg[255]), .B(n2537), .Z(n2539) );
  NANDN U3196 ( .A(sreg[254]), .B(n2532), .Z(n2536) );
  NAND U3197 ( .A(n2534), .B(n2533), .Z(n2535) );
  NAND U3198 ( .A(n2536), .B(n2535), .Z(n2538) );
  XNOR U3199 ( .A(n2539), .B(n2538), .Z(c[255]) );
  NANDN U3200 ( .A(sreg[255]), .B(n2537), .Z(n2541) );
  NAND U3201 ( .A(n2539), .B(n2538), .Z(n2540) );
  NAND U3202 ( .A(n2541), .B(n2540), .Z(n2826) );
  XNOR U3203 ( .A(sreg[256]), .B(n2826), .Z(n2828) );
  NANDN U3204 ( .A(n2543), .B(n2542), .Z(n2547) );
  NANDN U3205 ( .A(n2545), .B(n2544), .Z(n2546) );
  AND U3206 ( .A(n2547), .B(n2546), .Z(n2684) );
  NANDN U3207 ( .A(n2549), .B(n2548), .Z(n2553) );
  NAND U3208 ( .A(n2551), .B(n2550), .Z(n2552) );
  AND U3209 ( .A(n2553), .B(n2552), .Z(n2822) );
  NANDN U3210 ( .A(n2555), .B(n2554), .Z(n2559) );
  NANDN U3211 ( .A(n2557), .B(n2556), .Z(n2558) );
  AND U3212 ( .A(n2559), .B(n2558), .Z(n2821) );
  NANDN U3213 ( .A(n2561), .B(n2560), .Z(n2565) );
  OR U3214 ( .A(n2563), .B(n2562), .Z(n2564) );
  AND U3215 ( .A(n2565), .B(n2564), .Z(n2721) );
  NAND U3216 ( .A(n38289), .B(n2566), .Z(n2568) );
  XOR U3217 ( .A(b[25]), .B(a[8]), .Z(n2745) );
  NAND U3218 ( .A(n38247), .B(n2745), .Z(n2567) );
  AND U3219 ( .A(n2568), .B(n2567), .Z(n2765) );
  NAND U3220 ( .A(n38385), .B(n2569), .Z(n2571) );
  XOR U3221 ( .A(b[27]), .B(a[6]), .Z(n2754) );
  NAND U3222 ( .A(n38343), .B(n2754), .Z(n2570) );
  AND U3223 ( .A(n2571), .B(n2570), .Z(n2764) );
  OR U3224 ( .A(n2572), .B(n176), .Z(n2574) );
  XOR U3225 ( .A(b[11]), .B(a[22]), .Z(n2739) );
  NAND U3226 ( .A(n37097), .B(n2739), .Z(n2573) );
  NAND U3227 ( .A(n2574), .B(n2573), .Z(n2763) );
  XOR U3228 ( .A(n2764), .B(n2763), .Z(n2766) );
  XOR U3229 ( .A(n2765), .B(n2766), .Z(n2701) );
  NAND U3230 ( .A(n184), .B(n2575), .Z(n2577) );
  XOR U3231 ( .A(b[7]), .B(a[26]), .Z(n2730) );
  NAND U3232 ( .A(n36592), .B(n2730), .Z(n2576) );
  AND U3233 ( .A(n2577), .B(n2576), .Z(n2792) );
  NAND U3234 ( .A(n183), .B(n2578), .Z(n2580) );
  XOR U3235 ( .A(b[5]), .B(a[28]), .Z(n2733) );
  NAND U3236 ( .A(n36296), .B(n2733), .Z(n2579) );
  AND U3237 ( .A(n2580), .B(n2579), .Z(n2791) );
  NAND U3238 ( .A(n190), .B(n2581), .Z(n2583) );
  XOR U3239 ( .A(b[19]), .B(a[14]), .Z(n2781) );
  NAND U3240 ( .A(n37821), .B(n2781), .Z(n2582) );
  NAND U3241 ( .A(n2583), .B(n2582), .Z(n2790) );
  XOR U3242 ( .A(n2791), .B(n2790), .Z(n2793) );
  XNOR U3243 ( .A(n2792), .B(n2793), .Z(n2700) );
  XNOR U3244 ( .A(n2701), .B(n2700), .Z(n2703) );
  NANDN U3245 ( .A(n2585), .B(n2584), .Z(n2589) );
  OR U3246 ( .A(n2587), .B(n2586), .Z(n2588) );
  AND U3247 ( .A(n2589), .B(n2588), .Z(n2702) );
  XOR U3248 ( .A(n2703), .B(n2702), .Z(n2719) );
  NANDN U3249 ( .A(n2591), .B(n2590), .Z(n2595) );
  NANDN U3250 ( .A(n2593), .B(n2592), .Z(n2594) );
  AND U3251 ( .A(n2595), .B(n2594), .Z(n2709) );
  NOR U3252 ( .A(n2597), .B(n2596), .Z(n2727) );
  NANDN U3253 ( .A(n180), .B(n2598), .Z(n2600) );
  XNOR U3254 ( .A(b[3]), .B(a[30]), .Z(n2742) );
  OR U3255 ( .A(n2742), .B(n172), .Z(n2599) );
  AND U3256 ( .A(n2600), .B(n2599), .Z(n2725) );
  NANDN U3257 ( .A(n170), .B(n2601), .Z(n2603) );
  XNOR U3258 ( .A(b[17]), .B(a[16]), .Z(n2760) );
  OR U3259 ( .A(n2760), .B(n36922), .Z(n2602) );
  AND U3260 ( .A(n2603), .B(n2602), .Z(n2724) );
  XOR U3261 ( .A(n2725), .B(n2724), .Z(n2726) );
  XOR U3262 ( .A(n2727), .B(n2726), .Z(n2707) );
  NAND U3263 ( .A(n185), .B(n2604), .Z(n2606) );
  XOR U3264 ( .A(b[9]), .B(a[24]), .Z(n2736) );
  NAND U3265 ( .A(n36805), .B(n2736), .Z(n2605) );
  AND U3266 ( .A(n2606), .B(n2605), .Z(n2805) );
  NAND U3267 ( .A(n38470), .B(n2607), .Z(n2609) );
  XOR U3268 ( .A(b[31]), .B(a[2]), .Z(n2757) );
  NAND U3269 ( .A(n38453), .B(n2757), .Z(n2608) );
  AND U3270 ( .A(n2609), .B(n2608), .Z(n2803) );
  NAND U3271 ( .A(n38185), .B(n2610), .Z(n2612) );
  XOR U3272 ( .A(b[23]), .B(a[10]), .Z(n2778) );
  NAND U3273 ( .A(n38132), .B(n2778), .Z(n2611) );
  NAND U3274 ( .A(n2612), .B(n2611), .Z(n2802) );
  XNOR U3275 ( .A(n2803), .B(n2802), .Z(n2804) );
  XNOR U3276 ( .A(n2805), .B(n2804), .Z(n2706) );
  XOR U3277 ( .A(n2707), .B(n2706), .Z(n2708) );
  XNOR U3278 ( .A(n2709), .B(n2708), .Z(n2718) );
  XNOR U3279 ( .A(n2719), .B(n2718), .Z(n2720) );
  XOR U3280 ( .A(n2721), .B(n2720), .Z(n2689) );
  NANDN U3281 ( .A(n2614), .B(n2613), .Z(n2618) );
  NANDN U3282 ( .A(n2616), .B(n2615), .Z(n2617) );
  AND U3283 ( .A(n2618), .B(n2617), .Z(n2688) );
  XNOR U3284 ( .A(n2689), .B(n2688), .Z(n2691) );
  NANDN U3285 ( .A(n2620), .B(n2619), .Z(n2624) );
  NANDN U3286 ( .A(n2622), .B(n2621), .Z(n2623) );
  AND U3287 ( .A(n2624), .B(n2623), .Z(n2713) );
  NANDN U3288 ( .A(n2626), .B(n2625), .Z(n2630) );
  OR U3289 ( .A(n2628), .B(n2627), .Z(n2629) );
  AND U3290 ( .A(n2630), .B(n2629), .Z(n2712) );
  XNOR U3291 ( .A(n2713), .B(n2712), .Z(n2715) );
  NAND U3292 ( .A(n38064), .B(n2631), .Z(n2633) );
  XOR U3293 ( .A(b[21]), .B(a[12]), .Z(n2775) );
  NAND U3294 ( .A(n37993), .B(n2775), .Z(n2632) );
  AND U3295 ( .A(n2633), .B(n2632), .Z(n2772) );
  OR U3296 ( .A(n2634), .B(n178), .Z(n2636) );
  XOR U3297 ( .A(b[15]), .B(a[18]), .Z(n2784) );
  NAND U3298 ( .A(n37382), .B(n2784), .Z(n2635) );
  AND U3299 ( .A(n2636), .B(n2635), .Z(n2770) );
  NAND U3300 ( .A(n187), .B(n2637), .Z(n2639) );
  XOR U3301 ( .A(b[13]), .B(a[20]), .Z(n2751) );
  NAND U3302 ( .A(n37295), .B(n2751), .Z(n2638) );
  NAND U3303 ( .A(n2639), .B(n2638), .Z(n2769) );
  XNOR U3304 ( .A(n2770), .B(n2769), .Z(n2771) );
  XNOR U3305 ( .A(n2772), .B(n2771), .Z(n2809) );
  NAND U3306 ( .A(b[0]), .B(a[32]), .Z(n2640) );
  XNOR U3307 ( .A(b[1]), .B(n2640), .Z(n2642) );
  NANDN U3308 ( .A(b[0]), .B(a[31]), .Z(n2641) );
  NAND U3309 ( .A(n2642), .B(n2641), .Z(n2799) );
  NAND U3310 ( .A(n194), .B(n2643), .Z(n2645) );
  XOR U3311 ( .A(b[29]), .B(a[4]), .Z(n2787) );
  NAND U3312 ( .A(n38456), .B(n2787), .Z(n2644) );
  AND U3313 ( .A(n2645), .B(n2644), .Z(n2797) );
  AND U3314 ( .A(b[31]), .B(a[0]), .Z(n2796) );
  XOR U3315 ( .A(n2797), .B(n2796), .Z(n2798) );
  XOR U3316 ( .A(n2799), .B(n2798), .Z(n2808) );
  XOR U3317 ( .A(n2809), .B(n2808), .Z(n2811) );
  NANDN U3318 ( .A(n2647), .B(n2646), .Z(n2651) );
  OR U3319 ( .A(n2649), .B(n2648), .Z(n2650) );
  NAND U3320 ( .A(n2651), .B(n2650), .Z(n2810) );
  XOR U3321 ( .A(n2811), .B(n2810), .Z(n2714) );
  XOR U3322 ( .A(n2715), .B(n2714), .Z(n2695) );
  NANDN U3323 ( .A(n2653), .B(n2652), .Z(n2657) );
  NANDN U3324 ( .A(n2655), .B(n2654), .Z(n2656) );
  AND U3325 ( .A(n2657), .B(n2656), .Z(n2694) );
  XNOR U3326 ( .A(n2695), .B(n2694), .Z(n2696) );
  NANDN U3327 ( .A(n2659), .B(n2658), .Z(n2663) );
  NANDN U3328 ( .A(n2661), .B(n2660), .Z(n2662) );
  NAND U3329 ( .A(n2663), .B(n2662), .Z(n2697) );
  XNOR U3330 ( .A(n2696), .B(n2697), .Z(n2690) );
  XOR U3331 ( .A(n2691), .B(n2690), .Z(n2817) );
  NANDN U3332 ( .A(n2665), .B(n2664), .Z(n2669) );
  NANDN U3333 ( .A(n2667), .B(n2666), .Z(n2668) );
  AND U3334 ( .A(n2669), .B(n2668), .Z(n2815) );
  NANDN U3335 ( .A(n2671), .B(n2670), .Z(n2675) );
  NANDN U3336 ( .A(n2673), .B(n2672), .Z(n2674) );
  NAND U3337 ( .A(n2675), .B(n2674), .Z(n2814) );
  XNOR U3338 ( .A(n2815), .B(n2814), .Z(n2816) );
  XNOR U3339 ( .A(n2817), .B(n2816), .Z(n2820) );
  XOR U3340 ( .A(n2821), .B(n2820), .Z(n2823) );
  XOR U3341 ( .A(n2822), .B(n2823), .Z(n2683) );
  NANDN U3342 ( .A(n2677), .B(n2676), .Z(n2681) );
  NANDN U3343 ( .A(n2679), .B(n2678), .Z(n2680) );
  NAND U3344 ( .A(n2681), .B(n2680), .Z(n2682) );
  XOR U3345 ( .A(n2683), .B(n2682), .Z(n2685) );
  XNOR U3346 ( .A(n2684), .B(n2685), .Z(n2827) );
  XOR U3347 ( .A(n2828), .B(n2827), .Z(c[256]) );
  NANDN U3348 ( .A(n2683), .B(n2682), .Z(n2687) );
  OR U3349 ( .A(n2685), .B(n2684), .Z(n2686) );
  AND U3350 ( .A(n2687), .B(n2686), .Z(n2834) );
  NANDN U3351 ( .A(n2689), .B(n2688), .Z(n2693) );
  NAND U3352 ( .A(n2691), .B(n2690), .Z(n2692) );
  AND U3353 ( .A(n2693), .B(n2692), .Z(n2846) );
  NANDN U3354 ( .A(n2695), .B(n2694), .Z(n2699) );
  NANDN U3355 ( .A(n2697), .B(n2696), .Z(n2698) );
  AND U3356 ( .A(n2699), .B(n2698), .Z(n2844) );
  NANDN U3357 ( .A(n2701), .B(n2700), .Z(n2705) );
  NAND U3358 ( .A(n2703), .B(n2702), .Z(n2704) );
  AND U3359 ( .A(n2705), .B(n2704), .Z(n2856) );
  NAND U3360 ( .A(n2707), .B(n2706), .Z(n2711) );
  NANDN U3361 ( .A(n2709), .B(n2708), .Z(n2710) );
  AND U3362 ( .A(n2711), .B(n2710), .Z(n2855) );
  XNOR U3363 ( .A(n2856), .B(n2855), .Z(n2857) );
  NANDN U3364 ( .A(n2713), .B(n2712), .Z(n2717) );
  NAND U3365 ( .A(n2715), .B(n2714), .Z(n2716) );
  NAND U3366 ( .A(n2717), .B(n2716), .Z(n2858) );
  XNOR U3367 ( .A(n2857), .B(n2858), .Z(n2843) );
  XNOR U3368 ( .A(n2844), .B(n2843), .Z(n2845) );
  XNOR U3369 ( .A(n2846), .B(n2845), .Z(n2837) );
  NANDN U3370 ( .A(n2719), .B(n2718), .Z(n2723) );
  NAND U3371 ( .A(n2721), .B(n2720), .Z(n2722) );
  AND U3372 ( .A(n2723), .B(n2722), .Z(n2971) );
  NAND U3373 ( .A(n2725), .B(n2724), .Z(n2729) );
  NANDN U3374 ( .A(n2727), .B(n2726), .Z(n2728) );
  AND U3375 ( .A(n2729), .B(n2728), .Z(n2849) );
  NAND U3376 ( .A(n184), .B(n2730), .Z(n2732) );
  XOR U3377 ( .A(b[7]), .B(a[27]), .Z(n2948) );
  NAND U3378 ( .A(n36592), .B(n2948), .Z(n2731) );
  AND U3379 ( .A(n2732), .B(n2731), .Z(n2880) );
  NAND U3380 ( .A(n183), .B(n2733), .Z(n2735) );
  XOR U3381 ( .A(b[5]), .B(a[29]), .Z(n2897) );
  NAND U3382 ( .A(n36296), .B(n2897), .Z(n2734) );
  NAND U3383 ( .A(n2735), .B(n2734), .Z(n2879) );
  XNOR U3384 ( .A(n2880), .B(n2879), .Z(n2882) );
  NAND U3385 ( .A(n185), .B(n2736), .Z(n2738) );
  XOR U3386 ( .A(b[9]), .B(a[25]), .Z(n2966) );
  NAND U3387 ( .A(n36805), .B(n2966), .Z(n2737) );
  AND U3388 ( .A(n2738), .B(n2737), .Z(n2876) );
  NAND U3389 ( .A(n186), .B(n2739), .Z(n2741) );
  XOR U3390 ( .A(b[11]), .B(a[23]), .Z(n2957) );
  NAND U3391 ( .A(n37097), .B(n2957), .Z(n2740) );
  AND U3392 ( .A(n2741), .B(n2740), .Z(n2874) );
  OR U3393 ( .A(n2742), .B(n180), .Z(n2744) );
  XOR U3394 ( .A(b[3]), .B(a[31]), .Z(n2888) );
  NAND U3395 ( .A(n182), .B(n2888), .Z(n2743) );
  NAND U3396 ( .A(n2744), .B(n2743), .Z(n2873) );
  XNOR U3397 ( .A(n2874), .B(n2873), .Z(n2875) );
  XNOR U3398 ( .A(n2876), .B(n2875), .Z(n2881) );
  XOR U3399 ( .A(n2882), .B(n2881), .Z(n2923) );
  NAND U3400 ( .A(n38289), .B(n2745), .Z(n2747) );
  XOR U3401 ( .A(b[25]), .B(a[9]), .Z(n2951) );
  NAND U3402 ( .A(n38247), .B(n2951), .Z(n2746) );
  AND U3403 ( .A(n2747), .B(n2746), .Z(n2929) );
  NAND U3404 ( .A(b[0]), .B(a[33]), .Z(n2748) );
  XNOR U3405 ( .A(b[1]), .B(n2748), .Z(n2750) );
  NANDN U3406 ( .A(b[0]), .B(a[32]), .Z(n2749) );
  NAND U3407 ( .A(n2750), .B(n2749), .Z(n2928) );
  NAND U3408 ( .A(n187), .B(n2751), .Z(n2753) );
  XOR U3409 ( .A(b[13]), .B(a[21]), .Z(n2954) );
  NAND U3410 ( .A(n37295), .B(n2954), .Z(n2752) );
  NAND U3411 ( .A(n2753), .B(n2752), .Z(n2927) );
  XOR U3412 ( .A(n2928), .B(n2927), .Z(n2930) );
  XOR U3413 ( .A(n2929), .B(n2930), .Z(n2922) );
  NAND U3414 ( .A(n38385), .B(n2754), .Z(n2756) );
  XOR U3415 ( .A(b[27]), .B(a[7]), .Z(n2894) );
  NAND U3416 ( .A(n38343), .B(n2894), .Z(n2755) );
  AND U3417 ( .A(n2756), .B(n2755), .Z(n2869) );
  NAND U3418 ( .A(n38470), .B(n2757), .Z(n2759) );
  XOR U3419 ( .A(b[31]), .B(a[3]), .Z(n2885) );
  NAND U3420 ( .A(n38453), .B(n2885), .Z(n2758) );
  AND U3421 ( .A(n2759), .B(n2758), .Z(n2868) );
  OR U3422 ( .A(n2760), .B(n170), .Z(n2762) );
  XOR U3423 ( .A(b[17]), .B(a[17]), .Z(n2891) );
  NAND U3424 ( .A(n37652), .B(n2891), .Z(n2761) );
  NAND U3425 ( .A(n2762), .B(n2761), .Z(n2867) );
  XOR U3426 ( .A(n2868), .B(n2867), .Z(n2870) );
  XNOR U3427 ( .A(n2869), .B(n2870), .Z(n2921) );
  XOR U3428 ( .A(n2922), .B(n2921), .Z(n2924) );
  XOR U3429 ( .A(n2923), .B(n2924), .Z(n2912) );
  NANDN U3430 ( .A(n2764), .B(n2763), .Z(n2768) );
  OR U3431 ( .A(n2766), .B(n2765), .Z(n2767) );
  AND U3432 ( .A(n2768), .B(n2767), .Z(n2910) );
  NANDN U3433 ( .A(n2770), .B(n2769), .Z(n2774) );
  NANDN U3434 ( .A(n2772), .B(n2771), .Z(n2773) );
  NAND U3435 ( .A(n2774), .B(n2773), .Z(n2909) );
  XNOR U3436 ( .A(n2910), .B(n2909), .Z(n2911) );
  XOR U3437 ( .A(n2912), .B(n2911), .Z(n2850) );
  XNOR U3438 ( .A(n2849), .B(n2850), .Z(n2852) );
  NAND U3439 ( .A(n38064), .B(n2775), .Z(n2777) );
  XOR U3440 ( .A(b[21]), .B(a[13]), .Z(n2963) );
  NAND U3441 ( .A(n37993), .B(n2963), .Z(n2776) );
  AND U3442 ( .A(n2777), .B(n2776), .Z(n2935) );
  NAND U3443 ( .A(n38185), .B(n2778), .Z(n2780) );
  XOR U3444 ( .A(b[23]), .B(a[11]), .Z(n2945) );
  NAND U3445 ( .A(n38132), .B(n2945), .Z(n2779) );
  AND U3446 ( .A(n2780), .B(n2779), .Z(n2934) );
  NAND U3447 ( .A(n190), .B(n2781), .Z(n2783) );
  XOR U3448 ( .A(b[19]), .B(a[15]), .Z(n2900) );
  NAND U3449 ( .A(n37821), .B(n2900), .Z(n2782) );
  NAND U3450 ( .A(n2783), .B(n2782), .Z(n2933) );
  XOR U3451 ( .A(n2934), .B(n2933), .Z(n2936) );
  XOR U3452 ( .A(n2935), .B(n2936), .Z(n2862) );
  NAND U3453 ( .A(n188), .B(n2784), .Z(n2786) );
  XOR U3454 ( .A(b[15]), .B(a[19]), .Z(n2960) );
  NAND U3455 ( .A(n37382), .B(n2960), .Z(n2785) );
  AND U3456 ( .A(n2786), .B(n2785), .Z(n2905) );
  NAND U3457 ( .A(n194), .B(n2787), .Z(n2789) );
  XOR U3458 ( .A(b[29]), .B(a[5]), .Z(n2942) );
  NAND U3459 ( .A(n38456), .B(n2942), .Z(n2788) );
  AND U3460 ( .A(n2789), .B(n2788), .Z(n2904) );
  AND U3461 ( .A(b[31]), .B(a[1]), .Z(n2903) );
  XOR U3462 ( .A(n2904), .B(n2903), .Z(n2906) );
  XNOR U3463 ( .A(n2905), .B(n2906), .Z(n2861) );
  XNOR U3464 ( .A(n2862), .B(n2861), .Z(n2864) );
  NANDN U3465 ( .A(n2791), .B(n2790), .Z(n2795) );
  OR U3466 ( .A(n2793), .B(n2792), .Z(n2794) );
  AND U3467 ( .A(n2795), .B(n2794), .Z(n2863) );
  XOR U3468 ( .A(n2864), .B(n2863), .Z(n2918) );
  NANDN U3469 ( .A(n2797), .B(n2796), .Z(n2801) );
  OR U3470 ( .A(n2799), .B(n2798), .Z(n2800) );
  AND U3471 ( .A(n2801), .B(n2800), .Z(n2916) );
  NANDN U3472 ( .A(n2803), .B(n2802), .Z(n2807) );
  NANDN U3473 ( .A(n2805), .B(n2804), .Z(n2806) );
  NAND U3474 ( .A(n2807), .B(n2806), .Z(n2915) );
  XNOR U3475 ( .A(n2916), .B(n2915), .Z(n2917) );
  XNOR U3476 ( .A(n2918), .B(n2917), .Z(n2851) );
  XOR U3477 ( .A(n2852), .B(n2851), .Z(n2970) );
  NAND U3478 ( .A(n2809), .B(n2808), .Z(n2813) );
  NAND U3479 ( .A(n2811), .B(n2810), .Z(n2812) );
  AND U3480 ( .A(n2813), .B(n2812), .Z(n2969) );
  XOR U3481 ( .A(n2970), .B(n2969), .Z(n2972) );
  XOR U3482 ( .A(n2971), .B(n2972), .Z(n2838) );
  XNOR U3483 ( .A(n2837), .B(n2838), .Z(n2839) );
  NANDN U3484 ( .A(n2815), .B(n2814), .Z(n2819) );
  NANDN U3485 ( .A(n2817), .B(n2816), .Z(n2818) );
  NAND U3486 ( .A(n2819), .B(n2818), .Z(n2840) );
  XNOR U3487 ( .A(n2839), .B(n2840), .Z(n2831) );
  NANDN U3488 ( .A(n2821), .B(n2820), .Z(n2825) );
  OR U3489 ( .A(n2823), .B(n2822), .Z(n2824) );
  NAND U3490 ( .A(n2825), .B(n2824), .Z(n2832) );
  XNOR U3491 ( .A(n2831), .B(n2832), .Z(n2833) );
  XNOR U3492 ( .A(n2834), .B(n2833), .Z(n2975) );
  XNOR U3493 ( .A(sreg[257]), .B(n2975), .Z(n2977) );
  NANDN U3494 ( .A(n2826), .B(sreg[256]), .Z(n2830) );
  NAND U3495 ( .A(n2828), .B(n2827), .Z(n2829) );
  AND U3496 ( .A(n2830), .B(n2829), .Z(n2976) );
  XNOR U3497 ( .A(n2977), .B(n2976), .Z(c[257]) );
  NANDN U3498 ( .A(n2832), .B(n2831), .Z(n2836) );
  NANDN U3499 ( .A(n2834), .B(n2833), .Z(n2835) );
  AND U3500 ( .A(n2836), .B(n2835), .Z(n2983) );
  NANDN U3501 ( .A(n2838), .B(n2837), .Z(n2842) );
  NANDN U3502 ( .A(n2840), .B(n2839), .Z(n2841) );
  AND U3503 ( .A(n2842), .B(n2841), .Z(n2981) );
  NANDN U3504 ( .A(n2844), .B(n2843), .Z(n2848) );
  NANDN U3505 ( .A(n2846), .B(n2845), .Z(n2847) );
  AND U3506 ( .A(n2848), .B(n2847), .Z(n2989) );
  NANDN U3507 ( .A(n2850), .B(n2849), .Z(n2854) );
  NAND U3508 ( .A(n2852), .B(n2851), .Z(n2853) );
  AND U3509 ( .A(n2854), .B(n2853), .Z(n3119) );
  NANDN U3510 ( .A(n2856), .B(n2855), .Z(n2860) );
  NANDN U3511 ( .A(n2858), .B(n2857), .Z(n2859) );
  AND U3512 ( .A(n2860), .B(n2859), .Z(n3118) );
  XNOR U3513 ( .A(n3119), .B(n3118), .Z(n3121) );
  NANDN U3514 ( .A(n2862), .B(n2861), .Z(n2866) );
  NAND U3515 ( .A(n2864), .B(n2863), .Z(n2865) );
  AND U3516 ( .A(n2866), .B(n2865), .Z(n3000) );
  NANDN U3517 ( .A(n2868), .B(n2867), .Z(n2872) );
  OR U3518 ( .A(n2870), .B(n2869), .Z(n2871) );
  AND U3519 ( .A(n2872), .B(n2871), .Z(n3106) );
  NANDN U3520 ( .A(n2874), .B(n2873), .Z(n2878) );
  NANDN U3521 ( .A(n2876), .B(n2875), .Z(n2877) );
  NAND U3522 ( .A(n2878), .B(n2877), .Z(n3107) );
  XNOR U3523 ( .A(n3106), .B(n3107), .Z(n3108) );
  NANDN U3524 ( .A(n2880), .B(n2879), .Z(n2884) );
  NAND U3525 ( .A(n2882), .B(n2881), .Z(n2883) );
  NAND U3526 ( .A(n2884), .B(n2883), .Z(n3109) );
  XNOR U3527 ( .A(n3108), .B(n3109), .Z(n2998) );
  NAND U3528 ( .A(n38470), .B(n2885), .Z(n2887) );
  XOR U3529 ( .A(b[31]), .B(a[4]), .Z(n3019) );
  NAND U3530 ( .A(n38453), .B(n3019), .Z(n2886) );
  AND U3531 ( .A(n2887), .B(n2886), .Z(n3030) );
  NAND U3532 ( .A(n181), .B(n2888), .Z(n2890) );
  XOR U3533 ( .A(b[3]), .B(a[32]), .Z(n3022) );
  NAND U3534 ( .A(n182), .B(n3022), .Z(n2889) );
  AND U3535 ( .A(n2890), .B(n2889), .Z(n3029) );
  NAND U3536 ( .A(n189), .B(n2891), .Z(n2893) );
  XOR U3537 ( .A(b[17]), .B(a[18]), .Z(n3025) );
  NAND U3538 ( .A(n37652), .B(n3025), .Z(n2892) );
  NAND U3539 ( .A(n2893), .B(n2892), .Z(n3028) );
  XOR U3540 ( .A(n3029), .B(n3028), .Z(n3031) );
  XOR U3541 ( .A(n3030), .B(n3031), .Z(n3095) );
  NAND U3542 ( .A(n38385), .B(n2894), .Z(n2896) );
  XOR U3543 ( .A(b[27]), .B(a[8]), .Z(n3010) );
  NAND U3544 ( .A(n38343), .B(n3010), .Z(n2895) );
  AND U3545 ( .A(n2896), .B(n2895), .Z(n3054) );
  NAND U3546 ( .A(n183), .B(n2897), .Z(n2899) );
  XOR U3547 ( .A(b[5]), .B(a[30]), .Z(n3013) );
  NAND U3548 ( .A(n36296), .B(n3013), .Z(n2898) );
  AND U3549 ( .A(n2899), .B(n2898), .Z(n3053) );
  NAND U3550 ( .A(n190), .B(n2900), .Z(n2902) );
  XOR U3551 ( .A(b[19]), .B(a[16]), .Z(n3016) );
  NAND U3552 ( .A(n37821), .B(n3016), .Z(n2901) );
  NAND U3553 ( .A(n2902), .B(n2901), .Z(n3052) );
  XOR U3554 ( .A(n3053), .B(n3052), .Z(n3055) );
  XNOR U3555 ( .A(n3054), .B(n3055), .Z(n3094) );
  XNOR U3556 ( .A(n3095), .B(n3094), .Z(n3096) );
  NANDN U3557 ( .A(n2904), .B(n2903), .Z(n2908) );
  OR U3558 ( .A(n2906), .B(n2905), .Z(n2907) );
  NAND U3559 ( .A(n2908), .B(n2907), .Z(n3097) );
  XOR U3560 ( .A(n3096), .B(n3097), .Z(n2999) );
  XOR U3561 ( .A(n2998), .B(n2999), .Z(n3001) );
  XOR U3562 ( .A(n3000), .B(n3001), .Z(n3115) );
  NANDN U3563 ( .A(n2910), .B(n2909), .Z(n2914) );
  NANDN U3564 ( .A(n2912), .B(n2911), .Z(n2913) );
  AND U3565 ( .A(n2914), .B(n2913), .Z(n3113) );
  NANDN U3566 ( .A(n2916), .B(n2915), .Z(n2920) );
  NANDN U3567 ( .A(n2918), .B(n2917), .Z(n2919) );
  AND U3568 ( .A(n2920), .B(n2919), .Z(n2995) );
  NANDN U3569 ( .A(n2922), .B(n2921), .Z(n2926) );
  OR U3570 ( .A(n2924), .B(n2923), .Z(n2925) );
  AND U3571 ( .A(n2926), .B(n2925), .Z(n2992) );
  NANDN U3572 ( .A(n2928), .B(n2927), .Z(n2932) );
  OR U3573 ( .A(n2930), .B(n2929), .Z(n2931) );
  AND U3574 ( .A(n2932), .B(n2931), .Z(n3101) );
  NANDN U3575 ( .A(n2934), .B(n2933), .Z(n2938) );
  OR U3576 ( .A(n2936), .B(n2935), .Z(n2937) );
  NAND U3577 ( .A(n2938), .B(n2937), .Z(n3100) );
  XNOR U3578 ( .A(n3101), .B(n3100), .Z(n3102) );
  NAND U3579 ( .A(b[0]), .B(a[34]), .Z(n2939) );
  XNOR U3580 ( .A(b[1]), .B(n2939), .Z(n2941) );
  NANDN U3581 ( .A(b[0]), .B(a[33]), .Z(n2940) );
  NAND U3582 ( .A(n2941), .B(n2940), .Z(n3007) );
  NAND U3583 ( .A(n194), .B(n2942), .Z(n2944) );
  XOR U3584 ( .A(b[29]), .B(a[6]), .Z(n3064) );
  NAND U3585 ( .A(n38456), .B(n3064), .Z(n2943) );
  AND U3586 ( .A(n2944), .B(n2943), .Z(n3005) );
  AND U3587 ( .A(b[31]), .B(a[2]), .Z(n3004) );
  XNOR U3588 ( .A(n3005), .B(n3004), .Z(n3006) );
  XNOR U3589 ( .A(n3007), .B(n3006), .Z(n3046) );
  NAND U3590 ( .A(n38185), .B(n2945), .Z(n2947) );
  XOR U3591 ( .A(b[23]), .B(a[12]), .Z(n3070) );
  NAND U3592 ( .A(n38132), .B(n3070), .Z(n2946) );
  AND U3593 ( .A(n2947), .B(n2946), .Z(n3061) );
  NAND U3594 ( .A(n184), .B(n2948), .Z(n2950) );
  XOR U3595 ( .A(b[7]), .B(a[28]), .Z(n3073) );
  NAND U3596 ( .A(n36592), .B(n3073), .Z(n2949) );
  AND U3597 ( .A(n2950), .B(n2949), .Z(n3059) );
  NAND U3598 ( .A(n38289), .B(n2951), .Z(n2953) );
  XOR U3599 ( .A(b[25]), .B(a[10]), .Z(n3076) );
  NAND U3600 ( .A(n38247), .B(n3076), .Z(n2952) );
  NAND U3601 ( .A(n2953), .B(n2952), .Z(n3058) );
  XNOR U3602 ( .A(n3059), .B(n3058), .Z(n3060) );
  XOR U3603 ( .A(n3061), .B(n3060), .Z(n3047) );
  XNOR U3604 ( .A(n3046), .B(n3047), .Z(n3048) );
  NAND U3605 ( .A(n187), .B(n2954), .Z(n2956) );
  XOR U3606 ( .A(b[13]), .B(a[22]), .Z(n3079) );
  NAND U3607 ( .A(n37295), .B(n3079), .Z(n2955) );
  AND U3608 ( .A(n2956), .B(n2955), .Z(n3041) );
  NAND U3609 ( .A(n186), .B(n2957), .Z(n2959) );
  XOR U3610 ( .A(b[11]), .B(a[24]), .Z(n3082) );
  NAND U3611 ( .A(n37097), .B(n3082), .Z(n2958) );
  NAND U3612 ( .A(n2959), .B(n2958), .Z(n3040) );
  XNOR U3613 ( .A(n3041), .B(n3040), .Z(n3042) );
  NAND U3614 ( .A(n188), .B(n2960), .Z(n2962) );
  XOR U3615 ( .A(b[15]), .B(a[20]), .Z(n3085) );
  NAND U3616 ( .A(n37382), .B(n3085), .Z(n2961) );
  AND U3617 ( .A(n2962), .B(n2961), .Z(n3037) );
  NAND U3618 ( .A(n38064), .B(n2963), .Z(n2965) );
  XOR U3619 ( .A(b[21]), .B(a[14]), .Z(n3088) );
  NAND U3620 ( .A(n37993), .B(n3088), .Z(n2964) );
  AND U3621 ( .A(n2965), .B(n2964), .Z(n3035) );
  NAND U3622 ( .A(n185), .B(n2966), .Z(n2968) );
  XOR U3623 ( .A(b[9]), .B(a[26]), .Z(n3091) );
  NAND U3624 ( .A(n36805), .B(n3091), .Z(n2967) );
  NAND U3625 ( .A(n2968), .B(n2967), .Z(n3034) );
  XNOR U3626 ( .A(n3035), .B(n3034), .Z(n3036) );
  XOR U3627 ( .A(n3037), .B(n3036), .Z(n3043) );
  XOR U3628 ( .A(n3042), .B(n3043), .Z(n3049) );
  XOR U3629 ( .A(n3048), .B(n3049), .Z(n3103) );
  XOR U3630 ( .A(n3102), .B(n3103), .Z(n2993) );
  XNOR U3631 ( .A(n2992), .B(n2993), .Z(n2994) );
  XNOR U3632 ( .A(n2995), .B(n2994), .Z(n3112) );
  XNOR U3633 ( .A(n3113), .B(n3112), .Z(n3114) );
  XNOR U3634 ( .A(n3115), .B(n3114), .Z(n3120) );
  XOR U3635 ( .A(n3121), .B(n3120), .Z(n2987) );
  NANDN U3636 ( .A(n2970), .B(n2969), .Z(n2974) );
  NANDN U3637 ( .A(n2972), .B(n2971), .Z(n2973) );
  NAND U3638 ( .A(n2974), .B(n2973), .Z(n2986) );
  XNOR U3639 ( .A(n2987), .B(n2986), .Z(n2988) );
  XNOR U3640 ( .A(n2989), .B(n2988), .Z(n2980) );
  XNOR U3641 ( .A(n2981), .B(n2980), .Z(n2982) );
  XNOR U3642 ( .A(n2983), .B(n2982), .Z(n3124) );
  XNOR U3643 ( .A(sreg[258]), .B(n3124), .Z(n3126) );
  NANDN U3644 ( .A(sreg[257]), .B(n2975), .Z(n2979) );
  NAND U3645 ( .A(n2977), .B(n2976), .Z(n2978) );
  NAND U3646 ( .A(n2979), .B(n2978), .Z(n3125) );
  XNOR U3647 ( .A(n3126), .B(n3125), .Z(c[258]) );
  NANDN U3648 ( .A(n2981), .B(n2980), .Z(n2985) );
  NANDN U3649 ( .A(n2983), .B(n2982), .Z(n2984) );
  AND U3650 ( .A(n2985), .B(n2984), .Z(n3136) );
  NANDN U3651 ( .A(n2987), .B(n2986), .Z(n2991) );
  NANDN U3652 ( .A(n2989), .B(n2988), .Z(n2990) );
  AND U3653 ( .A(n2991), .B(n2990), .Z(n3135) );
  NANDN U3654 ( .A(n2993), .B(n2992), .Z(n2997) );
  NANDN U3655 ( .A(n2995), .B(n2994), .Z(n2996) );
  AND U3656 ( .A(n2997), .B(n2996), .Z(n3273) );
  NANDN U3657 ( .A(n2999), .B(n2998), .Z(n3003) );
  OR U3658 ( .A(n3001), .B(n3000), .Z(n3002) );
  AND U3659 ( .A(n3003), .B(n3002), .Z(n3272) );
  XNOR U3660 ( .A(n3273), .B(n3272), .Z(n3275) );
  NANDN U3661 ( .A(n3005), .B(n3004), .Z(n3009) );
  NANDN U3662 ( .A(n3007), .B(n3006), .Z(n3008) );
  AND U3663 ( .A(n3009), .B(n3008), .Z(n3220) );
  NAND U3664 ( .A(n38385), .B(n3010), .Z(n3012) );
  XOR U3665 ( .A(b[27]), .B(a[9]), .Z(n3164) );
  NAND U3666 ( .A(n38343), .B(n3164), .Z(n3011) );
  AND U3667 ( .A(n3012), .B(n3011), .Z(n3227) );
  NAND U3668 ( .A(n183), .B(n3013), .Z(n3015) );
  XOR U3669 ( .A(b[5]), .B(a[31]), .Z(n3167) );
  NAND U3670 ( .A(n36296), .B(n3167), .Z(n3014) );
  AND U3671 ( .A(n3015), .B(n3014), .Z(n3225) );
  NAND U3672 ( .A(n190), .B(n3016), .Z(n3018) );
  XOR U3673 ( .A(b[19]), .B(a[17]), .Z(n3170) );
  NAND U3674 ( .A(n37821), .B(n3170), .Z(n3017) );
  NAND U3675 ( .A(n3018), .B(n3017), .Z(n3224) );
  XNOR U3676 ( .A(n3225), .B(n3224), .Z(n3226) );
  XNOR U3677 ( .A(n3227), .B(n3226), .Z(n3218) );
  NAND U3678 ( .A(n38470), .B(n3019), .Z(n3021) );
  XOR U3679 ( .A(b[31]), .B(a[5]), .Z(n3173) );
  NAND U3680 ( .A(n38453), .B(n3173), .Z(n3020) );
  AND U3681 ( .A(n3021), .B(n3020), .Z(n3185) );
  NAND U3682 ( .A(n181), .B(n3022), .Z(n3024) );
  XOR U3683 ( .A(b[3]), .B(a[33]), .Z(n3176) );
  NAND U3684 ( .A(n182), .B(n3176), .Z(n3023) );
  AND U3685 ( .A(n3024), .B(n3023), .Z(n3183) );
  NAND U3686 ( .A(n189), .B(n3025), .Z(n3027) );
  XOR U3687 ( .A(b[17]), .B(a[19]), .Z(n3179) );
  NAND U3688 ( .A(n37652), .B(n3179), .Z(n3026) );
  NAND U3689 ( .A(n3027), .B(n3026), .Z(n3182) );
  XNOR U3690 ( .A(n3183), .B(n3182), .Z(n3184) );
  XOR U3691 ( .A(n3185), .B(n3184), .Z(n3219) );
  XOR U3692 ( .A(n3218), .B(n3219), .Z(n3221) );
  XOR U3693 ( .A(n3220), .B(n3221), .Z(n3147) );
  NANDN U3694 ( .A(n3029), .B(n3028), .Z(n3033) );
  OR U3695 ( .A(n3031), .B(n3030), .Z(n3032) );
  AND U3696 ( .A(n3033), .B(n3032), .Z(n3206) );
  NANDN U3697 ( .A(n3035), .B(n3034), .Z(n3039) );
  NANDN U3698 ( .A(n3037), .B(n3036), .Z(n3038) );
  NAND U3699 ( .A(n3039), .B(n3038), .Z(n3207) );
  XNOR U3700 ( .A(n3206), .B(n3207), .Z(n3208) );
  NANDN U3701 ( .A(n3041), .B(n3040), .Z(n3045) );
  NANDN U3702 ( .A(n3043), .B(n3042), .Z(n3044) );
  NAND U3703 ( .A(n3045), .B(n3044), .Z(n3209) );
  XNOR U3704 ( .A(n3208), .B(n3209), .Z(n3146) );
  XNOR U3705 ( .A(n3147), .B(n3146), .Z(n3149) );
  NANDN U3706 ( .A(n3047), .B(n3046), .Z(n3051) );
  NANDN U3707 ( .A(n3049), .B(n3048), .Z(n3050) );
  AND U3708 ( .A(n3051), .B(n3050), .Z(n3148) );
  XOR U3709 ( .A(n3149), .B(n3148), .Z(n3269) );
  NANDN U3710 ( .A(n3053), .B(n3052), .Z(n3057) );
  OR U3711 ( .A(n3055), .B(n3054), .Z(n3056) );
  AND U3712 ( .A(n3057), .B(n3056), .Z(n3213) );
  NANDN U3713 ( .A(n3059), .B(n3058), .Z(n3063) );
  NANDN U3714 ( .A(n3061), .B(n3060), .Z(n3062) );
  NAND U3715 ( .A(n3063), .B(n3062), .Z(n3212) );
  XNOR U3716 ( .A(n3213), .B(n3212), .Z(n3215) );
  NAND U3717 ( .A(n194), .B(n3064), .Z(n3066) );
  XOR U3718 ( .A(b[29]), .B(a[7]), .Z(n3239) );
  NAND U3719 ( .A(n38456), .B(n3239), .Z(n3065) );
  AND U3720 ( .A(n3066), .B(n3065), .Z(n3159) );
  AND U3721 ( .A(b[31]), .B(a[3]), .Z(n3158) );
  XNOR U3722 ( .A(n3159), .B(n3158), .Z(n3160) );
  NAND U3723 ( .A(b[0]), .B(a[35]), .Z(n3067) );
  XNOR U3724 ( .A(b[1]), .B(n3067), .Z(n3069) );
  NANDN U3725 ( .A(b[0]), .B(a[34]), .Z(n3068) );
  NAND U3726 ( .A(n3069), .B(n3068), .Z(n3161) );
  XNOR U3727 ( .A(n3160), .B(n3161), .Z(n3200) );
  NAND U3728 ( .A(n38185), .B(n3070), .Z(n3072) );
  XOR U3729 ( .A(b[23]), .B(a[13]), .Z(n3242) );
  NAND U3730 ( .A(n38132), .B(n3242), .Z(n3071) );
  AND U3731 ( .A(n3072), .B(n3071), .Z(n3233) );
  NAND U3732 ( .A(n184), .B(n3073), .Z(n3075) );
  XOR U3733 ( .A(b[7]), .B(a[29]), .Z(n3245) );
  NAND U3734 ( .A(n36592), .B(n3245), .Z(n3074) );
  AND U3735 ( .A(n3075), .B(n3074), .Z(n3231) );
  NAND U3736 ( .A(n38289), .B(n3076), .Z(n3078) );
  XOR U3737 ( .A(b[25]), .B(a[11]), .Z(n3248) );
  NAND U3738 ( .A(n38247), .B(n3248), .Z(n3077) );
  NAND U3739 ( .A(n3078), .B(n3077), .Z(n3230) );
  XNOR U3740 ( .A(n3231), .B(n3230), .Z(n3232) );
  XOR U3741 ( .A(n3233), .B(n3232), .Z(n3201) );
  XNOR U3742 ( .A(n3200), .B(n3201), .Z(n3202) );
  NAND U3743 ( .A(n187), .B(n3079), .Z(n3081) );
  XOR U3744 ( .A(b[13]), .B(a[23]), .Z(n3251) );
  NAND U3745 ( .A(n37295), .B(n3251), .Z(n3080) );
  AND U3746 ( .A(n3081), .B(n3080), .Z(n3195) );
  NAND U3747 ( .A(n186), .B(n3082), .Z(n3084) );
  XOR U3748 ( .A(b[11]), .B(a[25]), .Z(n3254) );
  NAND U3749 ( .A(n37097), .B(n3254), .Z(n3083) );
  NAND U3750 ( .A(n3084), .B(n3083), .Z(n3194) );
  XNOR U3751 ( .A(n3195), .B(n3194), .Z(n3196) );
  NAND U3752 ( .A(n188), .B(n3085), .Z(n3087) );
  XOR U3753 ( .A(b[15]), .B(a[21]), .Z(n3257) );
  NAND U3754 ( .A(n37382), .B(n3257), .Z(n3086) );
  AND U3755 ( .A(n3087), .B(n3086), .Z(n3191) );
  NAND U3756 ( .A(n38064), .B(n3088), .Z(n3090) );
  XOR U3757 ( .A(b[21]), .B(a[15]), .Z(n3260) );
  NAND U3758 ( .A(n37993), .B(n3260), .Z(n3089) );
  AND U3759 ( .A(n3090), .B(n3089), .Z(n3189) );
  NAND U3760 ( .A(n185), .B(n3091), .Z(n3093) );
  XOR U3761 ( .A(b[9]), .B(a[27]), .Z(n3263) );
  NAND U3762 ( .A(n36805), .B(n3263), .Z(n3092) );
  NAND U3763 ( .A(n3093), .B(n3092), .Z(n3188) );
  XNOR U3764 ( .A(n3189), .B(n3188), .Z(n3190) );
  XOR U3765 ( .A(n3191), .B(n3190), .Z(n3197) );
  XOR U3766 ( .A(n3196), .B(n3197), .Z(n3203) );
  XNOR U3767 ( .A(n3202), .B(n3203), .Z(n3214) );
  XOR U3768 ( .A(n3215), .B(n3214), .Z(n3153) );
  NANDN U3769 ( .A(n3095), .B(n3094), .Z(n3099) );
  NANDN U3770 ( .A(n3097), .B(n3096), .Z(n3098) );
  NAND U3771 ( .A(n3099), .B(n3098), .Z(n3152) );
  XNOR U3772 ( .A(n3153), .B(n3152), .Z(n3155) );
  NANDN U3773 ( .A(n3101), .B(n3100), .Z(n3105) );
  NANDN U3774 ( .A(n3103), .B(n3102), .Z(n3104) );
  AND U3775 ( .A(n3105), .B(n3104), .Z(n3154) );
  XOR U3776 ( .A(n3155), .B(n3154), .Z(n3267) );
  NANDN U3777 ( .A(n3107), .B(n3106), .Z(n3111) );
  NANDN U3778 ( .A(n3109), .B(n3108), .Z(n3110) );
  AND U3779 ( .A(n3111), .B(n3110), .Z(n3266) );
  XNOR U3780 ( .A(n3267), .B(n3266), .Z(n3268) );
  XNOR U3781 ( .A(n3269), .B(n3268), .Z(n3274) );
  XOR U3782 ( .A(n3275), .B(n3274), .Z(n3141) );
  NANDN U3783 ( .A(n3113), .B(n3112), .Z(n3117) );
  NANDN U3784 ( .A(n3115), .B(n3114), .Z(n3116) );
  AND U3785 ( .A(n3117), .B(n3116), .Z(n3140) );
  XNOR U3786 ( .A(n3141), .B(n3140), .Z(n3142) );
  NANDN U3787 ( .A(n3119), .B(n3118), .Z(n3123) );
  NAND U3788 ( .A(n3121), .B(n3120), .Z(n3122) );
  NAND U3789 ( .A(n3123), .B(n3122), .Z(n3143) );
  XNOR U3790 ( .A(n3142), .B(n3143), .Z(n3134) );
  XOR U3791 ( .A(n3135), .B(n3134), .Z(n3137) );
  XOR U3792 ( .A(n3136), .B(n3137), .Z(n3129) );
  XNOR U3793 ( .A(n3129), .B(sreg[259]), .Z(n3131) );
  NANDN U3794 ( .A(sreg[258]), .B(n3124), .Z(n3128) );
  NAND U3795 ( .A(n3126), .B(n3125), .Z(n3127) );
  AND U3796 ( .A(n3128), .B(n3127), .Z(n3130) );
  XOR U3797 ( .A(n3131), .B(n3130), .Z(c[259]) );
  NANDN U3798 ( .A(n3129), .B(sreg[259]), .Z(n3133) );
  NAND U3799 ( .A(n3131), .B(n3130), .Z(n3132) );
  AND U3800 ( .A(n3133), .B(n3132), .Z(n3422) );
  NANDN U3801 ( .A(n3135), .B(n3134), .Z(n3139) );
  OR U3802 ( .A(n3137), .B(n3136), .Z(n3138) );
  AND U3803 ( .A(n3139), .B(n3138), .Z(n3281) );
  NANDN U3804 ( .A(n3141), .B(n3140), .Z(n3145) );
  NANDN U3805 ( .A(n3143), .B(n3142), .Z(n3144) );
  AND U3806 ( .A(n3145), .B(n3144), .Z(n3279) );
  NANDN U3807 ( .A(n3147), .B(n3146), .Z(n3151) );
  NAND U3808 ( .A(n3149), .B(n3148), .Z(n3150) );
  AND U3809 ( .A(n3151), .B(n3150), .Z(n3414) );
  NANDN U3810 ( .A(n3153), .B(n3152), .Z(n3157) );
  NAND U3811 ( .A(n3155), .B(n3154), .Z(n3156) );
  NAND U3812 ( .A(n3157), .B(n3156), .Z(n3415) );
  XNOR U3813 ( .A(n3414), .B(n3415), .Z(n3417) );
  NANDN U3814 ( .A(n3159), .B(n3158), .Z(n3163) );
  NANDN U3815 ( .A(n3161), .B(n3160), .Z(n3162) );
  AND U3816 ( .A(n3163), .B(n3162), .Z(n3362) );
  NAND U3817 ( .A(n38385), .B(n3164), .Z(n3166) );
  XOR U3818 ( .A(b[27]), .B(a[10]), .Z(n3308) );
  NAND U3819 ( .A(n38343), .B(n3308), .Z(n3165) );
  AND U3820 ( .A(n3166), .B(n3165), .Z(n3369) );
  NAND U3821 ( .A(n183), .B(n3167), .Z(n3169) );
  XOR U3822 ( .A(b[5]), .B(a[32]), .Z(n3311) );
  NAND U3823 ( .A(n36296), .B(n3311), .Z(n3168) );
  AND U3824 ( .A(n3169), .B(n3168), .Z(n3367) );
  NAND U3825 ( .A(n190), .B(n3170), .Z(n3172) );
  XOR U3826 ( .A(b[19]), .B(a[18]), .Z(n3314) );
  NAND U3827 ( .A(n37821), .B(n3314), .Z(n3171) );
  NAND U3828 ( .A(n3172), .B(n3171), .Z(n3366) );
  XNOR U3829 ( .A(n3367), .B(n3366), .Z(n3368) );
  XNOR U3830 ( .A(n3369), .B(n3368), .Z(n3360) );
  NAND U3831 ( .A(n38470), .B(n3173), .Z(n3175) );
  XOR U3832 ( .A(b[31]), .B(a[6]), .Z(n3317) );
  NAND U3833 ( .A(n38453), .B(n3317), .Z(n3174) );
  AND U3834 ( .A(n3175), .B(n3174), .Z(n3329) );
  NAND U3835 ( .A(n181), .B(n3176), .Z(n3178) );
  XOR U3836 ( .A(b[3]), .B(a[34]), .Z(n3320) );
  NAND U3837 ( .A(n182), .B(n3320), .Z(n3177) );
  AND U3838 ( .A(n3178), .B(n3177), .Z(n3327) );
  NAND U3839 ( .A(n189), .B(n3179), .Z(n3181) );
  XOR U3840 ( .A(b[17]), .B(a[20]), .Z(n3323) );
  NAND U3841 ( .A(n37652), .B(n3323), .Z(n3180) );
  NAND U3842 ( .A(n3181), .B(n3180), .Z(n3326) );
  XNOR U3843 ( .A(n3327), .B(n3326), .Z(n3328) );
  XOR U3844 ( .A(n3329), .B(n3328), .Z(n3361) );
  XOR U3845 ( .A(n3360), .B(n3361), .Z(n3363) );
  XOR U3846 ( .A(n3362), .B(n3363), .Z(n3297) );
  NANDN U3847 ( .A(n3183), .B(n3182), .Z(n3187) );
  NANDN U3848 ( .A(n3185), .B(n3184), .Z(n3186) );
  AND U3849 ( .A(n3187), .B(n3186), .Z(n3350) );
  NANDN U3850 ( .A(n3189), .B(n3188), .Z(n3193) );
  NANDN U3851 ( .A(n3191), .B(n3190), .Z(n3192) );
  NAND U3852 ( .A(n3193), .B(n3192), .Z(n3351) );
  XNOR U3853 ( .A(n3350), .B(n3351), .Z(n3352) );
  NANDN U3854 ( .A(n3195), .B(n3194), .Z(n3199) );
  NANDN U3855 ( .A(n3197), .B(n3196), .Z(n3198) );
  NAND U3856 ( .A(n3199), .B(n3198), .Z(n3353) );
  XNOR U3857 ( .A(n3352), .B(n3353), .Z(n3296) );
  XNOR U3858 ( .A(n3297), .B(n3296), .Z(n3299) );
  NANDN U3859 ( .A(n3201), .B(n3200), .Z(n3205) );
  NANDN U3860 ( .A(n3203), .B(n3202), .Z(n3204) );
  AND U3861 ( .A(n3205), .B(n3204), .Z(n3298) );
  XOR U3862 ( .A(n3299), .B(n3298), .Z(n3411) );
  NANDN U3863 ( .A(n3207), .B(n3206), .Z(n3211) );
  NANDN U3864 ( .A(n3209), .B(n3208), .Z(n3210) );
  AND U3865 ( .A(n3211), .B(n3210), .Z(n3408) );
  NANDN U3866 ( .A(n3213), .B(n3212), .Z(n3217) );
  NAND U3867 ( .A(n3215), .B(n3214), .Z(n3216) );
  AND U3868 ( .A(n3217), .B(n3216), .Z(n3293) );
  NANDN U3869 ( .A(n3219), .B(n3218), .Z(n3223) );
  OR U3870 ( .A(n3221), .B(n3220), .Z(n3222) );
  AND U3871 ( .A(n3223), .B(n3222), .Z(n3291) );
  NANDN U3872 ( .A(n3225), .B(n3224), .Z(n3229) );
  NANDN U3873 ( .A(n3227), .B(n3226), .Z(n3228) );
  AND U3874 ( .A(n3229), .B(n3228), .Z(n3357) );
  NANDN U3875 ( .A(n3231), .B(n3230), .Z(n3235) );
  NANDN U3876 ( .A(n3233), .B(n3232), .Z(n3234) );
  NAND U3877 ( .A(n3235), .B(n3234), .Z(n3356) );
  XNOR U3878 ( .A(n3357), .B(n3356), .Z(n3359) );
  NAND U3879 ( .A(b[0]), .B(a[36]), .Z(n3236) );
  XNOR U3880 ( .A(b[1]), .B(n3236), .Z(n3238) );
  NANDN U3881 ( .A(b[0]), .B(a[35]), .Z(n3237) );
  NAND U3882 ( .A(n3238), .B(n3237), .Z(n3305) );
  NAND U3883 ( .A(n194), .B(n3239), .Z(n3241) );
  XOR U3884 ( .A(b[29]), .B(a[8]), .Z(n3378) );
  NAND U3885 ( .A(n38456), .B(n3378), .Z(n3240) );
  AND U3886 ( .A(n3241), .B(n3240), .Z(n3303) );
  AND U3887 ( .A(b[31]), .B(a[4]), .Z(n3302) );
  XNOR U3888 ( .A(n3303), .B(n3302), .Z(n3304) );
  XNOR U3889 ( .A(n3305), .B(n3304), .Z(n3345) );
  NAND U3890 ( .A(n38185), .B(n3242), .Z(n3244) );
  XOR U3891 ( .A(b[23]), .B(a[14]), .Z(n3384) );
  NAND U3892 ( .A(n38132), .B(n3384), .Z(n3243) );
  AND U3893 ( .A(n3244), .B(n3243), .Z(n3374) );
  NAND U3894 ( .A(n184), .B(n3245), .Z(n3247) );
  XOR U3895 ( .A(b[7]), .B(a[30]), .Z(n3387) );
  NAND U3896 ( .A(n36592), .B(n3387), .Z(n3246) );
  AND U3897 ( .A(n3247), .B(n3246), .Z(n3373) );
  NAND U3898 ( .A(n38289), .B(n3248), .Z(n3250) );
  XOR U3899 ( .A(b[25]), .B(a[12]), .Z(n3390) );
  NAND U3900 ( .A(n38247), .B(n3390), .Z(n3249) );
  NAND U3901 ( .A(n3250), .B(n3249), .Z(n3372) );
  XOR U3902 ( .A(n3373), .B(n3372), .Z(n3375) );
  XOR U3903 ( .A(n3374), .B(n3375), .Z(n3344) );
  XOR U3904 ( .A(n3345), .B(n3344), .Z(n3347) );
  NAND U3905 ( .A(n187), .B(n3251), .Z(n3253) );
  XOR U3906 ( .A(b[13]), .B(a[24]), .Z(n3393) );
  NAND U3907 ( .A(n37295), .B(n3393), .Z(n3252) );
  AND U3908 ( .A(n3253), .B(n3252), .Z(n3339) );
  NAND U3909 ( .A(n186), .B(n3254), .Z(n3256) );
  XOR U3910 ( .A(b[11]), .B(a[26]), .Z(n3396) );
  NAND U3911 ( .A(n37097), .B(n3396), .Z(n3255) );
  NAND U3912 ( .A(n3256), .B(n3255), .Z(n3338) );
  XNOR U3913 ( .A(n3339), .B(n3338), .Z(n3341) );
  NAND U3914 ( .A(n188), .B(n3257), .Z(n3259) );
  XOR U3915 ( .A(b[15]), .B(a[22]), .Z(n3399) );
  NAND U3916 ( .A(n37382), .B(n3399), .Z(n3258) );
  AND U3917 ( .A(n3259), .B(n3258), .Z(n3335) );
  NAND U3918 ( .A(n38064), .B(n3260), .Z(n3262) );
  XOR U3919 ( .A(b[21]), .B(a[16]), .Z(n3402) );
  NAND U3920 ( .A(n37993), .B(n3402), .Z(n3261) );
  AND U3921 ( .A(n3262), .B(n3261), .Z(n3333) );
  NAND U3922 ( .A(n185), .B(n3263), .Z(n3265) );
  XOR U3923 ( .A(b[9]), .B(a[28]), .Z(n3405) );
  NAND U3924 ( .A(n36805), .B(n3405), .Z(n3264) );
  NAND U3925 ( .A(n3265), .B(n3264), .Z(n3332) );
  XNOR U3926 ( .A(n3333), .B(n3332), .Z(n3334) );
  XNOR U3927 ( .A(n3335), .B(n3334), .Z(n3340) );
  XOR U3928 ( .A(n3341), .B(n3340), .Z(n3346) );
  XNOR U3929 ( .A(n3347), .B(n3346), .Z(n3358) );
  XNOR U3930 ( .A(n3359), .B(n3358), .Z(n3290) );
  XNOR U3931 ( .A(n3291), .B(n3290), .Z(n3292) );
  XOR U3932 ( .A(n3293), .B(n3292), .Z(n3409) );
  XNOR U3933 ( .A(n3408), .B(n3409), .Z(n3410) );
  XNOR U3934 ( .A(n3411), .B(n3410), .Z(n3416) );
  XOR U3935 ( .A(n3417), .B(n3416), .Z(n3285) );
  NANDN U3936 ( .A(n3267), .B(n3266), .Z(n3271) );
  NANDN U3937 ( .A(n3269), .B(n3268), .Z(n3270) );
  AND U3938 ( .A(n3271), .B(n3270), .Z(n3284) );
  XNOR U3939 ( .A(n3285), .B(n3284), .Z(n3286) );
  NANDN U3940 ( .A(n3273), .B(n3272), .Z(n3277) );
  NAND U3941 ( .A(n3275), .B(n3274), .Z(n3276) );
  NAND U3942 ( .A(n3277), .B(n3276), .Z(n3287) );
  XNOR U3943 ( .A(n3286), .B(n3287), .Z(n3278) );
  XNOR U3944 ( .A(n3279), .B(n3278), .Z(n3280) );
  XNOR U3945 ( .A(n3281), .B(n3280), .Z(n3420) );
  XNOR U3946 ( .A(sreg[260]), .B(n3420), .Z(n3421) );
  XNOR U3947 ( .A(n3422), .B(n3421), .Z(c[260]) );
  NANDN U3948 ( .A(n3279), .B(n3278), .Z(n3283) );
  NANDN U3949 ( .A(n3281), .B(n3280), .Z(n3282) );
  AND U3950 ( .A(n3283), .B(n3282), .Z(n3428) );
  NANDN U3951 ( .A(n3285), .B(n3284), .Z(n3289) );
  NANDN U3952 ( .A(n3287), .B(n3286), .Z(n3288) );
  AND U3953 ( .A(n3289), .B(n3288), .Z(n3426) );
  NANDN U3954 ( .A(n3291), .B(n3290), .Z(n3295) );
  NANDN U3955 ( .A(n3293), .B(n3292), .Z(n3294) );
  AND U3956 ( .A(n3295), .B(n3294), .Z(n3562) );
  NANDN U3957 ( .A(n3297), .B(n3296), .Z(n3301) );
  NAND U3958 ( .A(n3299), .B(n3298), .Z(n3300) );
  AND U3959 ( .A(n3301), .B(n3300), .Z(n3561) );
  XNOR U3960 ( .A(n3562), .B(n3561), .Z(n3564) );
  NANDN U3961 ( .A(n3303), .B(n3302), .Z(n3307) );
  NANDN U3962 ( .A(n3305), .B(n3304), .Z(n3306) );
  AND U3963 ( .A(n3307), .B(n3306), .Z(n3497) );
  NAND U3964 ( .A(n38385), .B(n3308), .Z(n3310) );
  XOR U3965 ( .A(b[27]), .B(a[11]), .Z(n3443) );
  NAND U3966 ( .A(n38343), .B(n3443), .Z(n3309) );
  AND U3967 ( .A(n3310), .B(n3309), .Z(n3504) );
  NAND U3968 ( .A(n183), .B(n3311), .Z(n3313) );
  XOR U3969 ( .A(b[5]), .B(a[33]), .Z(n3446) );
  NAND U3970 ( .A(n36296), .B(n3446), .Z(n3312) );
  AND U3971 ( .A(n3313), .B(n3312), .Z(n3502) );
  NAND U3972 ( .A(n190), .B(n3314), .Z(n3316) );
  XOR U3973 ( .A(b[19]), .B(a[19]), .Z(n3449) );
  NAND U3974 ( .A(n37821), .B(n3449), .Z(n3315) );
  NAND U3975 ( .A(n3316), .B(n3315), .Z(n3501) );
  XNOR U3976 ( .A(n3502), .B(n3501), .Z(n3503) );
  XNOR U3977 ( .A(n3504), .B(n3503), .Z(n3495) );
  NAND U3978 ( .A(n38470), .B(n3317), .Z(n3319) );
  XOR U3979 ( .A(b[31]), .B(a[7]), .Z(n3452) );
  NAND U3980 ( .A(n38453), .B(n3452), .Z(n3318) );
  AND U3981 ( .A(n3319), .B(n3318), .Z(n3464) );
  NAND U3982 ( .A(n181), .B(n3320), .Z(n3322) );
  XOR U3983 ( .A(b[3]), .B(a[35]), .Z(n3455) );
  NAND U3984 ( .A(n182), .B(n3455), .Z(n3321) );
  AND U3985 ( .A(n3322), .B(n3321), .Z(n3462) );
  NAND U3986 ( .A(n189), .B(n3323), .Z(n3325) );
  XOR U3987 ( .A(b[17]), .B(a[21]), .Z(n3458) );
  NAND U3988 ( .A(n37652), .B(n3458), .Z(n3324) );
  NAND U3989 ( .A(n3325), .B(n3324), .Z(n3461) );
  XNOR U3990 ( .A(n3462), .B(n3461), .Z(n3463) );
  XOR U3991 ( .A(n3464), .B(n3463), .Z(n3496) );
  XOR U3992 ( .A(n3495), .B(n3496), .Z(n3498) );
  XOR U3993 ( .A(n3497), .B(n3498), .Z(n3544) );
  NANDN U3994 ( .A(n3327), .B(n3326), .Z(n3331) );
  NANDN U3995 ( .A(n3329), .B(n3328), .Z(n3330) );
  AND U3996 ( .A(n3331), .B(n3330), .Z(n3485) );
  NANDN U3997 ( .A(n3333), .B(n3332), .Z(n3337) );
  NANDN U3998 ( .A(n3335), .B(n3334), .Z(n3336) );
  NAND U3999 ( .A(n3337), .B(n3336), .Z(n3486) );
  XNOR U4000 ( .A(n3485), .B(n3486), .Z(n3487) );
  NANDN U4001 ( .A(n3339), .B(n3338), .Z(n3343) );
  NAND U4002 ( .A(n3341), .B(n3340), .Z(n3342) );
  NAND U4003 ( .A(n3343), .B(n3342), .Z(n3488) );
  XNOR U4004 ( .A(n3487), .B(n3488), .Z(n3543) );
  XNOR U4005 ( .A(n3544), .B(n3543), .Z(n3546) );
  NAND U4006 ( .A(n3345), .B(n3344), .Z(n3349) );
  NAND U4007 ( .A(n3347), .B(n3346), .Z(n3348) );
  AND U4008 ( .A(n3349), .B(n3348), .Z(n3545) );
  XOR U4009 ( .A(n3546), .B(n3545), .Z(n3558) );
  NANDN U4010 ( .A(n3351), .B(n3350), .Z(n3355) );
  NANDN U4011 ( .A(n3353), .B(n3352), .Z(n3354) );
  AND U4012 ( .A(n3355), .B(n3354), .Z(n3555) );
  NANDN U4013 ( .A(n3361), .B(n3360), .Z(n3365) );
  OR U4014 ( .A(n3363), .B(n3362), .Z(n3364) );
  AND U4015 ( .A(n3365), .B(n3364), .Z(n3550) );
  NANDN U4016 ( .A(n3367), .B(n3366), .Z(n3371) );
  NANDN U4017 ( .A(n3369), .B(n3368), .Z(n3370) );
  AND U4018 ( .A(n3371), .B(n3370), .Z(n3492) );
  NANDN U4019 ( .A(n3373), .B(n3372), .Z(n3377) );
  OR U4020 ( .A(n3375), .B(n3374), .Z(n3376) );
  NAND U4021 ( .A(n3377), .B(n3376), .Z(n3491) );
  XNOR U4022 ( .A(n3492), .B(n3491), .Z(n3494) );
  NAND U4023 ( .A(n194), .B(n3378), .Z(n3380) );
  XOR U4024 ( .A(b[29]), .B(a[9]), .Z(n3516) );
  NAND U4025 ( .A(n38456), .B(n3516), .Z(n3379) );
  AND U4026 ( .A(n3380), .B(n3379), .Z(n3438) );
  AND U4027 ( .A(b[31]), .B(a[5]), .Z(n3437) );
  XNOR U4028 ( .A(n3438), .B(n3437), .Z(n3439) );
  NAND U4029 ( .A(b[0]), .B(a[37]), .Z(n3381) );
  XNOR U4030 ( .A(b[1]), .B(n3381), .Z(n3383) );
  NANDN U4031 ( .A(b[0]), .B(a[36]), .Z(n3382) );
  NAND U4032 ( .A(n3383), .B(n3382), .Z(n3440) );
  XNOR U4033 ( .A(n3439), .B(n3440), .Z(n3480) );
  NAND U4034 ( .A(n38185), .B(n3384), .Z(n3386) );
  XOR U4035 ( .A(b[23]), .B(a[15]), .Z(n3519) );
  NAND U4036 ( .A(n38132), .B(n3519), .Z(n3385) );
  AND U4037 ( .A(n3386), .B(n3385), .Z(n3509) );
  NAND U4038 ( .A(n184), .B(n3387), .Z(n3389) );
  XOR U4039 ( .A(b[7]), .B(a[31]), .Z(n3522) );
  NAND U4040 ( .A(n36592), .B(n3522), .Z(n3388) );
  AND U4041 ( .A(n3389), .B(n3388), .Z(n3508) );
  NAND U4042 ( .A(n38289), .B(n3390), .Z(n3392) );
  XOR U4043 ( .A(b[25]), .B(a[13]), .Z(n3525) );
  NAND U4044 ( .A(n38247), .B(n3525), .Z(n3391) );
  NAND U4045 ( .A(n3392), .B(n3391), .Z(n3507) );
  XOR U4046 ( .A(n3508), .B(n3507), .Z(n3510) );
  XOR U4047 ( .A(n3509), .B(n3510), .Z(n3479) );
  XOR U4048 ( .A(n3480), .B(n3479), .Z(n3482) );
  NAND U4049 ( .A(n187), .B(n3393), .Z(n3395) );
  XOR U4050 ( .A(b[13]), .B(a[25]), .Z(n3528) );
  NAND U4051 ( .A(n37295), .B(n3528), .Z(n3394) );
  AND U4052 ( .A(n3395), .B(n3394), .Z(n3474) );
  NAND U4053 ( .A(n186), .B(n3396), .Z(n3398) );
  XOR U4054 ( .A(b[11]), .B(a[27]), .Z(n3531) );
  NAND U4055 ( .A(n37097), .B(n3531), .Z(n3397) );
  NAND U4056 ( .A(n3398), .B(n3397), .Z(n3473) );
  XNOR U4057 ( .A(n3474), .B(n3473), .Z(n3476) );
  NAND U4058 ( .A(n188), .B(n3399), .Z(n3401) );
  XOR U4059 ( .A(b[15]), .B(a[23]), .Z(n3534) );
  NAND U4060 ( .A(n37382), .B(n3534), .Z(n3400) );
  AND U4061 ( .A(n3401), .B(n3400), .Z(n3470) );
  NAND U4062 ( .A(n38064), .B(n3402), .Z(n3404) );
  XOR U4063 ( .A(b[21]), .B(a[17]), .Z(n3537) );
  NAND U4064 ( .A(n37993), .B(n3537), .Z(n3403) );
  AND U4065 ( .A(n3404), .B(n3403), .Z(n3468) );
  NAND U4066 ( .A(n185), .B(n3405), .Z(n3407) );
  XOR U4067 ( .A(b[9]), .B(a[29]), .Z(n3540) );
  NAND U4068 ( .A(n36805), .B(n3540), .Z(n3406) );
  NAND U4069 ( .A(n3407), .B(n3406), .Z(n3467) );
  XNOR U4070 ( .A(n3468), .B(n3467), .Z(n3469) );
  XNOR U4071 ( .A(n3470), .B(n3469), .Z(n3475) );
  XOR U4072 ( .A(n3476), .B(n3475), .Z(n3481) );
  XNOR U4073 ( .A(n3482), .B(n3481), .Z(n3493) );
  XNOR U4074 ( .A(n3494), .B(n3493), .Z(n3549) );
  XNOR U4075 ( .A(n3550), .B(n3549), .Z(n3551) );
  XOR U4076 ( .A(n3552), .B(n3551), .Z(n3556) );
  XNOR U4077 ( .A(n3555), .B(n3556), .Z(n3557) );
  XNOR U4078 ( .A(n3558), .B(n3557), .Z(n3563) );
  XOR U4079 ( .A(n3564), .B(n3563), .Z(n3432) );
  NANDN U4080 ( .A(n3409), .B(n3408), .Z(n3413) );
  NANDN U4081 ( .A(n3411), .B(n3410), .Z(n3412) );
  AND U4082 ( .A(n3413), .B(n3412), .Z(n3431) );
  XNOR U4083 ( .A(n3432), .B(n3431), .Z(n3433) );
  NANDN U4084 ( .A(n3415), .B(n3414), .Z(n3419) );
  NAND U4085 ( .A(n3417), .B(n3416), .Z(n3418) );
  NAND U4086 ( .A(n3419), .B(n3418), .Z(n3434) );
  XNOR U4087 ( .A(n3433), .B(n3434), .Z(n3425) );
  XNOR U4088 ( .A(n3426), .B(n3425), .Z(n3427) );
  XNOR U4089 ( .A(n3428), .B(n3427), .Z(n3567) );
  XNOR U4090 ( .A(sreg[261]), .B(n3567), .Z(n3569) );
  NANDN U4091 ( .A(sreg[260]), .B(n3420), .Z(n3424) );
  NAND U4092 ( .A(n3422), .B(n3421), .Z(n3423) );
  NAND U4093 ( .A(n3424), .B(n3423), .Z(n3568) );
  XNOR U4094 ( .A(n3569), .B(n3568), .Z(c[261]) );
  NANDN U4095 ( .A(n3426), .B(n3425), .Z(n3430) );
  NANDN U4096 ( .A(n3428), .B(n3427), .Z(n3429) );
  AND U4097 ( .A(n3430), .B(n3429), .Z(n3575) );
  NANDN U4098 ( .A(n3432), .B(n3431), .Z(n3436) );
  NANDN U4099 ( .A(n3434), .B(n3433), .Z(n3435) );
  AND U4100 ( .A(n3436), .B(n3435), .Z(n3573) );
  NANDN U4101 ( .A(n3438), .B(n3437), .Z(n3442) );
  NANDN U4102 ( .A(n3440), .B(n3439), .Z(n3441) );
  AND U4103 ( .A(n3442), .B(n3441), .Z(n3650) );
  NAND U4104 ( .A(n38385), .B(n3443), .Z(n3445) );
  XOR U4105 ( .A(b[27]), .B(a[12]), .Z(n3596) );
  NAND U4106 ( .A(n38343), .B(n3596), .Z(n3444) );
  AND U4107 ( .A(n3445), .B(n3444), .Z(n3657) );
  NAND U4108 ( .A(n183), .B(n3446), .Z(n3448) );
  XOR U4109 ( .A(b[5]), .B(a[34]), .Z(n3599) );
  NAND U4110 ( .A(n36296), .B(n3599), .Z(n3447) );
  AND U4111 ( .A(n3448), .B(n3447), .Z(n3655) );
  NAND U4112 ( .A(n190), .B(n3449), .Z(n3451) );
  XOR U4113 ( .A(b[19]), .B(a[20]), .Z(n3602) );
  NAND U4114 ( .A(n37821), .B(n3602), .Z(n3450) );
  NAND U4115 ( .A(n3451), .B(n3450), .Z(n3654) );
  XNOR U4116 ( .A(n3655), .B(n3654), .Z(n3656) );
  XNOR U4117 ( .A(n3657), .B(n3656), .Z(n3648) );
  NAND U4118 ( .A(n38470), .B(n3452), .Z(n3454) );
  XOR U4119 ( .A(b[31]), .B(a[8]), .Z(n3605) );
  NAND U4120 ( .A(n38453), .B(n3605), .Z(n3453) );
  AND U4121 ( .A(n3454), .B(n3453), .Z(n3617) );
  NAND U4122 ( .A(n181), .B(n3455), .Z(n3457) );
  XOR U4123 ( .A(b[3]), .B(a[36]), .Z(n3608) );
  NAND U4124 ( .A(n182), .B(n3608), .Z(n3456) );
  AND U4125 ( .A(n3457), .B(n3456), .Z(n3615) );
  NAND U4126 ( .A(n189), .B(n3458), .Z(n3460) );
  XOR U4127 ( .A(b[17]), .B(a[22]), .Z(n3611) );
  NAND U4128 ( .A(n37652), .B(n3611), .Z(n3459) );
  NAND U4129 ( .A(n3460), .B(n3459), .Z(n3614) );
  XNOR U4130 ( .A(n3615), .B(n3614), .Z(n3616) );
  XOR U4131 ( .A(n3617), .B(n3616), .Z(n3649) );
  XOR U4132 ( .A(n3648), .B(n3649), .Z(n3651) );
  XOR U4133 ( .A(n3650), .B(n3651), .Z(n3697) );
  NANDN U4134 ( .A(n3462), .B(n3461), .Z(n3466) );
  NANDN U4135 ( .A(n3464), .B(n3463), .Z(n3465) );
  AND U4136 ( .A(n3466), .B(n3465), .Z(n3638) );
  NANDN U4137 ( .A(n3468), .B(n3467), .Z(n3472) );
  NANDN U4138 ( .A(n3470), .B(n3469), .Z(n3471) );
  NAND U4139 ( .A(n3472), .B(n3471), .Z(n3639) );
  XNOR U4140 ( .A(n3638), .B(n3639), .Z(n3640) );
  NANDN U4141 ( .A(n3474), .B(n3473), .Z(n3478) );
  NAND U4142 ( .A(n3476), .B(n3475), .Z(n3477) );
  NAND U4143 ( .A(n3478), .B(n3477), .Z(n3641) );
  XNOR U4144 ( .A(n3640), .B(n3641), .Z(n3696) );
  XNOR U4145 ( .A(n3697), .B(n3696), .Z(n3699) );
  NAND U4146 ( .A(n3480), .B(n3479), .Z(n3484) );
  NAND U4147 ( .A(n3482), .B(n3481), .Z(n3483) );
  AND U4148 ( .A(n3484), .B(n3483), .Z(n3698) );
  XOR U4149 ( .A(n3699), .B(n3698), .Z(n3710) );
  NANDN U4150 ( .A(n3486), .B(n3485), .Z(n3490) );
  NANDN U4151 ( .A(n3488), .B(n3487), .Z(n3489) );
  AND U4152 ( .A(n3490), .B(n3489), .Z(n3708) );
  NANDN U4153 ( .A(n3496), .B(n3495), .Z(n3500) );
  OR U4154 ( .A(n3498), .B(n3497), .Z(n3499) );
  AND U4155 ( .A(n3500), .B(n3499), .Z(n3703) );
  NANDN U4156 ( .A(n3502), .B(n3501), .Z(n3506) );
  NANDN U4157 ( .A(n3504), .B(n3503), .Z(n3505) );
  AND U4158 ( .A(n3506), .B(n3505), .Z(n3645) );
  NANDN U4159 ( .A(n3508), .B(n3507), .Z(n3512) );
  OR U4160 ( .A(n3510), .B(n3509), .Z(n3511) );
  NAND U4161 ( .A(n3512), .B(n3511), .Z(n3644) );
  XNOR U4162 ( .A(n3645), .B(n3644), .Z(n3647) );
  AND U4163 ( .A(b[0]), .B(a[38]), .Z(n3513) );
  XOR U4164 ( .A(b[1]), .B(n3513), .Z(n3515) );
  NANDN U4165 ( .A(b[0]), .B(a[37]), .Z(n3514) );
  AND U4166 ( .A(n3515), .B(n3514), .Z(n3592) );
  NAND U4167 ( .A(n194), .B(n3516), .Z(n3518) );
  XOR U4168 ( .A(b[29]), .B(a[10]), .Z(n3669) );
  NAND U4169 ( .A(n38456), .B(n3669), .Z(n3517) );
  AND U4170 ( .A(n3518), .B(n3517), .Z(n3591) );
  AND U4171 ( .A(b[31]), .B(a[6]), .Z(n3590) );
  XOR U4172 ( .A(n3591), .B(n3590), .Z(n3593) );
  XNOR U4173 ( .A(n3592), .B(n3593), .Z(n3633) );
  NAND U4174 ( .A(n38185), .B(n3519), .Z(n3521) );
  XOR U4175 ( .A(b[23]), .B(a[16]), .Z(n3672) );
  NAND U4176 ( .A(n38132), .B(n3672), .Z(n3520) );
  AND U4177 ( .A(n3521), .B(n3520), .Z(n3662) );
  NAND U4178 ( .A(n184), .B(n3522), .Z(n3524) );
  XOR U4179 ( .A(b[7]), .B(a[32]), .Z(n3675) );
  NAND U4180 ( .A(n36592), .B(n3675), .Z(n3523) );
  AND U4181 ( .A(n3524), .B(n3523), .Z(n3661) );
  NAND U4182 ( .A(n38289), .B(n3525), .Z(n3527) );
  XOR U4183 ( .A(b[25]), .B(a[14]), .Z(n3678) );
  NAND U4184 ( .A(n38247), .B(n3678), .Z(n3526) );
  NAND U4185 ( .A(n3527), .B(n3526), .Z(n3660) );
  XOR U4186 ( .A(n3661), .B(n3660), .Z(n3663) );
  XOR U4187 ( .A(n3662), .B(n3663), .Z(n3632) );
  XOR U4188 ( .A(n3633), .B(n3632), .Z(n3635) );
  NAND U4189 ( .A(n187), .B(n3528), .Z(n3530) );
  XOR U4190 ( .A(b[13]), .B(a[26]), .Z(n3681) );
  NAND U4191 ( .A(n37295), .B(n3681), .Z(n3529) );
  AND U4192 ( .A(n3530), .B(n3529), .Z(n3627) );
  NAND U4193 ( .A(n186), .B(n3531), .Z(n3533) );
  XOR U4194 ( .A(b[11]), .B(a[28]), .Z(n3684) );
  NAND U4195 ( .A(n37097), .B(n3684), .Z(n3532) );
  NAND U4196 ( .A(n3533), .B(n3532), .Z(n3626) );
  XNOR U4197 ( .A(n3627), .B(n3626), .Z(n3629) );
  NAND U4198 ( .A(n188), .B(n3534), .Z(n3536) );
  XOR U4199 ( .A(b[15]), .B(a[24]), .Z(n3687) );
  NAND U4200 ( .A(n37382), .B(n3687), .Z(n3535) );
  AND U4201 ( .A(n3536), .B(n3535), .Z(n3623) );
  NAND U4202 ( .A(n38064), .B(n3537), .Z(n3539) );
  XOR U4203 ( .A(b[21]), .B(a[18]), .Z(n3690) );
  NAND U4204 ( .A(n37993), .B(n3690), .Z(n3538) );
  AND U4205 ( .A(n3539), .B(n3538), .Z(n3621) );
  NAND U4206 ( .A(n185), .B(n3540), .Z(n3542) );
  XOR U4207 ( .A(b[9]), .B(a[30]), .Z(n3693) );
  NAND U4208 ( .A(n36805), .B(n3693), .Z(n3541) );
  NAND U4209 ( .A(n3542), .B(n3541), .Z(n3620) );
  XNOR U4210 ( .A(n3621), .B(n3620), .Z(n3622) );
  XNOR U4211 ( .A(n3623), .B(n3622), .Z(n3628) );
  XOR U4212 ( .A(n3629), .B(n3628), .Z(n3634) );
  XNOR U4213 ( .A(n3635), .B(n3634), .Z(n3646) );
  XNOR U4214 ( .A(n3647), .B(n3646), .Z(n3702) );
  XNOR U4215 ( .A(n3703), .B(n3702), .Z(n3704) );
  XOR U4216 ( .A(n3705), .B(n3704), .Z(n3709) );
  XOR U4217 ( .A(n3708), .B(n3709), .Z(n3711) );
  XOR U4218 ( .A(n3710), .B(n3711), .Z(n3587) );
  NANDN U4219 ( .A(n3544), .B(n3543), .Z(n3548) );
  NAND U4220 ( .A(n3546), .B(n3545), .Z(n3547) );
  AND U4221 ( .A(n3548), .B(n3547), .Z(n3585) );
  NANDN U4222 ( .A(n3550), .B(n3549), .Z(n3554) );
  NANDN U4223 ( .A(n3552), .B(n3551), .Z(n3553) );
  AND U4224 ( .A(n3554), .B(n3553), .Z(n3584) );
  XNOR U4225 ( .A(n3585), .B(n3584), .Z(n3586) );
  XNOR U4226 ( .A(n3587), .B(n3586), .Z(n3578) );
  NANDN U4227 ( .A(n3556), .B(n3555), .Z(n3560) );
  NANDN U4228 ( .A(n3558), .B(n3557), .Z(n3559) );
  NAND U4229 ( .A(n3560), .B(n3559), .Z(n3579) );
  XNOR U4230 ( .A(n3578), .B(n3579), .Z(n3580) );
  NANDN U4231 ( .A(n3562), .B(n3561), .Z(n3566) );
  NAND U4232 ( .A(n3564), .B(n3563), .Z(n3565) );
  NAND U4233 ( .A(n3566), .B(n3565), .Z(n3581) );
  XNOR U4234 ( .A(n3580), .B(n3581), .Z(n3572) );
  XNOR U4235 ( .A(n3573), .B(n3572), .Z(n3574) );
  XNOR U4236 ( .A(n3575), .B(n3574), .Z(n3714) );
  XNOR U4237 ( .A(sreg[262]), .B(n3714), .Z(n3716) );
  NANDN U4238 ( .A(sreg[261]), .B(n3567), .Z(n3571) );
  NAND U4239 ( .A(n3569), .B(n3568), .Z(n3570) );
  NAND U4240 ( .A(n3571), .B(n3570), .Z(n3715) );
  XNOR U4241 ( .A(n3716), .B(n3715), .Z(c[262]) );
  NANDN U4242 ( .A(n3573), .B(n3572), .Z(n3577) );
  NANDN U4243 ( .A(n3575), .B(n3574), .Z(n3576) );
  AND U4244 ( .A(n3577), .B(n3576), .Z(n3722) );
  NANDN U4245 ( .A(n3579), .B(n3578), .Z(n3583) );
  NANDN U4246 ( .A(n3581), .B(n3580), .Z(n3582) );
  AND U4247 ( .A(n3583), .B(n3582), .Z(n3720) );
  NANDN U4248 ( .A(n3585), .B(n3584), .Z(n3589) );
  NANDN U4249 ( .A(n3587), .B(n3586), .Z(n3588) );
  AND U4250 ( .A(n3589), .B(n3588), .Z(n3728) );
  NANDN U4251 ( .A(n3591), .B(n3590), .Z(n3595) );
  NANDN U4252 ( .A(n3593), .B(n3592), .Z(n3594) );
  AND U4253 ( .A(n3595), .B(n3594), .Z(n3799) );
  NAND U4254 ( .A(n38385), .B(n3596), .Z(n3598) );
  XOR U4255 ( .A(b[27]), .B(a[13]), .Z(n3743) );
  NAND U4256 ( .A(n38343), .B(n3743), .Z(n3597) );
  AND U4257 ( .A(n3598), .B(n3597), .Z(n3806) );
  NAND U4258 ( .A(n183), .B(n3599), .Z(n3601) );
  XOR U4259 ( .A(b[5]), .B(a[35]), .Z(n3746) );
  NAND U4260 ( .A(n36296), .B(n3746), .Z(n3600) );
  AND U4261 ( .A(n3601), .B(n3600), .Z(n3804) );
  NAND U4262 ( .A(n190), .B(n3602), .Z(n3604) );
  XOR U4263 ( .A(b[19]), .B(a[21]), .Z(n3749) );
  NAND U4264 ( .A(n37821), .B(n3749), .Z(n3603) );
  NAND U4265 ( .A(n3604), .B(n3603), .Z(n3803) );
  XNOR U4266 ( .A(n3804), .B(n3803), .Z(n3805) );
  XNOR U4267 ( .A(n3806), .B(n3805), .Z(n3797) );
  NAND U4268 ( .A(n38470), .B(n3605), .Z(n3607) );
  XOR U4269 ( .A(b[31]), .B(a[9]), .Z(n3752) );
  NAND U4270 ( .A(n38453), .B(n3752), .Z(n3606) );
  AND U4271 ( .A(n3607), .B(n3606), .Z(n3764) );
  NAND U4272 ( .A(n181), .B(n3608), .Z(n3610) );
  XOR U4273 ( .A(b[3]), .B(a[37]), .Z(n3755) );
  NAND U4274 ( .A(n182), .B(n3755), .Z(n3609) );
  AND U4275 ( .A(n3610), .B(n3609), .Z(n3762) );
  NAND U4276 ( .A(n189), .B(n3611), .Z(n3613) );
  XOR U4277 ( .A(b[17]), .B(a[23]), .Z(n3758) );
  NAND U4278 ( .A(n37652), .B(n3758), .Z(n3612) );
  NAND U4279 ( .A(n3613), .B(n3612), .Z(n3761) );
  XNOR U4280 ( .A(n3762), .B(n3761), .Z(n3763) );
  XOR U4281 ( .A(n3764), .B(n3763), .Z(n3798) );
  XOR U4282 ( .A(n3797), .B(n3798), .Z(n3800) );
  XOR U4283 ( .A(n3799), .B(n3800), .Z(n3846) );
  NANDN U4284 ( .A(n3615), .B(n3614), .Z(n3619) );
  NANDN U4285 ( .A(n3617), .B(n3616), .Z(n3618) );
  AND U4286 ( .A(n3619), .B(n3618), .Z(n3785) );
  NANDN U4287 ( .A(n3621), .B(n3620), .Z(n3625) );
  NANDN U4288 ( .A(n3623), .B(n3622), .Z(n3624) );
  NAND U4289 ( .A(n3625), .B(n3624), .Z(n3786) );
  XNOR U4290 ( .A(n3785), .B(n3786), .Z(n3787) );
  NANDN U4291 ( .A(n3627), .B(n3626), .Z(n3631) );
  NAND U4292 ( .A(n3629), .B(n3628), .Z(n3630) );
  NAND U4293 ( .A(n3631), .B(n3630), .Z(n3788) );
  XNOR U4294 ( .A(n3787), .B(n3788), .Z(n3845) );
  XNOR U4295 ( .A(n3846), .B(n3845), .Z(n3848) );
  NAND U4296 ( .A(n3633), .B(n3632), .Z(n3637) );
  NAND U4297 ( .A(n3635), .B(n3634), .Z(n3636) );
  AND U4298 ( .A(n3637), .B(n3636), .Z(n3847) );
  XOR U4299 ( .A(n3848), .B(n3847), .Z(n3859) );
  NANDN U4300 ( .A(n3639), .B(n3638), .Z(n3643) );
  NANDN U4301 ( .A(n3641), .B(n3640), .Z(n3642) );
  AND U4302 ( .A(n3643), .B(n3642), .Z(n3857) );
  NANDN U4303 ( .A(n3649), .B(n3648), .Z(n3653) );
  OR U4304 ( .A(n3651), .B(n3650), .Z(n3652) );
  AND U4305 ( .A(n3653), .B(n3652), .Z(n3852) );
  NANDN U4306 ( .A(n3655), .B(n3654), .Z(n3659) );
  NANDN U4307 ( .A(n3657), .B(n3656), .Z(n3658) );
  AND U4308 ( .A(n3659), .B(n3658), .Z(n3792) );
  NANDN U4309 ( .A(n3661), .B(n3660), .Z(n3665) );
  OR U4310 ( .A(n3663), .B(n3662), .Z(n3664) );
  NAND U4311 ( .A(n3665), .B(n3664), .Z(n3791) );
  XNOR U4312 ( .A(n3792), .B(n3791), .Z(n3793) );
  NAND U4313 ( .A(b[0]), .B(a[39]), .Z(n3666) );
  XNOR U4314 ( .A(b[1]), .B(n3666), .Z(n3668) );
  NANDN U4315 ( .A(b[0]), .B(a[38]), .Z(n3667) );
  NAND U4316 ( .A(n3668), .B(n3667), .Z(n3740) );
  NAND U4317 ( .A(n194), .B(n3669), .Z(n3671) );
  XOR U4318 ( .A(b[29]), .B(a[11]), .Z(n3815) );
  NAND U4319 ( .A(n38456), .B(n3815), .Z(n3670) );
  AND U4320 ( .A(n3671), .B(n3670), .Z(n3738) );
  AND U4321 ( .A(b[31]), .B(a[7]), .Z(n3737) );
  XNOR U4322 ( .A(n3738), .B(n3737), .Z(n3739) );
  XNOR U4323 ( .A(n3740), .B(n3739), .Z(n3779) );
  NAND U4324 ( .A(n38185), .B(n3672), .Z(n3674) );
  XOR U4325 ( .A(b[23]), .B(a[17]), .Z(n3821) );
  NAND U4326 ( .A(n38132), .B(n3821), .Z(n3673) );
  AND U4327 ( .A(n3674), .B(n3673), .Z(n3812) );
  NAND U4328 ( .A(n184), .B(n3675), .Z(n3677) );
  XOR U4329 ( .A(b[7]), .B(a[33]), .Z(n3824) );
  NAND U4330 ( .A(n36592), .B(n3824), .Z(n3676) );
  AND U4331 ( .A(n3677), .B(n3676), .Z(n3810) );
  NAND U4332 ( .A(n38289), .B(n3678), .Z(n3680) );
  XOR U4333 ( .A(b[25]), .B(a[15]), .Z(n3827) );
  NAND U4334 ( .A(n38247), .B(n3827), .Z(n3679) );
  NAND U4335 ( .A(n3680), .B(n3679), .Z(n3809) );
  XNOR U4336 ( .A(n3810), .B(n3809), .Z(n3811) );
  XOR U4337 ( .A(n3812), .B(n3811), .Z(n3780) );
  XNOR U4338 ( .A(n3779), .B(n3780), .Z(n3781) );
  NAND U4339 ( .A(n187), .B(n3681), .Z(n3683) );
  XOR U4340 ( .A(b[13]), .B(a[27]), .Z(n3830) );
  NAND U4341 ( .A(n37295), .B(n3830), .Z(n3682) );
  AND U4342 ( .A(n3683), .B(n3682), .Z(n3774) );
  NAND U4343 ( .A(n186), .B(n3684), .Z(n3686) );
  XOR U4344 ( .A(b[11]), .B(a[29]), .Z(n3833) );
  NAND U4345 ( .A(n37097), .B(n3833), .Z(n3685) );
  NAND U4346 ( .A(n3686), .B(n3685), .Z(n3773) );
  XNOR U4347 ( .A(n3774), .B(n3773), .Z(n3775) );
  NAND U4348 ( .A(n188), .B(n3687), .Z(n3689) );
  XOR U4349 ( .A(b[15]), .B(a[25]), .Z(n3836) );
  NAND U4350 ( .A(n37382), .B(n3836), .Z(n3688) );
  AND U4351 ( .A(n3689), .B(n3688), .Z(n3770) );
  NAND U4352 ( .A(n38064), .B(n3690), .Z(n3692) );
  XOR U4353 ( .A(b[21]), .B(a[19]), .Z(n3839) );
  NAND U4354 ( .A(n37993), .B(n3839), .Z(n3691) );
  AND U4355 ( .A(n3692), .B(n3691), .Z(n3768) );
  NAND U4356 ( .A(n185), .B(n3693), .Z(n3695) );
  XOR U4357 ( .A(b[9]), .B(a[31]), .Z(n3842) );
  NAND U4358 ( .A(n36805), .B(n3842), .Z(n3694) );
  NAND U4359 ( .A(n3695), .B(n3694), .Z(n3767) );
  XNOR U4360 ( .A(n3768), .B(n3767), .Z(n3769) );
  XOR U4361 ( .A(n3770), .B(n3769), .Z(n3776) );
  XOR U4362 ( .A(n3775), .B(n3776), .Z(n3782) );
  XOR U4363 ( .A(n3781), .B(n3782), .Z(n3794) );
  XNOR U4364 ( .A(n3793), .B(n3794), .Z(n3851) );
  XNOR U4365 ( .A(n3852), .B(n3851), .Z(n3853) );
  XOR U4366 ( .A(n3854), .B(n3853), .Z(n3858) );
  XOR U4367 ( .A(n3857), .B(n3858), .Z(n3860) );
  XOR U4368 ( .A(n3859), .B(n3860), .Z(n3734) );
  NANDN U4369 ( .A(n3697), .B(n3696), .Z(n3701) );
  NAND U4370 ( .A(n3699), .B(n3698), .Z(n3700) );
  AND U4371 ( .A(n3701), .B(n3700), .Z(n3732) );
  NANDN U4372 ( .A(n3703), .B(n3702), .Z(n3707) );
  NANDN U4373 ( .A(n3705), .B(n3704), .Z(n3706) );
  AND U4374 ( .A(n3707), .B(n3706), .Z(n3731) );
  XNOR U4375 ( .A(n3732), .B(n3731), .Z(n3733) );
  XNOR U4376 ( .A(n3734), .B(n3733), .Z(n3725) );
  NANDN U4377 ( .A(n3709), .B(n3708), .Z(n3713) );
  OR U4378 ( .A(n3711), .B(n3710), .Z(n3712) );
  NAND U4379 ( .A(n3713), .B(n3712), .Z(n3726) );
  XNOR U4380 ( .A(n3725), .B(n3726), .Z(n3727) );
  XNOR U4381 ( .A(n3728), .B(n3727), .Z(n3719) );
  XNOR U4382 ( .A(n3720), .B(n3719), .Z(n3721) );
  XNOR U4383 ( .A(n3722), .B(n3721), .Z(n3863) );
  XNOR U4384 ( .A(sreg[263]), .B(n3863), .Z(n3865) );
  NANDN U4385 ( .A(sreg[262]), .B(n3714), .Z(n3718) );
  NAND U4386 ( .A(n3716), .B(n3715), .Z(n3717) );
  NAND U4387 ( .A(n3718), .B(n3717), .Z(n3864) );
  XNOR U4388 ( .A(n3865), .B(n3864), .Z(c[263]) );
  NANDN U4389 ( .A(n3720), .B(n3719), .Z(n3724) );
  NANDN U4390 ( .A(n3722), .B(n3721), .Z(n3723) );
  AND U4391 ( .A(n3724), .B(n3723), .Z(n3871) );
  NANDN U4392 ( .A(n3726), .B(n3725), .Z(n3730) );
  NANDN U4393 ( .A(n3728), .B(n3727), .Z(n3729) );
  AND U4394 ( .A(n3730), .B(n3729), .Z(n3869) );
  NANDN U4395 ( .A(n3732), .B(n3731), .Z(n3736) );
  NANDN U4396 ( .A(n3734), .B(n3733), .Z(n3735) );
  AND U4397 ( .A(n3736), .B(n3735), .Z(n3877) );
  NANDN U4398 ( .A(n3738), .B(n3737), .Z(n3742) );
  NANDN U4399 ( .A(n3740), .B(n3739), .Z(n3741) );
  AND U4400 ( .A(n3742), .B(n3741), .Z(n3960) );
  NAND U4401 ( .A(n38385), .B(n3743), .Z(n3745) );
  XOR U4402 ( .A(b[27]), .B(a[14]), .Z(n3904) );
  NAND U4403 ( .A(n38343), .B(n3904), .Z(n3744) );
  AND U4404 ( .A(n3745), .B(n3744), .Z(n3967) );
  NAND U4405 ( .A(n183), .B(n3746), .Z(n3748) );
  XOR U4406 ( .A(b[5]), .B(a[36]), .Z(n3907) );
  NAND U4407 ( .A(n36296), .B(n3907), .Z(n3747) );
  AND U4408 ( .A(n3748), .B(n3747), .Z(n3965) );
  NAND U4409 ( .A(n190), .B(n3749), .Z(n3751) );
  XOR U4410 ( .A(b[19]), .B(a[22]), .Z(n3910) );
  NAND U4411 ( .A(n37821), .B(n3910), .Z(n3750) );
  NAND U4412 ( .A(n3751), .B(n3750), .Z(n3964) );
  XNOR U4413 ( .A(n3965), .B(n3964), .Z(n3966) );
  XNOR U4414 ( .A(n3967), .B(n3966), .Z(n3958) );
  NAND U4415 ( .A(n38470), .B(n3752), .Z(n3754) );
  XOR U4416 ( .A(b[31]), .B(a[10]), .Z(n3913) );
  NAND U4417 ( .A(n38453), .B(n3913), .Z(n3753) );
  AND U4418 ( .A(n3754), .B(n3753), .Z(n3925) );
  NAND U4419 ( .A(n181), .B(n3755), .Z(n3757) );
  XOR U4420 ( .A(b[3]), .B(a[38]), .Z(n3916) );
  NAND U4421 ( .A(n182), .B(n3916), .Z(n3756) );
  AND U4422 ( .A(n3757), .B(n3756), .Z(n3923) );
  NAND U4423 ( .A(n189), .B(n3758), .Z(n3760) );
  XOR U4424 ( .A(b[17]), .B(a[24]), .Z(n3919) );
  NAND U4425 ( .A(n37652), .B(n3919), .Z(n3759) );
  NAND U4426 ( .A(n3760), .B(n3759), .Z(n3922) );
  XNOR U4427 ( .A(n3923), .B(n3922), .Z(n3924) );
  XOR U4428 ( .A(n3925), .B(n3924), .Z(n3959) );
  XOR U4429 ( .A(n3958), .B(n3959), .Z(n3961) );
  XOR U4430 ( .A(n3960), .B(n3961), .Z(n3893) );
  NANDN U4431 ( .A(n3762), .B(n3761), .Z(n3766) );
  NANDN U4432 ( .A(n3764), .B(n3763), .Z(n3765) );
  AND U4433 ( .A(n3766), .B(n3765), .Z(n3946) );
  NANDN U4434 ( .A(n3768), .B(n3767), .Z(n3772) );
  NANDN U4435 ( .A(n3770), .B(n3769), .Z(n3771) );
  NAND U4436 ( .A(n3772), .B(n3771), .Z(n3947) );
  XNOR U4437 ( .A(n3946), .B(n3947), .Z(n3948) );
  NANDN U4438 ( .A(n3774), .B(n3773), .Z(n3778) );
  NANDN U4439 ( .A(n3776), .B(n3775), .Z(n3777) );
  NAND U4440 ( .A(n3778), .B(n3777), .Z(n3949) );
  XNOR U4441 ( .A(n3948), .B(n3949), .Z(n3892) );
  XNOR U4442 ( .A(n3893), .B(n3892), .Z(n3895) );
  NANDN U4443 ( .A(n3780), .B(n3779), .Z(n3784) );
  NANDN U4444 ( .A(n3782), .B(n3781), .Z(n3783) );
  AND U4445 ( .A(n3784), .B(n3783), .Z(n3894) );
  XOR U4446 ( .A(n3895), .B(n3894), .Z(n4008) );
  NANDN U4447 ( .A(n3786), .B(n3785), .Z(n3790) );
  NANDN U4448 ( .A(n3788), .B(n3787), .Z(n3789) );
  AND U4449 ( .A(n3790), .B(n3789), .Z(n4006) );
  NANDN U4450 ( .A(n3792), .B(n3791), .Z(n3796) );
  NANDN U4451 ( .A(n3794), .B(n3793), .Z(n3795) );
  AND U4452 ( .A(n3796), .B(n3795), .Z(n3889) );
  NANDN U4453 ( .A(n3798), .B(n3797), .Z(n3802) );
  OR U4454 ( .A(n3800), .B(n3799), .Z(n3801) );
  AND U4455 ( .A(n3802), .B(n3801), .Z(n3887) );
  NANDN U4456 ( .A(n3804), .B(n3803), .Z(n3808) );
  NANDN U4457 ( .A(n3806), .B(n3805), .Z(n3807) );
  AND U4458 ( .A(n3808), .B(n3807), .Z(n3953) );
  NANDN U4459 ( .A(n3810), .B(n3809), .Z(n3814) );
  NANDN U4460 ( .A(n3812), .B(n3811), .Z(n3813) );
  NAND U4461 ( .A(n3814), .B(n3813), .Z(n3952) );
  XNOR U4462 ( .A(n3953), .B(n3952), .Z(n3954) );
  NAND U4463 ( .A(n194), .B(n3815), .Z(n3817) );
  XOR U4464 ( .A(b[29]), .B(a[12]), .Z(n3979) );
  NAND U4465 ( .A(n38456), .B(n3979), .Z(n3816) );
  AND U4466 ( .A(n3817), .B(n3816), .Z(n3899) );
  AND U4467 ( .A(b[31]), .B(a[8]), .Z(n3898) );
  XNOR U4468 ( .A(n3899), .B(n3898), .Z(n3900) );
  NAND U4469 ( .A(b[0]), .B(a[40]), .Z(n3818) );
  XNOR U4470 ( .A(b[1]), .B(n3818), .Z(n3820) );
  NANDN U4471 ( .A(b[0]), .B(a[39]), .Z(n3819) );
  NAND U4472 ( .A(n3820), .B(n3819), .Z(n3901) );
  XNOR U4473 ( .A(n3900), .B(n3901), .Z(n3940) );
  NAND U4474 ( .A(n38185), .B(n3821), .Z(n3823) );
  XOR U4475 ( .A(b[23]), .B(a[18]), .Z(n3982) );
  NAND U4476 ( .A(n38132), .B(n3982), .Z(n3822) );
  AND U4477 ( .A(n3823), .B(n3822), .Z(n3973) );
  NAND U4478 ( .A(n184), .B(n3824), .Z(n3826) );
  XOR U4479 ( .A(b[7]), .B(a[34]), .Z(n3985) );
  NAND U4480 ( .A(n36592), .B(n3985), .Z(n3825) );
  AND U4481 ( .A(n3826), .B(n3825), .Z(n3971) );
  NAND U4482 ( .A(n38289), .B(n3827), .Z(n3829) );
  XOR U4483 ( .A(b[25]), .B(a[16]), .Z(n3988) );
  NAND U4484 ( .A(n38247), .B(n3988), .Z(n3828) );
  NAND U4485 ( .A(n3829), .B(n3828), .Z(n3970) );
  XNOR U4486 ( .A(n3971), .B(n3970), .Z(n3972) );
  XOR U4487 ( .A(n3973), .B(n3972), .Z(n3941) );
  XNOR U4488 ( .A(n3940), .B(n3941), .Z(n3942) );
  NAND U4489 ( .A(n187), .B(n3830), .Z(n3832) );
  XOR U4490 ( .A(b[13]), .B(a[28]), .Z(n3991) );
  NAND U4491 ( .A(n37295), .B(n3991), .Z(n3831) );
  AND U4492 ( .A(n3832), .B(n3831), .Z(n3935) );
  NAND U4493 ( .A(n186), .B(n3833), .Z(n3835) );
  XOR U4494 ( .A(b[11]), .B(a[30]), .Z(n3994) );
  NAND U4495 ( .A(n37097), .B(n3994), .Z(n3834) );
  NAND U4496 ( .A(n3835), .B(n3834), .Z(n3934) );
  XNOR U4497 ( .A(n3935), .B(n3934), .Z(n3936) );
  NAND U4498 ( .A(n188), .B(n3836), .Z(n3838) );
  XOR U4499 ( .A(b[15]), .B(a[26]), .Z(n3997) );
  NAND U4500 ( .A(n37382), .B(n3997), .Z(n3837) );
  AND U4501 ( .A(n3838), .B(n3837), .Z(n3931) );
  NAND U4502 ( .A(n38064), .B(n3839), .Z(n3841) );
  XOR U4503 ( .A(b[21]), .B(a[20]), .Z(n4000) );
  NAND U4504 ( .A(n37993), .B(n4000), .Z(n3840) );
  AND U4505 ( .A(n3841), .B(n3840), .Z(n3929) );
  NAND U4506 ( .A(n185), .B(n3842), .Z(n3844) );
  XOR U4507 ( .A(b[9]), .B(a[32]), .Z(n4003) );
  NAND U4508 ( .A(n36805), .B(n4003), .Z(n3843) );
  NAND U4509 ( .A(n3844), .B(n3843), .Z(n3928) );
  XNOR U4510 ( .A(n3929), .B(n3928), .Z(n3930) );
  XOR U4511 ( .A(n3931), .B(n3930), .Z(n3937) );
  XOR U4512 ( .A(n3936), .B(n3937), .Z(n3943) );
  XOR U4513 ( .A(n3942), .B(n3943), .Z(n3955) );
  XNOR U4514 ( .A(n3954), .B(n3955), .Z(n3886) );
  XNOR U4515 ( .A(n3887), .B(n3886), .Z(n3888) );
  XOR U4516 ( .A(n3889), .B(n3888), .Z(n4007) );
  XOR U4517 ( .A(n4006), .B(n4007), .Z(n4009) );
  XOR U4518 ( .A(n4008), .B(n4009), .Z(n3883) );
  NANDN U4519 ( .A(n3846), .B(n3845), .Z(n3850) );
  NAND U4520 ( .A(n3848), .B(n3847), .Z(n3849) );
  AND U4521 ( .A(n3850), .B(n3849), .Z(n3881) );
  NANDN U4522 ( .A(n3852), .B(n3851), .Z(n3856) );
  NANDN U4523 ( .A(n3854), .B(n3853), .Z(n3855) );
  AND U4524 ( .A(n3856), .B(n3855), .Z(n3880) );
  XNOR U4525 ( .A(n3881), .B(n3880), .Z(n3882) );
  XNOR U4526 ( .A(n3883), .B(n3882), .Z(n3874) );
  NANDN U4527 ( .A(n3858), .B(n3857), .Z(n3862) );
  OR U4528 ( .A(n3860), .B(n3859), .Z(n3861) );
  NAND U4529 ( .A(n3862), .B(n3861), .Z(n3875) );
  XNOR U4530 ( .A(n3874), .B(n3875), .Z(n3876) );
  XNOR U4531 ( .A(n3877), .B(n3876), .Z(n3868) );
  XNOR U4532 ( .A(n3869), .B(n3868), .Z(n3870) );
  XNOR U4533 ( .A(n3871), .B(n3870), .Z(n4012) );
  XNOR U4534 ( .A(sreg[264]), .B(n4012), .Z(n4014) );
  NANDN U4535 ( .A(sreg[263]), .B(n3863), .Z(n3867) );
  NAND U4536 ( .A(n3865), .B(n3864), .Z(n3866) );
  NAND U4537 ( .A(n3867), .B(n3866), .Z(n4013) );
  XNOR U4538 ( .A(n4014), .B(n4013), .Z(c[264]) );
  NANDN U4539 ( .A(n3869), .B(n3868), .Z(n3873) );
  NANDN U4540 ( .A(n3871), .B(n3870), .Z(n3872) );
  AND U4541 ( .A(n3873), .B(n3872), .Z(n4020) );
  NANDN U4542 ( .A(n3875), .B(n3874), .Z(n3879) );
  NANDN U4543 ( .A(n3877), .B(n3876), .Z(n3878) );
  AND U4544 ( .A(n3879), .B(n3878), .Z(n4018) );
  NANDN U4545 ( .A(n3881), .B(n3880), .Z(n3885) );
  NANDN U4546 ( .A(n3883), .B(n3882), .Z(n3884) );
  AND U4547 ( .A(n3885), .B(n3884), .Z(n4026) );
  NANDN U4548 ( .A(n3887), .B(n3886), .Z(n3891) );
  NANDN U4549 ( .A(n3889), .B(n3888), .Z(n3890) );
  AND U4550 ( .A(n3891), .B(n3890), .Z(n4030) );
  NANDN U4551 ( .A(n3893), .B(n3892), .Z(n3897) );
  NAND U4552 ( .A(n3895), .B(n3894), .Z(n3896) );
  AND U4553 ( .A(n3897), .B(n3896), .Z(n4029) );
  XNOR U4554 ( .A(n4030), .B(n4029), .Z(n4032) );
  NANDN U4555 ( .A(n3899), .B(n3898), .Z(n3903) );
  NANDN U4556 ( .A(n3901), .B(n3900), .Z(n3902) );
  AND U4557 ( .A(n3903), .B(n3902), .Z(n4107) );
  NAND U4558 ( .A(n38385), .B(n3904), .Z(n3906) );
  XOR U4559 ( .A(b[27]), .B(a[15]), .Z(n4053) );
  NAND U4560 ( .A(n38343), .B(n4053), .Z(n3905) );
  AND U4561 ( .A(n3906), .B(n3905), .Z(n4114) );
  NAND U4562 ( .A(n183), .B(n3907), .Z(n3909) );
  XOR U4563 ( .A(b[5]), .B(a[37]), .Z(n4056) );
  NAND U4564 ( .A(n36296), .B(n4056), .Z(n3908) );
  AND U4565 ( .A(n3909), .B(n3908), .Z(n4112) );
  NAND U4566 ( .A(n190), .B(n3910), .Z(n3912) );
  XOR U4567 ( .A(b[19]), .B(a[23]), .Z(n4059) );
  NAND U4568 ( .A(n37821), .B(n4059), .Z(n3911) );
  NAND U4569 ( .A(n3912), .B(n3911), .Z(n4111) );
  XNOR U4570 ( .A(n4112), .B(n4111), .Z(n4113) );
  XNOR U4571 ( .A(n4114), .B(n4113), .Z(n4105) );
  NAND U4572 ( .A(n38470), .B(n3913), .Z(n3915) );
  XOR U4573 ( .A(b[31]), .B(a[11]), .Z(n4062) );
  NAND U4574 ( .A(n38453), .B(n4062), .Z(n3914) );
  AND U4575 ( .A(n3915), .B(n3914), .Z(n4074) );
  NAND U4576 ( .A(n181), .B(n3916), .Z(n3918) );
  XOR U4577 ( .A(b[3]), .B(a[39]), .Z(n4065) );
  NAND U4578 ( .A(n182), .B(n4065), .Z(n3917) );
  AND U4579 ( .A(n3918), .B(n3917), .Z(n4072) );
  NAND U4580 ( .A(n189), .B(n3919), .Z(n3921) );
  XOR U4581 ( .A(b[17]), .B(a[25]), .Z(n4068) );
  NAND U4582 ( .A(n37652), .B(n4068), .Z(n3920) );
  NAND U4583 ( .A(n3921), .B(n3920), .Z(n4071) );
  XNOR U4584 ( .A(n4072), .B(n4071), .Z(n4073) );
  XOR U4585 ( .A(n4074), .B(n4073), .Z(n4106) );
  XOR U4586 ( .A(n4105), .B(n4106), .Z(n4108) );
  XOR U4587 ( .A(n4107), .B(n4108), .Z(n4042) );
  NANDN U4588 ( .A(n3923), .B(n3922), .Z(n3927) );
  NANDN U4589 ( .A(n3925), .B(n3924), .Z(n3926) );
  AND U4590 ( .A(n3927), .B(n3926), .Z(n4095) );
  NANDN U4591 ( .A(n3929), .B(n3928), .Z(n3933) );
  NANDN U4592 ( .A(n3931), .B(n3930), .Z(n3932) );
  NAND U4593 ( .A(n3933), .B(n3932), .Z(n4096) );
  XNOR U4594 ( .A(n4095), .B(n4096), .Z(n4097) );
  NANDN U4595 ( .A(n3935), .B(n3934), .Z(n3939) );
  NANDN U4596 ( .A(n3937), .B(n3936), .Z(n3938) );
  NAND U4597 ( .A(n3939), .B(n3938), .Z(n4098) );
  XNOR U4598 ( .A(n4097), .B(n4098), .Z(n4041) );
  XNOR U4599 ( .A(n4042), .B(n4041), .Z(n4044) );
  NANDN U4600 ( .A(n3941), .B(n3940), .Z(n3945) );
  NANDN U4601 ( .A(n3943), .B(n3942), .Z(n3944) );
  AND U4602 ( .A(n3945), .B(n3944), .Z(n4043) );
  XOR U4603 ( .A(n4044), .B(n4043), .Z(n4156) );
  NANDN U4604 ( .A(n3947), .B(n3946), .Z(n3951) );
  NANDN U4605 ( .A(n3949), .B(n3948), .Z(n3950) );
  AND U4606 ( .A(n3951), .B(n3950), .Z(n4153) );
  NANDN U4607 ( .A(n3953), .B(n3952), .Z(n3957) );
  NANDN U4608 ( .A(n3955), .B(n3954), .Z(n3956) );
  AND U4609 ( .A(n3957), .B(n3956), .Z(n4038) );
  NANDN U4610 ( .A(n3959), .B(n3958), .Z(n3963) );
  OR U4611 ( .A(n3961), .B(n3960), .Z(n3962) );
  AND U4612 ( .A(n3963), .B(n3962), .Z(n4036) );
  NANDN U4613 ( .A(n3965), .B(n3964), .Z(n3969) );
  NANDN U4614 ( .A(n3967), .B(n3966), .Z(n3968) );
  AND U4615 ( .A(n3969), .B(n3968), .Z(n4102) );
  NANDN U4616 ( .A(n3971), .B(n3970), .Z(n3975) );
  NANDN U4617 ( .A(n3973), .B(n3972), .Z(n3974) );
  NAND U4618 ( .A(n3975), .B(n3974), .Z(n4101) );
  XNOR U4619 ( .A(n4102), .B(n4101), .Z(n4104) );
  NAND U4620 ( .A(b[0]), .B(a[41]), .Z(n3976) );
  XNOR U4621 ( .A(b[1]), .B(n3976), .Z(n3978) );
  NANDN U4622 ( .A(b[0]), .B(a[40]), .Z(n3977) );
  NAND U4623 ( .A(n3978), .B(n3977), .Z(n4050) );
  NAND U4624 ( .A(n194), .B(n3979), .Z(n3981) );
  XOR U4625 ( .A(b[29]), .B(a[13]), .Z(n4126) );
  NAND U4626 ( .A(n38456), .B(n4126), .Z(n3980) );
  AND U4627 ( .A(n3981), .B(n3980), .Z(n4048) );
  AND U4628 ( .A(b[31]), .B(a[9]), .Z(n4047) );
  XNOR U4629 ( .A(n4048), .B(n4047), .Z(n4049) );
  XNOR U4630 ( .A(n4050), .B(n4049), .Z(n4090) );
  NAND U4631 ( .A(n38185), .B(n3982), .Z(n3984) );
  XOR U4632 ( .A(b[23]), .B(a[19]), .Z(n4129) );
  NAND U4633 ( .A(n38132), .B(n4129), .Z(n3983) );
  AND U4634 ( .A(n3984), .B(n3983), .Z(n4119) );
  NAND U4635 ( .A(n184), .B(n3985), .Z(n3987) );
  XOR U4636 ( .A(b[7]), .B(a[35]), .Z(n4132) );
  NAND U4637 ( .A(n36592), .B(n4132), .Z(n3986) );
  AND U4638 ( .A(n3987), .B(n3986), .Z(n4118) );
  NAND U4639 ( .A(n38289), .B(n3988), .Z(n3990) );
  XOR U4640 ( .A(b[25]), .B(a[17]), .Z(n4135) );
  NAND U4641 ( .A(n38247), .B(n4135), .Z(n3989) );
  NAND U4642 ( .A(n3990), .B(n3989), .Z(n4117) );
  XOR U4643 ( .A(n4118), .B(n4117), .Z(n4120) );
  XOR U4644 ( .A(n4119), .B(n4120), .Z(n4089) );
  XOR U4645 ( .A(n4090), .B(n4089), .Z(n4092) );
  NAND U4646 ( .A(n187), .B(n3991), .Z(n3993) );
  XOR U4647 ( .A(b[13]), .B(a[29]), .Z(n4138) );
  NAND U4648 ( .A(n37295), .B(n4138), .Z(n3992) );
  AND U4649 ( .A(n3993), .B(n3992), .Z(n4084) );
  NAND U4650 ( .A(n186), .B(n3994), .Z(n3996) );
  XOR U4651 ( .A(b[11]), .B(a[31]), .Z(n4141) );
  NAND U4652 ( .A(n37097), .B(n4141), .Z(n3995) );
  NAND U4653 ( .A(n3996), .B(n3995), .Z(n4083) );
  XNOR U4654 ( .A(n4084), .B(n4083), .Z(n4086) );
  NAND U4655 ( .A(n188), .B(n3997), .Z(n3999) );
  XOR U4656 ( .A(b[15]), .B(a[27]), .Z(n4144) );
  NAND U4657 ( .A(n37382), .B(n4144), .Z(n3998) );
  AND U4658 ( .A(n3999), .B(n3998), .Z(n4080) );
  NAND U4659 ( .A(n38064), .B(n4000), .Z(n4002) );
  XOR U4660 ( .A(b[21]), .B(a[21]), .Z(n4147) );
  NAND U4661 ( .A(n37993), .B(n4147), .Z(n4001) );
  AND U4662 ( .A(n4002), .B(n4001), .Z(n4078) );
  NAND U4663 ( .A(n185), .B(n4003), .Z(n4005) );
  XOR U4664 ( .A(b[9]), .B(a[33]), .Z(n4150) );
  NAND U4665 ( .A(n36805), .B(n4150), .Z(n4004) );
  NAND U4666 ( .A(n4005), .B(n4004), .Z(n4077) );
  XNOR U4667 ( .A(n4078), .B(n4077), .Z(n4079) );
  XNOR U4668 ( .A(n4080), .B(n4079), .Z(n4085) );
  XOR U4669 ( .A(n4086), .B(n4085), .Z(n4091) );
  XNOR U4670 ( .A(n4092), .B(n4091), .Z(n4103) );
  XNOR U4671 ( .A(n4104), .B(n4103), .Z(n4035) );
  XNOR U4672 ( .A(n4036), .B(n4035), .Z(n4037) );
  XOR U4673 ( .A(n4038), .B(n4037), .Z(n4154) );
  XNOR U4674 ( .A(n4153), .B(n4154), .Z(n4155) );
  XNOR U4675 ( .A(n4156), .B(n4155), .Z(n4031) );
  XOR U4676 ( .A(n4032), .B(n4031), .Z(n4024) );
  NANDN U4677 ( .A(n4007), .B(n4006), .Z(n4011) );
  OR U4678 ( .A(n4009), .B(n4008), .Z(n4010) );
  AND U4679 ( .A(n4011), .B(n4010), .Z(n4023) );
  XNOR U4680 ( .A(n4024), .B(n4023), .Z(n4025) );
  XNOR U4681 ( .A(n4026), .B(n4025), .Z(n4017) );
  XNOR U4682 ( .A(n4018), .B(n4017), .Z(n4019) );
  XNOR U4683 ( .A(n4020), .B(n4019), .Z(n4159) );
  XNOR U4684 ( .A(sreg[265]), .B(n4159), .Z(n4161) );
  NANDN U4685 ( .A(sreg[264]), .B(n4012), .Z(n4016) );
  NAND U4686 ( .A(n4014), .B(n4013), .Z(n4015) );
  NAND U4687 ( .A(n4016), .B(n4015), .Z(n4160) );
  XNOR U4688 ( .A(n4161), .B(n4160), .Z(c[265]) );
  NANDN U4689 ( .A(n4018), .B(n4017), .Z(n4022) );
  NANDN U4690 ( .A(n4020), .B(n4019), .Z(n4021) );
  AND U4691 ( .A(n4022), .B(n4021), .Z(n4167) );
  NANDN U4692 ( .A(n4024), .B(n4023), .Z(n4028) );
  NANDN U4693 ( .A(n4026), .B(n4025), .Z(n4027) );
  AND U4694 ( .A(n4028), .B(n4027), .Z(n4165) );
  NANDN U4695 ( .A(n4030), .B(n4029), .Z(n4034) );
  NAND U4696 ( .A(n4032), .B(n4031), .Z(n4033) );
  AND U4697 ( .A(n4034), .B(n4033), .Z(n4172) );
  NANDN U4698 ( .A(n4036), .B(n4035), .Z(n4040) );
  NANDN U4699 ( .A(n4038), .B(n4037), .Z(n4039) );
  AND U4700 ( .A(n4040), .B(n4039), .Z(n4177) );
  NANDN U4701 ( .A(n4042), .B(n4041), .Z(n4046) );
  NAND U4702 ( .A(n4044), .B(n4043), .Z(n4045) );
  AND U4703 ( .A(n4046), .B(n4045), .Z(n4176) );
  XNOR U4704 ( .A(n4177), .B(n4176), .Z(n4179) );
  NANDN U4705 ( .A(n4048), .B(n4047), .Z(n4052) );
  NANDN U4706 ( .A(n4050), .B(n4049), .Z(n4051) );
  AND U4707 ( .A(n4052), .B(n4051), .Z(n4244) );
  NAND U4708 ( .A(n38385), .B(n4053), .Z(n4055) );
  XOR U4709 ( .A(b[27]), .B(a[16]), .Z(n4188) );
  NAND U4710 ( .A(n38343), .B(n4188), .Z(n4054) );
  AND U4711 ( .A(n4055), .B(n4054), .Z(n4251) );
  NAND U4712 ( .A(n183), .B(n4056), .Z(n4058) );
  XOR U4713 ( .A(b[5]), .B(a[38]), .Z(n4191) );
  NAND U4714 ( .A(n36296), .B(n4191), .Z(n4057) );
  AND U4715 ( .A(n4058), .B(n4057), .Z(n4249) );
  NAND U4716 ( .A(n190), .B(n4059), .Z(n4061) );
  XOR U4717 ( .A(b[19]), .B(a[24]), .Z(n4194) );
  NAND U4718 ( .A(n37821), .B(n4194), .Z(n4060) );
  NAND U4719 ( .A(n4061), .B(n4060), .Z(n4248) );
  XNOR U4720 ( .A(n4249), .B(n4248), .Z(n4250) );
  XNOR U4721 ( .A(n4251), .B(n4250), .Z(n4242) );
  NAND U4722 ( .A(n38470), .B(n4062), .Z(n4064) );
  XOR U4723 ( .A(b[31]), .B(a[12]), .Z(n4197) );
  NAND U4724 ( .A(n38453), .B(n4197), .Z(n4063) );
  AND U4725 ( .A(n4064), .B(n4063), .Z(n4209) );
  NAND U4726 ( .A(n181), .B(n4065), .Z(n4067) );
  XOR U4727 ( .A(b[3]), .B(a[40]), .Z(n4200) );
  NAND U4728 ( .A(n182), .B(n4200), .Z(n4066) );
  AND U4729 ( .A(n4067), .B(n4066), .Z(n4207) );
  NAND U4730 ( .A(n189), .B(n4068), .Z(n4070) );
  XOR U4731 ( .A(b[17]), .B(a[26]), .Z(n4203) );
  NAND U4732 ( .A(n37652), .B(n4203), .Z(n4069) );
  NAND U4733 ( .A(n4070), .B(n4069), .Z(n4206) );
  XNOR U4734 ( .A(n4207), .B(n4206), .Z(n4208) );
  XOR U4735 ( .A(n4209), .B(n4208), .Z(n4243) );
  XOR U4736 ( .A(n4242), .B(n4243), .Z(n4245) );
  XOR U4737 ( .A(n4244), .B(n4245), .Z(n4291) );
  NANDN U4738 ( .A(n4072), .B(n4071), .Z(n4076) );
  NANDN U4739 ( .A(n4074), .B(n4073), .Z(n4075) );
  AND U4740 ( .A(n4076), .B(n4075), .Z(n4230) );
  NANDN U4741 ( .A(n4078), .B(n4077), .Z(n4082) );
  NANDN U4742 ( .A(n4080), .B(n4079), .Z(n4081) );
  NAND U4743 ( .A(n4082), .B(n4081), .Z(n4231) );
  XNOR U4744 ( .A(n4230), .B(n4231), .Z(n4232) );
  NANDN U4745 ( .A(n4084), .B(n4083), .Z(n4088) );
  NAND U4746 ( .A(n4086), .B(n4085), .Z(n4087) );
  NAND U4747 ( .A(n4088), .B(n4087), .Z(n4233) );
  XNOR U4748 ( .A(n4232), .B(n4233), .Z(n4290) );
  XNOR U4749 ( .A(n4291), .B(n4290), .Z(n4293) );
  NAND U4750 ( .A(n4090), .B(n4089), .Z(n4094) );
  NAND U4751 ( .A(n4092), .B(n4091), .Z(n4093) );
  AND U4752 ( .A(n4094), .B(n4093), .Z(n4292) );
  XOR U4753 ( .A(n4293), .B(n4292), .Z(n4305) );
  NANDN U4754 ( .A(n4096), .B(n4095), .Z(n4100) );
  NANDN U4755 ( .A(n4098), .B(n4097), .Z(n4099) );
  AND U4756 ( .A(n4100), .B(n4099), .Z(n4302) );
  NANDN U4757 ( .A(n4106), .B(n4105), .Z(n4110) );
  OR U4758 ( .A(n4108), .B(n4107), .Z(n4109) );
  AND U4759 ( .A(n4110), .B(n4109), .Z(n4297) );
  NANDN U4760 ( .A(n4112), .B(n4111), .Z(n4116) );
  NANDN U4761 ( .A(n4114), .B(n4113), .Z(n4115) );
  AND U4762 ( .A(n4116), .B(n4115), .Z(n4237) );
  NANDN U4763 ( .A(n4118), .B(n4117), .Z(n4122) );
  OR U4764 ( .A(n4120), .B(n4119), .Z(n4121) );
  NAND U4765 ( .A(n4122), .B(n4121), .Z(n4236) );
  XNOR U4766 ( .A(n4237), .B(n4236), .Z(n4238) );
  NAND U4767 ( .A(b[0]), .B(a[42]), .Z(n4123) );
  XNOR U4768 ( .A(b[1]), .B(n4123), .Z(n4125) );
  NANDN U4769 ( .A(b[0]), .B(a[41]), .Z(n4124) );
  NAND U4770 ( .A(n4125), .B(n4124), .Z(n4185) );
  NAND U4771 ( .A(n194), .B(n4126), .Z(n4128) );
  XOR U4772 ( .A(b[29]), .B(a[14]), .Z(n4263) );
  NAND U4773 ( .A(n38456), .B(n4263), .Z(n4127) );
  AND U4774 ( .A(n4128), .B(n4127), .Z(n4183) );
  AND U4775 ( .A(b[31]), .B(a[10]), .Z(n4182) );
  XNOR U4776 ( .A(n4183), .B(n4182), .Z(n4184) );
  XNOR U4777 ( .A(n4185), .B(n4184), .Z(n4224) );
  NAND U4778 ( .A(n38185), .B(n4129), .Z(n4131) );
  XOR U4779 ( .A(b[23]), .B(a[20]), .Z(n4266) );
  NAND U4780 ( .A(n38132), .B(n4266), .Z(n4130) );
  AND U4781 ( .A(n4131), .B(n4130), .Z(n4257) );
  NAND U4782 ( .A(n184), .B(n4132), .Z(n4134) );
  XOR U4783 ( .A(b[7]), .B(a[36]), .Z(n4269) );
  NAND U4784 ( .A(n36592), .B(n4269), .Z(n4133) );
  AND U4785 ( .A(n4134), .B(n4133), .Z(n4255) );
  NAND U4786 ( .A(n38289), .B(n4135), .Z(n4137) );
  XOR U4787 ( .A(b[25]), .B(a[18]), .Z(n4272) );
  NAND U4788 ( .A(n38247), .B(n4272), .Z(n4136) );
  NAND U4789 ( .A(n4137), .B(n4136), .Z(n4254) );
  XNOR U4790 ( .A(n4255), .B(n4254), .Z(n4256) );
  XOR U4791 ( .A(n4257), .B(n4256), .Z(n4225) );
  XNOR U4792 ( .A(n4224), .B(n4225), .Z(n4226) );
  NAND U4793 ( .A(n187), .B(n4138), .Z(n4140) );
  XOR U4794 ( .A(b[13]), .B(a[30]), .Z(n4275) );
  NAND U4795 ( .A(n37295), .B(n4275), .Z(n4139) );
  AND U4796 ( .A(n4140), .B(n4139), .Z(n4219) );
  NAND U4797 ( .A(n186), .B(n4141), .Z(n4143) );
  XOR U4798 ( .A(b[11]), .B(a[32]), .Z(n4278) );
  NAND U4799 ( .A(n37097), .B(n4278), .Z(n4142) );
  NAND U4800 ( .A(n4143), .B(n4142), .Z(n4218) );
  XNOR U4801 ( .A(n4219), .B(n4218), .Z(n4220) );
  NAND U4802 ( .A(n188), .B(n4144), .Z(n4146) );
  XOR U4803 ( .A(b[15]), .B(a[28]), .Z(n4281) );
  NAND U4804 ( .A(n37382), .B(n4281), .Z(n4145) );
  AND U4805 ( .A(n4146), .B(n4145), .Z(n4215) );
  NAND U4806 ( .A(n38064), .B(n4147), .Z(n4149) );
  XOR U4807 ( .A(b[21]), .B(a[22]), .Z(n4284) );
  NAND U4808 ( .A(n37993), .B(n4284), .Z(n4148) );
  AND U4809 ( .A(n4149), .B(n4148), .Z(n4213) );
  NAND U4810 ( .A(n185), .B(n4150), .Z(n4152) );
  XOR U4811 ( .A(b[9]), .B(a[34]), .Z(n4287) );
  NAND U4812 ( .A(n36805), .B(n4287), .Z(n4151) );
  NAND U4813 ( .A(n4152), .B(n4151), .Z(n4212) );
  XNOR U4814 ( .A(n4213), .B(n4212), .Z(n4214) );
  XOR U4815 ( .A(n4215), .B(n4214), .Z(n4221) );
  XOR U4816 ( .A(n4220), .B(n4221), .Z(n4227) );
  XOR U4817 ( .A(n4226), .B(n4227), .Z(n4239) );
  XNOR U4818 ( .A(n4238), .B(n4239), .Z(n4296) );
  XNOR U4819 ( .A(n4297), .B(n4296), .Z(n4298) );
  XOR U4820 ( .A(n4299), .B(n4298), .Z(n4303) );
  XNOR U4821 ( .A(n4302), .B(n4303), .Z(n4304) );
  XNOR U4822 ( .A(n4305), .B(n4304), .Z(n4178) );
  XOR U4823 ( .A(n4179), .B(n4178), .Z(n4171) );
  NANDN U4824 ( .A(n4154), .B(n4153), .Z(n4158) );
  NANDN U4825 ( .A(n4156), .B(n4155), .Z(n4157) );
  AND U4826 ( .A(n4158), .B(n4157), .Z(n4170) );
  XOR U4827 ( .A(n4171), .B(n4170), .Z(n4173) );
  XNOR U4828 ( .A(n4172), .B(n4173), .Z(n4164) );
  XNOR U4829 ( .A(n4165), .B(n4164), .Z(n4166) );
  XNOR U4830 ( .A(n4167), .B(n4166), .Z(n4308) );
  XNOR U4831 ( .A(sreg[266]), .B(n4308), .Z(n4310) );
  NANDN U4832 ( .A(sreg[265]), .B(n4159), .Z(n4163) );
  NAND U4833 ( .A(n4161), .B(n4160), .Z(n4162) );
  NAND U4834 ( .A(n4163), .B(n4162), .Z(n4309) );
  XNOR U4835 ( .A(n4310), .B(n4309), .Z(c[266]) );
  NANDN U4836 ( .A(n4165), .B(n4164), .Z(n4169) );
  NANDN U4837 ( .A(n4167), .B(n4166), .Z(n4168) );
  AND U4838 ( .A(n4169), .B(n4168), .Z(n4316) );
  NANDN U4839 ( .A(n4171), .B(n4170), .Z(n4175) );
  NANDN U4840 ( .A(n4173), .B(n4172), .Z(n4174) );
  AND U4841 ( .A(n4175), .B(n4174), .Z(n4314) );
  NANDN U4842 ( .A(n4177), .B(n4176), .Z(n4181) );
  NAND U4843 ( .A(n4179), .B(n4178), .Z(n4180) );
  AND U4844 ( .A(n4181), .B(n4180), .Z(n4321) );
  NANDN U4845 ( .A(n4183), .B(n4182), .Z(n4187) );
  NANDN U4846 ( .A(n4185), .B(n4184), .Z(n4186) );
  AND U4847 ( .A(n4187), .B(n4186), .Z(n4405) );
  NAND U4848 ( .A(n38385), .B(n4188), .Z(n4190) );
  XOR U4849 ( .A(b[27]), .B(a[17]), .Z(n4349) );
  NAND U4850 ( .A(n38343), .B(n4349), .Z(n4189) );
  AND U4851 ( .A(n4190), .B(n4189), .Z(n4412) );
  NAND U4852 ( .A(n183), .B(n4191), .Z(n4193) );
  XOR U4853 ( .A(b[5]), .B(a[39]), .Z(n4352) );
  NAND U4854 ( .A(n36296), .B(n4352), .Z(n4192) );
  AND U4855 ( .A(n4193), .B(n4192), .Z(n4410) );
  NAND U4856 ( .A(n190), .B(n4194), .Z(n4196) );
  XOR U4857 ( .A(b[19]), .B(a[25]), .Z(n4355) );
  NAND U4858 ( .A(n37821), .B(n4355), .Z(n4195) );
  NAND U4859 ( .A(n4196), .B(n4195), .Z(n4409) );
  XNOR U4860 ( .A(n4410), .B(n4409), .Z(n4411) );
  XNOR U4861 ( .A(n4412), .B(n4411), .Z(n4403) );
  NAND U4862 ( .A(n38470), .B(n4197), .Z(n4199) );
  XOR U4863 ( .A(b[31]), .B(a[13]), .Z(n4358) );
  NAND U4864 ( .A(n38453), .B(n4358), .Z(n4198) );
  AND U4865 ( .A(n4199), .B(n4198), .Z(n4370) );
  NAND U4866 ( .A(n181), .B(n4200), .Z(n4202) );
  XOR U4867 ( .A(b[3]), .B(a[41]), .Z(n4361) );
  NAND U4868 ( .A(n182), .B(n4361), .Z(n4201) );
  AND U4869 ( .A(n4202), .B(n4201), .Z(n4368) );
  NAND U4870 ( .A(n189), .B(n4203), .Z(n4205) );
  XOR U4871 ( .A(b[17]), .B(a[27]), .Z(n4364) );
  NAND U4872 ( .A(n37652), .B(n4364), .Z(n4204) );
  NAND U4873 ( .A(n4205), .B(n4204), .Z(n4367) );
  XNOR U4874 ( .A(n4368), .B(n4367), .Z(n4369) );
  XOR U4875 ( .A(n4370), .B(n4369), .Z(n4404) );
  XOR U4876 ( .A(n4403), .B(n4404), .Z(n4406) );
  XOR U4877 ( .A(n4405), .B(n4406), .Z(n4338) );
  NANDN U4878 ( .A(n4207), .B(n4206), .Z(n4211) );
  NANDN U4879 ( .A(n4209), .B(n4208), .Z(n4210) );
  AND U4880 ( .A(n4211), .B(n4210), .Z(n4391) );
  NANDN U4881 ( .A(n4213), .B(n4212), .Z(n4217) );
  NANDN U4882 ( .A(n4215), .B(n4214), .Z(n4216) );
  NAND U4883 ( .A(n4217), .B(n4216), .Z(n4392) );
  XNOR U4884 ( .A(n4391), .B(n4392), .Z(n4393) );
  NANDN U4885 ( .A(n4219), .B(n4218), .Z(n4223) );
  NANDN U4886 ( .A(n4221), .B(n4220), .Z(n4222) );
  NAND U4887 ( .A(n4223), .B(n4222), .Z(n4394) );
  XNOR U4888 ( .A(n4393), .B(n4394), .Z(n4337) );
  XNOR U4889 ( .A(n4338), .B(n4337), .Z(n4340) );
  NANDN U4890 ( .A(n4225), .B(n4224), .Z(n4229) );
  NANDN U4891 ( .A(n4227), .B(n4226), .Z(n4228) );
  AND U4892 ( .A(n4229), .B(n4228), .Z(n4339) );
  XOR U4893 ( .A(n4340), .B(n4339), .Z(n4453) );
  NANDN U4894 ( .A(n4231), .B(n4230), .Z(n4235) );
  NANDN U4895 ( .A(n4233), .B(n4232), .Z(n4234) );
  AND U4896 ( .A(n4235), .B(n4234), .Z(n4451) );
  NANDN U4897 ( .A(n4237), .B(n4236), .Z(n4241) );
  NANDN U4898 ( .A(n4239), .B(n4238), .Z(n4240) );
  AND U4899 ( .A(n4241), .B(n4240), .Z(n4334) );
  NANDN U4900 ( .A(n4243), .B(n4242), .Z(n4247) );
  OR U4901 ( .A(n4245), .B(n4244), .Z(n4246) );
  AND U4902 ( .A(n4247), .B(n4246), .Z(n4332) );
  NANDN U4903 ( .A(n4249), .B(n4248), .Z(n4253) );
  NANDN U4904 ( .A(n4251), .B(n4250), .Z(n4252) );
  AND U4905 ( .A(n4253), .B(n4252), .Z(n4398) );
  NANDN U4906 ( .A(n4255), .B(n4254), .Z(n4259) );
  NANDN U4907 ( .A(n4257), .B(n4256), .Z(n4258) );
  NAND U4908 ( .A(n4259), .B(n4258), .Z(n4397) );
  XNOR U4909 ( .A(n4398), .B(n4397), .Z(n4399) );
  NAND U4910 ( .A(b[0]), .B(a[43]), .Z(n4260) );
  XNOR U4911 ( .A(b[1]), .B(n4260), .Z(n4262) );
  NANDN U4912 ( .A(b[0]), .B(a[42]), .Z(n4261) );
  NAND U4913 ( .A(n4262), .B(n4261), .Z(n4346) );
  NAND U4914 ( .A(n194), .B(n4263), .Z(n4265) );
  XOR U4915 ( .A(b[29]), .B(a[15]), .Z(n4424) );
  NAND U4916 ( .A(n38456), .B(n4424), .Z(n4264) );
  AND U4917 ( .A(n4265), .B(n4264), .Z(n4344) );
  AND U4918 ( .A(b[31]), .B(a[11]), .Z(n4343) );
  XNOR U4919 ( .A(n4344), .B(n4343), .Z(n4345) );
  XNOR U4920 ( .A(n4346), .B(n4345), .Z(n4385) );
  NAND U4921 ( .A(n38185), .B(n4266), .Z(n4268) );
  XOR U4922 ( .A(b[23]), .B(a[21]), .Z(n4427) );
  NAND U4923 ( .A(n38132), .B(n4427), .Z(n4267) );
  AND U4924 ( .A(n4268), .B(n4267), .Z(n4418) );
  NAND U4925 ( .A(n184), .B(n4269), .Z(n4271) );
  XOR U4926 ( .A(b[7]), .B(a[37]), .Z(n4430) );
  NAND U4927 ( .A(n36592), .B(n4430), .Z(n4270) );
  AND U4928 ( .A(n4271), .B(n4270), .Z(n4416) );
  NAND U4929 ( .A(n38289), .B(n4272), .Z(n4274) );
  XOR U4930 ( .A(b[25]), .B(a[19]), .Z(n4433) );
  NAND U4931 ( .A(n38247), .B(n4433), .Z(n4273) );
  NAND U4932 ( .A(n4274), .B(n4273), .Z(n4415) );
  XNOR U4933 ( .A(n4416), .B(n4415), .Z(n4417) );
  XOR U4934 ( .A(n4418), .B(n4417), .Z(n4386) );
  XNOR U4935 ( .A(n4385), .B(n4386), .Z(n4387) );
  NAND U4936 ( .A(n187), .B(n4275), .Z(n4277) );
  XOR U4937 ( .A(b[13]), .B(a[31]), .Z(n4436) );
  NAND U4938 ( .A(n37295), .B(n4436), .Z(n4276) );
  AND U4939 ( .A(n4277), .B(n4276), .Z(n4380) );
  NAND U4940 ( .A(n186), .B(n4278), .Z(n4280) );
  XOR U4941 ( .A(b[11]), .B(a[33]), .Z(n4439) );
  NAND U4942 ( .A(n37097), .B(n4439), .Z(n4279) );
  NAND U4943 ( .A(n4280), .B(n4279), .Z(n4379) );
  XNOR U4944 ( .A(n4380), .B(n4379), .Z(n4381) );
  NAND U4945 ( .A(n188), .B(n4281), .Z(n4283) );
  XOR U4946 ( .A(b[15]), .B(a[29]), .Z(n4442) );
  NAND U4947 ( .A(n37382), .B(n4442), .Z(n4282) );
  AND U4948 ( .A(n4283), .B(n4282), .Z(n4376) );
  NAND U4949 ( .A(n38064), .B(n4284), .Z(n4286) );
  XOR U4950 ( .A(b[21]), .B(a[23]), .Z(n4445) );
  NAND U4951 ( .A(n37993), .B(n4445), .Z(n4285) );
  AND U4952 ( .A(n4286), .B(n4285), .Z(n4374) );
  NAND U4953 ( .A(n185), .B(n4287), .Z(n4289) );
  XOR U4954 ( .A(b[9]), .B(a[35]), .Z(n4448) );
  NAND U4955 ( .A(n36805), .B(n4448), .Z(n4288) );
  NAND U4956 ( .A(n4289), .B(n4288), .Z(n4373) );
  XNOR U4957 ( .A(n4374), .B(n4373), .Z(n4375) );
  XOR U4958 ( .A(n4376), .B(n4375), .Z(n4382) );
  XOR U4959 ( .A(n4381), .B(n4382), .Z(n4388) );
  XOR U4960 ( .A(n4387), .B(n4388), .Z(n4400) );
  XNOR U4961 ( .A(n4399), .B(n4400), .Z(n4331) );
  XNOR U4962 ( .A(n4332), .B(n4331), .Z(n4333) );
  XOR U4963 ( .A(n4334), .B(n4333), .Z(n4452) );
  XOR U4964 ( .A(n4451), .B(n4452), .Z(n4454) );
  XOR U4965 ( .A(n4453), .B(n4454), .Z(n4328) );
  NANDN U4966 ( .A(n4291), .B(n4290), .Z(n4295) );
  NAND U4967 ( .A(n4293), .B(n4292), .Z(n4294) );
  AND U4968 ( .A(n4295), .B(n4294), .Z(n4326) );
  NANDN U4969 ( .A(n4297), .B(n4296), .Z(n4301) );
  NANDN U4970 ( .A(n4299), .B(n4298), .Z(n4300) );
  AND U4971 ( .A(n4301), .B(n4300), .Z(n4325) );
  XNOR U4972 ( .A(n4326), .B(n4325), .Z(n4327) );
  XNOR U4973 ( .A(n4328), .B(n4327), .Z(n4319) );
  NANDN U4974 ( .A(n4303), .B(n4302), .Z(n4307) );
  NANDN U4975 ( .A(n4305), .B(n4304), .Z(n4306) );
  NAND U4976 ( .A(n4307), .B(n4306), .Z(n4320) );
  XOR U4977 ( .A(n4319), .B(n4320), .Z(n4322) );
  XNOR U4978 ( .A(n4321), .B(n4322), .Z(n4313) );
  XNOR U4979 ( .A(n4314), .B(n4313), .Z(n4315) );
  XNOR U4980 ( .A(n4316), .B(n4315), .Z(n4457) );
  XNOR U4981 ( .A(sreg[267]), .B(n4457), .Z(n4459) );
  NANDN U4982 ( .A(sreg[266]), .B(n4308), .Z(n4312) );
  NAND U4983 ( .A(n4310), .B(n4309), .Z(n4311) );
  NAND U4984 ( .A(n4312), .B(n4311), .Z(n4458) );
  XNOR U4985 ( .A(n4459), .B(n4458), .Z(c[267]) );
  NANDN U4986 ( .A(n4314), .B(n4313), .Z(n4318) );
  NANDN U4987 ( .A(n4316), .B(n4315), .Z(n4317) );
  AND U4988 ( .A(n4318), .B(n4317), .Z(n4465) );
  NANDN U4989 ( .A(n4320), .B(n4319), .Z(n4324) );
  NANDN U4990 ( .A(n4322), .B(n4321), .Z(n4323) );
  AND U4991 ( .A(n4324), .B(n4323), .Z(n4463) );
  NANDN U4992 ( .A(n4326), .B(n4325), .Z(n4330) );
  NANDN U4993 ( .A(n4328), .B(n4327), .Z(n4329) );
  AND U4994 ( .A(n4330), .B(n4329), .Z(n4471) );
  NANDN U4995 ( .A(n4332), .B(n4331), .Z(n4336) );
  NANDN U4996 ( .A(n4334), .B(n4333), .Z(n4335) );
  AND U4997 ( .A(n4336), .B(n4335), .Z(n4475) );
  NANDN U4998 ( .A(n4338), .B(n4337), .Z(n4342) );
  NAND U4999 ( .A(n4340), .B(n4339), .Z(n4341) );
  AND U5000 ( .A(n4342), .B(n4341), .Z(n4474) );
  XNOR U5001 ( .A(n4475), .B(n4474), .Z(n4477) );
  NANDN U5002 ( .A(n4344), .B(n4343), .Z(n4348) );
  NANDN U5003 ( .A(n4346), .B(n4345), .Z(n4347) );
  AND U5004 ( .A(n4348), .B(n4347), .Z(n4554) );
  NAND U5005 ( .A(n38385), .B(n4349), .Z(n4351) );
  XOR U5006 ( .A(b[27]), .B(a[18]), .Z(n4498) );
  NAND U5007 ( .A(n38343), .B(n4498), .Z(n4350) );
  AND U5008 ( .A(n4351), .B(n4350), .Z(n4561) );
  NAND U5009 ( .A(n183), .B(n4352), .Z(n4354) );
  XOR U5010 ( .A(b[5]), .B(a[40]), .Z(n4501) );
  NAND U5011 ( .A(n36296), .B(n4501), .Z(n4353) );
  AND U5012 ( .A(n4354), .B(n4353), .Z(n4559) );
  NAND U5013 ( .A(n190), .B(n4355), .Z(n4357) );
  XOR U5014 ( .A(b[19]), .B(a[26]), .Z(n4504) );
  NAND U5015 ( .A(n37821), .B(n4504), .Z(n4356) );
  NAND U5016 ( .A(n4357), .B(n4356), .Z(n4558) );
  XNOR U5017 ( .A(n4559), .B(n4558), .Z(n4560) );
  XNOR U5018 ( .A(n4561), .B(n4560), .Z(n4552) );
  NAND U5019 ( .A(n38470), .B(n4358), .Z(n4360) );
  XOR U5020 ( .A(b[31]), .B(a[14]), .Z(n4507) );
  NAND U5021 ( .A(n38453), .B(n4507), .Z(n4359) );
  AND U5022 ( .A(n4360), .B(n4359), .Z(n4519) );
  NAND U5023 ( .A(n181), .B(n4361), .Z(n4363) );
  XOR U5024 ( .A(b[3]), .B(a[42]), .Z(n4510) );
  NAND U5025 ( .A(n182), .B(n4510), .Z(n4362) );
  AND U5026 ( .A(n4363), .B(n4362), .Z(n4517) );
  NAND U5027 ( .A(n189), .B(n4364), .Z(n4366) );
  XOR U5028 ( .A(b[17]), .B(a[28]), .Z(n4513) );
  NAND U5029 ( .A(n37652), .B(n4513), .Z(n4365) );
  NAND U5030 ( .A(n4366), .B(n4365), .Z(n4516) );
  XNOR U5031 ( .A(n4517), .B(n4516), .Z(n4518) );
  XOR U5032 ( .A(n4519), .B(n4518), .Z(n4553) );
  XOR U5033 ( .A(n4552), .B(n4553), .Z(n4555) );
  XOR U5034 ( .A(n4554), .B(n4555), .Z(n4487) );
  NANDN U5035 ( .A(n4368), .B(n4367), .Z(n4372) );
  NANDN U5036 ( .A(n4370), .B(n4369), .Z(n4371) );
  AND U5037 ( .A(n4372), .B(n4371), .Z(n4540) );
  NANDN U5038 ( .A(n4374), .B(n4373), .Z(n4378) );
  NANDN U5039 ( .A(n4376), .B(n4375), .Z(n4377) );
  NAND U5040 ( .A(n4378), .B(n4377), .Z(n4541) );
  XNOR U5041 ( .A(n4540), .B(n4541), .Z(n4542) );
  NANDN U5042 ( .A(n4380), .B(n4379), .Z(n4384) );
  NANDN U5043 ( .A(n4382), .B(n4381), .Z(n4383) );
  NAND U5044 ( .A(n4384), .B(n4383), .Z(n4543) );
  XNOR U5045 ( .A(n4542), .B(n4543), .Z(n4486) );
  XNOR U5046 ( .A(n4487), .B(n4486), .Z(n4489) );
  NANDN U5047 ( .A(n4386), .B(n4385), .Z(n4390) );
  NANDN U5048 ( .A(n4388), .B(n4387), .Z(n4389) );
  AND U5049 ( .A(n4390), .B(n4389), .Z(n4488) );
  XOR U5050 ( .A(n4489), .B(n4488), .Z(n4603) );
  NANDN U5051 ( .A(n4392), .B(n4391), .Z(n4396) );
  NANDN U5052 ( .A(n4394), .B(n4393), .Z(n4395) );
  AND U5053 ( .A(n4396), .B(n4395), .Z(n4600) );
  NANDN U5054 ( .A(n4398), .B(n4397), .Z(n4402) );
  NANDN U5055 ( .A(n4400), .B(n4399), .Z(n4401) );
  AND U5056 ( .A(n4402), .B(n4401), .Z(n4483) );
  NANDN U5057 ( .A(n4404), .B(n4403), .Z(n4408) );
  OR U5058 ( .A(n4406), .B(n4405), .Z(n4407) );
  AND U5059 ( .A(n4408), .B(n4407), .Z(n4481) );
  NANDN U5060 ( .A(n4410), .B(n4409), .Z(n4414) );
  NANDN U5061 ( .A(n4412), .B(n4411), .Z(n4413) );
  AND U5062 ( .A(n4414), .B(n4413), .Z(n4547) );
  NANDN U5063 ( .A(n4416), .B(n4415), .Z(n4420) );
  NANDN U5064 ( .A(n4418), .B(n4417), .Z(n4419) );
  NAND U5065 ( .A(n4420), .B(n4419), .Z(n4546) );
  XNOR U5066 ( .A(n4547), .B(n4546), .Z(n4548) );
  NAND U5067 ( .A(b[0]), .B(a[44]), .Z(n4421) );
  XNOR U5068 ( .A(b[1]), .B(n4421), .Z(n4423) );
  NANDN U5069 ( .A(b[0]), .B(a[43]), .Z(n4422) );
  NAND U5070 ( .A(n4423), .B(n4422), .Z(n4495) );
  NAND U5071 ( .A(n194), .B(n4424), .Z(n4426) );
  XOR U5072 ( .A(b[29]), .B(a[16]), .Z(n4573) );
  NAND U5073 ( .A(n38456), .B(n4573), .Z(n4425) );
  AND U5074 ( .A(n4426), .B(n4425), .Z(n4493) );
  AND U5075 ( .A(b[31]), .B(a[12]), .Z(n4492) );
  XNOR U5076 ( .A(n4493), .B(n4492), .Z(n4494) );
  XNOR U5077 ( .A(n4495), .B(n4494), .Z(n4534) );
  NAND U5078 ( .A(n38185), .B(n4427), .Z(n4429) );
  XOR U5079 ( .A(b[23]), .B(a[22]), .Z(n4576) );
  NAND U5080 ( .A(n38132), .B(n4576), .Z(n4428) );
  AND U5081 ( .A(n4429), .B(n4428), .Z(n4567) );
  NAND U5082 ( .A(n184), .B(n4430), .Z(n4432) );
  XOR U5083 ( .A(b[7]), .B(a[38]), .Z(n4579) );
  NAND U5084 ( .A(n36592), .B(n4579), .Z(n4431) );
  AND U5085 ( .A(n4432), .B(n4431), .Z(n4565) );
  NAND U5086 ( .A(n38289), .B(n4433), .Z(n4435) );
  XOR U5087 ( .A(b[25]), .B(a[20]), .Z(n4582) );
  NAND U5088 ( .A(n38247), .B(n4582), .Z(n4434) );
  NAND U5089 ( .A(n4435), .B(n4434), .Z(n4564) );
  XNOR U5090 ( .A(n4565), .B(n4564), .Z(n4566) );
  XOR U5091 ( .A(n4567), .B(n4566), .Z(n4535) );
  XNOR U5092 ( .A(n4534), .B(n4535), .Z(n4536) );
  NAND U5093 ( .A(n187), .B(n4436), .Z(n4438) );
  XOR U5094 ( .A(b[13]), .B(a[32]), .Z(n4585) );
  NAND U5095 ( .A(n37295), .B(n4585), .Z(n4437) );
  AND U5096 ( .A(n4438), .B(n4437), .Z(n4529) );
  NAND U5097 ( .A(n186), .B(n4439), .Z(n4441) );
  XOR U5098 ( .A(b[11]), .B(a[34]), .Z(n4588) );
  NAND U5099 ( .A(n37097), .B(n4588), .Z(n4440) );
  NAND U5100 ( .A(n4441), .B(n4440), .Z(n4528) );
  XNOR U5101 ( .A(n4529), .B(n4528), .Z(n4530) );
  NAND U5102 ( .A(n188), .B(n4442), .Z(n4444) );
  XOR U5103 ( .A(b[15]), .B(a[30]), .Z(n4591) );
  NAND U5104 ( .A(n37382), .B(n4591), .Z(n4443) );
  AND U5105 ( .A(n4444), .B(n4443), .Z(n4525) );
  NAND U5106 ( .A(n38064), .B(n4445), .Z(n4447) );
  XOR U5107 ( .A(b[21]), .B(a[24]), .Z(n4594) );
  NAND U5108 ( .A(n37993), .B(n4594), .Z(n4446) );
  AND U5109 ( .A(n4447), .B(n4446), .Z(n4523) );
  NAND U5110 ( .A(n185), .B(n4448), .Z(n4450) );
  XOR U5111 ( .A(b[9]), .B(a[36]), .Z(n4597) );
  NAND U5112 ( .A(n36805), .B(n4597), .Z(n4449) );
  NAND U5113 ( .A(n4450), .B(n4449), .Z(n4522) );
  XNOR U5114 ( .A(n4523), .B(n4522), .Z(n4524) );
  XOR U5115 ( .A(n4525), .B(n4524), .Z(n4531) );
  XOR U5116 ( .A(n4530), .B(n4531), .Z(n4537) );
  XOR U5117 ( .A(n4536), .B(n4537), .Z(n4549) );
  XNOR U5118 ( .A(n4548), .B(n4549), .Z(n4480) );
  XNOR U5119 ( .A(n4481), .B(n4480), .Z(n4482) );
  XOR U5120 ( .A(n4483), .B(n4482), .Z(n4601) );
  XNOR U5121 ( .A(n4600), .B(n4601), .Z(n4602) );
  XNOR U5122 ( .A(n4603), .B(n4602), .Z(n4476) );
  XOR U5123 ( .A(n4477), .B(n4476), .Z(n4469) );
  NANDN U5124 ( .A(n4452), .B(n4451), .Z(n4456) );
  OR U5125 ( .A(n4454), .B(n4453), .Z(n4455) );
  AND U5126 ( .A(n4456), .B(n4455), .Z(n4468) );
  XNOR U5127 ( .A(n4469), .B(n4468), .Z(n4470) );
  XNOR U5128 ( .A(n4471), .B(n4470), .Z(n4462) );
  XNOR U5129 ( .A(n4463), .B(n4462), .Z(n4464) );
  XNOR U5130 ( .A(n4465), .B(n4464), .Z(n4606) );
  XNOR U5131 ( .A(sreg[268]), .B(n4606), .Z(n4608) );
  NANDN U5132 ( .A(sreg[267]), .B(n4457), .Z(n4461) );
  NAND U5133 ( .A(n4459), .B(n4458), .Z(n4460) );
  NAND U5134 ( .A(n4461), .B(n4460), .Z(n4607) );
  XNOR U5135 ( .A(n4608), .B(n4607), .Z(c[268]) );
  NANDN U5136 ( .A(n4463), .B(n4462), .Z(n4467) );
  NANDN U5137 ( .A(n4465), .B(n4464), .Z(n4466) );
  AND U5138 ( .A(n4467), .B(n4466), .Z(n4614) );
  NANDN U5139 ( .A(n4469), .B(n4468), .Z(n4473) );
  NANDN U5140 ( .A(n4471), .B(n4470), .Z(n4472) );
  AND U5141 ( .A(n4473), .B(n4472), .Z(n4612) );
  NANDN U5142 ( .A(n4475), .B(n4474), .Z(n4479) );
  NAND U5143 ( .A(n4477), .B(n4476), .Z(n4478) );
  AND U5144 ( .A(n4479), .B(n4478), .Z(n4619) );
  NANDN U5145 ( .A(n4481), .B(n4480), .Z(n4485) );
  NANDN U5146 ( .A(n4483), .B(n4482), .Z(n4484) );
  AND U5147 ( .A(n4485), .B(n4484), .Z(n4750) );
  NANDN U5148 ( .A(n4487), .B(n4486), .Z(n4491) );
  NAND U5149 ( .A(n4489), .B(n4488), .Z(n4490) );
  AND U5150 ( .A(n4491), .B(n4490), .Z(n4749) );
  XNOR U5151 ( .A(n4750), .B(n4749), .Z(n4752) );
  NANDN U5152 ( .A(n4493), .B(n4492), .Z(n4497) );
  NANDN U5153 ( .A(n4495), .B(n4494), .Z(n4496) );
  AND U5154 ( .A(n4497), .B(n4496), .Z(n4697) );
  NAND U5155 ( .A(n38385), .B(n4498), .Z(n4500) );
  XOR U5156 ( .A(b[27]), .B(a[19]), .Z(n4641) );
  NAND U5157 ( .A(n38343), .B(n4641), .Z(n4499) );
  AND U5158 ( .A(n4500), .B(n4499), .Z(n4704) );
  NAND U5159 ( .A(n183), .B(n4501), .Z(n4503) );
  XOR U5160 ( .A(b[5]), .B(a[41]), .Z(n4644) );
  NAND U5161 ( .A(n36296), .B(n4644), .Z(n4502) );
  AND U5162 ( .A(n4503), .B(n4502), .Z(n4702) );
  NAND U5163 ( .A(n190), .B(n4504), .Z(n4506) );
  XOR U5164 ( .A(b[19]), .B(a[27]), .Z(n4647) );
  NAND U5165 ( .A(n37821), .B(n4647), .Z(n4505) );
  NAND U5166 ( .A(n4506), .B(n4505), .Z(n4701) );
  XNOR U5167 ( .A(n4702), .B(n4701), .Z(n4703) );
  XNOR U5168 ( .A(n4704), .B(n4703), .Z(n4695) );
  NAND U5169 ( .A(n38470), .B(n4507), .Z(n4509) );
  XOR U5170 ( .A(b[31]), .B(a[15]), .Z(n4650) );
  NAND U5171 ( .A(n38453), .B(n4650), .Z(n4508) );
  AND U5172 ( .A(n4509), .B(n4508), .Z(n4662) );
  NAND U5173 ( .A(n181), .B(n4510), .Z(n4512) );
  XOR U5174 ( .A(b[3]), .B(a[43]), .Z(n4653) );
  NAND U5175 ( .A(n182), .B(n4653), .Z(n4511) );
  AND U5176 ( .A(n4512), .B(n4511), .Z(n4660) );
  NAND U5177 ( .A(n189), .B(n4513), .Z(n4515) );
  XOR U5178 ( .A(b[17]), .B(a[29]), .Z(n4656) );
  NAND U5179 ( .A(n37652), .B(n4656), .Z(n4514) );
  NAND U5180 ( .A(n4515), .B(n4514), .Z(n4659) );
  XNOR U5181 ( .A(n4660), .B(n4659), .Z(n4661) );
  XOR U5182 ( .A(n4662), .B(n4661), .Z(n4696) );
  XOR U5183 ( .A(n4695), .B(n4696), .Z(n4698) );
  XOR U5184 ( .A(n4697), .B(n4698), .Z(n4630) );
  NANDN U5185 ( .A(n4517), .B(n4516), .Z(n4521) );
  NANDN U5186 ( .A(n4519), .B(n4518), .Z(n4520) );
  AND U5187 ( .A(n4521), .B(n4520), .Z(n4683) );
  NANDN U5188 ( .A(n4523), .B(n4522), .Z(n4527) );
  NANDN U5189 ( .A(n4525), .B(n4524), .Z(n4526) );
  NAND U5190 ( .A(n4527), .B(n4526), .Z(n4684) );
  XNOR U5191 ( .A(n4683), .B(n4684), .Z(n4685) );
  NANDN U5192 ( .A(n4529), .B(n4528), .Z(n4533) );
  NANDN U5193 ( .A(n4531), .B(n4530), .Z(n4532) );
  NAND U5194 ( .A(n4533), .B(n4532), .Z(n4686) );
  XNOR U5195 ( .A(n4685), .B(n4686), .Z(n4629) );
  XNOR U5196 ( .A(n4630), .B(n4629), .Z(n4632) );
  NANDN U5197 ( .A(n4535), .B(n4534), .Z(n4539) );
  NANDN U5198 ( .A(n4537), .B(n4536), .Z(n4538) );
  AND U5199 ( .A(n4539), .B(n4538), .Z(n4631) );
  XOR U5200 ( .A(n4632), .B(n4631), .Z(n4746) );
  NANDN U5201 ( .A(n4541), .B(n4540), .Z(n4545) );
  NANDN U5202 ( .A(n4543), .B(n4542), .Z(n4544) );
  AND U5203 ( .A(n4545), .B(n4544), .Z(n4743) );
  NANDN U5204 ( .A(n4547), .B(n4546), .Z(n4551) );
  NANDN U5205 ( .A(n4549), .B(n4548), .Z(n4550) );
  AND U5206 ( .A(n4551), .B(n4550), .Z(n4626) );
  NANDN U5207 ( .A(n4553), .B(n4552), .Z(n4557) );
  OR U5208 ( .A(n4555), .B(n4554), .Z(n4556) );
  AND U5209 ( .A(n4557), .B(n4556), .Z(n4624) );
  NANDN U5210 ( .A(n4559), .B(n4558), .Z(n4563) );
  NANDN U5211 ( .A(n4561), .B(n4560), .Z(n4562) );
  AND U5212 ( .A(n4563), .B(n4562), .Z(n4690) );
  NANDN U5213 ( .A(n4565), .B(n4564), .Z(n4569) );
  NANDN U5214 ( .A(n4567), .B(n4566), .Z(n4568) );
  NAND U5215 ( .A(n4569), .B(n4568), .Z(n4689) );
  XNOR U5216 ( .A(n4690), .B(n4689), .Z(n4691) );
  NAND U5217 ( .A(b[0]), .B(a[45]), .Z(n4570) );
  XNOR U5218 ( .A(b[1]), .B(n4570), .Z(n4572) );
  NANDN U5219 ( .A(b[0]), .B(a[44]), .Z(n4571) );
  NAND U5220 ( .A(n4572), .B(n4571), .Z(n4638) );
  NAND U5221 ( .A(n194), .B(n4573), .Z(n4575) );
  XOR U5222 ( .A(b[29]), .B(a[17]), .Z(n4713) );
  NAND U5223 ( .A(n38456), .B(n4713), .Z(n4574) );
  AND U5224 ( .A(n4575), .B(n4574), .Z(n4636) );
  AND U5225 ( .A(b[31]), .B(a[13]), .Z(n4635) );
  XNOR U5226 ( .A(n4636), .B(n4635), .Z(n4637) );
  XNOR U5227 ( .A(n4638), .B(n4637), .Z(n4677) );
  NAND U5228 ( .A(n38185), .B(n4576), .Z(n4578) );
  XOR U5229 ( .A(b[23]), .B(a[23]), .Z(n4719) );
  NAND U5230 ( .A(n38132), .B(n4719), .Z(n4577) );
  AND U5231 ( .A(n4578), .B(n4577), .Z(n4710) );
  NAND U5232 ( .A(n184), .B(n4579), .Z(n4581) );
  XOR U5233 ( .A(b[7]), .B(a[39]), .Z(n4722) );
  NAND U5234 ( .A(n36592), .B(n4722), .Z(n4580) );
  AND U5235 ( .A(n4581), .B(n4580), .Z(n4708) );
  NAND U5236 ( .A(n38289), .B(n4582), .Z(n4584) );
  XOR U5237 ( .A(b[25]), .B(a[21]), .Z(n4725) );
  NAND U5238 ( .A(n38247), .B(n4725), .Z(n4583) );
  NAND U5239 ( .A(n4584), .B(n4583), .Z(n4707) );
  XNOR U5240 ( .A(n4708), .B(n4707), .Z(n4709) );
  XOR U5241 ( .A(n4710), .B(n4709), .Z(n4678) );
  XNOR U5242 ( .A(n4677), .B(n4678), .Z(n4679) );
  NAND U5243 ( .A(n187), .B(n4585), .Z(n4587) );
  XOR U5244 ( .A(b[13]), .B(a[33]), .Z(n4728) );
  NAND U5245 ( .A(n37295), .B(n4728), .Z(n4586) );
  AND U5246 ( .A(n4587), .B(n4586), .Z(n4672) );
  NAND U5247 ( .A(n186), .B(n4588), .Z(n4590) );
  XOR U5248 ( .A(b[11]), .B(a[35]), .Z(n4731) );
  NAND U5249 ( .A(n37097), .B(n4731), .Z(n4589) );
  NAND U5250 ( .A(n4590), .B(n4589), .Z(n4671) );
  XNOR U5251 ( .A(n4672), .B(n4671), .Z(n4673) );
  NAND U5252 ( .A(n188), .B(n4591), .Z(n4593) );
  XOR U5253 ( .A(b[15]), .B(a[31]), .Z(n4734) );
  NAND U5254 ( .A(n37382), .B(n4734), .Z(n4592) );
  AND U5255 ( .A(n4593), .B(n4592), .Z(n4668) );
  NAND U5256 ( .A(n38064), .B(n4594), .Z(n4596) );
  XOR U5257 ( .A(b[21]), .B(a[25]), .Z(n4737) );
  NAND U5258 ( .A(n37993), .B(n4737), .Z(n4595) );
  AND U5259 ( .A(n4596), .B(n4595), .Z(n4666) );
  NAND U5260 ( .A(n185), .B(n4597), .Z(n4599) );
  XOR U5261 ( .A(b[9]), .B(a[37]), .Z(n4740) );
  NAND U5262 ( .A(n36805), .B(n4740), .Z(n4598) );
  NAND U5263 ( .A(n4599), .B(n4598), .Z(n4665) );
  XNOR U5264 ( .A(n4666), .B(n4665), .Z(n4667) );
  XOR U5265 ( .A(n4668), .B(n4667), .Z(n4674) );
  XOR U5266 ( .A(n4673), .B(n4674), .Z(n4680) );
  XOR U5267 ( .A(n4679), .B(n4680), .Z(n4692) );
  XNOR U5268 ( .A(n4691), .B(n4692), .Z(n4623) );
  XNOR U5269 ( .A(n4624), .B(n4623), .Z(n4625) );
  XOR U5270 ( .A(n4626), .B(n4625), .Z(n4744) );
  XNOR U5271 ( .A(n4743), .B(n4744), .Z(n4745) );
  XNOR U5272 ( .A(n4746), .B(n4745), .Z(n4751) );
  XOR U5273 ( .A(n4752), .B(n4751), .Z(n4618) );
  NANDN U5274 ( .A(n4601), .B(n4600), .Z(n4605) );
  NANDN U5275 ( .A(n4603), .B(n4602), .Z(n4604) );
  AND U5276 ( .A(n4605), .B(n4604), .Z(n4617) );
  XOR U5277 ( .A(n4618), .B(n4617), .Z(n4620) );
  XNOR U5278 ( .A(n4619), .B(n4620), .Z(n4611) );
  XNOR U5279 ( .A(n4612), .B(n4611), .Z(n4613) );
  XNOR U5280 ( .A(n4614), .B(n4613), .Z(n4755) );
  XNOR U5281 ( .A(sreg[269]), .B(n4755), .Z(n4757) );
  NANDN U5282 ( .A(sreg[268]), .B(n4606), .Z(n4610) );
  NAND U5283 ( .A(n4608), .B(n4607), .Z(n4609) );
  NAND U5284 ( .A(n4610), .B(n4609), .Z(n4756) );
  XNOR U5285 ( .A(n4757), .B(n4756), .Z(c[269]) );
  NANDN U5286 ( .A(n4612), .B(n4611), .Z(n4616) );
  NANDN U5287 ( .A(n4614), .B(n4613), .Z(n4615) );
  AND U5288 ( .A(n4616), .B(n4615), .Z(n4763) );
  NANDN U5289 ( .A(n4618), .B(n4617), .Z(n4622) );
  NANDN U5290 ( .A(n4620), .B(n4619), .Z(n4621) );
  AND U5291 ( .A(n4622), .B(n4621), .Z(n4761) );
  NANDN U5292 ( .A(n4624), .B(n4623), .Z(n4628) );
  NANDN U5293 ( .A(n4626), .B(n4625), .Z(n4627) );
  AND U5294 ( .A(n4628), .B(n4627), .Z(n4773) );
  NANDN U5295 ( .A(n4630), .B(n4629), .Z(n4634) );
  NAND U5296 ( .A(n4632), .B(n4631), .Z(n4633) );
  AND U5297 ( .A(n4634), .B(n4633), .Z(n4772) );
  XNOR U5298 ( .A(n4773), .B(n4772), .Z(n4775) );
  NANDN U5299 ( .A(n4636), .B(n4635), .Z(n4640) );
  NANDN U5300 ( .A(n4638), .B(n4637), .Z(n4639) );
  AND U5301 ( .A(n4640), .B(n4639), .Z(n4852) );
  NAND U5302 ( .A(n38385), .B(n4641), .Z(n4643) );
  XOR U5303 ( .A(b[27]), .B(a[20]), .Z(n4796) );
  NAND U5304 ( .A(n38343), .B(n4796), .Z(n4642) );
  AND U5305 ( .A(n4643), .B(n4642), .Z(n4859) );
  NAND U5306 ( .A(n183), .B(n4644), .Z(n4646) );
  XOR U5307 ( .A(b[5]), .B(a[42]), .Z(n4799) );
  NAND U5308 ( .A(n36296), .B(n4799), .Z(n4645) );
  AND U5309 ( .A(n4646), .B(n4645), .Z(n4857) );
  NAND U5310 ( .A(n190), .B(n4647), .Z(n4649) );
  XOR U5311 ( .A(b[19]), .B(a[28]), .Z(n4802) );
  NAND U5312 ( .A(n37821), .B(n4802), .Z(n4648) );
  NAND U5313 ( .A(n4649), .B(n4648), .Z(n4856) );
  XNOR U5314 ( .A(n4857), .B(n4856), .Z(n4858) );
  XNOR U5315 ( .A(n4859), .B(n4858), .Z(n4850) );
  NAND U5316 ( .A(n38470), .B(n4650), .Z(n4652) );
  XOR U5317 ( .A(b[31]), .B(a[16]), .Z(n4805) );
  NAND U5318 ( .A(n38453), .B(n4805), .Z(n4651) );
  AND U5319 ( .A(n4652), .B(n4651), .Z(n4817) );
  NAND U5320 ( .A(n181), .B(n4653), .Z(n4655) );
  XOR U5321 ( .A(b[3]), .B(a[44]), .Z(n4808) );
  NAND U5322 ( .A(n182), .B(n4808), .Z(n4654) );
  AND U5323 ( .A(n4655), .B(n4654), .Z(n4815) );
  NAND U5324 ( .A(n189), .B(n4656), .Z(n4658) );
  XOR U5325 ( .A(b[17]), .B(a[30]), .Z(n4811) );
  NAND U5326 ( .A(n37652), .B(n4811), .Z(n4657) );
  NAND U5327 ( .A(n4658), .B(n4657), .Z(n4814) );
  XNOR U5328 ( .A(n4815), .B(n4814), .Z(n4816) );
  XOR U5329 ( .A(n4817), .B(n4816), .Z(n4851) );
  XOR U5330 ( .A(n4850), .B(n4851), .Z(n4853) );
  XOR U5331 ( .A(n4852), .B(n4853), .Z(n4785) );
  NANDN U5332 ( .A(n4660), .B(n4659), .Z(n4664) );
  NANDN U5333 ( .A(n4662), .B(n4661), .Z(n4663) );
  AND U5334 ( .A(n4664), .B(n4663), .Z(n4838) );
  NANDN U5335 ( .A(n4666), .B(n4665), .Z(n4670) );
  NANDN U5336 ( .A(n4668), .B(n4667), .Z(n4669) );
  NAND U5337 ( .A(n4670), .B(n4669), .Z(n4839) );
  XNOR U5338 ( .A(n4838), .B(n4839), .Z(n4840) );
  NANDN U5339 ( .A(n4672), .B(n4671), .Z(n4676) );
  NANDN U5340 ( .A(n4674), .B(n4673), .Z(n4675) );
  NAND U5341 ( .A(n4676), .B(n4675), .Z(n4841) );
  XNOR U5342 ( .A(n4840), .B(n4841), .Z(n4784) );
  XNOR U5343 ( .A(n4785), .B(n4784), .Z(n4787) );
  NANDN U5344 ( .A(n4678), .B(n4677), .Z(n4682) );
  NANDN U5345 ( .A(n4680), .B(n4679), .Z(n4681) );
  AND U5346 ( .A(n4682), .B(n4681), .Z(n4786) );
  XOR U5347 ( .A(n4787), .B(n4786), .Z(n4901) );
  NANDN U5348 ( .A(n4684), .B(n4683), .Z(n4688) );
  NANDN U5349 ( .A(n4686), .B(n4685), .Z(n4687) );
  AND U5350 ( .A(n4688), .B(n4687), .Z(n4898) );
  NANDN U5351 ( .A(n4690), .B(n4689), .Z(n4694) );
  NANDN U5352 ( .A(n4692), .B(n4691), .Z(n4693) );
  AND U5353 ( .A(n4694), .B(n4693), .Z(n4781) );
  NANDN U5354 ( .A(n4696), .B(n4695), .Z(n4700) );
  OR U5355 ( .A(n4698), .B(n4697), .Z(n4699) );
  AND U5356 ( .A(n4700), .B(n4699), .Z(n4779) );
  NANDN U5357 ( .A(n4702), .B(n4701), .Z(n4706) );
  NANDN U5358 ( .A(n4704), .B(n4703), .Z(n4705) );
  AND U5359 ( .A(n4706), .B(n4705), .Z(n4845) );
  NANDN U5360 ( .A(n4708), .B(n4707), .Z(n4712) );
  NANDN U5361 ( .A(n4710), .B(n4709), .Z(n4711) );
  NAND U5362 ( .A(n4712), .B(n4711), .Z(n4844) );
  XNOR U5363 ( .A(n4845), .B(n4844), .Z(n4846) );
  NAND U5364 ( .A(n194), .B(n4713), .Z(n4715) );
  XOR U5365 ( .A(b[29]), .B(a[18]), .Z(n4871) );
  NAND U5366 ( .A(n38456), .B(n4871), .Z(n4714) );
  AND U5367 ( .A(n4715), .B(n4714), .Z(n4791) );
  AND U5368 ( .A(b[31]), .B(a[14]), .Z(n4790) );
  XNOR U5369 ( .A(n4791), .B(n4790), .Z(n4792) );
  NAND U5370 ( .A(b[0]), .B(a[46]), .Z(n4716) );
  XNOR U5371 ( .A(b[1]), .B(n4716), .Z(n4718) );
  NANDN U5372 ( .A(b[0]), .B(a[45]), .Z(n4717) );
  NAND U5373 ( .A(n4718), .B(n4717), .Z(n4793) );
  XNOR U5374 ( .A(n4792), .B(n4793), .Z(n4832) );
  NAND U5375 ( .A(n38185), .B(n4719), .Z(n4721) );
  XOR U5376 ( .A(b[23]), .B(a[24]), .Z(n4874) );
  NAND U5377 ( .A(n38132), .B(n4874), .Z(n4720) );
  AND U5378 ( .A(n4721), .B(n4720), .Z(n4865) );
  NAND U5379 ( .A(n184), .B(n4722), .Z(n4724) );
  XOR U5380 ( .A(b[7]), .B(a[40]), .Z(n4877) );
  NAND U5381 ( .A(n36592), .B(n4877), .Z(n4723) );
  AND U5382 ( .A(n4724), .B(n4723), .Z(n4863) );
  NAND U5383 ( .A(n38289), .B(n4725), .Z(n4727) );
  XOR U5384 ( .A(b[25]), .B(a[22]), .Z(n4880) );
  NAND U5385 ( .A(n38247), .B(n4880), .Z(n4726) );
  NAND U5386 ( .A(n4727), .B(n4726), .Z(n4862) );
  XNOR U5387 ( .A(n4863), .B(n4862), .Z(n4864) );
  XOR U5388 ( .A(n4865), .B(n4864), .Z(n4833) );
  XNOR U5389 ( .A(n4832), .B(n4833), .Z(n4834) );
  NAND U5390 ( .A(n187), .B(n4728), .Z(n4730) );
  XOR U5391 ( .A(b[13]), .B(a[34]), .Z(n4883) );
  NAND U5392 ( .A(n37295), .B(n4883), .Z(n4729) );
  AND U5393 ( .A(n4730), .B(n4729), .Z(n4827) );
  NAND U5394 ( .A(n186), .B(n4731), .Z(n4733) );
  XOR U5395 ( .A(b[11]), .B(a[36]), .Z(n4886) );
  NAND U5396 ( .A(n37097), .B(n4886), .Z(n4732) );
  NAND U5397 ( .A(n4733), .B(n4732), .Z(n4826) );
  XNOR U5398 ( .A(n4827), .B(n4826), .Z(n4828) );
  NAND U5399 ( .A(n188), .B(n4734), .Z(n4736) );
  XOR U5400 ( .A(b[15]), .B(a[32]), .Z(n4889) );
  NAND U5401 ( .A(n37382), .B(n4889), .Z(n4735) );
  AND U5402 ( .A(n4736), .B(n4735), .Z(n4823) );
  NAND U5403 ( .A(n38064), .B(n4737), .Z(n4739) );
  XOR U5404 ( .A(b[21]), .B(a[26]), .Z(n4892) );
  NAND U5405 ( .A(n37993), .B(n4892), .Z(n4738) );
  AND U5406 ( .A(n4739), .B(n4738), .Z(n4821) );
  NAND U5407 ( .A(n185), .B(n4740), .Z(n4742) );
  XOR U5408 ( .A(b[9]), .B(a[38]), .Z(n4895) );
  NAND U5409 ( .A(n36805), .B(n4895), .Z(n4741) );
  NAND U5410 ( .A(n4742), .B(n4741), .Z(n4820) );
  XNOR U5411 ( .A(n4821), .B(n4820), .Z(n4822) );
  XOR U5412 ( .A(n4823), .B(n4822), .Z(n4829) );
  XOR U5413 ( .A(n4828), .B(n4829), .Z(n4835) );
  XOR U5414 ( .A(n4834), .B(n4835), .Z(n4847) );
  XNOR U5415 ( .A(n4846), .B(n4847), .Z(n4778) );
  XNOR U5416 ( .A(n4779), .B(n4778), .Z(n4780) );
  XOR U5417 ( .A(n4781), .B(n4780), .Z(n4899) );
  XNOR U5418 ( .A(n4898), .B(n4899), .Z(n4900) );
  XNOR U5419 ( .A(n4901), .B(n4900), .Z(n4774) );
  XOR U5420 ( .A(n4775), .B(n4774), .Z(n4767) );
  NANDN U5421 ( .A(n4744), .B(n4743), .Z(n4748) );
  NANDN U5422 ( .A(n4746), .B(n4745), .Z(n4747) );
  AND U5423 ( .A(n4748), .B(n4747), .Z(n4766) );
  XNOR U5424 ( .A(n4767), .B(n4766), .Z(n4768) );
  NANDN U5425 ( .A(n4750), .B(n4749), .Z(n4754) );
  NAND U5426 ( .A(n4752), .B(n4751), .Z(n4753) );
  NAND U5427 ( .A(n4754), .B(n4753), .Z(n4769) );
  XNOR U5428 ( .A(n4768), .B(n4769), .Z(n4760) );
  XNOR U5429 ( .A(n4761), .B(n4760), .Z(n4762) );
  XNOR U5430 ( .A(n4763), .B(n4762), .Z(n4904) );
  XNOR U5431 ( .A(sreg[270]), .B(n4904), .Z(n4906) );
  NANDN U5432 ( .A(sreg[269]), .B(n4755), .Z(n4759) );
  NAND U5433 ( .A(n4757), .B(n4756), .Z(n4758) );
  NAND U5434 ( .A(n4759), .B(n4758), .Z(n4905) );
  XNOR U5435 ( .A(n4906), .B(n4905), .Z(c[270]) );
  NANDN U5436 ( .A(n4761), .B(n4760), .Z(n4765) );
  NANDN U5437 ( .A(n4763), .B(n4762), .Z(n4764) );
  AND U5438 ( .A(n4765), .B(n4764), .Z(n4912) );
  NANDN U5439 ( .A(n4767), .B(n4766), .Z(n4771) );
  NANDN U5440 ( .A(n4769), .B(n4768), .Z(n4770) );
  AND U5441 ( .A(n4771), .B(n4770), .Z(n4910) );
  NANDN U5442 ( .A(n4773), .B(n4772), .Z(n4777) );
  NAND U5443 ( .A(n4775), .B(n4774), .Z(n4776) );
  AND U5444 ( .A(n4777), .B(n4776), .Z(n4917) );
  NANDN U5445 ( .A(n4779), .B(n4778), .Z(n4783) );
  NANDN U5446 ( .A(n4781), .B(n4780), .Z(n4782) );
  AND U5447 ( .A(n4783), .B(n4782), .Z(n4922) );
  NANDN U5448 ( .A(n4785), .B(n4784), .Z(n4789) );
  NAND U5449 ( .A(n4787), .B(n4786), .Z(n4788) );
  AND U5450 ( .A(n4789), .B(n4788), .Z(n4921) );
  XNOR U5451 ( .A(n4922), .B(n4921), .Z(n4924) );
  NANDN U5452 ( .A(n4791), .B(n4790), .Z(n4795) );
  NANDN U5453 ( .A(n4793), .B(n4792), .Z(n4794) );
  AND U5454 ( .A(n4795), .B(n4794), .Z(n4999) );
  NAND U5455 ( .A(n38385), .B(n4796), .Z(n4798) );
  XOR U5456 ( .A(b[27]), .B(a[21]), .Z(n4945) );
  NAND U5457 ( .A(n38343), .B(n4945), .Z(n4797) );
  AND U5458 ( .A(n4798), .B(n4797), .Z(n5006) );
  NAND U5459 ( .A(n183), .B(n4799), .Z(n4801) );
  XOR U5460 ( .A(b[5]), .B(a[43]), .Z(n4948) );
  NAND U5461 ( .A(n36296), .B(n4948), .Z(n4800) );
  AND U5462 ( .A(n4801), .B(n4800), .Z(n5004) );
  NAND U5463 ( .A(n190), .B(n4802), .Z(n4804) );
  XOR U5464 ( .A(b[19]), .B(a[29]), .Z(n4951) );
  NAND U5465 ( .A(n37821), .B(n4951), .Z(n4803) );
  NAND U5466 ( .A(n4804), .B(n4803), .Z(n5003) );
  XNOR U5467 ( .A(n5004), .B(n5003), .Z(n5005) );
  XNOR U5468 ( .A(n5006), .B(n5005), .Z(n4997) );
  NAND U5469 ( .A(n38470), .B(n4805), .Z(n4807) );
  XOR U5470 ( .A(b[31]), .B(a[17]), .Z(n4954) );
  NAND U5471 ( .A(n38453), .B(n4954), .Z(n4806) );
  AND U5472 ( .A(n4807), .B(n4806), .Z(n4966) );
  NAND U5473 ( .A(n181), .B(n4808), .Z(n4810) );
  XOR U5474 ( .A(b[3]), .B(a[45]), .Z(n4957) );
  NAND U5475 ( .A(n182), .B(n4957), .Z(n4809) );
  AND U5476 ( .A(n4810), .B(n4809), .Z(n4964) );
  NAND U5477 ( .A(n189), .B(n4811), .Z(n4813) );
  XOR U5478 ( .A(b[17]), .B(a[31]), .Z(n4960) );
  NAND U5479 ( .A(n37652), .B(n4960), .Z(n4812) );
  NAND U5480 ( .A(n4813), .B(n4812), .Z(n4963) );
  XNOR U5481 ( .A(n4964), .B(n4963), .Z(n4965) );
  XOR U5482 ( .A(n4966), .B(n4965), .Z(n4998) );
  XOR U5483 ( .A(n4997), .B(n4998), .Z(n5000) );
  XOR U5484 ( .A(n4999), .B(n5000), .Z(n4934) );
  NANDN U5485 ( .A(n4815), .B(n4814), .Z(n4819) );
  NANDN U5486 ( .A(n4817), .B(n4816), .Z(n4818) );
  AND U5487 ( .A(n4819), .B(n4818), .Z(n4987) );
  NANDN U5488 ( .A(n4821), .B(n4820), .Z(n4825) );
  NANDN U5489 ( .A(n4823), .B(n4822), .Z(n4824) );
  NAND U5490 ( .A(n4825), .B(n4824), .Z(n4988) );
  XNOR U5491 ( .A(n4987), .B(n4988), .Z(n4989) );
  NANDN U5492 ( .A(n4827), .B(n4826), .Z(n4831) );
  NANDN U5493 ( .A(n4829), .B(n4828), .Z(n4830) );
  NAND U5494 ( .A(n4831), .B(n4830), .Z(n4990) );
  XNOR U5495 ( .A(n4989), .B(n4990), .Z(n4933) );
  XNOR U5496 ( .A(n4934), .B(n4933), .Z(n4936) );
  NANDN U5497 ( .A(n4833), .B(n4832), .Z(n4837) );
  NANDN U5498 ( .A(n4835), .B(n4834), .Z(n4836) );
  AND U5499 ( .A(n4837), .B(n4836), .Z(n4935) );
  XOR U5500 ( .A(n4936), .B(n4935), .Z(n5048) );
  NANDN U5501 ( .A(n4839), .B(n4838), .Z(n4843) );
  NANDN U5502 ( .A(n4841), .B(n4840), .Z(n4842) );
  AND U5503 ( .A(n4843), .B(n4842), .Z(n5045) );
  NANDN U5504 ( .A(n4845), .B(n4844), .Z(n4849) );
  NANDN U5505 ( .A(n4847), .B(n4846), .Z(n4848) );
  AND U5506 ( .A(n4849), .B(n4848), .Z(n4930) );
  NANDN U5507 ( .A(n4851), .B(n4850), .Z(n4855) );
  OR U5508 ( .A(n4853), .B(n4852), .Z(n4854) );
  AND U5509 ( .A(n4855), .B(n4854), .Z(n4928) );
  NANDN U5510 ( .A(n4857), .B(n4856), .Z(n4861) );
  NANDN U5511 ( .A(n4859), .B(n4858), .Z(n4860) );
  AND U5512 ( .A(n4861), .B(n4860), .Z(n4994) );
  NANDN U5513 ( .A(n4863), .B(n4862), .Z(n4867) );
  NANDN U5514 ( .A(n4865), .B(n4864), .Z(n4866) );
  NAND U5515 ( .A(n4867), .B(n4866), .Z(n4993) );
  XNOR U5516 ( .A(n4994), .B(n4993), .Z(n4996) );
  NAND U5517 ( .A(b[0]), .B(a[47]), .Z(n4868) );
  XNOR U5518 ( .A(b[1]), .B(n4868), .Z(n4870) );
  NANDN U5519 ( .A(b[0]), .B(a[46]), .Z(n4869) );
  NAND U5520 ( .A(n4870), .B(n4869), .Z(n4942) );
  NAND U5521 ( .A(n194), .B(n4871), .Z(n4873) );
  XOR U5522 ( .A(b[29]), .B(a[19]), .Z(n5018) );
  NAND U5523 ( .A(n38456), .B(n5018), .Z(n4872) );
  AND U5524 ( .A(n4873), .B(n4872), .Z(n4940) );
  AND U5525 ( .A(b[31]), .B(a[15]), .Z(n4939) );
  XNOR U5526 ( .A(n4940), .B(n4939), .Z(n4941) );
  XNOR U5527 ( .A(n4942), .B(n4941), .Z(n4982) );
  NAND U5528 ( .A(n38185), .B(n4874), .Z(n4876) );
  XOR U5529 ( .A(b[23]), .B(a[25]), .Z(n5021) );
  NAND U5530 ( .A(n38132), .B(n5021), .Z(n4875) );
  AND U5531 ( .A(n4876), .B(n4875), .Z(n5011) );
  NAND U5532 ( .A(n184), .B(n4877), .Z(n4879) );
  XOR U5533 ( .A(b[7]), .B(a[41]), .Z(n5024) );
  NAND U5534 ( .A(n36592), .B(n5024), .Z(n4878) );
  AND U5535 ( .A(n4879), .B(n4878), .Z(n5010) );
  NAND U5536 ( .A(n38289), .B(n4880), .Z(n4882) );
  XOR U5537 ( .A(b[25]), .B(a[23]), .Z(n5027) );
  NAND U5538 ( .A(n38247), .B(n5027), .Z(n4881) );
  NAND U5539 ( .A(n4882), .B(n4881), .Z(n5009) );
  XOR U5540 ( .A(n5010), .B(n5009), .Z(n5012) );
  XOR U5541 ( .A(n5011), .B(n5012), .Z(n4981) );
  XOR U5542 ( .A(n4982), .B(n4981), .Z(n4984) );
  NAND U5543 ( .A(n187), .B(n4883), .Z(n4885) );
  XOR U5544 ( .A(b[13]), .B(a[35]), .Z(n5030) );
  NAND U5545 ( .A(n37295), .B(n5030), .Z(n4884) );
  AND U5546 ( .A(n4885), .B(n4884), .Z(n4976) );
  NAND U5547 ( .A(n186), .B(n4886), .Z(n4888) );
  XOR U5548 ( .A(b[11]), .B(a[37]), .Z(n5033) );
  NAND U5549 ( .A(n37097), .B(n5033), .Z(n4887) );
  NAND U5550 ( .A(n4888), .B(n4887), .Z(n4975) );
  XNOR U5551 ( .A(n4976), .B(n4975), .Z(n4978) );
  NAND U5552 ( .A(n188), .B(n4889), .Z(n4891) );
  XOR U5553 ( .A(b[15]), .B(a[33]), .Z(n5036) );
  NAND U5554 ( .A(n37382), .B(n5036), .Z(n4890) );
  AND U5555 ( .A(n4891), .B(n4890), .Z(n4972) );
  NAND U5556 ( .A(n38064), .B(n4892), .Z(n4894) );
  XOR U5557 ( .A(b[21]), .B(a[27]), .Z(n5039) );
  NAND U5558 ( .A(n37993), .B(n5039), .Z(n4893) );
  AND U5559 ( .A(n4894), .B(n4893), .Z(n4970) );
  NAND U5560 ( .A(n185), .B(n4895), .Z(n4897) );
  XOR U5561 ( .A(b[9]), .B(a[39]), .Z(n5042) );
  NAND U5562 ( .A(n36805), .B(n5042), .Z(n4896) );
  NAND U5563 ( .A(n4897), .B(n4896), .Z(n4969) );
  XNOR U5564 ( .A(n4970), .B(n4969), .Z(n4971) );
  XNOR U5565 ( .A(n4972), .B(n4971), .Z(n4977) );
  XOR U5566 ( .A(n4978), .B(n4977), .Z(n4983) );
  XNOR U5567 ( .A(n4984), .B(n4983), .Z(n4995) );
  XNOR U5568 ( .A(n4996), .B(n4995), .Z(n4927) );
  XNOR U5569 ( .A(n4928), .B(n4927), .Z(n4929) );
  XOR U5570 ( .A(n4930), .B(n4929), .Z(n5046) );
  XNOR U5571 ( .A(n5045), .B(n5046), .Z(n5047) );
  XNOR U5572 ( .A(n5048), .B(n5047), .Z(n4923) );
  XOR U5573 ( .A(n4924), .B(n4923), .Z(n4916) );
  NANDN U5574 ( .A(n4899), .B(n4898), .Z(n4903) );
  NANDN U5575 ( .A(n4901), .B(n4900), .Z(n4902) );
  AND U5576 ( .A(n4903), .B(n4902), .Z(n4915) );
  XOR U5577 ( .A(n4916), .B(n4915), .Z(n4918) );
  XNOR U5578 ( .A(n4917), .B(n4918), .Z(n4909) );
  XNOR U5579 ( .A(n4910), .B(n4909), .Z(n4911) );
  XNOR U5580 ( .A(n4912), .B(n4911), .Z(n5051) );
  XNOR U5581 ( .A(sreg[271]), .B(n5051), .Z(n5053) );
  NANDN U5582 ( .A(sreg[270]), .B(n4904), .Z(n4908) );
  NAND U5583 ( .A(n4906), .B(n4905), .Z(n4907) );
  NAND U5584 ( .A(n4908), .B(n4907), .Z(n5052) );
  XNOR U5585 ( .A(n5053), .B(n5052), .Z(c[271]) );
  NANDN U5586 ( .A(n4910), .B(n4909), .Z(n4914) );
  NANDN U5587 ( .A(n4912), .B(n4911), .Z(n4913) );
  AND U5588 ( .A(n4914), .B(n4913), .Z(n5059) );
  NANDN U5589 ( .A(n4916), .B(n4915), .Z(n4920) );
  NANDN U5590 ( .A(n4918), .B(n4917), .Z(n4919) );
  AND U5591 ( .A(n4920), .B(n4919), .Z(n5057) );
  NANDN U5592 ( .A(n4922), .B(n4921), .Z(n4926) );
  NAND U5593 ( .A(n4924), .B(n4923), .Z(n4925) );
  AND U5594 ( .A(n4926), .B(n4925), .Z(n5064) );
  NANDN U5595 ( .A(n4928), .B(n4927), .Z(n4932) );
  NANDN U5596 ( .A(n4930), .B(n4929), .Z(n4931) );
  AND U5597 ( .A(n4932), .B(n4931), .Z(n5193) );
  NANDN U5598 ( .A(n4934), .B(n4933), .Z(n4938) );
  NAND U5599 ( .A(n4936), .B(n4935), .Z(n4937) );
  AND U5600 ( .A(n4938), .B(n4937), .Z(n5192) );
  XNOR U5601 ( .A(n5193), .B(n5192), .Z(n5195) );
  NANDN U5602 ( .A(n4940), .B(n4939), .Z(n4944) );
  NANDN U5603 ( .A(n4942), .B(n4941), .Z(n4943) );
  AND U5604 ( .A(n4944), .B(n4943), .Z(n5128) );
  NAND U5605 ( .A(n38385), .B(n4945), .Z(n4947) );
  XOR U5606 ( .A(b[27]), .B(a[22]), .Z(n5074) );
  NAND U5607 ( .A(n38343), .B(n5074), .Z(n4946) );
  AND U5608 ( .A(n4947), .B(n4946), .Z(n5135) );
  NAND U5609 ( .A(n183), .B(n4948), .Z(n4950) );
  XOR U5610 ( .A(b[5]), .B(a[44]), .Z(n5077) );
  NAND U5611 ( .A(n36296), .B(n5077), .Z(n4949) );
  AND U5612 ( .A(n4950), .B(n4949), .Z(n5133) );
  NAND U5613 ( .A(n190), .B(n4951), .Z(n4953) );
  XOR U5614 ( .A(b[19]), .B(a[30]), .Z(n5080) );
  NAND U5615 ( .A(n37821), .B(n5080), .Z(n4952) );
  NAND U5616 ( .A(n4953), .B(n4952), .Z(n5132) );
  XNOR U5617 ( .A(n5133), .B(n5132), .Z(n5134) );
  XNOR U5618 ( .A(n5135), .B(n5134), .Z(n5126) );
  NAND U5619 ( .A(n38470), .B(n4954), .Z(n4956) );
  XOR U5620 ( .A(b[31]), .B(a[18]), .Z(n5083) );
  NAND U5621 ( .A(n38453), .B(n5083), .Z(n4955) );
  AND U5622 ( .A(n4956), .B(n4955), .Z(n5095) );
  NAND U5623 ( .A(n181), .B(n4957), .Z(n4959) );
  XOR U5624 ( .A(b[3]), .B(a[46]), .Z(n5086) );
  NAND U5625 ( .A(n182), .B(n5086), .Z(n4958) );
  AND U5626 ( .A(n4959), .B(n4958), .Z(n5093) );
  NAND U5627 ( .A(n189), .B(n4960), .Z(n4962) );
  XOR U5628 ( .A(b[17]), .B(a[32]), .Z(n5089) );
  NAND U5629 ( .A(n37652), .B(n5089), .Z(n4961) );
  NAND U5630 ( .A(n4962), .B(n4961), .Z(n5092) );
  XNOR U5631 ( .A(n5093), .B(n5092), .Z(n5094) );
  XOR U5632 ( .A(n5095), .B(n5094), .Z(n5127) );
  XOR U5633 ( .A(n5126), .B(n5127), .Z(n5129) );
  XOR U5634 ( .A(n5128), .B(n5129), .Z(n5175) );
  NANDN U5635 ( .A(n4964), .B(n4963), .Z(n4968) );
  NANDN U5636 ( .A(n4966), .B(n4965), .Z(n4967) );
  AND U5637 ( .A(n4968), .B(n4967), .Z(n5116) );
  NANDN U5638 ( .A(n4970), .B(n4969), .Z(n4974) );
  NANDN U5639 ( .A(n4972), .B(n4971), .Z(n4973) );
  NAND U5640 ( .A(n4974), .B(n4973), .Z(n5117) );
  XNOR U5641 ( .A(n5116), .B(n5117), .Z(n5118) );
  NANDN U5642 ( .A(n4976), .B(n4975), .Z(n4980) );
  NAND U5643 ( .A(n4978), .B(n4977), .Z(n4979) );
  NAND U5644 ( .A(n4980), .B(n4979), .Z(n5119) );
  XNOR U5645 ( .A(n5118), .B(n5119), .Z(n5174) );
  XNOR U5646 ( .A(n5175), .B(n5174), .Z(n5177) );
  NAND U5647 ( .A(n4982), .B(n4981), .Z(n4986) );
  NAND U5648 ( .A(n4984), .B(n4983), .Z(n4985) );
  AND U5649 ( .A(n4986), .B(n4985), .Z(n5176) );
  XOR U5650 ( .A(n5177), .B(n5176), .Z(n5189) );
  NANDN U5651 ( .A(n4988), .B(n4987), .Z(n4992) );
  NANDN U5652 ( .A(n4990), .B(n4989), .Z(n4991) );
  AND U5653 ( .A(n4992), .B(n4991), .Z(n5186) );
  NANDN U5654 ( .A(n4998), .B(n4997), .Z(n5002) );
  OR U5655 ( .A(n5000), .B(n4999), .Z(n5001) );
  AND U5656 ( .A(n5002), .B(n5001), .Z(n5181) );
  NANDN U5657 ( .A(n5004), .B(n5003), .Z(n5008) );
  NANDN U5658 ( .A(n5006), .B(n5005), .Z(n5007) );
  AND U5659 ( .A(n5008), .B(n5007), .Z(n5123) );
  NANDN U5660 ( .A(n5010), .B(n5009), .Z(n5014) );
  OR U5661 ( .A(n5012), .B(n5011), .Z(n5013) );
  NAND U5662 ( .A(n5014), .B(n5013), .Z(n5122) );
  XNOR U5663 ( .A(n5123), .B(n5122), .Z(n5125) );
  NAND U5664 ( .A(b[0]), .B(a[48]), .Z(n5015) );
  XNOR U5665 ( .A(b[1]), .B(n5015), .Z(n5017) );
  NANDN U5666 ( .A(b[0]), .B(a[47]), .Z(n5016) );
  NAND U5667 ( .A(n5017), .B(n5016), .Z(n5071) );
  NAND U5668 ( .A(n194), .B(n5018), .Z(n5020) );
  XOR U5669 ( .A(b[29]), .B(a[20]), .Z(n5144) );
  NAND U5670 ( .A(n38456), .B(n5144), .Z(n5019) );
  AND U5671 ( .A(n5020), .B(n5019), .Z(n5069) );
  AND U5672 ( .A(b[31]), .B(a[16]), .Z(n5068) );
  XNOR U5673 ( .A(n5069), .B(n5068), .Z(n5070) );
  XNOR U5674 ( .A(n5071), .B(n5070), .Z(n5111) );
  NAND U5675 ( .A(n38185), .B(n5021), .Z(n5023) );
  XOR U5676 ( .A(b[23]), .B(a[26]), .Z(n5150) );
  NAND U5677 ( .A(n38132), .B(n5150), .Z(n5022) );
  AND U5678 ( .A(n5023), .B(n5022), .Z(n5140) );
  NAND U5679 ( .A(n184), .B(n5024), .Z(n5026) );
  XOR U5680 ( .A(b[7]), .B(a[42]), .Z(n5153) );
  NAND U5681 ( .A(n36592), .B(n5153), .Z(n5025) );
  AND U5682 ( .A(n5026), .B(n5025), .Z(n5139) );
  NAND U5683 ( .A(n38289), .B(n5027), .Z(n5029) );
  XOR U5684 ( .A(b[25]), .B(a[24]), .Z(n5156) );
  NAND U5685 ( .A(n38247), .B(n5156), .Z(n5028) );
  NAND U5686 ( .A(n5029), .B(n5028), .Z(n5138) );
  XOR U5687 ( .A(n5139), .B(n5138), .Z(n5141) );
  XOR U5688 ( .A(n5140), .B(n5141), .Z(n5110) );
  XOR U5689 ( .A(n5111), .B(n5110), .Z(n5113) );
  NAND U5690 ( .A(n187), .B(n5030), .Z(n5032) );
  XOR U5691 ( .A(b[13]), .B(a[36]), .Z(n5159) );
  NAND U5692 ( .A(n37295), .B(n5159), .Z(n5031) );
  AND U5693 ( .A(n5032), .B(n5031), .Z(n5105) );
  NAND U5694 ( .A(n186), .B(n5033), .Z(n5035) );
  XOR U5695 ( .A(b[11]), .B(a[38]), .Z(n5162) );
  NAND U5696 ( .A(n37097), .B(n5162), .Z(n5034) );
  NAND U5697 ( .A(n5035), .B(n5034), .Z(n5104) );
  XNOR U5698 ( .A(n5105), .B(n5104), .Z(n5107) );
  NAND U5699 ( .A(n188), .B(n5036), .Z(n5038) );
  XOR U5700 ( .A(b[15]), .B(a[34]), .Z(n5165) );
  NAND U5701 ( .A(n37382), .B(n5165), .Z(n5037) );
  AND U5702 ( .A(n5038), .B(n5037), .Z(n5101) );
  NAND U5703 ( .A(n38064), .B(n5039), .Z(n5041) );
  XOR U5704 ( .A(b[21]), .B(a[28]), .Z(n5168) );
  NAND U5705 ( .A(n37993), .B(n5168), .Z(n5040) );
  AND U5706 ( .A(n5041), .B(n5040), .Z(n5099) );
  NAND U5707 ( .A(n185), .B(n5042), .Z(n5044) );
  XOR U5708 ( .A(b[9]), .B(a[40]), .Z(n5171) );
  NAND U5709 ( .A(n36805), .B(n5171), .Z(n5043) );
  NAND U5710 ( .A(n5044), .B(n5043), .Z(n5098) );
  XNOR U5711 ( .A(n5099), .B(n5098), .Z(n5100) );
  XNOR U5712 ( .A(n5101), .B(n5100), .Z(n5106) );
  XOR U5713 ( .A(n5107), .B(n5106), .Z(n5112) );
  XNOR U5714 ( .A(n5113), .B(n5112), .Z(n5124) );
  XNOR U5715 ( .A(n5125), .B(n5124), .Z(n5180) );
  XNOR U5716 ( .A(n5181), .B(n5180), .Z(n5182) );
  XOR U5717 ( .A(n5183), .B(n5182), .Z(n5187) );
  XNOR U5718 ( .A(n5186), .B(n5187), .Z(n5188) );
  XNOR U5719 ( .A(n5189), .B(n5188), .Z(n5194) );
  XOR U5720 ( .A(n5195), .B(n5194), .Z(n5063) );
  NANDN U5721 ( .A(n5046), .B(n5045), .Z(n5050) );
  NANDN U5722 ( .A(n5048), .B(n5047), .Z(n5049) );
  AND U5723 ( .A(n5050), .B(n5049), .Z(n5062) );
  XOR U5724 ( .A(n5063), .B(n5062), .Z(n5065) );
  XNOR U5725 ( .A(n5064), .B(n5065), .Z(n5056) );
  XNOR U5726 ( .A(n5057), .B(n5056), .Z(n5058) );
  XNOR U5727 ( .A(n5059), .B(n5058), .Z(n5198) );
  XNOR U5728 ( .A(sreg[272]), .B(n5198), .Z(n5200) );
  NANDN U5729 ( .A(sreg[271]), .B(n5051), .Z(n5055) );
  NAND U5730 ( .A(n5053), .B(n5052), .Z(n5054) );
  NAND U5731 ( .A(n5055), .B(n5054), .Z(n5199) );
  XNOR U5732 ( .A(n5200), .B(n5199), .Z(c[272]) );
  NANDN U5733 ( .A(n5057), .B(n5056), .Z(n5061) );
  NANDN U5734 ( .A(n5059), .B(n5058), .Z(n5060) );
  AND U5735 ( .A(n5061), .B(n5060), .Z(n5206) );
  NANDN U5736 ( .A(n5063), .B(n5062), .Z(n5067) );
  NANDN U5737 ( .A(n5065), .B(n5064), .Z(n5066) );
  AND U5738 ( .A(n5067), .B(n5066), .Z(n5204) );
  NANDN U5739 ( .A(n5069), .B(n5068), .Z(n5073) );
  NANDN U5740 ( .A(n5071), .B(n5070), .Z(n5072) );
  AND U5741 ( .A(n5073), .B(n5072), .Z(n5283) );
  NAND U5742 ( .A(n38385), .B(n5074), .Z(n5076) );
  XOR U5743 ( .A(b[27]), .B(a[23]), .Z(n5227) );
  NAND U5744 ( .A(n38343), .B(n5227), .Z(n5075) );
  AND U5745 ( .A(n5076), .B(n5075), .Z(n5290) );
  NAND U5746 ( .A(n183), .B(n5077), .Z(n5079) );
  XOR U5747 ( .A(b[5]), .B(a[45]), .Z(n5230) );
  NAND U5748 ( .A(n36296), .B(n5230), .Z(n5078) );
  AND U5749 ( .A(n5079), .B(n5078), .Z(n5288) );
  NAND U5750 ( .A(n190), .B(n5080), .Z(n5082) );
  XOR U5751 ( .A(b[19]), .B(a[31]), .Z(n5233) );
  NAND U5752 ( .A(n37821), .B(n5233), .Z(n5081) );
  NAND U5753 ( .A(n5082), .B(n5081), .Z(n5287) );
  XNOR U5754 ( .A(n5288), .B(n5287), .Z(n5289) );
  XNOR U5755 ( .A(n5290), .B(n5289), .Z(n5281) );
  NAND U5756 ( .A(n38470), .B(n5083), .Z(n5085) );
  XOR U5757 ( .A(b[31]), .B(a[19]), .Z(n5236) );
  NAND U5758 ( .A(n38453), .B(n5236), .Z(n5084) );
  AND U5759 ( .A(n5085), .B(n5084), .Z(n5248) );
  NAND U5760 ( .A(n181), .B(n5086), .Z(n5088) );
  XOR U5761 ( .A(b[3]), .B(a[47]), .Z(n5239) );
  NAND U5762 ( .A(n182), .B(n5239), .Z(n5087) );
  AND U5763 ( .A(n5088), .B(n5087), .Z(n5246) );
  NAND U5764 ( .A(n189), .B(n5089), .Z(n5091) );
  XOR U5765 ( .A(b[17]), .B(a[33]), .Z(n5242) );
  NAND U5766 ( .A(n37652), .B(n5242), .Z(n5090) );
  NAND U5767 ( .A(n5091), .B(n5090), .Z(n5245) );
  XNOR U5768 ( .A(n5246), .B(n5245), .Z(n5247) );
  XOR U5769 ( .A(n5248), .B(n5247), .Z(n5282) );
  XOR U5770 ( .A(n5281), .B(n5282), .Z(n5284) );
  XOR U5771 ( .A(n5283), .B(n5284), .Z(n5330) );
  NANDN U5772 ( .A(n5093), .B(n5092), .Z(n5097) );
  NANDN U5773 ( .A(n5095), .B(n5094), .Z(n5096) );
  AND U5774 ( .A(n5097), .B(n5096), .Z(n5269) );
  NANDN U5775 ( .A(n5099), .B(n5098), .Z(n5103) );
  NANDN U5776 ( .A(n5101), .B(n5100), .Z(n5102) );
  NAND U5777 ( .A(n5103), .B(n5102), .Z(n5270) );
  XNOR U5778 ( .A(n5269), .B(n5270), .Z(n5271) );
  NANDN U5779 ( .A(n5105), .B(n5104), .Z(n5109) );
  NAND U5780 ( .A(n5107), .B(n5106), .Z(n5108) );
  NAND U5781 ( .A(n5109), .B(n5108), .Z(n5272) );
  XNOR U5782 ( .A(n5271), .B(n5272), .Z(n5329) );
  XNOR U5783 ( .A(n5330), .B(n5329), .Z(n5332) );
  NAND U5784 ( .A(n5111), .B(n5110), .Z(n5115) );
  NAND U5785 ( .A(n5113), .B(n5112), .Z(n5114) );
  AND U5786 ( .A(n5115), .B(n5114), .Z(n5331) );
  XOR U5787 ( .A(n5332), .B(n5331), .Z(n5343) );
  NANDN U5788 ( .A(n5117), .B(n5116), .Z(n5121) );
  NANDN U5789 ( .A(n5119), .B(n5118), .Z(n5120) );
  AND U5790 ( .A(n5121), .B(n5120), .Z(n5341) );
  NANDN U5791 ( .A(n5127), .B(n5126), .Z(n5131) );
  OR U5792 ( .A(n5129), .B(n5128), .Z(n5130) );
  AND U5793 ( .A(n5131), .B(n5130), .Z(n5336) );
  NANDN U5794 ( .A(n5133), .B(n5132), .Z(n5137) );
  NANDN U5795 ( .A(n5135), .B(n5134), .Z(n5136) );
  AND U5796 ( .A(n5137), .B(n5136), .Z(n5276) );
  NANDN U5797 ( .A(n5139), .B(n5138), .Z(n5143) );
  OR U5798 ( .A(n5141), .B(n5140), .Z(n5142) );
  NAND U5799 ( .A(n5143), .B(n5142), .Z(n5275) );
  XNOR U5800 ( .A(n5276), .B(n5275), .Z(n5277) );
  NAND U5801 ( .A(n194), .B(n5144), .Z(n5146) );
  XOR U5802 ( .A(b[29]), .B(a[21]), .Z(n5302) );
  NAND U5803 ( .A(n38456), .B(n5302), .Z(n5145) );
  AND U5804 ( .A(n5146), .B(n5145), .Z(n5222) );
  AND U5805 ( .A(b[31]), .B(a[17]), .Z(n5221) );
  XNOR U5806 ( .A(n5222), .B(n5221), .Z(n5223) );
  NAND U5807 ( .A(b[0]), .B(a[49]), .Z(n5147) );
  XNOR U5808 ( .A(b[1]), .B(n5147), .Z(n5149) );
  NANDN U5809 ( .A(b[0]), .B(a[48]), .Z(n5148) );
  NAND U5810 ( .A(n5149), .B(n5148), .Z(n5224) );
  XNOR U5811 ( .A(n5223), .B(n5224), .Z(n5263) );
  NAND U5812 ( .A(n38185), .B(n5150), .Z(n5152) );
  XOR U5813 ( .A(b[23]), .B(a[27]), .Z(n5305) );
  NAND U5814 ( .A(n38132), .B(n5305), .Z(n5151) );
  AND U5815 ( .A(n5152), .B(n5151), .Z(n5296) );
  NAND U5816 ( .A(n184), .B(n5153), .Z(n5155) );
  XOR U5817 ( .A(b[7]), .B(a[43]), .Z(n5308) );
  NAND U5818 ( .A(n36592), .B(n5308), .Z(n5154) );
  AND U5819 ( .A(n5155), .B(n5154), .Z(n5294) );
  NAND U5820 ( .A(n38289), .B(n5156), .Z(n5158) );
  XOR U5821 ( .A(b[25]), .B(a[25]), .Z(n5311) );
  NAND U5822 ( .A(n38247), .B(n5311), .Z(n5157) );
  NAND U5823 ( .A(n5158), .B(n5157), .Z(n5293) );
  XNOR U5824 ( .A(n5294), .B(n5293), .Z(n5295) );
  XOR U5825 ( .A(n5296), .B(n5295), .Z(n5264) );
  XNOR U5826 ( .A(n5263), .B(n5264), .Z(n5265) );
  NAND U5827 ( .A(n187), .B(n5159), .Z(n5161) );
  XOR U5828 ( .A(b[13]), .B(a[37]), .Z(n5314) );
  NAND U5829 ( .A(n37295), .B(n5314), .Z(n5160) );
  AND U5830 ( .A(n5161), .B(n5160), .Z(n5258) );
  NAND U5831 ( .A(n186), .B(n5162), .Z(n5164) );
  XOR U5832 ( .A(b[11]), .B(a[39]), .Z(n5317) );
  NAND U5833 ( .A(n37097), .B(n5317), .Z(n5163) );
  NAND U5834 ( .A(n5164), .B(n5163), .Z(n5257) );
  XNOR U5835 ( .A(n5258), .B(n5257), .Z(n5259) );
  NAND U5836 ( .A(n188), .B(n5165), .Z(n5167) );
  XOR U5837 ( .A(b[15]), .B(a[35]), .Z(n5320) );
  NAND U5838 ( .A(n37382), .B(n5320), .Z(n5166) );
  AND U5839 ( .A(n5167), .B(n5166), .Z(n5254) );
  NAND U5840 ( .A(n38064), .B(n5168), .Z(n5170) );
  XOR U5841 ( .A(b[21]), .B(a[29]), .Z(n5323) );
  NAND U5842 ( .A(n37993), .B(n5323), .Z(n5169) );
  AND U5843 ( .A(n5170), .B(n5169), .Z(n5252) );
  NAND U5844 ( .A(n185), .B(n5171), .Z(n5173) );
  XOR U5845 ( .A(b[9]), .B(a[41]), .Z(n5326) );
  NAND U5846 ( .A(n36805), .B(n5326), .Z(n5172) );
  NAND U5847 ( .A(n5173), .B(n5172), .Z(n5251) );
  XNOR U5848 ( .A(n5252), .B(n5251), .Z(n5253) );
  XOR U5849 ( .A(n5254), .B(n5253), .Z(n5260) );
  XOR U5850 ( .A(n5259), .B(n5260), .Z(n5266) );
  XOR U5851 ( .A(n5265), .B(n5266), .Z(n5278) );
  XNOR U5852 ( .A(n5277), .B(n5278), .Z(n5335) );
  XNOR U5853 ( .A(n5336), .B(n5335), .Z(n5337) );
  XOR U5854 ( .A(n5338), .B(n5337), .Z(n5342) );
  XOR U5855 ( .A(n5341), .B(n5342), .Z(n5344) );
  XOR U5856 ( .A(n5343), .B(n5344), .Z(n5218) );
  NANDN U5857 ( .A(n5175), .B(n5174), .Z(n5179) );
  NAND U5858 ( .A(n5177), .B(n5176), .Z(n5178) );
  AND U5859 ( .A(n5179), .B(n5178), .Z(n5216) );
  NANDN U5860 ( .A(n5181), .B(n5180), .Z(n5185) );
  NANDN U5861 ( .A(n5183), .B(n5182), .Z(n5184) );
  AND U5862 ( .A(n5185), .B(n5184), .Z(n5215) );
  XNOR U5863 ( .A(n5216), .B(n5215), .Z(n5217) );
  XNOR U5864 ( .A(n5218), .B(n5217), .Z(n5209) );
  NANDN U5865 ( .A(n5187), .B(n5186), .Z(n5191) );
  NANDN U5866 ( .A(n5189), .B(n5188), .Z(n5190) );
  NAND U5867 ( .A(n5191), .B(n5190), .Z(n5210) );
  XNOR U5868 ( .A(n5209), .B(n5210), .Z(n5211) );
  NANDN U5869 ( .A(n5193), .B(n5192), .Z(n5197) );
  NAND U5870 ( .A(n5195), .B(n5194), .Z(n5196) );
  NAND U5871 ( .A(n5197), .B(n5196), .Z(n5212) );
  XNOR U5872 ( .A(n5211), .B(n5212), .Z(n5203) );
  XNOR U5873 ( .A(n5204), .B(n5203), .Z(n5205) );
  XNOR U5874 ( .A(n5206), .B(n5205), .Z(n5347) );
  XNOR U5875 ( .A(sreg[273]), .B(n5347), .Z(n5349) );
  NANDN U5876 ( .A(sreg[272]), .B(n5198), .Z(n5202) );
  NAND U5877 ( .A(n5200), .B(n5199), .Z(n5201) );
  NAND U5878 ( .A(n5202), .B(n5201), .Z(n5348) );
  XNOR U5879 ( .A(n5349), .B(n5348), .Z(c[273]) );
  NANDN U5880 ( .A(n5204), .B(n5203), .Z(n5208) );
  NANDN U5881 ( .A(n5206), .B(n5205), .Z(n5207) );
  AND U5882 ( .A(n5208), .B(n5207), .Z(n5355) );
  NANDN U5883 ( .A(n5210), .B(n5209), .Z(n5214) );
  NANDN U5884 ( .A(n5212), .B(n5211), .Z(n5213) );
  AND U5885 ( .A(n5214), .B(n5213), .Z(n5353) );
  NANDN U5886 ( .A(n5216), .B(n5215), .Z(n5220) );
  NANDN U5887 ( .A(n5218), .B(n5217), .Z(n5219) );
  AND U5888 ( .A(n5220), .B(n5219), .Z(n5361) );
  NANDN U5889 ( .A(n5222), .B(n5221), .Z(n5226) );
  NANDN U5890 ( .A(n5224), .B(n5223), .Z(n5225) );
  AND U5891 ( .A(n5226), .B(n5225), .Z(n5444) );
  NAND U5892 ( .A(n38385), .B(n5227), .Z(n5229) );
  XOR U5893 ( .A(b[27]), .B(a[24]), .Z(n5388) );
  NAND U5894 ( .A(n38343), .B(n5388), .Z(n5228) );
  AND U5895 ( .A(n5229), .B(n5228), .Z(n5451) );
  NAND U5896 ( .A(n183), .B(n5230), .Z(n5232) );
  XOR U5897 ( .A(b[5]), .B(a[46]), .Z(n5391) );
  NAND U5898 ( .A(n36296), .B(n5391), .Z(n5231) );
  AND U5899 ( .A(n5232), .B(n5231), .Z(n5449) );
  NAND U5900 ( .A(n190), .B(n5233), .Z(n5235) );
  XOR U5901 ( .A(b[19]), .B(a[32]), .Z(n5394) );
  NAND U5902 ( .A(n37821), .B(n5394), .Z(n5234) );
  NAND U5903 ( .A(n5235), .B(n5234), .Z(n5448) );
  XNOR U5904 ( .A(n5449), .B(n5448), .Z(n5450) );
  XNOR U5905 ( .A(n5451), .B(n5450), .Z(n5442) );
  NAND U5906 ( .A(n38470), .B(n5236), .Z(n5238) );
  XOR U5907 ( .A(b[31]), .B(a[20]), .Z(n5397) );
  NAND U5908 ( .A(n38453), .B(n5397), .Z(n5237) );
  AND U5909 ( .A(n5238), .B(n5237), .Z(n5409) );
  NAND U5910 ( .A(n181), .B(n5239), .Z(n5241) );
  XOR U5911 ( .A(b[3]), .B(a[48]), .Z(n5400) );
  NAND U5912 ( .A(n182), .B(n5400), .Z(n5240) );
  AND U5913 ( .A(n5241), .B(n5240), .Z(n5407) );
  NAND U5914 ( .A(n189), .B(n5242), .Z(n5244) );
  XOR U5915 ( .A(b[17]), .B(a[34]), .Z(n5403) );
  NAND U5916 ( .A(n37652), .B(n5403), .Z(n5243) );
  NAND U5917 ( .A(n5244), .B(n5243), .Z(n5406) );
  XNOR U5918 ( .A(n5407), .B(n5406), .Z(n5408) );
  XOR U5919 ( .A(n5409), .B(n5408), .Z(n5443) );
  XOR U5920 ( .A(n5442), .B(n5443), .Z(n5445) );
  XOR U5921 ( .A(n5444), .B(n5445), .Z(n5377) );
  NANDN U5922 ( .A(n5246), .B(n5245), .Z(n5250) );
  NANDN U5923 ( .A(n5248), .B(n5247), .Z(n5249) );
  AND U5924 ( .A(n5250), .B(n5249), .Z(n5430) );
  NANDN U5925 ( .A(n5252), .B(n5251), .Z(n5256) );
  NANDN U5926 ( .A(n5254), .B(n5253), .Z(n5255) );
  NAND U5927 ( .A(n5256), .B(n5255), .Z(n5431) );
  XNOR U5928 ( .A(n5430), .B(n5431), .Z(n5432) );
  NANDN U5929 ( .A(n5258), .B(n5257), .Z(n5262) );
  NANDN U5930 ( .A(n5260), .B(n5259), .Z(n5261) );
  NAND U5931 ( .A(n5262), .B(n5261), .Z(n5433) );
  XNOR U5932 ( .A(n5432), .B(n5433), .Z(n5376) );
  XNOR U5933 ( .A(n5377), .B(n5376), .Z(n5379) );
  NANDN U5934 ( .A(n5264), .B(n5263), .Z(n5268) );
  NANDN U5935 ( .A(n5266), .B(n5265), .Z(n5267) );
  AND U5936 ( .A(n5268), .B(n5267), .Z(n5378) );
  XOR U5937 ( .A(n5379), .B(n5378), .Z(n5492) );
  NANDN U5938 ( .A(n5270), .B(n5269), .Z(n5274) );
  NANDN U5939 ( .A(n5272), .B(n5271), .Z(n5273) );
  AND U5940 ( .A(n5274), .B(n5273), .Z(n5490) );
  NANDN U5941 ( .A(n5276), .B(n5275), .Z(n5280) );
  NANDN U5942 ( .A(n5278), .B(n5277), .Z(n5279) );
  AND U5943 ( .A(n5280), .B(n5279), .Z(n5373) );
  NANDN U5944 ( .A(n5282), .B(n5281), .Z(n5286) );
  OR U5945 ( .A(n5284), .B(n5283), .Z(n5285) );
  AND U5946 ( .A(n5286), .B(n5285), .Z(n5371) );
  NANDN U5947 ( .A(n5288), .B(n5287), .Z(n5292) );
  NANDN U5948 ( .A(n5290), .B(n5289), .Z(n5291) );
  AND U5949 ( .A(n5292), .B(n5291), .Z(n5437) );
  NANDN U5950 ( .A(n5294), .B(n5293), .Z(n5298) );
  NANDN U5951 ( .A(n5296), .B(n5295), .Z(n5297) );
  NAND U5952 ( .A(n5298), .B(n5297), .Z(n5436) );
  XNOR U5953 ( .A(n5437), .B(n5436), .Z(n5438) );
  NAND U5954 ( .A(b[0]), .B(a[50]), .Z(n5299) );
  XNOR U5955 ( .A(b[1]), .B(n5299), .Z(n5301) );
  NANDN U5956 ( .A(b[0]), .B(a[49]), .Z(n5300) );
  NAND U5957 ( .A(n5301), .B(n5300), .Z(n5385) );
  NAND U5958 ( .A(n194), .B(n5302), .Z(n5304) );
  XOR U5959 ( .A(b[29]), .B(a[22]), .Z(n5460) );
  NAND U5960 ( .A(n38456), .B(n5460), .Z(n5303) );
  AND U5961 ( .A(n5304), .B(n5303), .Z(n5383) );
  AND U5962 ( .A(b[31]), .B(a[18]), .Z(n5382) );
  XNOR U5963 ( .A(n5383), .B(n5382), .Z(n5384) );
  XNOR U5964 ( .A(n5385), .B(n5384), .Z(n5424) );
  NAND U5965 ( .A(n38185), .B(n5305), .Z(n5307) );
  XOR U5966 ( .A(b[23]), .B(a[28]), .Z(n5466) );
  NAND U5967 ( .A(n38132), .B(n5466), .Z(n5306) );
  AND U5968 ( .A(n5307), .B(n5306), .Z(n5457) );
  NAND U5969 ( .A(n184), .B(n5308), .Z(n5310) );
  XOR U5970 ( .A(b[7]), .B(a[44]), .Z(n5469) );
  NAND U5971 ( .A(n36592), .B(n5469), .Z(n5309) );
  AND U5972 ( .A(n5310), .B(n5309), .Z(n5455) );
  NAND U5973 ( .A(n38289), .B(n5311), .Z(n5313) );
  XOR U5974 ( .A(b[25]), .B(a[26]), .Z(n5472) );
  NAND U5975 ( .A(n38247), .B(n5472), .Z(n5312) );
  NAND U5976 ( .A(n5313), .B(n5312), .Z(n5454) );
  XNOR U5977 ( .A(n5455), .B(n5454), .Z(n5456) );
  XOR U5978 ( .A(n5457), .B(n5456), .Z(n5425) );
  XNOR U5979 ( .A(n5424), .B(n5425), .Z(n5426) );
  NAND U5980 ( .A(n187), .B(n5314), .Z(n5316) );
  XOR U5981 ( .A(b[13]), .B(a[38]), .Z(n5475) );
  NAND U5982 ( .A(n37295), .B(n5475), .Z(n5315) );
  AND U5983 ( .A(n5316), .B(n5315), .Z(n5419) );
  NAND U5984 ( .A(n186), .B(n5317), .Z(n5319) );
  XOR U5985 ( .A(b[11]), .B(a[40]), .Z(n5478) );
  NAND U5986 ( .A(n37097), .B(n5478), .Z(n5318) );
  NAND U5987 ( .A(n5319), .B(n5318), .Z(n5418) );
  XNOR U5988 ( .A(n5419), .B(n5418), .Z(n5420) );
  NAND U5989 ( .A(n188), .B(n5320), .Z(n5322) );
  XOR U5990 ( .A(b[15]), .B(a[36]), .Z(n5481) );
  NAND U5991 ( .A(n37382), .B(n5481), .Z(n5321) );
  AND U5992 ( .A(n5322), .B(n5321), .Z(n5415) );
  NAND U5993 ( .A(n38064), .B(n5323), .Z(n5325) );
  XOR U5994 ( .A(b[21]), .B(a[30]), .Z(n5484) );
  NAND U5995 ( .A(n37993), .B(n5484), .Z(n5324) );
  AND U5996 ( .A(n5325), .B(n5324), .Z(n5413) );
  NAND U5997 ( .A(n185), .B(n5326), .Z(n5328) );
  XOR U5998 ( .A(b[9]), .B(a[42]), .Z(n5487) );
  NAND U5999 ( .A(n36805), .B(n5487), .Z(n5327) );
  NAND U6000 ( .A(n5328), .B(n5327), .Z(n5412) );
  XNOR U6001 ( .A(n5413), .B(n5412), .Z(n5414) );
  XOR U6002 ( .A(n5415), .B(n5414), .Z(n5421) );
  XOR U6003 ( .A(n5420), .B(n5421), .Z(n5427) );
  XOR U6004 ( .A(n5426), .B(n5427), .Z(n5439) );
  XNOR U6005 ( .A(n5438), .B(n5439), .Z(n5370) );
  XNOR U6006 ( .A(n5371), .B(n5370), .Z(n5372) );
  XOR U6007 ( .A(n5373), .B(n5372), .Z(n5491) );
  XOR U6008 ( .A(n5490), .B(n5491), .Z(n5493) );
  XOR U6009 ( .A(n5492), .B(n5493), .Z(n5367) );
  NANDN U6010 ( .A(n5330), .B(n5329), .Z(n5334) );
  NAND U6011 ( .A(n5332), .B(n5331), .Z(n5333) );
  AND U6012 ( .A(n5334), .B(n5333), .Z(n5365) );
  NANDN U6013 ( .A(n5336), .B(n5335), .Z(n5340) );
  NANDN U6014 ( .A(n5338), .B(n5337), .Z(n5339) );
  AND U6015 ( .A(n5340), .B(n5339), .Z(n5364) );
  XNOR U6016 ( .A(n5365), .B(n5364), .Z(n5366) );
  XNOR U6017 ( .A(n5367), .B(n5366), .Z(n5358) );
  NANDN U6018 ( .A(n5342), .B(n5341), .Z(n5346) );
  OR U6019 ( .A(n5344), .B(n5343), .Z(n5345) );
  NAND U6020 ( .A(n5346), .B(n5345), .Z(n5359) );
  XNOR U6021 ( .A(n5358), .B(n5359), .Z(n5360) );
  XNOR U6022 ( .A(n5361), .B(n5360), .Z(n5352) );
  XNOR U6023 ( .A(n5353), .B(n5352), .Z(n5354) );
  XNOR U6024 ( .A(n5355), .B(n5354), .Z(n5496) );
  XNOR U6025 ( .A(sreg[274]), .B(n5496), .Z(n5498) );
  NANDN U6026 ( .A(sreg[273]), .B(n5347), .Z(n5351) );
  NAND U6027 ( .A(n5349), .B(n5348), .Z(n5350) );
  NAND U6028 ( .A(n5351), .B(n5350), .Z(n5497) );
  XNOR U6029 ( .A(n5498), .B(n5497), .Z(c[274]) );
  NANDN U6030 ( .A(n5353), .B(n5352), .Z(n5357) );
  NANDN U6031 ( .A(n5355), .B(n5354), .Z(n5356) );
  AND U6032 ( .A(n5357), .B(n5356), .Z(n5504) );
  NANDN U6033 ( .A(n5359), .B(n5358), .Z(n5363) );
  NANDN U6034 ( .A(n5361), .B(n5360), .Z(n5362) );
  AND U6035 ( .A(n5363), .B(n5362), .Z(n5502) );
  NANDN U6036 ( .A(n5365), .B(n5364), .Z(n5369) );
  NANDN U6037 ( .A(n5367), .B(n5366), .Z(n5368) );
  AND U6038 ( .A(n5369), .B(n5368), .Z(n5510) );
  NANDN U6039 ( .A(n5371), .B(n5370), .Z(n5375) );
  NANDN U6040 ( .A(n5373), .B(n5372), .Z(n5374) );
  AND U6041 ( .A(n5375), .B(n5374), .Z(n5514) );
  NANDN U6042 ( .A(n5377), .B(n5376), .Z(n5381) );
  NAND U6043 ( .A(n5379), .B(n5378), .Z(n5380) );
  AND U6044 ( .A(n5381), .B(n5380), .Z(n5513) );
  XNOR U6045 ( .A(n5514), .B(n5513), .Z(n5516) );
  NANDN U6046 ( .A(n5383), .B(n5382), .Z(n5387) );
  NANDN U6047 ( .A(n5385), .B(n5384), .Z(n5386) );
  AND U6048 ( .A(n5387), .B(n5386), .Z(n5591) );
  NAND U6049 ( .A(n38385), .B(n5388), .Z(n5390) );
  XOR U6050 ( .A(b[27]), .B(a[25]), .Z(n5537) );
  NAND U6051 ( .A(n38343), .B(n5537), .Z(n5389) );
  AND U6052 ( .A(n5390), .B(n5389), .Z(n5598) );
  NAND U6053 ( .A(n183), .B(n5391), .Z(n5393) );
  XOR U6054 ( .A(b[5]), .B(a[47]), .Z(n5540) );
  NAND U6055 ( .A(n36296), .B(n5540), .Z(n5392) );
  AND U6056 ( .A(n5393), .B(n5392), .Z(n5596) );
  NAND U6057 ( .A(n190), .B(n5394), .Z(n5396) );
  XOR U6058 ( .A(b[19]), .B(a[33]), .Z(n5543) );
  NAND U6059 ( .A(n37821), .B(n5543), .Z(n5395) );
  NAND U6060 ( .A(n5396), .B(n5395), .Z(n5595) );
  XNOR U6061 ( .A(n5596), .B(n5595), .Z(n5597) );
  XNOR U6062 ( .A(n5598), .B(n5597), .Z(n5589) );
  NAND U6063 ( .A(n38470), .B(n5397), .Z(n5399) );
  XOR U6064 ( .A(b[31]), .B(a[21]), .Z(n5546) );
  NAND U6065 ( .A(n38453), .B(n5546), .Z(n5398) );
  AND U6066 ( .A(n5399), .B(n5398), .Z(n5558) );
  NAND U6067 ( .A(n181), .B(n5400), .Z(n5402) );
  XOR U6068 ( .A(b[3]), .B(a[49]), .Z(n5549) );
  NAND U6069 ( .A(n182), .B(n5549), .Z(n5401) );
  AND U6070 ( .A(n5402), .B(n5401), .Z(n5556) );
  NAND U6071 ( .A(n189), .B(n5403), .Z(n5405) );
  XOR U6072 ( .A(b[17]), .B(a[35]), .Z(n5552) );
  NAND U6073 ( .A(n37652), .B(n5552), .Z(n5404) );
  NAND U6074 ( .A(n5405), .B(n5404), .Z(n5555) );
  XNOR U6075 ( .A(n5556), .B(n5555), .Z(n5557) );
  XOR U6076 ( .A(n5558), .B(n5557), .Z(n5590) );
  XOR U6077 ( .A(n5589), .B(n5590), .Z(n5592) );
  XOR U6078 ( .A(n5591), .B(n5592), .Z(n5526) );
  NANDN U6079 ( .A(n5407), .B(n5406), .Z(n5411) );
  NANDN U6080 ( .A(n5409), .B(n5408), .Z(n5410) );
  AND U6081 ( .A(n5411), .B(n5410), .Z(n5579) );
  NANDN U6082 ( .A(n5413), .B(n5412), .Z(n5417) );
  NANDN U6083 ( .A(n5415), .B(n5414), .Z(n5416) );
  NAND U6084 ( .A(n5417), .B(n5416), .Z(n5580) );
  XNOR U6085 ( .A(n5579), .B(n5580), .Z(n5581) );
  NANDN U6086 ( .A(n5419), .B(n5418), .Z(n5423) );
  NANDN U6087 ( .A(n5421), .B(n5420), .Z(n5422) );
  NAND U6088 ( .A(n5423), .B(n5422), .Z(n5582) );
  XNOR U6089 ( .A(n5581), .B(n5582), .Z(n5525) );
  XNOR U6090 ( .A(n5526), .B(n5525), .Z(n5528) );
  NANDN U6091 ( .A(n5425), .B(n5424), .Z(n5429) );
  NANDN U6092 ( .A(n5427), .B(n5426), .Z(n5428) );
  AND U6093 ( .A(n5429), .B(n5428), .Z(n5527) );
  XOR U6094 ( .A(n5528), .B(n5527), .Z(n5640) );
  NANDN U6095 ( .A(n5431), .B(n5430), .Z(n5435) );
  NANDN U6096 ( .A(n5433), .B(n5432), .Z(n5434) );
  AND U6097 ( .A(n5435), .B(n5434), .Z(n5637) );
  NANDN U6098 ( .A(n5437), .B(n5436), .Z(n5441) );
  NANDN U6099 ( .A(n5439), .B(n5438), .Z(n5440) );
  AND U6100 ( .A(n5441), .B(n5440), .Z(n5522) );
  NANDN U6101 ( .A(n5443), .B(n5442), .Z(n5447) );
  OR U6102 ( .A(n5445), .B(n5444), .Z(n5446) );
  AND U6103 ( .A(n5447), .B(n5446), .Z(n5520) );
  NANDN U6104 ( .A(n5449), .B(n5448), .Z(n5453) );
  NANDN U6105 ( .A(n5451), .B(n5450), .Z(n5452) );
  AND U6106 ( .A(n5453), .B(n5452), .Z(n5586) );
  NANDN U6107 ( .A(n5455), .B(n5454), .Z(n5459) );
  NANDN U6108 ( .A(n5457), .B(n5456), .Z(n5458) );
  NAND U6109 ( .A(n5459), .B(n5458), .Z(n5585) );
  XNOR U6110 ( .A(n5586), .B(n5585), .Z(n5588) );
  NAND U6111 ( .A(n194), .B(n5460), .Z(n5462) );
  XOR U6112 ( .A(b[29]), .B(a[23]), .Z(n5607) );
  NAND U6113 ( .A(n38456), .B(n5607), .Z(n5461) );
  AND U6114 ( .A(n5462), .B(n5461), .Z(n5532) );
  AND U6115 ( .A(b[31]), .B(a[19]), .Z(n5531) );
  XNOR U6116 ( .A(n5532), .B(n5531), .Z(n5533) );
  NAND U6117 ( .A(b[0]), .B(a[51]), .Z(n5463) );
  XNOR U6118 ( .A(b[1]), .B(n5463), .Z(n5465) );
  NANDN U6119 ( .A(b[0]), .B(a[50]), .Z(n5464) );
  NAND U6120 ( .A(n5465), .B(n5464), .Z(n5534) );
  XNOR U6121 ( .A(n5533), .B(n5534), .Z(n5574) );
  NAND U6122 ( .A(n38185), .B(n5466), .Z(n5468) );
  XOR U6123 ( .A(b[23]), .B(a[29]), .Z(n5613) );
  NAND U6124 ( .A(n38132), .B(n5613), .Z(n5467) );
  AND U6125 ( .A(n5468), .B(n5467), .Z(n5603) );
  NAND U6126 ( .A(n184), .B(n5469), .Z(n5471) );
  XOR U6127 ( .A(b[7]), .B(a[45]), .Z(n5616) );
  NAND U6128 ( .A(n36592), .B(n5616), .Z(n5470) );
  AND U6129 ( .A(n5471), .B(n5470), .Z(n5602) );
  NAND U6130 ( .A(n38289), .B(n5472), .Z(n5474) );
  XOR U6131 ( .A(b[25]), .B(a[27]), .Z(n5619) );
  NAND U6132 ( .A(n38247), .B(n5619), .Z(n5473) );
  NAND U6133 ( .A(n5474), .B(n5473), .Z(n5601) );
  XOR U6134 ( .A(n5602), .B(n5601), .Z(n5604) );
  XOR U6135 ( .A(n5603), .B(n5604), .Z(n5573) );
  XOR U6136 ( .A(n5574), .B(n5573), .Z(n5576) );
  NAND U6137 ( .A(n187), .B(n5475), .Z(n5477) );
  XOR U6138 ( .A(b[13]), .B(a[39]), .Z(n5622) );
  NAND U6139 ( .A(n37295), .B(n5622), .Z(n5476) );
  AND U6140 ( .A(n5477), .B(n5476), .Z(n5568) );
  NAND U6141 ( .A(n186), .B(n5478), .Z(n5480) );
  XOR U6142 ( .A(b[11]), .B(a[41]), .Z(n5625) );
  NAND U6143 ( .A(n37097), .B(n5625), .Z(n5479) );
  NAND U6144 ( .A(n5480), .B(n5479), .Z(n5567) );
  XNOR U6145 ( .A(n5568), .B(n5567), .Z(n5570) );
  NAND U6146 ( .A(n188), .B(n5481), .Z(n5483) );
  XOR U6147 ( .A(b[15]), .B(a[37]), .Z(n5628) );
  NAND U6148 ( .A(n37382), .B(n5628), .Z(n5482) );
  AND U6149 ( .A(n5483), .B(n5482), .Z(n5564) );
  NAND U6150 ( .A(n38064), .B(n5484), .Z(n5486) );
  XOR U6151 ( .A(b[21]), .B(a[31]), .Z(n5631) );
  NAND U6152 ( .A(n37993), .B(n5631), .Z(n5485) );
  AND U6153 ( .A(n5486), .B(n5485), .Z(n5562) );
  NAND U6154 ( .A(n185), .B(n5487), .Z(n5489) );
  XOR U6155 ( .A(b[9]), .B(a[43]), .Z(n5634) );
  NAND U6156 ( .A(n36805), .B(n5634), .Z(n5488) );
  NAND U6157 ( .A(n5489), .B(n5488), .Z(n5561) );
  XNOR U6158 ( .A(n5562), .B(n5561), .Z(n5563) );
  XNOR U6159 ( .A(n5564), .B(n5563), .Z(n5569) );
  XOR U6160 ( .A(n5570), .B(n5569), .Z(n5575) );
  XNOR U6161 ( .A(n5576), .B(n5575), .Z(n5587) );
  XNOR U6162 ( .A(n5588), .B(n5587), .Z(n5519) );
  XNOR U6163 ( .A(n5520), .B(n5519), .Z(n5521) );
  XOR U6164 ( .A(n5522), .B(n5521), .Z(n5638) );
  XNOR U6165 ( .A(n5637), .B(n5638), .Z(n5639) );
  XNOR U6166 ( .A(n5640), .B(n5639), .Z(n5515) );
  XOR U6167 ( .A(n5516), .B(n5515), .Z(n5508) );
  NANDN U6168 ( .A(n5491), .B(n5490), .Z(n5495) );
  OR U6169 ( .A(n5493), .B(n5492), .Z(n5494) );
  AND U6170 ( .A(n5495), .B(n5494), .Z(n5507) );
  XNOR U6171 ( .A(n5508), .B(n5507), .Z(n5509) );
  XNOR U6172 ( .A(n5510), .B(n5509), .Z(n5501) );
  XNOR U6173 ( .A(n5502), .B(n5501), .Z(n5503) );
  XNOR U6174 ( .A(n5504), .B(n5503), .Z(n5643) );
  XNOR U6175 ( .A(sreg[275]), .B(n5643), .Z(n5645) );
  NANDN U6176 ( .A(sreg[274]), .B(n5496), .Z(n5500) );
  NAND U6177 ( .A(n5498), .B(n5497), .Z(n5499) );
  NAND U6178 ( .A(n5500), .B(n5499), .Z(n5644) );
  XNOR U6179 ( .A(n5645), .B(n5644), .Z(c[275]) );
  NANDN U6180 ( .A(n5502), .B(n5501), .Z(n5506) );
  NANDN U6181 ( .A(n5504), .B(n5503), .Z(n5505) );
  AND U6182 ( .A(n5506), .B(n5505), .Z(n5651) );
  NANDN U6183 ( .A(n5508), .B(n5507), .Z(n5512) );
  NANDN U6184 ( .A(n5510), .B(n5509), .Z(n5511) );
  AND U6185 ( .A(n5512), .B(n5511), .Z(n5649) );
  NANDN U6186 ( .A(n5514), .B(n5513), .Z(n5518) );
  NAND U6187 ( .A(n5516), .B(n5515), .Z(n5517) );
  AND U6188 ( .A(n5518), .B(n5517), .Z(n5656) );
  NANDN U6189 ( .A(n5520), .B(n5519), .Z(n5524) );
  NANDN U6190 ( .A(n5522), .B(n5521), .Z(n5523) );
  AND U6191 ( .A(n5524), .B(n5523), .Z(n5787) );
  NANDN U6192 ( .A(n5526), .B(n5525), .Z(n5530) );
  NAND U6193 ( .A(n5528), .B(n5527), .Z(n5529) );
  AND U6194 ( .A(n5530), .B(n5529), .Z(n5786) );
  XNOR U6195 ( .A(n5787), .B(n5786), .Z(n5789) );
  NANDN U6196 ( .A(n5532), .B(n5531), .Z(n5536) );
  NANDN U6197 ( .A(n5534), .B(n5533), .Z(n5535) );
  AND U6198 ( .A(n5536), .B(n5535), .Z(n5722) );
  NAND U6199 ( .A(n38385), .B(n5537), .Z(n5539) );
  XOR U6200 ( .A(b[27]), .B(a[26]), .Z(n5666) );
  NAND U6201 ( .A(n38343), .B(n5666), .Z(n5538) );
  AND U6202 ( .A(n5539), .B(n5538), .Z(n5729) );
  NAND U6203 ( .A(n183), .B(n5540), .Z(n5542) );
  XOR U6204 ( .A(b[5]), .B(a[48]), .Z(n5669) );
  NAND U6205 ( .A(n36296), .B(n5669), .Z(n5541) );
  AND U6206 ( .A(n5542), .B(n5541), .Z(n5727) );
  NAND U6207 ( .A(n190), .B(n5543), .Z(n5545) );
  XOR U6208 ( .A(b[19]), .B(a[34]), .Z(n5672) );
  NAND U6209 ( .A(n37821), .B(n5672), .Z(n5544) );
  NAND U6210 ( .A(n5545), .B(n5544), .Z(n5726) );
  XNOR U6211 ( .A(n5727), .B(n5726), .Z(n5728) );
  XNOR U6212 ( .A(n5729), .B(n5728), .Z(n5720) );
  NAND U6213 ( .A(n38470), .B(n5546), .Z(n5548) );
  XOR U6214 ( .A(b[31]), .B(a[22]), .Z(n5675) );
  NAND U6215 ( .A(n38453), .B(n5675), .Z(n5547) );
  AND U6216 ( .A(n5548), .B(n5547), .Z(n5687) );
  NAND U6217 ( .A(n181), .B(n5549), .Z(n5551) );
  XOR U6218 ( .A(b[3]), .B(a[50]), .Z(n5678) );
  NAND U6219 ( .A(n182), .B(n5678), .Z(n5550) );
  AND U6220 ( .A(n5551), .B(n5550), .Z(n5685) );
  NAND U6221 ( .A(n189), .B(n5552), .Z(n5554) );
  XOR U6222 ( .A(b[17]), .B(a[36]), .Z(n5681) );
  NAND U6223 ( .A(n37652), .B(n5681), .Z(n5553) );
  NAND U6224 ( .A(n5554), .B(n5553), .Z(n5684) );
  XNOR U6225 ( .A(n5685), .B(n5684), .Z(n5686) );
  XOR U6226 ( .A(n5687), .B(n5686), .Z(n5721) );
  XOR U6227 ( .A(n5720), .B(n5721), .Z(n5723) );
  XOR U6228 ( .A(n5722), .B(n5723), .Z(n5769) );
  NANDN U6229 ( .A(n5556), .B(n5555), .Z(n5560) );
  NANDN U6230 ( .A(n5558), .B(n5557), .Z(n5559) );
  AND U6231 ( .A(n5560), .B(n5559), .Z(n5708) );
  NANDN U6232 ( .A(n5562), .B(n5561), .Z(n5566) );
  NANDN U6233 ( .A(n5564), .B(n5563), .Z(n5565) );
  NAND U6234 ( .A(n5566), .B(n5565), .Z(n5709) );
  XNOR U6235 ( .A(n5708), .B(n5709), .Z(n5710) );
  NANDN U6236 ( .A(n5568), .B(n5567), .Z(n5572) );
  NAND U6237 ( .A(n5570), .B(n5569), .Z(n5571) );
  NAND U6238 ( .A(n5572), .B(n5571), .Z(n5711) );
  XNOR U6239 ( .A(n5710), .B(n5711), .Z(n5768) );
  XNOR U6240 ( .A(n5769), .B(n5768), .Z(n5771) );
  NAND U6241 ( .A(n5574), .B(n5573), .Z(n5578) );
  NAND U6242 ( .A(n5576), .B(n5575), .Z(n5577) );
  AND U6243 ( .A(n5578), .B(n5577), .Z(n5770) );
  XOR U6244 ( .A(n5771), .B(n5770), .Z(n5783) );
  NANDN U6245 ( .A(n5580), .B(n5579), .Z(n5584) );
  NANDN U6246 ( .A(n5582), .B(n5581), .Z(n5583) );
  AND U6247 ( .A(n5584), .B(n5583), .Z(n5780) );
  NANDN U6248 ( .A(n5590), .B(n5589), .Z(n5594) );
  OR U6249 ( .A(n5592), .B(n5591), .Z(n5593) );
  AND U6250 ( .A(n5594), .B(n5593), .Z(n5775) );
  NANDN U6251 ( .A(n5596), .B(n5595), .Z(n5600) );
  NANDN U6252 ( .A(n5598), .B(n5597), .Z(n5599) );
  AND U6253 ( .A(n5600), .B(n5599), .Z(n5715) );
  NANDN U6254 ( .A(n5602), .B(n5601), .Z(n5606) );
  OR U6255 ( .A(n5604), .B(n5603), .Z(n5605) );
  NAND U6256 ( .A(n5606), .B(n5605), .Z(n5714) );
  XNOR U6257 ( .A(n5715), .B(n5714), .Z(n5716) );
  NAND U6258 ( .A(n194), .B(n5607), .Z(n5609) );
  XOR U6259 ( .A(b[29]), .B(a[24]), .Z(n5741) );
  NAND U6260 ( .A(n38456), .B(n5741), .Z(n5608) );
  AND U6261 ( .A(n5609), .B(n5608), .Z(n5661) );
  AND U6262 ( .A(b[31]), .B(a[20]), .Z(n5660) );
  XNOR U6263 ( .A(n5661), .B(n5660), .Z(n5662) );
  NAND U6264 ( .A(b[0]), .B(a[52]), .Z(n5610) );
  XNOR U6265 ( .A(b[1]), .B(n5610), .Z(n5612) );
  NANDN U6266 ( .A(b[0]), .B(a[51]), .Z(n5611) );
  NAND U6267 ( .A(n5612), .B(n5611), .Z(n5663) );
  XNOR U6268 ( .A(n5662), .B(n5663), .Z(n5702) );
  NAND U6269 ( .A(n38185), .B(n5613), .Z(n5615) );
  XOR U6270 ( .A(b[23]), .B(a[30]), .Z(n5744) );
  NAND U6271 ( .A(n38132), .B(n5744), .Z(n5614) );
  AND U6272 ( .A(n5615), .B(n5614), .Z(n5735) );
  NAND U6273 ( .A(n184), .B(n5616), .Z(n5618) );
  XOR U6274 ( .A(b[7]), .B(a[46]), .Z(n5747) );
  NAND U6275 ( .A(n36592), .B(n5747), .Z(n5617) );
  AND U6276 ( .A(n5618), .B(n5617), .Z(n5733) );
  NAND U6277 ( .A(n38289), .B(n5619), .Z(n5621) );
  XOR U6278 ( .A(b[25]), .B(a[28]), .Z(n5750) );
  NAND U6279 ( .A(n38247), .B(n5750), .Z(n5620) );
  NAND U6280 ( .A(n5621), .B(n5620), .Z(n5732) );
  XNOR U6281 ( .A(n5733), .B(n5732), .Z(n5734) );
  XOR U6282 ( .A(n5735), .B(n5734), .Z(n5703) );
  XNOR U6283 ( .A(n5702), .B(n5703), .Z(n5704) );
  NAND U6284 ( .A(n187), .B(n5622), .Z(n5624) );
  XOR U6285 ( .A(b[13]), .B(a[40]), .Z(n5753) );
  NAND U6286 ( .A(n37295), .B(n5753), .Z(n5623) );
  AND U6287 ( .A(n5624), .B(n5623), .Z(n5697) );
  NAND U6288 ( .A(n186), .B(n5625), .Z(n5627) );
  XOR U6289 ( .A(b[11]), .B(a[42]), .Z(n5756) );
  NAND U6290 ( .A(n37097), .B(n5756), .Z(n5626) );
  NAND U6291 ( .A(n5627), .B(n5626), .Z(n5696) );
  XNOR U6292 ( .A(n5697), .B(n5696), .Z(n5698) );
  NAND U6293 ( .A(n188), .B(n5628), .Z(n5630) );
  XOR U6294 ( .A(b[15]), .B(a[38]), .Z(n5759) );
  NAND U6295 ( .A(n37382), .B(n5759), .Z(n5629) );
  AND U6296 ( .A(n5630), .B(n5629), .Z(n5693) );
  NAND U6297 ( .A(n38064), .B(n5631), .Z(n5633) );
  XOR U6298 ( .A(b[21]), .B(a[32]), .Z(n5762) );
  NAND U6299 ( .A(n37993), .B(n5762), .Z(n5632) );
  AND U6300 ( .A(n5633), .B(n5632), .Z(n5691) );
  NAND U6301 ( .A(n185), .B(n5634), .Z(n5636) );
  XOR U6302 ( .A(b[9]), .B(a[44]), .Z(n5765) );
  NAND U6303 ( .A(n36805), .B(n5765), .Z(n5635) );
  NAND U6304 ( .A(n5636), .B(n5635), .Z(n5690) );
  XNOR U6305 ( .A(n5691), .B(n5690), .Z(n5692) );
  XOR U6306 ( .A(n5693), .B(n5692), .Z(n5699) );
  XOR U6307 ( .A(n5698), .B(n5699), .Z(n5705) );
  XOR U6308 ( .A(n5704), .B(n5705), .Z(n5717) );
  XNOR U6309 ( .A(n5716), .B(n5717), .Z(n5774) );
  XNOR U6310 ( .A(n5775), .B(n5774), .Z(n5776) );
  XOR U6311 ( .A(n5777), .B(n5776), .Z(n5781) );
  XNOR U6312 ( .A(n5780), .B(n5781), .Z(n5782) );
  XNOR U6313 ( .A(n5783), .B(n5782), .Z(n5788) );
  XOR U6314 ( .A(n5789), .B(n5788), .Z(n5655) );
  NANDN U6315 ( .A(n5638), .B(n5637), .Z(n5642) );
  NANDN U6316 ( .A(n5640), .B(n5639), .Z(n5641) );
  AND U6317 ( .A(n5642), .B(n5641), .Z(n5654) );
  XOR U6318 ( .A(n5655), .B(n5654), .Z(n5657) );
  XNOR U6319 ( .A(n5656), .B(n5657), .Z(n5648) );
  XNOR U6320 ( .A(n5649), .B(n5648), .Z(n5650) );
  XNOR U6321 ( .A(n5651), .B(n5650), .Z(n5792) );
  XNOR U6322 ( .A(sreg[276]), .B(n5792), .Z(n5794) );
  NANDN U6323 ( .A(sreg[275]), .B(n5643), .Z(n5647) );
  NAND U6324 ( .A(n5645), .B(n5644), .Z(n5646) );
  NAND U6325 ( .A(n5647), .B(n5646), .Z(n5793) );
  XNOR U6326 ( .A(n5794), .B(n5793), .Z(c[276]) );
  NANDN U6327 ( .A(n5649), .B(n5648), .Z(n5653) );
  NANDN U6328 ( .A(n5651), .B(n5650), .Z(n5652) );
  AND U6329 ( .A(n5653), .B(n5652), .Z(n5800) );
  NANDN U6330 ( .A(n5655), .B(n5654), .Z(n5659) );
  NANDN U6331 ( .A(n5657), .B(n5656), .Z(n5658) );
  AND U6332 ( .A(n5659), .B(n5658), .Z(n5798) );
  NANDN U6333 ( .A(n5661), .B(n5660), .Z(n5665) );
  NANDN U6334 ( .A(n5663), .B(n5662), .Z(n5664) );
  AND U6335 ( .A(n5665), .B(n5664), .Z(n5889) );
  NAND U6336 ( .A(n38385), .B(n5666), .Z(n5668) );
  XOR U6337 ( .A(b[27]), .B(a[27]), .Z(n5833) );
  NAND U6338 ( .A(n38343), .B(n5833), .Z(n5667) );
  AND U6339 ( .A(n5668), .B(n5667), .Z(n5896) );
  NAND U6340 ( .A(n183), .B(n5669), .Z(n5671) );
  XOR U6341 ( .A(b[5]), .B(a[49]), .Z(n5836) );
  NAND U6342 ( .A(n36296), .B(n5836), .Z(n5670) );
  AND U6343 ( .A(n5671), .B(n5670), .Z(n5894) );
  NAND U6344 ( .A(n190), .B(n5672), .Z(n5674) );
  XOR U6345 ( .A(b[19]), .B(a[35]), .Z(n5839) );
  NAND U6346 ( .A(n37821), .B(n5839), .Z(n5673) );
  NAND U6347 ( .A(n5674), .B(n5673), .Z(n5893) );
  XNOR U6348 ( .A(n5894), .B(n5893), .Z(n5895) );
  XNOR U6349 ( .A(n5896), .B(n5895), .Z(n5887) );
  NAND U6350 ( .A(n38470), .B(n5675), .Z(n5677) );
  XOR U6351 ( .A(b[31]), .B(a[23]), .Z(n5842) );
  NAND U6352 ( .A(n38453), .B(n5842), .Z(n5676) );
  AND U6353 ( .A(n5677), .B(n5676), .Z(n5854) );
  NAND U6354 ( .A(n181), .B(n5678), .Z(n5680) );
  XOR U6355 ( .A(b[3]), .B(a[51]), .Z(n5845) );
  NAND U6356 ( .A(n182), .B(n5845), .Z(n5679) );
  AND U6357 ( .A(n5680), .B(n5679), .Z(n5852) );
  NAND U6358 ( .A(n189), .B(n5681), .Z(n5683) );
  XOR U6359 ( .A(b[17]), .B(a[37]), .Z(n5848) );
  NAND U6360 ( .A(n37652), .B(n5848), .Z(n5682) );
  NAND U6361 ( .A(n5683), .B(n5682), .Z(n5851) );
  XNOR U6362 ( .A(n5852), .B(n5851), .Z(n5853) );
  XOR U6363 ( .A(n5854), .B(n5853), .Z(n5888) );
  XOR U6364 ( .A(n5887), .B(n5888), .Z(n5890) );
  XOR U6365 ( .A(n5889), .B(n5890), .Z(n5822) );
  NANDN U6366 ( .A(n5685), .B(n5684), .Z(n5689) );
  NANDN U6367 ( .A(n5687), .B(n5686), .Z(n5688) );
  AND U6368 ( .A(n5689), .B(n5688), .Z(n5875) );
  NANDN U6369 ( .A(n5691), .B(n5690), .Z(n5695) );
  NANDN U6370 ( .A(n5693), .B(n5692), .Z(n5694) );
  NAND U6371 ( .A(n5695), .B(n5694), .Z(n5876) );
  XNOR U6372 ( .A(n5875), .B(n5876), .Z(n5877) );
  NANDN U6373 ( .A(n5697), .B(n5696), .Z(n5701) );
  NANDN U6374 ( .A(n5699), .B(n5698), .Z(n5700) );
  NAND U6375 ( .A(n5701), .B(n5700), .Z(n5878) );
  XNOR U6376 ( .A(n5877), .B(n5878), .Z(n5821) );
  XNOR U6377 ( .A(n5822), .B(n5821), .Z(n5824) );
  NANDN U6378 ( .A(n5703), .B(n5702), .Z(n5707) );
  NANDN U6379 ( .A(n5705), .B(n5704), .Z(n5706) );
  AND U6380 ( .A(n5707), .B(n5706), .Z(n5823) );
  XOR U6381 ( .A(n5824), .B(n5823), .Z(n5937) );
  NANDN U6382 ( .A(n5709), .B(n5708), .Z(n5713) );
  NANDN U6383 ( .A(n5711), .B(n5710), .Z(n5712) );
  AND U6384 ( .A(n5713), .B(n5712), .Z(n5935) );
  NANDN U6385 ( .A(n5715), .B(n5714), .Z(n5719) );
  NANDN U6386 ( .A(n5717), .B(n5716), .Z(n5718) );
  AND U6387 ( .A(n5719), .B(n5718), .Z(n5818) );
  NANDN U6388 ( .A(n5721), .B(n5720), .Z(n5725) );
  OR U6389 ( .A(n5723), .B(n5722), .Z(n5724) );
  AND U6390 ( .A(n5725), .B(n5724), .Z(n5816) );
  NANDN U6391 ( .A(n5727), .B(n5726), .Z(n5731) );
  NANDN U6392 ( .A(n5729), .B(n5728), .Z(n5730) );
  AND U6393 ( .A(n5731), .B(n5730), .Z(n5882) );
  NANDN U6394 ( .A(n5733), .B(n5732), .Z(n5737) );
  NANDN U6395 ( .A(n5735), .B(n5734), .Z(n5736) );
  NAND U6396 ( .A(n5737), .B(n5736), .Z(n5881) );
  XNOR U6397 ( .A(n5882), .B(n5881), .Z(n5883) );
  NAND U6398 ( .A(b[0]), .B(a[53]), .Z(n5738) );
  XNOR U6399 ( .A(b[1]), .B(n5738), .Z(n5740) );
  NANDN U6400 ( .A(b[0]), .B(a[52]), .Z(n5739) );
  NAND U6401 ( .A(n5740), .B(n5739), .Z(n5830) );
  NAND U6402 ( .A(n194), .B(n5741), .Z(n5743) );
  XOR U6403 ( .A(b[29]), .B(a[25]), .Z(n5908) );
  NAND U6404 ( .A(n38456), .B(n5908), .Z(n5742) );
  AND U6405 ( .A(n5743), .B(n5742), .Z(n5828) );
  AND U6406 ( .A(b[31]), .B(a[21]), .Z(n5827) );
  XNOR U6407 ( .A(n5828), .B(n5827), .Z(n5829) );
  XNOR U6408 ( .A(n5830), .B(n5829), .Z(n5869) );
  NAND U6409 ( .A(n38185), .B(n5744), .Z(n5746) );
  XOR U6410 ( .A(b[23]), .B(a[31]), .Z(n5911) );
  NAND U6411 ( .A(n38132), .B(n5911), .Z(n5745) );
  AND U6412 ( .A(n5746), .B(n5745), .Z(n5902) );
  NAND U6413 ( .A(n184), .B(n5747), .Z(n5749) );
  XOR U6414 ( .A(b[7]), .B(a[47]), .Z(n5914) );
  NAND U6415 ( .A(n36592), .B(n5914), .Z(n5748) );
  AND U6416 ( .A(n5749), .B(n5748), .Z(n5900) );
  NAND U6417 ( .A(n38289), .B(n5750), .Z(n5752) );
  XOR U6418 ( .A(b[25]), .B(a[29]), .Z(n5917) );
  NAND U6419 ( .A(n38247), .B(n5917), .Z(n5751) );
  NAND U6420 ( .A(n5752), .B(n5751), .Z(n5899) );
  XNOR U6421 ( .A(n5900), .B(n5899), .Z(n5901) );
  XOR U6422 ( .A(n5902), .B(n5901), .Z(n5870) );
  XNOR U6423 ( .A(n5869), .B(n5870), .Z(n5871) );
  NAND U6424 ( .A(n187), .B(n5753), .Z(n5755) );
  XOR U6425 ( .A(b[13]), .B(a[41]), .Z(n5920) );
  NAND U6426 ( .A(n37295), .B(n5920), .Z(n5754) );
  AND U6427 ( .A(n5755), .B(n5754), .Z(n5864) );
  NAND U6428 ( .A(n186), .B(n5756), .Z(n5758) );
  XOR U6429 ( .A(b[11]), .B(a[43]), .Z(n5923) );
  NAND U6430 ( .A(n37097), .B(n5923), .Z(n5757) );
  NAND U6431 ( .A(n5758), .B(n5757), .Z(n5863) );
  XNOR U6432 ( .A(n5864), .B(n5863), .Z(n5865) );
  NAND U6433 ( .A(n188), .B(n5759), .Z(n5761) );
  XOR U6434 ( .A(b[15]), .B(a[39]), .Z(n5926) );
  NAND U6435 ( .A(n37382), .B(n5926), .Z(n5760) );
  AND U6436 ( .A(n5761), .B(n5760), .Z(n5860) );
  NAND U6437 ( .A(n38064), .B(n5762), .Z(n5764) );
  XOR U6438 ( .A(b[21]), .B(a[33]), .Z(n5929) );
  NAND U6439 ( .A(n37993), .B(n5929), .Z(n5763) );
  AND U6440 ( .A(n5764), .B(n5763), .Z(n5858) );
  NAND U6441 ( .A(n185), .B(n5765), .Z(n5767) );
  XOR U6442 ( .A(b[9]), .B(a[45]), .Z(n5932) );
  NAND U6443 ( .A(n36805), .B(n5932), .Z(n5766) );
  NAND U6444 ( .A(n5767), .B(n5766), .Z(n5857) );
  XNOR U6445 ( .A(n5858), .B(n5857), .Z(n5859) );
  XOR U6446 ( .A(n5860), .B(n5859), .Z(n5866) );
  XOR U6447 ( .A(n5865), .B(n5866), .Z(n5872) );
  XOR U6448 ( .A(n5871), .B(n5872), .Z(n5884) );
  XNOR U6449 ( .A(n5883), .B(n5884), .Z(n5815) );
  XNOR U6450 ( .A(n5816), .B(n5815), .Z(n5817) );
  XOR U6451 ( .A(n5818), .B(n5817), .Z(n5936) );
  XOR U6452 ( .A(n5935), .B(n5936), .Z(n5938) );
  XOR U6453 ( .A(n5937), .B(n5938), .Z(n5812) );
  NANDN U6454 ( .A(n5769), .B(n5768), .Z(n5773) );
  NAND U6455 ( .A(n5771), .B(n5770), .Z(n5772) );
  AND U6456 ( .A(n5773), .B(n5772), .Z(n5810) );
  NANDN U6457 ( .A(n5775), .B(n5774), .Z(n5779) );
  NANDN U6458 ( .A(n5777), .B(n5776), .Z(n5778) );
  AND U6459 ( .A(n5779), .B(n5778), .Z(n5809) );
  XNOR U6460 ( .A(n5810), .B(n5809), .Z(n5811) );
  XNOR U6461 ( .A(n5812), .B(n5811), .Z(n5803) );
  NANDN U6462 ( .A(n5781), .B(n5780), .Z(n5785) );
  NANDN U6463 ( .A(n5783), .B(n5782), .Z(n5784) );
  NAND U6464 ( .A(n5785), .B(n5784), .Z(n5804) );
  XNOR U6465 ( .A(n5803), .B(n5804), .Z(n5805) );
  NANDN U6466 ( .A(n5787), .B(n5786), .Z(n5791) );
  NAND U6467 ( .A(n5789), .B(n5788), .Z(n5790) );
  NAND U6468 ( .A(n5791), .B(n5790), .Z(n5806) );
  XNOR U6469 ( .A(n5805), .B(n5806), .Z(n5797) );
  XNOR U6470 ( .A(n5798), .B(n5797), .Z(n5799) );
  XNOR U6471 ( .A(n5800), .B(n5799), .Z(n5941) );
  XNOR U6472 ( .A(sreg[277]), .B(n5941), .Z(n5943) );
  NANDN U6473 ( .A(sreg[276]), .B(n5792), .Z(n5796) );
  NAND U6474 ( .A(n5794), .B(n5793), .Z(n5795) );
  NAND U6475 ( .A(n5796), .B(n5795), .Z(n5942) );
  XNOR U6476 ( .A(n5943), .B(n5942), .Z(c[277]) );
  NANDN U6477 ( .A(n5798), .B(n5797), .Z(n5802) );
  NANDN U6478 ( .A(n5800), .B(n5799), .Z(n5801) );
  AND U6479 ( .A(n5802), .B(n5801), .Z(n5949) );
  NANDN U6480 ( .A(n5804), .B(n5803), .Z(n5808) );
  NANDN U6481 ( .A(n5806), .B(n5805), .Z(n5807) );
  AND U6482 ( .A(n5808), .B(n5807), .Z(n5947) );
  NANDN U6483 ( .A(n5810), .B(n5809), .Z(n5814) );
  NANDN U6484 ( .A(n5812), .B(n5811), .Z(n5813) );
  AND U6485 ( .A(n5814), .B(n5813), .Z(n5955) );
  NANDN U6486 ( .A(n5816), .B(n5815), .Z(n5820) );
  NANDN U6487 ( .A(n5818), .B(n5817), .Z(n5819) );
  AND U6488 ( .A(n5820), .B(n5819), .Z(n5959) );
  NANDN U6489 ( .A(n5822), .B(n5821), .Z(n5826) );
  NAND U6490 ( .A(n5824), .B(n5823), .Z(n5825) );
  AND U6491 ( .A(n5826), .B(n5825), .Z(n5958) );
  XNOR U6492 ( .A(n5959), .B(n5958), .Z(n5961) );
  NANDN U6493 ( .A(n5828), .B(n5827), .Z(n5832) );
  NANDN U6494 ( .A(n5830), .B(n5829), .Z(n5831) );
  AND U6495 ( .A(n5832), .B(n5831), .Z(n6038) );
  NAND U6496 ( .A(n38385), .B(n5833), .Z(n5835) );
  XOR U6497 ( .A(b[27]), .B(a[28]), .Z(n5982) );
  NAND U6498 ( .A(n38343), .B(n5982), .Z(n5834) );
  AND U6499 ( .A(n5835), .B(n5834), .Z(n6045) );
  NAND U6500 ( .A(n183), .B(n5836), .Z(n5838) );
  XOR U6501 ( .A(b[5]), .B(a[50]), .Z(n5985) );
  NAND U6502 ( .A(n36296), .B(n5985), .Z(n5837) );
  AND U6503 ( .A(n5838), .B(n5837), .Z(n6043) );
  NAND U6504 ( .A(n190), .B(n5839), .Z(n5841) );
  XOR U6505 ( .A(b[19]), .B(a[36]), .Z(n5988) );
  NAND U6506 ( .A(n37821), .B(n5988), .Z(n5840) );
  NAND U6507 ( .A(n5841), .B(n5840), .Z(n6042) );
  XNOR U6508 ( .A(n6043), .B(n6042), .Z(n6044) );
  XNOR U6509 ( .A(n6045), .B(n6044), .Z(n6036) );
  NAND U6510 ( .A(n38470), .B(n5842), .Z(n5844) );
  XOR U6511 ( .A(b[31]), .B(a[24]), .Z(n5991) );
  NAND U6512 ( .A(n38453), .B(n5991), .Z(n5843) );
  AND U6513 ( .A(n5844), .B(n5843), .Z(n6003) );
  NAND U6514 ( .A(n181), .B(n5845), .Z(n5847) );
  XOR U6515 ( .A(b[3]), .B(a[52]), .Z(n5994) );
  NAND U6516 ( .A(n182), .B(n5994), .Z(n5846) );
  AND U6517 ( .A(n5847), .B(n5846), .Z(n6001) );
  NAND U6518 ( .A(n189), .B(n5848), .Z(n5850) );
  XOR U6519 ( .A(b[17]), .B(a[38]), .Z(n5997) );
  NAND U6520 ( .A(n37652), .B(n5997), .Z(n5849) );
  NAND U6521 ( .A(n5850), .B(n5849), .Z(n6000) );
  XNOR U6522 ( .A(n6001), .B(n6000), .Z(n6002) );
  XOR U6523 ( .A(n6003), .B(n6002), .Z(n6037) );
  XOR U6524 ( .A(n6036), .B(n6037), .Z(n6039) );
  XOR U6525 ( .A(n6038), .B(n6039), .Z(n5971) );
  NANDN U6526 ( .A(n5852), .B(n5851), .Z(n5856) );
  NANDN U6527 ( .A(n5854), .B(n5853), .Z(n5855) );
  AND U6528 ( .A(n5856), .B(n5855), .Z(n6024) );
  NANDN U6529 ( .A(n5858), .B(n5857), .Z(n5862) );
  NANDN U6530 ( .A(n5860), .B(n5859), .Z(n5861) );
  NAND U6531 ( .A(n5862), .B(n5861), .Z(n6025) );
  XNOR U6532 ( .A(n6024), .B(n6025), .Z(n6026) );
  NANDN U6533 ( .A(n5864), .B(n5863), .Z(n5868) );
  NANDN U6534 ( .A(n5866), .B(n5865), .Z(n5867) );
  NAND U6535 ( .A(n5868), .B(n5867), .Z(n6027) );
  XNOR U6536 ( .A(n6026), .B(n6027), .Z(n5970) );
  XNOR U6537 ( .A(n5971), .B(n5970), .Z(n5973) );
  NANDN U6538 ( .A(n5870), .B(n5869), .Z(n5874) );
  NANDN U6539 ( .A(n5872), .B(n5871), .Z(n5873) );
  AND U6540 ( .A(n5874), .B(n5873), .Z(n5972) );
  XOR U6541 ( .A(n5973), .B(n5972), .Z(n6087) );
  NANDN U6542 ( .A(n5876), .B(n5875), .Z(n5880) );
  NANDN U6543 ( .A(n5878), .B(n5877), .Z(n5879) );
  AND U6544 ( .A(n5880), .B(n5879), .Z(n6084) );
  NANDN U6545 ( .A(n5882), .B(n5881), .Z(n5886) );
  NANDN U6546 ( .A(n5884), .B(n5883), .Z(n5885) );
  AND U6547 ( .A(n5886), .B(n5885), .Z(n5967) );
  NANDN U6548 ( .A(n5888), .B(n5887), .Z(n5892) );
  OR U6549 ( .A(n5890), .B(n5889), .Z(n5891) );
  AND U6550 ( .A(n5892), .B(n5891), .Z(n5965) );
  NANDN U6551 ( .A(n5894), .B(n5893), .Z(n5898) );
  NANDN U6552 ( .A(n5896), .B(n5895), .Z(n5897) );
  AND U6553 ( .A(n5898), .B(n5897), .Z(n6031) );
  NANDN U6554 ( .A(n5900), .B(n5899), .Z(n5904) );
  NANDN U6555 ( .A(n5902), .B(n5901), .Z(n5903) );
  NAND U6556 ( .A(n5904), .B(n5903), .Z(n6030) );
  XNOR U6557 ( .A(n6031), .B(n6030), .Z(n6032) );
  NAND U6558 ( .A(b[0]), .B(a[54]), .Z(n5905) );
  XNOR U6559 ( .A(b[1]), .B(n5905), .Z(n5907) );
  NANDN U6560 ( .A(b[0]), .B(a[53]), .Z(n5906) );
  NAND U6561 ( .A(n5907), .B(n5906), .Z(n5979) );
  NAND U6562 ( .A(n194), .B(n5908), .Z(n5910) );
  XOR U6563 ( .A(b[29]), .B(a[26]), .Z(n6054) );
  NAND U6564 ( .A(n38456), .B(n6054), .Z(n5909) );
  AND U6565 ( .A(n5910), .B(n5909), .Z(n5977) );
  AND U6566 ( .A(b[31]), .B(a[22]), .Z(n5976) );
  XNOR U6567 ( .A(n5977), .B(n5976), .Z(n5978) );
  XNOR U6568 ( .A(n5979), .B(n5978), .Z(n6018) );
  NAND U6569 ( .A(n38185), .B(n5911), .Z(n5913) );
  XOR U6570 ( .A(b[23]), .B(a[32]), .Z(n6060) );
  NAND U6571 ( .A(n38132), .B(n6060), .Z(n5912) );
  AND U6572 ( .A(n5913), .B(n5912), .Z(n6051) );
  NAND U6573 ( .A(n184), .B(n5914), .Z(n5916) );
  XOR U6574 ( .A(b[7]), .B(a[48]), .Z(n6063) );
  NAND U6575 ( .A(n36592), .B(n6063), .Z(n5915) );
  AND U6576 ( .A(n5916), .B(n5915), .Z(n6049) );
  NAND U6577 ( .A(n38289), .B(n5917), .Z(n5919) );
  XOR U6578 ( .A(b[25]), .B(a[30]), .Z(n6066) );
  NAND U6579 ( .A(n38247), .B(n6066), .Z(n5918) );
  NAND U6580 ( .A(n5919), .B(n5918), .Z(n6048) );
  XNOR U6581 ( .A(n6049), .B(n6048), .Z(n6050) );
  XOR U6582 ( .A(n6051), .B(n6050), .Z(n6019) );
  XNOR U6583 ( .A(n6018), .B(n6019), .Z(n6020) );
  NAND U6584 ( .A(n187), .B(n5920), .Z(n5922) );
  XOR U6585 ( .A(b[13]), .B(a[42]), .Z(n6069) );
  NAND U6586 ( .A(n37295), .B(n6069), .Z(n5921) );
  AND U6587 ( .A(n5922), .B(n5921), .Z(n6013) );
  NAND U6588 ( .A(n186), .B(n5923), .Z(n5925) );
  XOR U6589 ( .A(b[11]), .B(a[44]), .Z(n6072) );
  NAND U6590 ( .A(n37097), .B(n6072), .Z(n5924) );
  NAND U6591 ( .A(n5925), .B(n5924), .Z(n6012) );
  XNOR U6592 ( .A(n6013), .B(n6012), .Z(n6014) );
  NAND U6593 ( .A(n188), .B(n5926), .Z(n5928) );
  XOR U6594 ( .A(b[15]), .B(a[40]), .Z(n6075) );
  NAND U6595 ( .A(n37382), .B(n6075), .Z(n5927) );
  AND U6596 ( .A(n5928), .B(n5927), .Z(n6009) );
  NAND U6597 ( .A(n38064), .B(n5929), .Z(n5931) );
  XOR U6598 ( .A(b[21]), .B(a[34]), .Z(n6078) );
  NAND U6599 ( .A(n37993), .B(n6078), .Z(n5930) );
  AND U6600 ( .A(n5931), .B(n5930), .Z(n6007) );
  NAND U6601 ( .A(n185), .B(n5932), .Z(n5934) );
  XOR U6602 ( .A(b[9]), .B(a[46]), .Z(n6081) );
  NAND U6603 ( .A(n36805), .B(n6081), .Z(n5933) );
  NAND U6604 ( .A(n5934), .B(n5933), .Z(n6006) );
  XNOR U6605 ( .A(n6007), .B(n6006), .Z(n6008) );
  XOR U6606 ( .A(n6009), .B(n6008), .Z(n6015) );
  XOR U6607 ( .A(n6014), .B(n6015), .Z(n6021) );
  XOR U6608 ( .A(n6020), .B(n6021), .Z(n6033) );
  XNOR U6609 ( .A(n6032), .B(n6033), .Z(n5964) );
  XNOR U6610 ( .A(n5965), .B(n5964), .Z(n5966) );
  XOR U6611 ( .A(n5967), .B(n5966), .Z(n6085) );
  XNOR U6612 ( .A(n6084), .B(n6085), .Z(n6086) );
  XNOR U6613 ( .A(n6087), .B(n6086), .Z(n5960) );
  XOR U6614 ( .A(n5961), .B(n5960), .Z(n5953) );
  NANDN U6615 ( .A(n5936), .B(n5935), .Z(n5940) );
  OR U6616 ( .A(n5938), .B(n5937), .Z(n5939) );
  AND U6617 ( .A(n5940), .B(n5939), .Z(n5952) );
  XNOR U6618 ( .A(n5953), .B(n5952), .Z(n5954) );
  XNOR U6619 ( .A(n5955), .B(n5954), .Z(n5946) );
  XNOR U6620 ( .A(n5947), .B(n5946), .Z(n5948) );
  XNOR U6621 ( .A(n5949), .B(n5948), .Z(n6090) );
  XNOR U6622 ( .A(sreg[278]), .B(n6090), .Z(n6092) );
  NANDN U6623 ( .A(sreg[277]), .B(n5941), .Z(n5945) );
  NAND U6624 ( .A(n5943), .B(n5942), .Z(n5944) );
  NAND U6625 ( .A(n5945), .B(n5944), .Z(n6091) );
  XNOR U6626 ( .A(n6092), .B(n6091), .Z(c[278]) );
  NANDN U6627 ( .A(n5947), .B(n5946), .Z(n5951) );
  NANDN U6628 ( .A(n5949), .B(n5948), .Z(n5950) );
  AND U6629 ( .A(n5951), .B(n5950), .Z(n6098) );
  NANDN U6630 ( .A(n5953), .B(n5952), .Z(n5957) );
  NANDN U6631 ( .A(n5955), .B(n5954), .Z(n5956) );
  AND U6632 ( .A(n5957), .B(n5956), .Z(n6096) );
  NANDN U6633 ( .A(n5959), .B(n5958), .Z(n5963) );
  NAND U6634 ( .A(n5961), .B(n5960), .Z(n5962) );
  AND U6635 ( .A(n5963), .B(n5962), .Z(n6103) );
  NANDN U6636 ( .A(n5965), .B(n5964), .Z(n5969) );
  NANDN U6637 ( .A(n5967), .B(n5966), .Z(n5968) );
  AND U6638 ( .A(n5969), .B(n5968), .Z(n6108) );
  NANDN U6639 ( .A(n5971), .B(n5970), .Z(n5975) );
  NAND U6640 ( .A(n5973), .B(n5972), .Z(n5974) );
  AND U6641 ( .A(n5975), .B(n5974), .Z(n6107) );
  XNOR U6642 ( .A(n6108), .B(n6107), .Z(n6110) );
  NANDN U6643 ( .A(n5977), .B(n5976), .Z(n5981) );
  NANDN U6644 ( .A(n5979), .B(n5978), .Z(n5980) );
  AND U6645 ( .A(n5981), .B(n5980), .Z(n6185) );
  NAND U6646 ( .A(n38385), .B(n5982), .Z(n5984) );
  XOR U6647 ( .A(b[27]), .B(a[29]), .Z(n6131) );
  NAND U6648 ( .A(n38343), .B(n6131), .Z(n5983) );
  AND U6649 ( .A(n5984), .B(n5983), .Z(n6192) );
  NAND U6650 ( .A(n183), .B(n5985), .Z(n5987) );
  XOR U6651 ( .A(b[5]), .B(a[51]), .Z(n6134) );
  NAND U6652 ( .A(n36296), .B(n6134), .Z(n5986) );
  AND U6653 ( .A(n5987), .B(n5986), .Z(n6190) );
  NAND U6654 ( .A(n190), .B(n5988), .Z(n5990) );
  XOR U6655 ( .A(b[19]), .B(a[37]), .Z(n6137) );
  NAND U6656 ( .A(n37821), .B(n6137), .Z(n5989) );
  NAND U6657 ( .A(n5990), .B(n5989), .Z(n6189) );
  XNOR U6658 ( .A(n6190), .B(n6189), .Z(n6191) );
  XNOR U6659 ( .A(n6192), .B(n6191), .Z(n6183) );
  NAND U6660 ( .A(n38470), .B(n5991), .Z(n5993) );
  XOR U6661 ( .A(b[31]), .B(a[25]), .Z(n6140) );
  NAND U6662 ( .A(n38453), .B(n6140), .Z(n5992) );
  AND U6663 ( .A(n5993), .B(n5992), .Z(n6152) );
  NAND U6664 ( .A(n181), .B(n5994), .Z(n5996) );
  XOR U6665 ( .A(b[3]), .B(a[53]), .Z(n6143) );
  NAND U6666 ( .A(n182), .B(n6143), .Z(n5995) );
  AND U6667 ( .A(n5996), .B(n5995), .Z(n6150) );
  NAND U6668 ( .A(n189), .B(n5997), .Z(n5999) );
  XOR U6669 ( .A(b[17]), .B(a[39]), .Z(n6146) );
  NAND U6670 ( .A(n37652), .B(n6146), .Z(n5998) );
  NAND U6671 ( .A(n5999), .B(n5998), .Z(n6149) );
  XNOR U6672 ( .A(n6150), .B(n6149), .Z(n6151) );
  XOR U6673 ( .A(n6152), .B(n6151), .Z(n6184) );
  XOR U6674 ( .A(n6183), .B(n6184), .Z(n6186) );
  XOR U6675 ( .A(n6185), .B(n6186), .Z(n6120) );
  NANDN U6676 ( .A(n6001), .B(n6000), .Z(n6005) );
  NANDN U6677 ( .A(n6003), .B(n6002), .Z(n6004) );
  AND U6678 ( .A(n6005), .B(n6004), .Z(n6173) );
  NANDN U6679 ( .A(n6007), .B(n6006), .Z(n6011) );
  NANDN U6680 ( .A(n6009), .B(n6008), .Z(n6010) );
  NAND U6681 ( .A(n6011), .B(n6010), .Z(n6174) );
  XNOR U6682 ( .A(n6173), .B(n6174), .Z(n6175) );
  NANDN U6683 ( .A(n6013), .B(n6012), .Z(n6017) );
  NANDN U6684 ( .A(n6015), .B(n6014), .Z(n6016) );
  NAND U6685 ( .A(n6017), .B(n6016), .Z(n6176) );
  XNOR U6686 ( .A(n6175), .B(n6176), .Z(n6119) );
  XNOR U6687 ( .A(n6120), .B(n6119), .Z(n6122) );
  NANDN U6688 ( .A(n6019), .B(n6018), .Z(n6023) );
  NANDN U6689 ( .A(n6021), .B(n6020), .Z(n6022) );
  AND U6690 ( .A(n6023), .B(n6022), .Z(n6121) );
  XOR U6691 ( .A(n6122), .B(n6121), .Z(n6234) );
  NANDN U6692 ( .A(n6025), .B(n6024), .Z(n6029) );
  NANDN U6693 ( .A(n6027), .B(n6026), .Z(n6028) );
  AND U6694 ( .A(n6029), .B(n6028), .Z(n6231) );
  NANDN U6695 ( .A(n6031), .B(n6030), .Z(n6035) );
  NANDN U6696 ( .A(n6033), .B(n6032), .Z(n6034) );
  AND U6697 ( .A(n6035), .B(n6034), .Z(n6116) );
  NANDN U6698 ( .A(n6037), .B(n6036), .Z(n6041) );
  OR U6699 ( .A(n6039), .B(n6038), .Z(n6040) );
  AND U6700 ( .A(n6041), .B(n6040), .Z(n6114) );
  NANDN U6701 ( .A(n6043), .B(n6042), .Z(n6047) );
  NANDN U6702 ( .A(n6045), .B(n6044), .Z(n6046) );
  AND U6703 ( .A(n6047), .B(n6046), .Z(n6180) );
  NANDN U6704 ( .A(n6049), .B(n6048), .Z(n6053) );
  NANDN U6705 ( .A(n6051), .B(n6050), .Z(n6052) );
  NAND U6706 ( .A(n6053), .B(n6052), .Z(n6179) );
  XNOR U6707 ( .A(n6180), .B(n6179), .Z(n6182) );
  NAND U6708 ( .A(n194), .B(n6054), .Z(n6056) );
  XOR U6709 ( .A(b[29]), .B(a[27]), .Z(n6201) );
  NAND U6710 ( .A(n38456), .B(n6201), .Z(n6055) );
  AND U6711 ( .A(n6056), .B(n6055), .Z(n6126) );
  AND U6712 ( .A(b[31]), .B(a[23]), .Z(n6125) );
  XNOR U6713 ( .A(n6126), .B(n6125), .Z(n6127) );
  NAND U6714 ( .A(b[0]), .B(a[55]), .Z(n6057) );
  XNOR U6715 ( .A(b[1]), .B(n6057), .Z(n6059) );
  NANDN U6716 ( .A(b[0]), .B(a[54]), .Z(n6058) );
  NAND U6717 ( .A(n6059), .B(n6058), .Z(n6128) );
  XNOR U6718 ( .A(n6127), .B(n6128), .Z(n6168) );
  NAND U6719 ( .A(n38185), .B(n6060), .Z(n6062) );
  XOR U6720 ( .A(b[23]), .B(a[33]), .Z(n6207) );
  NAND U6721 ( .A(n38132), .B(n6207), .Z(n6061) );
  AND U6722 ( .A(n6062), .B(n6061), .Z(n6197) );
  NAND U6723 ( .A(n184), .B(n6063), .Z(n6065) );
  XOR U6724 ( .A(b[7]), .B(a[49]), .Z(n6210) );
  NAND U6725 ( .A(n36592), .B(n6210), .Z(n6064) );
  AND U6726 ( .A(n6065), .B(n6064), .Z(n6196) );
  NAND U6727 ( .A(n38289), .B(n6066), .Z(n6068) );
  XOR U6728 ( .A(b[25]), .B(a[31]), .Z(n6213) );
  NAND U6729 ( .A(n38247), .B(n6213), .Z(n6067) );
  NAND U6730 ( .A(n6068), .B(n6067), .Z(n6195) );
  XOR U6731 ( .A(n6196), .B(n6195), .Z(n6198) );
  XOR U6732 ( .A(n6197), .B(n6198), .Z(n6167) );
  XOR U6733 ( .A(n6168), .B(n6167), .Z(n6170) );
  NAND U6734 ( .A(n187), .B(n6069), .Z(n6071) );
  XOR U6735 ( .A(b[13]), .B(a[43]), .Z(n6216) );
  NAND U6736 ( .A(n37295), .B(n6216), .Z(n6070) );
  AND U6737 ( .A(n6071), .B(n6070), .Z(n6162) );
  NAND U6738 ( .A(n186), .B(n6072), .Z(n6074) );
  XOR U6739 ( .A(b[11]), .B(a[45]), .Z(n6219) );
  NAND U6740 ( .A(n37097), .B(n6219), .Z(n6073) );
  NAND U6741 ( .A(n6074), .B(n6073), .Z(n6161) );
  XNOR U6742 ( .A(n6162), .B(n6161), .Z(n6164) );
  NAND U6743 ( .A(n188), .B(n6075), .Z(n6077) );
  XOR U6744 ( .A(b[15]), .B(a[41]), .Z(n6222) );
  NAND U6745 ( .A(n37382), .B(n6222), .Z(n6076) );
  AND U6746 ( .A(n6077), .B(n6076), .Z(n6158) );
  NAND U6747 ( .A(n38064), .B(n6078), .Z(n6080) );
  XOR U6748 ( .A(b[21]), .B(a[35]), .Z(n6225) );
  NAND U6749 ( .A(n37993), .B(n6225), .Z(n6079) );
  AND U6750 ( .A(n6080), .B(n6079), .Z(n6156) );
  NAND U6751 ( .A(n185), .B(n6081), .Z(n6083) );
  XOR U6752 ( .A(b[9]), .B(a[47]), .Z(n6228) );
  NAND U6753 ( .A(n36805), .B(n6228), .Z(n6082) );
  NAND U6754 ( .A(n6083), .B(n6082), .Z(n6155) );
  XNOR U6755 ( .A(n6156), .B(n6155), .Z(n6157) );
  XNOR U6756 ( .A(n6158), .B(n6157), .Z(n6163) );
  XOR U6757 ( .A(n6164), .B(n6163), .Z(n6169) );
  XNOR U6758 ( .A(n6170), .B(n6169), .Z(n6181) );
  XNOR U6759 ( .A(n6182), .B(n6181), .Z(n6113) );
  XNOR U6760 ( .A(n6114), .B(n6113), .Z(n6115) );
  XOR U6761 ( .A(n6116), .B(n6115), .Z(n6232) );
  XNOR U6762 ( .A(n6231), .B(n6232), .Z(n6233) );
  XNOR U6763 ( .A(n6234), .B(n6233), .Z(n6109) );
  XOR U6764 ( .A(n6110), .B(n6109), .Z(n6102) );
  NANDN U6765 ( .A(n6085), .B(n6084), .Z(n6089) );
  NANDN U6766 ( .A(n6087), .B(n6086), .Z(n6088) );
  AND U6767 ( .A(n6089), .B(n6088), .Z(n6101) );
  XOR U6768 ( .A(n6102), .B(n6101), .Z(n6104) );
  XNOR U6769 ( .A(n6103), .B(n6104), .Z(n6095) );
  XNOR U6770 ( .A(n6096), .B(n6095), .Z(n6097) );
  XNOR U6771 ( .A(n6098), .B(n6097), .Z(n6237) );
  XNOR U6772 ( .A(sreg[279]), .B(n6237), .Z(n6239) );
  NANDN U6773 ( .A(sreg[278]), .B(n6090), .Z(n6094) );
  NAND U6774 ( .A(n6092), .B(n6091), .Z(n6093) );
  NAND U6775 ( .A(n6094), .B(n6093), .Z(n6238) );
  XNOR U6776 ( .A(n6239), .B(n6238), .Z(c[279]) );
  NANDN U6777 ( .A(n6096), .B(n6095), .Z(n6100) );
  NANDN U6778 ( .A(n6098), .B(n6097), .Z(n6099) );
  AND U6779 ( .A(n6100), .B(n6099), .Z(n6245) );
  NANDN U6780 ( .A(n6102), .B(n6101), .Z(n6106) );
  NANDN U6781 ( .A(n6104), .B(n6103), .Z(n6105) );
  AND U6782 ( .A(n6106), .B(n6105), .Z(n6243) );
  NANDN U6783 ( .A(n6108), .B(n6107), .Z(n6112) );
  NAND U6784 ( .A(n6110), .B(n6109), .Z(n6111) );
  AND U6785 ( .A(n6112), .B(n6111), .Z(n6250) );
  NANDN U6786 ( .A(n6114), .B(n6113), .Z(n6118) );
  NANDN U6787 ( .A(n6116), .B(n6115), .Z(n6117) );
  AND U6788 ( .A(n6118), .B(n6117), .Z(n6255) );
  NANDN U6789 ( .A(n6120), .B(n6119), .Z(n6124) );
  NAND U6790 ( .A(n6122), .B(n6121), .Z(n6123) );
  AND U6791 ( .A(n6124), .B(n6123), .Z(n6254) );
  XNOR U6792 ( .A(n6255), .B(n6254), .Z(n6257) );
  NANDN U6793 ( .A(n6126), .B(n6125), .Z(n6130) );
  NANDN U6794 ( .A(n6128), .B(n6127), .Z(n6129) );
  AND U6795 ( .A(n6130), .B(n6129), .Z(n6322) );
  NAND U6796 ( .A(n38385), .B(n6131), .Z(n6133) );
  XOR U6797 ( .A(b[27]), .B(a[30]), .Z(n6266) );
  NAND U6798 ( .A(n38343), .B(n6266), .Z(n6132) );
  AND U6799 ( .A(n6133), .B(n6132), .Z(n6329) );
  NAND U6800 ( .A(n183), .B(n6134), .Z(n6136) );
  XOR U6801 ( .A(b[5]), .B(a[52]), .Z(n6269) );
  NAND U6802 ( .A(n36296), .B(n6269), .Z(n6135) );
  AND U6803 ( .A(n6136), .B(n6135), .Z(n6327) );
  NAND U6804 ( .A(n190), .B(n6137), .Z(n6139) );
  XOR U6805 ( .A(b[19]), .B(a[38]), .Z(n6272) );
  NAND U6806 ( .A(n37821), .B(n6272), .Z(n6138) );
  NAND U6807 ( .A(n6139), .B(n6138), .Z(n6326) );
  XNOR U6808 ( .A(n6327), .B(n6326), .Z(n6328) );
  XNOR U6809 ( .A(n6329), .B(n6328), .Z(n6320) );
  NAND U6810 ( .A(n38470), .B(n6140), .Z(n6142) );
  XOR U6811 ( .A(b[31]), .B(a[26]), .Z(n6275) );
  NAND U6812 ( .A(n38453), .B(n6275), .Z(n6141) );
  AND U6813 ( .A(n6142), .B(n6141), .Z(n6287) );
  NAND U6814 ( .A(n181), .B(n6143), .Z(n6145) );
  XOR U6815 ( .A(b[3]), .B(a[54]), .Z(n6278) );
  NAND U6816 ( .A(n182), .B(n6278), .Z(n6144) );
  AND U6817 ( .A(n6145), .B(n6144), .Z(n6285) );
  NAND U6818 ( .A(n189), .B(n6146), .Z(n6148) );
  XOR U6819 ( .A(b[17]), .B(a[40]), .Z(n6281) );
  NAND U6820 ( .A(n37652), .B(n6281), .Z(n6147) );
  NAND U6821 ( .A(n6148), .B(n6147), .Z(n6284) );
  XNOR U6822 ( .A(n6285), .B(n6284), .Z(n6286) );
  XOR U6823 ( .A(n6287), .B(n6286), .Z(n6321) );
  XOR U6824 ( .A(n6320), .B(n6321), .Z(n6323) );
  XOR U6825 ( .A(n6322), .B(n6323), .Z(n6369) );
  NANDN U6826 ( .A(n6150), .B(n6149), .Z(n6154) );
  NANDN U6827 ( .A(n6152), .B(n6151), .Z(n6153) );
  AND U6828 ( .A(n6154), .B(n6153), .Z(n6308) );
  NANDN U6829 ( .A(n6156), .B(n6155), .Z(n6160) );
  NANDN U6830 ( .A(n6158), .B(n6157), .Z(n6159) );
  NAND U6831 ( .A(n6160), .B(n6159), .Z(n6309) );
  XNOR U6832 ( .A(n6308), .B(n6309), .Z(n6310) );
  NANDN U6833 ( .A(n6162), .B(n6161), .Z(n6166) );
  NAND U6834 ( .A(n6164), .B(n6163), .Z(n6165) );
  NAND U6835 ( .A(n6166), .B(n6165), .Z(n6311) );
  XNOR U6836 ( .A(n6310), .B(n6311), .Z(n6368) );
  XNOR U6837 ( .A(n6369), .B(n6368), .Z(n6371) );
  NAND U6838 ( .A(n6168), .B(n6167), .Z(n6172) );
  NAND U6839 ( .A(n6170), .B(n6169), .Z(n6171) );
  AND U6840 ( .A(n6172), .B(n6171), .Z(n6370) );
  XOR U6841 ( .A(n6371), .B(n6370), .Z(n6383) );
  NANDN U6842 ( .A(n6174), .B(n6173), .Z(n6178) );
  NANDN U6843 ( .A(n6176), .B(n6175), .Z(n6177) );
  AND U6844 ( .A(n6178), .B(n6177), .Z(n6380) );
  NANDN U6845 ( .A(n6184), .B(n6183), .Z(n6188) );
  OR U6846 ( .A(n6186), .B(n6185), .Z(n6187) );
  AND U6847 ( .A(n6188), .B(n6187), .Z(n6375) );
  NANDN U6848 ( .A(n6190), .B(n6189), .Z(n6194) );
  NANDN U6849 ( .A(n6192), .B(n6191), .Z(n6193) );
  AND U6850 ( .A(n6194), .B(n6193), .Z(n6315) );
  NANDN U6851 ( .A(n6196), .B(n6195), .Z(n6200) );
  OR U6852 ( .A(n6198), .B(n6197), .Z(n6199) );
  NAND U6853 ( .A(n6200), .B(n6199), .Z(n6314) );
  XNOR U6854 ( .A(n6315), .B(n6314), .Z(n6316) );
  NAND U6855 ( .A(n194), .B(n6201), .Z(n6203) );
  XOR U6856 ( .A(b[29]), .B(a[28]), .Z(n6341) );
  NAND U6857 ( .A(n38456), .B(n6341), .Z(n6202) );
  AND U6858 ( .A(n6203), .B(n6202), .Z(n6261) );
  AND U6859 ( .A(b[31]), .B(a[24]), .Z(n6260) );
  XNOR U6860 ( .A(n6261), .B(n6260), .Z(n6262) );
  NAND U6861 ( .A(b[0]), .B(a[56]), .Z(n6204) );
  XNOR U6862 ( .A(b[1]), .B(n6204), .Z(n6206) );
  NANDN U6863 ( .A(b[0]), .B(a[55]), .Z(n6205) );
  NAND U6864 ( .A(n6206), .B(n6205), .Z(n6263) );
  XNOR U6865 ( .A(n6262), .B(n6263), .Z(n6302) );
  NAND U6866 ( .A(n38185), .B(n6207), .Z(n6209) );
  XOR U6867 ( .A(b[23]), .B(a[34]), .Z(n6344) );
  NAND U6868 ( .A(n38132), .B(n6344), .Z(n6208) );
  AND U6869 ( .A(n6209), .B(n6208), .Z(n6335) );
  NAND U6870 ( .A(n184), .B(n6210), .Z(n6212) );
  XOR U6871 ( .A(b[7]), .B(a[50]), .Z(n6347) );
  NAND U6872 ( .A(n36592), .B(n6347), .Z(n6211) );
  AND U6873 ( .A(n6212), .B(n6211), .Z(n6333) );
  NAND U6874 ( .A(n38289), .B(n6213), .Z(n6215) );
  XOR U6875 ( .A(b[25]), .B(a[32]), .Z(n6350) );
  NAND U6876 ( .A(n38247), .B(n6350), .Z(n6214) );
  NAND U6877 ( .A(n6215), .B(n6214), .Z(n6332) );
  XNOR U6878 ( .A(n6333), .B(n6332), .Z(n6334) );
  XOR U6879 ( .A(n6335), .B(n6334), .Z(n6303) );
  XNOR U6880 ( .A(n6302), .B(n6303), .Z(n6304) );
  NAND U6881 ( .A(n187), .B(n6216), .Z(n6218) );
  XOR U6882 ( .A(b[13]), .B(a[44]), .Z(n6353) );
  NAND U6883 ( .A(n37295), .B(n6353), .Z(n6217) );
  AND U6884 ( .A(n6218), .B(n6217), .Z(n6297) );
  NAND U6885 ( .A(n186), .B(n6219), .Z(n6221) );
  XOR U6886 ( .A(b[11]), .B(a[46]), .Z(n6356) );
  NAND U6887 ( .A(n37097), .B(n6356), .Z(n6220) );
  NAND U6888 ( .A(n6221), .B(n6220), .Z(n6296) );
  XNOR U6889 ( .A(n6297), .B(n6296), .Z(n6298) );
  NAND U6890 ( .A(n188), .B(n6222), .Z(n6224) );
  XOR U6891 ( .A(b[15]), .B(a[42]), .Z(n6359) );
  NAND U6892 ( .A(n37382), .B(n6359), .Z(n6223) );
  AND U6893 ( .A(n6224), .B(n6223), .Z(n6293) );
  NAND U6894 ( .A(n38064), .B(n6225), .Z(n6227) );
  XOR U6895 ( .A(b[21]), .B(a[36]), .Z(n6362) );
  NAND U6896 ( .A(n37993), .B(n6362), .Z(n6226) );
  AND U6897 ( .A(n6227), .B(n6226), .Z(n6291) );
  NAND U6898 ( .A(n185), .B(n6228), .Z(n6230) );
  XOR U6899 ( .A(b[9]), .B(a[48]), .Z(n6365) );
  NAND U6900 ( .A(n36805), .B(n6365), .Z(n6229) );
  NAND U6901 ( .A(n6230), .B(n6229), .Z(n6290) );
  XNOR U6902 ( .A(n6291), .B(n6290), .Z(n6292) );
  XOR U6903 ( .A(n6293), .B(n6292), .Z(n6299) );
  XOR U6904 ( .A(n6298), .B(n6299), .Z(n6305) );
  XOR U6905 ( .A(n6304), .B(n6305), .Z(n6317) );
  XNOR U6906 ( .A(n6316), .B(n6317), .Z(n6374) );
  XNOR U6907 ( .A(n6375), .B(n6374), .Z(n6376) );
  XOR U6908 ( .A(n6377), .B(n6376), .Z(n6381) );
  XNOR U6909 ( .A(n6380), .B(n6381), .Z(n6382) );
  XNOR U6910 ( .A(n6383), .B(n6382), .Z(n6256) );
  XOR U6911 ( .A(n6257), .B(n6256), .Z(n6249) );
  NANDN U6912 ( .A(n6232), .B(n6231), .Z(n6236) );
  NANDN U6913 ( .A(n6234), .B(n6233), .Z(n6235) );
  AND U6914 ( .A(n6236), .B(n6235), .Z(n6248) );
  XOR U6915 ( .A(n6249), .B(n6248), .Z(n6251) );
  XNOR U6916 ( .A(n6250), .B(n6251), .Z(n6242) );
  XNOR U6917 ( .A(n6243), .B(n6242), .Z(n6244) );
  XNOR U6918 ( .A(n6245), .B(n6244), .Z(n6386) );
  XNOR U6919 ( .A(sreg[280]), .B(n6386), .Z(n6388) );
  NANDN U6920 ( .A(sreg[279]), .B(n6237), .Z(n6241) );
  NAND U6921 ( .A(n6239), .B(n6238), .Z(n6240) );
  NAND U6922 ( .A(n6241), .B(n6240), .Z(n6387) );
  XNOR U6923 ( .A(n6388), .B(n6387), .Z(c[280]) );
  NANDN U6924 ( .A(n6243), .B(n6242), .Z(n6247) );
  NANDN U6925 ( .A(n6245), .B(n6244), .Z(n6246) );
  AND U6926 ( .A(n6247), .B(n6246), .Z(n6394) );
  NANDN U6927 ( .A(n6249), .B(n6248), .Z(n6253) );
  NANDN U6928 ( .A(n6251), .B(n6250), .Z(n6252) );
  AND U6929 ( .A(n6253), .B(n6252), .Z(n6392) );
  NANDN U6930 ( .A(n6255), .B(n6254), .Z(n6259) );
  NAND U6931 ( .A(n6257), .B(n6256), .Z(n6258) );
  AND U6932 ( .A(n6259), .B(n6258), .Z(n6399) );
  NANDN U6933 ( .A(n6261), .B(n6260), .Z(n6265) );
  NANDN U6934 ( .A(n6263), .B(n6262), .Z(n6264) );
  AND U6935 ( .A(n6265), .B(n6264), .Z(n6483) );
  NAND U6936 ( .A(n38385), .B(n6266), .Z(n6268) );
  XOR U6937 ( .A(b[27]), .B(a[31]), .Z(n6427) );
  NAND U6938 ( .A(n38343), .B(n6427), .Z(n6267) );
  AND U6939 ( .A(n6268), .B(n6267), .Z(n6490) );
  NAND U6940 ( .A(n183), .B(n6269), .Z(n6271) );
  XOR U6941 ( .A(b[5]), .B(a[53]), .Z(n6430) );
  NAND U6942 ( .A(n36296), .B(n6430), .Z(n6270) );
  AND U6943 ( .A(n6271), .B(n6270), .Z(n6488) );
  NAND U6944 ( .A(n190), .B(n6272), .Z(n6274) );
  XOR U6945 ( .A(b[19]), .B(a[39]), .Z(n6433) );
  NAND U6946 ( .A(n37821), .B(n6433), .Z(n6273) );
  NAND U6947 ( .A(n6274), .B(n6273), .Z(n6487) );
  XNOR U6948 ( .A(n6488), .B(n6487), .Z(n6489) );
  XNOR U6949 ( .A(n6490), .B(n6489), .Z(n6481) );
  NAND U6950 ( .A(n38470), .B(n6275), .Z(n6277) );
  XOR U6951 ( .A(b[31]), .B(a[27]), .Z(n6436) );
  NAND U6952 ( .A(n38453), .B(n6436), .Z(n6276) );
  AND U6953 ( .A(n6277), .B(n6276), .Z(n6448) );
  NAND U6954 ( .A(n181), .B(n6278), .Z(n6280) );
  XOR U6955 ( .A(b[3]), .B(a[55]), .Z(n6439) );
  NAND U6956 ( .A(n182), .B(n6439), .Z(n6279) );
  AND U6957 ( .A(n6280), .B(n6279), .Z(n6446) );
  NAND U6958 ( .A(n189), .B(n6281), .Z(n6283) );
  XOR U6959 ( .A(b[17]), .B(a[41]), .Z(n6442) );
  NAND U6960 ( .A(n37652), .B(n6442), .Z(n6282) );
  NAND U6961 ( .A(n6283), .B(n6282), .Z(n6445) );
  XNOR U6962 ( .A(n6446), .B(n6445), .Z(n6447) );
  XOR U6963 ( .A(n6448), .B(n6447), .Z(n6482) );
  XOR U6964 ( .A(n6481), .B(n6482), .Z(n6484) );
  XOR U6965 ( .A(n6483), .B(n6484), .Z(n6416) );
  NANDN U6966 ( .A(n6285), .B(n6284), .Z(n6289) );
  NANDN U6967 ( .A(n6287), .B(n6286), .Z(n6288) );
  AND U6968 ( .A(n6289), .B(n6288), .Z(n6469) );
  NANDN U6969 ( .A(n6291), .B(n6290), .Z(n6295) );
  NANDN U6970 ( .A(n6293), .B(n6292), .Z(n6294) );
  NAND U6971 ( .A(n6295), .B(n6294), .Z(n6470) );
  XNOR U6972 ( .A(n6469), .B(n6470), .Z(n6471) );
  NANDN U6973 ( .A(n6297), .B(n6296), .Z(n6301) );
  NANDN U6974 ( .A(n6299), .B(n6298), .Z(n6300) );
  NAND U6975 ( .A(n6301), .B(n6300), .Z(n6472) );
  XNOR U6976 ( .A(n6471), .B(n6472), .Z(n6415) );
  XNOR U6977 ( .A(n6416), .B(n6415), .Z(n6418) );
  NANDN U6978 ( .A(n6303), .B(n6302), .Z(n6307) );
  NANDN U6979 ( .A(n6305), .B(n6304), .Z(n6306) );
  AND U6980 ( .A(n6307), .B(n6306), .Z(n6417) );
  XOR U6981 ( .A(n6418), .B(n6417), .Z(n6531) );
  NANDN U6982 ( .A(n6309), .B(n6308), .Z(n6313) );
  NANDN U6983 ( .A(n6311), .B(n6310), .Z(n6312) );
  AND U6984 ( .A(n6313), .B(n6312), .Z(n6529) );
  NANDN U6985 ( .A(n6315), .B(n6314), .Z(n6319) );
  NANDN U6986 ( .A(n6317), .B(n6316), .Z(n6318) );
  AND U6987 ( .A(n6319), .B(n6318), .Z(n6412) );
  NANDN U6988 ( .A(n6321), .B(n6320), .Z(n6325) );
  OR U6989 ( .A(n6323), .B(n6322), .Z(n6324) );
  AND U6990 ( .A(n6325), .B(n6324), .Z(n6410) );
  NANDN U6991 ( .A(n6327), .B(n6326), .Z(n6331) );
  NANDN U6992 ( .A(n6329), .B(n6328), .Z(n6330) );
  AND U6993 ( .A(n6331), .B(n6330), .Z(n6476) );
  NANDN U6994 ( .A(n6333), .B(n6332), .Z(n6337) );
  NANDN U6995 ( .A(n6335), .B(n6334), .Z(n6336) );
  NAND U6996 ( .A(n6337), .B(n6336), .Z(n6475) );
  XNOR U6997 ( .A(n6476), .B(n6475), .Z(n6477) );
  NAND U6998 ( .A(b[0]), .B(a[57]), .Z(n6338) );
  XNOR U6999 ( .A(b[1]), .B(n6338), .Z(n6340) );
  NANDN U7000 ( .A(b[0]), .B(a[56]), .Z(n6339) );
  NAND U7001 ( .A(n6340), .B(n6339), .Z(n6424) );
  NAND U7002 ( .A(n194), .B(n6341), .Z(n6343) );
  XOR U7003 ( .A(b[29]), .B(a[29]), .Z(n6502) );
  NAND U7004 ( .A(n38456), .B(n6502), .Z(n6342) );
  AND U7005 ( .A(n6343), .B(n6342), .Z(n6422) );
  AND U7006 ( .A(b[31]), .B(a[25]), .Z(n6421) );
  XNOR U7007 ( .A(n6422), .B(n6421), .Z(n6423) );
  XNOR U7008 ( .A(n6424), .B(n6423), .Z(n6463) );
  NAND U7009 ( .A(n38185), .B(n6344), .Z(n6346) );
  XOR U7010 ( .A(b[23]), .B(a[35]), .Z(n6505) );
  NAND U7011 ( .A(n38132), .B(n6505), .Z(n6345) );
  AND U7012 ( .A(n6346), .B(n6345), .Z(n6496) );
  NAND U7013 ( .A(n184), .B(n6347), .Z(n6349) );
  XOR U7014 ( .A(b[7]), .B(a[51]), .Z(n6508) );
  NAND U7015 ( .A(n36592), .B(n6508), .Z(n6348) );
  AND U7016 ( .A(n6349), .B(n6348), .Z(n6494) );
  NAND U7017 ( .A(n38289), .B(n6350), .Z(n6352) );
  XOR U7018 ( .A(b[25]), .B(a[33]), .Z(n6511) );
  NAND U7019 ( .A(n38247), .B(n6511), .Z(n6351) );
  NAND U7020 ( .A(n6352), .B(n6351), .Z(n6493) );
  XNOR U7021 ( .A(n6494), .B(n6493), .Z(n6495) );
  XOR U7022 ( .A(n6496), .B(n6495), .Z(n6464) );
  XNOR U7023 ( .A(n6463), .B(n6464), .Z(n6465) );
  NAND U7024 ( .A(n187), .B(n6353), .Z(n6355) );
  XOR U7025 ( .A(b[13]), .B(a[45]), .Z(n6514) );
  NAND U7026 ( .A(n37295), .B(n6514), .Z(n6354) );
  AND U7027 ( .A(n6355), .B(n6354), .Z(n6458) );
  NAND U7028 ( .A(n186), .B(n6356), .Z(n6358) );
  XOR U7029 ( .A(b[11]), .B(a[47]), .Z(n6517) );
  NAND U7030 ( .A(n37097), .B(n6517), .Z(n6357) );
  NAND U7031 ( .A(n6358), .B(n6357), .Z(n6457) );
  XNOR U7032 ( .A(n6458), .B(n6457), .Z(n6459) );
  NAND U7033 ( .A(n188), .B(n6359), .Z(n6361) );
  XOR U7034 ( .A(b[15]), .B(a[43]), .Z(n6520) );
  NAND U7035 ( .A(n37382), .B(n6520), .Z(n6360) );
  AND U7036 ( .A(n6361), .B(n6360), .Z(n6454) );
  NAND U7037 ( .A(n38064), .B(n6362), .Z(n6364) );
  XOR U7038 ( .A(b[21]), .B(a[37]), .Z(n6523) );
  NAND U7039 ( .A(n37993), .B(n6523), .Z(n6363) );
  AND U7040 ( .A(n6364), .B(n6363), .Z(n6452) );
  NAND U7041 ( .A(n185), .B(n6365), .Z(n6367) );
  XOR U7042 ( .A(b[9]), .B(a[49]), .Z(n6526) );
  NAND U7043 ( .A(n36805), .B(n6526), .Z(n6366) );
  NAND U7044 ( .A(n6367), .B(n6366), .Z(n6451) );
  XNOR U7045 ( .A(n6452), .B(n6451), .Z(n6453) );
  XOR U7046 ( .A(n6454), .B(n6453), .Z(n6460) );
  XOR U7047 ( .A(n6459), .B(n6460), .Z(n6466) );
  XOR U7048 ( .A(n6465), .B(n6466), .Z(n6478) );
  XNOR U7049 ( .A(n6477), .B(n6478), .Z(n6409) );
  XNOR U7050 ( .A(n6410), .B(n6409), .Z(n6411) );
  XOR U7051 ( .A(n6412), .B(n6411), .Z(n6530) );
  XOR U7052 ( .A(n6529), .B(n6530), .Z(n6532) );
  XOR U7053 ( .A(n6531), .B(n6532), .Z(n6406) );
  NANDN U7054 ( .A(n6369), .B(n6368), .Z(n6373) );
  NAND U7055 ( .A(n6371), .B(n6370), .Z(n6372) );
  AND U7056 ( .A(n6373), .B(n6372), .Z(n6404) );
  NANDN U7057 ( .A(n6375), .B(n6374), .Z(n6379) );
  NANDN U7058 ( .A(n6377), .B(n6376), .Z(n6378) );
  AND U7059 ( .A(n6379), .B(n6378), .Z(n6403) );
  XNOR U7060 ( .A(n6404), .B(n6403), .Z(n6405) );
  XNOR U7061 ( .A(n6406), .B(n6405), .Z(n6397) );
  NANDN U7062 ( .A(n6381), .B(n6380), .Z(n6385) );
  NANDN U7063 ( .A(n6383), .B(n6382), .Z(n6384) );
  NAND U7064 ( .A(n6385), .B(n6384), .Z(n6398) );
  XOR U7065 ( .A(n6397), .B(n6398), .Z(n6400) );
  XNOR U7066 ( .A(n6399), .B(n6400), .Z(n6391) );
  XNOR U7067 ( .A(n6392), .B(n6391), .Z(n6393) );
  XNOR U7068 ( .A(n6394), .B(n6393), .Z(n6535) );
  XNOR U7069 ( .A(sreg[281]), .B(n6535), .Z(n6537) );
  NANDN U7070 ( .A(sreg[280]), .B(n6386), .Z(n6390) );
  NAND U7071 ( .A(n6388), .B(n6387), .Z(n6389) );
  NAND U7072 ( .A(n6390), .B(n6389), .Z(n6536) );
  XNOR U7073 ( .A(n6537), .B(n6536), .Z(c[281]) );
  NANDN U7074 ( .A(n6392), .B(n6391), .Z(n6396) );
  NANDN U7075 ( .A(n6394), .B(n6393), .Z(n6395) );
  AND U7076 ( .A(n6396), .B(n6395), .Z(n6543) );
  NANDN U7077 ( .A(n6398), .B(n6397), .Z(n6402) );
  NANDN U7078 ( .A(n6400), .B(n6399), .Z(n6401) );
  AND U7079 ( .A(n6402), .B(n6401), .Z(n6541) );
  NANDN U7080 ( .A(n6404), .B(n6403), .Z(n6408) );
  NANDN U7081 ( .A(n6406), .B(n6405), .Z(n6407) );
  AND U7082 ( .A(n6408), .B(n6407), .Z(n6549) );
  NANDN U7083 ( .A(n6410), .B(n6409), .Z(n6414) );
  NANDN U7084 ( .A(n6412), .B(n6411), .Z(n6413) );
  AND U7085 ( .A(n6414), .B(n6413), .Z(n6553) );
  NANDN U7086 ( .A(n6416), .B(n6415), .Z(n6420) );
  NAND U7087 ( .A(n6418), .B(n6417), .Z(n6419) );
  AND U7088 ( .A(n6420), .B(n6419), .Z(n6552) );
  XNOR U7089 ( .A(n6553), .B(n6552), .Z(n6555) );
  NANDN U7090 ( .A(n6422), .B(n6421), .Z(n6426) );
  NANDN U7091 ( .A(n6424), .B(n6423), .Z(n6425) );
  AND U7092 ( .A(n6426), .B(n6425), .Z(n6632) );
  NAND U7093 ( .A(n38385), .B(n6427), .Z(n6429) );
  XOR U7094 ( .A(b[27]), .B(a[32]), .Z(n6576) );
  NAND U7095 ( .A(n38343), .B(n6576), .Z(n6428) );
  AND U7096 ( .A(n6429), .B(n6428), .Z(n6639) );
  NAND U7097 ( .A(n183), .B(n6430), .Z(n6432) );
  XOR U7098 ( .A(b[5]), .B(a[54]), .Z(n6579) );
  NAND U7099 ( .A(n36296), .B(n6579), .Z(n6431) );
  AND U7100 ( .A(n6432), .B(n6431), .Z(n6637) );
  NAND U7101 ( .A(n190), .B(n6433), .Z(n6435) );
  XOR U7102 ( .A(b[19]), .B(a[40]), .Z(n6582) );
  NAND U7103 ( .A(n37821), .B(n6582), .Z(n6434) );
  NAND U7104 ( .A(n6435), .B(n6434), .Z(n6636) );
  XNOR U7105 ( .A(n6637), .B(n6636), .Z(n6638) );
  XNOR U7106 ( .A(n6639), .B(n6638), .Z(n6630) );
  NAND U7107 ( .A(n38470), .B(n6436), .Z(n6438) );
  XOR U7108 ( .A(b[31]), .B(a[28]), .Z(n6585) );
  NAND U7109 ( .A(n38453), .B(n6585), .Z(n6437) );
  AND U7110 ( .A(n6438), .B(n6437), .Z(n6597) );
  NAND U7111 ( .A(n181), .B(n6439), .Z(n6441) );
  XOR U7112 ( .A(b[3]), .B(a[56]), .Z(n6588) );
  NAND U7113 ( .A(n182), .B(n6588), .Z(n6440) );
  AND U7114 ( .A(n6441), .B(n6440), .Z(n6595) );
  NAND U7115 ( .A(n189), .B(n6442), .Z(n6444) );
  XOR U7116 ( .A(b[17]), .B(a[42]), .Z(n6591) );
  NAND U7117 ( .A(n37652), .B(n6591), .Z(n6443) );
  NAND U7118 ( .A(n6444), .B(n6443), .Z(n6594) );
  XNOR U7119 ( .A(n6595), .B(n6594), .Z(n6596) );
  XOR U7120 ( .A(n6597), .B(n6596), .Z(n6631) );
  XOR U7121 ( .A(n6630), .B(n6631), .Z(n6633) );
  XOR U7122 ( .A(n6632), .B(n6633), .Z(n6565) );
  NANDN U7123 ( .A(n6446), .B(n6445), .Z(n6450) );
  NANDN U7124 ( .A(n6448), .B(n6447), .Z(n6449) );
  AND U7125 ( .A(n6450), .B(n6449), .Z(n6618) );
  NANDN U7126 ( .A(n6452), .B(n6451), .Z(n6456) );
  NANDN U7127 ( .A(n6454), .B(n6453), .Z(n6455) );
  NAND U7128 ( .A(n6456), .B(n6455), .Z(n6619) );
  XNOR U7129 ( .A(n6618), .B(n6619), .Z(n6620) );
  NANDN U7130 ( .A(n6458), .B(n6457), .Z(n6462) );
  NANDN U7131 ( .A(n6460), .B(n6459), .Z(n6461) );
  NAND U7132 ( .A(n6462), .B(n6461), .Z(n6621) );
  XNOR U7133 ( .A(n6620), .B(n6621), .Z(n6564) );
  XNOR U7134 ( .A(n6565), .B(n6564), .Z(n6567) );
  NANDN U7135 ( .A(n6464), .B(n6463), .Z(n6468) );
  NANDN U7136 ( .A(n6466), .B(n6465), .Z(n6467) );
  AND U7137 ( .A(n6468), .B(n6467), .Z(n6566) );
  XOR U7138 ( .A(n6567), .B(n6566), .Z(n6681) );
  NANDN U7139 ( .A(n6470), .B(n6469), .Z(n6474) );
  NANDN U7140 ( .A(n6472), .B(n6471), .Z(n6473) );
  AND U7141 ( .A(n6474), .B(n6473), .Z(n6678) );
  NANDN U7142 ( .A(n6476), .B(n6475), .Z(n6480) );
  NANDN U7143 ( .A(n6478), .B(n6477), .Z(n6479) );
  AND U7144 ( .A(n6480), .B(n6479), .Z(n6561) );
  NANDN U7145 ( .A(n6482), .B(n6481), .Z(n6486) );
  OR U7146 ( .A(n6484), .B(n6483), .Z(n6485) );
  AND U7147 ( .A(n6486), .B(n6485), .Z(n6559) );
  NANDN U7148 ( .A(n6488), .B(n6487), .Z(n6492) );
  NANDN U7149 ( .A(n6490), .B(n6489), .Z(n6491) );
  AND U7150 ( .A(n6492), .B(n6491), .Z(n6625) );
  NANDN U7151 ( .A(n6494), .B(n6493), .Z(n6498) );
  NANDN U7152 ( .A(n6496), .B(n6495), .Z(n6497) );
  NAND U7153 ( .A(n6498), .B(n6497), .Z(n6624) );
  XNOR U7154 ( .A(n6625), .B(n6624), .Z(n6626) );
  NAND U7155 ( .A(b[0]), .B(a[58]), .Z(n6499) );
  XNOR U7156 ( .A(b[1]), .B(n6499), .Z(n6501) );
  NANDN U7157 ( .A(b[0]), .B(a[57]), .Z(n6500) );
  NAND U7158 ( .A(n6501), .B(n6500), .Z(n6573) );
  NAND U7159 ( .A(n194), .B(n6502), .Z(n6504) );
  XOR U7160 ( .A(b[29]), .B(a[30]), .Z(n6651) );
  NAND U7161 ( .A(n38456), .B(n6651), .Z(n6503) );
  AND U7162 ( .A(n6504), .B(n6503), .Z(n6571) );
  AND U7163 ( .A(b[31]), .B(a[26]), .Z(n6570) );
  XNOR U7164 ( .A(n6571), .B(n6570), .Z(n6572) );
  XNOR U7165 ( .A(n6573), .B(n6572), .Z(n6612) );
  NAND U7166 ( .A(n38185), .B(n6505), .Z(n6507) );
  XOR U7167 ( .A(b[23]), .B(a[36]), .Z(n6654) );
  NAND U7168 ( .A(n38132), .B(n6654), .Z(n6506) );
  AND U7169 ( .A(n6507), .B(n6506), .Z(n6645) );
  NAND U7170 ( .A(n184), .B(n6508), .Z(n6510) );
  XOR U7171 ( .A(b[7]), .B(a[52]), .Z(n6657) );
  NAND U7172 ( .A(n36592), .B(n6657), .Z(n6509) );
  AND U7173 ( .A(n6510), .B(n6509), .Z(n6643) );
  NAND U7174 ( .A(n38289), .B(n6511), .Z(n6513) );
  XOR U7175 ( .A(b[25]), .B(a[34]), .Z(n6660) );
  NAND U7176 ( .A(n38247), .B(n6660), .Z(n6512) );
  NAND U7177 ( .A(n6513), .B(n6512), .Z(n6642) );
  XNOR U7178 ( .A(n6643), .B(n6642), .Z(n6644) );
  XOR U7179 ( .A(n6645), .B(n6644), .Z(n6613) );
  XNOR U7180 ( .A(n6612), .B(n6613), .Z(n6614) );
  NAND U7181 ( .A(n187), .B(n6514), .Z(n6516) );
  XOR U7182 ( .A(b[13]), .B(a[46]), .Z(n6663) );
  NAND U7183 ( .A(n37295), .B(n6663), .Z(n6515) );
  AND U7184 ( .A(n6516), .B(n6515), .Z(n6607) );
  NAND U7185 ( .A(n186), .B(n6517), .Z(n6519) );
  XOR U7186 ( .A(b[11]), .B(a[48]), .Z(n6666) );
  NAND U7187 ( .A(n37097), .B(n6666), .Z(n6518) );
  NAND U7188 ( .A(n6519), .B(n6518), .Z(n6606) );
  XNOR U7189 ( .A(n6607), .B(n6606), .Z(n6608) );
  NAND U7190 ( .A(n188), .B(n6520), .Z(n6522) );
  XOR U7191 ( .A(b[15]), .B(a[44]), .Z(n6669) );
  NAND U7192 ( .A(n37382), .B(n6669), .Z(n6521) );
  AND U7193 ( .A(n6522), .B(n6521), .Z(n6603) );
  NAND U7194 ( .A(n38064), .B(n6523), .Z(n6525) );
  XOR U7195 ( .A(b[21]), .B(a[38]), .Z(n6672) );
  NAND U7196 ( .A(n37993), .B(n6672), .Z(n6524) );
  AND U7197 ( .A(n6525), .B(n6524), .Z(n6601) );
  NAND U7198 ( .A(n185), .B(n6526), .Z(n6528) );
  XOR U7199 ( .A(b[9]), .B(a[50]), .Z(n6675) );
  NAND U7200 ( .A(n36805), .B(n6675), .Z(n6527) );
  NAND U7201 ( .A(n6528), .B(n6527), .Z(n6600) );
  XNOR U7202 ( .A(n6601), .B(n6600), .Z(n6602) );
  XOR U7203 ( .A(n6603), .B(n6602), .Z(n6609) );
  XOR U7204 ( .A(n6608), .B(n6609), .Z(n6615) );
  XOR U7205 ( .A(n6614), .B(n6615), .Z(n6627) );
  XNOR U7206 ( .A(n6626), .B(n6627), .Z(n6558) );
  XNOR U7207 ( .A(n6559), .B(n6558), .Z(n6560) );
  XOR U7208 ( .A(n6561), .B(n6560), .Z(n6679) );
  XNOR U7209 ( .A(n6678), .B(n6679), .Z(n6680) );
  XNOR U7210 ( .A(n6681), .B(n6680), .Z(n6554) );
  XOR U7211 ( .A(n6555), .B(n6554), .Z(n6547) );
  NANDN U7212 ( .A(n6530), .B(n6529), .Z(n6534) );
  OR U7213 ( .A(n6532), .B(n6531), .Z(n6533) );
  AND U7214 ( .A(n6534), .B(n6533), .Z(n6546) );
  XNOR U7215 ( .A(n6547), .B(n6546), .Z(n6548) );
  XNOR U7216 ( .A(n6549), .B(n6548), .Z(n6540) );
  XNOR U7217 ( .A(n6541), .B(n6540), .Z(n6542) );
  XNOR U7218 ( .A(n6543), .B(n6542), .Z(n6684) );
  XNOR U7219 ( .A(sreg[282]), .B(n6684), .Z(n6686) );
  NANDN U7220 ( .A(sreg[281]), .B(n6535), .Z(n6539) );
  NAND U7221 ( .A(n6537), .B(n6536), .Z(n6538) );
  NAND U7222 ( .A(n6539), .B(n6538), .Z(n6685) );
  XNOR U7223 ( .A(n6686), .B(n6685), .Z(c[282]) );
  NANDN U7224 ( .A(n6541), .B(n6540), .Z(n6545) );
  NANDN U7225 ( .A(n6543), .B(n6542), .Z(n6544) );
  AND U7226 ( .A(n6545), .B(n6544), .Z(n6692) );
  NANDN U7227 ( .A(n6547), .B(n6546), .Z(n6551) );
  NANDN U7228 ( .A(n6549), .B(n6548), .Z(n6550) );
  AND U7229 ( .A(n6551), .B(n6550), .Z(n6690) );
  NANDN U7230 ( .A(n6553), .B(n6552), .Z(n6557) );
  NAND U7231 ( .A(n6555), .B(n6554), .Z(n6556) );
  AND U7232 ( .A(n6557), .B(n6556), .Z(n6697) );
  NANDN U7233 ( .A(n6559), .B(n6558), .Z(n6563) );
  NANDN U7234 ( .A(n6561), .B(n6560), .Z(n6562) );
  AND U7235 ( .A(n6563), .B(n6562), .Z(n6702) );
  NANDN U7236 ( .A(n6565), .B(n6564), .Z(n6569) );
  NAND U7237 ( .A(n6567), .B(n6566), .Z(n6568) );
  AND U7238 ( .A(n6569), .B(n6568), .Z(n6701) );
  XNOR U7239 ( .A(n6702), .B(n6701), .Z(n6704) );
  NANDN U7240 ( .A(n6571), .B(n6570), .Z(n6575) );
  NANDN U7241 ( .A(n6573), .B(n6572), .Z(n6574) );
  AND U7242 ( .A(n6575), .B(n6574), .Z(n6781) );
  NAND U7243 ( .A(n38385), .B(n6576), .Z(n6578) );
  XOR U7244 ( .A(b[27]), .B(a[33]), .Z(n6725) );
  NAND U7245 ( .A(n38343), .B(n6725), .Z(n6577) );
  AND U7246 ( .A(n6578), .B(n6577), .Z(n6788) );
  NAND U7247 ( .A(n183), .B(n6579), .Z(n6581) );
  XOR U7248 ( .A(b[5]), .B(a[55]), .Z(n6728) );
  NAND U7249 ( .A(n36296), .B(n6728), .Z(n6580) );
  AND U7250 ( .A(n6581), .B(n6580), .Z(n6786) );
  NAND U7251 ( .A(n190), .B(n6582), .Z(n6584) );
  XOR U7252 ( .A(b[19]), .B(a[41]), .Z(n6731) );
  NAND U7253 ( .A(n37821), .B(n6731), .Z(n6583) );
  NAND U7254 ( .A(n6584), .B(n6583), .Z(n6785) );
  XNOR U7255 ( .A(n6786), .B(n6785), .Z(n6787) );
  XNOR U7256 ( .A(n6788), .B(n6787), .Z(n6779) );
  NAND U7257 ( .A(n38470), .B(n6585), .Z(n6587) );
  XOR U7258 ( .A(b[31]), .B(a[29]), .Z(n6734) );
  NAND U7259 ( .A(n38453), .B(n6734), .Z(n6586) );
  AND U7260 ( .A(n6587), .B(n6586), .Z(n6746) );
  NAND U7261 ( .A(n181), .B(n6588), .Z(n6590) );
  XOR U7262 ( .A(b[3]), .B(a[57]), .Z(n6737) );
  NAND U7263 ( .A(n182), .B(n6737), .Z(n6589) );
  AND U7264 ( .A(n6590), .B(n6589), .Z(n6744) );
  NAND U7265 ( .A(n189), .B(n6591), .Z(n6593) );
  XOR U7266 ( .A(b[17]), .B(a[43]), .Z(n6740) );
  NAND U7267 ( .A(n37652), .B(n6740), .Z(n6592) );
  NAND U7268 ( .A(n6593), .B(n6592), .Z(n6743) );
  XNOR U7269 ( .A(n6744), .B(n6743), .Z(n6745) );
  XOR U7270 ( .A(n6746), .B(n6745), .Z(n6780) );
  XOR U7271 ( .A(n6779), .B(n6780), .Z(n6782) );
  XOR U7272 ( .A(n6781), .B(n6782), .Z(n6714) );
  NANDN U7273 ( .A(n6595), .B(n6594), .Z(n6599) );
  NANDN U7274 ( .A(n6597), .B(n6596), .Z(n6598) );
  AND U7275 ( .A(n6599), .B(n6598), .Z(n6767) );
  NANDN U7276 ( .A(n6601), .B(n6600), .Z(n6605) );
  NANDN U7277 ( .A(n6603), .B(n6602), .Z(n6604) );
  NAND U7278 ( .A(n6605), .B(n6604), .Z(n6768) );
  XNOR U7279 ( .A(n6767), .B(n6768), .Z(n6769) );
  NANDN U7280 ( .A(n6607), .B(n6606), .Z(n6611) );
  NANDN U7281 ( .A(n6609), .B(n6608), .Z(n6610) );
  NAND U7282 ( .A(n6611), .B(n6610), .Z(n6770) );
  XNOR U7283 ( .A(n6769), .B(n6770), .Z(n6713) );
  XNOR U7284 ( .A(n6714), .B(n6713), .Z(n6716) );
  NANDN U7285 ( .A(n6613), .B(n6612), .Z(n6617) );
  NANDN U7286 ( .A(n6615), .B(n6614), .Z(n6616) );
  AND U7287 ( .A(n6617), .B(n6616), .Z(n6715) );
  XOR U7288 ( .A(n6716), .B(n6715), .Z(n6830) );
  NANDN U7289 ( .A(n6619), .B(n6618), .Z(n6623) );
  NANDN U7290 ( .A(n6621), .B(n6620), .Z(n6622) );
  AND U7291 ( .A(n6623), .B(n6622), .Z(n6827) );
  NANDN U7292 ( .A(n6625), .B(n6624), .Z(n6629) );
  NANDN U7293 ( .A(n6627), .B(n6626), .Z(n6628) );
  AND U7294 ( .A(n6629), .B(n6628), .Z(n6710) );
  NANDN U7295 ( .A(n6631), .B(n6630), .Z(n6635) );
  OR U7296 ( .A(n6633), .B(n6632), .Z(n6634) );
  AND U7297 ( .A(n6635), .B(n6634), .Z(n6708) );
  NANDN U7298 ( .A(n6637), .B(n6636), .Z(n6641) );
  NANDN U7299 ( .A(n6639), .B(n6638), .Z(n6640) );
  AND U7300 ( .A(n6641), .B(n6640), .Z(n6774) );
  NANDN U7301 ( .A(n6643), .B(n6642), .Z(n6647) );
  NANDN U7302 ( .A(n6645), .B(n6644), .Z(n6646) );
  NAND U7303 ( .A(n6647), .B(n6646), .Z(n6773) );
  XNOR U7304 ( .A(n6774), .B(n6773), .Z(n6775) );
  NAND U7305 ( .A(b[0]), .B(a[59]), .Z(n6648) );
  XNOR U7306 ( .A(b[1]), .B(n6648), .Z(n6650) );
  NANDN U7307 ( .A(b[0]), .B(a[58]), .Z(n6649) );
  NAND U7308 ( .A(n6650), .B(n6649), .Z(n6722) );
  NAND U7309 ( .A(n194), .B(n6651), .Z(n6653) );
  XOR U7310 ( .A(b[29]), .B(a[31]), .Z(n6800) );
  NAND U7311 ( .A(n38456), .B(n6800), .Z(n6652) );
  AND U7312 ( .A(n6653), .B(n6652), .Z(n6720) );
  AND U7313 ( .A(b[31]), .B(a[27]), .Z(n6719) );
  XNOR U7314 ( .A(n6720), .B(n6719), .Z(n6721) );
  XNOR U7315 ( .A(n6722), .B(n6721), .Z(n6761) );
  NAND U7316 ( .A(n38185), .B(n6654), .Z(n6656) );
  XOR U7317 ( .A(b[23]), .B(a[37]), .Z(n6803) );
  NAND U7318 ( .A(n38132), .B(n6803), .Z(n6655) );
  AND U7319 ( .A(n6656), .B(n6655), .Z(n6794) );
  NAND U7320 ( .A(n184), .B(n6657), .Z(n6659) );
  XOR U7321 ( .A(b[7]), .B(a[53]), .Z(n6806) );
  NAND U7322 ( .A(n36592), .B(n6806), .Z(n6658) );
  AND U7323 ( .A(n6659), .B(n6658), .Z(n6792) );
  NAND U7324 ( .A(n38289), .B(n6660), .Z(n6662) );
  XOR U7325 ( .A(b[25]), .B(a[35]), .Z(n6809) );
  NAND U7326 ( .A(n38247), .B(n6809), .Z(n6661) );
  NAND U7327 ( .A(n6662), .B(n6661), .Z(n6791) );
  XNOR U7328 ( .A(n6792), .B(n6791), .Z(n6793) );
  XOR U7329 ( .A(n6794), .B(n6793), .Z(n6762) );
  XNOR U7330 ( .A(n6761), .B(n6762), .Z(n6763) );
  NAND U7331 ( .A(n187), .B(n6663), .Z(n6665) );
  XOR U7332 ( .A(b[13]), .B(a[47]), .Z(n6812) );
  NAND U7333 ( .A(n37295), .B(n6812), .Z(n6664) );
  AND U7334 ( .A(n6665), .B(n6664), .Z(n6756) );
  NAND U7335 ( .A(n186), .B(n6666), .Z(n6668) );
  XOR U7336 ( .A(b[11]), .B(a[49]), .Z(n6815) );
  NAND U7337 ( .A(n37097), .B(n6815), .Z(n6667) );
  NAND U7338 ( .A(n6668), .B(n6667), .Z(n6755) );
  XNOR U7339 ( .A(n6756), .B(n6755), .Z(n6757) );
  NAND U7340 ( .A(n188), .B(n6669), .Z(n6671) );
  XOR U7341 ( .A(b[15]), .B(a[45]), .Z(n6818) );
  NAND U7342 ( .A(n37382), .B(n6818), .Z(n6670) );
  AND U7343 ( .A(n6671), .B(n6670), .Z(n6752) );
  NAND U7344 ( .A(n38064), .B(n6672), .Z(n6674) );
  XOR U7345 ( .A(b[21]), .B(a[39]), .Z(n6821) );
  NAND U7346 ( .A(n37993), .B(n6821), .Z(n6673) );
  AND U7347 ( .A(n6674), .B(n6673), .Z(n6750) );
  NAND U7348 ( .A(n185), .B(n6675), .Z(n6677) );
  XOR U7349 ( .A(b[9]), .B(a[51]), .Z(n6824) );
  NAND U7350 ( .A(n36805), .B(n6824), .Z(n6676) );
  NAND U7351 ( .A(n6677), .B(n6676), .Z(n6749) );
  XNOR U7352 ( .A(n6750), .B(n6749), .Z(n6751) );
  XOR U7353 ( .A(n6752), .B(n6751), .Z(n6758) );
  XOR U7354 ( .A(n6757), .B(n6758), .Z(n6764) );
  XOR U7355 ( .A(n6763), .B(n6764), .Z(n6776) );
  XNOR U7356 ( .A(n6775), .B(n6776), .Z(n6707) );
  XNOR U7357 ( .A(n6708), .B(n6707), .Z(n6709) );
  XOR U7358 ( .A(n6710), .B(n6709), .Z(n6828) );
  XNOR U7359 ( .A(n6827), .B(n6828), .Z(n6829) );
  XNOR U7360 ( .A(n6830), .B(n6829), .Z(n6703) );
  XOR U7361 ( .A(n6704), .B(n6703), .Z(n6696) );
  NANDN U7362 ( .A(n6679), .B(n6678), .Z(n6683) );
  NANDN U7363 ( .A(n6681), .B(n6680), .Z(n6682) );
  AND U7364 ( .A(n6683), .B(n6682), .Z(n6695) );
  XOR U7365 ( .A(n6696), .B(n6695), .Z(n6698) );
  XNOR U7366 ( .A(n6697), .B(n6698), .Z(n6689) );
  XNOR U7367 ( .A(n6690), .B(n6689), .Z(n6691) );
  XNOR U7368 ( .A(n6692), .B(n6691), .Z(n6833) );
  XNOR U7369 ( .A(sreg[283]), .B(n6833), .Z(n6835) );
  NANDN U7370 ( .A(sreg[282]), .B(n6684), .Z(n6688) );
  NAND U7371 ( .A(n6686), .B(n6685), .Z(n6687) );
  NAND U7372 ( .A(n6688), .B(n6687), .Z(n6834) );
  XNOR U7373 ( .A(n6835), .B(n6834), .Z(c[283]) );
  NANDN U7374 ( .A(n6690), .B(n6689), .Z(n6694) );
  NANDN U7375 ( .A(n6692), .B(n6691), .Z(n6693) );
  AND U7376 ( .A(n6694), .B(n6693), .Z(n6841) );
  NANDN U7377 ( .A(n6696), .B(n6695), .Z(n6700) );
  NANDN U7378 ( .A(n6698), .B(n6697), .Z(n6699) );
  AND U7379 ( .A(n6700), .B(n6699), .Z(n6839) );
  NANDN U7380 ( .A(n6702), .B(n6701), .Z(n6706) );
  NAND U7381 ( .A(n6704), .B(n6703), .Z(n6705) );
  AND U7382 ( .A(n6706), .B(n6705), .Z(n6846) );
  NANDN U7383 ( .A(n6708), .B(n6707), .Z(n6712) );
  NANDN U7384 ( .A(n6710), .B(n6709), .Z(n6711) );
  AND U7385 ( .A(n6712), .B(n6711), .Z(n6975) );
  NANDN U7386 ( .A(n6714), .B(n6713), .Z(n6718) );
  NAND U7387 ( .A(n6716), .B(n6715), .Z(n6717) );
  AND U7388 ( .A(n6718), .B(n6717), .Z(n6974) );
  XNOR U7389 ( .A(n6975), .B(n6974), .Z(n6977) );
  NANDN U7390 ( .A(n6720), .B(n6719), .Z(n6724) );
  NANDN U7391 ( .A(n6722), .B(n6721), .Z(n6723) );
  AND U7392 ( .A(n6724), .B(n6723), .Z(n6922) );
  NAND U7393 ( .A(n38385), .B(n6725), .Z(n6727) );
  XOR U7394 ( .A(b[27]), .B(a[34]), .Z(n6868) );
  NAND U7395 ( .A(n38343), .B(n6868), .Z(n6726) );
  AND U7396 ( .A(n6727), .B(n6726), .Z(n6929) );
  NAND U7397 ( .A(n183), .B(n6728), .Z(n6730) );
  XOR U7398 ( .A(b[5]), .B(a[56]), .Z(n6871) );
  NAND U7399 ( .A(n36296), .B(n6871), .Z(n6729) );
  AND U7400 ( .A(n6730), .B(n6729), .Z(n6927) );
  NAND U7401 ( .A(n190), .B(n6731), .Z(n6733) );
  XOR U7402 ( .A(b[19]), .B(a[42]), .Z(n6874) );
  NAND U7403 ( .A(n37821), .B(n6874), .Z(n6732) );
  NAND U7404 ( .A(n6733), .B(n6732), .Z(n6926) );
  XNOR U7405 ( .A(n6927), .B(n6926), .Z(n6928) );
  XNOR U7406 ( .A(n6929), .B(n6928), .Z(n6920) );
  NAND U7407 ( .A(n38470), .B(n6734), .Z(n6736) );
  XOR U7408 ( .A(b[31]), .B(a[30]), .Z(n6877) );
  NAND U7409 ( .A(n38453), .B(n6877), .Z(n6735) );
  AND U7410 ( .A(n6736), .B(n6735), .Z(n6889) );
  NAND U7411 ( .A(n181), .B(n6737), .Z(n6739) );
  XOR U7412 ( .A(b[3]), .B(a[58]), .Z(n6880) );
  NAND U7413 ( .A(n182), .B(n6880), .Z(n6738) );
  AND U7414 ( .A(n6739), .B(n6738), .Z(n6887) );
  NAND U7415 ( .A(n189), .B(n6740), .Z(n6742) );
  XOR U7416 ( .A(b[17]), .B(a[44]), .Z(n6883) );
  NAND U7417 ( .A(n37652), .B(n6883), .Z(n6741) );
  NAND U7418 ( .A(n6742), .B(n6741), .Z(n6886) );
  XNOR U7419 ( .A(n6887), .B(n6886), .Z(n6888) );
  XOR U7420 ( .A(n6889), .B(n6888), .Z(n6921) );
  XOR U7421 ( .A(n6920), .B(n6921), .Z(n6923) );
  XOR U7422 ( .A(n6922), .B(n6923), .Z(n6857) );
  NANDN U7423 ( .A(n6744), .B(n6743), .Z(n6748) );
  NANDN U7424 ( .A(n6746), .B(n6745), .Z(n6747) );
  AND U7425 ( .A(n6748), .B(n6747), .Z(n6910) );
  NANDN U7426 ( .A(n6750), .B(n6749), .Z(n6754) );
  NANDN U7427 ( .A(n6752), .B(n6751), .Z(n6753) );
  NAND U7428 ( .A(n6754), .B(n6753), .Z(n6911) );
  XNOR U7429 ( .A(n6910), .B(n6911), .Z(n6912) );
  NANDN U7430 ( .A(n6756), .B(n6755), .Z(n6760) );
  NANDN U7431 ( .A(n6758), .B(n6757), .Z(n6759) );
  NAND U7432 ( .A(n6760), .B(n6759), .Z(n6913) );
  XNOR U7433 ( .A(n6912), .B(n6913), .Z(n6856) );
  XNOR U7434 ( .A(n6857), .B(n6856), .Z(n6859) );
  NANDN U7435 ( .A(n6762), .B(n6761), .Z(n6766) );
  NANDN U7436 ( .A(n6764), .B(n6763), .Z(n6765) );
  AND U7437 ( .A(n6766), .B(n6765), .Z(n6858) );
  XOR U7438 ( .A(n6859), .B(n6858), .Z(n6971) );
  NANDN U7439 ( .A(n6768), .B(n6767), .Z(n6772) );
  NANDN U7440 ( .A(n6770), .B(n6769), .Z(n6771) );
  AND U7441 ( .A(n6772), .B(n6771), .Z(n6968) );
  NANDN U7442 ( .A(n6774), .B(n6773), .Z(n6778) );
  NANDN U7443 ( .A(n6776), .B(n6775), .Z(n6777) );
  AND U7444 ( .A(n6778), .B(n6777), .Z(n6853) );
  NANDN U7445 ( .A(n6780), .B(n6779), .Z(n6784) );
  OR U7446 ( .A(n6782), .B(n6781), .Z(n6783) );
  AND U7447 ( .A(n6784), .B(n6783), .Z(n6851) );
  NANDN U7448 ( .A(n6786), .B(n6785), .Z(n6790) );
  NANDN U7449 ( .A(n6788), .B(n6787), .Z(n6789) );
  AND U7450 ( .A(n6790), .B(n6789), .Z(n6917) );
  NANDN U7451 ( .A(n6792), .B(n6791), .Z(n6796) );
  NANDN U7452 ( .A(n6794), .B(n6793), .Z(n6795) );
  NAND U7453 ( .A(n6796), .B(n6795), .Z(n6916) );
  XNOR U7454 ( .A(n6917), .B(n6916), .Z(n6919) );
  NAND U7455 ( .A(b[0]), .B(a[60]), .Z(n6797) );
  XNOR U7456 ( .A(b[1]), .B(n6797), .Z(n6799) );
  NANDN U7457 ( .A(b[0]), .B(a[59]), .Z(n6798) );
  NAND U7458 ( .A(n6799), .B(n6798), .Z(n6865) );
  NAND U7459 ( .A(n194), .B(n6800), .Z(n6802) );
  XOR U7460 ( .A(b[29]), .B(a[32]), .Z(n6941) );
  NAND U7461 ( .A(n38456), .B(n6941), .Z(n6801) );
  AND U7462 ( .A(n6802), .B(n6801), .Z(n6863) );
  AND U7463 ( .A(b[31]), .B(a[28]), .Z(n6862) );
  XNOR U7464 ( .A(n6863), .B(n6862), .Z(n6864) );
  XNOR U7465 ( .A(n6865), .B(n6864), .Z(n6905) );
  NAND U7466 ( .A(n38185), .B(n6803), .Z(n6805) );
  XOR U7467 ( .A(b[23]), .B(a[38]), .Z(n6944) );
  NAND U7468 ( .A(n38132), .B(n6944), .Z(n6804) );
  AND U7469 ( .A(n6805), .B(n6804), .Z(n6934) );
  NAND U7470 ( .A(n184), .B(n6806), .Z(n6808) );
  XOR U7471 ( .A(b[7]), .B(a[54]), .Z(n6947) );
  NAND U7472 ( .A(n36592), .B(n6947), .Z(n6807) );
  AND U7473 ( .A(n6808), .B(n6807), .Z(n6933) );
  NAND U7474 ( .A(n38289), .B(n6809), .Z(n6811) );
  XOR U7475 ( .A(b[25]), .B(a[36]), .Z(n6950) );
  NAND U7476 ( .A(n38247), .B(n6950), .Z(n6810) );
  NAND U7477 ( .A(n6811), .B(n6810), .Z(n6932) );
  XOR U7478 ( .A(n6933), .B(n6932), .Z(n6935) );
  XOR U7479 ( .A(n6934), .B(n6935), .Z(n6904) );
  XOR U7480 ( .A(n6905), .B(n6904), .Z(n6907) );
  NAND U7481 ( .A(n187), .B(n6812), .Z(n6814) );
  XOR U7482 ( .A(b[13]), .B(a[48]), .Z(n6953) );
  NAND U7483 ( .A(n37295), .B(n6953), .Z(n6813) );
  AND U7484 ( .A(n6814), .B(n6813), .Z(n6899) );
  NAND U7485 ( .A(n186), .B(n6815), .Z(n6817) );
  XOR U7486 ( .A(b[11]), .B(a[50]), .Z(n6956) );
  NAND U7487 ( .A(n37097), .B(n6956), .Z(n6816) );
  NAND U7488 ( .A(n6817), .B(n6816), .Z(n6898) );
  XNOR U7489 ( .A(n6899), .B(n6898), .Z(n6901) );
  NAND U7490 ( .A(n188), .B(n6818), .Z(n6820) );
  XOR U7491 ( .A(b[15]), .B(a[46]), .Z(n6959) );
  NAND U7492 ( .A(n37382), .B(n6959), .Z(n6819) );
  AND U7493 ( .A(n6820), .B(n6819), .Z(n6895) );
  NAND U7494 ( .A(n38064), .B(n6821), .Z(n6823) );
  XOR U7495 ( .A(b[21]), .B(a[40]), .Z(n6962) );
  NAND U7496 ( .A(n37993), .B(n6962), .Z(n6822) );
  AND U7497 ( .A(n6823), .B(n6822), .Z(n6893) );
  NAND U7498 ( .A(n185), .B(n6824), .Z(n6826) );
  XOR U7499 ( .A(b[9]), .B(a[52]), .Z(n6965) );
  NAND U7500 ( .A(n36805), .B(n6965), .Z(n6825) );
  NAND U7501 ( .A(n6826), .B(n6825), .Z(n6892) );
  XNOR U7502 ( .A(n6893), .B(n6892), .Z(n6894) );
  XNOR U7503 ( .A(n6895), .B(n6894), .Z(n6900) );
  XOR U7504 ( .A(n6901), .B(n6900), .Z(n6906) );
  XNOR U7505 ( .A(n6907), .B(n6906), .Z(n6918) );
  XNOR U7506 ( .A(n6919), .B(n6918), .Z(n6850) );
  XNOR U7507 ( .A(n6851), .B(n6850), .Z(n6852) );
  XOR U7508 ( .A(n6853), .B(n6852), .Z(n6969) );
  XNOR U7509 ( .A(n6968), .B(n6969), .Z(n6970) );
  XNOR U7510 ( .A(n6971), .B(n6970), .Z(n6976) );
  XOR U7511 ( .A(n6977), .B(n6976), .Z(n6845) );
  NANDN U7512 ( .A(n6828), .B(n6827), .Z(n6832) );
  NANDN U7513 ( .A(n6830), .B(n6829), .Z(n6831) );
  AND U7514 ( .A(n6832), .B(n6831), .Z(n6844) );
  XOR U7515 ( .A(n6845), .B(n6844), .Z(n6847) );
  XNOR U7516 ( .A(n6846), .B(n6847), .Z(n6838) );
  XNOR U7517 ( .A(n6839), .B(n6838), .Z(n6840) );
  XNOR U7518 ( .A(n6841), .B(n6840), .Z(n6980) );
  XNOR U7519 ( .A(sreg[284]), .B(n6980), .Z(n6982) );
  NANDN U7520 ( .A(sreg[283]), .B(n6833), .Z(n6837) );
  NAND U7521 ( .A(n6835), .B(n6834), .Z(n6836) );
  NAND U7522 ( .A(n6837), .B(n6836), .Z(n6981) );
  XNOR U7523 ( .A(n6982), .B(n6981), .Z(c[284]) );
  NANDN U7524 ( .A(n6839), .B(n6838), .Z(n6843) );
  NANDN U7525 ( .A(n6841), .B(n6840), .Z(n6842) );
  AND U7526 ( .A(n6843), .B(n6842), .Z(n6988) );
  NANDN U7527 ( .A(n6845), .B(n6844), .Z(n6849) );
  NANDN U7528 ( .A(n6847), .B(n6846), .Z(n6848) );
  AND U7529 ( .A(n6849), .B(n6848), .Z(n6986) );
  NANDN U7530 ( .A(n6851), .B(n6850), .Z(n6855) );
  NANDN U7531 ( .A(n6853), .B(n6852), .Z(n6854) );
  AND U7532 ( .A(n6855), .B(n6854), .Z(n7124) );
  NANDN U7533 ( .A(n6857), .B(n6856), .Z(n6861) );
  NAND U7534 ( .A(n6859), .B(n6858), .Z(n6860) );
  AND U7535 ( .A(n6861), .B(n6860), .Z(n7123) );
  XNOR U7536 ( .A(n7124), .B(n7123), .Z(n7126) );
  NANDN U7537 ( .A(n6863), .B(n6862), .Z(n6867) );
  NANDN U7538 ( .A(n6865), .B(n6864), .Z(n6866) );
  AND U7539 ( .A(n6867), .B(n6866), .Z(n7059) );
  NAND U7540 ( .A(n38385), .B(n6868), .Z(n6870) );
  XOR U7541 ( .A(b[27]), .B(a[35]), .Z(n7003) );
  NAND U7542 ( .A(n38343), .B(n7003), .Z(n6869) );
  AND U7543 ( .A(n6870), .B(n6869), .Z(n7066) );
  NAND U7544 ( .A(n183), .B(n6871), .Z(n6873) );
  XOR U7545 ( .A(b[5]), .B(a[57]), .Z(n7006) );
  NAND U7546 ( .A(n36296), .B(n7006), .Z(n6872) );
  AND U7547 ( .A(n6873), .B(n6872), .Z(n7064) );
  NAND U7548 ( .A(n190), .B(n6874), .Z(n6876) );
  XOR U7549 ( .A(b[19]), .B(a[43]), .Z(n7009) );
  NAND U7550 ( .A(n37821), .B(n7009), .Z(n6875) );
  NAND U7551 ( .A(n6876), .B(n6875), .Z(n7063) );
  XNOR U7552 ( .A(n7064), .B(n7063), .Z(n7065) );
  XNOR U7553 ( .A(n7066), .B(n7065), .Z(n7057) );
  NAND U7554 ( .A(n38470), .B(n6877), .Z(n6879) );
  XOR U7555 ( .A(b[31]), .B(a[31]), .Z(n7012) );
  NAND U7556 ( .A(n38453), .B(n7012), .Z(n6878) );
  AND U7557 ( .A(n6879), .B(n6878), .Z(n7024) );
  NAND U7558 ( .A(n181), .B(n6880), .Z(n6882) );
  XOR U7559 ( .A(b[3]), .B(a[59]), .Z(n7015) );
  NAND U7560 ( .A(n182), .B(n7015), .Z(n6881) );
  AND U7561 ( .A(n6882), .B(n6881), .Z(n7022) );
  NAND U7562 ( .A(n189), .B(n6883), .Z(n6885) );
  XOR U7563 ( .A(b[17]), .B(a[45]), .Z(n7018) );
  NAND U7564 ( .A(n37652), .B(n7018), .Z(n6884) );
  NAND U7565 ( .A(n6885), .B(n6884), .Z(n7021) );
  XNOR U7566 ( .A(n7022), .B(n7021), .Z(n7023) );
  XOR U7567 ( .A(n7024), .B(n7023), .Z(n7058) );
  XOR U7568 ( .A(n7057), .B(n7058), .Z(n7060) );
  XOR U7569 ( .A(n7059), .B(n7060), .Z(n7106) );
  NANDN U7570 ( .A(n6887), .B(n6886), .Z(n6891) );
  NANDN U7571 ( .A(n6889), .B(n6888), .Z(n6890) );
  AND U7572 ( .A(n6891), .B(n6890), .Z(n7045) );
  NANDN U7573 ( .A(n6893), .B(n6892), .Z(n6897) );
  NANDN U7574 ( .A(n6895), .B(n6894), .Z(n6896) );
  NAND U7575 ( .A(n6897), .B(n6896), .Z(n7046) );
  XNOR U7576 ( .A(n7045), .B(n7046), .Z(n7047) );
  NANDN U7577 ( .A(n6899), .B(n6898), .Z(n6903) );
  NAND U7578 ( .A(n6901), .B(n6900), .Z(n6902) );
  NAND U7579 ( .A(n6903), .B(n6902), .Z(n7048) );
  XNOR U7580 ( .A(n7047), .B(n7048), .Z(n7105) );
  XNOR U7581 ( .A(n7106), .B(n7105), .Z(n7108) );
  NAND U7582 ( .A(n6905), .B(n6904), .Z(n6909) );
  NAND U7583 ( .A(n6907), .B(n6906), .Z(n6908) );
  AND U7584 ( .A(n6909), .B(n6908), .Z(n7107) );
  XOR U7585 ( .A(n7108), .B(n7107), .Z(n7120) );
  NANDN U7586 ( .A(n6911), .B(n6910), .Z(n6915) );
  NANDN U7587 ( .A(n6913), .B(n6912), .Z(n6914) );
  AND U7588 ( .A(n6915), .B(n6914), .Z(n7117) );
  NANDN U7589 ( .A(n6921), .B(n6920), .Z(n6925) );
  OR U7590 ( .A(n6923), .B(n6922), .Z(n6924) );
  AND U7591 ( .A(n6925), .B(n6924), .Z(n7112) );
  NANDN U7592 ( .A(n6927), .B(n6926), .Z(n6931) );
  NANDN U7593 ( .A(n6929), .B(n6928), .Z(n6930) );
  AND U7594 ( .A(n6931), .B(n6930), .Z(n7052) );
  NANDN U7595 ( .A(n6933), .B(n6932), .Z(n6937) );
  OR U7596 ( .A(n6935), .B(n6934), .Z(n6936) );
  NAND U7597 ( .A(n6937), .B(n6936), .Z(n7051) );
  XNOR U7598 ( .A(n7052), .B(n7051), .Z(n7053) );
  NAND U7599 ( .A(b[0]), .B(a[61]), .Z(n6938) );
  XNOR U7600 ( .A(b[1]), .B(n6938), .Z(n6940) );
  NANDN U7601 ( .A(b[0]), .B(a[60]), .Z(n6939) );
  NAND U7602 ( .A(n6940), .B(n6939), .Z(n7000) );
  NAND U7603 ( .A(n194), .B(n6941), .Z(n6943) );
  XOR U7604 ( .A(b[29]), .B(a[33]), .Z(n7078) );
  NAND U7605 ( .A(n38456), .B(n7078), .Z(n6942) );
  AND U7606 ( .A(n6943), .B(n6942), .Z(n6998) );
  AND U7607 ( .A(b[31]), .B(a[29]), .Z(n6997) );
  XNOR U7608 ( .A(n6998), .B(n6997), .Z(n6999) );
  XNOR U7609 ( .A(n7000), .B(n6999), .Z(n7039) );
  NAND U7610 ( .A(n38185), .B(n6944), .Z(n6946) );
  XOR U7611 ( .A(b[23]), .B(a[39]), .Z(n7081) );
  NAND U7612 ( .A(n38132), .B(n7081), .Z(n6945) );
  AND U7613 ( .A(n6946), .B(n6945), .Z(n7072) );
  NAND U7614 ( .A(n184), .B(n6947), .Z(n6949) );
  XOR U7615 ( .A(b[7]), .B(a[55]), .Z(n7084) );
  NAND U7616 ( .A(n36592), .B(n7084), .Z(n6948) );
  AND U7617 ( .A(n6949), .B(n6948), .Z(n7070) );
  NAND U7618 ( .A(n38289), .B(n6950), .Z(n6952) );
  XOR U7619 ( .A(b[25]), .B(a[37]), .Z(n7087) );
  NAND U7620 ( .A(n38247), .B(n7087), .Z(n6951) );
  NAND U7621 ( .A(n6952), .B(n6951), .Z(n7069) );
  XNOR U7622 ( .A(n7070), .B(n7069), .Z(n7071) );
  XOR U7623 ( .A(n7072), .B(n7071), .Z(n7040) );
  XNOR U7624 ( .A(n7039), .B(n7040), .Z(n7041) );
  NAND U7625 ( .A(n187), .B(n6953), .Z(n6955) );
  XOR U7626 ( .A(b[13]), .B(a[49]), .Z(n7090) );
  NAND U7627 ( .A(n37295), .B(n7090), .Z(n6954) );
  AND U7628 ( .A(n6955), .B(n6954), .Z(n7034) );
  NAND U7629 ( .A(n186), .B(n6956), .Z(n6958) );
  XOR U7630 ( .A(b[11]), .B(a[51]), .Z(n7093) );
  NAND U7631 ( .A(n37097), .B(n7093), .Z(n6957) );
  NAND U7632 ( .A(n6958), .B(n6957), .Z(n7033) );
  XNOR U7633 ( .A(n7034), .B(n7033), .Z(n7035) );
  NAND U7634 ( .A(n188), .B(n6959), .Z(n6961) );
  XOR U7635 ( .A(b[15]), .B(a[47]), .Z(n7096) );
  NAND U7636 ( .A(n37382), .B(n7096), .Z(n6960) );
  AND U7637 ( .A(n6961), .B(n6960), .Z(n7030) );
  NAND U7638 ( .A(n38064), .B(n6962), .Z(n6964) );
  XOR U7639 ( .A(b[21]), .B(a[41]), .Z(n7099) );
  NAND U7640 ( .A(n37993), .B(n7099), .Z(n6963) );
  AND U7641 ( .A(n6964), .B(n6963), .Z(n7028) );
  NAND U7642 ( .A(n185), .B(n6965), .Z(n6967) );
  XOR U7643 ( .A(b[9]), .B(a[53]), .Z(n7102) );
  NAND U7644 ( .A(n36805), .B(n7102), .Z(n6966) );
  NAND U7645 ( .A(n6967), .B(n6966), .Z(n7027) );
  XNOR U7646 ( .A(n7028), .B(n7027), .Z(n7029) );
  XOR U7647 ( .A(n7030), .B(n7029), .Z(n7036) );
  XOR U7648 ( .A(n7035), .B(n7036), .Z(n7042) );
  XOR U7649 ( .A(n7041), .B(n7042), .Z(n7054) );
  XNOR U7650 ( .A(n7053), .B(n7054), .Z(n7111) );
  XNOR U7651 ( .A(n7112), .B(n7111), .Z(n7113) );
  XOR U7652 ( .A(n7114), .B(n7113), .Z(n7118) );
  XNOR U7653 ( .A(n7117), .B(n7118), .Z(n7119) );
  XNOR U7654 ( .A(n7120), .B(n7119), .Z(n7125) );
  XOR U7655 ( .A(n7126), .B(n7125), .Z(n6992) );
  NANDN U7656 ( .A(n6969), .B(n6968), .Z(n6973) );
  NANDN U7657 ( .A(n6971), .B(n6970), .Z(n6972) );
  AND U7658 ( .A(n6973), .B(n6972), .Z(n6991) );
  XNOR U7659 ( .A(n6992), .B(n6991), .Z(n6993) );
  NANDN U7660 ( .A(n6975), .B(n6974), .Z(n6979) );
  NAND U7661 ( .A(n6977), .B(n6976), .Z(n6978) );
  NAND U7662 ( .A(n6979), .B(n6978), .Z(n6994) );
  XNOR U7663 ( .A(n6993), .B(n6994), .Z(n6985) );
  XNOR U7664 ( .A(n6986), .B(n6985), .Z(n6987) );
  XNOR U7665 ( .A(n6988), .B(n6987), .Z(n7129) );
  XNOR U7666 ( .A(sreg[285]), .B(n7129), .Z(n7131) );
  NANDN U7667 ( .A(sreg[284]), .B(n6980), .Z(n6984) );
  NAND U7668 ( .A(n6982), .B(n6981), .Z(n6983) );
  NAND U7669 ( .A(n6984), .B(n6983), .Z(n7130) );
  XNOR U7670 ( .A(n7131), .B(n7130), .Z(c[285]) );
  NANDN U7671 ( .A(n6986), .B(n6985), .Z(n6990) );
  NANDN U7672 ( .A(n6988), .B(n6987), .Z(n6989) );
  AND U7673 ( .A(n6990), .B(n6989), .Z(n7137) );
  NANDN U7674 ( .A(n6992), .B(n6991), .Z(n6996) );
  NANDN U7675 ( .A(n6994), .B(n6993), .Z(n6995) );
  AND U7676 ( .A(n6996), .B(n6995), .Z(n7135) );
  NANDN U7677 ( .A(n6998), .B(n6997), .Z(n7002) );
  NANDN U7678 ( .A(n7000), .B(n6999), .Z(n7001) );
  AND U7679 ( .A(n7002), .B(n7001), .Z(n7226) );
  NAND U7680 ( .A(n38385), .B(n7003), .Z(n7005) );
  XOR U7681 ( .A(b[27]), .B(a[36]), .Z(n7170) );
  NAND U7682 ( .A(n38343), .B(n7170), .Z(n7004) );
  AND U7683 ( .A(n7005), .B(n7004), .Z(n7233) );
  NAND U7684 ( .A(n183), .B(n7006), .Z(n7008) );
  XOR U7685 ( .A(b[5]), .B(a[58]), .Z(n7173) );
  NAND U7686 ( .A(n36296), .B(n7173), .Z(n7007) );
  AND U7687 ( .A(n7008), .B(n7007), .Z(n7231) );
  NAND U7688 ( .A(n190), .B(n7009), .Z(n7011) );
  XOR U7689 ( .A(b[19]), .B(a[44]), .Z(n7176) );
  NAND U7690 ( .A(n37821), .B(n7176), .Z(n7010) );
  NAND U7691 ( .A(n7011), .B(n7010), .Z(n7230) );
  XNOR U7692 ( .A(n7231), .B(n7230), .Z(n7232) );
  XNOR U7693 ( .A(n7233), .B(n7232), .Z(n7224) );
  NAND U7694 ( .A(n38470), .B(n7012), .Z(n7014) );
  XOR U7695 ( .A(b[31]), .B(a[32]), .Z(n7179) );
  NAND U7696 ( .A(n38453), .B(n7179), .Z(n7013) );
  AND U7697 ( .A(n7014), .B(n7013), .Z(n7191) );
  NAND U7698 ( .A(n181), .B(n7015), .Z(n7017) );
  XOR U7699 ( .A(b[3]), .B(a[60]), .Z(n7182) );
  NAND U7700 ( .A(n182), .B(n7182), .Z(n7016) );
  AND U7701 ( .A(n7017), .B(n7016), .Z(n7189) );
  NAND U7702 ( .A(n189), .B(n7018), .Z(n7020) );
  XOR U7703 ( .A(b[17]), .B(a[46]), .Z(n7185) );
  NAND U7704 ( .A(n37652), .B(n7185), .Z(n7019) );
  NAND U7705 ( .A(n7020), .B(n7019), .Z(n7188) );
  XNOR U7706 ( .A(n7189), .B(n7188), .Z(n7190) );
  XOR U7707 ( .A(n7191), .B(n7190), .Z(n7225) );
  XOR U7708 ( .A(n7224), .B(n7225), .Z(n7227) );
  XOR U7709 ( .A(n7226), .B(n7227), .Z(n7159) );
  NANDN U7710 ( .A(n7022), .B(n7021), .Z(n7026) );
  NANDN U7711 ( .A(n7024), .B(n7023), .Z(n7025) );
  AND U7712 ( .A(n7026), .B(n7025), .Z(n7212) );
  NANDN U7713 ( .A(n7028), .B(n7027), .Z(n7032) );
  NANDN U7714 ( .A(n7030), .B(n7029), .Z(n7031) );
  NAND U7715 ( .A(n7032), .B(n7031), .Z(n7213) );
  XNOR U7716 ( .A(n7212), .B(n7213), .Z(n7214) );
  NANDN U7717 ( .A(n7034), .B(n7033), .Z(n7038) );
  NANDN U7718 ( .A(n7036), .B(n7035), .Z(n7037) );
  NAND U7719 ( .A(n7038), .B(n7037), .Z(n7215) );
  XNOR U7720 ( .A(n7214), .B(n7215), .Z(n7158) );
  XNOR U7721 ( .A(n7159), .B(n7158), .Z(n7161) );
  NANDN U7722 ( .A(n7040), .B(n7039), .Z(n7044) );
  NANDN U7723 ( .A(n7042), .B(n7041), .Z(n7043) );
  AND U7724 ( .A(n7044), .B(n7043), .Z(n7160) );
  XOR U7725 ( .A(n7161), .B(n7160), .Z(n7274) );
  NANDN U7726 ( .A(n7046), .B(n7045), .Z(n7050) );
  NANDN U7727 ( .A(n7048), .B(n7047), .Z(n7049) );
  AND U7728 ( .A(n7050), .B(n7049), .Z(n7272) );
  NANDN U7729 ( .A(n7052), .B(n7051), .Z(n7056) );
  NANDN U7730 ( .A(n7054), .B(n7053), .Z(n7055) );
  AND U7731 ( .A(n7056), .B(n7055), .Z(n7155) );
  NANDN U7732 ( .A(n7058), .B(n7057), .Z(n7062) );
  OR U7733 ( .A(n7060), .B(n7059), .Z(n7061) );
  AND U7734 ( .A(n7062), .B(n7061), .Z(n7153) );
  NANDN U7735 ( .A(n7064), .B(n7063), .Z(n7068) );
  NANDN U7736 ( .A(n7066), .B(n7065), .Z(n7067) );
  AND U7737 ( .A(n7068), .B(n7067), .Z(n7219) );
  NANDN U7738 ( .A(n7070), .B(n7069), .Z(n7074) );
  NANDN U7739 ( .A(n7072), .B(n7071), .Z(n7073) );
  NAND U7740 ( .A(n7074), .B(n7073), .Z(n7218) );
  XNOR U7741 ( .A(n7219), .B(n7218), .Z(n7220) );
  NAND U7742 ( .A(b[0]), .B(a[62]), .Z(n7075) );
  XNOR U7743 ( .A(b[1]), .B(n7075), .Z(n7077) );
  NANDN U7744 ( .A(b[0]), .B(a[61]), .Z(n7076) );
  NAND U7745 ( .A(n7077), .B(n7076), .Z(n7167) );
  NAND U7746 ( .A(n194), .B(n7078), .Z(n7080) );
  XOR U7747 ( .A(b[29]), .B(a[34]), .Z(n7245) );
  NAND U7748 ( .A(n38456), .B(n7245), .Z(n7079) );
  AND U7749 ( .A(n7080), .B(n7079), .Z(n7165) );
  AND U7750 ( .A(b[31]), .B(a[30]), .Z(n7164) );
  XNOR U7751 ( .A(n7165), .B(n7164), .Z(n7166) );
  XNOR U7752 ( .A(n7167), .B(n7166), .Z(n7206) );
  NAND U7753 ( .A(n38185), .B(n7081), .Z(n7083) );
  XOR U7754 ( .A(b[23]), .B(a[40]), .Z(n7248) );
  NAND U7755 ( .A(n38132), .B(n7248), .Z(n7082) );
  AND U7756 ( .A(n7083), .B(n7082), .Z(n7239) );
  NAND U7757 ( .A(n184), .B(n7084), .Z(n7086) );
  XOR U7758 ( .A(b[7]), .B(a[56]), .Z(n7251) );
  NAND U7759 ( .A(n36592), .B(n7251), .Z(n7085) );
  AND U7760 ( .A(n7086), .B(n7085), .Z(n7237) );
  NAND U7761 ( .A(n38289), .B(n7087), .Z(n7089) );
  XOR U7762 ( .A(b[25]), .B(a[38]), .Z(n7254) );
  NAND U7763 ( .A(n38247), .B(n7254), .Z(n7088) );
  NAND U7764 ( .A(n7089), .B(n7088), .Z(n7236) );
  XNOR U7765 ( .A(n7237), .B(n7236), .Z(n7238) );
  XOR U7766 ( .A(n7239), .B(n7238), .Z(n7207) );
  XNOR U7767 ( .A(n7206), .B(n7207), .Z(n7208) );
  NAND U7768 ( .A(n187), .B(n7090), .Z(n7092) );
  XOR U7769 ( .A(b[13]), .B(a[50]), .Z(n7257) );
  NAND U7770 ( .A(n37295), .B(n7257), .Z(n7091) );
  AND U7771 ( .A(n7092), .B(n7091), .Z(n7201) );
  NAND U7772 ( .A(n186), .B(n7093), .Z(n7095) );
  XOR U7773 ( .A(b[11]), .B(a[52]), .Z(n7260) );
  NAND U7774 ( .A(n37097), .B(n7260), .Z(n7094) );
  NAND U7775 ( .A(n7095), .B(n7094), .Z(n7200) );
  XNOR U7776 ( .A(n7201), .B(n7200), .Z(n7202) );
  NAND U7777 ( .A(n188), .B(n7096), .Z(n7098) );
  XOR U7778 ( .A(b[15]), .B(a[48]), .Z(n7263) );
  NAND U7779 ( .A(n37382), .B(n7263), .Z(n7097) );
  AND U7780 ( .A(n7098), .B(n7097), .Z(n7197) );
  NAND U7781 ( .A(n38064), .B(n7099), .Z(n7101) );
  XOR U7782 ( .A(b[21]), .B(a[42]), .Z(n7266) );
  NAND U7783 ( .A(n37993), .B(n7266), .Z(n7100) );
  AND U7784 ( .A(n7101), .B(n7100), .Z(n7195) );
  NAND U7785 ( .A(n185), .B(n7102), .Z(n7104) );
  XOR U7786 ( .A(b[9]), .B(a[54]), .Z(n7269) );
  NAND U7787 ( .A(n36805), .B(n7269), .Z(n7103) );
  NAND U7788 ( .A(n7104), .B(n7103), .Z(n7194) );
  XNOR U7789 ( .A(n7195), .B(n7194), .Z(n7196) );
  XOR U7790 ( .A(n7197), .B(n7196), .Z(n7203) );
  XOR U7791 ( .A(n7202), .B(n7203), .Z(n7209) );
  XOR U7792 ( .A(n7208), .B(n7209), .Z(n7221) );
  XNOR U7793 ( .A(n7220), .B(n7221), .Z(n7152) );
  XNOR U7794 ( .A(n7153), .B(n7152), .Z(n7154) );
  XOR U7795 ( .A(n7155), .B(n7154), .Z(n7273) );
  XOR U7796 ( .A(n7272), .B(n7273), .Z(n7275) );
  XOR U7797 ( .A(n7274), .B(n7275), .Z(n7149) );
  NANDN U7798 ( .A(n7106), .B(n7105), .Z(n7110) );
  NAND U7799 ( .A(n7108), .B(n7107), .Z(n7109) );
  AND U7800 ( .A(n7110), .B(n7109), .Z(n7147) );
  NANDN U7801 ( .A(n7112), .B(n7111), .Z(n7116) );
  NANDN U7802 ( .A(n7114), .B(n7113), .Z(n7115) );
  AND U7803 ( .A(n7116), .B(n7115), .Z(n7146) );
  XNOR U7804 ( .A(n7147), .B(n7146), .Z(n7148) );
  XNOR U7805 ( .A(n7149), .B(n7148), .Z(n7140) );
  NANDN U7806 ( .A(n7118), .B(n7117), .Z(n7122) );
  NANDN U7807 ( .A(n7120), .B(n7119), .Z(n7121) );
  NAND U7808 ( .A(n7122), .B(n7121), .Z(n7141) );
  XNOR U7809 ( .A(n7140), .B(n7141), .Z(n7142) );
  NANDN U7810 ( .A(n7124), .B(n7123), .Z(n7128) );
  NAND U7811 ( .A(n7126), .B(n7125), .Z(n7127) );
  NAND U7812 ( .A(n7128), .B(n7127), .Z(n7143) );
  XNOR U7813 ( .A(n7142), .B(n7143), .Z(n7134) );
  XNOR U7814 ( .A(n7135), .B(n7134), .Z(n7136) );
  XNOR U7815 ( .A(n7137), .B(n7136), .Z(n7278) );
  XNOR U7816 ( .A(sreg[286]), .B(n7278), .Z(n7280) );
  NANDN U7817 ( .A(sreg[285]), .B(n7129), .Z(n7133) );
  NAND U7818 ( .A(n7131), .B(n7130), .Z(n7132) );
  NAND U7819 ( .A(n7133), .B(n7132), .Z(n7279) );
  XNOR U7820 ( .A(n7280), .B(n7279), .Z(c[286]) );
  NANDN U7821 ( .A(n7135), .B(n7134), .Z(n7139) );
  NANDN U7822 ( .A(n7137), .B(n7136), .Z(n7138) );
  AND U7823 ( .A(n7139), .B(n7138), .Z(n7286) );
  NANDN U7824 ( .A(n7141), .B(n7140), .Z(n7145) );
  NANDN U7825 ( .A(n7143), .B(n7142), .Z(n7144) );
  AND U7826 ( .A(n7145), .B(n7144), .Z(n7284) );
  NANDN U7827 ( .A(n7147), .B(n7146), .Z(n7151) );
  NANDN U7828 ( .A(n7149), .B(n7148), .Z(n7150) );
  AND U7829 ( .A(n7151), .B(n7150), .Z(n7292) );
  NANDN U7830 ( .A(n7153), .B(n7152), .Z(n7157) );
  NANDN U7831 ( .A(n7155), .B(n7154), .Z(n7156) );
  AND U7832 ( .A(n7157), .B(n7156), .Z(n7296) );
  NANDN U7833 ( .A(n7159), .B(n7158), .Z(n7163) );
  NAND U7834 ( .A(n7161), .B(n7160), .Z(n7162) );
  AND U7835 ( .A(n7163), .B(n7162), .Z(n7295) );
  XNOR U7836 ( .A(n7296), .B(n7295), .Z(n7298) );
  NANDN U7837 ( .A(n7165), .B(n7164), .Z(n7169) );
  NANDN U7838 ( .A(n7167), .B(n7166), .Z(n7168) );
  AND U7839 ( .A(n7169), .B(n7168), .Z(n7375) );
  NAND U7840 ( .A(n38385), .B(n7170), .Z(n7172) );
  XOR U7841 ( .A(b[27]), .B(a[37]), .Z(n7319) );
  NAND U7842 ( .A(n38343), .B(n7319), .Z(n7171) );
  AND U7843 ( .A(n7172), .B(n7171), .Z(n7382) );
  NAND U7844 ( .A(n183), .B(n7173), .Z(n7175) );
  XOR U7845 ( .A(b[5]), .B(a[59]), .Z(n7322) );
  NAND U7846 ( .A(n36296), .B(n7322), .Z(n7174) );
  AND U7847 ( .A(n7175), .B(n7174), .Z(n7380) );
  NAND U7848 ( .A(n190), .B(n7176), .Z(n7178) );
  XOR U7849 ( .A(b[19]), .B(a[45]), .Z(n7325) );
  NAND U7850 ( .A(n37821), .B(n7325), .Z(n7177) );
  NAND U7851 ( .A(n7178), .B(n7177), .Z(n7379) );
  XNOR U7852 ( .A(n7380), .B(n7379), .Z(n7381) );
  XNOR U7853 ( .A(n7382), .B(n7381), .Z(n7373) );
  NAND U7854 ( .A(n38470), .B(n7179), .Z(n7181) );
  XOR U7855 ( .A(b[31]), .B(a[33]), .Z(n7328) );
  NAND U7856 ( .A(n38453), .B(n7328), .Z(n7180) );
  AND U7857 ( .A(n7181), .B(n7180), .Z(n7340) );
  NAND U7858 ( .A(n181), .B(n7182), .Z(n7184) );
  XOR U7859 ( .A(b[3]), .B(a[61]), .Z(n7331) );
  NAND U7860 ( .A(n182), .B(n7331), .Z(n7183) );
  AND U7861 ( .A(n7184), .B(n7183), .Z(n7338) );
  NAND U7862 ( .A(n189), .B(n7185), .Z(n7187) );
  XOR U7863 ( .A(b[17]), .B(a[47]), .Z(n7334) );
  NAND U7864 ( .A(n37652), .B(n7334), .Z(n7186) );
  NAND U7865 ( .A(n7187), .B(n7186), .Z(n7337) );
  XNOR U7866 ( .A(n7338), .B(n7337), .Z(n7339) );
  XOR U7867 ( .A(n7340), .B(n7339), .Z(n7374) );
  XOR U7868 ( .A(n7373), .B(n7374), .Z(n7376) );
  XOR U7869 ( .A(n7375), .B(n7376), .Z(n7308) );
  NANDN U7870 ( .A(n7189), .B(n7188), .Z(n7193) );
  NANDN U7871 ( .A(n7191), .B(n7190), .Z(n7192) );
  AND U7872 ( .A(n7193), .B(n7192), .Z(n7361) );
  NANDN U7873 ( .A(n7195), .B(n7194), .Z(n7199) );
  NANDN U7874 ( .A(n7197), .B(n7196), .Z(n7198) );
  NAND U7875 ( .A(n7199), .B(n7198), .Z(n7362) );
  XNOR U7876 ( .A(n7361), .B(n7362), .Z(n7363) );
  NANDN U7877 ( .A(n7201), .B(n7200), .Z(n7205) );
  NANDN U7878 ( .A(n7203), .B(n7202), .Z(n7204) );
  NAND U7879 ( .A(n7205), .B(n7204), .Z(n7364) );
  XNOR U7880 ( .A(n7363), .B(n7364), .Z(n7307) );
  XNOR U7881 ( .A(n7308), .B(n7307), .Z(n7310) );
  NANDN U7882 ( .A(n7207), .B(n7206), .Z(n7211) );
  NANDN U7883 ( .A(n7209), .B(n7208), .Z(n7210) );
  AND U7884 ( .A(n7211), .B(n7210), .Z(n7309) );
  XOR U7885 ( .A(n7310), .B(n7309), .Z(n7424) );
  NANDN U7886 ( .A(n7213), .B(n7212), .Z(n7217) );
  NANDN U7887 ( .A(n7215), .B(n7214), .Z(n7216) );
  AND U7888 ( .A(n7217), .B(n7216), .Z(n7421) );
  NANDN U7889 ( .A(n7219), .B(n7218), .Z(n7223) );
  NANDN U7890 ( .A(n7221), .B(n7220), .Z(n7222) );
  AND U7891 ( .A(n7223), .B(n7222), .Z(n7304) );
  NANDN U7892 ( .A(n7225), .B(n7224), .Z(n7229) );
  OR U7893 ( .A(n7227), .B(n7226), .Z(n7228) );
  AND U7894 ( .A(n7229), .B(n7228), .Z(n7302) );
  NANDN U7895 ( .A(n7231), .B(n7230), .Z(n7235) );
  NANDN U7896 ( .A(n7233), .B(n7232), .Z(n7234) );
  AND U7897 ( .A(n7235), .B(n7234), .Z(n7368) );
  NANDN U7898 ( .A(n7237), .B(n7236), .Z(n7241) );
  NANDN U7899 ( .A(n7239), .B(n7238), .Z(n7240) );
  NAND U7900 ( .A(n7241), .B(n7240), .Z(n7367) );
  XNOR U7901 ( .A(n7368), .B(n7367), .Z(n7369) );
  NAND U7902 ( .A(b[0]), .B(a[63]), .Z(n7242) );
  XNOR U7903 ( .A(b[1]), .B(n7242), .Z(n7244) );
  NANDN U7904 ( .A(b[0]), .B(a[62]), .Z(n7243) );
  NAND U7905 ( .A(n7244), .B(n7243), .Z(n7316) );
  NAND U7906 ( .A(n194), .B(n7245), .Z(n7247) );
  XOR U7907 ( .A(b[29]), .B(a[35]), .Z(n7394) );
  NAND U7908 ( .A(n38456), .B(n7394), .Z(n7246) );
  AND U7909 ( .A(n7247), .B(n7246), .Z(n7314) );
  AND U7910 ( .A(b[31]), .B(a[31]), .Z(n7313) );
  XNOR U7911 ( .A(n7314), .B(n7313), .Z(n7315) );
  XNOR U7912 ( .A(n7316), .B(n7315), .Z(n7355) );
  NAND U7913 ( .A(n38185), .B(n7248), .Z(n7250) );
  XOR U7914 ( .A(b[23]), .B(a[41]), .Z(n7397) );
  NAND U7915 ( .A(n38132), .B(n7397), .Z(n7249) );
  AND U7916 ( .A(n7250), .B(n7249), .Z(n7388) );
  NAND U7917 ( .A(n184), .B(n7251), .Z(n7253) );
  XOR U7918 ( .A(b[7]), .B(a[57]), .Z(n7400) );
  NAND U7919 ( .A(n36592), .B(n7400), .Z(n7252) );
  AND U7920 ( .A(n7253), .B(n7252), .Z(n7386) );
  NAND U7921 ( .A(n38289), .B(n7254), .Z(n7256) );
  XOR U7922 ( .A(b[25]), .B(a[39]), .Z(n7403) );
  NAND U7923 ( .A(n38247), .B(n7403), .Z(n7255) );
  NAND U7924 ( .A(n7256), .B(n7255), .Z(n7385) );
  XNOR U7925 ( .A(n7386), .B(n7385), .Z(n7387) );
  XOR U7926 ( .A(n7388), .B(n7387), .Z(n7356) );
  XNOR U7927 ( .A(n7355), .B(n7356), .Z(n7357) );
  NAND U7928 ( .A(n187), .B(n7257), .Z(n7259) );
  XOR U7929 ( .A(b[13]), .B(a[51]), .Z(n7406) );
  NAND U7930 ( .A(n37295), .B(n7406), .Z(n7258) );
  AND U7931 ( .A(n7259), .B(n7258), .Z(n7350) );
  NAND U7932 ( .A(n186), .B(n7260), .Z(n7262) );
  XOR U7933 ( .A(b[11]), .B(a[53]), .Z(n7409) );
  NAND U7934 ( .A(n37097), .B(n7409), .Z(n7261) );
  NAND U7935 ( .A(n7262), .B(n7261), .Z(n7349) );
  XNOR U7936 ( .A(n7350), .B(n7349), .Z(n7351) );
  NAND U7937 ( .A(n188), .B(n7263), .Z(n7265) );
  XOR U7938 ( .A(b[15]), .B(a[49]), .Z(n7412) );
  NAND U7939 ( .A(n37382), .B(n7412), .Z(n7264) );
  AND U7940 ( .A(n7265), .B(n7264), .Z(n7346) );
  NAND U7941 ( .A(n38064), .B(n7266), .Z(n7268) );
  XOR U7942 ( .A(b[21]), .B(a[43]), .Z(n7415) );
  NAND U7943 ( .A(n37993), .B(n7415), .Z(n7267) );
  AND U7944 ( .A(n7268), .B(n7267), .Z(n7344) );
  NAND U7945 ( .A(n185), .B(n7269), .Z(n7271) );
  XOR U7946 ( .A(b[9]), .B(a[55]), .Z(n7418) );
  NAND U7947 ( .A(n36805), .B(n7418), .Z(n7270) );
  NAND U7948 ( .A(n7271), .B(n7270), .Z(n7343) );
  XNOR U7949 ( .A(n7344), .B(n7343), .Z(n7345) );
  XOR U7950 ( .A(n7346), .B(n7345), .Z(n7352) );
  XOR U7951 ( .A(n7351), .B(n7352), .Z(n7358) );
  XOR U7952 ( .A(n7357), .B(n7358), .Z(n7370) );
  XNOR U7953 ( .A(n7369), .B(n7370), .Z(n7301) );
  XNOR U7954 ( .A(n7302), .B(n7301), .Z(n7303) );
  XOR U7955 ( .A(n7304), .B(n7303), .Z(n7422) );
  XNOR U7956 ( .A(n7421), .B(n7422), .Z(n7423) );
  XNOR U7957 ( .A(n7424), .B(n7423), .Z(n7297) );
  XOR U7958 ( .A(n7298), .B(n7297), .Z(n7290) );
  NANDN U7959 ( .A(n7273), .B(n7272), .Z(n7277) );
  OR U7960 ( .A(n7275), .B(n7274), .Z(n7276) );
  AND U7961 ( .A(n7277), .B(n7276), .Z(n7289) );
  XNOR U7962 ( .A(n7290), .B(n7289), .Z(n7291) );
  XNOR U7963 ( .A(n7292), .B(n7291), .Z(n7283) );
  XNOR U7964 ( .A(n7284), .B(n7283), .Z(n7285) );
  XNOR U7965 ( .A(n7286), .B(n7285), .Z(n7427) );
  XNOR U7966 ( .A(sreg[287]), .B(n7427), .Z(n7429) );
  NANDN U7967 ( .A(sreg[286]), .B(n7278), .Z(n7282) );
  NAND U7968 ( .A(n7280), .B(n7279), .Z(n7281) );
  NAND U7969 ( .A(n7282), .B(n7281), .Z(n7428) );
  XNOR U7970 ( .A(n7429), .B(n7428), .Z(c[287]) );
  NANDN U7971 ( .A(n7284), .B(n7283), .Z(n7288) );
  NANDN U7972 ( .A(n7286), .B(n7285), .Z(n7287) );
  AND U7973 ( .A(n7288), .B(n7287), .Z(n7435) );
  NANDN U7974 ( .A(n7290), .B(n7289), .Z(n7294) );
  NANDN U7975 ( .A(n7292), .B(n7291), .Z(n7293) );
  AND U7976 ( .A(n7294), .B(n7293), .Z(n7433) );
  NANDN U7977 ( .A(n7296), .B(n7295), .Z(n7300) );
  NAND U7978 ( .A(n7298), .B(n7297), .Z(n7299) );
  AND U7979 ( .A(n7300), .B(n7299), .Z(n7440) );
  NANDN U7980 ( .A(n7302), .B(n7301), .Z(n7306) );
  NANDN U7981 ( .A(n7304), .B(n7303), .Z(n7305) );
  AND U7982 ( .A(n7306), .B(n7305), .Z(n7445) );
  NANDN U7983 ( .A(n7308), .B(n7307), .Z(n7312) );
  NAND U7984 ( .A(n7310), .B(n7309), .Z(n7311) );
  AND U7985 ( .A(n7312), .B(n7311), .Z(n7444) );
  XNOR U7986 ( .A(n7445), .B(n7444), .Z(n7447) );
  NANDN U7987 ( .A(n7314), .B(n7313), .Z(n7318) );
  NANDN U7988 ( .A(n7316), .B(n7315), .Z(n7317) );
  AND U7989 ( .A(n7318), .B(n7317), .Z(n7524) );
  NAND U7990 ( .A(n38385), .B(n7319), .Z(n7321) );
  XOR U7991 ( .A(b[27]), .B(a[38]), .Z(n7468) );
  NAND U7992 ( .A(n38343), .B(n7468), .Z(n7320) );
  AND U7993 ( .A(n7321), .B(n7320), .Z(n7531) );
  NAND U7994 ( .A(n183), .B(n7322), .Z(n7324) );
  XOR U7995 ( .A(b[5]), .B(a[60]), .Z(n7471) );
  NAND U7996 ( .A(n36296), .B(n7471), .Z(n7323) );
  AND U7997 ( .A(n7324), .B(n7323), .Z(n7529) );
  NAND U7998 ( .A(n190), .B(n7325), .Z(n7327) );
  XOR U7999 ( .A(b[19]), .B(a[46]), .Z(n7474) );
  NAND U8000 ( .A(n37821), .B(n7474), .Z(n7326) );
  NAND U8001 ( .A(n7327), .B(n7326), .Z(n7528) );
  XNOR U8002 ( .A(n7529), .B(n7528), .Z(n7530) );
  XNOR U8003 ( .A(n7531), .B(n7530), .Z(n7522) );
  NAND U8004 ( .A(n38470), .B(n7328), .Z(n7330) );
  XOR U8005 ( .A(b[31]), .B(a[34]), .Z(n7477) );
  NAND U8006 ( .A(n38453), .B(n7477), .Z(n7329) );
  AND U8007 ( .A(n7330), .B(n7329), .Z(n7489) );
  NAND U8008 ( .A(n181), .B(n7331), .Z(n7333) );
  XOR U8009 ( .A(b[3]), .B(a[62]), .Z(n7480) );
  NAND U8010 ( .A(n182), .B(n7480), .Z(n7332) );
  AND U8011 ( .A(n7333), .B(n7332), .Z(n7487) );
  NAND U8012 ( .A(n189), .B(n7334), .Z(n7336) );
  XOR U8013 ( .A(b[17]), .B(a[48]), .Z(n7483) );
  NAND U8014 ( .A(n37652), .B(n7483), .Z(n7335) );
  NAND U8015 ( .A(n7336), .B(n7335), .Z(n7486) );
  XNOR U8016 ( .A(n7487), .B(n7486), .Z(n7488) );
  XOR U8017 ( .A(n7489), .B(n7488), .Z(n7523) );
  XOR U8018 ( .A(n7522), .B(n7523), .Z(n7525) );
  XOR U8019 ( .A(n7524), .B(n7525), .Z(n7457) );
  NANDN U8020 ( .A(n7338), .B(n7337), .Z(n7342) );
  NANDN U8021 ( .A(n7340), .B(n7339), .Z(n7341) );
  AND U8022 ( .A(n7342), .B(n7341), .Z(n7510) );
  NANDN U8023 ( .A(n7344), .B(n7343), .Z(n7348) );
  NANDN U8024 ( .A(n7346), .B(n7345), .Z(n7347) );
  NAND U8025 ( .A(n7348), .B(n7347), .Z(n7511) );
  XNOR U8026 ( .A(n7510), .B(n7511), .Z(n7512) );
  NANDN U8027 ( .A(n7350), .B(n7349), .Z(n7354) );
  NANDN U8028 ( .A(n7352), .B(n7351), .Z(n7353) );
  NAND U8029 ( .A(n7354), .B(n7353), .Z(n7513) );
  XNOR U8030 ( .A(n7512), .B(n7513), .Z(n7456) );
  XNOR U8031 ( .A(n7457), .B(n7456), .Z(n7459) );
  NANDN U8032 ( .A(n7356), .B(n7355), .Z(n7360) );
  NANDN U8033 ( .A(n7358), .B(n7357), .Z(n7359) );
  AND U8034 ( .A(n7360), .B(n7359), .Z(n7458) );
  XOR U8035 ( .A(n7459), .B(n7458), .Z(n7573) );
  NANDN U8036 ( .A(n7362), .B(n7361), .Z(n7366) );
  NANDN U8037 ( .A(n7364), .B(n7363), .Z(n7365) );
  AND U8038 ( .A(n7366), .B(n7365), .Z(n7570) );
  NANDN U8039 ( .A(n7368), .B(n7367), .Z(n7372) );
  NANDN U8040 ( .A(n7370), .B(n7369), .Z(n7371) );
  AND U8041 ( .A(n7372), .B(n7371), .Z(n7453) );
  NANDN U8042 ( .A(n7374), .B(n7373), .Z(n7378) );
  OR U8043 ( .A(n7376), .B(n7375), .Z(n7377) );
  AND U8044 ( .A(n7378), .B(n7377), .Z(n7451) );
  NANDN U8045 ( .A(n7380), .B(n7379), .Z(n7384) );
  NANDN U8046 ( .A(n7382), .B(n7381), .Z(n7383) );
  AND U8047 ( .A(n7384), .B(n7383), .Z(n7517) );
  NANDN U8048 ( .A(n7386), .B(n7385), .Z(n7390) );
  NANDN U8049 ( .A(n7388), .B(n7387), .Z(n7389) );
  NAND U8050 ( .A(n7390), .B(n7389), .Z(n7516) );
  XNOR U8051 ( .A(n7517), .B(n7516), .Z(n7518) );
  NAND U8052 ( .A(b[0]), .B(a[64]), .Z(n7391) );
  XNOR U8053 ( .A(b[1]), .B(n7391), .Z(n7393) );
  NANDN U8054 ( .A(b[0]), .B(a[63]), .Z(n7392) );
  NAND U8055 ( .A(n7393), .B(n7392), .Z(n7465) );
  NAND U8056 ( .A(n194), .B(n7394), .Z(n7396) );
  XOR U8057 ( .A(b[29]), .B(a[36]), .Z(n7543) );
  NAND U8058 ( .A(n38456), .B(n7543), .Z(n7395) );
  AND U8059 ( .A(n7396), .B(n7395), .Z(n7463) );
  AND U8060 ( .A(b[31]), .B(a[32]), .Z(n7462) );
  XNOR U8061 ( .A(n7463), .B(n7462), .Z(n7464) );
  XNOR U8062 ( .A(n7465), .B(n7464), .Z(n7504) );
  NAND U8063 ( .A(n38185), .B(n7397), .Z(n7399) );
  XOR U8064 ( .A(b[23]), .B(a[42]), .Z(n7546) );
  NAND U8065 ( .A(n38132), .B(n7546), .Z(n7398) );
  AND U8066 ( .A(n7399), .B(n7398), .Z(n7537) );
  NAND U8067 ( .A(n184), .B(n7400), .Z(n7402) );
  XOR U8068 ( .A(b[7]), .B(a[58]), .Z(n7549) );
  NAND U8069 ( .A(n36592), .B(n7549), .Z(n7401) );
  AND U8070 ( .A(n7402), .B(n7401), .Z(n7535) );
  NAND U8071 ( .A(n38289), .B(n7403), .Z(n7405) );
  XOR U8072 ( .A(b[25]), .B(a[40]), .Z(n7552) );
  NAND U8073 ( .A(n38247), .B(n7552), .Z(n7404) );
  NAND U8074 ( .A(n7405), .B(n7404), .Z(n7534) );
  XNOR U8075 ( .A(n7535), .B(n7534), .Z(n7536) );
  XOR U8076 ( .A(n7537), .B(n7536), .Z(n7505) );
  XNOR U8077 ( .A(n7504), .B(n7505), .Z(n7506) );
  NAND U8078 ( .A(n187), .B(n7406), .Z(n7408) );
  XOR U8079 ( .A(b[13]), .B(a[52]), .Z(n7555) );
  NAND U8080 ( .A(n37295), .B(n7555), .Z(n7407) );
  AND U8081 ( .A(n7408), .B(n7407), .Z(n7499) );
  NAND U8082 ( .A(n186), .B(n7409), .Z(n7411) );
  XOR U8083 ( .A(b[11]), .B(a[54]), .Z(n7558) );
  NAND U8084 ( .A(n37097), .B(n7558), .Z(n7410) );
  NAND U8085 ( .A(n7411), .B(n7410), .Z(n7498) );
  XNOR U8086 ( .A(n7499), .B(n7498), .Z(n7500) );
  NAND U8087 ( .A(n188), .B(n7412), .Z(n7414) );
  XOR U8088 ( .A(b[15]), .B(a[50]), .Z(n7561) );
  NAND U8089 ( .A(n37382), .B(n7561), .Z(n7413) );
  AND U8090 ( .A(n7414), .B(n7413), .Z(n7495) );
  NAND U8091 ( .A(n38064), .B(n7415), .Z(n7417) );
  XOR U8092 ( .A(b[21]), .B(a[44]), .Z(n7564) );
  NAND U8093 ( .A(n37993), .B(n7564), .Z(n7416) );
  AND U8094 ( .A(n7417), .B(n7416), .Z(n7493) );
  NAND U8095 ( .A(n185), .B(n7418), .Z(n7420) );
  XOR U8096 ( .A(b[9]), .B(a[56]), .Z(n7567) );
  NAND U8097 ( .A(n36805), .B(n7567), .Z(n7419) );
  NAND U8098 ( .A(n7420), .B(n7419), .Z(n7492) );
  XNOR U8099 ( .A(n7493), .B(n7492), .Z(n7494) );
  XOR U8100 ( .A(n7495), .B(n7494), .Z(n7501) );
  XOR U8101 ( .A(n7500), .B(n7501), .Z(n7507) );
  XOR U8102 ( .A(n7506), .B(n7507), .Z(n7519) );
  XNOR U8103 ( .A(n7518), .B(n7519), .Z(n7450) );
  XNOR U8104 ( .A(n7451), .B(n7450), .Z(n7452) );
  XOR U8105 ( .A(n7453), .B(n7452), .Z(n7571) );
  XNOR U8106 ( .A(n7570), .B(n7571), .Z(n7572) );
  XNOR U8107 ( .A(n7573), .B(n7572), .Z(n7446) );
  XOR U8108 ( .A(n7447), .B(n7446), .Z(n7439) );
  NANDN U8109 ( .A(n7422), .B(n7421), .Z(n7426) );
  NANDN U8110 ( .A(n7424), .B(n7423), .Z(n7425) );
  AND U8111 ( .A(n7426), .B(n7425), .Z(n7438) );
  XOR U8112 ( .A(n7439), .B(n7438), .Z(n7441) );
  XNOR U8113 ( .A(n7440), .B(n7441), .Z(n7432) );
  XNOR U8114 ( .A(n7433), .B(n7432), .Z(n7434) );
  XNOR U8115 ( .A(n7435), .B(n7434), .Z(n7576) );
  XNOR U8116 ( .A(sreg[288]), .B(n7576), .Z(n7578) );
  NANDN U8117 ( .A(sreg[287]), .B(n7427), .Z(n7431) );
  NAND U8118 ( .A(n7429), .B(n7428), .Z(n7430) );
  NAND U8119 ( .A(n7431), .B(n7430), .Z(n7577) );
  XNOR U8120 ( .A(n7578), .B(n7577), .Z(c[288]) );
  NANDN U8121 ( .A(n7433), .B(n7432), .Z(n7437) );
  NANDN U8122 ( .A(n7435), .B(n7434), .Z(n7436) );
  AND U8123 ( .A(n7437), .B(n7436), .Z(n7584) );
  NANDN U8124 ( .A(n7439), .B(n7438), .Z(n7443) );
  NANDN U8125 ( .A(n7441), .B(n7440), .Z(n7442) );
  AND U8126 ( .A(n7443), .B(n7442), .Z(n7582) );
  NANDN U8127 ( .A(n7445), .B(n7444), .Z(n7449) );
  NAND U8128 ( .A(n7447), .B(n7446), .Z(n7448) );
  AND U8129 ( .A(n7449), .B(n7448), .Z(n7589) );
  NANDN U8130 ( .A(n7451), .B(n7450), .Z(n7455) );
  NANDN U8131 ( .A(n7453), .B(n7452), .Z(n7454) );
  AND U8132 ( .A(n7455), .B(n7454), .Z(n7720) );
  NANDN U8133 ( .A(n7457), .B(n7456), .Z(n7461) );
  NAND U8134 ( .A(n7459), .B(n7458), .Z(n7460) );
  AND U8135 ( .A(n7461), .B(n7460), .Z(n7719) );
  XNOR U8136 ( .A(n7720), .B(n7719), .Z(n7722) );
  NANDN U8137 ( .A(n7463), .B(n7462), .Z(n7467) );
  NANDN U8138 ( .A(n7465), .B(n7464), .Z(n7466) );
  AND U8139 ( .A(n7467), .B(n7466), .Z(n7667) );
  NAND U8140 ( .A(n38385), .B(n7468), .Z(n7470) );
  XOR U8141 ( .A(b[27]), .B(a[39]), .Z(n7611) );
  NAND U8142 ( .A(n38343), .B(n7611), .Z(n7469) );
  AND U8143 ( .A(n7470), .B(n7469), .Z(n7674) );
  NAND U8144 ( .A(n183), .B(n7471), .Z(n7473) );
  XOR U8145 ( .A(b[5]), .B(a[61]), .Z(n7614) );
  NAND U8146 ( .A(n36296), .B(n7614), .Z(n7472) );
  AND U8147 ( .A(n7473), .B(n7472), .Z(n7672) );
  NAND U8148 ( .A(n190), .B(n7474), .Z(n7476) );
  XOR U8149 ( .A(b[19]), .B(a[47]), .Z(n7617) );
  NAND U8150 ( .A(n37821), .B(n7617), .Z(n7475) );
  NAND U8151 ( .A(n7476), .B(n7475), .Z(n7671) );
  XNOR U8152 ( .A(n7672), .B(n7671), .Z(n7673) );
  XNOR U8153 ( .A(n7674), .B(n7673), .Z(n7665) );
  NAND U8154 ( .A(n38470), .B(n7477), .Z(n7479) );
  XOR U8155 ( .A(b[31]), .B(a[35]), .Z(n7620) );
  NAND U8156 ( .A(n38453), .B(n7620), .Z(n7478) );
  AND U8157 ( .A(n7479), .B(n7478), .Z(n7632) );
  NAND U8158 ( .A(n181), .B(n7480), .Z(n7482) );
  XOR U8159 ( .A(b[3]), .B(a[63]), .Z(n7623) );
  NAND U8160 ( .A(n182), .B(n7623), .Z(n7481) );
  AND U8161 ( .A(n7482), .B(n7481), .Z(n7630) );
  NAND U8162 ( .A(n189), .B(n7483), .Z(n7485) );
  XOR U8163 ( .A(b[17]), .B(a[49]), .Z(n7626) );
  NAND U8164 ( .A(n37652), .B(n7626), .Z(n7484) );
  NAND U8165 ( .A(n7485), .B(n7484), .Z(n7629) );
  XNOR U8166 ( .A(n7630), .B(n7629), .Z(n7631) );
  XOR U8167 ( .A(n7632), .B(n7631), .Z(n7666) );
  XOR U8168 ( .A(n7665), .B(n7666), .Z(n7668) );
  XOR U8169 ( .A(n7667), .B(n7668), .Z(n7600) );
  NANDN U8170 ( .A(n7487), .B(n7486), .Z(n7491) );
  NANDN U8171 ( .A(n7489), .B(n7488), .Z(n7490) );
  AND U8172 ( .A(n7491), .B(n7490), .Z(n7653) );
  NANDN U8173 ( .A(n7493), .B(n7492), .Z(n7497) );
  NANDN U8174 ( .A(n7495), .B(n7494), .Z(n7496) );
  NAND U8175 ( .A(n7497), .B(n7496), .Z(n7654) );
  XNOR U8176 ( .A(n7653), .B(n7654), .Z(n7655) );
  NANDN U8177 ( .A(n7499), .B(n7498), .Z(n7503) );
  NANDN U8178 ( .A(n7501), .B(n7500), .Z(n7502) );
  NAND U8179 ( .A(n7503), .B(n7502), .Z(n7656) );
  XNOR U8180 ( .A(n7655), .B(n7656), .Z(n7599) );
  XNOR U8181 ( .A(n7600), .B(n7599), .Z(n7602) );
  NANDN U8182 ( .A(n7505), .B(n7504), .Z(n7509) );
  NANDN U8183 ( .A(n7507), .B(n7506), .Z(n7508) );
  AND U8184 ( .A(n7509), .B(n7508), .Z(n7601) );
  XOR U8185 ( .A(n7602), .B(n7601), .Z(n7716) );
  NANDN U8186 ( .A(n7511), .B(n7510), .Z(n7515) );
  NANDN U8187 ( .A(n7513), .B(n7512), .Z(n7514) );
  AND U8188 ( .A(n7515), .B(n7514), .Z(n7713) );
  NANDN U8189 ( .A(n7517), .B(n7516), .Z(n7521) );
  NANDN U8190 ( .A(n7519), .B(n7518), .Z(n7520) );
  AND U8191 ( .A(n7521), .B(n7520), .Z(n7596) );
  NANDN U8192 ( .A(n7523), .B(n7522), .Z(n7527) );
  OR U8193 ( .A(n7525), .B(n7524), .Z(n7526) );
  AND U8194 ( .A(n7527), .B(n7526), .Z(n7594) );
  NANDN U8195 ( .A(n7529), .B(n7528), .Z(n7533) );
  NANDN U8196 ( .A(n7531), .B(n7530), .Z(n7532) );
  AND U8197 ( .A(n7533), .B(n7532), .Z(n7660) );
  NANDN U8198 ( .A(n7535), .B(n7534), .Z(n7539) );
  NANDN U8199 ( .A(n7537), .B(n7536), .Z(n7538) );
  NAND U8200 ( .A(n7539), .B(n7538), .Z(n7659) );
  XNOR U8201 ( .A(n7660), .B(n7659), .Z(n7661) );
  NAND U8202 ( .A(b[0]), .B(a[65]), .Z(n7540) );
  XNOR U8203 ( .A(b[1]), .B(n7540), .Z(n7542) );
  NANDN U8204 ( .A(b[0]), .B(a[64]), .Z(n7541) );
  NAND U8205 ( .A(n7542), .B(n7541), .Z(n7608) );
  NAND U8206 ( .A(n194), .B(n7543), .Z(n7545) );
  XOR U8207 ( .A(b[29]), .B(a[37]), .Z(n7686) );
  NAND U8208 ( .A(n38456), .B(n7686), .Z(n7544) );
  AND U8209 ( .A(n7545), .B(n7544), .Z(n7606) );
  AND U8210 ( .A(b[31]), .B(a[33]), .Z(n7605) );
  XNOR U8211 ( .A(n7606), .B(n7605), .Z(n7607) );
  XNOR U8212 ( .A(n7608), .B(n7607), .Z(n7647) );
  NAND U8213 ( .A(n38185), .B(n7546), .Z(n7548) );
  XOR U8214 ( .A(b[23]), .B(a[43]), .Z(n7689) );
  NAND U8215 ( .A(n38132), .B(n7689), .Z(n7547) );
  AND U8216 ( .A(n7548), .B(n7547), .Z(n7680) );
  NAND U8217 ( .A(n184), .B(n7549), .Z(n7551) );
  XOR U8218 ( .A(b[7]), .B(a[59]), .Z(n7692) );
  NAND U8219 ( .A(n36592), .B(n7692), .Z(n7550) );
  AND U8220 ( .A(n7551), .B(n7550), .Z(n7678) );
  NAND U8221 ( .A(n38289), .B(n7552), .Z(n7554) );
  XOR U8222 ( .A(b[25]), .B(a[41]), .Z(n7695) );
  NAND U8223 ( .A(n38247), .B(n7695), .Z(n7553) );
  NAND U8224 ( .A(n7554), .B(n7553), .Z(n7677) );
  XNOR U8225 ( .A(n7678), .B(n7677), .Z(n7679) );
  XOR U8226 ( .A(n7680), .B(n7679), .Z(n7648) );
  XNOR U8227 ( .A(n7647), .B(n7648), .Z(n7649) );
  NAND U8228 ( .A(n187), .B(n7555), .Z(n7557) );
  XOR U8229 ( .A(b[13]), .B(a[53]), .Z(n7698) );
  NAND U8230 ( .A(n37295), .B(n7698), .Z(n7556) );
  AND U8231 ( .A(n7557), .B(n7556), .Z(n7642) );
  NAND U8232 ( .A(n186), .B(n7558), .Z(n7560) );
  XOR U8233 ( .A(b[11]), .B(a[55]), .Z(n7701) );
  NAND U8234 ( .A(n37097), .B(n7701), .Z(n7559) );
  NAND U8235 ( .A(n7560), .B(n7559), .Z(n7641) );
  XNOR U8236 ( .A(n7642), .B(n7641), .Z(n7643) );
  NAND U8237 ( .A(n188), .B(n7561), .Z(n7563) );
  XOR U8238 ( .A(b[15]), .B(a[51]), .Z(n7704) );
  NAND U8239 ( .A(n37382), .B(n7704), .Z(n7562) );
  AND U8240 ( .A(n7563), .B(n7562), .Z(n7638) );
  NAND U8241 ( .A(n38064), .B(n7564), .Z(n7566) );
  XOR U8242 ( .A(b[21]), .B(a[45]), .Z(n7707) );
  NAND U8243 ( .A(n37993), .B(n7707), .Z(n7565) );
  AND U8244 ( .A(n7566), .B(n7565), .Z(n7636) );
  NAND U8245 ( .A(n185), .B(n7567), .Z(n7569) );
  XOR U8246 ( .A(b[9]), .B(a[57]), .Z(n7710) );
  NAND U8247 ( .A(n36805), .B(n7710), .Z(n7568) );
  NAND U8248 ( .A(n7569), .B(n7568), .Z(n7635) );
  XNOR U8249 ( .A(n7636), .B(n7635), .Z(n7637) );
  XOR U8250 ( .A(n7638), .B(n7637), .Z(n7644) );
  XOR U8251 ( .A(n7643), .B(n7644), .Z(n7650) );
  XOR U8252 ( .A(n7649), .B(n7650), .Z(n7662) );
  XNOR U8253 ( .A(n7661), .B(n7662), .Z(n7593) );
  XNOR U8254 ( .A(n7594), .B(n7593), .Z(n7595) );
  XOR U8255 ( .A(n7596), .B(n7595), .Z(n7714) );
  XNOR U8256 ( .A(n7713), .B(n7714), .Z(n7715) );
  XNOR U8257 ( .A(n7716), .B(n7715), .Z(n7721) );
  XOR U8258 ( .A(n7722), .B(n7721), .Z(n7588) );
  NANDN U8259 ( .A(n7571), .B(n7570), .Z(n7575) );
  NANDN U8260 ( .A(n7573), .B(n7572), .Z(n7574) );
  AND U8261 ( .A(n7575), .B(n7574), .Z(n7587) );
  XOR U8262 ( .A(n7588), .B(n7587), .Z(n7590) );
  XNOR U8263 ( .A(n7589), .B(n7590), .Z(n7581) );
  XNOR U8264 ( .A(n7582), .B(n7581), .Z(n7583) );
  XNOR U8265 ( .A(n7584), .B(n7583), .Z(n7725) );
  XNOR U8266 ( .A(sreg[289]), .B(n7725), .Z(n7727) );
  NANDN U8267 ( .A(sreg[288]), .B(n7576), .Z(n7580) );
  NAND U8268 ( .A(n7578), .B(n7577), .Z(n7579) );
  NAND U8269 ( .A(n7580), .B(n7579), .Z(n7726) );
  XNOR U8270 ( .A(n7727), .B(n7726), .Z(c[289]) );
  NANDN U8271 ( .A(n7582), .B(n7581), .Z(n7586) );
  NANDN U8272 ( .A(n7584), .B(n7583), .Z(n7585) );
  AND U8273 ( .A(n7586), .B(n7585), .Z(n7733) );
  NANDN U8274 ( .A(n7588), .B(n7587), .Z(n7592) );
  NANDN U8275 ( .A(n7590), .B(n7589), .Z(n7591) );
  AND U8276 ( .A(n7592), .B(n7591), .Z(n7731) );
  NANDN U8277 ( .A(n7594), .B(n7593), .Z(n7598) );
  NANDN U8278 ( .A(n7596), .B(n7595), .Z(n7597) );
  AND U8279 ( .A(n7598), .B(n7597), .Z(n7869) );
  NANDN U8280 ( .A(n7600), .B(n7599), .Z(n7604) );
  NAND U8281 ( .A(n7602), .B(n7601), .Z(n7603) );
  AND U8282 ( .A(n7604), .B(n7603), .Z(n7868) );
  XNOR U8283 ( .A(n7869), .B(n7868), .Z(n7871) );
  NANDN U8284 ( .A(n7606), .B(n7605), .Z(n7610) );
  NANDN U8285 ( .A(n7608), .B(n7607), .Z(n7609) );
  AND U8286 ( .A(n7610), .B(n7609), .Z(n7816) );
  NAND U8287 ( .A(n38385), .B(n7611), .Z(n7613) );
  XOR U8288 ( .A(b[27]), .B(a[40]), .Z(n7760) );
  NAND U8289 ( .A(n38343), .B(n7760), .Z(n7612) );
  AND U8290 ( .A(n7613), .B(n7612), .Z(n7823) );
  NAND U8291 ( .A(n183), .B(n7614), .Z(n7616) );
  XOR U8292 ( .A(b[5]), .B(a[62]), .Z(n7763) );
  NAND U8293 ( .A(n36296), .B(n7763), .Z(n7615) );
  AND U8294 ( .A(n7616), .B(n7615), .Z(n7821) );
  NAND U8295 ( .A(n190), .B(n7617), .Z(n7619) );
  XOR U8296 ( .A(b[19]), .B(a[48]), .Z(n7766) );
  NAND U8297 ( .A(n37821), .B(n7766), .Z(n7618) );
  NAND U8298 ( .A(n7619), .B(n7618), .Z(n7820) );
  XNOR U8299 ( .A(n7821), .B(n7820), .Z(n7822) );
  XNOR U8300 ( .A(n7823), .B(n7822), .Z(n7814) );
  NAND U8301 ( .A(n38470), .B(n7620), .Z(n7622) );
  XOR U8302 ( .A(b[31]), .B(a[36]), .Z(n7769) );
  NAND U8303 ( .A(n38453), .B(n7769), .Z(n7621) );
  AND U8304 ( .A(n7622), .B(n7621), .Z(n7781) );
  NAND U8305 ( .A(n181), .B(n7623), .Z(n7625) );
  XOR U8306 ( .A(b[3]), .B(a[64]), .Z(n7772) );
  NAND U8307 ( .A(n182), .B(n7772), .Z(n7624) );
  AND U8308 ( .A(n7625), .B(n7624), .Z(n7779) );
  NAND U8309 ( .A(n189), .B(n7626), .Z(n7628) );
  XOR U8310 ( .A(b[17]), .B(a[50]), .Z(n7775) );
  NAND U8311 ( .A(n37652), .B(n7775), .Z(n7627) );
  NAND U8312 ( .A(n7628), .B(n7627), .Z(n7778) );
  XNOR U8313 ( .A(n7779), .B(n7778), .Z(n7780) );
  XOR U8314 ( .A(n7781), .B(n7780), .Z(n7815) );
  XOR U8315 ( .A(n7814), .B(n7815), .Z(n7817) );
  XOR U8316 ( .A(n7816), .B(n7817), .Z(n7749) );
  NANDN U8317 ( .A(n7630), .B(n7629), .Z(n7634) );
  NANDN U8318 ( .A(n7632), .B(n7631), .Z(n7633) );
  AND U8319 ( .A(n7634), .B(n7633), .Z(n7802) );
  NANDN U8320 ( .A(n7636), .B(n7635), .Z(n7640) );
  NANDN U8321 ( .A(n7638), .B(n7637), .Z(n7639) );
  NAND U8322 ( .A(n7640), .B(n7639), .Z(n7803) );
  XNOR U8323 ( .A(n7802), .B(n7803), .Z(n7804) );
  NANDN U8324 ( .A(n7642), .B(n7641), .Z(n7646) );
  NANDN U8325 ( .A(n7644), .B(n7643), .Z(n7645) );
  NAND U8326 ( .A(n7646), .B(n7645), .Z(n7805) );
  XNOR U8327 ( .A(n7804), .B(n7805), .Z(n7748) );
  XNOR U8328 ( .A(n7749), .B(n7748), .Z(n7751) );
  NANDN U8329 ( .A(n7648), .B(n7647), .Z(n7652) );
  NANDN U8330 ( .A(n7650), .B(n7649), .Z(n7651) );
  AND U8331 ( .A(n7652), .B(n7651), .Z(n7750) );
  XOR U8332 ( .A(n7751), .B(n7750), .Z(n7865) );
  NANDN U8333 ( .A(n7654), .B(n7653), .Z(n7658) );
  NANDN U8334 ( .A(n7656), .B(n7655), .Z(n7657) );
  AND U8335 ( .A(n7658), .B(n7657), .Z(n7862) );
  NANDN U8336 ( .A(n7660), .B(n7659), .Z(n7664) );
  NANDN U8337 ( .A(n7662), .B(n7661), .Z(n7663) );
  AND U8338 ( .A(n7664), .B(n7663), .Z(n7745) );
  NANDN U8339 ( .A(n7666), .B(n7665), .Z(n7670) );
  OR U8340 ( .A(n7668), .B(n7667), .Z(n7669) );
  AND U8341 ( .A(n7670), .B(n7669), .Z(n7743) );
  NANDN U8342 ( .A(n7672), .B(n7671), .Z(n7676) );
  NANDN U8343 ( .A(n7674), .B(n7673), .Z(n7675) );
  AND U8344 ( .A(n7676), .B(n7675), .Z(n7809) );
  NANDN U8345 ( .A(n7678), .B(n7677), .Z(n7682) );
  NANDN U8346 ( .A(n7680), .B(n7679), .Z(n7681) );
  NAND U8347 ( .A(n7682), .B(n7681), .Z(n7808) );
  XNOR U8348 ( .A(n7809), .B(n7808), .Z(n7810) );
  NAND U8349 ( .A(b[0]), .B(a[66]), .Z(n7683) );
  XNOR U8350 ( .A(b[1]), .B(n7683), .Z(n7685) );
  NANDN U8351 ( .A(b[0]), .B(a[65]), .Z(n7684) );
  NAND U8352 ( .A(n7685), .B(n7684), .Z(n7757) );
  NAND U8353 ( .A(n194), .B(n7686), .Z(n7688) );
  XOR U8354 ( .A(b[29]), .B(a[38]), .Z(n7832) );
  NAND U8355 ( .A(n38456), .B(n7832), .Z(n7687) );
  AND U8356 ( .A(n7688), .B(n7687), .Z(n7755) );
  AND U8357 ( .A(b[31]), .B(a[34]), .Z(n7754) );
  XNOR U8358 ( .A(n7755), .B(n7754), .Z(n7756) );
  XNOR U8359 ( .A(n7757), .B(n7756), .Z(n7796) );
  NAND U8360 ( .A(n38185), .B(n7689), .Z(n7691) );
  XOR U8361 ( .A(b[23]), .B(a[44]), .Z(n7838) );
  NAND U8362 ( .A(n38132), .B(n7838), .Z(n7690) );
  AND U8363 ( .A(n7691), .B(n7690), .Z(n7829) );
  NAND U8364 ( .A(n184), .B(n7692), .Z(n7694) );
  XOR U8365 ( .A(b[7]), .B(a[60]), .Z(n7841) );
  NAND U8366 ( .A(n36592), .B(n7841), .Z(n7693) );
  AND U8367 ( .A(n7694), .B(n7693), .Z(n7827) );
  NAND U8368 ( .A(n38289), .B(n7695), .Z(n7697) );
  XOR U8369 ( .A(b[25]), .B(a[42]), .Z(n7844) );
  NAND U8370 ( .A(n38247), .B(n7844), .Z(n7696) );
  NAND U8371 ( .A(n7697), .B(n7696), .Z(n7826) );
  XNOR U8372 ( .A(n7827), .B(n7826), .Z(n7828) );
  XOR U8373 ( .A(n7829), .B(n7828), .Z(n7797) );
  XNOR U8374 ( .A(n7796), .B(n7797), .Z(n7798) );
  NAND U8375 ( .A(n187), .B(n7698), .Z(n7700) );
  XOR U8376 ( .A(b[13]), .B(a[54]), .Z(n7847) );
  NAND U8377 ( .A(n37295), .B(n7847), .Z(n7699) );
  AND U8378 ( .A(n7700), .B(n7699), .Z(n7791) );
  NAND U8379 ( .A(n186), .B(n7701), .Z(n7703) );
  XOR U8380 ( .A(b[11]), .B(a[56]), .Z(n7850) );
  NAND U8381 ( .A(n37097), .B(n7850), .Z(n7702) );
  NAND U8382 ( .A(n7703), .B(n7702), .Z(n7790) );
  XNOR U8383 ( .A(n7791), .B(n7790), .Z(n7792) );
  NAND U8384 ( .A(n188), .B(n7704), .Z(n7706) );
  XOR U8385 ( .A(b[15]), .B(a[52]), .Z(n7853) );
  NAND U8386 ( .A(n37382), .B(n7853), .Z(n7705) );
  AND U8387 ( .A(n7706), .B(n7705), .Z(n7787) );
  NAND U8388 ( .A(n38064), .B(n7707), .Z(n7709) );
  XOR U8389 ( .A(b[21]), .B(a[46]), .Z(n7856) );
  NAND U8390 ( .A(n37993), .B(n7856), .Z(n7708) );
  AND U8391 ( .A(n7709), .B(n7708), .Z(n7785) );
  NAND U8392 ( .A(n185), .B(n7710), .Z(n7712) );
  XOR U8393 ( .A(b[9]), .B(a[58]), .Z(n7859) );
  NAND U8394 ( .A(n36805), .B(n7859), .Z(n7711) );
  NAND U8395 ( .A(n7712), .B(n7711), .Z(n7784) );
  XNOR U8396 ( .A(n7785), .B(n7784), .Z(n7786) );
  XOR U8397 ( .A(n7787), .B(n7786), .Z(n7793) );
  XOR U8398 ( .A(n7792), .B(n7793), .Z(n7799) );
  XOR U8399 ( .A(n7798), .B(n7799), .Z(n7811) );
  XNOR U8400 ( .A(n7810), .B(n7811), .Z(n7742) );
  XNOR U8401 ( .A(n7743), .B(n7742), .Z(n7744) );
  XOR U8402 ( .A(n7745), .B(n7744), .Z(n7863) );
  XNOR U8403 ( .A(n7862), .B(n7863), .Z(n7864) );
  XNOR U8404 ( .A(n7865), .B(n7864), .Z(n7870) );
  XOR U8405 ( .A(n7871), .B(n7870), .Z(n7737) );
  NANDN U8406 ( .A(n7714), .B(n7713), .Z(n7718) );
  NANDN U8407 ( .A(n7716), .B(n7715), .Z(n7717) );
  AND U8408 ( .A(n7718), .B(n7717), .Z(n7736) );
  XNOR U8409 ( .A(n7737), .B(n7736), .Z(n7738) );
  NANDN U8410 ( .A(n7720), .B(n7719), .Z(n7724) );
  NAND U8411 ( .A(n7722), .B(n7721), .Z(n7723) );
  NAND U8412 ( .A(n7724), .B(n7723), .Z(n7739) );
  XNOR U8413 ( .A(n7738), .B(n7739), .Z(n7730) );
  XNOR U8414 ( .A(n7731), .B(n7730), .Z(n7732) );
  XNOR U8415 ( .A(n7733), .B(n7732), .Z(n7874) );
  XNOR U8416 ( .A(sreg[290]), .B(n7874), .Z(n7876) );
  NANDN U8417 ( .A(sreg[289]), .B(n7725), .Z(n7729) );
  NAND U8418 ( .A(n7727), .B(n7726), .Z(n7728) );
  NAND U8419 ( .A(n7729), .B(n7728), .Z(n7875) );
  XNOR U8420 ( .A(n7876), .B(n7875), .Z(c[290]) );
  NANDN U8421 ( .A(n7731), .B(n7730), .Z(n7735) );
  NANDN U8422 ( .A(n7733), .B(n7732), .Z(n7734) );
  AND U8423 ( .A(n7735), .B(n7734), .Z(n7882) );
  NANDN U8424 ( .A(n7737), .B(n7736), .Z(n7741) );
  NANDN U8425 ( .A(n7739), .B(n7738), .Z(n7740) );
  AND U8426 ( .A(n7741), .B(n7740), .Z(n7880) );
  NANDN U8427 ( .A(n7743), .B(n7742), .Z(n7747) );
  NANDN U8428 ( .A(n7745), .B(n7744), .Z(n7746) );
  AND U8429 ( .A(n7747), .B(n7746), .Z(n7892) );
  NANDN U8430 ( .A(n7749), .B(n7748), .Z(n7753) );
  NAND U8431 ( .A(n7751), .B(n7750), .Z(n7752) );
  AND U8432 ( .A(n7753), .B(n7752), .Z(n7891) );
  XNOR U8433 ( .A(n7892), .B(n7891), .Z(n7894) );
  NANDN U8434 ( .A(n7755), .B(n7754), .Z(n7759) );
  NANDN U8435 ( .A(n7757), .B(n7756), .Z(n7758) );
  AND U8436 ( .A(n7759), .B(n7758), .Z(n7969) );
  NAND U8437 ( .A(n38385), .B(n7760), .Z(n7762) );
  XOR U8438 ( .A(b[27]), .B(a[41]), .Z(n7915) );
  NAND U8439 ( .A(n38343), .B(n7915), .Z(n7761) );
  AND U8440 ( .A(n7762), .B(n7761), .Z(n7976) );
  NAND U8441 ( .A(n183), .B(n7763), .Z(n7765) );
  XOR U8442 ( .A(b[5]), .B(a[63]), .Z(n7918) );
  NAND U8443 ( .A(n36296), .B(n7918), .Z(n7764) );
  AND U8444 ( .A(n7765), .B(n7764), .Z(n7974) );
  NAND U8445 ( .A(n190), .B(n7766), .Z(n7768) );
  XOR U8446 ( .A(b[19]), .B(a[49]), .Z(n7921) );
  NAND U8447 ( .A(n37821), .B(n7921), .Z(n7767) );
  NAND U8448 ( .A(n7768), .B(n7767), .Z(n7973) );
  XNOR U8449 ( .A(n7974), .B(n7973), .Z(n7975) );
  XNOR U8450 ( .A(n7976), .B(n7975), .Z(n7967) );
  NAND U8451 ( .A(n38470), .B(n7769), .Z(n7771) );
  XOR U8452 ( .A(b[31]), .B(a[37]), .Z(n7924) );
  NAND U8453 ( .A(n38453), .B(n7924), .Z(n7770) );
  AND U8454 ( .A(n7771), .B(n7770), .Z(n7936) );
  NAND U8455 ( .A(n181), .B(n7772), .Z(n7774) );
  XOR U8456 ( .A(b[3]), .B(a[65]), .Z(n7927) );
  NAND U8457 ( .A(n182), .B(n7927), .Z(n7773) );
  AND U8458 ( .A(n7774), .B(n7773), .Z(n7934) );
  NAND U8459 ( .A(n189), .B(n7775), .Z(n7777) );
  XOR U8460 ( .A(b[17]), .B(a[51]), .Z(n7930) );
  NAND U8461 ( .A(n37652), .B(n7930), .Z(n7776) );
  NAND U8462 ( .A(n7777), .B(n7776), .Z(n7933) );
  XNOR U8463 ( .A(n7934), .B(n7933), .Z(n7935) );
  XOR U8464 ( .A(n7936), .B(n7935), .Z(n7968) );
  XOR U8465 ( .A(n7967), .B(n7968), .Z(n7970) );
  XOR U8466 ( .A(n7969), .B(n7970), .Z(n7904) );
  NANDN U8467 ( .A(n7779), .B(n7778), .Z(n7783) );
  NANDN U8468 ( .A(n7781), .B(n7780), .Z(n7782) );
  AND U8469 ( .A(n7783), .B(n7782), .Z(n7957) );
  NANDN U8470 ( .A(n7785), .B(n7784), .Z(n7789) );
  NANDN U8471 ( .A(n7787), .B(n7786), .Z(n7788) );
  NAND U8472 ( .A(n7789), .B(n7788), .Z(n7958) );
  XNOR U8473 ( .A(n7957), .B(n7958), .Z(n7959) );
  NANDN U8474 ( .A(n7791), .B(n7790), .Z(n7795) );
  NANDN U8475 ( .A(n7793), .B(n7792), .Z(n7794) );
  NAND U8476 ( .A(n7795), .B(n7794), .Z(n7960) );
  XNOR U8477 ( .A(n7959), .B(n7960), .Z(n7903) );
  XNOR U8478 ( .A(n7904), .B(n7903), .Z(n7906) );
  NANDN U8479 ( .A(n7797), .B(n7796), .Z(n7801) );
  NANDN U8480 ( .A(n7799), .B(n7798), .Z(n7800) );
  AND U8481 ( .A(n7801), .B(n7800), .Z(n7905) );
  XOR U8482 ( .A(n7906), .B(n7905), .Z(n8018) );
  NANDN U8483 ( .A(n7803), .B(n7802), .Z(n7807) );
  NANDN U8484 ( .A(n7805), .B(n7804), .Z(n7806) );
  AND U8485 ( .A(n7807), .B(n7806), .Z(n8015) );
  NANDN U8486 ( .A(n7809), .B(n7808), .Z(n7813) );
  NANDN U8487 ( .A(n7811), .B(n7810), .Z(n7812) );
  AND U8488 ( .A(n7813), .B(n7812), .Z(n7900) );
  NANDN U8489 ( .A(n7815), .B(n7814), .Z(n7819) );
  OR U8490 ( .A(n7817), .B(n7816), .Z(n7818) );
  AND U8491 ( .A(n7819), .B(n7818), .Z(n7898) );
  NANDN U8492 ( .A(n7821), .B(n7820), .Z(n7825) );
  NANDN U8493 ( .A(n7823), .B(n7822), .Z(n7824) );
  AND U8494 ( .A(n7825), .B(n7824), .Z(n7964) );
  NANDN U8495 ( .A(n7827), .B(n7826), .Z(n7831) );
  NANDN U8496 ( .A(n7829), .B(n7828), .Z(n7830) );
  NAND U8497 ( .A(n7831), .B(n7830), .Z(n7963) );
  XNOR U8498 ( .A(n7964), .B(n7963), .Z(n7966) );
  NAND U8499 ( .A(n194), .B(n7832), .Z(n7834) );
  XOR U8500 ( .A(b[29]), .B(a[39]), .Z(n7988) );
  NAND U8501 ( .A(n38456), .B(n7988), .Z(n7833) );
  AND U8502 ( .A(n7834), .B(n7833), .Z(n7910) );
  AND U8503 ( .A(b[31]), .B(a[35]), .Z(n7909) );
  XNOR U8504 ( .A(n7910), .B(n7909), .Z(n7911) );
  NAND U8505 ( .A(b[0]), .B(a[67]), .Z(n7835) );
  XNOR U8506 ( .A(b[1]), .B(n7835), .Z(n7837) );
  NANDN U8507 ( .A(b[0]), .B(a[66]), .Z(n7836) );
  NAND U8508 ( .A(n7837), .B(n7836), .Z(n7912) );
  XNOR U8509 ( .A(n7911), .B(n7912), .Z(n7952) );
  NAND U8510 ( .A(n38185), .B(n7838), .Z(n7840) );
  XOR U8511 ( .A(b[23]), .B(a[45]), .Z(n7991) );
  NAND U8512 ( .A(n38132), .B(n7991), .Z(n7839) );
  AND U8513 ( .A(n7840), .B(n7839), .Z(n7981) );
  NAND U8514 ( .A(n184), .B(n7841), .Z(n7843) );
  XOR U8515 ( .A(b[7]), .B(a[61]), .Z(n7994) );
  NAND U8516 ( .A(n36592), .B(n7994), .Z(n7842) );
  AND U8517 ( .A(n7843), .B(n7842), .Z(n7980) );
  NAND U8518 ( .A(n38289), .B(n7844), .Z(n7846) );
  XOR U8519 ( .A(b[25]), .B(a[43]), .Z(n7997) );
  NAND U8520 ( .A(n38247), .B(n7997), .Z(n7845) );
  NAND U8521 ( .A(n7846), .B(n7845), .Z(n7979) );
  XOR U8522 ( .A(n7980), .B(n7979), .Z(n7982) );
  XOR U8523 ( .A(n7981), .B(n7982), .Z(n7951) );
  XOR U8524 ( .A(n7952), .B(n7951), .Z(n7954) );
  NAND U8525 ( .A(n187), .B(n7847), .Z(n7849) );
  XOR U8526 ( .A(b[13]), .B(a[55]), .Z(n8000) );
  NAND U8527 ( .A(n37295), .B(n8000), .Z(n7848) );
  AND U8528 ( .A(n7849), .B(n7848), .Z(n7946) );
  NAND U8529 ( .A(n186), .B(n7850), .Z(n7852) );
  XOR U8530 ( .A(b[11]), .B(a[57]), .Z(n8003) );
  NAND U8531 ( .A(n37097), .B(n8003), .Z(n7851) );
  NAND U8532 ( .A(n7852), .B(n7851), .Z(n7945) );
  XNOR U8533 ( .A(n7946), .B(n7945), .Z(n7948) );
  NAND U8534 ( .A(n188), .B(n7853), .Z(n7855) );
  XOR U8535 ( .A(b[15]), .B(a[53]), .Z(n8006) );
  NAND U8536 ( .A(n37382), .B(n8006), .Z(n7854) );
  AND U8537 ( .A(n7855), .B(n7854), .Z(n7942) );
  NAND U8538 ( .A(n38064), .B(n7856), .Z(n7858) );
  XOR U8539 ( .A(b[21]), .B(a[47]), .Z(n8009) );
  NAND U8540 ( .A(n37993), .B(n8009), .Z(n7857) );
  AND U8541 ( .A(n7858), .B(n7857), .Z(n7940) );
  NAND U8542 ( .A(n185), .B(n7859), .Z(n7861) );
  XOR U8543 ( .A(b[9]), .B(a[59]), .Z(n8012) );
  NAND U8544 ( .A(n36805), .B(n8012), .Z(n7860) );
  NAND U8545 ( .A(n7861), .B(n7860), .Z(n7939) );
  XNOR U8546 ( .A(n7940), .B(n7939), .Z(n7941) );
  XNOR U8547 ( .A(n7942), .B(n7941), .Z(n7947) );
  XOR U8548 ( .A(n7948), .B(n7947), .Z(n7953) );
  XNOR U8549 ( .A(n7954), .B(n7953), .Z(n7965) );
  XNOR U8550 ( .A(n7966), .B(n7965), .Z(n7897) );
  XNOR U8551 ( .A(n7898), .B(n7897), .Z(n7899) );
  XOR U8552 ( .A(n7900), .B(n7899), .Z(n8016) );
  XNOR U8553 ( .A(n8015), .B(n8016), .Z(n8017) );
  XNOR U8554 ( .A(n8018), .B(n8017), .Z(n7893) );
  XOR U8555 ( .A(n7894), .B(n7893), .Z(n7886) );
  NANDN U8556 ( .A(n7863), .B(n7862), .Z(n7867) );
  NANDN U8557 ( .A(n7865), .B(n7864), .Z(n7866) );
  AND U8558 ( .A(n7867), .B(n7866), .Z(n7885) );
  XNOR U8559 ( .A(n7886), .B(n7885), .Z(n7887) );
  NANDN U8560 ( .A(n7869), .B(n7868), .Z(n7873) );
  NAND U8561 ( .A(n7871), .B(n7870), .Z(n7872) );
  NAND U8562 ( .A(n7873), .B(n7872), .Z(n7888) );
  XNOR U8563 ( .A(n7887), .B(n7888), .Z(n7879) );
  XNOR U8564 ( .A(n7880), .B(n7879), .Z(n7881) );
  XNOR U8565 ( .A(n7882), .B(n7881), .Z(n8021) );
  XNOR U8566 ( .A(sreg[291]), .B(n8021), .Z(n8023) );
  NANDN U8567 ( .A(sreg[290]), .B(n7874), .Z(n7878) );
  NAND U8568 ( .A(n7876), .B(n7875), .Z(n7877) );
  NAND U8569 ( .A(n7878), .B(n7877), .Z(n8022) );
  XNOR U8570 ( .A(n8023), .B(n8022), .Z(c[291]) );
  NANDN U8571 ( .A(n7880), .B(n7879), .Z(n7884) );
  NANDN U8572 ( .A(n7882), .B(n7881), .Z(n7883) );
  AND U8573 ( .A(n7884), .B(n7883), .Z(n8029) );
  NANDN U8574 ( .A(n7886), .B(n7885), .Z(n7890) );
  NANDN U8575 ( .A(n7888), .B(n7887), .Z(n7889) );
  AND U8576 ( .A(n7890), .B(n7889), .Z(n8027) );
  NANDN U8577 ( .A(n7892), .B(n7891), .Z(n7896) );
  NAND U8578 ( .A(n7894), .B(n7893), .Z(n7895) );
  AND U8579 ( .A(n7896), .B(n7895), .Z(n8034) );
  NANDN U8580 ( .A(n7898), .B(n7897), .Z(n7902) );
  NANDN U8581 ( .A(n7900), .B(n7899), .Z(n7901) );
  AND U8582 ( .A(n7902), .B(n7901), .Z(n8165) );
  NANDN U8583 ( .A(n7904), .B(n7903), .Z(n7908) );
  NAND U8584 ( .A(n7906), .B(n7905), .Z(n7907) );
  AND U8585 ( .A(n7908), .B(n7907), .Z(n8164) );
  XNOR U8586 ( .A(n8165), .B(n8164), .Z(n8167) );
  NANDN U8587 ( .A(n7910), .B(n7909), .Z(n7914) );
  NANDN U8588 ( .A(n7912), .B(n7911), .Z(n7913) );
  AND U8589 ( .A(n7914), .B(n7913), .Z(n8100) );
  NAND U8590 ( .A(n38385), .B(n7915), .Z(n7917) );
  XOR U8591 ( .A(b[27]), .B(a[42]), .Z(n8044) );
  NAND U8592 ( .A(n38343), .B(n8044), .Z(n7916) );
  AND U8593 ( .A(n7917), .B(n7916), .Z(n8107) );
  NAND U8594 ( .A(n183), .B(n7918), .Z(n7920) );
  XOR U8595 ( .A(b[5]), .B(a[64]), .Z(n8047) );
  NAND U8596 ( .A(n36296), .B(n8047), .Z(n7919) );
  AND U8597 ( .A(n7920), .B(n7919), .Z(n8105) );
  NAND U8598 ( .A(n190), .B(n7921), .Z(n7923) );
  XOR U8599 ( .A(b[19]), .B(a[50]), .Z(n8050) );
  NAND U8600 ( .A(n37821), .B(n8050), .Z(n7922) );
  NAND U8601 ( .A(n7923), .B(n7922), .Z(n8104) );
  XNOR U8602 ( .A(n8105), .B(n8104), .Z(n8106) );
  XNOR U8603 ( .A(n8107), .B(n8106), .Z(n8098) );
  NAND U8604 ( .A(n38470), .B(n7924), .Z(n7926) );
  XOR U8605 ( .A(b[31]), .B(a[38]), .Z(n8053) );
  NAND U8606 ( .A(n38453), .B(n8053), .Z(n7925) );
  AND U8607 ( .A(n7926), .B(n7925), .Z(n8065) );
  NAND U8608 ( .A(n181), .B(n7927), .Z(n7929) );
  XOR U8609 ( .A(b[3]), .B(a[66]), .Z(n8056) );
  NAND U8610 ( .A(n182), .B(n8056), .Z(n7928) );
  AND U8611 ( .A(n7929), .B(n7928), .Z(n8063) );
  NAND U8612 ( .A(n189), .B(n7930), .Z(n7932) );
  XOR U8613 ( .A(b[17]), .B(a[52]), .Z(n8059) );
  NAND U8614 ( .A(n37652), .B(n8059), .Z(n7931) );
  NAND U8615 ( .A(n7932), .B(n7931), .Z(n8062) );
  XNOR U8616 ( .A(n8063), .B(n8062), .Z(n8064) );
  XOR U8617 ( .A(n8065), .B(n8064), .Z(n8099) );
  XOR U8618 ( .A(n8098), .B(n8099), .Z(n8101) );
  XOR U8619 ( .A(n8100), .B(n8101), .Z(n8147) );
  NANDN U8620 ( .A(n7934), .B(n7933), .Z(n7938) );
  NANDN U8621 ( .A(n7936), .B(n7935), .Z(n7937) );
  AND U8622 ( .A(n7938), .B(n7937), .Z(n8086) );
  NANDN U8623 ( .A(n7940), .B(n7939), .Z(n7944) );
  NANDN U8624 ( .A(n7942), .B(n7941), .Z(n7943) );
  NAND U8625 ( .A(n7944), .B(n7943), .Z(n8087) );
  XNOR U8626 ( .A(n8086), .B(n8087), .Z(n8088) );
  NANDN U8627 ( .A(n7946), .B(n7945), .Z(n7950) );
  NAND U8628 ( .A(n7948), .B(n7947), .Z(n7949) );
  NAND U8629 ( .A(n7950), .B(n7949), .Z(n8089) );
  XNOR U8630 ( .A(n8088), .B(n8089), .Z(n8146) );
  XNOR U8631 ( .A(n8147), .B(n8146), .Z(n8149) );
  NAND U8632 ( .A(n7952), .B(n7951), .Z(n7956) );
  NAND U8633 ( .A(n7954), .B(n7953), .Z(n7955) );
  AND U8634 ( .A(n7956), .B(n7955), .Z(n8148) );
  XOR U8635 ( .A(n8149), .B(n8148), .Z(n8161) );
  NANDN U8636 ( .A(n7958), .B(n7957), .Z(n7962) );
  NANDN U8637 ( .A(n7960), .B(n7959), .Z(n7961) );
  AND U8638 ( .A(n7962), .B(n7961), .Z(n8158) );
  NANDN U8639 ( .A(n7968), .B(n7967), .Z(n7972) );
  OR U8640 ( .A(n7970), .B(n7969), .Z(n7971) );
  AND U8641 ( .A(n7972), .B(n7971), .Z(n8153) );
  NANDN U8642 ( .A(n7974), .B(n7973), .Z(n7978) );
  NANDN U8643 ( .A(n7976), .B(n7975), .Z(n7977) );
  AND U8644 ( .A(n7978), .B(n7977), .Z(n8093) );
  NANDN U8645 ( .A(n7980), .B(n7979), .Z(n7984) );
  OR U8646 ( .A(n7982), .B(n7981), .Z(n7983) );
  NAND U8647 ( .A(n7984), .B(n7983), .Z(n8092) );
  XNOR U8648 ( .A(n8093), .B(n8092), .Z(n8094) );
  NAND U8649 ( .A(b[0]), .B(a[68]), .Z(n7985) );
  XNOR U8650 ( .A(b[1]), .B(n7985), .Z(n7987) );
  NANDN U8651 ( .A(b[0]), .B(a[67]), .Z(n7986) );
  NAND U8652 ( .A(n7987), .B(n7986), .Z(n8041) );
  NAND U8653 ( .A(n194), .B(n7988), .Z(n7990) );
  XOR U8654 ( .A(b[29]), .B(a[40]), .Z(n8116) );
  NAND U8655 ( .A(n38456), .B(n8116), .Z(n7989) );
  AND U8656 ( .A(n7990), .B(n7989), .Z(n8039) );
  AND U8657 ( .A(b[31]), .B(a[36]), .Z(n8038) );
  XNOR U8658 ( .A(n8039), .B(n8038), .Z(n8040) );
  XNOR U8659 ( .A(n8041), .B(n8040), .Z(n8080) );
  NAND U8660 ( .A(n38185), .B(n7991), .Z(n7993) );
  XOR U8661 ( .A(b[23]), .B(a[46]), .Z(n8122) );
  NAND U8662 ( .A(n38132), .B(n8122), .Z(n7992) );
  AND U8663 ( .A(n7993), .B(n7992), .Z(n8113) );
  NAND U8664 ( .A(n184), .B(n7994), .Z(n7996) );
  XOR U8665 ( .A(b[7]), .B(a[62]), .Z(n8125) );
  NAND U8666 ( .A(n36592), .B(n8125), .Z(n7995) );
  AND U8667 ( .A(n7996), .B(n7995), .Z(n8111) );
  NAND U8668 ( .A(n38289), .B(n7997), .Z(n7999) );
  XOR U8669 ( .A(b[25]), .B(a[44]), .Z(n8128) );
  NAND U8670 ( .A(n38247), .B(n8128), .Z(n7998) );
  NAND U8671 ( .A(n7999), .B(n7998), .Z(n8110) );
  XNOR U8672 ( .A(n8111), .B(n8110), .Z(n8112) );
  XOR U8673 ( .A(n8113), .B(n8112), .Z(n8081) );
  XNOR U8674 ( .A(n8080), .B(n8081), .Z(n8082) );
  NAND U8675 ( .A(n187), .B(n8000), .Z(n8002) );
  XOR U8676 ( .A(b[13]), .B(a[56]), .Z(n8131) );
  NAND U8677 ( .A(n37295), .B(n8131), .Z(n8001) );
  AND U8678 ( .A(n8002), .B(n8001), .Z(n8075) );
  NAND U8679 ( .A(n186), .B(n8003), .Z(n8005) );
  XOR U8680 ( .A(b[11]), .B(a[58]), .Z(n8134) );
  NAND U8681 ( .A(n37097), .B(n8134), .Z(n8004) );
  NAND U8682 ( .A(n8005), .B(n8004), .Z(n8074) );
  XNOR U8683 ( .A(n8075), .B(n8074), .Z(n8076) );
  NAND U8684 ( .A(n188), .B(n8006), .Z(n8008) );
  XOR U8685 ( .A(b[15]), .B(a[54]), .Z(n8137) );
  NAND U8686 ( .A(n37382), .B(n8137), .Z(n8007) );
  AND U8687 ( .A(n8008), .B(n8007), .Z(n8071) );
  NAND U8688 ( .A(n38064), .B(n8009), .Z(n8011) );
  XOR U8689 ( .A(b[21]), .B(a[48]), .Z(n8140) );
  NAND U8690 ( .A(n37993), .B(n8140), .Z(n8010) );
  AND U8691 ( .A(n8011), .B(n8010), .Z(n8069) );
  NAND U8692 ( .A(n185), .B(n8012), .Z(n8014) );
  XOR U8693 ( .A(b[9]), .B(a[60]), .Z(n8143) );
  NAND U8694 ( .A(n36805), .B(n8143), .Z(n8013) );
  NAND U8695 ( .A(n8014), .B(n8013), .Z(n8068) );
  XNOR U8696 ( .A(n8069), .B(n8068), .Z(n8070) );
  XOR U8697 ( .A(n8071), .B(n8070), .Z(n8077) );
  XOR U8698 ( .A(n8076), .B(n8077), .Z(n8083) );
  XOR U8699 ( .A(n8082), .B(n8083), .Z(n8095) );
  XNOR U8700 ( .A(n8094), .B(n8095), .Z(n8152) );
  XNOR U8701 ( .A(n8153), .B(n8152), .Z(n8154) );
  XOR U8702 ( .A(n8155), .B(n8154), .Z(n8159) );
  XNOR U8703 ( .A(n8158), .B(n8159), .Z(n8160) );
  XNOR U8704 ( .A(n8161), .B(n8160), .Z(n8166) );
  XOR U8705 ( .A(n8167), .B(n8166), .Z(n8033) );
  NANDN U8706 ( .A(n8016), .B(n8015), .Z(n8020) );
  NANDN U8707 ( .A(n8018), .B(n8017), .Z(n8019) );
  AND U8708 ( .A(n8020), .B(n8019), .Z(n8032) );
  XOR U8709 ( .A(n8033), .B(n8032), .Z(n8035) );
  XNOR U8710 ( .A(n8034), .B(n8035), .Z(n8026) );
  XNOR U8711 ( .A(n8027), .B(n8026), .Z(n8028) );
  XNOR U8712 ( .A(n8029), .B(n8028), .Z(n8170) );
  XNOR U8713 ( .A(sreg[292]), .B(n8170), .Z(n8172) );
  NANDN U8714 ( .A(sreg[291]), .B(n8021), .Z(n8025) );
  NAND U8715 ( .A(n8023), .B(n8022), .Z(n8024) );
  NAND U8716 ( .A(n8025), .B(n8024), .Z(n8171) );
  XNOR U8717 ( .A(n8172), .B(n8171), .Z(c[292]) );
  NANDN U8718 ( .A(n8027), .B(n8026), .Z(n8031) );
  NANDN U8719 ( .A(n8029), .B(n8028), .Z(n8030) );
  AND U8720 ( .A(n8031), .B(n8030), .Z(n8178) );
  NANDN U8721 ( .A(n8033), .B(n8032), .Z(n8037) );
  NANDN U8722 ( .A(n8035), .B(n8034), .Z(n8036) );
  AND U8723 ( .A(n8037), .B(n8036), .Z(n8176) );
  NANDN U8724 ( .A(n8039), .B(n8038), .Z(n8043) );
  NANDN U8725 ( .A(n8041), .B(n8040), .Z(n8042) );
  AND U8726 ( .A(n8043), .B(n8042), .Z(n8267) );
  NAND U8727 ( .A(n38385), .B(n8044), .Z(n8046) );
  XOR U8728 ( .A(b[27]), .B(a[43]), .Z(n8211) );
  NAND U8729 ( .A(n38343), .B(n8211), .Z(n8045) );
  AND U8730 ( .A(n8046), .B(n8045), .Z(n8274) );
  NAND U8731 ( .A(n183), .B(n8047), .Z(n8049) );
  XOR U8732 ( .A(b[5]), .B(a[65]), .Z(n8214) );
  NAND U8733 ( .A(n36296), .B(n8214), .Z(n8048) );
  AND U8734 ( .A(n8049), .B(n8048), .Z(n8272) );
  NAND U8735 ( .A(n190), .B(n8050), .Z(n8052) );
  XOR U8736 ( .A(b[19]), .B(a[51]), .Z(n8217) );
  NAND U8737 ( .A(n37821), .B(n8217), .Z(n8051) );
  NAND U8738 ( .A(n8052), .B(n8051), .Z(n8271) );
  XNOR U8739 ( .A(n8272), .B(n8271), .Z(n8273) );
  XNOR U8740 ( .A(n8274), .B(n8273), .Z(n8265) );
  NAND U8741 ( .A(n38470), .B(n8053), .Z(n8055) );
  XOR U8742 ( .A(b[31]), .B(a[39]), .Z(n8220) );
  NAND U8743 ( .A(n38453), .B(n8220), .Z(n8054) );
  AND U8744 ( .A(n8055), .B(n8054), .Z(n8232) );
  NAND U8745 ( .A(n181), .B(n8056), .Z(n8058) );
  XOR U8746 ( .A(b[3]), .B(a[67]), .Z(n8223) );
  NAND U8747 ( .A(n182), .B(n8223), .Z(n8057) );
  AND U8748 ( .A(n8058), .B(n8057), .Z(n8230) );
  NAND U8749 ( .A(n189), .B(n8059), .Z(n8061) );
  XOR U8750 ( .A(b[17]), .B(a[53]), .Z(n8226) );
  NAND U8751 ( .A(n37652), .B(n8226), .Z(n8060) );
  NAND U8752 ( .A(n8061), .B(n8060), .Z(n8229) );
  XNOR U8753 ( .A(n8230), .B(n8229), .Z(n8231) );
  XOR U8754 ( .A(n8232), .B(n8231), .Z(n8266) );
  XOR U8755 ( .A(n8265), .B(n8266), .Z(n8268) );
  XOR U8756 ( .A(n8267), .B(n8268), .Z(n8200) );
  NANDN U8757 ( .A(n8063), .B(n8062), .Z(n8067) );
  NANDN U8758 ( .A(n8065), .B(n8064), .Z(n8066) );
  AND U8759 ( .A(n8067), .B(n8066), .Z(n8253) );
  NANDN U8760 ( .A(n8069), .B(n8068), .Z(n8073) );
  NANDN U8761 ( .A(n8071), .B(n8070), .Z(n8072) );
  NAND U8762 ( .A(n8073), .B(n8072), .Z(n8254) );
  XNOR U8763 ( .A(n8253), .B(n8254), .Z(n8255) );
  NANDN U8764 ( .A(n8075), .B(n8074), .Z(n8079) );
  NANDN U8765 ( .A(n8077), .B(n8076), .Z(n8078) );
  NAND U8766 ( .A(n8079), .B(n8078), .Z(n8256) );
  XNOR U8767 ( .A(n8255), .B(n8256), .Z(n8199) );
  XNOR U8768 ( .A(n8200), .B(n8199), .Z(n8202) );
  NANDN U8769 ( .A(n8081), .B(n8080), .Z(n8085) );
  NANDN U8770 ( .A(n8083), .B(n8082), .Z(n8084) );
  AND U8771 ( .A(n8085), .B(n8084), .Z(n8201) );
  XOR U8772 ( .A(n8202), .B(n8201), .Z(n8315) );
  NANDN U8773 ( .A(n8087), .B(n8086), .Z(n8091) );
  NANDN U8774 ( .A(n8089), .B(n8088), .Z(n8090) );
  AND U8775 ( .A(n8091), .B(n8090), .Z(n8313) );
  NANDN U8776 ( .A(n8093), .B(n8092), .Z(n8097) );
  NANDN U8777 ( .A(n8095), .B(n8094), .Z(n8096) );
  AND U8778 ( .A(n8097), .B(n8096), .Z(n8196) );
  NANDN U8779 ( .A(n8099), .B(n8098), .Z(n8103) );
  OR U8780 ( .A(n8101), .B(n8100), .Z(n8102) );
  AND U8781 ( .A(n8103), .B(n8102), .Z(n8194) );
  NANDN U8782 ( .A(n8105), .B(n8104), .Z(n8109) );
  NANDN U8783 ( .A(n8107), .B(n8106), .Z(n8108) );
  AND U8784 ( .A(n8109), .B(n8108), .Z(n8260) );
  NANDN U8785 ( .A(n8111), .B(n8110), .Z(n8115) );
  NANDN U8786 ( .A(n8113), .B(n8112), .Z(n8114) );
  NAND U8787 ( .A(n8115), .B(n8114), .Z(n8259) );
  XNOR U8788 ( .A(n8260), .B(n8259), .Z(n8261) );
  NAND U8789 ( .A(n194), .B(n8116), .Z(n8118) );
  XOR U8790 ( .A(b[29]), .B(a[41]), .Z(n8286) );
  NAND U8791 ( .A(n38456), .B(n8286), .Z(n8117) );
  AND U8792 ( .A(n8118), .B(n8117), .Z(n8206) );
  AND U8793 ( .A(b[31]), .B(a[37]), .Z(n8205) );
  XNOR U8794 ( .A(n8206), .B(n8205), .Z(n8207) );
  NAND U8795 ( .A(b[0]), .B(a[69]), .Z(n8119) );
  XNOR U8796 ( .A(b[1]), .B(n8119), .Z(n8121) );
  NANDN U8797 ( .A(b[0]), .B(a[68]), .Z(n8120) );
  NAND U8798 ( .A(n8121), .B(n8120), .Z(n8208) );
  XNOR U8799 ( .A(n8207), .B(n8208), .Z(n8247) );
  NAND U8800 ( .A(n38185), .B(n8122), .Z(n8124) );
  XOR U8801 ( .A(b[23]), .B(a[47]), .Z(n8289) );
  NAND U8802 ( .A(n38132), .B(n8289), .Z(n8123) );
  AND U8803 ( .A(n8124), .B(n8123), .Z(n8280) );
  NAND U8804 ( .A(n184), .B(n8125), .Z(n8127) );
  XOR U8805 ( .A(b[7]), .B(a[63]), .Z(n8292) );
  NAND U8806 ( .A(n36592), .B(n8292), .Z(n8126) );
  AND U8807 ( .A(n8127), .B(n8126), .Z(n8278) );
  NAND U8808 ( .A(n38289), .B(n8128), .Z(n8130) );
  XOR U8809 ( .A(b[25]), .B(a[45]), .Z(n8295) );
  NAND U8810 ( .A(n38247), .B(n8295), .Z(n8129) );
  NAND U8811 ( .A(n8130), .B(n8129), .Z(n8277) );
  XNOR U8812 ( .A(n8278), .B(n8277), .Z(n8279) );
  XOR U8813 ( .A(n8280), .B(n8279), .Z(n8248) );
  XNOR U8814 ( .A(n8247), .B(n8248), .Z(n8249) );
  NAND U8815 ( .A(n187), .B(n8131), .Z(n8133) );
  XOR U8816 ( .A(b[13]), .B(a[57]), .Z(n8298) );
  NAND U8817 ( .A(n37295), .B(n8298), .Z(n8132) );
  AND U8818 ( .A(n8133), .B(n8132), .Z(n8242) );
  NAND U8819 ( .A(n186), .B(n8134), .Z(n8136) );
  XOR U8820 ( .A(b[11]), .B(a[59]), .Z(n8301) );
  NAND U8821 ( .A(n37097), .B(n8301), .Z(n8135) );
  NAND U8822 ( .A(n8136), .B(n8135), .Z(n8241) );
  XNOR U8823 ( .A(n8242), .B(n8241), .Z(n8243) );
  NAND U8824 ( .A(n188), .B(n8137), .Z(n8139) );
  XOR U8825 ( .A(b[15]), .B(a[55]), .Z(n8304) );
  NAND U8826 ( .A(n37382), .B(n8304), .Z(n8138) );
  AND U8827 ( .A(n8139), .B(n8138), .Z(n8238) );
  NAND U8828 ( .A(n38064), .B(n8140), .Z(n8142) );
  XOR U8829 ( .A(b[21]), .B(a[49]), .Z(n8307) );
  NAND U8830 ( .A(n37993), .B(n8307), .Z(n8141) );
  AND U8831 ( .A(n8142), .B(n8141), .Z(n8236) );
  NAND U8832 ( .A(n185), .B(n8143), .Z(n8145) );
  XOR U8833 ( .A(b[9]), .B(a[61]), .Z(n8310) );
  NAND U8834 ( .A(n36805), .B(n8310), .Z(n8144) );
  NAND U8835 ( .A(n8145), .B(n8144), .Z(n8235) );
  XNOR U8836 ( .A(n8236), .B(n8235), .Z(n8237) );
  XOR U8837 ( .A(n8238), .B(n8237), .Z(n8244) );
  XOR U8838 ( .A(n8243), .B(n8244), .Z(n8250) );
  XOR U8839 ( .A(n8249), .B(n8250), .Z(n8262) );
  XNOR U8840 ( .A(n8261), .B(n8262), .Z(n8193) );
  XNOR U8841 ( .A(n8194), .B(n8193), .Z(n8195) );
  XOR U8842 ( .A(n8196), .B(n8195), .Z(n8314) );
  XOR U8843 ( .A(n8313), .B(n8314), .Z(n8316) );
  XOR U8844 ( .A(n8315), .B(n8316), .Z(n8190) );
  NANDN U8845 ( .A(n8147), .B(n8146), .Z(n8151) );
  NAND U8846 ( .A(n8149), .B(n8148), .Z(n8150) );
  AND U8847 ( .A(n8151), .B(n8150), .Z(n8188) );
  NANDN U8848 ( .A(n8153), .B(n8152), .Z(n8157) );
  NANDN U8849 ( .A(n8155), .B(n8154), .Z(n8156) );
  AND U8850 ( .A(n8157), .B(n8156), .Z(n8187) );
  XNOR U8851 ( .A(n8188), .B(n8187), .Z(n8189) );
  XNOR U8852 ( .A(n8190), .B(n8189), .Z(n8181) );
  NANDN U8853 ( .A(n8159), .B(n8158), .Z(n8163) );
  NANDN U8854 ( .A(n8161), .B(n8160), .Z(n8162) );
  NAND U8855 ( .A(n8163), .B(n8162), .Z(n8182) );
  XNOR U8856 ( .A(n8181), .B(n8182), .Z(n8183) );
  NANDN U8857 ( .A(n8165), .B(n8164), .Z(n8169) );
  NAND U8858 ( .A(n8167), .B(n8166), .Z(n8168) );
  NAND U8859 ( .A(n8169), .B(n8168), .Z(n8184) );
  XNOR U8860 ( .A(n8183), .B(n8184), .Z(n8175) );
  XNOR U8861 ( .A(n8176), .B(n8175), .Z(n8177) );
  XNOR U8862 ( .A(n8178), .B(n8177), .Z(n8319) );
  XNOR U8863 ( .A(sreg[293]), .B(n8319), .Z(n8321) );
  NANDN U8864 ( .A(sreg[292]), .B(n8170), .Z(n8174) );
  NAND U8865 ( .A(n8172), .B(n8171), .Z(n8173) );
  NAND U8866 ( .A(n8174), .B(n8173), .Z(n8320) );
  XNOR U8867 ( .A(n8321), .B(n8320), .Z(c[293]) );
  NANDN U8868 ( .A(n8176), .B(n8175), .Z(n8180) );
  NANDN U8869 ( .A(n8178), .B(n8177), .Z(n8179) );
  AND U8870 ( .A(n8180), .B(n8179), .Z(n8327) );
  NANDN U8871 ( .A(n8182), .B(n8181), .Z(n8186) );
  NANDN U8872 ( .A(n8184), .B(n8183), .Z(n8185) );
  AND U8873 ( .A(n8186), .B(n8185), .Z(n8325) );
  NANDN U8874 ( .A(n8188), .B(n8187), .Z(n8192) );
  NANDN U8875 ( .A(n8190), .B(n8189), .Z(n8191) );
  AND U8876 ( .A(n8192), .B(n8191), .Z(n8333) );
  NANDN U8877 ( .A(n8194), .B(n8193), .Z(n8198) );
  NANDN U8878 ( .A(n8196), .B(n8195), .Z(n8197) );
  AND U8879 ( .A(n8198), .B(n8197), .Z(n8337) );
  NANDN U8880 ( .A(n8200), .B(n8199), .Z(n8204) );
  NAND U8881 ( .A(n8202), .B(n8201), .Z(n8203) );
  AND U8882 ( .A(n8204), .B(n8203), .Z(n8336) );
  XNOR U8883 ( .A(n8337), .B(n8336), .Z(n8339) );
  NANDN U8884 ( .A(n8206), .B(n8205), .Z(n8210) );
  NANDN U8885 ( .A(n8208), .B(n8207), .Z(n8209) );
  AND U8886 ( .A(n8210), .B(n8209), .Z(n8416) );
  NAND U8887 ( .A(n38385), .B(n8211), .Z(n8213) );
  XOR U8888 ( .A(b[27]), .B(a[44]), .Z(n8360) );
  NAND U8889 ( .A(n38343), .B(n8360), .Z(n8212) );
  AND U8890 ( .A(n8213), .B(n8212), .Z(n8423) );
  NAND U8891 ( .A(n183), .B(n8214), .Z(n8216) );
  XOR U8892 ( .A(b[5]), .B(a[66]), .Z(n8363) );
  NAND U8893 ( .A(n36296), .B(n8363), .Z(n8215) );
  AND U8894 ( .A(n8216), .B(n8215), .Z(n8421) );
  NAND U8895 ( .A(n190), .B(n8217), .Z(n8219) );
  XOR U8896 ( .A(b[19]), .B(a[52]), .Z(n8366) );
  NAND U8897 ( .A(n37821), .B(n8366), .Z(n8218) );
  NAND U8898 ( .A(n8219), .B(n8218), .Z(n8420) );
  XNOR U8899 ( .A(n8421), .B(n8420), .Z(n8422) );
  XNOR U8900 ( .A(n8423), .B(n8422), .Z(n8414) );
  NAND U8901 ( .A(n38470), .B(n8220), .Z(n8222) );
  XOR U8902 ( .A(b[31]), .B(a[40]), .Z(n8369) );
  NAND U8903 ( .A(n38453), .B(n8369), .Z(n8221) );
  AND U8904 ( .A(n8222), .B(n8221), .Z(n8381) );
  NAND U8905 ( .A(n181), .B(n8223), .Z(n8225) );
  XOR U8906 ( .A(b[3]), .B(a[68]), .Z(n8372) );
  NAND U8907 ( .A(n182), .B(n8372), .Z(n8224) );
  AND U8908 ( .A(n8225), .B(n8224), .Z(n8379) );
  NAND U8909 ( .A(n189), .B(n8226), .Z(n8228) );
  XOR U8910 ( .A(b[17]), .B(a[54]), .Z(n8375) );
  NAND U8911 ( .A(n37652), .B(n8375), .Z(n8227) );
  NAND U8912 ( .A(n8228), .B(n8227), .Z(n8378) );
  XNOR U8913 ( .A(n8379), .B(n8378), .Z(n8380) );
  XOR U8914 ( .A(n8381), .B(n8380), .Z(n8415) );
  XOR U8915 ( .A(n8414), .B(n8415), .Z(n8417) );
  XOR U8916 ( .A(n8416), .B(n8417), .Z(n8349) );
  NANDN U8917 ( .A(n8230), .B(n8229), .Z(n8234) );
  NANDN U8918 ( .A(n8232), .B(n8231), .Z(n8233) );
  AND U8919 ( .A(n8234), .B(n8233), .Z(n8402) );
  NANDN U8920 ( .A(n8236), .B(n8235), .Z(n8240) );
  NANDN U8921 ( .A(n8238), .B(n8237), .Z(n8239) );
  NAND U8922 ( .A(n8240), .B(n8239), .Z(n8403) );
  XNOR U8923 ( .A(n8402), .B(n8403), .Z(n8404) );
  NANDN U8924 ( .A(n8242), .B(n8241), .Z(n8246) );
  NANDN U8925 ( .A(n8244), .B(n8243), .Z(n8245) );
  NAND U8926 ( .A(n8246), .B(n8245), .Z(n8405) );
  XNOR U8927 ( .A(n8404), .B(n8405), .Z(n8348) );
  XNOR U8928 ( .A(n8349), .B(n8348), .Z(n8351) );
  NANDN U8929 ( .A(n8248), .B(n8247), .Z(n8252) );
  NANDN U8930 ( .A(n8250), .B(n8249), .Z(n8251) );
  AND U8931 ( .A(n8252), .B(n8251), .Z(n8350) );
  XOR U8932 ( .A(n8351), .B(n8350), .Z(n8465) );
  NANDN U8933 ( .A(n8254), .B(n8253), .Z(n8258) );
  NANDN U8934 ( .A(n8256), .B(n8255), .Z(n8257) );
  AND U8935 ( .A(n8258), .B(n8257), .Z(n8462) );
  NANDN U8936 ( .A(n8260), .B(n8259), .Z(n8264) );
  NANDN U8937 ( .A(n8262), .B(n8261), .Z(n8263) );
  AND U8938 ( .A(n8264), .B(n8263), .Z(n8345) );
  NANDN U8939 ( .A(n8266), .B(n8265), .Z(n8270) );
  OR U8940 ( .A(n8268), .B(n8267), .Z(n8269) );
  AND U8941 ( .A(n8270), .B(n8269), .Z(n8343) );
  NANDN U8942 ( .A(n8272), .B(n8271), .Z(n8276) );
  NANDN U8943 ( .A(n8274), .B(n8273), .Z(n8275) );
  AND U8944 ( .A(n8276), .B(n8275), .Z(n8409) );
  NANDN U8945 ( .A(n8278), .B(n8277), .Z(n8282) );
  NANDN U8946 ( .A(n8280), .B(n8279), .Z(n8281) );
  NAND U8947 ( .A(n8282), .B(n8281), .Z(n8408) );
  XNOR U8948 ( .A(n8409), .B(n8408), .Z(n8410) );
  NAND U8949 ( .A(b[0]), .B(a[70]), .Z(n8283) );
  XNOR U8950 ( .A(b[1]), .B(n8283), .Z(n8285) );
  NANDN U8951 ( .A(b[0]), .B(a[69]), .Z(n8284) );
  NAND U8952 ( .A(n8285), .B(n8284), .Z(n8357) );
  NAND U8953 ( .A(n194), .B(n8286), .Z(n8288) );
  XOR U8954 ( .A(b[29]), .B(a[42]), .Z(n8435) );
  NAND U8955 ( .A(n38456), .B(n8435), .Z(n8287) );
  AND U8956 ( .A(n8288), .B(n8287), .Z(n8355) );
  AND U8957 ( .A(b[31]), .B(a[38]), .Z(n8354) );
  XNOR U8958 ( .A(n8355), .B(n8354), .Z(n8356) );
  XNOR U8959 ( .A(n8357), .B(n8356), .Z(n8396) );
  NAND U8960 ( .A(n38185), .B(n8289), .Z(n8291) );
  XOR U8961 ( .A(b[23]), .B(a[48]), .Z(n8438) );
  NAND U8962 ( .A(n38132), .B(n8438), .Z(n8290) );
  AND U8963 ( .A(n8291), .B(n8290), .Z(n8429) );
  NAND U8964 ( .A(n184), .B(n8292), .Z(n8294) );
  XOR U8965 ( .A(b[7]), .B(a[64]), .Z(n8441) );
  NAND U8966 ( .A(n36592), .B(n8441), .Z(n8293) );
  AND U8967 ( .A(n8294), .B(n8293), .Z(n8427) );
  NAND U8968 ( .A(n38289), .B(n8295), .Z(n8297) );
  XOR U8969 ( .A(b[25]), .B(a[46]), .Z(n8444) );
  NAND U8970 ( .A(n38247), .B(n8444), .Z(n8296) );
  NAND U8971 ( .A(n8297), .B(n8296), .Z(n8426) );
  XNOR U8972 ( .A(n8427), .B(n8426), .Z(n8428) );
  XOR U8973 ( .A(n8429), .B(n8428), .Z(n8397) );
  XNOR U8974 ( .A(n8396), .B(n8397), .Z(n8398) );
  NAND U8975 ( .A(n187), .B(n8298), .Z(n8300) );
  XOR U8976 ( .A(b[13]), .B(a[58]), .Z(n8447) );
  NAND U8977 ( .A(n37295), .B(n8447), .Z(n8299) );
  AND U8978 ( .A(n8300), .B(n8299), .Z(n8391) );
  NAND U8979 ( .A(n186), .B(n8301), .Z(n8303) );
  XOR U8980 ( .A(b[11]), .B(a[60]), .Z(n8450) );
  NAND U8981 ( .A(n37097), .B(n8450), .Z(n8302) );
  NAND U8982 ( .A(n8303), .B(n8302), .Z(n8390) );
  XNOR U8983 ( .A(n8391), .B(n8390), .Z(n8392) );
  NAND U8984 ( .A(n188), .B(n8304), .Z(n8306) );
  XOR U8985 ( .A(b[15]), .B(a[56]), .Z(n8453) );
  NAND U8986 ( .A(n37382), .B(n8453), .Z(n8305) );
  AND U8987 ( .A(n8306), .B(n8305), .Z(n8387) );
  NAND U8988 ( .A(n38064), .B(n8307), .Z(n8309) );
  XOR U8989 ( .A(b[21]), .B(a[50]), .Z(n8456) );
  NAND U8990 ( .A(n37993), .B(n8456), .Z(n8308) );
  AND U8991 ( .A(n8309), .B(n8308), .Z(n8385) );
  NAND U8992 ( .A(n185), .B(n8310), .Z(n8312) );
  XOR U8993 ( .A(b[9]), .B(a[62]), .Z(n8459) );
  NAND U8994 ( .A(n36805), .B(n8459), .Z(n8311) );
  NAND U8995 ( .A(n8312), .B(n8311), .Z(n8384) );
  XNOR U8996 ( .A(n8385), .B(n8384), .Z(n8386) );
  XOR U8997 ( .A(n8387), .B(n8386), .Z(n8393) );
  XOR U8998 ( .A(n8392), .B(n8393), .Z(n8399) );
  XOR U8999 ( .A(n8398), .B(n8399), .Z(n8411) );
  XNOR U9000 ( .A(n8410), .B(n8411), .Z(n8342) );
  XNOR U9001 ( .A(n8343), .B(n8342), .Z(n8344) );
  XOR U9002 ( .A(n8345), .B(n8344), .Z(n8463) );
  XNOR U9003 ( .A(n8462), .B(n8463), .Z(n8464) );
  XNOR U9004 ( .A(n8465), .B(n8464), .Z(n8338) );
  XOR U9005 ( .A(n8339), .B(n8338), .Z(n8331) );
  NANDN U9006 ( .A(n8314), .B(n8313), .Z(n8318) );
  OR U9007 ( .A(n8316), .B(n8315), .Z(n8317) );
  AND U9008 ( .A(n8318), .B(n8317), .Z(n8330) );
  XNOR U9009 ( .A(n8331), .B(n8330), .Z(n8332) );
  XNOR U9010 ( .A(n8333), .B(n8332), .Z(n8324) );
  XNOR U9011 ( .A(n8325), .B(n8324), .Z(n8326) );
  XNOR U9012 ( .A(n8327), .B(n8326), .Z(n8468) );
  XNOR U9013 ( .A(sreg[294]), .B(n8468), .Z(n8470) );
  NANDN U9014 ( .A(sreg[293]), .B(n8319), .Z(n8323) );
  NAND U9015 ( .A(n8321), .B(n8320), .Z(n8322) );
  NAND U9016 ( .A(n8323), .B(n8322), .Z(n8469) );
  XNOR U9017 ( .A(n8470), .B(n8469), .Z(c[294]) );
  NANDN U9018 ( .A(n8325), .B(n8324), .Z(n8329) );
  NANDN U9019 ( .A(n8327), .B(n8326), .Z(n8328) );
  AND U9020 ( .A(n8329), .B(n8328), .Z(n8476) );
  NANDN U9021 ( .A(n8331), .B(n8330), .Z(n8335) );
  NANDN U9022 ( .A(n8333), .B(n8332), .Z(n8334) );
  AND U9023 ( .A(n8335), .B(n8334), .Z(n8474) );
  NANDN U9024 ( .A(n8337), .B(n8336), .Z(n8341) );
  NAND U9025 ( .A(n8339), .B(n8338), .Z(n8340) );
  AND U9026 ( .A(n8341), .B(n8340), .Z(n8481) );
  NANDN U9027 ( .A(n8343), .B(n8342), .Z(n8347) );
  NANDN U9028 ( .A(n8345), .B(n8344), .Z(n8346) );
  AND U9029 ( .A(n8347), .B(n8346), .Z(n8486) );
  NANDN U9030 ( .A(n8349), .B(n8348), .Z(n8353) );
  NAND U9031 ( .A(n8351), .B(n8350), .Z(n8352) );
  AND U9032 ( .A(n8353), .B(n8352), .Z(n8485) );
  XNOR U9033 ( .A(n8486), .B(n8485), .Z(n8488) );
  NANDN U9034 ( .A(n8355), .B(n8354), .Z(n8359) );
  NANDN U9035 ( .A(n8357), .B(n8356), .Z(n8358) );
  AND U9036 ( .A(n8359), .B(n8358), .Z(n8565) );
  NAND U9037 ( .A(n38385), .B(n8360), .Z(n8362) );
  XOR U9038 ( .A(b[27]), .B(a[45]), .Z(n8509) );
  NAND U9039 ( .A(n38343), .B(n8509), .Z(n8361) );
  AND U9040 ( .A(n8362), .B(n8361), .Z(n8572) );
  NAND U9041 ( .A(n183), .B(n8363), .Z(n8365) );
  XOR U9042 ( .A(b[5]), .B(a[67]), .Z(n8512) );
  NAND U9043 ( .A(n36296), .B(n8512), .Z(n8364) );
  AND U9044 ( .A(n8365), .B(n8364), .Z(n8570) );
  NAND U9045 ( .A(n190), .B(n8366), .Z(n8368) );
  XOR U9046 ( .A(b[19]), .B(a[53]), .Z(n8515) );
  NAND U9047 ( .A(n37821), .B(n8515), .Z(n8367) );
  NAND U9048 ( .A(n8368), .B(n8367), .Z(n8569) );
  XNOR U9049 ( .A(n8570), .B(n8569), .Z(n8571) );
  XNOR U9050 ( .A(n8572), .B(n8571), .Z(n8563) );
  NAND U9051 ( .A(n38470), .B(n8369), .Z(n8371) );
  XOR U9052 ( .A(b[31]), .B(a[41]), .Z(n8518) );
  NAND U9053 ( .A(n38453), .B(n8518), .Z(n8370) );
  AND U9054 ( .A(n8371), .B(n8370), .Z(n8530) );
  NAND U9055 ( .A(n181), .B(n8372), .Z(n8374) );
  XOR U9056 ( .A(b[3]), .B(a[69]), .Z(n8521) );
  NAND U9057 ( .A(n182), .B(n8521), .Z(n8373) );
  AND U9058 ( .A(n8374), .B(n8373), .Z(n8528) );
  NAND U9059 ( .A(n189), .B(n8375), .Z(n8377) );
  XOR U9060 ( .A(b[17]), .B(a[55]), .Z(n8524) );
  NAND U9061 ( .A(n37652), .B(n8524), .Z(n8376) );
  NAND U9062 ( .A(n8377), .B(n8376), .Z(n8527) );
  XNOR U9063 ( .A(n8528), .B(n8527), .Z(n8529) );
  XOR U9064 ( .A(n8530), .B(n8529), .Z(n8564) );
  XOR U9065 ( .A(n8563), .B(n8564), .Z(n8566) );
  XOR U9066 ( .A(n8565), .B(n8566), .Z(n8498) );
  NANDN U9067 ( .A(n8379), .B(n8378), .Z(n8383) );
  NANDN U9068 ( .A(n8381), .B(n8380), .Z(n8382) );
  AND U9069 ( .A(n8383), .B(n8382), .Z(n8551) );
  NANDN U9070 ( .A(n8385), .B(n8384), .Z(n8389) );
  NANDN U9071 ( .A(n8387), .B(n8386), .Z(n8388) );
  NAND U9072 ( .A(n8389), .B(n8388), .Z(n8552) );
  XNOR U9073 ( .A(n8551), .B(n8552), .Z(n8553) );
  NANDN U9074 ( .A(n8391), .B(n8390), .Z(n8395) );
  NANDN U9075 ( .A(n8393), .B(n8392), .Z(n8394) );
  NAND U9076 ( .A(n8395), .B(n8394), .Z(n8554) );
  XNOR U9077 ( .A(n8553), .B(n8554), .Z(n8497) );
  XNOR U9078 ( .A(n8498), .B(n8497), .Z(n8500) );
  NANDN U9079 ( .A(n8397), .B(n8396), .Z(n8401) );
  NANDN U9080 ( .A(n8399), .B(n8398), .Z(n8400) );
  AND U9081 ( .A(n8401), .B(n8400), .Z(n8499) );
  XOR U9082 ( .A(n8500), .B(n8499), .Z(n8614) );
  NANDN U9083 ( .A(n8403), .B(n8402), .Z(n8407) );
  NANDN U9084 ( .A(n8405), .B(n8404), .Z(n8406) );
  AND U9085 ( .A(n8407), .B(n8406), .Z(n8611) );
  NANDN U9086 ( .A(n8409), .B(n8408), .Z(n8413) );
  NANDN U9087 ( .A(n8411), .B(n8410), .Z(n8412) );
  AND U9088 ( .A(n8413), .B(n8412), .Z(n8494) );
  NANDN U9089 ( .A(n8415), .B(n8414), .Z(n8419) );
  OR U9090 ( .A(n8417), .B(n8416), .Z(n8418) );
  AND U9091 ( .A(n8419), .B(n8418), .Z(n8492) );
  NANDN U9092 ( .A(n8421), .B(n8420), .Z(n8425) );
  NANDN U9093 ( .A(n8423), .B(n8422), .Z(n8424) );
  AND U9094 ( .A(n8425), .B(n8424), .Z(n8558) );
  NANDN U9095 ( .A(n8427), .B(n8426), .Z(n8431) );
  NANDN U9096 ( .A(n8429), .B(n8428), .Z(n8430) );
  NAND U9097 ( .A(n8431), .B(n8430), .Z(n8557) );
  XNOR U9098 ( .A(n8558), .B(n8557), .Z(n8559) );
  NAND U9099 ( .A(b[0]), .B(a[71]), .Z(n8432) );
  XNOR U9100 ( .A(b[1]), .B(n8432), .Z(n8434) );
  NANDN U9101 ( .A(b[0]), .B(a[70]), .Z(n8433) );
  NAND U9102 ( .A(n8434), .B(n8433), .Z(n8506) );
  NAND U9103 ( .A(n194), .B(n8435), .Z(n8437) );
  XOR U9104 ( .A(b[29]), .B(a[43]), .Z(n8584) );
  NAND U9105 ( .A(n38456), .B(n8584), .Z(n8436) );
  AND U9106 ( .A(n8437), .B(n8436), .Z(n8504) );
  AND U9107 ( .A(b[31]), .B(a[39]), .Z(n8503) );
  XNOR U9108 ( .A(n8504), .B(n8503), .Z(n8505) );
  XNOR U9109 ( .A(n8506), .B(n8505), .Z(n8545) );
  NAND U9110 ( .A(n38185), .B(n8438), .Z(n8440) );
  XOR U9111 ( .A(b[23]), .B(a[49]), .Z(n8587) );
  NAND U9112 ( .A(n38132), .B(n8587), .Z(n8439) );
  AND U9113 ( .A(n8440), .B(n8439), .Z(n8578) );
  NAND U9114 ( .A(n184), .B(n8441), .Z(n8443) );
  XOR U9115 ( .A(b[7]), .B(a[65]), .Z(n8590) );
  NAND U9116 ( .A(n36592), .B(n8590), .Z(n8442) );
  AND U9117 ( .A(n8443), .B(n8442), .Z(n8576) );
  NAND U9118 ( .A(n38289), .B(n8444), .Z(n8446) );
  XOR U9119 ( .A(b[25]), .B(a[47]), .Z(n8593) );
  NAND U9120 ( .A(n38247), .B(n8593), .Z(n8445) );
  NAND U9121 ( .A(n8446), .B(n8445), .Z(n8575) );
  XNOR U9122 ( .A(n8576), .B(n8575), .Z(n8577) );
  XOR U9123 ( .A(n8578), .B(n8577), .Z(n8546) );
  XNOR U9124 ( .A(n8545), .B(n8546), .Z(n8547) );
  NAND U9125 ( .A(n187), .B(n8447), .Z(n8449) );
  XOR U9126 ( .A(b[13]), .B(a[59]), .Z(n8596) );
  NAND U9127 ( .A(n37295), .B(n8596), .Z(n8448) );
  AND U9128 ( .A(n8449), .B(n8448), .Z(n8540) );
  NAND U9129 ( .A(n186), .B(n8450), .Z(n8452) );
  XOR U9130 ( .A(b[11]), .B(a[61]), .Z(n8599) );
  NAND U9131 ( .A(n37097), .B(n8599), .Z(n8451) );
  NAND U9132 ( .A(n8452), .B(n8451), .Z(n8539) );
  XNOR U9133 ( .A(n8540), .B(n8539), .Z(n8541) );
  NAND U9134 ( .A(n188), .B(n8453), .Z(n8455) );
  XOR U9135 ( .A(b[15]), .B(a[57]), .Z(n8602) );
  NAND U9136 ( .A(n37382), .B(n8602), .Z(n8454) );
  AND U9137 ( .A(n8455), .B(n8454), .Z(n8536) );
  NAND U9138 ( .A(n38064), .B(n8456), .Z(n8458) );
  XOR U9139 ( .A(b[21]), .B(a[51]), .Z(n8605) );
  NAND U9140 ( .A(n37993), .B(n8605), .Z(n8457) );
  AND U9141 ( .A(n8458), .B(n8457), .Z(n8534) );
  NAND U9142 ( .A(n185), .B(n8459), .Z(n8461) );
  XOR U9143 ( .A(b[9]), .B(a[63]), .Z(n8608) );
  NAND U9144 ( .A(n36805), .B(n8608), .Z(n8460) );
  NAND U9145 ( .A(n8461), .B(n8460), .Z(n8533) );
  XNOR U9146 ( .A(n8534), .B(n8533), .Z(n8535) );
  XOR U9147 ( .A(n8536), .B(n8535), .Z(n8542) );
  XOR U9148 ( .A(n8541), .B(n8542), .Z(n8548) );
  XOR U9149 ( .A(n8547), .B(n8548), .Z(n8560) );
  XNOR U9150 ( .A(n8559), .B(n8560), .Z(n8491) );
  XNOR U9151 ( .A(n8492), .B(n8491), .Z(n8493) );
  XOR U9152 ( .A(n8494), .B(n8493), .Z(n8612) );
  XNOR U9153 ( .A(n8611), .B(n8612), .Z(n8613) );
  XNOR U9154 ( .A(n8614), .B(n8613), .Z(n8487) );
  XOR U9155 ( .A(n8488), .B(n8487), .Z(n8480) );
  NANDN U9156 ( .A(n8463), .B(n8462), .Z(n8467) );
  NANDN U9157 ( .A(n8465), .B(n8464), .Z(n8466) );
  AND U9158 ( .A(n8467), .B(n8466), .Z(n8479) );
  XOR U9159 ( .A(n8480), .B(n8479), .Z(n8482) );
  XNOR U9160 ( .A(n8481), .B(n8482), .Z(n8473) );
  XNOR U9161 ( .A(n8474), .B(n8473), .Z(n8475) );
  XNOR U9162 ( .A(n8476), .B(n8475), .Z(n8617) );
  XNOR U9163 ( .A(sreg[295]), .B(n8617), .Z(n8619) );
  NANDN U9164 ( .A(sreg[294]), .B(n8468), .Z(n8472) );
  NAND U9165 ( .A(n8470), .B(n8469), .Z(n8471) );
  NAND U9166 ( .A(n8472), .B(n8471), .Z(n8618) );
  XNOR U9167 ( .A(n8619), .B(n8618), .Z(c[295]) );
  NANDN U9168 ( .A(n8474), .B(n8473), .Z(n8478) );
  NANDN U9169 ( .A(n8476), .B(n8475), .Z(n8477) );
  AND U9170 ( .A(n8478), .B(n8477), .Z(n8625) );
  NANDN U9171 ( .A(n8480), .B(n8479), .Z(n8484) );
  NANDN U9172 ( .A(n8482), .B(n8481), .Z(n8483) );
  AND U9173 ( .A(n8484), .B(n8483), .Z(n8623) );
  NANDN U9174 ( .A(n8486), .B(n8485), .Z(n8490) );
  NAND U9175 ( .A(n8488), .B(n8487), .Z(n8489) );
  AND U9176 ( .A(n8490), .B(n8489), .Z(n8630) );
  NANDN U9177 ( .A(n8492), .B(n8491), .Z(n8496) );
  NANDN U9178 ( .A(n8494), .B(n8493), .Z(n8495) );
  AND U9179 ( .A(n8496), .B(n8495), .Z(n8635) );
  NANDN U9180 ( .A(n8498), .B(n8497), .Z(n8502) );
  NAND U9181 ( .A(n8500), .B(n8499), .Z(n8501) );
  AND U9182 ( .A(n8502), .B(n8501), .Z(n8634) );
  XNOR U9183 ( .A(n8635), .B(n8634), .Z(n8637) );
  NANDN U9184 ( .A(n8504), .B(n8503), .Z(n8508) );
  NANDN U9185 ( .A(n8506), .B(n8505), .Z(n8507) );
  AND U9186 ( .A(n8508), .B(n8507), .Z(n8714) );
  NAND U9187 ( .A(n38385), .B(n8509), .Z(n8511) );
  XOR U9188 ( .A(b[27]), .B(a[46]), .Z(n8658) );
  NAND U9189 ( .A(n38343), .B(n8658), .Z(n8510) );
  AND U9190 ( .A(n8511), .B(n8510), .Z(n8721) );
  NAND U9191 ( .A(n183), .B(n8512), .Z(n8514) );
  XOR U9192 ( .A(b[5]), .B(a[68]), .Z(n8661) );
  NAND U9193 ( .A(n36296), .B(n8661), .Z(n8513) );
  AND U9194 ( .A(n8514), .B(n8513), .Z(n8719) );
  NAND U9195 ( .A(n190), .B(n8515), .Z(n8517) );
  XOR U9196 ( .A(b[19]), .B(a[54]), .Z(n8664) );
  NAND U9197 ( .A(n37821), .B(n8664), .Z(n8516) );
  NAND U9198 ( .A(n8517), .B(n8516), .Z(n8718) );
  XNOR U9199 ( .A(n8719), .B(n8718), .Z(n8720) );
  XNOR U9200 ( .A(n8721), .B(n8720), .Z(n8712) );
  NAND U9201 ( .A(n38470), .B(n8518), .Z(n8520) );
  XOR U9202 ( .A(b[31]), .B(a[42]), .Z(n8667) );
  NAND U9203 ( .A(n38453), .B(n8667), .Z(n8519) );
  AND U9204 ( .A(n8520), .B(n8519), .Z(n8679) );
  NAND U9205 ( .A(n181), .B(n8521), .Z(n8523) );
  XOR U9206 ( .A(b[3]), .B(a[70]), .Z(n8670) );
  NAND U9207 ( .A(n182), .B(n8670), .Z(n8522) );
  AND U9208 ( .A(n8523), .B(n8522), .Z(n8677) );
  NAND U9209 ( .A(n189), .B(n8524), .Z(n8526) );
  XOR U9210 ( .A(b[17]), .B(a[56]), .Z(n8673) );
  NAND U9211 ( .A(n37652), .B(n8673), .Z(n8525) );
  NAND U9212 ( .A(n8526), .B(n8525), .Z(n8676) );
  XNOR U9213 ( .A(n8677), .B(n8676), .Z(n8678) );
  XOR U9214 ( .A(n8679), .B(n8678), .Z(n8713) );
  XOR U9215 ( .A(n8712), .B(n8713), .Z(n8715) );
  XOR U9216 ( .A(n8714), .B(n8715), .Z(n8647) );
  NANDN U9217 ( .A(n8528), .B(n8527), .Z(n8532) );
  NANDN U9218 ( .A(n8530), .B(n8529), .Z(n8531) );
  AND U9219 ( .A(n8532), .B(n8531), .Z(n8700) );
  NANDN U9220 ( .A(n8534), .B(n8533), .Z(n8538) );
  NANDN U9221 ( .A(n8536), .B(n8535), .Z(n8537) );
  NAND U9222 ( .A(n8538), .B(n8537), .Z(n8701) );
  XNOR U9223 ( .A(n8700), .B(n8701), .Z(n8702) );
  NANDN U9224 ( .A(n8540), .B(n8539), .Z(n8544) );
  NANDN U9225 ( .A(n8542), .B(n8541), .Z(n8543) );
  NAND U9226 ( .A(n8544), .B(n8543), .Z(n8703) );
  XNOR U9227 ( .A(n8702), .B(n8703), .Z(n8646) );
  XNOR U9228 ( .A(n8647), .B(n8646), .Z(n8649) );
  NANDN U9229 ( .A(n8546), .B(n8545), .Z(n8550) );
  NANDN U9230 ( .A(n8548), .B(n8547), .Z(n8549) );
  AND U9231 ( .A(n8550), .B(n8549), .Z(n8648) );
  XOR U9232 ( .A(n8649), .B(n8648), .Z(n8763) );
  NANDN U9233 ( .A(n8552), .B(n8551), .Z(n8556) );
  NANDN U9234 ( .A(n8554), .B(n8553), .Z(n8555) );
  AND U9235 ( .A(n8556), .B(n8555), .Z(n8760) );
  NANDN U9236 ( .A(n8558), .B(n8557), .Z(n8562) );
  NANDN U9237 ( .A(n8560), .B(n8559), .Z(n8561) );
  AND U9238 ( .A(n8562), .B(n8561), .Z(n8643) );
  NANDN U9239 ( .A(n8564), .B(n8563), .Z(n8568) );
  OR U9240 ( .A(n8566), .B(n8565), .Z(n8567) );
  AND U9241 ( .A(n8568), .B(n8567), .Z(n8641) );
  NANDN U9242 ( .A(n8570), .B(n8569), .Z(n8574) );
  NANDN U9243 ( .A(n8572), .B(n8571), .Z(n8573) );
  AND U9244 ( .A(n8574), .B(n8573), .Z(n8707) );
  NANDN U9245 ( .A(n8576), .B(n8575), .Z(n8580) );
  NANDN U9246 ( .A(n8578), .B(n8577), .Z(n8579) );
  NAND U9247 ( .A(n8580), .B(n8579), .Z(n8706) );
  XNOR U9248 ( .A(n8707), .B(n8706), .Z(n8708) );
  NAND U9249 ( .A(b[0]), .B(a[72]), .Z(n8581) );
  XNOR U9250 ( .A(b[1]), .B(n8581), .Z(n8583) );
  NANDN U9251 ( .A(b[0]), .B(a[71]), .Z(n8582) );
  NAND U9252 ( .A(n8583), .B(n8582), .Z(n8655) );
  NAND U9253 ( .A(n194), .B(n8584), .Z(n8586) );
  XOR U9254 ( .A(b[29]), .B(a[44]), .Z(n8733) );
  NAND U9255 ( .A(n38456), .B(n8733), .Z(n8585) );
  AND U9256 ( .A(n8586), .B(n8585), .Z(n8653) );
  AND U9257 ( .A(b[31]), .B(a[40]), .Z(n8652) );
  XNOR U9258 ( .A(n8653), .B(n8652), .Z(n8654) );
  XNOR U9259 ( .A(n8655), .B(n8654), .Z(n8694) );
  NAND U9260 ( .A(n38185), .B(n8587), .Z(n8589) );
  XOR U9261 ( .A(b[23]), .B(a[50]), .Z(n8736) );
  NAND U9262 ( .A(n38132), .B(n8736), .Z(n8588) );
  AND U9263 ( .A(n8589), .B(n8588), .Z(n8727) );
  NAND U9264 ( .A(n184), .B(n8590), .Z(n8592) );
  XOR U9265 ( .A(b[7]), .B(a[66]), .Z(n8739) );
  NAND U9266 ( .A(n36592), .B(n8739), .Z(n8591) );
  AND U9267 ( .A(n8592), .B(n8591), .Z(n8725) );
  NAND U9268 ( .A(n38289), .B(n8593), .Z(n8595) );
  XOR U9269 ( .A(b[25]), .B(a[48]), .Z(n8742) );
  NAND U9270 ( .A(n38247), .B(n8742), .Z(n8594) );
  NAND U9271 ( .A(n8595), .B(n8594), .Z(n8724) );
  XNOR U9272 ( .A(n8725), .B(n8724), .Z(n8726) );
  XOR U9273 ( .A(n8727), .B(n8726), .Z(n8695) );
  XNOR U9274 ( .A(n8694), .B(n8695), .Z(n8696) );
  NAND U9275 ( .A(n187), .B(n8596), .Z(n8598) );
  XOR U9276 ( .A(b[13]), .B(a[60]), .Z(n8745) );
  NAND U9277 ( .A(n37295), .B(n8745), .Z(n8597) );
  AND U9278 ( .A(n8598), .B(n8597), .Z(n8689) );
  NAND U9279 ( .A(n186), .B(n8599), .Z(n8601) );
  XOR U9280 ( .A(b[11]), .B(a[62]), .Z(n8748) );
  NAND U9281 ( .A(n37097), .B(n8748), .Z(n8600) );
  NAND U9282 ( .A(n8601), .B(n8600), .Z(n8688) );
  XNOR U9283 ( .A(n8689), .B(n8688), .Z(n8690) );
  NAND U9284 ( .A(n188), .B(n8602), .Z(n8604) );
  XOR U9285 ( .A(b[15]), .B(a[58]), .Z(n8751) );
  NAND U9286 ( .A(n37382), .B(n8751), .Z(n8603) );
  AND U9287 ( .A(n8604), .B(n8603), .Z(n8685) );
  NAND U9288 ( .A(n38064), .B(n8605), .Z(n8607) );
  XOR U9289 ( .A(b[21]), .B(a[52]), .Z(n8754) );
  NAND U9290 ( .A(n37993), .B(n8754), .Z(n8606) );
  AND U9291 ( .A(n8607), .B(n8606), .Z(n8683) );
  NAND U9292 ( .A(n185), .B(n8608), .Z(n8610) );
  XOR U9293 ( .A(b[9]), .B(a[64]), .Z(n8757) );
  NAND U9294 ( .A(n36805), .B(n8757), .Z(n8609) );
  NAND U9295 ( .A(n8610), .B(n8609), .Z(n8682) );
  XNOR U9296 ( .A(n8683), .B(n8682), .Z(n8684) );
  XOR U9297 ( .A(n8685), .B(n8684), .Z(n8691) );
  XOR U9298 ( .A(n8690), .B(n8691), .Z(n8697) );
  XOR U9299 ( .A(n8696), .B(n8697), .Z(n8709) );
  XNOR U9300 ( .A(n8708), .B(n8709), .Z(n8640) );
  XNOR U9301 ( .A(n8641), .B(n8640), .Z(n8642) );
  XOR U9302 ( .A(n8643), .B(n8642), .Z(n8761) );
  XNOR U9303 ( .A(n8760), .B(n8761), .Z(n8762) );
  XNOR U9304 ( .A(n8763), .B(n8762), .Z(n8636) );
  XOR U9305 ( .A(n8637), .B(n8636), .Z(n8629) );
  NANDN U9306 ( .A(n8612), .B(n8611), .Z(n8616) );
  NANDN U9307 ( .A(n8614), .B(n8613), .Z(n8615) );
  AND U9308 ( .A(n8616), .B(n8615), .Z(n8628) );
  XOR U9309 ( .A(n8629), .B(n8628), .Z(n8631) );
  XNOR U9310 ( .A(n8630), .B(n8631), .Z(n8622) );
  XNOR U9311 ( .A(n8623), .B(n8622), .Z(n8624) );
  XNOR U9312 ( .A(n8625), .B(n8624), .Z(n8766) );
  XNOR U9313 ( .A(sreg[296]), .B(n8766), .Z(n8768) );
  NANDN U9314 ( .A(sreg[295]), .B(n8617), .Z(n8621) );
  NAND U9315 ( .A(n8619), .B(n8618), .Z(n8620) );
  NAND U9316 ( .A(n8621), .B(n8620), .Z(n8767) );
  XNOR U9317 ( .A(n8768), .B(n8767), .Z(c[296]) );
  NANDN U9318 ( .A(n8623), .B(n8622), .Z(n8627) );
  NANDN U9319 ( .A(n8625), .B(n8624), .Z(n8626) );
  AND U9320 ( .A(n8627), .B(n8626), .Z(n8774) );
  NANDN U9321 ( .A(n8629), .B(n8628), .Z(n8633) );
  NANDN U9322 ( .A(n8631), .B(n8630), .Z(n8632) );
  AND U9323 ( .A(n8633), .B(n8632), .Z(n8772) );
  NANDN U9324 ( .A(n8635), .B(n8634), .Z(n8639) );
  NAND U9325 ( .A(n8637), .B(n8636), .Z(n8638) );
  AND U9326 ( .A(n8639), .B(n8638), .Z(n8779) );
  NANDN U9327 ( .A(n8641), .B(n8640), .Z(n8645) );
  NANDN U9328 ( .A(n8643), .B(n8642), .Z(n8644) );
  AND U9329 ( .A(n8645), .B(n8644), .Z(n8910) );
  NANDN U9330 ( .A(n8647), .B(n8646), .Z(n8651) );
  NAND U9331 ( .A(n8649), .B(n8648), .Z(n8650) );
  AND U9332 ( .A(n8651), .B(n8650), .Z(n8909) );
  XNOR U9333 ( .A(n8910), .B(n8909), .Z(n8912) );
  NANDN U9334 ( .A(n8653), .B(n8652), .Z(n8657) );
  NANDN U9335 ( .A(n8655), .B(n8654), .Z(n8656) );
  AND U9336 ( .A(n8657), .B(n8656), .Z(n8857) );
  NAND U9337 ( .A(n38385), .B(n8658), .Z(n8660) );
  XOR U9338 ( .A(b[27]), .B(a[47]), .Z(n8801) );
  NAND U9339 ( .A(n38343), .B(n8801), .Z(n8659) );
  AND U9340 ( .A(n8660), .B(n8659), .Z(n8864) );
  NAND U9341 ( .A(n183), .B(n8661), .Z(n8663) );
  XOR U9342 ( .A(b[5]), .B(a[69]), .Z(n8804) );
  NAND U9343 ( .A(n36296), .B(n8804), .Z(n8662) );
  AND U9344 ( .A(n8663), .B(n8662), .Z(n8862) );
  NAND U9345 ( .A(n190), .B(n8664), .Z(n8666) );
  XOR U9346 ( .A(b[19]), .B(a[55]), .Z(n8807) );
  NAND U9347 ( .A(n37821), .B(n8807), .Z(n8665) );
  NAND U9348 ( .A(n8666), .B(n8665), .Z(n8861) );
  XNOR U9349 ( .A(n8862), .B(n8861), .Z(n8863) );
  XNOR U9350 ( .A(n8864), .B(n8863), .Z(n8855) );
  NAND U9351 ( .A(n38470), .B(n8667), .Z(n8669) );
  XOR U9352 ( .A(b[31]), .B(a[43]), .Z(n8810) );
  NAND U9353 ( .A(n38453), .B(n8810), .Z(n8668) );
  AND U9354 ( .A(n8669), .B(n8668), .Z(n8822) );
  NAND U9355 ( .A(n181), .B(n8670), .Z(n8672) );
  XOR U9356 ( .A(b[3]), .B(a[71]), .Z(n8813) );
  NAND U9357 ( .A(n182), .B(n8813), .Z(n8671) );
  AND U9358 ( .A(n8672), .B(n8671), .Z(n8820) );
  NAND U9359 ( .A(n189), .B(n8673), .Z(n8675) );
  XOR U9360 ( .A(b[17]), .B(a[57]), .Z(n8816) );
  NAND U9361 ( .A(n37652), .B(n8816), .Z(n8674) );
  NAND U9362 ( .A(n8675), .B(n8674), .Z(n8819) );
  XNOR U9363 ( .A(n8820), .B(n8819), .Z(n8821) );
  XOR U9364 ( .A(n8822), .B(n8821), .Z(n8856) );
  XOR U9365 ( .A(n8855), .B(n8856), .Z(n8858) );
  XOR U9366 ( .A(n8857), .B(n8858), .Z(n8790) );
  NANDN U9367 ( .A(n8677), .B(n8676), .Z(n8681) );
  NANDN U9368 ( .A(n8679), .B(n8678), .Z(n8680) );
  AND U9369 ( .A(n8681), .B(n8680), .Z(n8843) );
  NANDN U9370 ( .A(n8683), .B(n8682), .Z(n8687) );
  NANDN U9371 ( .A(n8685), .B(n8684), .Z(n8686) );
  NAND U9372 ( .A(n8687), .B(n8686), .Z(n8844) );
  XNOR U9373 ( .A(n8843), .B(n8844), .Z(n8845) );
  NANDN U9374 ( .A(n8689), .B(n8688), .Z(n8693) );
  NANDN U9375 ( .A(n8691), .B(n8690), .Z(n8692) );
  NAND U9376 ( .A(n8693), .B(n8692), .Z(n8846) );
  XNOR U9377 ( .A(n8845), .B(n8846), .Z(n8789) );
  XNOR U9378 ( .A(n8790), .B(n8789), .Z(n8792) );
  NANDN U9379 ( .A(n8695), .B(n8694), .Z(n8699) );
  NANDN U9380 ( .A(n8697), .B(n8696), .Z(n8698) );
  AND U9381 ( .A(n8699), .B(n8698), .Z(n8791) );
  XOR U9382 ( .A(n8792), .B(n8791), .Z(n8906) );
  NANDN U9383 ( .A(n8701), .B(n8700), .Z(n8705) );
  NANDN U9384 ( .A(n8703), .B(n8702), .Z(n8704) );
  AND U9385 ( .A(n8705), .B(n8704), .Z(n8903) );
  NANDN U9386 ( .A(n8707), .B(n8706), .Z(n8711) );
  NANDN U9387 ( .A(n8709), .B(n8708), .Z(n8710) );
  AND U9388 ( .A(n8711), .B(n8710), .Z(n8786) );
  NANDN U9389 ( .A(n8713), .B(n8712), .Z(n8717) );
  OR U9390 ( .A(n8715), .B(n8714), .Z(n8716) );
  AND U9391 ( .A(n8717), .B(n8716), .Z(n8784) );
  NANDN U9392 ( .A(n8719), .B(n8718), .Z(n8723) );
  NANDN U9393 ( .A(n8721), .B(n8720), .Z(n8722) );
  AND U9394 ( .A(n8723), .B(n8722), .Z(n8850) );
  NANDN U9395 ( .A(n8725), .B(n8724), .Z(n8729) );
  NANDN U9396 ( .A(n8727), .B(n8726), .Z(n8728) );
  NAND U9397 ( .A(n8729), .B(n8728), .Z(n8849) );
  XNOR U9398 ( .A(n8850), .B(n8849), .Z(n8851) );
  NAND U9399 ( .A(b[0]), .B(a[73]), .Z(n8730) );
  XNOR U9400 ( .A(b[1]), .B(n8730), .Z(n8732) );
  NANDN U9401 ( .A(b[0]), .B(a[72]), .Z(n8731) );
  NAND U9402 ( .A(n8732), .B(n8731), .Z(n8798) );
  NAND U9403 ( .A(n194), .B(n8733), .Z(n8735) );
  XOR U9404 ( .A(b[29]), .B(a[45]), .Z(n8873) );
  NAND U9405 ( .A(n38456), .B(n8873), .Z(n8734) );
  AND U9406 ( .A(n8735), .B(n8734), .Z(n8796) );
  AND U9407 ( .A(b[31]), .B(a[41]), .Z(n8795) );
  XNOR U9408 ( .A(n8796), .B(n8795), .Z(n8797) );
  XNOR U9409 ( .A(n8798), .B(n8797), .Z(n8837) );
  NAND U9410 ( .A(n38185), .B(n8736), .Z(n8738) );
  XOR U9411 ( .A(b[23]), .B(a[51]), .Z(n8879) );
  NAND U9412 ( .A(n38132), .B(n8879), .Z(n8737) );
  AND U9413 ( .A(n8738), .B(n8737), .Z(n8870) );
  NAND U9414 ( .A(n184), .B(n8739), .Z(n8741) );
  XOR U9415 ( .A(b[7]), .B(a[67]), .Z(n8882) );
  NAND U9416 ( .A(n36592), .B(n8882), .Z(n8740) );
  AND U9417 ( .A(n8741), .B(n8740), .Z(n8868) );
  NAND U9418 ( .A(n38289), .B(n8742), .Z(n8744) );
  XOR U9419 ( .A(b[25]), .B(a[49]), .Z(n8885) );
  NAND U9420 ( .A(n38247), .B(n8885), .Z(n8743) );
  NAND U9421 ( .A(n8744), .B(n8743), .Z(n8867) );
  XNOR U9422 ( .A(n8868), .B(n8867), .Z(n8869) );
  XOR U9423 ( .A(n8870), .B(n8869), .Z(n8838) );
  XNOR U9424 ( .A(n8837), .B(n8838), .Z(n8839) );
  NAND U9425 ( .A(n187), .B(n8745), .Z(n8747) );
  XOR U9426 ( .A(b[13]), .B(a[61]), .Z(n8888) );
  NAND U9427 ( .A(n37295), .B(n8888), .Z(n8746) );
  AND U9428 ( .A(n8747), .B(n8746), .Z(n8832) );
  NAND U9429 ( .A(n186), .B(n8748), .Z(n8750) );
  XOR U9430 ( .A(b[11]), .B(a[63]), .Z(n8891) );
  NAND U9431 ( .A(n37097), .B(n8891), .Z(n8749) );
  NAND U9432 ( .A(n8750), .B(n8749), .Z(n8831) );
  XNOR U9433 ( .A(n8832), .B(n8831), .Z(n8833) );
  NAND U9434 ( .A(n188), .B(n8751), .Z(n8753) );
  XOR U9435 ( .A(b[15]), .B(a[59]), .Z(n8894) );
  NAND U9436 ( .A(n37382), .B(n8894), .Z(n8752) );
  AND U9437 ( .A(n8753), .B(n8752), .Z(n8828) );
  NAND U9438 ( .A(n38064), .B(n8754), .Z(n8756) );
  XOR U9439 ( .A(b[21]), .B(a[53]), .Z(n8897) );
  NAND U9440 ( .A(n37993), .B(n8897), .Z(n8755) );
  AND U9441 ( .A(n8756), .B(n8755), .Z(n8826) );
  NAND U9442 ( .A(n185), .B(n8757), .Z(n8759) );
  XOR U9443 ( .A(b[9]), .B(a[65]), .Z(n8900) );
  NAND U9444 ( .A(n36805), .B(n8900), .Z(n8758) );
  NAND U9445 ( .A(n8759), .B(n8758), .Z(n8825) );
  XNOR U9446 ( .A(n8826), .B(n8825), .Z(n8827) );
  XOR U9447 ( .A(n8828), .B(n8827), .Z(n8834) );
  XOR U9448 ( .A(n8833), .B(n8834), .Z(n8840) );
  XOR U9449 ( .A(n8839), .B(n8840), .Z(n8852) );
  XNOR U9450 ( .A(n8851), .B(n8852), .Z(n8783) );
  XNOR U9451 ( .A(n8784), .B(n8783), .Z(n8785) );
  XOR U9452 ( .A(n8786), .B(n8785), .Z(n8904) );
  XNOR U9453 ( .A(n8903), .B(n8904), .Z(n8905) );
  XNOR U9454 ( .A(n8906), .B(n8905), .Z(n8911) );
  XOR U9455 ( .A(n8912), .B(n8911), .Z(n8778) );
  NANDN U9456 ( .A(n8761), .B(n8760), .Z(n8765) );
  NANDN U9457 ( .A(n8763), .B(n8762), .Z(n8764) );
  AND U9458 ( .A(n8765), .B(n8764), .Z(n8777) );
  XOR U9459 ( .A(n8778), .B(n8777), .Z(n8780) );
  XNOR U9460 ( .A(n8779), .B(n8780), .Z(n8771) );
  XNOR U9461 ( .A(n8772), .B(n8771), .Z(n8773) );
  XNOR U9462 ( .A(n8774), .B(n8773), .Z(n8915) );
  XNOR U9463 ( .A(sreg[297]), .B(n8915), .Z(n8917) );
  NANDN U9464 ( .A(sreg[296]), .B(n8766), .Z(n8770) );
  NAND U9465 ( .A(n8768), .B(n8767), .Z(n8769) );
  NAND U9466 ( .A(n8770), .B(n8769), .Z(n8916) );
  XNOR U9467 ( .A(n8917), .B(n8916), .Z(c[297]) );
  NANDN U9468 ( .A(n8772), .B(n8771), .Z(n8776) );
  NANDN U9469 ( .A(n8774), .B(n8773), .Z(n8775) );
  AND U9470 ( .A(n8776), .B(n8775), .Z(n8923) );
  NANDN U9471 ( .A(n8778), .B(n8777), .Z(n8782) );
  NANDN U9472 ( .A(n8780), .B(n8779), .Z(n8781) );
  AND U9473 ( .A(n8782), .B(n8781), .Z(n8921) );
  NANDN U9474 ( .A(n8784), .B(n8783), .Z(n8788) );
  NANDN U9475 ( .A(n8786), .B(n8785), .Z(n8787) );
  AND U9476 ( .A(n8788), .B(n8787), .Z(n9059) );
  NANDN U9477 ( .A(n8790), .B(n8789), .Z(n8794) );
  NAND U9478 ( .A(n8792), .B(n8791), .Z(n8793) );
  AND U9479 ( .A(n8794), .B(n8793), .Z(n9058) );
  XNOR U9480 ( .A(n9059), .B(n9058), .Z(n9061) );
  NANDN U9481 ( .A(n8796), .B(n8795), .Z(n8800) );
  NANDN U9482 ( .A(n8798), .B(n8797), .Z(n8799) );
  AND U9483 ( .A(n8800), .B(n8799), .Z(n9006) );
  NAND U9484 ( .A(n38385), .B(n8801), .Z(n8803) );
  XOR U9485 ( .A(b[27]), .B(a[48]), .Z(n8950) );
  NAND U9486 ( .A(n38343), .B(n8950), .Z(n8802) );
  AND U9487 ( .A(n8803), .B(n8802), .Z(n9013) );
  NAND U9488 ( .A(n183), .B(n8804), .Z(n8806) );
  XOR U9489 ( .A(b[5]), .B(a[70]), .Z(n8953) );
  NAND U9490 ( .A(n36296), .B(n8953), .Z(n8805) );
  AND U9491 ( .A(n8806), .B(n8805), .Z(n9011) );
  NAND U9492 ( .A(n190), .B(n8807), .Z(n8809) );
  XOR U9493 ( .A(b[19]), .B(a[56]), .Z(n8956) );
  NAND U9494 ( .A(n37821), .B(n8956), .Z(n8808) );
  NAND U9495 ( .A(n8809), .B(n8808), .Z(n9010) );
  XNOR U9496 ( .A(n9011), .B(n9010), .Z(n9012) );
  XNOR U9497 ( .A(n9013), .B(n9012), .Z(n9004) );
  NAND U9498 ( .A(n38470), .B(n8810), .Z(n8812) );
  XOR U9499 ( .A(b[31]), .B(a[44]), .Z(n8959) );
  NAND U9500 ( .A(n38453), .B(n8959), .Z(n8811) );
  AND U9501 ( .A(n8812), .B(n8811), .Z(n8971) );
  NAND U9502 ( .A(n181), .B(n8813), .Z(n8815) );
  XOR U9503 ( .A(b[3]), .B(a[72]), .Z(n8962) );
  NAND U9504 ( .A(n182), .B(n8962), .Z(n8814) );
  AND U9505 ( .A(n8815), .B(n8814), .Z(n8969) );
  NAND U9506 ( .A(n189), .B(n8816), .Z(n8818) );
  XOR U9507 ( .A(b[17]), .B(a[58]), .Z(n8965) );
  NAND U9508 ( .A(n37652), .B(n8965), .Z(n8817) );
  NAND U9509 ( .A(n8818), .B(n8817), .Z(n8968) );
  XNOR U9510 ( .A(n8969), .B(n8968), .Z(n8970) );
  XOR U9511 ( .A(n8971), .B(n8970), .Z(n9005) );
  XOR U9512 ( .A(n9004), .B(n9005), .Z(n9007) );
  XOR U9513 ( .A(n9006), .B(n9007), .Z(n8939) );
  NANDN U9514 ( .A(n8820), .B(n8819), .Z(n8824) );
  NANDN U9515 ( .A(n8822), .B(n8821), .Z(n8823) );
  AND U9516 ( .A(n8824), .B(n8823), .Z(n8992) );
  NANDN U9517 ( .A(n8826), .B(n8825), .Z(n8830) );
  NANDN U9518 ( .A(n8828), .B(n8827), .Z(n8829) );
  NAND U9519 ( .A(n8830), .B(n8829), .Z(n8993) );
  XNOR U9520 ( .A(n8992), .B(n8993), .Z(n8994) );
  NANDN U9521 ( .A(n8832), .B(n8831), .Z(n8836) );
  NANDN U9522 ( .A(n8834), .B(n8833), .Z(n8835) );
  NAND U9523 ( .A(n8836), .B(n8835), .Z(n8995) );
  XNOR U9524 ( .A(n8994), .B(n8995), .Z(n8938) );
  XNOR U9525 ( .A(n8939), .B(n8938), .Z(n8941) );
  NANDN U9526 ( .A(n8838), .B(n8837), .Z(n8842) );
  NANDN U9527 ( .A(n8840), .B(n8839), .Z(n8841) );
  AND U9528 ( .A(n8842), .B(n8841), .Z(n8940) );
  XOR U9529 ( .A(n8941), .B(n8940), .Z(n9055) );
  NANDN U9530 ( .A(n8844), .B(n8843), .Z(n8848) );
  NANDN U9531 ( .A(n8846), .B(n8845), .Z(n8847) );
  AND U9532 ( .A(n8848), .B(n8847), .Z(n9052) );
  NANDN U9533 ( .A(n8850), .B(n8849), .Z(n8854) );
  NANDN U9534 ( .A(n8852), .B(n8851), .Z(n8853) );
  AND U9535 ( .A(n8854), .B(n8853), .Z(n8935) );
  NANDN U9536 ( .A(n8856), .B(n8855), .Z(n8860) );
  OR U9537 ( .A(n8858), .B(n8857), .Z(n8859) );
  AND U9538 ( .A(n8860), .B(n8859), .Z(n8933) );
  NANDN U9539 ( .A(n8862), .B(n8861), .Z(n8866) );
  NANDN U9540 ( .A(n8864), .B(n8863), .Z(n8865) );
  AND U9541 ( .A(n8866), .B(n8865), .Z(n8999) );
  NANDN U9542 ( .A(n8868), .B(n8867), .Z(n8872) );
  NANDN U9543 ( .A(n8870), .B(n8869), .Z(n8871) );
  NAND U9544 ( .A(n8872), .B(n8871), .Z(n8998) );
  XNOR U9545 ( .A(n8999), .B(n8998), .Z(n9000) );
  NAND U9546 ( .A(n194), .B(n8873), .Z(n8875) );
  XOR U9547 ( .A(b[29]), .B(a[46]), .Z(n9025) );
  NAND U9548 ( .A(n38456), .B(n9025), .Z(n8874) );
  AND U9549 ( .A(n8875), .B(n8874), .Z(n8945) );
  AND U9550 ( .A(b[31]), .B(a[42]), .Z(n8944) );
  XNOR U9551 ( .A(n8945), .B(n8944), .Z(n8946) );
  NAND U9552 ( .A(b[0]), .B(a[74]), .Z(n8876) );
  XNOR U9553 ( .A(b[1]), .B(n8876), .Z(n8878) );
  NANDN U9554 ( .A(b[0]), .B(a[73]), .Z(n8877) );
  NAND U9555 ( .A(n8878), .B(n8877), .Z(n8947) );
  XNOR U9556 ( .A(n8946), .B(n8947), .Z(n8986) );
  NAND U9557 ( .A(n38185), .B(n8879), .Z(n8881) );
  XOR U9558 ( .A(b[23]), .B(a[52]), .Z(n9028) );
  NAND U9559 ( .A(n38132), .B(n9028), .Z(n8880) );
  AND U9560 ( .A(n8881), .B(n8880), .Z(n9019) );
  NAND U9561 ( .A(n184), .B(n8882), .Z(n8884) );
  XOR U9562 ( .A(b[7]), .B(a[68]), .Z(n9031) );
  NAND U9563 ( .A(n36592), .B(n9031), .Z(n8883) );
  AND U9564 ( .A(n8884), .B(n8883), .Z(n9017) );
  NAND U9565 ( .A(n38289), .B(n8885), .Z(n8887) );
  XOR U9566 ( .A(b[25]), .B(a[50]), .Z(n9034) );
  NAND U9567 ( .A(n38247), .B(n9034), .Z(n8886) );
  NAND U9568 ( .A(n8887), .B(n8886), .Z(n9016) );
  XNOR U9569 ( .A(n9017), .B(n9016), .Z(n9018) );
  XOR U9570 ( .A(n9019), .B(n9018), .Z(n8987) );
  XNOR U9571 ( .A(n8986), .B(n8987), .Z(n8988) );
  NAND U9572 ( .A(n187), .B(n8888), .Z(n8890) );
  XOR U9573 ( .A(b[13]), .B(a[62]), .Z(n9037) );
  NAND U9574 ( .A(n37295), .B(n9037), .Z(n8889) );
  AND U9575 ( .A(n8890), .B(n8889), .Z(n8981) );
  NAND U9576 ( .A(n186), .B(n8891), .Z(n8893) );
  XOR U9577 ( .A(b[11]), .B(a[64]), .Z(n9040) );
  NAND U9578 ( .A(n37097), .B(n9040), .Z(n8892) );
  NAND U9579 ( .A(n8893), .B(n8892), .Z(n8980) );
  XNOR U9580 ( .A(n8981), .B(n8980), .Z(n8982) );
  NAND U9581 ( .A(n188), .B(n8894), .Z(n8896) );
  XOR U9582 ( .A(b[15]), .B(a[60]), .Z(n9043) );
  NAND U9583 ( .A(n37382), .B(n9043), .Z(n8895) );
  AND U9584 ( .A(n8896), .B(n8895), .Z(n8977) );
  NAND U9585 ( .A(n38064), .B(n8897), .Z(n8899) );
  XOR U9586 ( .A(b[21]), .B(a[54]), .Z(n9046) );
  NAND U9587 ( .A(n37993), .B(n9046), .Z(n8898) );
  AND U9588 ( .A(n8899), .B(n8898), .Z(n8975) );
  NAND U9589 ( .A(n185), .B(n8900), .Z(n8902) );
  XOR U9590 ( .A(b[9]), .B(a[66]), .Z(n9049) );
  NAND U9591 ( .A(n36805), .B(n9049), .Z(n8901) );
  NAND U9592 ( .A(n8902), .B(n8901), .Z(n8974) );
  XNOR U9593 ( .A(n8975), .B(n8974), .Z(n8976) );
  XOR U9594 ( .A(n8977), .B(n8976), .Z(n8983) );
  XOR U9595 ( .A(n8982), .B(n8983), .Z(n8989) );
  XOR U9596 ( .A(n8988), .B(n8989), .Z(n9001) );
  XNOR U9597 ( .A(n9000), .B(n9001), .Z(n8932) );
  XNOR U9598 ( .A(n8933), .B(n8932), .Z(n8934) );
  XOR U9599 ( .A(n8935), .B(n8934), .Z(n9053) );
  XNOR U9600 ( .A(n9052), .B(n9053), .Z(n9054) );
  XNOR U9601 ( .A(n9055), .B(n9054), .Z(n9060) );
  XOR U9602 ( .A(n9061), .B(n9060), .Z(n8927) );
  NANDN U9603 ( .A(n8904), .B(n8903), .Z(n8908) );
  NANDN U9604 ( .A(n8906), .B(n8905), .Z(n8907) );
  AND U9605 ( .A(n8908), .B(n8907), .Z(n8926) );
  XNOR U9606 ( .A(n8927), .B(n8926), .Z(n8928) );
  NANDN U9607 ( .A(n8910), .B(n8909), .Z(n8914) );
  NAND U9608 ( .A(n8912), .B(n8911), .Z(n8913) );
  NAND U9609 ( .A(n8914), .B(n8913), .Z(n8929) );
  XNOR U9610 ( .A(n8928), .B(n8929), .Z(n8920) );
  XNOR U9611 ( .A(n8921), .B(n8920), .Z(n8922) );
  XNOR U9612 ( .A(n8923), .B(n8922), .Z(n9064) );
  XNOR U9613 ( .A(sreg[298]), .B(n9064), .Z(n9066) );
  NANDN U9614 ( .A(sreg[297]), .B(n8915), .Z(n8919) );
  NAND U9615 ( .A(n8917), .B(n8916), .Z(n8918) );
  NAND U9616 ( .A(n8919), .B(n8918), .Z(n9065) );
  XNOR U9617 ( .A(n9066), .B(n9065), .Z(c[298]) );
  NANDN U9618 ( .A(n8921), .B(n8920), .Z(n8925) );
  NANDN U9619 ( .A(n8923), .B(n8922), .Z(n8924) );
  AND U9620 ( .A(n8925), .B(n8924), .Z(n9072) );
  NANDN U9621 ( .A(n8927), .B(n8926), .Z(n8931) );
  NANDN U9622 ( .A(n8929), .B(n8928), .Z(n8930) );
  AND U9623 ( .A(n8931), .B(n8930), .Z(n9070) );
  NANDN U9624 ( .A(n8933), .B(n8932), .Z(n8937) );
  NANDN U9625 ( .A(n8935), .B(n8934), .Z(n8936) );
  AND U9626 ( .A(n8937), .B(n8936), .Z(n9208) );
  NANDN U9627 ( .A(n8939), .B(n8938), .Z(n8943) );
  NAND U9628 ( .A(n8941), .B(n8940), .Z(n8942) );
  AND U9629 ( .A(n8943), .B(n8942), .Z(n9207) );
  XNOR U9630 ( .A(n9208), .B(n9207), .Z(n9210) );
  NANDN U9631 ( .A(n8945), .B(n8944), .Z(n8949) );
  NANDN U9632 ( .A(n8947), .B(n8946), .Z(n8948) );
  AND U9633 ( .A(n8949), .B(n8948), .Z(n9155) );
  NAND U9634 ( .A(n38385), .B(n8950), .Z(n8952) );
  XOR U9635 ( .A(b[27]), .B(a[49]), .Z(n9099) );
  NAND U9636 ( .A(n38343), .B(n9099), .Z(n8951) );
  AND U9637 ( .A(n8952), .B(n8951), .Z(n9162) );
  NAND U9638 ( .A(n183), .B(n8953), .Z(n8955) );
  XOR U9639 ( .A(b[5]), .B(a[71]), .Z(n9102) );
  NAND U9640 ( .A(n36296), .B(n9102), .Z(n8954) );
  AND U9641 ( .A(n8955), .B(n8954), .Z(n9160) );
  NAND U9642 ( .A(n190), .B(n8956), .Z(n8958) );
  XOR U9643 ( .A(b[19]), .B(a[57]), .Z(n9105) );
  NAND U9644 ( .A(n37821), .B(n9105), .Z(n8957) );
  NAND U9645 ( .A(n8958), .B(n8957), .Z(n9159) );
  XNOR U9646 ( .A(n9160), .B(n9159), .Z(n9161) );
  XNOR U9647 ( .A(n9162), .B(n9161), .Z(n9153) );
  NAND U9648 ( .A(n38470), .B(n8959), .Z(n8961) );
  XOR U9649 ( .A(b[31]), .B(a[45]), .Z(n9108) );
  NAND U9650 ( .A(n38453), .B(n9108), .Z(n8960) );
  AND U9651 ( .A(n8961), .B(n8960), .Z(n9120) );
  NAND U9652 ( .A(n181), .B(n8962), .Z(n8964) );
  XOR U9653 ( .A(b[3]), .B(a[73]), .Z(n9111) );
  NAND U9654 ( .A(n182), .B(n9111), .Z(n8963) );
  AND U9655 ( .A(n8964), .B(n8963), .Z(n9118) );
  NAND U9656 ( .A(n189), .B(n8965), .Z(n8967) );
  XOR U9657 ( .A(b[17]), .B(a[59]), .Z(n9114) );
  NAND U9658 ( .A(n37652), .B(n9114), .Z(n8966) );
  NAND U9659 ( .A(n8967), .B(n8966), .Z(n9117) );
  XNOR U9660 ( .A(n9118), .B(n9117), .Z(n9119) );
  XOR U9661 ( .A(n9120), .B(n9119), .Z(n9154) );
  XOR U9662 ( .A(n9153), .B(n9154), .Z(n9156) );
  XOR U9663 ( .A(n9155), .B(n9156), .Z(n9088) );
  NANDN U9664 ( .A(n8969), .B(n8968), .Z(n8973) );
  NANDN U9665 ( .A(n8971), .B(n8970), .Z(n8972) );
  AND U9666 ( .A(n8973), .B(n8972), .Z(n9141) );
  NANDN U9667 ( .A(n8975), .B(n8974), .Z(n8979) );
  NANDN U9668 ( .A(n8977), .B(n8976), .Z(n8978) );
  NAND U9669 ( .A(n8979), .B(n8978), .Z(n9142) );
  XNOR U9670 ( .A(n9141), .B(n9142), .Z(n9143) );
  NANDN U9671 ( .A(n8981), .B(n8980), .Z(n8985) );
  NANDN U9672 ( .A(n8983), .B(n8982), .Z(n8984) );
  NAND U9673 ( .A(n8985), .B(n8984), .Z(n9144) );
  XNOR U9674 ( .A(n9143), .B(n9144), .Z(n9087) );
  XNOR U9675 ( .A(n9088), .B(n9087), .Z(n9090) );
  NANDN U9676 ( .A(n8987), .B(n8986), .Z(n8991) );
  NANDN U9677 ( .A(n8989), .B(n8988), .Z(n8990) );
  AND U9678 ( .A(n8991), .B(n8990), .Z(n9089) );
  XOR U9679 ( .A(n9090), .B(n9089), .Z(n9204) );
  NANDN U9680 ( .A(n8993), .B(n8992), .Z(n8997) );
  NANDN U9681 ( .A(n8995), .B(n8994), .Z(n8996) );
  AND U9682 ( .A(n8997), .B(n8996), .Z(n9201) );
  NANDN U9683 ( .A(n8999), .B(n8998), .Z(n9003) );
  NANDN U9684 ( .A(n9001), .B(n9000), .Z(n9002) );
  AND U9685 ( .A(n9003), .B(n9002), .Z(n9084) );
  NANDN U9686 ( .A(n9005), .B(n9004), .Z(n9009) );
  OR U9687 ( .A(n9007), .B(n9006), .Z(n9008) );
  AND U9688 ( .A(n9009), .B(n9008), .Z(n9082) );
  NANDN U9689 ( .A(n9011), .B(n9010), .Z(n9015) );
  NANDN U9690 ( .A(n9013), .B(n9012), .Z(n9014) );
  AND U9691 ( .A(n9015), .B(n9014), .Z(n9148) );
  NANDN U9692 ( .A(n9017), .B(n9016), .Z(n9021) );
  NANDN U9693 ( .A(n9019), .B(n9018), .Z(n9020) );
  NAND U9694 ( .A(n9021), .B(n9020), .Z(n9147) );
  XNOR U9695 ( .A(n9148), .B(n9147), .Z(n9149) );
  NAND U9696 ( .A(b[0]), .B(a[75]), .Z(n9022) );
  XNOR U9697 ( .A(b[1]), .B(n9022), .Z(n9024) );
  NANDN U9698 ( .A(b[0]), .B(a[74]), .Z(n9023) );
  NAND U9699 ( .A(n9024), .B(n9023), .Z(n9096) );
  NAND U9700 ( .A(n194), .B(n9025), .Z(n9027) );
  XOR U9701 ( .A(b[29]), .B(a[47]), .Z(n9171) );
  NAND U9702 ( .A(n38456), .B(n9171), .Z(n9026) );
  AND U9703 ( .A(n9027), .B(n9026), .Z(n9094) );
  AND U9704 ( .A(b[31]), .B(a[43]), .Z(n9093) );
  XNOR U9705 ( .A(n9094), .B(n9093), .Z(n9095) );
  XNOR U9706 ( .A(n9096), .B(n9095), .Z(n9135) );
  NAND U9707 ( .A(n38185), .B(n9028), .Z(n9030) );
  XOR U9708 ( .A(b[23]), .B(a[53]), .Z(n9177) );
  NAND U9709 ( .A(n38132), .B(n9177), .Z(n9029) );
  AND U9710 ( .A(n9030), .B(n9029), .Z(n9168) );
  NAND U9711 ( .A(n184), .B(n9031), .Z(n9033) );
  XOR U9712 ( .A(b[7]), .B(a[69]), .Z(n9180) );
  NAND U9713 ( .A(n36592), .B(n9180), .Z(n9032) );
  AND U9714 ( .A(n9033), .B(n9032), .Z(n9166) );
  NAND U9715 ( .A(n38289), .B(n9034), .Z(n9036) );
  XOR U9716 ( .A(b[25]), .B(a[51]), .Z(n9183) );
  NAND U9717 ( .A(n38247), .B(n9183), .Z(n9035) );
  NAND U9718 ( .A(n9036), .B(n9035), .Z(n9165) );
  XNOR U9719 ( .A(n9166), .B(n9165), .Z(n9167) );
  XOR U9720 ( .A(n9168), .B(n9167), .Z(n9136) );
  XNOR U9721 ( .A(n9135), .B(n9136), .Z(n9137) );
  NAND U9722 ( .A(n187), .B(n9037), .Z(n9039) );
  XOR U9723 ( .A(b[13]), .B(a[63]), .Z(n9186) );
  NAND U9724 ( .A(n37295), .B(n9186), .Z(n9038) );
  AND U9725 ( .A(n9039), .B(n9038), .Z(n9130) );
  NAND U9726 ( .A(n186), .B(n9040), .Z(n9042) );
  XOR U9727 ( .A(b[11]), .B(a[65]), .Z(n9189) );
  NAND U9728 ( .A(n37097), .B(n9189), .Z(n9041) );
  NAND U9729 ( .A(n9042), .B(n9041), .Z(n9129) );
  XNOR U9730 ( .A(n9130), .B(n9129), .Z(n9131) );
  NAND U9731 ( .A(n188), .B(n9043), .Z(n9045) );
  XOR U9732 ( .A(b[15]), .B(a[61]), .Z(n9192) );
  NAND U9733 ( .A(n37382), .B(n9192), .Z(n9044) );
  AND U9734 ( .A(n9045), .B(n9044), .Z(n9126) );
  NAND U9735 ( .A(n38064), .B(n9046), .Z(n9048) );
  XOR U9736 ( .A(b[21]), .B(a[55]), .Z(n9195) );
  NAND U9737 ( .A(n37993), .B(n9195), .Z(n9047) );
  AND U9738 ( .A(n9048), .B(n9047), .Z(n9124) );
  NAND U9739 ( .A(n185), .B(n9049), .Z(n9051) );
  XOR U9740 ( .A(b[9]), .B(a[67]), .Z(n9198) );
  NAND U9741 ( .A(n36805), .B(n9198), .Z(n9050) );
  NAND U9742 ( .A(n9051), .B(n9050), .Z(n9123) );
  XNOR U9743 ( .A(n9124), .B(n9123), .Z(n9125) );
  XOR U9744 ( .A(n9126), .B(n9125), .Z(n9132) );
  XOR U9745 ( .A(n9131), .B(n9132), .Z(n9138) );
  XOR U9746 ( .A(n9137), .B(n9138), .Z(n9150) );
  XNOR U9747 ( .A(n9149), .B(n9150), .Z(n9081) );
  XNOR U9748 ( .A(n9082), .B(n9081), .Z(n9083) );
  XOR U9749 ( .A(n9084), .B(n9083), .Z(n9202) );
  XNOR U9750 ( .A(n9201), .B(n9202), .Z(n9203) );
  XNOR U9751 ( .A(n9204), .B(n9203), .Z(n9209) );
  XOR U9752 ( .A(n9210), .B(n9209), .Z(n9076) );
  NANDN U9753 ( .A(n9053), .B(n9052), .Z(n9057) );
  NANDN U9754 ( .A(n9055), .B(n9054), .Z(n9056) );
  AND U9755 ( .A(n9057), .B(n9056), .Z(n9075) );
  XNOR U9756 ( .A(n9076), .B(n9075), .Z(n9077) );
  NANDN U9757 ( .A(n9059), .B(n9058), .Z(n9063) );
  NAND U9758 ( .A(n9061), .B(n9060), .Z(n9062) );
  NAND U9759 ( .A(n9063), .B(n9062), .Z(n9078) );
  XNOR U9760 ( .A(n9077), .B(n9078), .Z(n9069) );
  XNOR U9761 ( .A(n9070), .B(n9069), .Z(n9071) );
  XNOR U9762 ( .A(n9072), .B(n9071), .Z(n9213) );
  XNOR U9763 ( .A(sreg[299]), .B(n9213), .Z(n9215) );
  NANDN U9764 ( .A(sreg[298]), .B(n9064), .Z(n9068) );
  NAND U9765 ( .A(n9066), .B(n9065), .Z(n9067) );
  NAND U9766 ( .A(n9068), .B(n9067), .Z(n9214) );
  XNOR U9767 ( .A(n9215), .B(n9214), .Z(c[299]) );
  NANDN U9768 ( .A(n9070), .B(n9069), .Z(n9074) );
  NANDN U9769 ( .A(n9072), .B(n9071), .Z(n9073) );
  AND U9770 ( .A(n9074), .B(n9073), .Z(n9221) );
  NANDN U9771 ( .A(n9076), .B(n9075), .Z(n9080) );
  NANDN U9772 ( .A(n9078), .B(n9077), .Z(n9079) );
  AND U9773 ( .A(n9080), .B(n9079), .Z(n9219) );
  NANDN U9774 ( .A(n9082), .B(n9081), .Z(n9086) );
  NANDN U9775 ( .A(n9084), .B(n9083), .Z(n9085) );
  AND U9776 ( .A(n9086), .B(n9085), .Z(n9231) );
  NANDN U9777 ( .A(n9088), .B(n9087), .Z(n9092) );
  NAND U9778 ( .A(n9090), .B(n9089), .Z(n9091) );
  AND U9779 ( .A(n9092), .B(n9091), .Z(n9230) );
  XNOR U9780 ( .A(n9231), .B(n9230), .Z(n9233) );
  NANDN U9781 ( .A(n9094), .B(n9093), .Z(n9098) );
  NANDN U9782 ( .A(n9096), .B(n9095), .Z(n9097) );
  AND U9783 ( .A(n9098), .B(n9097), .Z(n9308) );
  NAND U9784 ( .A(n38385), .B(n9099), .Z(n9101) );
  XOR U9785 ( .A(b[27]), .B(a[50]), .Z(n9254) );
  NAND U9786 ( .A(n38343), .B(n9254), .Z(n9100) );
  AND U9787 ( .A(n9101), .B(n9100), .Z(n9315) );
  NAND U9788 ( .A(n183), .B(n9102), .Z(n9104) );
  XOR U9789 ( .A(b[5]), .B(a[72]), .Z(n9257) );
  NAND U9790 ( .A(n36296), .B(n9257), .Z(n9103) );
  AND U9791 ( .A(n9104), .B(n9103), .Z(n9313) );
  NAND U9792 ( .A(n190), .B(n9105), .Z(n9107) );
  XOR U9793 ( .A(b[19]), .B(a[58]), .Z(n9260) );
  NAND U9794 ( .A(n37821), .B(n9260), .Z(n9106) );
  NAND U9795 ( .A(n9107), .B(n9106), .Z(n9312) );
  XNOR U9796 ( .A(n9313), .B(n9312), .Z(n9314) );
  XNOR U9797 ( .A(n9315), .B(n9314), .Z(n9306) );
  NAND U9798 ( .A(n38470), .B(n9108), .Z(n9110) );
  XOR U9799 ( .A(b[31]), .B(a[46]), .Z(n9263) );
  NAND U9800 ( .A(n38453), .B(n9263), .Z(n9109) );
  AND U9801 ( .A(n9110), .B(n9109), .Z(n9275) );
  NAND U9802 ( .A(n181), .B(n9111), .Z(n9113) );
  XOR U9803 ( .A(b[3]), .B(a[74]), .Z(n9266) );
  NAND U9804 ( .A(n182), .B(n9266), .Z(n9112) );
  AND U9805 ( .A(n9113), .B(n9112), .Z(n9273) );
  NAND U9806 ( .A(n189), .B(n9114), .Z(n9116) );
  XOR U9807 ( .A(b[17]), .B(a[60]), .Z(n9269) );
  NAND U9808 ( .A(n37652), .B(n9269), .Z(n9115) );
  NAND U9809 ( .A(n9116), .B(n9115), .Z(n9272) );
  XNOR U9810 ( .A(n9273), .B(n9272), .Z(n9274) );
  XOR U9811 ( .A(n9275), .B(n9274), .Z(n9307) );
  XOR U9812 ( .A(n9306), .B(n9307), .Z(n9309) );
  XOR U9813 ( .A(n9308), .B(n9309), .Z(n9243) );
  NANDN U9814 ( .A(n9118), .B(n9117), .Z(n9122) );
  NANDN U9815 ( .A(n9120), .B(n9119), .Z(n9121) );
  AND U9816 ( .A(n9122), .B(n9121), .Z(n9296) );
  NANDN U9817 ( .A(n9124), .B(n9123), .Z(n9128) );
  NANDN U9818 ( .A(n9126), .B(n9125), .Z(n9127) );
  NAND U9819 ( .A(n9128), .B(n9127), .Z(n9297) );
  XNOR U9820 ( .A(n9296), .B(n9297), .Z(n9298) );
  NANDN U9821 ( .A(n9130), .B(n9129), .Z(n9134) );
  NANDN U9822 ( .A(n9132), .B(n9131), .Z(n9133) );
  NAND U9823 ( .A(n9134), .B(n9133), .Z(n9299) );
  XNOR U9824 ( .A(n9298), .B(n9299), .Z(n9242) );
  XNOR U9825 ( .A(n9243), .B(n9242), .Z(n9245) );
  NANDN U9826 ( .A(n9136), .B(n9135), .Z(n9140) );
  NANDN U9827 ( .A(n9138), .B(n9137), .Z(n9139) );
  AND U9828 ( .A(n9140), .B(n9139), .Z(n9244) );
  XOR U9829 ( .A(n9245), .B(n9244), .Z(n9357) );
  NANDN U9830 ( .A(n9142), .B(n9141), .Z(n9146) );
  NANDN U9831 ( .A(n9144), .B(n9143), .Z(n9145) );
  AND U9832 ( .A(n9146), .B(n9145), .Z(n9354) );
  NANDN U9833 ( .A(n9148), .B(n9147), .Z(n9152) );
  NANDN U9834 ( .A(n9150), .B(n9149), .Z(n9151) );
  AND U9835 ( .A(n9152), .B(n9151), .Z(n9239) );
  NANDN U9836 ( .A(n9154), .B(n9153), .Z(n9158) );
  OR U9837 ( .A(n9156), .B(n9155), .Z(n9157) );
  AND U9838 ( .A(n9158), .B(n9157), .Z(n9237) );
  NANDN U9839 ( .A(n9160), .B(n9159), .Z(n9164) );
  NANDN U9840 ( .A(n9162), .B(n9161), .Z(n9163) );
  AND U9841 ( .A(n9164), .B(n9163), .Z(n9303) );
  NANDN U9842 ( .A(n9166), .B(n9165), .Z(n9170) );
  NANDN U9843 ( .A(n9168), .B(n9167), .Z(n9169) );
  NAND U9844 ( .A(n9170), .B(n9169), .Z(n9302) );
  XNOR U9845 ( .A(n9303), .B(n9302), .Z(n9305) );
  NAND U9846 ( .A(n194), .B(n9171), .Z(n9173) );
  XOR U9847 ( .A(b[29]), .B(a[48]), .Z(n9327) );
  NAND U9848 ( .A(n38456), .B(n9327), .Z(n9172) );
  AND U9849 ( .A(n9173), .B(n9172), .Z(n9249) );
  AND U9850 ( .A(b[31]), .B(a[44]), .Z(n9248) );
  XNOR U9851 ( .A(n9249), .B(n9248), .Z(n9250) );
  NAND U9852 ( .A(b[0]), .B(a[76]), .Z(n9174) );
  XNOR U9853 ( .A(b[1]), .B(n9174), .Z(n9176) );
  NANDN U9854 ( .A(b[0]), .B(a[75]), .Z(n9175) );
  NAND U9855 ( .A(n9176), .B(n9175), .Z(n9251) );
  XNOR U9856 ( .A(n9250), .B(n9251), .Z(n9291) );
  NAND U9857 ( .A(n38185), .B(n9177), .Z(n9179) );
  XOR U9858 ( .A(b[23]), .B(a[54]), .Z(n9330) );
  NAND U9859 ( .A(n38132), .B(n9330), .Z(n9178) );
  AND U9860 ( .A(n9179), .B(n9178), .Z(n9320) );
  NAND U9861 ( .A(n184), .B(n9180), .Z(n9182) );
  XOR U9862 ( .A(b[7]), .B(a[70]), .Z(n9333) );
  NAND U9863 ( .A(n36592), .B(n9333), .Z(n9181) );
  AND U9864 ( .A(n9182), .B(n9181), .Z(n9319) );
  NAND U9865 ( .A(n38289), .B(n9183), .Z(n9185) );
  XOR U9866 ( .A(b[25]), .B(a[52]), .Z(n9336) );
  NAND U9867 ( .A(n38247), .B(n9336), .Z(n9184) );
  NAND U9868 ( .A(n9185), .B(n9184), .Z(n9318) );
  XOR U9869 ( .A(n9319), .B(n9318), .Z(n9321) );
  XOR U9870 ( .A(n9320), .B(n9321), .Z(n9290) );
  XOR U9871 ( .A(n9291), .B(n9290), .Z(n9293) );
  NAND U9872 ( .A(n187), .B(n9186), .Z(n9188) );
  XOR U9873 ( .A(b[13]), .B(a[64]), .Z(n9339) );
  NAND U9874 ( .A(n37295), .B(n9339), .Z(n9187) );
  AND U9875 ( .A(n9188), .B(n9187), .Z(n9285) );
  NAND U9876 ( .A(n186), .B(n9189), .Z(n9191) );
  XOR U9877 ( .A(b[11]), .B(a[66]), .Z(n9342) );
  NAND U9878 ( .A(n37097), .B(n9342), .Z(n9190) );
  NAND U9879 ( .A(n9191), .B(n9190), .Z(n9284) );
  XNOR U9880 ( .A(n9285), .B(n9284), .Z(n9287) );
  NAND U9881 ( .A(n188), .B(n9192), .Z(n9194) );
  XOR U9882 ( .A(b[15]), .B(a[62]), .Z(n9345) );
  NAND U9883 ( .A(n37382), .B(n9345), .Z(n9193) );
  AND U9884 ( .A(n9194), .B(n9193), .Z(n9281) );
  NAND U9885 ( .A(n38064), .B(n9195), .Z(n9197) );
  XOR U9886 ( .A(b[21]), .B(a[56]), .Z(n9348) );
  NAND U9887 ( .A(n37993), .B(n9348), .Z(n9196) );
  AND U9888 ( .A(n9197), .B(n9196), .Z(n9279) );
  NAND U9889 ( .A(n185), .B(n9198), .Z(n9200) );
  XOR U9890 ( .A(b[9]), .B(a[68]), .Z(n9351) );
  NAND U9891 ( .A(n36805), .B(n9351), .Z(n9199) );
  NAND U9892 ( .A(n9200), .B(n9199), .Z(n9278) );
  XNOR U9893 ( .A(n9279), .B(n9278), .Z(n9280) );
  XNOR U9894 ( .A(n9281), .B(n9280), .Z(n9286) );
  XOR U9895 ( .A(n9287), .B(n9286), .Z(n9292) );
  XNOR U9896 ( .A(n9293), .B(n9292), .Z(n9304) );
  XNOR U9897 ( .A(n9305), .B(n9304), .Z(n9236) );
  XNOR U9898 ( .A(n9237), .B(n9236), .Z(n9238) );
  XOR U9899 ( .A(n9239), .B(n9238), .Z(n9355) );
  XNOR U9900 ( .A(n9354), .B(n9355), .Z(n9356) );
  XNOR U9901 ( .A(n9357), .B(n9356), .Z(n9232) );
  XOR U9902 ( .A(n9233), .B(n9232), .Z(n9225) );
  NANDN U9903 ( .A(n9202), .B(n9201), .Z(n9206) );
  NANDN U9904 ( .A(n9204), .B(n9203), .Z(n9205) );
  AND U9905 ( .A(n9206), .B(n9205), .Z(n9224) );
  XNOR U9906 ( .A(n9225), .B(n9224), .Z(n9226) );
  NANDN U9907 ( .A(n9208), .B(n9207), .Z(n9212) );
  NAND U9908 ( .A(n9210), .B(n9209), .Z(n9211) );
  NAND U9909 ( .A(n9212), .B(n9211), .Z(n9227) );
  XNOR U9910 ( .A(n9226), .B(n9227), .Z(n9218) );
  XNOR U9911 ( .A(n9219), .B(n9218), .Z(n9220) );
  XNOR U9912 ( .A(n9221), .B(n9220), .Z(n9360) );
  XNOR U9913 ( .A(sreg[300]), .B(n9360), .Z(n9362) );
  NANDN U9914 ( .A(sreg[299]), .B(n9213), .Z(n9217) );
  NAND U9915 ( .A(n9215), .B(n9214), .Z(n9216) );
  NAND U9916 ( .A(n9217), .B(n9216), .Z(n9361) );
  XNOR U9917 ( .A(n9362), .B(n9361), .Z(c[300]) );
  NANDN U9918 ( .A(n9219), .B(n9218), .Z(n9223) );
  NANDN U9919 ( .A(n9221), .B(n9220), .Z(n9222) );
  AND U9920 ( .A(n9223), .B(n9222), .Z(n9368) );
  NANDN U9921 ( .A(n9225), .B(n9224), .Z(n9229) );
  NANDN U9922 ( .A(n9227), .B(n9226), .Z(n9228) );
  AND U9923 ( .A(n9229), .B(n9228), .Z(n9366) );
  NANDN U9924 ( .A(n9231), .B(n9230), .Z(n9235) );
  NAND U9925 ( .A(n9233), .B(n9232), .Z(n9234) );
  AND U9926 ( .A(n9235), .B(n9234), .Z(n9373) );
  NANDN U9927 ( .A(n9237), .B(n9236), .Z(n9241) );
  NANDN U9928 ( .A(n9239), .B(n9238), .Z(n9240) );
  AND U9929 ( .A(n9241), .B(n9240), .Z(n9502) );
  NANDN U9930 ( .A(n9243), .B(n9242), .Z(n9247) );
  NAND U9931 ( .A(n9245), .B(n9244), .Z(n9246) );
  AND U9932 ( .A(n9247), .B(n9246), .Z(n9501) );
  XNOR U9933 ( .A(n9502), .B(n9501), .Z(n9504) );
  NANDN U9934 ( .A(n9249), .B(n9248), .Z(n9253) );
  NANDN U9935 ( .A(n9251), .B(n9250), .Z(n9252) );
  AND U9936 ( .A(n9253), .B(n9252), .Z(n9437) );
  NAND U9937 ( .A(n38385), .B(n9254), .Z(n9256) );
  XOR U9938 ( .A(b[27]), .B(a[51]), .Z(n9383) );
  NAND U9939 ( .A(n38343), .B(n9383), .Z(n9255) );
  AND U9940 ( .A(n9256), .B(n9255), .Z(n9444) );
  NAND U9941 ( .A(n183), .B(n9257), .Z(n9259) );
  XOR U9942 ( .A(b[5]), .B(a[73]), .Z(n9386) );
  NAND U9943 ( .A(n36296), .B(n9386), .Z(n9258) );
  AND U9944 ( .A(n9259), .B(n9258), .Z(n9442) );
  NAND U9945 ( .A(n190), .B(n9260), .Z(n9262) );
  XOR U9946 ( .A(b[19]), .B(a[59]), .Z(n9389) );
  NAND U9947 ( .A(n37821), .B(n9389), .Z(n9261) );
  NAND U9948 ( .A(n9262), .B(n9261), .Z(n9441) );
  XNOR U9949 ( .A(n9442), .B(n9441), .Z(n9443) );
  XNOR U9950 ( .A(n9444), .B(n9443), .Z(n9435) );
  NAND U9951 ( .A(n38470), .B(n9263), .Z(n9265) );
  XOR U9952 ( .A(b[31]), .B(a[47]), .Z(n9392) );
  NAND U9953 ( .A(n38453), .B(n9392), .Z(n9264) );
  AND U9954 ( .A(n9265), .B(n9264), .Z(n9404) );
  NAND U9955 ( .A(n181), .B(n9266), .Z(n9268) );
  XOR U9956 ( .A(b[3]), .B(a[75]), .Z(n9395) );
  NAND U9957 ( .A(n182), .B(n9395), .Z(n9267) );
  AND U9958 ( .A(n9268), .B(n9267), .Z(n9402) );
  NAND U9959 ( .A(n189), .B(n9269), .Z(n9271) );
  XOR U9960 ( .A(b[17]), .B(a[61]), .Z(n9398) );
  NAND U9961 ( .A(n37652), .B(n9398), .Z(n9270) );
  NAND U9962 ( .A(n9271), .B(n9270), .Z(n9401) );
  XNOR U9963 ( .A(n9402), .B(n9401), .Z(n9403) );
  XOR U9964 ( .A(n9404), .B(n9403), .Z(n9436) );
  XOR U9965 ( .A(n9435), .B(n9436), .Z(n9438) );
  XOR U9966 ( .A(n9437), .B(n9438), .Z(n9484) );
  NANDN U9967 ( .A(n9273), .B(n9272), .Z(n9277) );
  NANDN U9968 ( .A(n9275), .B(n9274), .Z(n9276) );
  AND U9969 ( .A(n9277), .B(n9276), .Z(n9425) );
  NANDN U9970 ( .A(n9279), .B(n9278), .Z(n9283) );
  NANDN U9971 ( .A(n9281), .B(n9280), .Z(n9282) );
  NAND U9972 ( .A(n9283), .B(n9282), .Z(n9426) );
  XNOR U9973 ( .A(n9425), .B(n9426), .Z(n9427) );
  NANDN U9974 ( .A(n9285), .B(n9284), .Z(n9289) );
  NAND U9975 ( .A(n9287), .B(n9286), .Z(n9288) );
  NAND U9976 ( .A(n9289), .B(n9288), .Z(n9428) );
  XNOR U9977 ( .A(n9427), .B(n9428), .Z(n9483) );
  XNOR U9978 ( .A(n9484), .B(n9483), .Z(n9486) );
  NAND U9979 ( .A(n9291), .B(n9290), .Z(n9295) );
  NAND U9980 ( .A(n9293), .B(n9292), .Z(n9294) );
  AND U9981 ( .A(n9295), .B(n9294), .Z(n9485) );
  XOR U9982 ( .A(n9486), .B(n9485), .Z(n9498) );
  NANDN U9983 ( .A(n9297), .B(n9296), .Z(n9301) );
  NANDN U9984 ( .A(n9299), .B(n9298), .Z(n9300) );
  AND U9985 ( .A(n9301), .B(n9300), .Z(n9495) );
  NANDN U9986 ( .A(n9307), .B(n9306), .Z(n9311) );
  OR U9987 ( .A(n9309), .B(n9308), .Z(n9310) );
  AND U9988 ( .A(n9311), .B(n9310), .Z(n9490) );
  NANDN U9989 ( .A(n9313), .B(n9312), .Z(n9317) );
  NANDN U9990 ( .A(n9315), .B(n9314), .Z(n9316) );
  AND U9991 ( .A(n9317), .B(n9316), .Z(n9432) );
  NANDN U9992 ( .A(n9319), .B(n9318), .Z(n9323) );
  OR U9993 ( .A(n9321), .B(n9320), .Z(n9322) );
  NAND U9994 ( .A(n9323), .B(n9322), .Z(n9431) );
  XNOR U9995 ( .A(n9432), .B(n9431), .Z(n9434) );
  NAND U9996 ( .A(b[0]), .B(a[77]), .Z(n9324) );
  XNOR U9997 ( .A(b[1]), .B(n9324), .Z(n9326) );
  NANDN U9998 ( .A(b[0]), .B(a[76]), .Z(n9325) );
  NAND U9999 ( .A(n9326), .B(n9325), .Z(n9380) );
  NAND U10000 ( .A(n194), .B(n9327), .Z(n9329) );
  XOR U10001 ( .A(b[29]), .B(a[49]), .Z(n9453) );
  NAND U10002 ( .A(n38456), .B(n9453), .Z(n9328) );
  AND U10003 ( .A(n9329), .B(n9328), .Z(n9378) );
  AND U10004 ( .A(b[31]), .B(a[45]), .Z(n9377) );
  XNOR U10005 ( .A(n9378), .B(n9377), .Z(n9379) );
  XNOR U10006 ( .A(n9380), .B(n9379), .Z(n9420) );
  NAND U10007 ( .A(n38185), .B(n9330), .Z(n9332) );
  XOR U10008 ( .A(b[23]), .B(a[55]), .Z(n9459) );
  NAND U10009 ( .A(n38132), .B(n9459), .Z(n9331) );
  AND U10010 ( .A(n9332), .B(n9331), .Z(n9449) );
  NAND U10011 ( .A(n184), .B(n9333), .Z(n9335) );
  XOR U10012 ( .A(b[7]), .B(a[71]), .Z(n9462) );
  NAND U10013 ( .A(n36592), .B(n9462), .Z(n9334) );
  AND U10014 ( .A(n9335), .B(n9334), .Z(n9448) );
  NAND U10015 ( .A(n38289), .B(n9336), .Z(n9338) );
  XOR U10016 ( .A(b[25]), .B(a[53]), .Z(n9465) );
  NAND U10017 ( .A(n38247), .B(n9465), .Z(n9337) );
  NAND U10018 ( .A(n9338), .B(n9337), .Z(n9447) );
  XOR U10019 ( .A(n9448), .B(n9447), .Z(n9450) );
  XOR U10020 ( .A(n9449), .B(n9450), .Z(n9419) );
  XOR U10021 ( .A(n9420), .B(n9419), .Z(n9422) );
  NAND U10022 ( .A(n187), .B(n9339), .Z(n9341) );
  XOR U10023 ( .A(b[13]), .B(a[65]), .Z(n9468) );
  NAND U10024 ( .A(n37295), .B(n9468), .Z(n9340) );
  AND U10025 ( .A(n9341), .B(n9340), .Z(n9414) );
  NAND U10026 ( .A(n186), .B(n9342), .Z(n9344) );
  XOR U10027 ( .A(b[11]), .B(a[67]), .Z(n9471) );
  NAND U10028 ( .A(n37097), .B(n9471), .Z(n9343) );
  NAND U10029 ( .A(n9344), .B(n9343), .Z(n9413) );
  XNOR U10030 ( .A(n9414), .B(n9413), .Z(n9416) );
  NAND U10031 ( .A(n188), .B(n9345), .Z(n9347) );
  XOR U10032 ( .A(b[15]), .B(a[63]), .Z(n9474) );
  NAND U10033 ( .A(n37382), .B(n9474), .Z(n9346) );
  AND U10034 ( .A(n9347), .B(n9346), .Z(n9410) );
  NAND U10035 ( .A(n38064), .B(n9348), .Z(n9350) );
  XOR U10036 ( .A(b[21]), .B(a[57]), .Z(n9477) );
  NAND U10037 ( .A(n37993), .B(n9477), .Z(n9349) );
  AND U10038 ( .A(n9350), .B(n9349), .Z(n9408) );
  NAND U10039 ( .A(n185), .B(n9351), .Z(n9353) );
  XOR U10040 ( .A(b[9]), .B(a[69]), .Z(n9480) );
  NAND U10041 ( .A(n36805), .B(n9480), .Z(n9352) );
  NAND U10042 ( .A(n9353), .B(n9352), .Z(n9407) );
  XNOR U10043 ( .A(n9408), .B(n9407), .Z(n9409) );
  XNOR U10044 ( .A(n9410), .B(n9409), .Z(n9415) );
  XOR U10045 ( .A(n9416), .B(n9415), .Z(n9421) );
  XNOR U10046 ( .A(n9422), .B(n9421), .Z(n9433) );
  XNOR U10047 ( .A(n9434), .B(n9433), .Z(n9489) );
  XNOR U10048 ( .A(n9490), .B(n9489), .Z(n9491) );
  XOR U10049 ( .A(n9492), .B(n9491), .Z(n9496) );
  XNOR U10050 ( .A(n9495), .B(n9496), .Z(n9497) );
  XNOR U10051 ( .A(n9498), .B(n9497), .Z(n9503) );
  XOR U10052 ( .A(n9504), .B(n9503), .Z(n9372) );
  NANDN U10053 ( .A(n9355), .B(n9354), .Z(n9359) );
  NANDN U10054 ( .A(n9357), .B(n9356), .Z(n9358) );
  AND U10055 ( .A(n9359), .B(n9358), .Z(n9371) );
  XOR U10056 ( .A(n9372), .B(n9371), .Z(n9374) );
  XNOR U10057 ( .A(n9373), .B(n9374), .Z(n9365) );
  XNOR U10058 ( .A(n9366), .B(n9365), .Z(n9367) );
  XNOR U10059 ( .A(n9368), .B(n9367), .Z(n9507) );
  XNOR U10060 ( .A(sreg[301]), .B(n9507), .Z(n9509) );
  NANDN U10061 ( .A(sreg[300]), .B(n9360), .Z(n9364) );
  NAND U10062 ( .A(n9362), .B(n9361), .Z(n9363) );
  NAND U10063 ( .A(n9364), .B(n9363), .Z(n9508) );
  XNOR U10064 ( .A(n9509), .B(n9508), .Z(c[301]) );
  NANDN U10065 ( .A(n9366), .B(n9365), .Z(n9370) );
  NANDN U10066 ( .A(n9368), .B(n9367), .Z(n9369) );
  AND U10067 ( .A(n9370), .B(n9369), .Z(n9515) );
  NANDN U10068 ( .A(n9372), .B(n9371), .Z(n9376) );
  NANDN U10069 ( .A(n9374), .B(n9373), .Z(n9375) );
  AND U10070 ( .A(n9376), .B(n9375), .Z(n9513) );
  NANDN U10071 ( .A(n9378), .B(n9377), .Z(n9382) );
  NANDN U10072 ( .A(n9380), .B(n9379), .Z(n9381) );
  AND U10073 ( .A(n9382), .B(n9381), .Z(n9590) );
  NAND U10074 ( .A(n38385), .B(n9383), .Z(n9385) );
  XOR U10075 ( .A(b[27]), .B(a[52]), .Z(n9536) );
  NAND U10076 ( .A(n38343), .B(n9536), .Z(n9384) );
  AND U10077 ( .A(n9385), .B(n9384), .Z(n9597) );
  NAND U10078 ( .A(n183), .B(n9386), .Z(n9388) );
  XOR U10079 ( .A(b[5]), .B(a[74]), .Z(n9539) );
  NAND U10080 ( .A(n36296), .B(n9539), .Z(n9387) );
  AND U10081 ( .A(n9388), .B(n9387), .Z(n9595) );
  NAND U10082 ( .A(n190), .B(n9389), .Z(n9391) );
  XOR U10083 ( .A(b[19]), .B(a[60]), .Z(n9542) );
  NAND U10084 ( .A(n37821), .B(n9542), .Z(n9390) );
  NAND U10085 ( .A(n9391), .B(n9390), .Z(n9594) );
  XNOR U10086 ( .A(n9595), .B(n9594), .Z(n9596) );
  XNOR U10087 ( .A(n9597), .B(n9596), .Z(n9588) );
  NAND U10088 ( .A(n38470), .B(n9392), .Z(n9394) );
  XOR U10089 ( .A(b[31]), .B(a[48]), .Z(n9545) );
  NAND U10090 ( .A(n38453), .B(n9545), .Z(n9393) );
  AND U10091 ( .A(n9394), .B(n9393), .Z(n9557) );
  NAND U10092 ( .A(n181), .B(n9395), .Z(n9397) );
  XOR U10093 ( .A(b[3]), .B(a[76]), .Z(n9548) );
  NAND U10094 ( .A(n182), .B(n9548), .Z(n9396) );
  AND U10095 ( .A(n9397), .B(n9396), .Z(n9555) );
  NAND U10096 ( .A(n189), .B(n9398), .Z(n9400) );
  XOR U10097 ( .A(b[17]), .B(a[62]), .Z(n9551) );
  NAND U10098 ( .A(n37652), .B(n9551), .Z(n9399) );
  NAND U10099 ( .A(n9400), .B(n9399), .Z(n9554) );
  XNOR U10100 ( .A(n9555), .B(n9554), .Z(n9556) );
  XOR U10101 ( .A(n9557), .B(n9556), .Z(n9589) );
  XOR U10102 ( .A(n9588), .B(n9589), .Z(n9591) );
  XOR U10103 ( .A(n9590), .B(n9591), .Z(n9637) );
  NANDN U10104 ( .A(n9402), .B(n9401), .Z(n9406) );
  NANDN U10105 ( .A(n9404), .B(n9403), .Z(n9405) );
  AND U10106 ( .A(n9406), .B(n9405), .Z(n9578) );
  NANDN U10107 ( .A(n9408), .B(n9407), .Z(n9412) );
  NANDN U10108 ( .A(n9410), .B(n9409), .Z(n9411) );
  NAND U10109 ( .A(n9412), .B(n9411), .Z(n9579) );
  XNOR U10110 ( .A(n9578), .B(n9579), .Z(n9580) );
  NANDN U10111 ( .A(n9414), .B(n9413), .Z(n9418) );
  NAND U10112 ( .A(n9416), .B(n9415), .Z(n9417) );
  NAND U10113 ( .A(n9418), .B(n9417), .Z(n9581) );
  XNOR U10114 ( .A(n9580), .B(n9581), .Z(n9636) );
  XNOR U10115 ( .A(n9637), .B(n9636), .Z(n9639) );
  NAND U10116 ( .A(n9420), .B(n9419), .Z(n9424) );
  NAND U10117 ( .A(n9422), .B(n9421), .Z(n9423) );
  AND U10118 ( .A(n9424), .B(n9423), .Z(n9638) );
  XOR U10119 ( .A(n9639), .B(n9638), .Z(n9650) );
  NANDN U10120 ( .A(n9426), .B(n9425), .Z(n9430) );
  NANDN U10121 ( .A(n9428), .B(n9427), .Z(n9429) );
  AND U10122 ( .A(n9430), .B(n9429), .Z(n9648) );
  NANDN U10123 ( .A(n9436), .B(n9435), .Z(n9440) );
  OR U10124 ( .A(n9438), .B(n9437), .Z(n9439) );
  AND U10125 ( .A(n9440), .B(n9439), .Z(n9643) );
  NANDN U10126 ( .A(n9442), .B(n9441), .Z(n9446) );
  NANDN U10127 ( .A(n9444), .B(n9443), .Z(n9445) );
  AND U10128 ( .A(n9446), .B(n9445), .Z(n9585) );
  NANDN U10129 ( .A(n9448), .B(n9447), .Z(n9452) );
  OR U10130 ( .A(n9450), .B(n9449), .Z(n9451) );
  NAND U10131 ( .A(n9452), .B(n9451), .Z(n9584) );
  XNOR U10132 ( .A(n9585), .B(n9584), .Z(n9587) );
  NAND U10133 ( .A(n194), .B(n9453), .Z(n9455) );
  XOR U10134 ( .A(b[29]), .B(a[50]), .Z(n9609) );
  NAND U10135 ( .A(n38456), .B(n9609), .Z(n9454) );
  AND U10136 ( .A(n9455), .B(n9454), .Z(n9531) );
  AND U10137 ( .A(b[31]), .B(a[46]), .Z(n9530) );
  XNOR U10138 ( .A(n9531), .B(n9530), .Z(n9532) );
  NAND U10139 ( .A(b[0]), .B(a[78]), .Z(n9456) );
  XNOR U10140 ( .A(b[1]), .B(n9456), .Z(n9458) );
  NANDN U10141 ( .A(b[0]), .B(a[77]), .Z(n9457) );
  NAND U10142 ( .A(n9458), .B(n9457), .Z(n9533) );
  XNOR U10143 ( .A(n9532), .B(n9533), .Z(n9573) );
  NAND U10144 ( .A(n38185), .B(n9459), .Z(n9461) );
  XOR U10145 ( .A(b[23]), .B(a[56]), .Z(n9612) );
  NAND U10146 ( .A(n38132), .B(n9612), .Z(n9460) );
  AND U10147 ( .A(n9461), .B(n9460), .Z(n9602) );
  NAND U10148 ( .A(n184), .B(n9462), .Z(n9464) );
  XOR U10149 ( .A(b[7]), .B(a[72]), .Z(n9615) );
  NAND U10150 ( .A(n36592), .B(n9615), .Z(n9463) );
  AND U10151 ( .A(n9464), .B(n9463), .Z(n9601) );
  NAND U10152 ( .A(n38289), .B(n9465), .Z(n9467) );
  XOR U10153 ( .A(b[25]), .B(a[54]), .Z(n9618) );
  NAND U10154 ( .A(n38247), .B(n9618), .Z(n9466) );
  NAND U10155 ( .A(n9467), .B(n9466), .Z(n9600) );
  XOR U10156 ( .A(n9601), .B(n9600), .Z(n9603) );
  XOR U10157 ( .A(n9602), .B(n9603), .Z(n9572) );
  XOR U10158 ( .A(n9573), .B(n9572), .Z(n9575) );
  NAND U10159 ( .A(n187), .B(n9468), .Z(n9470) );
  XOR U10160 ( .A(b[13]), .B(a[66]), .Z(n9621) );
  NAND U10161 ( .A(n37295), .B(n9621), .Z(n9469) );
  AND U10162 ( .A(n9470), .B(n9469), .Z(n9567) );
  NAND U10163 ( .A(n186), .B(n9471), .Z(n9473) );
  XOR U10164 ( .A(b[11]), .B(a[68]), .Z(n9624) );
  NAND U10165 ( .A(n37097), .B(n9624), .Z(n9472) );
  NAND U10166 ( .A(n9473), .B(n9472), .Z(n9566) );
  XNOR U10167 ( .A(n9567), .B(n9566), .Z(n9569) );
  NAND U10168 ( .A(n188), .B(n9474), .Z(n9476) );
  XOR U10169 ( .A(b[15]), .B(a[64]), .Z(n9627) );
  NAND U10170 ( .A(n37382), .B(n9627), .Z(n9475) );
  AND U10171 ( .A(n9476), .B(n9475), .Z(n9563) );
  NAND U10172 ( .A(n38064), .B(n9477), .Z(n9479) );
  XOR U10173 ( .A(b[21]), .B(a[58]), .Z(n9630) );
  NAND U10174 ( .A(n37993), .B(n9630), .Z(n9478) );
  AND U10175 ( .A(n9479), .B(n9478), .Z(n9561) );
  NAND U10176 ( .A(n185), .B(n9480), .Z(n9482) );
  XOR U10177 ( .A(b[9]), .B(a[70]), .Z(n9633) );
  NAND U10178 ( .A(n36805), .B(n9633), .Z(n9481) );
  NAND U10179 ( .A(n9482), .B(n9481), .Z(n9560) );
  XNOR U10180 ( .A(n9561), .B(n9560), .Z(n9562) );
  XNOR U10181 ( .A(n9563), .B(n9562), .Z(n9568) );
  XOR U10182 ( .A(n9569), .B(n9568), .Z(n9574) );
  XNOR U10183 ( .A(n9575), .B(n9574), .Z(n9586) );
  XNOR U10184 ( .A(n9587), .B(n9586), .Z(n9642) );
  XNOR U10185 ( .A(n9643), .B(n9642), .Z(n9644) );
  XOR U10186 ( .A(n9645), .B(n9644), .Z(n9649) );
  XOR U10187 ( .A(n9648), .B(n9649), .Z(n9651) );
  XOR U10188 ( .A(n9650), .B(n9651), .Z(n9527) );
  NANDN U10189 ( .A(n9484), .B(n9483), .Z(n9488) );
  NAND U10190 ( .A(n9486), .B(n9485), .Z(n9487) );
  AND U10191 ( .A(n9488), .B(n9487), .Z(n9525) );
  NANDN U10192 ( .A(n9490), .B(n9489), .Z(n9494) );
  NANDN U10193 ( .A(n9492), .B(n9491), .Z(n9493) );
  AND U10194 ( .A(n9494), .B(n9493), .Z(n9524) );
  XNOR U10195 ( .A(n9525), .B(n9524), .Z(n9526) );
  XNOR U10196 ( .A(n9527), .B(n9526), .Z(n9518) );
  NANDN U10197 ( .A(n9496), .B(n9495), .Z(n9500) );
  NANDN U10198 ( .A(n9498), .B(n9497), .Z(n9499) );
  NAND U10199 ( .A(n9500), .B(n9499), .Z(n9519) );
  XNOR U10200 ( .A(n9518), .B(n9519), .Z(n9520) );
  NANDN U10201 ( .A(n9502), .B(n9501), .Z(n9506) );
  NAND U10202 ( .A(n9504), .B(n9503), .Z(n9505) );
  NAND U10203 ( .A(n9506), .B(n9505), .Z(n9521) );
  XNOR U10204 ( .A(n9520), .B(n9521), .Z(n9512) );
  XNOR U10205 ( .A(n9513), .B(n9512), .Z(n9514) );
  XNOR U10206 ( .A(n9515), .B(n9514), .Z(n9654) );
  XNOR U10207 ( .A(sreg[302]), .B(n9654), .Z(n9656) );
  NANDN U10208 ( .A(sreg[301]), .B(n9507), .Z(n9511) );
  NAND U10209 ( .A(n9509), .B(n9508), .Z(n9510) );
  NAND U10210 ( .A(n9511), .B(n9510), .Z(n9655) );
  XNOR U10211 ( .A(n9656), .B(n9655), .Z(c[302]) );
  NANDN U10212 ( .A(n9513), .B(n9512), .Z(n9517) );
  NANDN U10213 ( .A(n9515), .B(n9514), .Z(n9516) );
  AND U10214 ( .A(n9517), .B(n9516), .Z(n9662) );
  NANDN U10215 ( .A(n9519), .B(n9518), .Z(n9523) );
  NANDN U10216 ( .A(n9521), .B(n9520), .Z(n9522) );
  AND U10217 ( .A(n9523), .B(n9522), .Z(n9660) );
  NANDN U10218 ( .A(n9525), .B(n9524), .Z(n9529) );
  NANDN U10219 ( .A(n9527), .B(n9526), .Z(n9528) );
  AND U10220 ( .A(n9529), .B(n9528), .Z(n9668) );
  NANDN U10221 ( .A(n9531), .B(n9530), .Z(n9535) );
  NANDN U10222 ( .A(n9533), .B(n9532), .Z(n9534) );
  AND U10223 ( .A(n9535), .B(n9534), .Z(n9737) );
  NAND U10224 ( .A(n38385), .B(n9536), .Z(n9538) );
  XOR U10225 ( .A(b[27]), .B(a[53]), .Z(n9683) );
  NAND U10226 ( .A(n38343), .B(n9683), .Z(n9537) );
  AND U10227 ( .A(n9538), .B(n9537), .Z(n9744) );
  NAND U10228 ( .A(n183), .B(n9539), .Z(n9541) );
  XOR U10229 ( .A(b[5]), .B(a[75]), .Z(n9686) );
  NAND U10230 ( .A(n36296), .B(n9686), .Z(n9540) );
  AND U10231 ( .A(n9541), .B(n9540), .Z(n9742) );
  NAND U10232 ( .A(n190), .B(n9542), .Z(n9544) );
  XOR U10233 ( .A(b[19]), .B(a[61]), .Z(n9689) );
  NAND U10234 ( .A(n37821), .B(n9689), .Z(n9543) );
  NAND U10235 ( .A(n9544), .B(n9543), .Z(n9741) );
  XNOR U10236 ( .A(n9742), .B(n9741), .Z(n9743) );
  XNOR U10237 ( .A(n9744), .B(n9743), .Z(n9735) );
  NAND U10238 ( .A(n38470), .B(n9545), .Z(n9547) );
  XOR U10239 ( .A(b[31]), .B(a[49]), .Z(n9692) );
  NAND U10240 ( .A(n38453), .B(n9692), .Z(n9546) );
  AND U10241 ( .A(n9547), .B(n9546), .Z(n9704) );
  NAND U10242 ( .A(n181), .B(n9548), .Z(n9550) );
  XOR U10243 ( .A(b[3]), .B(a[77]), .Z(n9695) );
  NAND U10244 ( .A(n182), .B(n9695), .Z(n9549) );
  AND U10245 ( .A(n9550), .B(n9549), .Z(n9702) );
  NAND U10246 ( .A(n189), .B(n9551), .Z(n9553) );
  XOR U10247 ( .A(b[17]), .B(a[63]), .Z(n9698) );
  NAND U10248 ( .A(n37652), .B(n9698), .Z(n9552) );
  NAND U10249 ( .A(n9553), .B(n9552), .Z(n9701) );
  XNOR U10250 ( .A(n9702), .B(n9701), .Z(n9703) );
  XOR U10251 ( .A(n9704), .B(n9703), .Z(n9736) );
  XOR U10252 ( .A(n9735), .B(n9736), .Z(n9738) );
  XOR U10253 ( .A(n9737), .B(n9738), .Z(n9784) );
  NANDN U10254 ( .A(n9555), .B(n9554), .Z(n9559) );
  NANDN U10255 ( .A(n9557), .B(n9556), .Z(n9558) );
  AND U10256 ( .A(n9559), .B(n9558), .Z(n9725) );
  NANDN U10257 ( .A(n9561), .B(n9560), .Z(n9565) );
  NANDN U10258 ( .A(n9563), .B(n9562), .Z(n9564) );
  NAND U10259 ( .A(n9565), .B(n9564), .Z(n9726) );
  XNOR U10260 ( .A(n9725), .B(n9726), .Z(n9727) );
  NANDN U10261 ( .A(n9567), .B(n9566), .Z(n9571) );
  NAND U10262 ( .A(n9569), .B(n9568), .Z(n9570) );
  NAND U10263 ( .A(n9571), .B(n9570), .Z(n9728) );
  XNOR U10264 ( .A(n9727), .B(n9728), .Z(n9783) );
  XNOR U10265 ( .A(n9784), .B(n9783), .Z(n9786) );
  NAND U10266 ( .A(n9573), .B(n9572), .Z(n9577) );
  NAND U10267 ( .A(n9575), .B(n9574), .Z(n9576) );
  AND U10268 ( .A(n9577), .B(n9576), .Z(n9785) );
  XOR U10269 ( .A(n9786), .B(n9785), .Z(n9797) );
  NANDN U10270 ( .A(n9579), .B(n9578), .Z(n9583) );
  NANDN U10271 ( .A(n9581), .B(n9580), .Z(n9582) );
  AND U10272 ( .A(n9583), .B(n9582), .Z(n9795) );
  NANDN U10273 ( .A(n9589), .B(n9588), .Z(n9593) );
  OR U10274 ( .A(n9591), .B(n9590), .Z(n9592) );
  AND U10275 ( .A(n9593), .B(n9592), .Z(n9790) );
  NANDN U10276 ( .A(n9595), .B(n9594), .Z(n9599) );
  NANDN U10277 ( .A(n9597), .B(n9596), .Z(n9598) );
  AND U10278 ( .A(n9599), .B(n9598), .Z(n9732) );
  NANDN U10279 ( .A(n9601), .B(n9600), .Z(n9605) );
  OR U10280 ( .A(n9603), .B(n9602), .Z(n9604) );
  NAND U10281 ( .A(n9605), .B(n9604), .Z(n9731) );
  XNOR U10282 ( .A(n9732), .B(n9731), .Z(n9734) );
  NAND U10283 ( .A(b[0]), .B(a[79]), .Z(n9606) );
  XNOR U10284 ( .A(b[1]), .B(n9606), .Z(n9608) );
  NANDN U10285 ( .A(b[0]), .B(a[78]), .Z(n9607) );
  NAND U10286 ( .A(n9608), .B(n9607), .Z(n9680) );
  NAND U10287 ( .A(n194), .B(n9609), .Z(n9611) );
  XOR U10288 ( .A(b[29]), .B(a[51]), .Z(n9753) );
  NAND U10289 ( .A(n38456), .B(n9753), .Z(n9610) );
  AND U10290 ( .A(n9611), .B(n9610), .Z(n9678) );
  AND U10291 ( .A(b[31]), .B(a[47]), .Z(n9677) );
  XNOR U10292 ( .A(n9678), .B(n9677), .Z(n9679) );
  XNOR U10293 ( .A(n9680), .B(n9679), .Z(n9720) );
  NAND U10294 ( .A(n38185), .B(n9612), .Z(n9614) );
  XOR U10295 ( .A(b[23]), .B(a[57]), .Z(n9759) );
  NAND U10296 ( .A(n38132), .B(n9759), .Z(n9613) );
  AND U10297 ( .A(n9614), .B(n9613), .Z(n9749) );
  NAND U10298 ( .A(n184), .B(n9615), .Z(n9617) );
  XOR U10299 ( .A(b[7]), .B(a[73]), .Z(n9762) );
  NAND U10300 ( .A(n36592), .B(n9762), .Z(n9616) );
  AND U10301 ( .A(n9617), .B(n9616), .Z(n9748) );
  NAND U10302 ( .A(n38289), .B(n9618), .Z(n9620) );
  XOR U10303 ( .A(b[25]), .B(a[55]), .Z(n9765) );
  NAND U10304 ( .A(n38247), .B(n9765), .Z(n9619) );
  NAND U10305 ( .A(n9620), .B(n9619), .Z(n9747) );
  XOR U10306 ( .A(n9748), .B(n9747), .Z(n9750) );
  XOR U10307 ( .A(n9749), .B(n9750), .Z(n9719) );
  XOR U10308 ( .A(n9720), .B(n9719), .Z(n9722) );
  NAND U10309 ( .A(n187), .B(n9621), .Z(n9623) );
  XOR U10310 ( .A(b[13]), .B(a[67]), .Z(n9768) );
  NAND U10311 ( .A(n37295), .B(n9768), .Z(n9622) );
  AND U10312 ( .A(n9623), .B(n9622), .Z(n9714) );
  NAND U10313 ( .A(n186), .B(n9624), .Z(n9626) );
  XOR U10314 ( .A(b[11]), .B(a[69]), .Z(n9771) );
  NAND U10315 ( .A(n37097), .B(n9771), .Z(n9625) );
  NAND U10316 ( .A(n9626), .B(n9625), .Z(n9713) );
  XNOR U10317 ( .A(n9714), .B(n9713), .Z(n9716) );
  NAND U10318 ( .A(n188), .B(n9627), .Z(n9629) );
  XOR U10319 ( .A(b[15]), .B(a[65]), .Z(n9774) );
  NAND U10320 ( .A(n37382), .B(n9774), .Z(n9628) );
  AND U10321 ( .A(n9629), .B(n9628), .Z(n9710) );
  NAND U10322 ( .A(n38064), .B(n9630), .Z(n9632) );
  XOR U10323 ( .A(b[21]), .B(a[59]), .Z(n9777) );
  NAND U10324 ( .A(n37993), .B(n9777), .Z(n9631) );
  AND U10325 ( .A(n9632), .B(n9631), .Z(n9708) );
  NAND U10326 ( .A(n185), .B(n9633), .Z(n9635) );
  XOR U10327 ( .A(b[9]), .B(a[71]), .Z(n9780) );
  NAND U10328 ( .A(n36805), .B(n9780), .Z(n9634) );
  NAND U10329 ( .A(n9635), .B(n9634), .Z(n9707) );
  XNOR U10330 ( .A(n9708), .B(n9707), .Z(n9709) );
  XNOR U10331 ( .A(n9710), .B(n9709), .Z(n9715) );
  XOR U10332 ( .A(n9716), .B(n9715), .Z(n9721) );
  XNOR U10333 ( .A(n9722), .B(n9721), .Z(n9733) );
  XNOR U10334 ( .A(n9734), .B(n9733), .Z(n9789) );
  XNOR U10335 ( .A(n9790), .B(n9789), .Z(n9791) );
  XOR U10336 ( .A(n9792), .B(n9791), .Z(n9796) );
  XOR U10337 ( .A(n9795), .B(n9796), .Z(n9798) );
  XOR U10338 ( .A(n9797), .B(n9798), .Z(n9674) );
  NANDN U10339 ( .A(n9637), .B(n9636), .Z(n9641) );
  NAND U10340 ( .A(n9639), .B(n9638), .Z(n9640) );
  AND U10341 ( .A(n9641), .B(n9640), .Z(n9672) );
  NANDN U10342 ( .A(n9643), .B(n9642), .Z(n9647) );
  NANDN U10343 ( .A(n9645), .B(n9644), .Z(n9646) );
  AND U10344 ( .A(n9647), .B(n9646), .Z(n9671) );
  XNOR U10345 ( .A(n9672), .B(n9671), .Z(n9673) );
  XNOR U10346 ( .A(n9674), .B(n9673), .Z(n9665) );
  NANDN U10347 ( .A(n9649), .B(n9648), .Z(n9653) );
  OR U10348 ( .A(n9651), .B(n9650), .Z(n9652) );
  NAND U10349 ( .A(n9653), .B(n9652), .Z(n9666) );
  XNOR U10350 ( .A(n9665), .B(n9666), .Z(n9667) );
  XNOR U10351 ( .A(n9668), .B(n9667), .Z(n9659) );
  XNOR U10352 ( .A(n9660), .B(n9659), .Z(n9661) );
  XNOR U10353 ( .A(n9662), .B(n9661), .Z(n9801) );
  XNOR U10354 ( .A(sreg[303]), .B(n9801), .Z(n9803) );
  NANDN U10355 ( .A(sreg[302]), .B(n9654), .Z(n9658) );
  NAND U10356 ( .A(n9656), .B(n9655), .Z(n9657) );
  NAND U10357 ( .A(n9658), .B(n9657), .Z(n9802) );
  XNOR U10358 ( .A(n9803), .B(n9802), .Z(c[303]) );
  NANDN U10359 ( .A(n9660), .B(n9659), .Z(n9664) );
  NANDN U10360 ( .A(n9662), .B(n9661), .Z(n9663) );
  AND U10361 ( .A(n9664), .B(n9663), .Z(n9809) );
  NANDN U10362 ( .A(n9666), .B(n9665), .Z(n9670) );
  NANDN U10363 ( .A(n9668), .B(n9667), .Z(n9669) );
  AND U10364 ( .A(n9670), .B(n9669), .Z(n9807) );
  NANDN U10365 ( .A(n9672), .B(n9671), .Z(n9676) );
  NANDN U10366 ( .A(n9674), .B(n9673), .Z(n9675) );
  AND U10367 ( .A(n9676), .B(n9675), .Z(n9815) );
  NANDN U10368 ( .A(n9678), .B(n9677), .Z(n9682) );
  NANDN U10369 ( .A(n9680), .B(n9679), .Z(n9681) );
  AND U10370 ( .A(n9682), .B(n9681), .Z(n9886) );
  NAND U10371 ( .A(n38385), .B(n9683), .Z(n9685) );
  XOR U10372 ( .A(b[27]), .B(a[54]), .Z(n9830) );
  NAND U10373 ( .A(n38343), .B(n9830), .Z(n9684) );
  AND U10374 ( .A(n9685), .B(n9684), .Z(n9893) );
  NAND U10375 ( .A(n183), .B(n9686), .Z(n9688) );
  XOR U10376 ( .A(b[5]), .B(a[76]), .Z(n9833) );
  NAND U10377 ( .A(n36296), .B(n9833), .Z(n9687) );
  AND U10378 ( .A(n9688), .B(n9687), .Z(n9891) );
  NAND U10379 ( .A(n190), .B(n9689), .Z(n9691) );
  XOR U10380 ( .A(b[19]), .B(a[62]), .Z(n9836) );
  NAND U10381 ( .A(n37821), .B(n9836), .Z(n9690) );
  NAND U10382 ( .A(n9691), .B(n9690), .Z(n9890) );
  XNOR U10383 ( .A(n9891), .B(n9890), .Z(n9892) );
  XNOR U10384 ( .A(n9893), .B(n9892), .Z(n9884) );
  NAND U10385 ( .A(n38470), .B(n9692), .Z(n9694) );
  XOR U10386 ( .A(b[31]), .B(a[50]), .Z(n9839) );
  NAND U10387 ( .A(n38453), .B(n9839), .Z(n9693) );
  AND U10388 ( .A(n9694), .B(n9693), .Z(n9851) );
  NAND U10389 ( .A(n181), .B(n9695), .Z(n9697) );
  XOR U10390 ( .A(b[3]), .B(a[78]), .Z(n9842) );
  NAND U10391 ( .A(n182), .B(n9842), .Z(n9696) );
  AND U10392 ( .A(n9697), .B(n9696), .Z(n9849) );
  NAND U10393 ( .A(n189), .B(n9698), .Z(n9700) );
  XOR U10394 ( .A(b[17]), .B(a[64]), .Z(n9845) );
  NAND U10395 ( .A(n37652), .B(n9845), .Z(n9699) );
  NAND U10396 ( .A(n9700), .B(n9699), .Z(n9848) );
  XNOR U10397 ( .A(n9849), .B(n9848), .Z(n9850) );
  XOR U10398 ( .A(n9851), .B(n9850), .Z(n9885) );
  XOR U10399 ( .A(n9884), .B(n9885), .Z(n9887) );
  XOR U10400 ( .A(n9886), .B(n9887), .Z(n9933) );
  NANDN U10401 ( .A(n9702), .B(n9701), .Z(n9706) );
  NANDN U10402 ( .A(n9704), .B(n9703), .Z(n9705) );
  AND U10403 ( .A(n9706), .B(n9705), .Z(n9872) );
  NANDN U10404 ( .A(n9708), .B(n9707), .Z(n9712) );
  NANDN U10405 ( .A(n9710), .B(n9709), .Z(n9711) );
  NAND U10406 ( .A(n9712), .B(n9711), .Z(n9873) );
  XNOR U10407 ( .A(n9872), .B(n9873), .Z(n9874) );
  NANDN U10408 ( .A(n9714), .B(n9713), .Z(n9718) );
  NAND U10409 ( .A(n9716), .B(n9715), .Z(n9717) );
  NAND U10410 ( .A(n9718), .B(n9717), .Z(n9875) );
  XNOR U10411 ( .A(n9874), .B(n9875), .Z(n9932) );
  XNOR U10412 ( .A(n9933), .B(n9932), .Z(n9935) );
  NAND U10413 ( .A(n9720), .B(n9719), .Z(n9724) );
  NAND U10414 ( .A(n9722), .B(n9721), .Z(n9723) );
  AND U10415 ( .A(n9724), .B(n9723), .Z(n9934) );
  XOR U10416 ( .A(n9935), .B(n9934), .Z(n9946) );
  NANDN U10417 ( .A(n9726), .B(n9725), .Z(n9730) );
  NANDN U10418 ( .A(n9728), .B(n9727), .Z(n9729) );
  AND U10419 ( .A(n9730), .B(n9729), .Z(n9944) );
  NANDN U10420 ( .A(n9736), .B(n9735), .Z(n9740) );
  OR U10421 ( .A(n9738), .B(n9737), .Z(n9739) );
  AND U10422 ( .A(n9740), .B(n9739), .Z(n9939) );
  NANDN U10423 ( .A(n9742), .B(n9741), .Z(n9746) );
  NANDN U10424 ( .A(n9744), .B(n9743), .Z(n9745) );
  AND U10425 ( .A(n9746), .B(n9745), .Z(n9879) );
  NANDN U10426 ( .A(n9748), .B(n9747), .Z(n9752) );
  OR U10427 ( .A(n9750), .B(n9749), .Z(n9751) );
  NAND U10428 ( .A(n9752), .B(n9751), .Z(n9878) );
  XNOR U10429 ( .A(n9879), .B(n9878), .Z(n9880) );
  NAND U10430 ( .A(n194), .B(n9753), .Z(n9755) );
  XOR U10431 ( .A(b[29]), .B(a[52]), .Z(n9905) );
  NAND U10432 ( .A(n38456), .B(n9905), .Z(n9754) );
  AND U10433 ( .A(n9755), .B(n9754), .Z(n9825) );
  AND U10434 ( .A(b[31]), .B(a[48]), .Z(n9824) );
  XNOR U10435 ( .A(n9825), .B(n9824), .Z(n9826) );
  NAND U10436 ( .A(b[0]), .B(a[80]), .Z(n9756) );
  XNOR U10437 ( .A(b[1]), .B(n9756), .Z(n9758) );
  NANDN U10438 ( .A(b[0]), .B(a[79]), .Z(n9757) );
  NAND U10439 ( .A(n9758), .B(n9757), .Z(n9827) );
  XNOR U10440 ( .A(n9826), .B(n9827), .Z(n9866) );
  NAND U10441 ( .A(n38185), .B(n9759), .Z(n9761) );
  XOR U10442 ( .A(b[23]), .B(a[58]), .Z(n9908) );
  NAND U10443 ( .A(n38132), .B(n9908), .Z(n9760) );
  AND U10444 ( .A(n9761), .B(n9760), .Z(n9899) );
  NAND U10445 ( .A(n184), .B(n9762), .Z(n9764) );
  XOR U10446 ( .A(b[7]), .B(a[74]), .Z(n9911) );
  NAND U10447 ( .A(n36592), .B(n9911), .Z(n9763) );
  AND U10448 ( .A(n9764), .B(n9763), .Z(n9897) );
  NAND U10449 ( .A(n38289), .B(n9765), .Z(n9767) );
  XOR U10450 ( .A(b[25]), .B(a[56]), .Z(n9914) );
  NAND U10451 ( .A(n38247), .B(n9914), .Z(n9766) );
  NAND U10452 ( .A(n9767), .B(n9766), .Z(n9896) );
  XNOR U10453 ( .A(n9897), .B(n9896), .Z(n9898) );
  XOR U10454 ( .A(n9899), .B(n9898), .Z(n9867) );
  XNOR U10455 ( .A(n9866), .B(n9867), .Z(n9868) );
  NAND U10456 ( .A(n187), .B(n9768), .Z(n9770) );
  XOR U10457 ( .A(b[13]), .B(a[68]), .Z(n9917) );
  NAND U10458 ( .A(n37295), .B(n9917), .Z(n9769) );
  AND U10459 ( .A(n9770), .B(n9769), .Z(n9861) );
  NAND U10460 ( .A(n186), .B(n9771), .Z(n9773) );
  XOR U10461 ( .A(b[11]), .B(a[70]), .Z(n9920) );
  NAND U10462 ( .A(n37097), .B(n9920), .Z(n9772) );
  NAND U10463 ( .A(n9773), .B(n9772), .Z(n9860) );
  XNOR U10464 ( .A(n9861), .B(n9860), .Z(n9862) );
  NAND U10465 ( .A(n188), .B(n9774), .Z(n9776) );
  XOR U10466 ( .A(b[15]), .B(a[66]), .Z(n9923) );
  NAND U10467 ( .A(n37382), .B(n9923), .Z(n9775) );
  AND U10468 ( .A(n9776), .B(n9775), .Z(n9857) );
  NAND U10469 ( .A(n38064), .B(n9777), .Z(n9779) );
  XOR U10470 ( .A(b[21]), .B(a[60]), .Z(n9926) );
  NAND U10471 ( .A(n37993), .B(n9926), .Z(n9778) );
  AND U10472 ( .A(n9779), .B(n9778), .Z(n9855) );
  NAND U10473 ( .A(n185), .B(n9780), .Z(n9782) );
  XOR U10474 ( .A(b[9]), .B(a[72]), .Z(n9929) );
  NAND U10475 ( .A(n36805), .B(n9929), .Z(n9781) );
  NAND U10476 ( .A(n9782), .B(n9781), .Z(n9854) );
  XNOR U10477 ( .A(n9855), .B(n9854), .Z(n9856) );
  XOR U10478 ( .A(n9857), .B(n9856), .Z(n9863) );
  XOR U10479 ( .A(n9862), .B(n9863), .Z(n9869) );
  XOR U10480 ( .A(n9868), .B(n9869), .Z(n9881) );
  XNOR U10481 ( .A(n9880), .B(n9881), .Z(n9938) );
  XNOR U10482 ( .A(n9939), .B(n9938), .Z(n9940) );
  XOR U10483 ( .A(n9941), .B(n9940), .Z(n9945) );
  XOR U10484 ( .A(n9944), .B(n9945), .Z(n9947) );
  XOR U10485 ( .A(n9946), .B(n9947), .Z(n9821) );
  NANDN U10486 ( .A(n9784), .B(n9783), .Z(n9788) );
  NAND U10487 ( .A(n9786), .B(n9785), .Z(n9787) );
  AND U10488 ( .A(n9788), .B(n9787), .Z(n9819) );
  NANDN U10489 ( .A(n9790), .B(n9789), .Z(n9794) );
  NANDN U10490 ( .A(n9792), .B(n9791), .Z(n9793) );
  AND U10491 ( .A(n9794), .B(n9793), .Z(n9818) );
  XNOR U10492 ( .A(n9819), .B(n9818), .Z(n9820) );
  XNOR U10493 ( .A(n9821), .B(n9820), .Z(n9812) );
  NANDN U10494 ( .A(n9796), .B(n9795), .Z(n9800) );
  OR U10495 ( .A(n9798), .B(n9797), .Z(n9799) );
  NAND U10496 ( .A(n9800), .B(n9799), .Z(n9813) );
  XNOR U10497 ( .A(n9812), .B(n9813), .Z(n9814) );
  XNOR U10498 ( .A(n9815), .B(n9814), .Z(n9806) );
  XNOR U10499 ( .A(n9807), .B(n9806), .Z(n9808) );
  XNOR U10500 ( .A(n9809), .B(n9808), .Z(n9950) );
  XNOR U10501 ( .A(sreg[304]), .B(n9950), .Z(n9952) );
  NANDN U10502 ( .A(sreg[303]), .B(n9801), .Z(n9805) );
  NAND U10503 ( .A(n9803), .B(n9802), .Z(n9804) );
  NAND U10504 ( .A(n9805), .B(n9804), .Z(n9951) );
  XNOR U10505 ( .A(n9952), .B(n9951), .Z(c[304]) );
  NANDN U10506 ( .A(n9807), .B(n9806), .Z(n9811) );
  NANDN U10507 ( .A(n9809), .B(n9808), .Z(n9810) );
  AND U10508 ( .A(n9811), .B(n9810), .Z(n9958) );
  NANDN U10509 ( .A(n9813), .B(n9812), .Z(n9817) );
  NANDN U10510 ( .A(n9815), .B(n9814), .Z(n9816) );
  AND U10511 ( .A(n9817), .B(n9816), .Z(n9956) );
  NANDN U10512 ( .A(n9819), .B(n9818), .Z(n9823) );
  NANDN U10513 ( .A(n9821), .B(n9820), .Z(n9822) );
  AND U10514 ( .A(n9823), .B(n9822), .Z(n9964) );
  NANDN U10515 ( .A(n9825), .B(n9824), .Z(n9829) );
  NANDN U10516 ( .A(n9827), .B(n9826), .Z(n9828) );
  AND U10517 ( .A(n9829), .B(n9828), .Z(n10045) );
  NAND U10518 ( .A(n38385), .B(n9830), .Z(n9832) );
  XOR U10519 ( .A(b[27]), .B(a[55]), .Z(n9991) );
  NAND U10520 ( .A(n38343), .B(n9991), .Z(n9831) );
  AND U10521 ( .A(n9832), .B(n9831), .Z(n10052) );
  NAND U10522 ( .A(n183), .B(n9833), .Z(n9835) );
  XOR U10523 ( .A(b[5]), .B(a[77]), .Z(n9994) );
  NAND U10524 ( .A(n36296), .B(n9994), .Z(n9834) );
  AND U10525 ( .A(n9835), .B(n9834), .Z(n10050) );
  NAND U10526 ( .A(n190), .B(n9836), .Z(n9838) );
  XOR U10527 ( .A(b[19]), .B(a[63]), .Z(n9997) );
  NAND U10528 ( .A(n37821), .B(n9997), .Z(n9837) );
  NAND U10529 ( .A(n9838), .B(n9837), .Z(n10049) );
  XNOR U10530 ( .A(n10050), .B(n10049), .Z(n10051) );
  XNOR U10531 ( .A(n10052), .B(n10051), .Z(n10043) );
  NAND U10532 ( .A(n38470), .B(n9839), .Z(n9841) );
  XOR U10533 ( .A(b[31]), .B(a[51]), .Z(n10000) );
  NAND U10534 ( .A(n38453), .B(n10000), .Z(n9840) );
  AND U10535 ( .A(n9841), .B(n9840), .Z(n10012) );
  NAND U10536 ( .A(n181), .B(n9842), .Z(n9844) );
  XOR U10537 ( .A(b[3]), .B(a[79]), .Z(n10003) );
  NAND U10538 ( .A(n182), .B(n10003), .Z(n9843) );
  AND U10539 ( .A(n9844), .B(n9843), .Z(n10010) );
  NAND U10540 ( .A(n189), .B(n9845), .Z(n9847) );
  XOR U10541 ( .A(b[17]), .B(a[65]), .Z(n10006) );
  NAND U10542 ( .A(n37652), .B(n10006), .Z(n9846) );
  NAND U10543 ( .A(n9847), .B(n9846), .Z(n10009) );
  XNOR U10544 ( .A(n10010), .B(n10009), .Z(n10011) );
  XOR U10545 ( .A(n10012), .B(n10011), .Z(n10044) );
  XOR U10546 ( .A(n10043), .B(n10044), .Z(n10046) );
  XOR U10547 ( .A(n10045), .B(n10046), .Z(n9980) );
  NANDN U10548 ( .A(n9849), .B(n9848), .Z(n9853) );
  NANDN U10549 ( .A(n9851), .B(n9850), .Z(n9852) );
  AND U10550 ( .A(n9853), .B(n9852), .Z(n10033) );
  NANDN U10551 ( .A(n9855), .B(n9854), .Z(n9859) );
  NANDN U10552 ( .A(n9857), .B(n9856), .Z(n9858) );
  NAND U10553 ( .A(n9859), .B(n9858), .Z(n10034) );
  XNOR U10554 ( .A(n10033), .B(n10034), .Z(n10035) );
  NANDN U10555 ( .A(n9861), .B(n9860), .Z(n9865) );
  NANDN U10556 ( .A(n9863), .B(n9862), .Z(n9864) );
  NAND U10557 ( .A(n9865), .B(n9864), .Z(n10036) );
  XNOR U10558 ( .A(n10035), .B(n10036), .Z(n9979) );
  XNOR U10559 ( .A(n9980), .B(n9979), .Z(n9982) );
  NANDN U10560 ( .A(n9867), .B(n9866), .Z(n9871) );
  NANDN U10561 ( .A(n9869), .B(n9868), .Z(n9870) );
  AND U10562 ( .A(n9871), .B(n9870), .Z(n9981) );
  XOR U10563 ( .A(n9982), .B(n9981), .Z(n10093) );
  NANDN U10564 ( .A(n9873), .B(n9872), .Z(n9877) );
  NANDN U10565 ( .A(n9875), .B(n9874), .Z(n9876) );
  AND U10566 ( .A(n9877), .B(n9876), .Z(n10091) );
  NANDN U10567 ( .A(n9879), .B(n9878), .Z(n9883) );
  NANDN U10568 ( .A(n9881), .B(n9880), .Z(n9882) );
  AND U10569 ( .A(n9883), .B(n9882), .Z(n9976) );
  NANDN U10570 ( .A(n9885), .B(n9884), .Z(n9889) );
  OR U10571 ( .A(n9887), .B(n9886), .Z(n9888) );
  AND U10572 ( .A(n9889), .B(n9888), .Z(n9974) );
  NANDN U10573 ( .A(n9891), .B(n9890), .Z(n9895) );
  NANDN U10574 ( .A(n9893), .B(n9892), .Z(n9894) );
  AND U10575 ( .A(n9895), .B(n9894), .Z(n10040) );
  NANDN U10576 ( .A(n9897), .B(n9896), .Z(n9901) );
  NANDN U10577 ( .A(n9899), .B(n9898), .Z(n9900) );
  NAND U10578 ( .A(n9901), .B(n9900), .Z(n10039) );
  XNOR U10579 ( .A(n10040), .B(n10039), .Z(n10042) );
  NAND U10580 ( .A(b[0]), .B(a[81]), .Z(n9902) );
  XNOR U10581 ( .A(b[1]), .B(n9902), .Z(n9904) );
  NANDN U10582 ( .A(b[0]), .B(a[80]), .Z(n9903) );
  NAND U10583 ( .A(n9904), .B(n9903), .Z(n9988) );
  NAND U10584 ( .A(n194), .B(n9905), .Z(n9907) );
  XOR U10585 ( .A(b[29]), .B(a[53]), .Z(n10064) );
  NAND U10586 ( .A(n38456), .B(n10064), .Z(n9906) );
  AND U10587 ( .A(n9907), .B(n9906), .Z(n9986) );
  AND U10588 ( .A(b[31]), .B(a[49]), .Z(n9985) );
  XNOR U10589 ( .A(n9986), .B(n9985), .Z(n9987) );
  XNOR U10590 ( .A(n9988), .B(n9987), .Z(n10028) );
  NAND U10591 ( .A(n38185), .B(n9908), .Z(n9910) );
  XOR U10592 ( .A(b[23]), .B(a[59]), .Z(n10067) );
  NAND U10593 ( .A(n38132), .B(n10067), .Z(n9909) );
  AND U10594 ( .A(n9910), .B(n9909), .Z(n10057) );
  NAND U10595 ( .A(n184), .B(n9911), .Z(n9913) );
  XOR U10596 ( .A(b[7]), .B(a[75]), .Z(n10070) );
  NAND U10597 ( .A(n36592), .B(n10070), .Z(n9912) );
  AND U10598 ( .A(n9913), .B(n9912), .Z(n10056) );
  NAND U10599 ( .A(n38289), .B(n9914), .Z(n9916) );
  XOR U10600 ( .A(b[25]), .B(a[57]), .Z(n10073) );
  NAND U10601 ( .A(n38247), .B(n10073), .Z(n9915) );
  NAND U10602 ( .A(n9916), .B(n9915), .Z(n10055) );
  XOR U10603 ( .A(n10056), .B(n10055), .Z(n10058) );
  XOR U10604 ( .A(n10057), .B(n10058), .Z(n10027) );
  XOR U10605 ( .A(n10028), .B(n10027), .Z(n10030) );
  NAND U10606 ( .A(n187), .B(n9917), .Z(n9919) );
  XOR U10607 ( .A(b[13]), .B(a[69]), .Z(n10076) );
  NAND U10608 ( .A(n37295), .B(n10076), .Z(n9918) );
  AND U10609 ( .A(n9919), .B(n9918), .Z(n10022) );
  NAND U10610 ( .A(n186), .B(n9920), .Z(n9922) );
  XOR U10611 ( .A(b[11]), .B(a[71]), .Z(n10079) );
  NAND U10612 ( .A(n37097), .B(n10079), .Z(n9921) );
  NAND U10613 ( .A(n9922), .B(n9921), .Z(n10021) );
  XNOR U10614 ( .A(n10022), .B(n10021), .Z(n10024) );
  NAND U10615 ( .A(n188), .B(n9923), .Z(n9925) );
  XOR U10616 ( .A(b[15]), .B(a[67]), .Z(n10082) );
  NAND U10617 ( .A(n37382), .B(n10082), .Z(n9924) );
  AND U10618 ( .A(n9925), .B(n9924), .Z(n10018) );
  NAND U10619 ( .A(n38064), .B(n9926), .Z(n9928) );
  XOR U10620 ( .A(b[21]), .B(a[61]), .Z(n10085) );
  NAND U10621 ( .A(n37993), .B(n10085), .Z(n9927) );
  AND U10622 ( .A(n9928), .B(n9927), .Z(n10016) );
  NAND U10623 ( .A(n185), .B(n9929), .Z(n9931) );
  XOR U10624 ( .A(b[9]), .B(a[73]), .Z(n10088) );
  NAND U10625 ( .A(n36805), .B(n10088), .Z(n9930) );
  NAND U10626 ( .A(n9931), .B(n9930), .Z(n10015) );
  XNOR U10627 ( .A(n10016), .B(n10015), .Z(n10017) );
  XNOR U10628 ( .A(n10018), .B(n10017), .Z(n10023) );
  XOR U10629 ( .A(n10024), .B(n10023), .Z(n10029) );
  XNOR U10630 ( .A(n10030), .B(n10029), .Z(n10041) );
  XNOR U10631 ( .A(n10042), .B(n10041), .Z(n9973) );
  XNOR U10632 ( .A(n9974), .B(n9973), .Z(n9975) );
  XOR U10633 ( .A(n9976), .B(n9975), .Z(n10092) );
  XOR U10634 ( .A(n10091), .B(n10092), .Z(n10094) );
  XOR U10635 ( .A(n10093), .B(n10094), .Z(n9970) );
  NANDN U10636 ( .A(n9933), .B(n9932), .Z(n9937) );
  NAND U10637 ( .A(n9935), .B(n9934), .Z(n9936) );
  AND U10638 ( .A(n9937), .B(n9936), .Z(n9968) );
  NANDN U10639 ( .A(n9939), .B(n9938), .Z(n9943) );
  NANDN U10640 ( .A(n9941), .B(n9940), .Z(n9942) );
  AND U10641 ( .A(n9943), .B(n9942), .Z(n9967) );
  XNOR U10642 ( .A(n9968), .B(n9967), .Z(n9969) );
  XNOR U10643 ( .A(n9970), .B(n9969), .Z(n9961) );
  NANDN U10644 ( .A(n9945), .B(n9944), .Z(n9949) );
  OR U10645 ( .A(n9947), .B(n9946), .Z(n9948) );
  NAND U10646 ( .A(n9949), .B(n9948), .Z(n9962) );
  XNOR U10647 ( .A(n9961), .B(n9962), .Z(n9963) );
  XNOR U10648 ( .A(n9964), .B(n9963), .Z(n9955) );
  XNOR U10649 ( .A(n9956), .B(n9955), .Z(n9957) );
  XNOR U10650 ( .A(n9958), .B(n9957), .Z(n10097) );
  XNOR U10651 ( .A(sreg[305]), .B(n10097), .Z(n10099) );
  NANDN U10652 ( .A(sreg[304]), .B(n9950), .Z(n9954) );
  NAND U10653 ( .A(n9952), .B(n9951), .Z(n9953) );
  NAND U10654 ( .A(n9954), .B(n9953), .Z(n10098) );
  XNOR U10655 ( .A(n10099), .B(n10098), .Z(c[305]) );
  NANDN U10656 ( .A(n9956), .B(n9955), .Z(n9960) );
  NANDN U10657 ( .A(n9958), .B(n9957), .Z(n9959) );
  AND U10658 ( .A(n9960), .B(n9959), .Z(n10105) );
  NANDN U10659 ( .A(n9962), .B(n9961), .Z(n9966) );
  NANDN U10660 ( .A(n9964), .B(n9963), .Z(n9965) );
  AND U10661 ( .A(n9966), .B(n9965), .Z(n10103) );
  NANDN U10662 ( .A(n9968), .B(n9967), .Z(n9972) );
  NANDN U10663 ( .A(n9970), .B(n9969), .Z(n9971) );
  AND U10664 ( .A(n9972), .B(n9971), .Z(n10111) );
  NANDN U10665 ( .A(n9974), .B(n9973), .Z(n9978) );
  NANDN U10666 ( .A(n9976), .B(n9975), .Z(n9977) );
  AND U10667 ( .A(n9978), .B(n9977), .Z(n10239) );
  NANDN U10668 ( .A(n9980), .B(n9979), .Z(n9984) );
  NAND U10669 ( .A(n9982), .B(n9981), .Z(n9983) );
  AND U10670 ( .A(n9984), .B(n9983), .Z(n10238) );
  XNOR U10671 ( .A(n10239), .B(n10238), .Z(n10241) );
  NANDN U10672 ( .A(n9986), .B(n9985), .Z(n9990) );
  NANDN U10673 ( .A(n9988), .B(n9987), .Z(n9989) );
  AND U10674 ( .A(n9990), .B(n9989), .Z(n10174) );
  NAND U10675 ( .A(n38385), .B(n9991), .Z(n9993) );
  XOR U10676 ( .A(b[27]), .B(a[56]), .Z(n10120) );
  NAND U10677 ( .A(n38343), .B(n10120), .Z(n9992) );
  AND U10678 ( .A(n9993), .B(n9992), .Z(n10181) );
  NAND U10679 ( .A(n183), .B(n9994), .Z(n9996) );
  XOR U10680 ( .A(b[5]), .B(a[78]), .Z(n10123) );
  NAND U10681 ( .A(n36296), .B(n10123), .Z(n9995) );
  AND U10682 ( .A(n9996), .B(n9995), .Z(n10179) );
  NAND U10683 ( .A(n190), .B(n9997), .Z(n9999) );
  XOR U10684 ( .A(b[19]), .B(a[64]), .Z(n10126) );
  NAND U10685 ( .A(n37821), .B(n10126), .Z(n9998) );
  NAND U10686 ( .A(n9999), .B(n9998), .Z(n10178) );
  XNOR U10687 ( .A(n10179), .B(n10178), .Z(n10180) );
  XNOR U10688 ( .A(n10181), .B(n10180), .Z(n10172) );
  NAND U10689 ( .A(n38470), .B(n10000), .Z(n10002) );
  XOR U10690 ( .A(b[31]), .B(a[52]), .Z(n10129) );
  NAND U10691 ( .A(n38453), .B(n10129), .Z(n10001) );
  AND U10692 ( .A(n10002), .B(n10001), .Z(n10141) );
  NAND U10693 ( .A(n181), .B(n10003), .Z(n10005) );
  XOR U10694 ( .A(b[3]), .B(a[80]), .Z(n10132) );
  NAND U10695 ( .A(n182), .B(n10132), .Z(n10004) );
  AND U10696 ( .A(n10005), .B(n10004), .Z(n10139) );
  NAND U10697 ( .A(n189), .B(n10006), .Z(n10008) );
  XOR U10698 ( .A(b[17]), .B(a[66]), .Z(n10135) );
  NAND U10699 ( .A(n37652), .B(n10135), .Z(n10007) );
  NAND U10700 ( .A(n10008), .B(n10007), .Z(n10138) );
  XNOR U10701 ( .A(n10139), .B(n10138), .Z(n10140) );
  XOR U10702 ( .A(n10141), .B(n10140), .Z(n10173) );
  XOR U10703 ( .A(n10172), .B(n10173), .Z(n10175) );
  XOR U10704 ( .A(n10174), .B(n10175), .Z(n10221) );
  NANDN U10705 ( .A(n10010), .B(n10009), .Z(n10014) );
  NANDN U10706 ( .A(n10012), .B(n10011), .Z(n10013) );
  AND U10707 ( .A(n10014), .B(n10013), .Z(n10162) );
  NANDN U10708 ( .A(n10016), .B(n10015), .Z(n10020) );
  NANDN U10709 ( .A(n10018), .B(n10017), .Z(n10019) );
  NAND U10710 ( .A(n10020), .B(n10019), .Z(n10163) );
  XNOR U10711 ( .A(n10162), .B(n10163), .Z(n10164) );
  NANDN U10712 ( .A(n10022), .B(n10021), .Z(n10026) );
  NAND U10713 ( .A(n10024), .B(n10023), .Z(n10025) );
  NAND U10714 ( .A(n10026), .B(n10025), .Z(n10165) );
  XNOR U10715 ( .A(n10164), .B(n10165), .Z(n10220) );
  XNOR U10716 ( .A(n10221), .B(n10220), .Z(n10223) );
  NAND U10717 ( .A(n10028), .B(n10027), .Z(n10032) );
  NAND U10718 ( .A(n10030), .B(n10029), .Z(n10031) );
  AND U10719 ( .A(n10032), .B(n10031), .Z(n10222) );
  XOR U10720 ( .A(n10223), .B(n10222), .Z(n10235) );
  NANDN U10721 ( .A(n10034), .B(n10033), .Z(n10038) );
  NANDN U10722 ( .A(n10036), .B(n10035), .Z(n10037) );
  AND U10723 ( .A(n10038), .B(n10037), .Z(n10232) );
  NANDN U10724 ( .A(n10044), .B(n10043), .Z(n10048) );
  OR U10725 ( .A(n10046), .B(n10045), .Z(n10047) );
  AND U10726 ( .A(n10048), .B(n10047), .Z(n10227) );
  NANDN U10727 ( .A(n10050), .B(n10049), .Z(n10054) );
  NANDN U10728 ( .A(n10052), .B(n10051), .Z(n10053) );
  AND U10729 ( .A(n10054), .B(n10053), .Z(n10169) );
  NANDN U10730 ( .A(n10056), .B(n10055), .Z(n10060) );
  OR U10731 ( .A(n10058), .B(n10057), .Z(n10059) );
  NAND U10732 ( .A(n10060), .B(n10059), .Z(n10168) );
  XNOR U10733 ( .A(n10169), .B(n10168), .Z(n10171) );
  NAND U10734 ( .A(b[0]), .B(a[82]), .Z(n10061) );
  XNOR U10735 ( .A(b[1]), .B(n10061), .Z(n10063) );
  NANDN U10736 ( .A(b[0]), .B(a[81]), .Z(n10062) );
  NAND U10737 ( .A(n10063), .B(n10062), .Z(n10117) );
  NAND U10738 ( .A(n194), .B(n10064), .Z(n10066) );
  XOR U10739 ( .A(b[29]), .B(a[54]), .Z(n10193) );
  NAND U10740 ( .A(n38456), .B(n10193), .Z(n10065) );
  AND U10741 ( .A(n10066), .B(n10065), .Z(n10115) );
  AND U10742 ( .A(b[31]), .B(a[50]), .Z(n10114) );
  XNOR U10743 ( .A(n10115), .B(n10114), .Z(n10116) );
  XNOR U10744 ( .A(n10117), .B(n10116), .Z(n10157) );
  NAND U10745 ( .A(n38185), .B(n10067), .Z(n10069) );
  XOR U10746 ( .A(b[23]), .B(a[60]), .Z(n10196) );
  NAND U10747 ( .A(n38132), .B(n10196), .Z(n10068) );
  AND U10748 ( .A(n10069), .B(n10068), .Z(n10186) );
  NAND U10749 ( .A(n184), .B(n10070), .Z(n10072) );
  XOR U10750 ( .A(b[7]), .B(a[76]), .Z(n10199) );
  NAND U10751 ( .A(n36592), .B(n10199), .Z(n10071) );
  AND U10752 ( .A(n10072), .B(n10071), .Z(n10185) );
  NAND U10753 ( .A(n38289), .B(n10073), .Z(n10075) );
  XOR U10754 ( .A(b[25]), .B(a[58]), .Z(n10202) );
  NAND U10755 ( .A(n38247), .B(n10202), .Z(n10074) );
  NAND U10756 ( .A(n10075), .B(n10074), .Z(n10184) );
  XOR U10757 ( .A(n10185), .B(n10184), .Z(n10187) );
  XOR U10758 ( .A(n10186), .B(n10187), .Z(n10156) );
  XOR U10759 ( .A(n10157), .B(n10156), .Z(n10159) );
  NAND U10760 ( .A(n187), .B(n10076), .Z(n10078) );
  XOR U10761 ( .A(b[13]), .B(a[70]), .Z(n10205) );
  NAND U10762 ( .A(n37295), .B(n10205), .Z(n10077) );
  AND U10763 ( .A(n10078), .B(n10077), .Z(n10151) );
  NAND U10764 ( .A(n186), .B(n10079), .Z(n10081) );
  XOR U10765 ( .A(b[11]), .B(a[72]), .Z(n10208) );
  NAND U10766 ( .A(n37097), .B(n10208), .Z(n10080) );
  NAND U10767 ( .A(n10081), .B(n10080), .Z(n10150) );
  XNOR U10768 ( .A(n10151), .B(n10150), .Z(n10153) );
  NAND U10769 ( .A(n188), .B(n10082), .Z(n10084) );
  XOR U10770 ( .A(b[15]), .B(a[68]), .Z(n10211) );
  NAND U10771 ( .A(n37382), .B(n10211), .Z(n10083) );
  AND U10772 ( .A(n10084), .B(n10083), .Z(n10147) );
  NAND U10773 ( .A(n38064), .B(n10085), .Z(n10087) );
  XOR U10774 ( .A(b[21]), .B(a[62]), .Z(n10214) );
  NAND U10775 ( .A(n37993), .B(n10214), .Z(n10086) );
  AND U10776 ( .A(n10087), .B(n10086), .Z(n10145) );
  NAND U10777 ( .A(n185), .B(n10088), .Z(n10090) );
  XOR U10778 ( .A(b[9]), .B(a[74]), .Z(n10217) );
  NAND U10779 ( .A(n36805), .B(n10217), .Z(n10089) );
  NAND U10780 ( .A(n10090), .B(n10089), .Z(n10144) );
  XNOR U10781 ( .A(n10145), .B(n10144), .Z(n10146) );
  XNOR U10782 ( .A(n10147), .B(n10146), .Z(n10152) );
  XOR U10783 ( .A(n10153), .B(n10152), .Z(n10158) );
  XNOR U10784 ( .A(n10159), .B(n10158), .Z(n10170) );
  XNOR U10785 ( .A(n10171), .B(n10170), .Z(n10226) );
  XNOR U10786 ( .A(n10227), .B(n10226), .Z(n10228) );
  XOR U10787 ( .A(n10229), .B(n10228), .Z(n10233) );
  XNOR U10788 ( .A(n10232), .B(n10233), .Z(n10234) );
  XNOR U10789 ( .A(n10235), .B(n10234), .Z(n10240) );
  XOR U10790 ( .A(n10241), .B(n10240), .Z(n10109) );
  NANDN U10791 ( .A(n10092), .B(n10091), .Z(n10096) );
  OR U10792 ( .A(n10094), .B(n10093), .Z(n10095) );
  AND U10793 ( .A(n10096), .B(n10095), .Z(n10108) );
  XNOR U10794 ( .A(n10109), .B(n10108), .Z(n10110) );
  XNOR U10795 ( .A(n10111), .B(n10110), .Z(n10102) );
  XNOR U10796 ( .A(n10103), .B(n10102), .Z(n10104) );
  XNOR U10797 ( .A(n10105), .B(n10104), .Z(n10244) );
  XNOR U10798 ( .A(sreg[306]), .B(n10244), .Z(n10246) );
  NANDN U10799 ( .A(sreg[305]), .B(n10097), .Z(n10101) );
  NAND U10800 ( .A(n10099), .B(n10098), .Z(n10100) );
  NAND U10801 ( .A(n10101), .B(n10100), .Z(n10245) );
  XNOR U10802 ( .A(n10246), .B(n10245), .Z(c[306]) );
  NANDN U10803 ( .A(n10103), .B(n10102), .Z(n10107) );
  NANDN U10804 ( .A(n10105), .B(n10104), .Z(n10106) );
  AND U10805 ( .A(n10107), .B(n10106), .Z(n10252) );
  NANDN U10806 ( .A(n10109), .B(n10108), .Z(n10113) );
  NANDN U10807 ( .A(n10111), .B(n10110), .Z(n10112) );
  AND U10808 ( .A(n10113), .B(n10112), .Z(n10250) );
  NANDN U10809 ( .A(n10115), .B(n10114), .Z(n10119) );
  NANDN U10810 ( .A(n10117), .B(n10116), .Z(n10118) );
  AND U10811 ( .A(n10119), .B(n10118), .Z(n10327) );
  NAND U10812 ( .A(n38385), .B(n10120), .Z(n10122) );
  XOR U10813 ( .A(b[27]), .B(a[57]), .Z(n10273) );
  NAND U10814 ( .A(n38343), .B(n10273), .Z(n10121) );
  AND U10815 ( .A(n10122), .B(n10121), .Z(n10334) );
  NAND U10816 ( .A(n183), .B(n10123), .Z(n10125) );
  XOR U10817 ( .A(b[5]), .B(a[79]), .Z(n10276) );
  NAND U10818 ( .A(n36296), .B(n10276), .Z(n10124) );
  AND U10819 ( .A(n10125), .B(n10124), .Z(n10332) );
  NAND U10820 ( .A(n190), .B(n10126), .Z(n10128) );
  XOR U10821 ( .A(b[19]), .B(a[65]), .Z(n10279) );
  NAND U10822 ( .A(n37821), .B(n10279), .Z(n10127) );
  NAND U10823 ( .A(n10128), .B(n10127), .Z(n10331) );
  XNOR U10824 ( .A(n10332), .B(n10331), .Z(n10333) );
  XNOR U10825 ( .A(n10334), .B(n10333), .Z(n10325) );
  NAND U10826 ( .A(n38470), .B(n10129), .Z(n10131) );
  XOR U10827 ( .A(b[31]), .B(a[53]), .Z(n10282) );
  NAND U10828 ( .A(n38453), .B(n10282), .Z(n10130) );
  AND U10829 ( .A(n10131), .B(n10130), .Z(n10294) );
  NAND U10830 ( .A(n181), .B(n10132), .Z(n10134) );
  XOR U10831 ( .A(b[3]), .B(a[81]), .Z(n10285) );
  NAND U10832 ( .A(n182), .B(n10285), .Z(n10133) );
  AND U10833 ( .A(n10134), .B(n10133), .Z(n10292) );
  NAND U10834 ( .A(n189), .B(n10135), .Z(n10137) );
  XOR U10835 ( .A(b[17]), .B(a[67]), .Z(n10288) );
  NAND U10836 ( .A(n37652), .B(n10288), .Z(n10136) );
  NAND U10837 ( .A(n10137), .B(n10136), .Z(n10291) );
  XNOR U10838 ( .A(n10292), .B(n10291), .Z(n10293) );
  XOR U10839 ( .A(n10294), .B(n10293), .Z(n10326) );
  XOR U10840 ( .A(n10325), .B(n10326), .Z(n10328) );
  XOR U10841 ( .A(n10327), .B(n10328), .Z(n10374) );
  NANDN U10842 ( .A(n10139), .B(n10138), .Z(n10143) );
  NANDN U10843 ( .A(n10141), .B(n10140), .Z(n10142) );
  AND U10844 ( .A(n10143), .B(n10142), .Z(n10315) );
  NANDN U10845 ( .A(n10145), .B(n10144), .Z(n10149) );
  NANDN U10846 ( .A(n10147), .B(n10146), .Z(n10148) );
  NAND U10847 ( .A(n10149), .B(n10148), .Z(n10316) );
  XNOR U10848 ( .A(n10315), .B(n10316), .Z(n10317) );
  NANDN U10849 ( .A(n10151), .B(n10150), .Z(n10155) );
  NAND U10850 ( .A(n10153), .B(n10152), .Z(n10154) );
  NAND U10851 ( .A(n10155), .B(n10154), .Z(n10318) );
  XNOR U10852 ( .A(n10317), .B(n10318), .Z(n10373) );
  XNOR U10853 ( .A(n10374), .B(n10373), .Z(n10376) );
  NAND U10854 ( .A(n10157), .B(n10156), .Z(n10161) );
  NAND U10855 ( .A(n10159), .B(n10158), .Z(n10160) );
  AND U10856 ( .A(n10161), .B(n10160), .Z(n10375) );
  XOR U10857 ( .A(n10376), .B(n10375), .Z(n10387) );
  NANDN U10858 ( .A(n10163), .B(n10162), .Z(n10167) );
  NANDN U10859 ( .A(n10165), .B(n10164), .Z(n10166) );
  AND U10860 ( .A(n10167), .B(n10166), .Z(n10385) );
  NANDN U10861 ( .A(n10173), .B(n10172), .Z(n10177) );
  OR U10862 ( .A(n10175), .B(n10174), .Z(n10176) );
  AND U10863 ( .A(n10177), .B(n10176), .Z(n10380) );
  NANDN U10864 ( .A(n10179), .B(n10178), .Z(n10183) );
  NANDN U10865 ( .A(n10181), .B(n10180), .Z(n10182) );
  AND U10866 ( .A(n10183), .B(n10182), .Z(n10322) );
  NANDN U10867 ( .A(n10185), .B(n10184), .Z(n10189) );
  OR U10868 ( .A(n10187), .B(n10186), .Z(n10188) );
  NAND U10869 ( .A(n10189), .B(n10188), .Z(n10321) );
  XNOR U10870 ( .A(n10322), .B(n10321), .Z(n10324) );
  NAND U10871 ( .A(b[0]), .B(a[83]), .Z(n10190) );
  XNOR U10872 ( .A(b[1]), .B(n10190), .Z(n10192) );
  NANDN U10873 ( .A(b[0]), .B(a[82]), .Z(n10191) );
  NAND U10874 ( .A(n10192), .B(n10191), .Z(n10270) );
  NAND U10875 ( .A(n194), .B(n10193), .Z(n10195) );
  XOR U10876 ( .A(b[29]), .B(a[55]), .Z(n10346) );
  NAND U10877 ( .A(n38456), .B(n10346), .Z(n10194) );
  AND U10878 ( .A(n10195), .B(n10194), .Z(n10268) );
  AND U10879 ( .A(b[31]), .B(a[51]), .Z(n10267) );
  XNOR U10880 ( .A(n10268), .B(n10267), .Z(n10269) );
  XNOR U10881 ( .A(n10270), .B(n10269), .Z(n10310) );
  NAND U10882 ( .A(n38185), .B(n10196), .Z(n10198) );
  XOR U10883 ( .A(b[23]), .B(a[61]), .Z(n10349) );
  NAND U10884 ( .A(n38132), .B(n10349), .Z(n10197) );
  AND U10885 ( .A(n10198), .B(n10197), .Z(n10339) );
  NAND U10886 ( .A(n184), .B(n10199), .Z(n10201) );
  XOR U10887 ( .A(b[7]), .B(a[77]), .Z(n10352) );
  NAND U10888 ( .A(n36592), .B(n10352), .Z(n10200) );
  AND U10889 ( .A(n10201), .B(n10200), .Z(n10338) );
  NAND U10890 ( .A(n38289), .B(n10202), .Z(n10204) );
  XOR U10891 ( .A(b[25]), .B(a[59]), .Z(n10355) );
  NAND U10892 ( .A(n38247), .B(n10355), .Z(n10203) );
  NAND U10893 ( .A(n10204), .B(n10203), .Z(n10337) );
  XOR U10894 ( .A(n10338), .B(n10337), .Z(n10340) );
  XOR U10895 ( .A(n10339), .B(n10340), .Z(n10309) );
  XOR U10896 ( .A(n10310), .B(n10309), .Z(n10312) );
  NAND U10897 ( .A(n187), .B(n10205), .Z(n10207) );
  XOR U10898 ( .A(b[13]), .B(a[71]), .Z(n10358) );
  NAND U10899 ( .A(n37295), .B(n10358), .Z(n10206) );
  AND U10900 ( .A(n10207), .B(n10206), .Z(n10304) );
  NAND U10901 ( .A(n186), .B(n10208), .Z(n10210) );
  XOR U10902 ( .A(b[11]), .B(a[73]), .Z(n10361) );
  NAND U10903 ( .A(n37097), .B(n10361), .Z(n10209) );
  NAND U10904 ( .A(n10210), .B(n10209), .Z(n10303) );
  XNOR U10905 ( .A(n10304), .B(n10303), .Z(n10306) );
  NAND U10906 ( .A(n188), .B(n10211), .Z(n10213) );
  XOR U10907 ( .A(b[15]), .B(a[69]), .Z(n10364) );
  NAND U10908 ( .A(n37382), .B(n10364), .Z(n10212) );
  AND U10909 ( .A(n10213), .B(n10212), .Z(n10300) );
  NAND U10910 ( .A(n38064), .B(n10214), .Z(n10216) );
  XOR U10911 ( .A(b[21]), .B(a[63]), .Z(n10367) );
  NAND U10912 ( .A(n37993), .B(n10367), .Z(n10215) );
  AND U10913 ( .A(n10216), .B(n10215), .Z(n10298) );
  NAND U10914 ( .A(n185), .B(n10217), .Z(n10219) );
  XOR U10915 ( .A(b[9]), .B(a[75]), .Z(n10370) );
  NAND U10916 ( .A(n36805), .B(n10370), .Z(n10218) );
  NAND U10917 ( .A(n10219), .B(n10218), .Z(n10297) );
  XNOR U10918 ( .A(n10298), .B(n10297), .Z(n10299) );
  XNOR U10919 ( .A(n10300), .B(n10299), .Z(n10305) );
  XOR U10920 ( .A(n10306), .B(n10305), .Z(n10311) );
  XNOR U10921 ( .A(n10312), .B(n10311), .Z(n10323) );
  XNOR U10922 ( .A(n10324), .B(n10323), .Z(n10379) );
  XNOR U10923 ( .A(n10380), .B(n10379), .Z(n10381) );
  XOR U10924 ( .A(n10382), .B(n10381), .Z(n10386) );
  XOR U10925 ( .A(n10385), .B(n10386), .Z(n10388) );
  XOR U10926 ( .A(n10387), .B(n10388), .Z(n10264) );
  NANDN U10927 ( .A(n10221), .B(n10220), .Z(n10225) );
  NAND U10928 ( .A(n10223), .B(n10222), .Z(n10224) );
  AND U10929 ( .A(n10225), .B(n10224), .Z(n10262) );
  NANDN U10930 ( .A(n10227), .B(n10226), .Z(n10231) );
  NANDN U10931 ( .A(n10229), .B(n10228), .Z(n10230) );
  AND U10932 ( .A(n10231), .B(n10230), .Z(n10261) );
  XNOR U10933 ( .A(n10262), .B(n10261), .Z(n10263) );
  XNOR U10934 ( .A(n10264), .B(n10263), .Z(n10255) );
  NANDN U10935 ( .A(n10233), .B(n10232), .Z(n10237) );
  NANDN U10936 ( .A(n10235), .B(n10234), .Z(n10236) );
  NAND U10937 ( .A(n10237), .B(n10236), .Z(n10256) );
  XNOR U10938 ( .A(n10255), .B(n10256), .Z(n10257) );
  NANDN U10939 ( .A(n10239), .B(n10238), .Z(n10243) );
  NAND U10940 ( .A(n10241), .B(n10240), .Z(n10242) );
  NAND U10941 ( .A(n10243), .B(n10242), .Z(n10258) );
  XNOR U10942 ( .A(n10257), .B(n10258), .Z(n10249) );
  XNOR U10943 ( .A(n10250), .B(n10249), .Z(n10251) );
  XNOR U10944 ( .A(n10252), .B(n10251), .Z(n10391) );
  XNOR U10945 ( .A(sreg[307]), .B(n10391), .Z(n10393) );
  NANDN U10946 ( .A(sreg[306]), .B(n10244), .Z(n10248) );
  NAND U10947 ( .A(n10246), .B(n10245), .Z(n10247) );
  NAND U10948 ( .A(n10248), .B(n10247), .Z(n10392) );
  XNOR U10949 ( .A(n10393), .B(n10392), .Z(c[307]) );
  NANDN U10950 ( .A(n10250), .B(n10249), .Z(n10254) );
  NANDN U10951 ( .A(n10252), .B(n10251), .Z(n10253) );
  AND U10952 ( .A(n10254), .B(n10253), .Z(n10399) );
  NANDN U10953 ( .A(n10256), .B(n10255), .Z(n10260) );
  NANDN U10954 ( .A(n10258), .B(n10257), .Z(n10259) );
  AND U10955 ( .A(n10260), .B(n10259), .Z(n10397) );
  NANDN U10956 ( .A(n10262), .B(n10261), .Z(n10266) );
  NANDN U10957 ( .A(n10264), .B(n10263), .Z(n10265) );
  AND U10958 ( .A(n10266), .B(n10265), .Z(n10405) );
  NANDN U10959 ( .A(n10268), .B(n10267), .Z(n10272) );
  NANDN U10960 ( .A(n10270), .B(n10269), .Z(n10271) );
  AND U10961 ( .A(n10272), .B(n10271), .Z(n10474) );
  NAND U10962 ( .A(n38385), .B(n10273), .Z(n10275) );
  XOR U10963 ( .A(b[27]), .B(a[58]), .Z(n10420) );
  NAND U10964 ( .A(n38343), .B(n10420), .Z(n10274) );
  AND U10965 ( .A(n10275), .B(n10274), .Z(n10481) );
  NAND U10966 ( .A(n183), .B(n10276), .Z(n10278) );
  XOR U10967 ( .A(b[5]), .B(a[80]), .Z(n10423) );
  NAND U10968 ( .A(n36296), .B(n10423), .Z(n10277) );
  AND U10969 ( .A(n10278), .B(n10277), .Z(n10479) );
  NAND U10970 ( .A(n190), .B(n10279), .Z(n10281) );
  XOR U10971 ( .A(b[19]), .B(a[66]), .Z(n10426) );
  NAND U10972 ( .A(n37821), .B(n10426), .Z(n10280) );
  NAND U10973 ( .A(n10281), .B(n10280), .Z(n10478) );
  XNOR U10974 ( .A(n10479), .B(n10478), .Z(n10480) );
  XNOR U10975 ( .A(n10481), .B(n10480), .Z(n10472) );
  NAND U10976 ( .A(n38470), .B(n10282), .Z(n10284) );
  XOR U10977 ( .A(b[31]), .B(a[54]), .Z(n10429) );
  NAND U10978 ( .A(n38453), .B(n10429), .Z(n10283) );
  AND U10979 ( .A(n10284), .B(n10283), .Z(n10441) );
  NAND U10980 ( .A(n181), .B(n10285), .Z(n10287) );
  XOR U10981 ( .A(b[3]), .B(a[82]), .Z(n10432) );
  NAND U10982 ( .A(n182), .B(n10432), .Z(n10286) );
  AND U10983 ( .A(n10287), .B(n10286), .Z(n10439) );
  NAND U10984 ( .A(n189), .B(n10288), .Z(n10290) );
  XOR U10985 ( .A(b[17]), .B(a[68]), .Z(n10435) );
  NAND U10986 ( .A(n37652), .B(n10435), .Z(n10289) );
  NAND U10987 ( .A(n10290), .B(n10289), .Z(n10438) );
  XNOR U10988 ( .A(n10439), .B(n10438), .Z(n10440) );
  XOR U10989 ( .A(n10441), .B(n10440), .Z(n10473) );
  XOR U10990 ( .A(n10472), .B(n10473), .Z(n10475) );
  XOR U10991 ( .A(n10474), .B(n10475), .Z(n10521) );
  NANDN U10992 ( .A(n10292), .B(n10291), .Z(n10296) );
  NANDN U10993 ( .A(n10294), .B(n10293), .Z(n10295) );
  AND U10994 ( .A(n10296), .B(n10295), .Z(n10462) );
  NANDN U10995 ( .A(n10298), .B(n10297), .Z(n10302) );
  NANDN U10996 ( .A(n10300), .B(n10299), .Z(n10301) );
  NAND U10997 ( .A(n10302), .B(n10301), .Z(n10463) );
  XNOR U10998 ( .A(n10462), .B(n10463), .Z(n10464) );
  NANDN U10999 ( .A(n10304), .B(n10303), .Z(n10308) );
  NAND U11000 ( .A(n10306), .B(n10305), .Z(n10307) );
  NAND U11001 ( .A(n10308), .B(n10307), .Z(n10465) );
  XNOR U11002 ( .A(n10464), .B(n10465), .Z(n10520) );
  XNOR U11003 ( .A(n10521), .B(n10520), .Z(n10523) );
  NAND U11004 ( .A(n10310), .B(n10309), .Z(n10314) );
  NAND U11005 ( .A(n10312), .B(n10311), .Z(n10313) );
  AND U11006 ( .A(n10314), .B(n10313), .Z(n10522) );
  XOR U11007 ( .A(n10523), .B(n10522), .Z(n10534) );
  NANDN U11008 ( .A(n10316), .B(n10315), .Z(n10320) );
  NANDN U11009 ( .A(n10318), .B(n10317), .Z(n10319) );
  AND U11010 ( .A(n10320), .B(n10319), .Z(n10532) );
  NANDN U11011 ( .A(n10326), .B(n10325), .Z(n10330) );
  OR U11012 ( .A(n10328), .B(n10327), .Z(n10329) );
  AND U11013 ( .A(n10330), .B(n10329), .Z(n10527) );
  NANDN U11014 ( .A(n10332), .B(n10331), .Z(n10336) );
  NANDN U11015 ( .A(n10334), .B(n10333), .Z(n10335) );
  AND U11016 ( .A(n10336), .B(n10335), .Z(n10469) );
  NANDN U11017 ( .A(n10338), .B(n10337), .Z(n10342) );
  OR U11018 ( .A(n10340), .B(n10339), .Z(n10341) );
  NAND U11019 ( .A(n10342), .B(n10341), .Z(n10468) );
  XNOR U11020 ( .A(n10469), .B(n10468), .Z(n10471) );
  NAND U11021 ( .A(b[0]), .B(a[84]), .Z(n10343) );
  XNOR U11022 ( .A(b[1]), .B(n10343), .Z(n10345) );
  NANDN U11023 ( .A(b[0]), .B(a[83]), .Z(n10344) );
  NAND U11024 ( .A(n10345), .B(n10344), .Z(n10417) );
  NAND U11025 ( .A(n194), .B(n10346), .Z(n10348) );
  XOR U11026 ( .A(b[29]), .B(a[56]), .Z(n10490) );
  NAND U11027 ( .A(n38456), .B(n10490), .Z(n10347) );
  AND U11028 ( .A(n10348), .B(n10347), .Z(n10415) );
  AND U11029 ( .A(b[31]), .B(a[52]), .Z(n10414) );
  XNOR U11030 ( .A(n10415), .B(n10414), .Z(n10416) );
  XNOR U11031 ( .A(n10417), .B(n10416), .Z(n10457) );
  NAND U11032 ( .A(n38185), .B(n10349), .Z(n10351) );
  XOR U11033 ( .A(b[23]), .B(a[62]), .Z(n10496) );
  NAND U11034 ( .A(n38132), .B(n10496), .Z(n10350) );
  AND U11035 ( .A(n10351), .B(n10350), .Z(n10486) );
  NAND U11036 ( .A(n184), .B(n10352), .Z(n10354) );
  XOR U11037 ( .A(b[7]), .B(a[78]), .Z(n10499) );
  NAND U11038 ( .A(n36592), .B(n10499), .Z(n10353) );
  AND U11039 ( .A(n10354), .B(n10353), .Z(n10485) );
  NAND U11040 ( .A(n38289), .B(n10355), .Z(n10357) );
  XOR U11041 ( .A(b[25]), .B(a[60]), .Z(n10502) );
  NAND U11042 ( .A(n38247), .B(n10502), .Z(n10356) );
  NAND U11043 ( .A(n10357), .B(n10356), .Z(n10484) );
  XOR U11044 ( .A(n10485), .B(n10484), .Z(n10487) );
  XOR U11045 ( .A(n10486), .B(n10487), .Z(n10456) );
  XOR U11046 ( .A(n10457), .B(n10456), .Z(n10459) );
  NAND U11047 ( .A(n187), .B(n10358), .Z(n10360) );
  XOR U11048 ( .A(b[13]), .B(a[72]), .Z(n10505) );
  NAND U11049 ( .A(n37295), .B(n10505), .Z(n10359) );
  AND U11050 ( .A(n10360), .B(n10359), .Z(n10451) );
  NAND U11051 ( .A(n186), .B(n10361), .Z(n10363) );
  XOR U11052 ( .A(b[11]), .B(a[74]), .Z(n10508) );
  NAND U11053 ( .A(n37097), .B(n10508), .Z(n10362) );
  NAND U11054 ( .A(n10363), .B(n10362), .Z(n10450) );
  XNOR U11055 ( .A(n10451), .B(n10450), .Z(n10453) );
  NAND U11056 ( .A(n188), .B(n10364), .Z(n10366) );
  XOR U11057 ( .A(b[15]), .B(a[70]), .Z(n10511) );
  NAND U11058 ( .A(n37382), .B(n10511), .Z(n10365) );
  AND U11059 ( .A(n10366), .B(n10365), .Z(n10447) );
  NAND U11060 ( .A(n38064), .B(n10367), .Z(n10369) );
  XOR U11061 ( .A(b[21]), .B(a[64]), .Z(n10514) );
  NAND U11062 ( .A(n37993), .B(n10514), .Z(n10368) );
  AND U11063 ( .A(n10369), .B(n10368), .Z(n10445) );
  NAND U11064 ( .A(n185), .B(n10370), .Z(n10372) );
  XOR U11065 ( .A(b[9]), .B(a[76]), .Z(n10517) );
  NAND U11066 ( .A(n36805), .B(n10517), .Z(n10371) );
  NAND U11067 ( .A(n10372), .B(n10371), .Z(n10444) );
  XNOR U11068 ( .A(n10445), .B(n10444), .Z(n10446) );
  XNOR U11069 ( .A(n10447), .B(n10446), .Z(n10452) );
  XOR U11070 ( .A(n10453), .B(n10452), .Z(n10458) );
  XNOR U11071 ( .A(n10459), .B(n10458), .Z(n10470) );
  XNOR U11072 ( .A(n10471), .B(n10470), .Z(n10526) );
  XNOR U11073 ( .A(n10527), .B(n10526), .Z(n10528) );
  XOR U11074 ( .A(n10529), .B(n10528), .Z(n10533) );
  XOR U11075 ( .A(n10532), .B(n10533), .Z(n10535) );
  XOR U11076 ( .A(n10534), .B(n10535), .Z(n10411) );
  NANDN U11077 ( .A(n10374), .B(n10373), .Z(n10378) );
  NAND U11078 ( .A(n10376), .B(n10375), .Z(n10377) );
  AND U11079 ( .A(n10378), .B(n10377), .Z(n10409) );
  NANDN U11080 ( .A(n10380), .B(n10379), .Z(n10384) );
  NANDN U11081 ( .A(n10382), .B(n10381), .Z(n10383) );
  AND U11082 ( .A(n10384), .B(n10383), .Z(n10408) );
  XNOR U11083 ( .A(n10409), .B(n10408), .Z(n10410) );
  XNOR U11084 ( .A(n10411), .B(n10410), .Z(n10402) );
  NANDN U11085 ( .A(n10386), .B(n10385), .Z(n10390) );
  OR U11086 ( .A(n10388), .B(n10387), .Z(n10389) );
  NAND U11087 ( .A(n10390), .B(n10389), .Z(n10403) );
  XNOR U11088 ( .A(n10402), .B(n10403), .Z(n10404) );
  XNOR U11089 ( .A(n10405), .B(n10404), .Z(n10396) );
  XNOR U11090 ( .A(n10397), .B(n10396), .Z(n10398) );
  XNOR U11091 ( .A(n10399), .B(n10398), .Z(n10538) );
  XNOR U11092 ( .A(sreg[308]), .B(n10538), .Z(n10540) );
  NANDN U11093 ( .A(sreg[307]), .B(n10391), .Z(n10395) );
  NAND U11094 ( .A(n10393), .B(n10392), .Z(n10394) );
  NAND U11095 ( .A(n10395), .B(n10394), .Z(n10539) );
  XNOR U11096 ( .A(n10540), .B(n10539), .Z(c[308]) );
  NANDN U11097 ( .A(n10397), .B(n10396), .Z(n10401) );
  NANDN U11098 ( .A(n10399), .B(n10398), .Z(n10400) );
  AND U11099 ( .A(n10401), .B(n10400), .Z(n10546) );
  NANDN U11100 ( .A(n10403), .B(n10402), .Z(n10407) );
  NANDN U11101 ( .A(n10405), .B(n10404), .Z(n10406) );
  AND U11102 ( .A(n10407), .B(n10406), .Z(n10544) );
  NANDN U11103 ( .A(n10409), .B(n10408), .Z(n10413) );
  NANDN U11104 ( .A(n10411), .B(n10410), .Z(n10412) );
  AND U11105 ( .A(n10413), .B(n10412), .Z(n10552) );
  NANDN U11106 ( .A(n10415), .B(n10414), .Z(n10419) );
  NANDN U11107 ( .A(n10417), .B(n10416), .Z(n10418) );
  AND U11108 ( .A(n10419), .B(n10418), .Z(n10623) );
  NAND U11109 ( .A(n38385), .B(n10420), .Z(n10422) );
  XOR U11110 ( .A(b[27]), .B(a[59]), .Z(n10567) );
  NAND U11111 ( .A(n38343), .B(n10567), .Z(n10421) );
  AND U11112 ( .A(n10422), .B(n10421), .Z(n10630) );
  NAND U11113 ( .A(n183), .B(n10423), .Z(n10425) );
  XOR U11114 ( .A(b[5]), .B(a[81]), .Z(n10570) );
  NAND U11115 ( .A(n36296), .B(n10570), .Z(n10424) );
  AND U11116 ( .A(n10425), .B(n10424), .Z(n10628) );
  NAND U11117 ( .A(n190), .B(n10426), .Z(n10428) );
  XOR U11118 ( .A(b[19]), .B(a[67]), .Z(n10573) );
  NAND U11119 ( .A(n37821), .B(n10573), .Z(n10427) );
  NAND U11120 ( .A(n10428), .B(n10427), .Z(n10627) );
  XNOR U11121 ( .A(n10628), .B(n10627), .Z(n10629) );
  XNOR U11122 ( .A(n10630), .B(n10629), .Z(n10621) );
  NAND U11123 ( .A(n38470), .B(n10429), .Z(n10431) );
  XOR U11124 ( .A(b[31]), .B(a[55]), .Z(n10576) );
  NAND U11125 ( .A(n38453), .B(n10576), .Z(n10430) );
  AND U11126 ( .A(n10431), .B(n10430), .Z(n10588) );
  NAND U11127 ( .A(n181), .B(n10432), .Z(n10434) );
  XOR U11128 ( .A(b[3]), .B(a[83]), .Z(n10579) );
  NAND U11129 ( .A(n182), .B(n10579), .Z(n10433) );
  AND U11130 ( .A(n10434), .B(n10433), .Z(n10586) );
  NAND U11131 ( .A(n189), .B(n10435), .Z(n10437) );
  XOR U11132 ( .A(b[17]), .B(a[69]), .Z(n10582) );
  NAND U11133 ( .A(n37652), .B(n10582), .Z(n10436) );
  NAND U11134 ( .A(n10437), .B(n10436), .Z(n10585) );
  XNOR U11135 ( .A(n10586), .B(n10585), .Z(n10587) );
  XOR U11136 ( .A(n10588), .B(n10587), .Z(n10622) );
  XOR U11137 ( .A(n10621), .B(n10622), .Z(n10624) );
  XOR U11138 ( .A(n10623), .B(n10624), .Z(n10670) );
  NANDN U11139 ( .A(n10439), .B(n10438), .Z(n10443) );
  NANDN U11140 ( .A(n10441), .B(n10440), .Z(n10442) );
  AND U11141 ( .A(n10443), .B(n10442), .Z(n10609) );
  NANDN U11142 ( .A(n10445), .B(n10444), .Z(n10449) );
  NANDN U11143 ( .A(n10447), .B(n10446), .Z(n10448) );
  NAND U11144 ( .A(n10449), .B(n10448), .Z(n10610) );
  XNOR U11145 ( .A(n10609), .B(n10610), .Z(n10611) );
  NANDN U11146 ( .A(n10451), .B(n10450), .Z(n10455) );
  NAND U11147 ( .A(n10453), .B(n10452), .Z(n10454) );
  NAND U11148 ( .A(n10455), .B(n10454), .Z(n10612) );
  XNOR U11149 ( .A(n10611), .B(n10612), .Z(n10669) );
  XNOR U11150 ( .A(n10670), .B(n10669), .Z(n10672) );
  NAND U11151 ( .A(n10457), .B(n10456), .Z(n10461) );
  NAND U11152 ( .A(n10459), .B(n10458), .Z(n10460) );
  AND U11153 ( .A(n10461), .B(n10460), .Z(n10671) );
  XOR U11154 ( .A(n10672), .B(n10671), .Z(n10683) );
  NANDN U11155 ( .A(n10463), .B(n10462), .Z(n10467) );
  NANDN U11156 ( .A(n10465), .B(n10464), .Z(n10466) );
  AND U11157 ( .A(n10467), .B(n10466), .Z(n10681) );
  NANDN U11158 ( .A(n10473), .B(n10472), .Z(n10477) );
  OR U11159 ( .A(n10475), .B(n10474), .Z(n10476) );
  AND U11160 ( .A(n10477), .B(n10476), .Z(n10676) );
  NANDN U11161 ( .A(n10479), .B(n10478), .Z(n10483) );
  NANDN U11162 ( .A(n10481), .B(n10480), .Z(n10482) );
  AND U11163 ( .A(n10483), .B(n10482), .Z(n10616) );
  NANDN U11164 ( .A(n10485), .B(n10484), .Z(n10489) );
  OR U11165 ( .A(n10487), .B(n10486), .Z(n10488) );
  NAND U11166 ( .A(n10489), .B(n10488), .Z(n10615) );
  XNOR U11167 ( .A(n10616), .B(n10615), .Z(n10617) );
  NAND U11168 ( .A(n194), .B(n10490), .Z(n10492) );
  XOR U11169 ( .A(b[29]), .B(a[57]), .Z(n10639) );
  NAND U11170 ( .A(n38456), .B(n10639), .Z(n10491) );
  AND U11171 ( .A(n10492), .B(n10491), .Z(n10562) );
  AND U11172 ( .A(b[31]), .B(a[53]), .Z(n10561) );
  XNOR U11173 ( .A(n10562), .B(n10561), .Z(n10563) );
  NAND U11174 ( .A(b[0]), .B(a[85]), .Z(n10493) );
  XNOR U11175 ( .A(b[1]), .B(n10493), .Z(n10495) );
  NANDN U11176 ( .A(b[0]), .B(a[84]), .Z(n10494) );
  NAND U11177 ( .A(n10495), .B(n10494), .Z(n10564) );
  XNOR U11178 ( .A(n10563), .B(n10564), .Z(n10603) );
  NAND U11179 ( .A(n38185), .B(n10496), .Z(n10498) );
  XOR U11180 ( .A(b[23]), .B(a[63]), .Z(n10645) );
  NAND U11181 ( .A(n38132), .B(n10645), .Z(n10497) );
  AND U11182 ( .A(n10498), .B(n10497), .Z(n10636) );
  NAND U11183 ( .A(n184), .B(n10499), .Z(n10501) );
  XOR U11184 ( .A(b[7]), .B(a[79]), .Z(n10648) );
  NAND U11185 ( .A(n36592), .B(n10648), .Z(n10500) );
  AND U11186 ( .A(n10501), .B(n10500), .Z(n10634) );
  NAND U11187 ( .A(n38289), .B(n10502), .Z(n10504) );
  XOR U11188 ( .A(b[25]), .B(a[61]), .Z(n10651) );
  NAND U11189 ( .A(n38247), .B(n10651), .Z(n10503) );
  NAND U11190 ( .A(n10504), .B(n10503), .Z(n10633) );
  XNOR U11191 ( .A(n10634), .B(n10633), .Z(n10635) );
  XOR U11192 ( .A(n10636), .B(n10635), .Z(n10604) );
  XNOR U11193 ( .A(n10603), .B(n10604), .Z(n10605) );
  NAND U11194 ( .A(n187), .B(n10505), .Z(n10507) );
  XOR U11195 ( .A(b[13]), .B(a[73]), .Z(n10654) );
  NAND U11196 ( .A(n37295), .B(n10654), .Z(n10506) );
  AND U11197 ( .A(n10507), .B(n10506), .Z(n10598) );
  NAND U11198 ( .A(n186), .B(n10508), .Z(n10510) );
  XOR U11199 ( .A(b[11]), .B(a[75]), .Z(n10657) );
  NAND U11200 ( .A(n37097), .B(n10657), .Z(n10509) );
  NAND U11201 ( .A(n10510), .B(n10509), .Z(n10597) );
  XNOR U11202 ( .A(n10598), .B(n10597), .Z(n10599) );
  NAND U11203 ( .A(n188), .B(n10511), .Z(n10513) );
  XOR U11204 ( .A(b[15]), .B(a[71]), .Z(n10660) );
  NAND U11205 ( .A(n37382), .B(n10660), .Z(n10512) );
  AND U11206 ( .A(n10513), .B(n10512), .Z(n10594) );
  NAND U11207 ( .A(n38064), .B(n10514), .Z(n10516) );
  XOR U11208 ( .A(b[21]), .B(a[65]), .Z(n10663) );
  NAND U11209 ( .A(n37993), .B(n10663), .Z(n10515) );
  AND U11210 ( .A(n10516), .B(n10515), .Z(n10592) );
  NAND U11211 ( .A(n185), .B(n10517), .Z(n10519) );
  XOR U11212 ( .A(b[9]), .B(a[77]), .Z(n10666) );
  NAND U11213 ( .A(n36805), .B(n10666), .Z(n10518) );
  NAND U11214 ( .A(n10519), .B(n10518), .Z(n10591) );
  XNOR U11215 ( .A(n10592), .B(n10591), .Z(n10593) );
  XOR U11216 ( .A(n10594), .B(n10593), .Z(n10600) );
  XOR U11217 ( .A(n10599), .B(n10600), .Z(n10606) );
  XOR U11218 ( .A(n10605), .B(n10606), .Z(n10618) );
  XNOR U11219 ( .A(n10617), .B(n10618), .Z(n10675) );
  XNOR U11220 ( .A(n10676), .B(n10675), .Z(n10677) );
  XOR U11221 ( .A(n10678), .B(n10677), .Z(n10682) );
  XOR U11222 ( .A(n10681), .B(n10682), .Z(n10684) );
  XOR U11223 ( .A(n10683), .B(n10684), .Z(n10558) );
  NANDN U11224 ( .A(n10521), .B(n10520), .Z(n10525) );
  NAND U11225 ( .A(n10523), .B(n10522), .Z(n10524) );
  AND U11226 ( .A(n10525), .B(n10524), .Z(n10556) );
  NANDN U11227 ( .A(n10527), .B(n10526), .Z(n10531) );
  NANDN U11228 ( .A(n10529), .B(n10528), .Z(n10530) );
  AND U11229 ( .A(n10531), .B(n10530), .Z(n10555) );
  XNOR U11230 ( .A(n10556), .B(n10555), .Z(n10557) );
  XNOR U11231 ( .A(n10558), .B(n10557), .Z(n10549) );
  NANDN U11232 ( .A(n10533), .B(n10532), .Z(n10537) );
  OR U11233 ( .A(n10535), .B(n10534), .Z(n10536) );
  NAND U11234 ( .A(n10537), .B(n10536), .Z(n10550) );
  XNOR U11235 ( .A(n10549), .B(n10550), .Z(n10551) );
  XNOR U11236 ( .A(n10552), .B(n10551), .Z(n10543) );
  XNOR U11237 ( .A(n10544), .B(n10543), .Z(n10545) );
  XNOR U11238 ( .A(n10546), .B(n10545), .Z(n10687) );
  XNOR U11239 ( .A(sreg[309]), .B(n10687), .Z(n10689) );
  NANDN U11240 ( .A(sreg[308]), .B(n10538), .Z(n10542) );
  NAND U11241 ( .A(n10540), .B(n10539), .Z(n10541) );
  NAND U11242 ( .A(n10542), .B(n10541), .Z(n10688) );
  XNOR U11243 ( .A(n10689), .B(n10688), .Z(c[309]) );
  NANDN U11244 ( .A(n10544), .B(n10543), .Z(n10548) );
  NANDN U11245 ( .A(n10546), .B(n10545), .Z(n10547) );
  AND U11246 ( .A(n10548), .B(n10547), .Z(n10695) );
  NANDN U11247 ( .A(n10550), .B(n10549), .Z(n10554) );
  NANDN U11248 ( .A(n10552), .B(n10551), .Z(n10553) );
  AND U11249 ( .A(n10554), .B(n10553), .Z(n10693) );
  NANDN U11250 ( .A(n10556), .B(n10555), .Z(n10560) );
  NANDN U11251 ( .A(n10558), .B(n10557), .Z(n10559) );
  AND U11252 ( .A(n10560), .B(n10559), .Z(n10701) );
  NANDN U11253 ( .A(n10562), .B(n10561), .Z(n10566) );
  NANDN U11254 ( .A(n10564), .B(n10563), .Z(n10565) );
  AND U11255 ( .A(n10566), .B(n10565), .Z(n10782) );
  NAND U11256 ( .A(n38385), .B(n10567), .Z(n10569) );
  XOR U11257 ( .A(b[27]), .B(a[60]), .Z(n10728) );
  NAND U11258 ( .A(n38343), .B(n10728), .Z(n10568) );
  AND U11259 ( .A(n10569), .B(n10568), .Z(n10789) );
  NAND U11260 ( .A(n183), .B(n10570), .Z(n10572) );
  XOR U11261 ( .A(b[5]), .B(a[82]), .Z(n10731) );
  NAND U11262 ( .A(n36296), .B(n10731), .Z(n10571) );
  AND U11263 ( .A(n10572), .B(n10571), .Z(n10787) );
  NAND U11264 ( .A(n190), .B(n10573), .Z(n10575) );
  XOR U11265 ( .A(b[19]), .B(a[68]), .Z(n10734) );
  NAND U11266 ( .A(n37821), .B(n10734), .Z(n10574) );
  NAND U11267 ( .A(n10575), .B(n10574), .Z(n10786) );
  XNOR U11268 ( .A(n10787), .B(n10786), .Z(n10788) );
  XNOR U11269 ( .A(n10789), .B(n10788), .Z(n10780) );
  NAND U11270 ( .A(n38470), .B(n10576), .Z(n10578) );
  XOR U11271 ( .A(b[31]), .B(a[56]), .Z(n10737) );
  NAND U11272 ( .A(n38453), .B(n10737), .Z(n10577) );
  AND U11273 ( .A(n10578), .B(n10577), .Z(n10749) );
  NAND U11274 ( .A(n181), .B(n10579), .Z(n10581) );
  XOR U11275 ( .A(b[3]), .B(a[84]), .Z(n10740) );
  NAND U11276 ( .A(n182), .B(n10740), .Z(n10580) );
  AND U11277 ( .A(n10581), .B(n10580), .Z(n10747) );
  NAND U11278 ( .A(n189), .B(n10582), .Z(n10584) );
  XOR U11279 ( .A(b[17]), .B(a[70]), .Z(n10743) );
  NAND U11280 ( .A(n37652), .B(n10743), .Z(n10583) );
  NAND U11281 ( .A(n10584), .B(n10583), .Z(n10746) );
  XNOR U11282 ( .A(n10747), .B(n10746), .Z(n10748) );
  XOR U11283 ( .A(n10749), .B(n10748), .Z(n10781) );
  XOR U11284 ( .A(n10780), .B(n10781), .Z(n10783) );
  XOR U11285 ( .A(n10782), .B(n10783), .Z(n10717) );
  NANDN U11286 ( .A(n10586), .B(n10585), .Z(n10590) );
  NANDN U11287 ( .A(n10588), .B(n10587), .Z(n10589) );
  AND U11288 ( .A(n10590), .B(n10589), .Z(n10770) );
  NANDN U11289 ( .A(n10592), .B(n10591), .Z(n10596) );
  NANDN U11290 ( .A(n10594), .B(n10593), .Z(n10595) );
  NAND U11291 ( .A(n10596), .B(n10595), .Z(n10771) );
  XNOR U11292 ( .A(n10770), .B(n10771), .Z(n10772) );
  NANDN U11293 ( .A(n10598), .B(n10597), .Z(n10602) );
  NANDN U11294 ( .A(n10600), .B(n10599), .Z(n10601) );
  NAND U11295 ( .A(n10602), .B(n10601), .Z(n10773) );
  XNOR U11296 ( .A(n10772), .B(n10773), .Z(n10716) );
  XNOR U11297 ( .A(n10717), .B(n10716), .Z(n10719) );
  NANDN U11298 ( .A(n10604), .B(n10603), .Z(n10608) );
  NANDN U11299 ( .A(n10606), .B(n10605), .Z(n10607) );
  AND U11300 ( .A(n10608), .B(n10607), .Z(n10718) );
  XOR U11301 ( .A(n10719), .B(n10718), .Z(n10830) );
  NANDN U11302 ( .A(n10610), .B(n10609), .Z(n10614) );
  NANDN U11303 ( .A(n10612), .B(n10611), .Z(n10613) );
  AND U11304 ( .A(n10614), .B(n10613), .Z(n10828) );
  NANDN U11305 ( .A(n10616), .B(n10615), .Z(n10620) );
  NANDN U11306 ( .A(n10618), .B(n10617), .Z(n10619) );
  AND U11307 ( .A(n10620), .B(n10619), .Z(n10713) );
  NANDN U11308 ( .A(n10622), .B(n10621), .Z(n10626) );
  OR U11309 ( .A(n10624), .B(n10623), .Z(n10625) );
  AND U11310 ( .A(n10626), .B(n10625), .Z(n10711) );
  NANDN U11311 ( .A(n10628), .B(n10627), .Z(n10632) );
  NANDN U11312 ( .A(n10630), .B(n10629), .Z(n10631) );
  AND U11313 ( .A(n10632), .B(n10631), .Z(n10777) );
  NANDN U11314 ( .A(n10634), .B(n10633), .Z(n10638) );
  NANDN U11315 ( .A(n10636), .B(n10635), .Z(n10637) );
  NAND U11316 ( .A(n10638), .B(n10637), .Z(n10776) );
  XNOR U11317 ( .A(n10777), .B(n10776), .Z(n10779) );
  NAND U11318 ( .A(n194), .B(n10639), .Z(n10641) );
  XOR U11319 ( .A(b[29]), .B(a[58]), .Z(n10798) );
  NAND U11320 ( .A(n38456), .B(n10798), .Z(n10640) );
  AND U11321 ( .A(n10641), .B(n10640), .Z(n10723) );
  AND U11322 ( .A(b[31]), .B(a[54]), .Z(n10722) );
  XNOR U11323 ( .A(n10723), .B(n10722), .Z(n10724) );
  NAND U11324 ( .A(b[0]), .B(a[86]), .Z(n10642) );
  XNOR U11325 ( .A(b[1]), .B(n10642), .Z(n10644) );
  NANDN U11326 ( .A(b[0]), .B(a[85]), .Z(n10643) );
  NAND U11327 ( .A(n10644), .B(n10643), .Z(n10725) );
  XNOR U11328 ( .A(n10724), .B(n10725), .Z(n10765) );
  NAND U11329 ( .A(n38185), .B(n10645), .Z(n10647) );
  XOR U11330 ( .A(b[23]), .B(a[64]), .Z(n10804) );
  NAND U11331 ( .A(n38132), .B(n10804), .Z(n10646) );
  AND U11332 ( .A(n10647), .B(n10646), .Z(n10794) );
  NAND U11333 ( .A(n184), .B(n10648), .Z(n10650) );
  XOR U11334 ( .A(b[7]), .B(a[80]), .Z(n10807) );
  NAND U11335 ( .A(n36592), .B(n10807), .Z(n10649) );
  AND U11336 ( .A(n10650), .B(n10649), .Z(n10793) );
  NAND U11337 ( .A(n38289), .B(n10651), .Z(n10653) );
  XOR U11338 ( .A(b[25]), .B(a[62]), .Z(n10810) );
  NAND U11339 ( .A(n38247), .B(n10810), .Z(n10652) );
  NAND U11340 ( .A(n10653), .B(n10652), .Z(n10792) );
  XOR U11341 ( .A(n10793), .B(n10792), .Z(n10795) );
  XOR U11342 ( .A(n10794), .B(n10795), .Z(n10764) );
  XOR U11343 ( .A(n10765), .B(n10764), .Z(n10767) );
  NAND U11344 ( .A(n187), .B(n10654), .Z(n10656) );
  XOR U11345 ( .A(b[13]), .B(a[74]), .Z(n10813) );
  NAND U11346 ( .A(n37295), .B(n10813), .Z(n10655) );
  AND U11347 ( .A(n10656), .B(n10655), .Z(n10759) );
  NAND U11348 ( .A(n186), .B(n10657), .Z(n10659) );
  XOR U11349 ( .A(b[11]), .B(a[76]), .Z(n10816) );
  NAND U11350 ( .A(n37097), .B(n10816), .Z(n10658) );
  NAND U11351 ( .A(n10659), .B(n10658), .Z(n10758) );
  XNOR U11352 ( .A(n10759), .B(n10758), .Z(n10761) );
  NAND U11353 ( .A(n188), .B(n10660), .Z(n10662) );
  XOR U11354 ( .A(b[15]), .B(a[72]), .Z(n10819) );
  NAND U11355 ( .A(n37382), .B(n10819), .Z(n10661) );
  AND U11356 ( .A(n10662), .B(n10661), .Z(n10755) );
  NAND U11357 ( .A(n38064), .B(n10663), .Z(n10665) );
  XOR U11358 ( .A(b[21]), .B(a[66]), .Z(n10822) );
  NAND U11359 ( .A(n37993), .B(n10822), .Z(n10664) );
  AND U11360 ( .A(n10665), .B(n10664), .Z(n10753) );
  NAND U11361 ( .A(n185), .B(n10666), .Z(n10668) );
  XOR U11362 ( .A(b[9]), .B(a[78]), .Z(n10825) );
  NAND U11363 ( .A(n36805), .B(n10825), .Z(n10667) );
  NAND U11364 ( .A(n10668), .B(n10667), .Z(n10752) );
  XNOR U11365 ( .A(n10753), .B(n10752), .Z(n10754) );
  XNOR U11366 ( .A(n10755), .B(n10754), .Z(n10760) );
  XOR U11367 ( .A(n10761), .B(n10760), .Z(n10766) );
  XNOR U11368 ( .A(n10767), .B(n10766), .Z(n10778) );
  XNOR U11369 ( .A(n10779), .B(n10778), .Z(n10710) );
  XNOR U11370 ( .A(n10711), .B(n10710), .Z(n10712) );
  XOR U11371 ( .A(n10713), .B(n10712), .Z(n10829) );
  XOR U11372 ( .A(n10828), .B(n10829), .Z(n10831) );
  XOR U11373 ( .A(n10830), .B(n10831), .Z(n10707) );
  NANDN U11374 ( .A(n10670), .B(n10669), .Z(n10674) );
  NAND U11375 ( .A(n10672), .B(n10671), .Z(n10673) );
  AND U11376 ( .A(n10674), .B(n10673), .Z(n10705) );
  NANDN U11377 ( .A(n10676), .B(n10675), .Z(n10680) );
  NANDN U11378 ( .A(n10678), .B(n10677), .Z(n10679) );
  AND U11379 ( .A(n10680), .B(n10679), .Z(n10704) );
  XNOR U11380 ( .A(n10705), .B(n10704), .Z(n10706) );
  XNOR U11381 ( .A(n10707), .B(n10706), .Z(n10698) );
  NANDN U11382 ( .A(n10682), .B(n10681), .Z(n10686) );
  OR U11383 ( .A(n10684), .B(n10683), .Z(n10685) );
  NAND U11384 ( .A(n10686), .B(n10685), .Z(n10699) );
  XNOR U11385 ( .A(n10698), .B(n10699), .Z(n10700) );
  XNOR U11386 ( .A(n10701), .B(n10700), .Z(n10692) );
  XNOR U11387 ( .A(n10693), .B(n10692), .Z(n10694) );
  XNOR U11388 ( .A(n10695), .B(n10694), .Z(n10834) );
  XNOR U11389 ( .A(sreg[310]), .B(n10834), .Z(n10836) );
  NANDN U11390 ( .A(sreg[309]), .B(n10687), .Z(n10691) );
  NAND U11391 ( .A(n10689), .B(n10688), .Z(n10690) );
  NAND U11392 ( .A(n10691), .B(n10690), .Z(n10835) );
  XNOR U11393 ( .A(n10836), .B(n10835), .Z(c[310]) );
  NANDN U11394 ( .A(n10693), .B(n10692), .Z(n10697) );
  NANDN U11395 ( .A(n10695), .B(n10694), .Z(n10696) );
  AND U11396 ( .A(n10697), .B(n10696), .Z(n10842) );
  NANDN U11397 ( .A(n10699), .B(n10698), .Z(n10703) );
  NANDN U11398 ( .A(n10701), .B(n10700), .Z(n10702) );
  AND U11399 ( .A(n10703), .B(n10702), .Z(n10840) );
  NANDN U11400 ( .A(n10705), .B(n10704), .Z(n10709) );
  NANDN U11401 ( .A(n10707), .B(n10706), .Z(n10708) );
  AND U11402 ( .A(n10709), .B(n10708), .Z(n10848) );
  NANDN U11403 ( .A(n10711), .B(n10710), .Z(n10715) );
  NANDN U11404 ( .A(n10713), .B(n10712), .Z(n10714) );
  AND U11405 ( .A(n10715), .B(n10714), .Z(n10976) );
  NANDN U11406 ( .A(n10717), .B(n10716), .Z(n10721) );
  NAND U11407 ( .A(n10719), .B(n10718), .Z(n10720) );
  AND U11408 ( .A(n10721), .B(n10720), .Z(n10975) );
  XNOR U11409 ( .A(n10976), .B(n10975), .Z(n10978) );
  NANDN U11410 ( .A(n10723), .B(n10722), .Z(n10727) );
  NANDN U11411 ( .A(n10725), .B(n10724), .Z(n10726) );
  AND U11412 ( .A(n10727), .B(n10726), .Z(n10911) );
  NAND U11413 ( .A(n38385), .B(n10728), .Z(n10730) );
  XOR U11414 ( .A(b[27]), .B(a[61]), .Z(n10857) );
  NAND U11415 ( .A(n38343), .B(n10857), .Z(n10729) );
  AND U11416 ( .A(n10730), .B(n10729), .Z(n10918) );
  NAND U11417 ( .A(n183), .B(n10731), .Z(n10733) );
  XOR U11418 ( .A(b[5]), .B(a[83]), .Z(n10860) );
  NAND U11419 ( .A(n36296), .B(n10860), .Z(n10732) );
  AND U11420 ( .A(n10733), .B(n10732), .Z(n10916) );
  NAND U11421 ( .A(n190), .B(n10734), .Z(n10736) );
  XOR U11422 ( .A(b[19]), .B(a[69]), .Z(n10863) );
  NAND U11423 ( .A(n37821), .B(n10863), .Z(n10735) );
  NAND U11424 ( .A(n10736), .B(n10735), .Z(n10915) );
  XNOR U11425 ( .A(n10916), .B(n10915), .Z(n10917) );
  XNOR U11426 ( .A(n10918), .B(n10917), .Z(n10909) );
  NAND U11427 ( .A(n38470), .B(n10737), .Z(n10739) );
  XOR U11428 ( .A(b[31]), .B(a[57]), .Z(n10866) );
  NAND U11429 ( .A(n38453), .B(n10866), .Z(n10738) );
  AND U11430 ( .A(n10739), .B(n10738), .Z(n10878) );
  NAND U11431 ( .A(n181), .B(n10740), .Z(n10742) );
  XOR U11432 ( .A(b[3]), .B(a[85]), .Z(n10869) );
  NAND U11433 ( .A(n182), .B(n10869), .Z(n10741) );
  AND U11434 ( .A(n10742), .B(n10741), .Z(n10876) );
  NAND U11435 ( .A(n189), .B(n10743), .Z(n10745) );
  XOR U11436 ( .A(b[17]), .B(a[71]), .Z(n10872) );
  NAND U11437 ( .A(n37652), .B(n10872), .Z(n10744) );
  NAND U11438 ( .A(n10745), .B(n10744), .Z(n10875) );
  XNOR U11439 ( .A(n10876), .B(n10875), .Z(n10877) );
  XOR U11440 ( .A(n10878), .B(n10877), .Z(n10910) );
  XOR U11441 ( .A(n10909), .B(n10910), .Z(n10912) );
  XOR U11442 ( .A(n10911), .B(n10912), .Z(n10958) );
  NANDN U11443 ( .A(n10747), .B(n10746), .Z(n10751) );
  NANDN U11444 ( .A(n10749), .B(n10748), .Z(n10750) );
  AND U11445 ( .A(n10751), .B(n10750), .Z(n10899) );
  NANDN U11446 ( .A(n10753), .B(n10752), .Z(n10757) );
  NANDN U11447 ( .A(n10755), .B(n10754), .Z(n10756) );
  NAND U11448 ( .A(n10757), .B(n10756), .Z(n10900) );
  XNOR U11449 ( .A(n10899), .B(n10900), .Z(n10901) );
  NANDN U11450 ( .A(n10759), .B(n10758), .Z(n10763) );
  NAND U11451 ( .A(n10761), .B(n10760), .Z(n10762) );
  NAND U11452 ( .A(n10763), .B(n10762), .Z(n10902) );
  XNOR U11453 ( .A(n10901), .B(n10902), .Z(n10957) );
  XNOR U11454 ( .A(n10958), .B(n10957), .Z(n10960) );
  NAND U11455 ( .A(n10765), .B(n10764), .Z(n10769) );
  NAND U11456 ( .A(n10767), .B(n10766), .Z(n10768) );
  AND U11457 ( .A(n10769), .B(n10768), .Z(n10959) );
  XOR U11458 ( .A(n10960), .B(n10959), .Z(n10972) );
  NANDN U11459 ( .A(n10771), .B(n10770), .Z(n10775) );
  NANDN U11460 ( .A(n10773), .B(n10772), .Z(n10774) );
  AND U11461 ( .A(n10775), .B(n10774), .Z(n10969) );
  NANDN U11462 ( .A(n10781), .B(n10780), .Z(n10785) );
  OR U11463 ( .A(n10783), .B(n10782), .Z(n10784) );
  AND U11464 ( .A(n10785), .B(n10784), .Z(n10964) );
  NANDN U11465 ( .A(n10787), .B(n10786), .Z(n10791) );
  NANDN U11466 ( .A(n10789), .B(n10788), .Z(n10790) );
  AND U11467 ( .A(n10791), .B(n10790), .Z(n10906) );
  NANDN U11468 ( .A(n10793), .B(n10792), .Z(n10797) );
  OR U11469 ( .A(n10795), .B(n10794), .Z(n10796) );
  NAND U11470 ( .A(n10797), .B(n10796), .Z(n10905) );
  XNOR U11471 ( .A(n10906), .B(n10905), .Z(n10908) );
  NAND U11472 ( .A(n194), .B(n10798), .Z(n10800) );
  XOR U11473 ( .A(b[29]), .B(a[59]), .Z(n10930) );
  NAND U11474 ( .A(n38456), .B(n10930), .Z(n10799) );
  AND U11475 ( .A(n10800), .B(n10799), .Z(n10852) );
  AND U11476 ( .A(b[31]), .B(a[55]), .Z(n10851) );
  XNOR U11477 ( .A(n10852), .B(n10851), .Z(n10853) );
  NAND U11478 ( .A(b[0]), .B(a[87]), .Z(n10801) );
  XNOR U11479 ( .A(b[1]), .B(n10801), .Z(n10803) );
  NANDN U11480 ( .A(b[0]), .B(a[86]), .Z(n10802) );
  NAND U11481 ( .A(n10803), .B(n10802), .Z(n10854) );
  XNOR U11482 ( .A(n10853), .B(n10854), .Z(n10894) );
  NAND U11483 ( .A(n38185), .B(n10804), .Z(n10806) );
  XOR U11484 ( .A(b[23]), .B(a[65]), .Z(n10933) );
  NAND U11485 ( .A(n38132), .B(n10933), .Z(n10805) );
  AND U11486 ( .A(n10806), .B(n10805), .Z(n10923) );
  NAND U11487 ( .A(n184), .B(n10807), .Z(n10809) );
  XOR U11488 ( .A(b[7]), .B(a[81]), .Z(n10936) );
  NAND U11489 ( .A(n36592), .B(n10936), .Z(n10808) );
  AND U11490 ( .A(n10809), .B(n10808), .Z(n10922) );
  NAND U11491 ( .A(n38289), .B(n10810), .Z(n10812) );
  XOR U11492 ( .A(b[25]), .B(a[63]), .Z(n10939) );
  NAND U11493 ( .A(n38247), .B(n10939), .Z(n10811) );
  NAND U11494 ( .A(n10812), .B(n10811), .Z(n10921) );
  XOR U11495 ( .A(n10922), .B(n10921), .Z(n10924) );
  XOR U11496 ( .A(n10923), .B(n10924), .Z(n10893) );
  XOR U11497 ( .A(n10894), .B(n10893), .Z(n10896) );
  NAND U11498 ( .A(n187), .B(n10813), .Z(n10815) );
  XOR U11499 ( .A(b[13]), .B(a[75]), .Z(n10942) );
  NAND U11500 ( .A(n37295), .B(n10942), .Z(n10814) );
  AND U11501 ( .A(n10815), .B(n10814), .Z(n10888) );
  NAND U11502 ( .A(n186), .B(n10816), .Z(n10818) );
  XOR U11503 ( .A(b[11]), .B(a[77]), .Z(n10945) );
  NAND U11504 ( .A(n37097), .B(n10945), .Z(n10817) );
  NAND U11505 ( .A(n10818), .B(n10817), .Z(n10887) );
  XNOR U11506 ( .A(n10888), .B(n10887), .Z(n10890) );
  NAND U11507 ( .A(n188), .B(n10819), .Z(n10821) );
  XOR U11508 ( .A(b[15]), .B(a[73]), .Z(n10948) );
  NAND U11509 ( .A(n37382), .B(n10948), .Z(n10820) );
  AND U11510 ( .A(n10821), .B(n10820), .Z(n10884) );
  NAND U11511 ( .A(n38064), .B(n10822), .Z(n10824) );
  XOR U11512 ( .A(b[21]), .B(a[67]), .Z(n10951) );
  NAND U11513 ( .A(n37993), .B(n10951), .Z(n10823) );
  AND U11514 ( .A(n10824), .B(n10823), .Z(n10882) );
  NAND U11515 ( .A(n185), .B(n10825), .Z(n10827) );
  XOR U11516 ( .A(b[9]), .B(a[79]), .Z(n10954) );
  NAND U11517 ( .A(n36805), .B(n10954), .Z(n10826) );
  NAND U11518 ( .A(n10827), .B(n10826), .Z(n10881) );
  XNOR U11519 ( .A(n10882), .B(n10881), .Z(n10883) );
  XNOR U11520 ( .A(n10884), .B(n10883), .Z(n10889) );
  XOR U11521 ( .A(n10890), .B(n10889), .Z(n10895) );
  XNOR U11522 ( .A(n10896), .B(n10895), .Z(n10907) );
  XNOR U11523 ( .A(n10908), .B(n10907), .Z(n10963) );
  XNOR U11524 ( .A(n10964), .B(n10963), .Z(n10965) );
  XOR U11525 ( .A(n10966), .B(n10965), .Z(n10970) );
  XNOR U11526 ( .A(n10969), .B(n10970), .Z(n10971) );
  XNOR U11527 ( .A(n10972), .B(n10971), .Z(n10977) );
  XOR U11528 ( .A(n10978), .B(n10977), .Z(n10846) );
  NANDN U11529 ( .A(n10829), .B(n10828), .Z(n10833) );
  OR U11530 ( .A(n10831), .B(n10830), .Z(n10832) );
  AND U11531 ( .A(n10833), .B(n10832), .Z(n10845) );
  XNOR U11532 ( .A(n10846), .B(n10845), .Z(n10847) );
  XNOR U11533 ( .A(n10848), .B(n10847), .Z(n10839) );
  XNOR U11534 ( .A(n10840), .B(n10839), .Z(n10841) );
  XNOR U11535 ( .A(n10842), .B(n10841), .Z(n10981) );
  XNOR U11536 ( .A(sreg[311]), .B(n10981), .Z(n10983) );
  NANDN U11537 ( .A(sreg[310]), .B(n10834), .Z(n10838) );
  NAND U11538 ( .A(n10836), .B(n10835), .Z(n10837) );
  NAND U11539 ( .A(n10838), .B(n10837), .Z(n10982) );
  XNOR U11540 ( .A(n10983), .B(n10982), .Z(c[311]) );
  NANDN U11541 ( .A(n10840), .B(n10839), .Z(n10844) );
  NANDN U11542 ( .A(n10842), .B(n10841), .Z(n10843) );
  AND U11543 ( .A(n10844), .B(n10843), .Z(n10989) );
  NANDN U11544 ( .A(n10846), .B(n10845), .Z(n10850) );
  NANDN U11545 ( .A(n10848), .B(n10847), .Z(n10849) );
  AND U11546 ( .A(n10850), .B(n10849), .Z(n10987) );
  NANDN U11547 ( .A(n10852), .B(n10851), .Z(n10856) );
  NANDN U11548 ( .A(n10854), .B(n10853), .Z(n10855) );
  AND U11549 ( .A(n10856), .B(n10855), .Z(n11066) );
  NAND U11550 ( .A(n38385), .B(n10857), .Z(n10859) );
  XOR U11551 ( .A(b[27]), .B(a[62]), .Z(n11010) );
  NAND U11552 ( .A(n38343), .B(n11010), .Z(n10858) );
  AND U11553 ( .A(n10859), .B(n10858), .Z(n11073) );
  NAND U11554 ( .A(n183), .B(n10860), .Z(n10862) );
  XOR U11555 ( .A(b[5]), .B(a[84]), .Z(n11013) );
  NAND U11556 ( .A(n36296), .B(n11013), .Z(n10861) );
  AND U11557 ( .A(n10862), .B(n10861), .Z(n11071) );
  NAND U11558 ( .A(n190), .B(n10863), .Z(n10865) );
  XOR U11559 ( .A(b[19]), .B(a[70]), .Z(n11016) );
  NAND U11560 ( .A(n37821), .B(n11016), .Z(n10864) );
  NAND U11561 ( .A(n10865), .B(n10864), .Z(n11070) );
  XNOR U11562 ( .A(n11071), .B(n11070), .Z(n11072) );
  XNOR U11563 ( .A(n11073), .B(n11072), .Z(n11064) );
  NAND U11564 ( .A(n38470), .B(n10866), .Z(n10868) );
  XOR U11565 ( .A(b[31]), .B(a[58]), .Z(n11019) );
  NAND U11566 ( .A(n38453), .B(n11019), .Z(n10867) );
  AND U11567 ( .A(n10868), .B(n10867), .Z(n11031) );
  NAND U11568 ( .A(n181), .B(n10869), .Z(n10871) );
  XOR U11569 ( .A(b[3]), .B(a[86]), .Z(n11022) );
  NAND U11570 ( .A(n182), .B(n11022), .Z(n10870) );
  AND U11571 ( .A(n10871), .B(n10870), .Z(n11029) );
  NAND U11572 ( .A(n189), .B(n10872), .Z(n10874) );
  XOR U11573 ( .A(b[17]), .B(a[72]), .Z(n11025) );
  NAND U11574 ( .A(n37652), .B(n11025), .Z(n10873) );
  NAND U11575 ( .A(n10874), .B(n10873), .Z(n11028) );
  XNOR U11576 ( .A(n11029), .B(n11028), .Z(n11030) );
  XOR U11577 ( .A(n11031), .B(n11030), .Z(n11065) );
  XOR U11578 ( .A(n11064), .B(n11065), .Z(n11067) );
  XOR U11579 ( .A(n11066), .B(n11067), .Z(n11113) );
  NANDN U11580 ( .A(n10876), .B(n10875), .Z(n10880) );
  NANDN U11581 ( .A(n10878), .B(n10877), .Z(n10879) );
  AND U11582 ( .A(n10880), .B(n10879), .Z(n11052) );
  NANDN U11583 ( .A(n10882), .B(n10881), .Z(n10886) );
  NANDN U11584 ( .A(n10884), .B(n10883), .Z(n10885) );
  NAND U11585 ( .A(n10886), .B(n10885), .Z(n11053) );
  XNOR U11586 ( .A(n11052), .B(n11053), .Z(n11054) );
  NANDN U11587 ( .A(n10888), .B(n10887), .Z(n10892) );
  NAND U11588 ( .A(n10890), .B(n10889), .Z(n10891) );
  NAND U11589 ( .A(n10892), .B(n10891), .Z(n11055) );
  XNOR U11590 ( .A(n11054), .B(n11055), .Z(n11112) );
  XNOR U11591 ( .A(n11113), .B(n11112), .Z(n11115) );
  NAND U11592 ( .A(n10894), .B(n10893), .Z(n10898) );
  NAND U11593 ( .A(n10896), .B(n10895), .Z(n10897) );
  AND U11594 ( .A(n10898), .B(n10897), .Z(n11114) );
  XOR U11595 ( .A(n11115), .B(n11114), .Z(n11126) );
  NANDN U11596 ( .A(n10900), .B(n10899), .Z(n10904) );
  NANDN U11597 ( .A(n10902), .B(n10901), .Z(n10903) );
  AND U11598 ( .A(n10904), .B(n10903), .Z(n11124) );
  NANDN U11599 ( .A(n10910), .B(n10909), .Z(n10914) );
  OR U11600 ( .A(n10912), .B(n10911), .Z(n10913) );
  AND U11601 ( .A(n10914), .B(n10913), .Z(n11119) );
  NANDN U11602 ( .A(n10916), .B(n10915), .Z(n10920) );
  NANDN U11603 ( .A(n10918), .B(n10917), .Z(n10919) );
  AND U11604 ( .A(n10920), .B(n10919), .Z(n11059) );
  NANDN U11605 ( .A(n10922), .B(n10921), .Z(n10926) );
  OR U11606 ( .A(n10924), .B(n10923), .Z(n10925) );
  NAND U11607 ( .A(n10926), .B(n10925), .Z(n11058) );
  XNOR U11608 ( .A(n11059), .B(n11058), .Z(n11060) );
  NAND U11609 ( .A(b[0]), .B(a[88]), .Z(n10927) );
  XNOR U11610 ( .A(b[1]), .B(n10927), .Z(n10929) );
  NANDN U11611 ( .A(b[0]), .B(a[87]), .Z(n10928) );
  NAND U11612 ( .A(n10929), .B(n10928), .Z(n11007) );
  NAND U11613 ( .A(n194), .B(n10930), .Z(n10932) );
  XOR U11614 ( .A(b[29]), .B(a[60]), .Z(n11085) );
  NAND U11615 ( .A(n38456), .B(n11085), .Z(n10931) );
  AND U11616 ( .A(n10932), .B(n10931), .Z(n11005) );
  AND U11617 ( .A(b[31]), .B(a[56]), .Z(n11004) );
  XNOR U11618 ( .A(n11005), .B(n11004), .Z(n11006) );
  XNOR U11619 ( .A(n11007), .B(n11006), .Z(n11046) );
  NAND U11620 ( .A(n38185), .B(n10933), .Z(n10935) );
  XOR U11621 ( .A(b[23]), .B(a[66]), .Z(n11088) );
  NAND U11622 ( .A(n38132), .B(n11088), .Z(n10934) );
  AND U11623 ( .A(n10935), .B(n10934), .Z(n11079) );
  NAND U11624 ( .A(n184), .B(n10936), .Z(n10938) );
  XOR U11625 ( .A(b[7]), .B(a[82]), .Z(n11091) );
  NAND U11626 ( .A(n36592), .B(n11091), .Z(n10937) );
  AND U11627 ( .A(n10938), .B(n10937), .Z(n11077) );
  NAND U11628 ( .A(n38289), .B(n10939), .Z(n10941) );
  XOR U11629 ( .A(b[25]), .B(a[64]), .Z(n11094) );
  NAND U11630 ( .A(n38247), .B(n11094), .Z(n10940) );
  NAND U11631 ( .A(n10941), .B(n10940), .Z(n11076) );
  XNOR U11632 ( .A(n11077), .B(n11076), .Z(n11078) );
  XOR U11633 ( .A(n11079), .B(n11078), .Z(n11047) );
  XNOR U11634 ( .A(n11046), .B(n11047), .Z(n11048) );
  NAND U11635 ( .A(n187), .B(n10942), .Z(n10944) );
  XOR U11636 ( .A(b[13]), .B(a[76]), .Z(n11097) );
  NAND U11637 ( .A(n37295), .B(n11097), .Z(n10943) );
  AND U11638 ( .A(n10944), .B(n10943), .Z(n11041) );
  NAND U11639 ( .A(n186), .B(n10945), .Z(n10947) );
  XOR U11640 ( .A(b[11]), .B(a[78]), .Z(n11100) );
  NAND U11641 ( .A(n37097), .B(n11100), .Z(n10946) );
  NAND U11642 ( .A(n10947), .B(n10946), .Z(n11040) );
  XNOR U11643 ( .A(n11041), .B(n11040), .Z(n11042) );
  NAND U11644 ( .A(n188), .B(n10948), .Z(n10950) );
  XOR U11645 ( .A(b[15]), .B(a[74]), .Z(n11103) );
  NAND U11646 ( .A(n37382), .B(n11103), .Z(n10949) );
  AND U11647 ( .A(n10950), .B(n10949), .Z(n11037) );
  NAND U11648 ( .A(n38064), .B(n10951), .Z(n10953) );
  XOR U11649 ( .A(b[21]), .B(a[68]), .Z(n11106) );
  NAND U11650 ( .A(n37993), .B(n11106), .Z(n10952) );
  AND U11651 ( .A(n10953), .B(n10952), .Z(n11035) );
  NAND U11652 ( .A(n185), .B(n10954), .Z(n10956) );
  XOR U11653 ( .A(b[9]), .B(a[80]), .Z(n11109) );
  NAND U11654 ( .A(n36805), .B(n11109), .Z(n10955) );
  NAND U11655 ( .A(n10956), .B(n10955), .Z(n11034) );
  XNOR U11656 ( .A(n11035), .B(n11034), .Z(n11036) );
  XOR U11657 ( .A(n11037), .B(n11036), .Z(n11043) );
  XOR U11658 ( .A(n11042), .B(n11043), .Z(n11049) );
  XOR U11659 ( .A(n11048), .B(n11049), .Z(n11061) );
  XNOR U11660 ( .A(n11060), .B(n11061), .Z(n11118) );
  XNOR U11661 ( .A(n11119), .B(n11118), .Z(n11120) );
  XOR U11662 ( .A(n11121), .B(n11120), .Z(n11125) );
  XOR U11663 ( .A(n11124), .B(n11125), .Z(n11127) );
  XOR U11664 ( .A(n11126), .B(n11127), .Z(n11001) );
  NANDN U11665 ( .A(n10958), .B(n10957), .Z(n10962) );
  NAND U11666 ( .A(n10960), .B(n10959), .Z(n10961) );
  AND U11667 ( .A(n10962), .B(n10961), .Z(n10999) );
  NANDN U11668 ( .A(n10964), .B(n10963), .Z(n10968) );
  NANDN U11669 ( .A(n10966), .B(n10965), .Z(n10967) );
  AND U11670 ( .A(n10968), .B(n10967), .Z(n10998) );
  XNOR U11671 ( .A(n10999), .B(n10998), .Z(n11000) );
  XNOR U11672 ( .A(n11001), .B(n11000), .Z(n10992) );
  NANDN U11673 ( .A(n10970), .B(n10969), .Z(n10974) );
  NANDN U11674 ( .A(n10972), .B(n10971), .Z(n10973) );
  NAND U11675 ( .A(n10974), .B(n10973), .Z(n10993) );
  XNOR U11676 ( .A(n10992), .B(n10993), .Z(n10994) );
  NANDN U11677 ( .A(n10976), .B(n10975), .Z(n10980) );
  NAND U11678 ( .A(n10978), .B(n10977), .Z(n10979) );
  NAND U11679 ( .A(n10980), .B(n10979), .Z(n10995) );
  XNOR U11680 ( .A(n10994), .B(n10995), .Z(n10986) );
  XNOR U11681 ( .A(n10987), .B(n10986), .Z(n10988) );
  XNOR U11682 ( .A(n10989), .B(n10988), .Z(n11130) );
  XNOR U11683 ( .A(sreg[312]), .B(n11130), .Z(n11132) );
  NANDN U11684 ( .A(sreg[311]), .B(n10981), .Z(n10985) );
  NAND U11685 ( .A(n10983), .B(n10982), .Z(n10984) );
  NAND U11686 ( .A(n10985), .B(n10984), .Z(n11131) );
  XNOR U11687 ( .A(n11132), .B(n11131), .Z(c[312]) );
  NANDN U11688 ( .A(n10987), .B(n10986), .Z(n10991) );
  NANDN U11689 ( .A(n10989), .B(n10988), .Z(n10990) );
  AND U11690 ( .A(n10991), .B(n10990), .Z(n11138) );
  NANDN U11691 ( .A(n10993), .B(n10992), .Z(n10997) );
  NANDN U11692 ( .A(n10995), .B(n10994), .Z(n10996) );
  AND U11693 ( .A(n10997), .B(n10996), .Z(n11136) );
  NANDN U11694 ( .A(n10999), .B(n10998), .Z(n11003) );
  NANDN U11695 ( .A(n11001), .B(n11000), .Z(n11002) );
  AND U11696 ( .A(n11003), .B(n11002), .Z(n11144) );
  NANDN U11697 ( .A(n11005), .B(n11004), .Z(n11009) );
  NANDN U11698 ( .A(n11007), .B(n11006), .Z(n11008) );
  AND U11699 ( .A(n11009), .B(n11008), .Z(n11227) );
  NAND U11700 ( .A(n38385), .B(n11010), .Z(n11012) );
  XOR U11701 ( .A(b[27]), .B(a[63]), .Z(n11171) );
  NAND U11702 ( .A(n38343), .B(n11171), .Z(n11011) );
  AND U11703 ( .A(n11012), .B(n11011), .Z(n11234) );
  NAND U11704 ( .A(n183), .B(n11013), .Z(n11015) );
  XOR U11705 ( .A(b[5]), .B(a[85]), .Z(n11174) );
  NAND U11706 ( .A(n36296), .B(n11174), .Z(n11014) );
  AND U11707 ( .A(n11015), .B(n11014), .Z(n11232) );
  NAND U11708 ( .A(n190), .B(n11016), .Z(n11018) );
  XOR U11709 ( .A(b[19]), .B(a[71]), .Z(n11177) );
  NAND U11710 ( .A(n37821), .B(n11177), .Z(n11017) );
  NAND U11711 ( .A(n11018), .B(n11017), .Z(n11231) );
  XNOR U11712 ( .A(n11232), .B(n11231), .Z(n11233) );
  XNOR U11713 ( .A(n11234), .B(n11233), .Z(n11225) );
  NAND U11714 ( .A(n38470), .B(n11019), .Z(n11021) );
  XOR U11715 ( .A(b[31]), .B(a[59]), .Z(n11180) );
  NAND U11716 ( .A(n38453), .B(n11180), .Z(n11020) );
  AND U11717 ( .A(n11021), .B(n11020), .Z(n11192) );
  NAND U11718 ( .A(n181), .B(n11022), .Z(n11024) );
  XOR U11719 ( .A(b[3]), .B(a[87]), .Z(n11183) );
  NAND U11720 ( .A(n182), .B(n11183), .Z(n11023) );
  AND U11721 ( .A(n11024), .B(n11023), .Z(n11190) );
  NAND U11722 ( .A(n189), .B(n11025), .Z(n11027) );
  XOR U11723 ( .A(b[17]), .B(a[73]), .Z(n11186) );
  NAND U11724 ( .A(n37652), .B(n11186), .Z(n11026) );
  NAND U11725 ( .A(n11027), .B(n11026), .Z(n11189) );
  XNOR U11726 ( .A(n11190), .B(n11189), .Z(n11191) );
  XOR U11727 ( .A(n11192), .B(n11191), .Z(n11226) );
  XOR U11728 ( .A(n11225), .B(n11226), .Z(n11228) );
  XOR U11729 ( .A(n11227), .B(n11228), .Z(n11160) );
  NANDN U11730 ( .A(n11029), .B(n11028), .Z(n11033) );
  NANDN U11731 ( .A(n11031), .B(n11030), .Z(n11032) );
  AND U11732 ( .A(n11033), .B(n11032), .Z(n11213) );
  NANDN U11733 ( .A(n11035), .B(n11034), .Z(n11039) );
  NANDN U11734 ( .A(n11037), .B(n11036), .Z(n11038) );
  NAND U11735 ( .A(n11039), .B(n11038), .Z(n11214) );
  XNOR U11736 ( .A(n11213), .B(n11214), .Z(n11215) );
  NANDN U11737 ( .A(n11041), .B(n11040), .Z(n11045) );
  NANDN U11738 ( .A(n11043), .B(n11042), .Z(n11044) );
  NAND U11739 ( .A(n11045), .B(n11044), .Z(n11216) );
  XNOR U11740 ( .A(n11215), .B(n11216), .Z(n11159) );
  XNOR U11741 ( .A(n11160), .B(n11159), .Z(n11162) );
  NANDN U11742 ( .A(n11047), .B(n11046), .Z(n11051) );
  NANDN U11743 ( .A(n11049), .B(n11048), .Z(n11050) );
  AND U11744 ( .A(n11051), .B(n11050), .Z(n11161) );
  XOR U11745 ( .A(n11162), .B(n11161), .Z(n11275) );
  NANDN U11746 ( .A(n11053), .B(n11052), .Z(n11057) );
  NANDN U11747 ( .A(n11055), .B(n11054), .Z(n11056) );
  AND U11748 ( .A(n11057), .B(n11056), .Z(n11273) );
  NANDN U11749 ( .A(n11059), .B(n11058), .Z(n11063) );
  NANDN U11750 ( .A(n11061), .B(n11060), .Z(n11062) );
  AND U11751 ( .A(n11063), .B(n11062), .Z(n11156) );
  NANDN U11752 ( .A(n11065), .B(n11064), .Z(n11069) );
  OR U11753 ( .A(n11067), .B(n11066), .Z(n11068) );
  AND U11754 ( .A(n11069), .B(n11068), .Z(n11154) );
  NANDN U11755 ( .A(n11071), .B(n11070), .Z(n11075) );
  NANDN U11756 ( .A(n11073), .B(n11072), .Z(n11074) );
  AND U11757 ( .A(n11075), .B(n11074), .Z(n11220) );
  NANDN U11758 ( .A(n11077), .B(n11076), .Z(n11081) );
  NANDN U11759 ( .A(n11079), .B(n11078), .Z(n11080) );
  NAND U11760 ( .A(n11081), .B(n11080), .Z(n11219) );
  XNOR U11761 ( .A(n11220), .B(n11219), .Z(n11221) );
  NAND U11762 ( .A(b[0]), .B(a[89]), .Z(n11082) );
  XNOR U11763 ( .A(b[1]), .B(n11082), .Z(n11084) );
  NANDN U11764 ( .A(b[0]), .B(a[88]), .Z(n11083) );
  NAND U11765 ( .A(n11084), .B(n11083), .Z(n11168) );
  NAND U11766 ( .A(n194), .B(n11085), .Z(n11087) );
  XOR U11767 ( .A(b[29]), .B(a[61]), .Z(n11246) );
  NAND U11768 ( .A(n38456), .B(n11246), .Z(n11086) );
  AND U11769 ( .A(n11087), .B(n11086), .Z(n11166) );
  AND U11770 ( .A(b[31]), .B(a[57]), .Z(n11165) );
  XNOR U11771 ( .A(n11166), .B(n11165), .Z(n11167) );
  XNOR U11772 ( .A(n11168), .B(n11167), .Z(n11207) );
  NAND U11773 ( .A(n38185), .B(n11088), .Z(n11090) );
  XOR U11774 ( .A(b[23]), .B(a[67]), .Z(n11249) );
  NAND U11775 ( .A(n38132), .B(n11249), .Z(n11089) );
  AND U11776 ( .A(n11090), .B(n11089), .Z(n11240) );
  NAND U11777 ( .A(n184), .B(n11091), .Z(n11093) );
  XOR U11778 ( .A(b[7]), .B(a[83]), .Z(n11252) );
  NAND U11779 ( .A(n36592), .B(n11252), .Z(n11092) );
  AND U11780 ( .A(n11093), .B(n11092), .Z(n11238) );
  NAND U11781 ( .A(n38289), .B(n11094), .Z(n11096) );
  XOR U11782 ( .A(b[25]), .B(a[65]), .Z(n11255) );
  NAND U11783 ( .A(n38247), .B(n11255), .Z(n11095) );
  NAND U11784 ( .A(n11096), .B(n11095), .Z(n11237) );
  XNOR U11785 ( .A(n11238), .B(n11237), .Z(n11239) );
  XOR U11786 ( .A(n11240), .B(n11239), .Z(n11208) );
  XNOR U11787 ( .A(n11207), .B(n11208), .Z(n11209) );
  NAND U11788 ( .A(n187), .B(n11097), .Z(n11099) );
  XOR U11789 ( .A(b[13]), .B(a[77]), .Z(n11258) );
  NAND U11790 ( .A(n37295), .B(n11258), .Z(n11098) );
  AND U11791 ( .A(n11099), .B(n11098), .Z(n11202) );
  NAND U11792 ( .A(n186), .B(n11100), .Z(n11102) );
  XOR U11793 ( .A(b[11]), .B(a[79]), .Z(n11261) );
  NAND U11794 ( .A(n37097), .B(n11261), .Z(n11101) );
  NAND U11795 ( .A(n11102), .B(n11101), .Z(n11201) );
  XNOR U11796 ( .A(n11202), .B(n11201), .Z(n11203) );
  NAND U11797 ( .A(n188), .B(n11103), .Z(n11105) );
  XOR U11798 ( .A(b[15]), .B(a[75]), .Z(n11264) );
  NAND U11799 ( .A(n37382), .B(n11264), .Z(n11104) );
  AND U11800 ( .A(n11105), .B(n11104), .Z(n11198) );
  NAND U11801 ( .A(n38064), .B(n11106), .Z(n11108) );
  XOR U11802 ( .A(b[21]), .B(a[69]), .Z(n11267) );
  NAND U11803 ( .A(n37993), .B(n11267), .Z(n11107) );
  AND U11804 ( .A(n11108), .B(n11107), .Z(n11196) );
  NAND U11805 ( .A(n185), .B(n11109), .Z(n11111) );
  XOR U11806 ( .A(b[9]), .B(a[81]), .Z(n11270) );
  NAND U11807 ( .A(n36805), .B(n11270), .Z(n11110) );
  NAND U11808 ( .A(n11111), .B(n11110), .Z(n11195) );
  XNOR U11809 ( .A(n11196), .B(n11195), .Z(n11197) );
  XOR U11810 ( .A(n11198), .B(n11197), .Z(n11204) );
  XOR U11811 ( .A(n11203), .B(n11204), .Z(n11210) );
  XOR U11812 ( .A(n11209), .B(n11210), .Z(n11222) );
  XNOR U11813 ( .A(n11221), .B(n11222), .Z(n11153) );
  XNOR U11814 ( .A(n11154), .B(n11153), .Z(n11155) );
  XOR U11815 ( .A(n11156), .B(n11155), .Z(n11274) );
  XOR U11816 ( .A(n11273), .B(n11274), .Z(n11276) );
  XOR U11817 ( .A(n11275), .B(n11276), .Z(n11150) );
  NANDN U11818 ( .A(n11113), .B(n11112), .Z(n11117) );
  NAND U11819 ( .A(n11115), .B(n11114), .Z(n11116) );
  AND U11820 ( .A(n11117), .B(n11116), .Z(n11148) );
  NANDN U11821 ( .A(n11119), .B(n11118), .Z(n11123) );
  NANDN U11822 ( .A(n11121), .B(n11120), .Z(n11122) );
  AND U11823 ( .A(n11123), .B(n11122), .Z(n11147) );
  XNOR U11824 ( .A(n11148), .B(n11147), .Z(n11149) );
  XNOR U11825 ( .A(n11150), .B(n11149), .Z(n11141) );
  NANDN U11826 ( .A(n11125), .B(n11124), .Z(n11129) );
  OR U11827 ( .A(n11127), .B(n11126), .Z(n11128) );
  NAND U11828 ( .A(n11129), .B(n11128), .Z(n11142) );
  XNOR U11829 ( .A(n11141), .B(n11142), .Z(n11143) );
  XNOR U11830 ( .A(n11144), .B(n11143), .Z(n11135) );
  XNOR U11831 ( .A(n11136), .B(n11135), .Z(n11137) );
  XNOR U11832 ( .A(n11138), .B(n11137), .Z(n11279) );
  XNOR U11833 ( .A(sreg[313]), .B(n11279), .Z(n11281) );
  NANDN U11834 ( .A(sreg[312]), .B(n11130), .Z(n11134) );
  NAND U11835 ( .A(n11132), .B(n11131), .Z(n11133) );
  NAND U11836 ( .A(n11134), .B(n11133), .Z(n11280) );
  XNOR U11837 ( .A(n11281), .B(n11280), .Z(c[313]) );
  NANDN U11838 ( .A(n11136), .B(n11135), .Z(n11140) );
  NANDN U11839 ( .A(n11138), .B(n11137), .Z(n11139) );
  AND U11840 ( .A(n11140), .B(n11139), .Z(n11287) );
  NANDN U11841 ( .A(n11142), .B(n11141), .Z(n11146) );
  NANDN U11842 ( .A(n11144), .B(n11143), .Z(n11145) );
  AND U11843 ( .A(n11146), .B(n11145), .Z(n11285) );
  NANDN U11844 ( .A(n11148), .B(n11147), .Z(n11152) );
  NANDN U11845 ( .A(n11150), .B(n11149), .Z(n11151) );
  AND U11846 ( .A(n11152), .B(n11151), .Z(n11293) );
  NANDN U11847 ( .A(n11154), .B(n11153), .Z(n11158) );
  NANDN U11848 ( .A(n11156), .B(n11155), .Z(n11157) );
  AND U11849 ( .A(n11158), .B(n11157), .Z(n11297) );
  NANDN U11850 ( .A(n11160), .B(n11159), .Z(n11164) );
  NAND U11851 ( .A(n11162), .B(n11161), .Z(n11163) );
  AND U11852 ( .A(n11164), .B(n11163), .Z(n11296) );
  XNOR U11853 ( .A(n11297), .B(n11296), .Z(n11299) );
  NANDN U11854 ( .A(n11166), .B(n11165), .Z(n11170) );
  NANDN U11855 ( .A(n11168), .B(n11167), .Z(n11169) );
  AND U11856 ( .A(n11170), .B(n11169), .Z(n11374) );
  NAND U11857 ( .A(n38385), .B(n11171), .Z(n11173) );
  XOR U11858 ( .A(b[27]), .B(a[64]), .Z(n11320) );
  NAND U11859 ( .A(n38343), .B(n11320), .Z(n11172) );
  AND U11860 ( .A(n11173), .B(n11172), .Z(n11381) );
  NAND U11861 ( .A(n183), .B(n11174), .Z(n11176) );
  XOR U11862 ( .A(b[5]), .B(a[86]), .Z(n11323) );
  NAND U11863 ( .A(n36296), .B(n11323), .Z(n11175) );
  AND U11864 ( .A(n11176), .B(n11175), .Z(n11379) );
  NAND U11865 ( .A(n190), .B(n11177), .Z(n11179) );
  XOR U11866 ( .A(b[19]), .B(a[72]), .Z(n11326) );
  NAND U11867 ( .A(n37821), .B(n11326), .Z(n11178) );
  NAND U11868 ( .A(n11179), .B(n11178), .Z(n11378) );
  XNOR U11869 ( .A(n11379), .B(n11378), .Z(n11380) );
  XNOR U11870 ( .A(n11381), .B(n11380), .Z(n11372) );
  NAND U11871 ( .A(n38470), .B(n11180), .Z(n11182) );
  XOR U11872 ( .A(b[31]), .B(a[60]), .Z(n11329) );
  NAND U11873 ( .A(n38453), .B(n11329), .Z(n11181) );
  AND U11874 ( .A(n11182), .B(n11181), .Z(n11341) );
  NAND U11875 ( .A(n181), .B(n11183), .Z(n11185) );
  XOR U11876 ( .A(b[3]), .B(a[88]), .Z(n11332) );
  NAND U11877 ( .A(n182), .B(n11332), .Z(n11184) );
  AND U11878 ( .A(n11185), .B(n11184), .Z(n11339) );
  NAND U11879 ( .A(n189), .B(n11186), .Z(n11188) );
  XOR U11880 ( .A(b[17]), .B(a[74]), .Z(n11335) );
  NAND U11881 ( .A(n37652), .B(n11335), .Z(n11187) );
  NAND U11882 ( .A(n11188), .B(n11187), .Z(n11338) );
  XNOR U11883 ( .A(n11339), .B(n11338), .Z(n11340) );
  XOR U11884 ( .A(n11341), .B(n11340), .Z(n11373) );
  XOR U11885 ( .A(n11372), .B(n11373), .Z(n11375) );
  XOR U11886 ( .A(n11374), .B(n11375), .Z(n11309) );
  NANDN U11887 ( .A(n11190), .B(n11189), .Z(n11194) );
  NANDN U11888 ( .A(n11192), .B(n11191), .Z(n11193) );
  AND U11889 ( .A(n11194), .B(n11193), .Z(n11362) );
  NANDN U11890 ( .A(n11196), .B(n11195), .Z(n11200) );
  NANDN U11891 ( .A(n11198), .B(n11197), .Z(n11199) );
  NAND U11892 ( .A(n11200), .B(n11199), .Z(n11363) );
  XNOR U11893 ( .A(n11362), .B(n11363), .Z(n11364) );
  NANDN U11894 ( .A(n11202), .B(n11201), .Z(n11206) );
  NANDN U11895 ( .A(n11204), .B(n11203), .Z(n11205) );
  NAND U11896 ( .A(n11206), .B(n11205), .Z(n11365) );
  XNOR U11897 ( .A(n11364), .B(n11365), .Z(n11308) );
  XNOR U11898 ( .A(n11309), .B(n11308), .Z(n11311) );
  NANDN U11899 ( .A(n11208), .B(n11207), .Z(n11212) );
  NANDN U11900 ( .A(n11210), .B(n11209), .Z(n11211) );
  AND U11901 ( .A(n11212), .B(n11211), .Z(n11310) );
  XOR U11902 ( .A(n11311), .B(n11310), .Z(n11423) );
  NANDN U11903 ( .A(n11214), .B(n11213), .Z(n11218) );
  NANDN U11904 ( .A(n11216), .B(n11215), .Z(n11217) );
  AND U11905 ( .A(n11218), .B(n11217), .Z(n11420) );
  NANDN U11906 ( .A(n11220), .B(n11219), .Z(n11224) );
  NANDN U11907 ( .A(n11222), .B(n11221), .Z(n11223) );
  AND U11908 ( .A(n11224), .B(n11223), .Z(n11305) );
  NANDN U11909 ( .A(n11226), .B(n11225), .Z(n11230) );
  OR U11910 ( .A(n11228), .B(n11227), .Z(n11229) );
  AND U11911 ( .A(n11230), .B(n11229), .Z(n11303) );
  NANDN U11912 ( .A(n11232), .B(n11231), .Z(n11236) );
  NANDN U11913 ( .A(n11234), .B(n11233), .Z(n11235) );
  AND U11914 ( .A(n11236), .B(n11235), .Z(n11369) );
  NANDN U11915 ( .A(n11238), .B(n11237), .Z(n11242) );
  NANDN U11916 ( .A(n11240), .B(n11239), .Z(n11241) );
  NAND U11917 ( .A(n11242), .B(n11241), .Z(n11368) );
  XNOR U11918 ( .A(n11369), .B(n11368), .Z(n11371) );
  NAND U11919 ( .A(b[0]), .B(a[90]), .Z(n11243) );
  XNOR U11920 ( .A(b[1]), .B(n11243), .Z(n11245) );
  NANDN U11921 ( .A(b[0]), .B(a[89]), .Z(n11244) );
  NAND U11922 ( .A(n11245), .B(n11244), .Z(n11317) );
  NAND U11923 ( .A(n194), .B(n11246), .Z(n11248) );
  XOR U11924 ( .A(b[29]), .B(a[62]), .Z(n11390) );
  NAND U11925 ( .A(n38456), .B(n11390), .Z(n11247) );
  AND U11926 ( .A(n11248), .B(n11247), .Z(n11315) );
  AND U11927 ( .A(b[31]), .B(a[58]), .Z(n11314) );
  XNOR U11928 ( .A(n11315), .B(n11314), .Z(n11316) );
  XNOR U11929 ( .A(n11317), .B(n11316), .Z(n11357) );
  NAND U11930 ( .A(n38185), .B(n11249), .Z(n11251) );
  XOR U11931 ( .A(b[23]), .B(a[68]), .Z(n11396) );
  NAND U11932 ( .A(n38132), .B(n11396), .Z(n11250) );
  AND U11933 ( .A(n11251), .B(n11250), .Z(n11386) );
  NAND U11934 ( .A(n184), .B(n11252), .Z(n11254) );
  XOR U11935 ( .A(b[7]), .B(a[84]), .Z(n11399) );
  NAND U11936 ( .A(n36592), .B(n11399), .Z(n11253) );
  AND U11937 ( .A(n11254), .B(n11253), .Z(n11385) );
  NAND U11938 ( .A(n38289), .B(n11255), .Z(n11257) );
  XOR U11939 ( .A(b[25]), .B(a[66]), .Z(n11402) );
  NAND U11940 ( .A(n38247), .B(n11402), .Z(n11256) );
  NAND U11941 ( .A(n11257), .B(n11256), .Z(n11384) );
  XOR U11942 ( .A(n11385), .B(n11384), .Z(n11387) );
  XOR U11943 ( .A(n11386), .B(n11387), .Z(n11356) );
  XOR U11944 ( .A(n11357), .B(n11356), .Z(n11359) );
  NAND U11945 ( .A(n187), .B(n11258), .Z(n11260) );
  XOR U11946 ( .A(b[13]), .B(a[78]), .Z(n11405) );
  NAND U11947 ( .A(n37295), .B(n11405), .Z(n11259) );
  AND U11948 ( .A(n11260), .B(n11259), .Z(n11351) );
  NAND U11949 ( .A(n186), .B(n11261), .Z(n11263) );
  XOR U11950 ( .A(b[11]), .B(a[80]), .Z(n11408) );
  NAND U11951 ( .A(n37097), .B(n11408), .Z(n11262) );
  NAND U11952 ( .A(n11263), .B(n11262), .Z(n11350) );
  XNOR U11953 ( .A(n11351), .B(n11350), .Z(n11353) );
  NAND U11954 ( .A(n188), .B(n11264), .Z(n11266) );
  XOR U11955 ( .A(b[15]), .B(a[76]), .Z(n11411) );
  NAND U11956 ( .A(n37382), .B(n11411), .Z(n11265) );
  AND U11957 ( .A(n11266), .B(n11265), .Z(n11347) );
  NAND U11958 ( .A(n38064), .B(n11267), .Z(n11269) );
  XOR U11959 ( .A(b[21]), .B(a[70]), .Z(n11414) );
  NAND U11960 ( .A(n37993), .B(n11414), .Z(n11268) );
  AND U11961 ( .A(n11269), .B(n11268), .Z(n11345) );
  NAND U11962 ( .A(n185), .B(n11270), .Z(n11272) );
  XOR U11963 ( .A(b[9]), .B(a[82]), .Z(n11417) );
  NAND U11964 ( .A(n36805), .B(n11417), .Z(n11271) );
  NAND U11965 ( .A(n11272), .B(n11271), .Z(n11344) );
  XNOR U11966 ( .A(n11345), .B(n11344), .Z(n11346) );
  XNOR U11967 ( .A(n11347), .B(n11346), .Z(n11352) );
  XOR U11968 ( .A(n11353), .B(n11352), .Z(n11358) );
  XNOR U11969 ( .A(n11359), .B(n11358), .Z(n11370) );
  XNOR U11970 ( .A(n11371), .B(n11370), .Z(n11302) );
  XNOR U11971 ( .A(n11303), .B(n11302), .Z(n11304) );
  XOR U11972 ( .A(n11305), .B(n11304), .Z(n11421) );
  XNOR U11973 ( .A(n11420), .B(n11421), .Z(n11422) );
  XNOR U11974 ( .A(n11423), .B(n11422), .Z(n11298) );
  XOR U11975 ( .A(n11299), .B(n11298), .Z(n11291) );
  NANDN U11976 ( .A(n11274), .B(n11273), .Z(n11278) );
  OR U11977 ( .A(n11276), .B(n11275), .Z(n11277) );
  AND U11978 ( .A(n11278), .B(n11277), .Z(n11290) );
  XNOR U11979 ( .A(n11291), .B(n11290), .Z(n11292) );
  XNOR U11980 ( .A(n11293), .B(n11292), .Z(n11284) );
  XNOR U11981 ( .A(n11285), .B(n11284), .Z(n11286) );
  XNOR U11982 ( .A(n11287), .B(n11286), .Z(n11426) );
  XNOR U11983 ( .A(sreg[314]), .B(n11426), .Z(n11428) );
  NANDN U11984 ( .A(sreg[313]), .B(n11279), .Z(n11283) );
  NAND U11985 ( .A(n11281), .B(n11280), .Z(n11282) );
  NAND U11986 ( .A(n11283), .B(n11282), .Z(n11427) );
  XNOR U11987 ( .A(n11428), .B(n11427), .Z(c[314]) );
  NANDN U11988 ( .A(n11285), .B(n11284), .Z(n11289) );
  NANDN U11989 ( .A(n11287), .B(n11286), .Z(n11288) );
  AND U11990 ( .A(n11289), .B(n11288), .Z(n11434) );
  NANDN U11991 ( .A(n11291), .B(n11290), .Z(n11295) );
  NANDN U11992 ( .A(n11293), .B(n11292), .Z(n11294) );
  AND U11993 ( .A(n11295), .B(n11294), .Z(n11432) );
  NANDN U11994 ( .A(n11297), .B(n11296), .Z(n11301) );
  NAND U11995 ( .A(n11299), .B(n11298), .Z(n11300) );
  AND U11996 ( .A(n11301), .B(n11300), .Z(n11439) );
  NANDN U11997 ( .A(n11303), .B(n11302), .Z(n11307) );
  NANDN U11998 ( .A(n11305), .B(n11304), .Z(n11306) );
  AND U11999 ( .A(n11307), .B(n11306), .Z(n11568) );
  NANDN U12000 ( .A(n11309), .B(n11308), .Z(n11313) );
  NAND U12001 ( .A(n11311), .B(n11310), .Z(n11312) );
  AND U12002 ( .A(n11313), .B(n11312), .Z(n11567) );
  XNOR U12003 ( .A(n11568), .B(n11567), .Z(n11570) );
  NANDN U12004 ( .A(n11315), .B(n11314), .Z(n11319) );
  NANDN U12005 ( .A(n11317), .B(n11316), .Z(n11318) );
  AND U12006 ( .A(n11319), .B(n11318), .Z(n11503) );
  NAND U12007 ( .A(n38385), .B(n11320), .Z(n11322) );
  XOR U12008 ( .A(b[27]), .B(a[65]), .Z(n11449) );
  NAND U12009 ( .A(n38343), .B(n11449), .Z(n11321) );
  AND U12010 ( .A(n11322), .B(n11321), .Z(n11510) );
  NAND U12011 ( .A(n183), .B(n11323), .Z(n11325) );
  XOR U12012 ( .A(b[5]), .B(a[87]), .Z(n11452) );
  NAND U12013 ( .A(n36296), .B(n11452), .Z(n11324) );
  AND U12014 ( .A(n11325), .B(n11324), .Z(n11508) );
  NAND U12015 ( .A(n190), .B(n11326), .Z(n11328) );
  XOR U12016 ( .A(b[19]), .B(a[73]), .Z(n11455) );
  NAND U12017 ( .A(n37821), .B(n11455), .Z(n11327) );
  NAND U12018 ( .A(n11328), .B(n11327), .Z(n11507) );
  XNOR U12019 ( .A(n11508), .B(n11507), .Z(n11509) );
  XNOR U12020 ( .A(n11510), .B(n11509), .Z(n11501) );
  NAND U12021 ( .A(n38470), .B(n11329), .Z(n11331) );
  XOR U12022 ( .A(b[31]), .B(a[61]), .Z(n11458) );
  NAND U12023 ( .A(n38453), .B(n11458), .Z(n11330) );
  AND U12024 ( .A(n11331), .B(n11330), .Z(n11470) );
  NAND U12025 ( .A(n181), .B(n11332), .Z(n11334) );
  XOR U12026 ( .A(b[3]), .B(a[89]), .Z(n11461) );
  NAND U12027 ( .A(n182), .B(n11461), .Z(n11333) );
  AND U12028 ( .A(n11334), .B(n11333), .Z(n11468) );
  NAND U12029 ( .A(n189), .B(n11335), .Z(n11337) );
  XOR U12030 ( .A(b[17]), .B(a[75]), .Z(n11464) );
  NAND U12031 ( .A(n37652), .B(n11464), .Z(n11336) );
  NAND U12032 ( .A(n11337), .B(n11336), .Z(n11467) );
  XNOR U12033 ( .A(n11468), .B(n11467), .Z(n11469) );
  XOR U12034 ( .A(n11470), .B(n11469), .Z(n11502) );
  XOR U12035 ( .A(n11501), .B(n11502), .Z(n11504) );
  XOR U12036 ( .A(n11503), .B(n11504), .Z(n11550) );
  NANDN U12037 ( .A(n11339), .B(n11338), .Z(n11343) );
  NANDN U12038 ( .A(n11341), .B(n11340), .Z(n11342) );
  AND U12039 ( .A(n11343), .B(n11342), .Z(n11491) );
  NANDN U12040 ( .A(n11345), .B(n11344), .Z(n11349) );
  NANDN U12041 ( .A(n11347), .B(n11346), .Z(n11348) );
  NAND U12042 ( .A(n11349), .B(n11348), .Z(n11492) );
  XNOR U12043 ( .A(n11491), .B(n11492), .Z(n11493) );
  NANDN U12044 ( .A(n11351), .B(n11350), .Z(n11355) );
  NAND U12045 ( .A(n11353), .B(n11352), .Z(n11354) );
  NAND U12046 ( .A(n11355), .B(n11354), .Z(n11494) );
  XNOR U12047 ( .A(n11493), .B(n11494), .Z(n11549) );
  XNOR U12048 ( .A(n11550), .B(n11549), .Z(n11552) );
  NAND U12049 ( .A(n11357), .B(n11356), .Z(n11361) );
  NAND U12050 ( .A(n11359), .B(n11358), .Z(n11360) );
  AND U12051 ( .A(n11361), .B(n11360), .Z(n11551) );
  XOR U12052 ( .A(n11552), .B(n11551), .Z(n11564) );
  NANDN U12053 ( .A(n11363), .B(n11362), .Z(n11367) );
  NANDN U12054 ( .A(n11365), .B(n11364), .Z(n11366) );
  AND U12055 ( .A(n11367), .B(n11366), .Z(n11561) );
  NANDN U12056 ( .A(n11373), .B(n11372), .Z(n11377) );
  OR U12057 ( .A(n11375), .B(n11374), .Z(n11376) );
  AND U12058 ( .A(n11377), .B(n11376), .Z(n11556) );
  NANDN U12059 ( .A(n11379), .B(n11378), .Z(n11383) );
  NANDN U12060 ( .A(n11381), .B(n11380), .Z(n11382) );
  AND U12061 ( .A(n11383), .B(n11382), .Z(n11498) );
  NANDN U12062 ( .A(n11385), .B(n11384), .Z(n11389) );
  OR U12063 ( .A(n11387), .B(n11386), .Z(n11388) );
  NAND U12064 ( .A(n11389), .B(n11388), .Z(n11497) );
  XNOR U12065 ( .A(n11498), .B(n11497), .Z(n11500) );
  NAND U12066 ( .A(n194), .B(n11390), .Z(n11392) );
  XOR U12067 ( .A(b[29]), .B(a[63]), .Z(n11522) );
  NAND U12068 ( .A(n38456), .B(n11522), .Z(n11391) );
  AND U12069 ( .A(n11392), .B(n11391), .Z(n11444) );
  AND U12070 ( .A(b[31]), .B(a[59]), .Z(n11443) );
  XNOR U12071 ( .A(n11444), .B(n11443), .Z(n11445) );
  NAND U12072 ( .A(b[0]), .B(a[91]), .Z(n11393) );
  XNOR U12073 ( .A(b[1]), .B(n11393), .Z(n11395) );
  NANDN U12074 ( .A(b[0]), .B(a[90]), .Z(n11394) );
  NAND U12075 ( .A(n11395), .B(n11394), .Z(n11446) );
  XNOR U12076 ( .A(n11445), .B(n11446), .Z(n11486) );
  NAND U12077 ( .A(n38185), .B(n11396), .Z(n11398) );
  XOR U12078 ( .A(b[23]), .B(a[69]), .Z(n11525) );
  NAND U12079 ( .A(n38132), .B(n11525), .Z(n11397) );
  AND U12080 ( .A(n11398), .B(n11397), .Z(n11515) );
  NAND U12081 ( .A(n184), .B(n11399), .Z(n11401) );
  XOR U12082 ( .A(b[7]), .B(a[85]), .Z(n11528) );
  NAND U12083 ( .A(n36592), .B(n11528), .Z(n11400) );
  AND U12084 ( .A(n11401), .B(n11400), .Z(n11514) );
  NAND U12085 ( .A(n38289), .B(n11402), .Z(n11404) );
  XOR U12086 ( .A(b[25]), .B(a[67]), .Z(n11531) );
  NAND U12087 ( .A(n38247), .B(n11531), .Z(n11403) );
  NAND U12088 ( .A(n11404), .B(n11403), .Z(n11513) );
  XOR U12089 ( .A(n11514), .B(n11513), .Z(n11516) );
  XOR U12090 ( .A(n11515), .B(n11516), .Z(n11485) );
  XOR U12091 ( .A(n11486), .B(n11485), .Z(n11488) );
  NAND U12092 ( .A(n187), .B(n11405), .Z(n11407) );
  XOR U12093 ( .A(b[13]), .B(a[79]), .Z(n11534) );
  NAND U12094 ( .A(n37295), .B(n11534), .Z(n11406) );
  AND U12095 ( .A(n11407), .B(n11406), .Z(n11480) );
  NAND U12096 ( .A(n186), .B(n11408), .Z(n11410) );
  XOR U12097 ( .A(b[11]), .B(a[81]), .Z(n11537) );
  NAND U12098 ( .A(n37097), .B(n11537), .Z(n11409) );
  NAND U12099 ( .A(n11410), .B(n11409), .Z(n11479) );
  XNOR U12100 ( .A(n11480), .B(n11479), .Z(n11482) );
  NAND U12101 ( .A(n188), .B(n11411), .Z(n11413) );
  XOR U12102 ( .A(b[15]), .B(a[77]), .Z(n11540) );
  NAND U12103 ( .A(n37382), .B(n11540), .Z(n11412) );
  AND U12104 ( .A(n11413), .B(n11412), .Z(n11476) );
  NAND U12105 ( .A(n38064), .B(n11414), .Z(n11416) );
  XOR U12106 ( .A(b[21]), .B(a[71]), .Z(n11543) );
  NAND U12107 ( .A(n37993), .B(n11543), .Z(n11415) );
  AND U12108 ( .A(n11416), .B(n11415), .Z(n11474) );
  NAND U12109 ( .A(n185), .B(n11417), .Z(n11419) );
  XOR U12110 ( .A(b[9]), .B(a[83]), .Z(n11546) );
  NAND U12111 ( .A(n36805), .B(n11546), .Z(n11418) );
  NAND U12112 ( .A(n11419), .B(n11418), .Z(n11473) );
  XNOR U12113 ( .A(n11474), .B(n11473), .Z(n11475) );
  XNOR U12114 ( .A(n11476), .B(n11475), .Z(n11481) );
  XOR U12115 ( .A(n11482), .B(n11481), .Z(n11487) );
  XNOR U12116 ( .A(n11488), .B(n11487), .Z(n11499) );
  XNOR U12117 ( .A(n11500), .B(n11499), .Z(n11555) );
  XNOR U12118 ( .A(n11556), .B(n11555), .Z(n11557) );
  XOR U12119 ( .A(n11558), .B(n11557), .Z(n11562) );
  XNOR U12120 ( .A(n11561), .B(n11562), .Z(n11563) );
  XNOR U12121 ( .A(n11564), .B(n11563), .Z(n11569) );
  XOR U12122 ( .A(n11570), .B(n11569), .Z(n11438) );
  NANDN U12123 ( .A(n11421), .B(n11420), .Z(n11425) );
  NANDN U12124 ( .A(n11423), .B(n11422), .Z(n11424) );
  AND U12125 ( .A(n11425), .B(n11424), .Z(n11437) );
  XOR U12126 ( .A(n11438), .B(n11437), .Z(n11440) );
  XNOR U12127 ( .A(n11439), .B(n11440), .Z(n11431) );
  XNOR U12128 ( .A(n11432), .B(n11431), .Z(n11433) );
  XNOR U12129 ( .A(n11434), .B(n11433), .Z(n11573) );
  XNOR U12130 ( .A(sreg[315]), .B(n11573), .Z(n11575) );
  NANDN U12131 ( .A(sreg[314]), .B(n11426), .Z(n11430) );
  NAND U12132 ( .A(n11428), .B(n11427), .Z(n11429) );
  NAND U12133 ( .A(n11430), .B(n11429), .Z(n11574) );
  XNOR U12134 ( .A(n11575), .B(n11574), .Z(c[315]) );
  NANDN U12135 ( .A(n11432), .B(n11431), .Z(n11436) );
  NANDN U12136 ( .A(n11434), .B(n11433), .Z(n11435) );
  AND U12137 ( .A(n11436), .B(n11435), .Z(n11581) );
  NANDN U12138 ( .A(n11438), .B(n11437), .Z(n11442) );
  NANDN U12139 ( .A(n11440), .B(n11439), .Z(n11441) );
  AND U12140 ( .A(n11442), .B(n11441), .Z(n11579) );
  NANDN U12141 ( .A(n11444), .B(n11443), .Z(n11448) );
  NANDN U12142 ( .A(n11446), .B(n11445), .Z(n11447) );
  AND U12143 ( .A(n11448), .B(n11447), .Z(n11656) );
  NAND U12144 ( .A(n38385), .B(n11449), .Z(n11451) );
  XOR U12145 ( .A(b[27]), .B(a[66]), .Z(n11602) );
  NAND U12146 ( .A(n38343), .B(n11602), .Z(n11450) );
  AND U12147 ( .A(n11451), .B(n11450), .Z(n11663) );
  NAND U12148 ( .A(n183), .B(n11452), .Z(n11454) );
  XOR U12149 ( .A(b[5]), .B(a[88]), .Z(n11605) );
  NAND U12150 ( .A(n36296), .B(n11605), .Z(n11453) );
  AND U12151 ( .A(n11454), .B(n11453), .Z(n11661) );
  NAND U12152 ( .A(n190), .B(n11455), .Z(n11457) );
  XOR U12153 ( .A(b[19]), .B(a[74]), .Z(n11608) );
  NAND U12154 ( .A(n37821), .B(n11608), .Z(n11456) );
  NAND U12155 ( .A(n11457), .B(n11456), .Z(n11660) );
  XNOR U12156 ( .A(n11661), .B(n11660), .Z(n11662) );
  XNOR U12157 ( .A(n11663), .B(n11662), .Z(n11654) );
  NAND U12158 ( .A(n38470), .B(n11458), .Z(n11460) );
  XOR U12159 ( .A(b[31]), .B(a[62]), .Z(n11611) );
  NAND U12160 ( .A(n38453), .B(n11611), .Z(n11459) );
  AND U12161 ( .A(n11460), .B(n11459), .Z(n11623) );
  NAND U12162 ( .A(n181), .B(n11461), .Z(n11463) );
  XOR U12163 ( .A(b[3]), .B(a[90]), .Z(n11614) );
  NAND U12164 ( .A(n182), .B(n11614), .Z(n11462) );
  AND U12165 ( .A(n11463), .B(n11462), .Z(n11621) );
  NAND U12166 ( .A(n189), .B(n11464), .Z(n11466) );
  XOR U12167 ( .A(b[17]), .B(a[76]), .Z(n11617) );
  NAND U12168 ( .A(n37652), .B(n11617), .Z(n11465) );
  NAND U12169 ( .A(n11466), .B(n11465), .Z(n11620) );
  XNOR U12170 ( .A(n11621), .B(n11620), .Z(n11622) );
  XOR U12171 ( .A(n11623), .B(n11622), .Z(n11655) );
  XOR U12172 ( .A(n11654), .B(n11655), .Z(n11657) );
  XOR U12173 ( .A(n11656), .B(n11657), .Z(n11703) );
  NANDN U12174 ( .A(n11468), .B(n11467), .Z(n11472) );
  NANDN U12175 ( .A(n11470), .B(n11469), .Z(n11471) );
  AND U12176 ( .A(n11472), .B(n11471), .Z(n11644) );
  NANDN U12177 ( .A(n11474), .B(n11473), .Z(n11478) );
  NANDN U12178 ( .A(n11476), .B(n11475), .Z(n11477) );
  NAND U12179 ( .A(n11478), .B(n11477), .Z(n11645) );
  XNOR U12180 ( .A(n11644), .B(n11645), .Z(n11646) );
  NANDN U12181 ( .A(n11480), .B(n11479), .Z(n11484) );
  NAND U12182 ( .A(n11482), .B(n11481), .Z(n11483) );
  NAND U12183 ( .A(n11484), .B(n11483), .Z(n11647) );
  XNOR U12184 ( .A(n11646), .B(n11647), .Z(n11702) );
  XNOR U12185 ( .A(n11703), .B(n11702), .Z(n11705) );
  NAND U12186 ( .A(n11486), .B(n11485), .Z(n11490) );
  NAND U12187 ( .A(n11488), .B(n11487), .Z(n11489) );
  AND U12188 ( .A(n11490), .B(n11489), .Z(n11704) );
  XOR U12189 ( .A(n11705), .B(n11704), .Z(n11716) );
  NANDN U12190 ( .A(n11492), .B(n11491), .Z(n11496) );
  NANDN U12191 ( .A(n11494), .B(n11493), .Z(n11495) );
  AND U12192 ( .A(n11496), .B(n11495), .Z(n11714) );
  NANDN U12193 ( .A(n11502), .B(n11501), .Z(n11506) );
  OR U12194 ( .A(n11504), .B(n11503), .Z(n11505) );
  AND U12195 ( .A(n11506), .B(n11505), .Z(n11709) );
  NANDN U12196 ( .A(n11508), .B(n11507), .Z(n11512) );
  NANDN U12197 ( .A(n11510), .B(n11509), .Z(n11511) );
  AND U12198 ( .A(n11512), .B(n11511), .Z(n11651) );
  NANDN U12199 ( .A(n11514), .B(n11513), .Z(n11518) );
  OR U12200 ( .A(n11516), .B(n11515), .Z(n11517) );
  NAND U12201 ( .A(n11518), .B(n11517), .Z(n11650) );
  XNOR U12202 ( .A(n11651), .B(n11650), .Z(n11653) );
  NAND U12203 ( .A(b[0]), .B(a[92]), .Z(n11519) );
  XNOR U12204 ( .A(b[1]), .B(n11519), .Z(n11521) );
  NANDN U12205 ( .A(b[0]), .B(a[91]), .Z(n11520) );
  NAND U12206 ( .A(n11521), .B(n11520), .Z(n11599) );
  NAND U12207 ( .A(n194), .B(n11522), .Z(n11524) );
  XOR U12208 ( .A(b[29]), .B(a[64]), .Z(n11675) );
  NAND U12209 ( .A(n38456), .B(n11675), .Z(n11523) );
  AND U12210 ( .A(n11524), .B(n11523), .Z(n11597) );
  AND U12211 ( .A(b[31]), .B(a[60]), .Z(n11596) );
  XNOR U12212 ( .A(n11597), .B(n11596), .Z(n11598) );
  XNOR U12213 ( .A(n11599), .B(n11598), .Z(n11639) );
  NAND U12214 ( .A(n38185), .B(n11525), .Z(n11527) );
  XOR U12215 ( .A(b[23]), .B(a[70]), .Z(n11678) );
  NAND U12216 ( .A(n38132), .B(n11678), .Z(n11526) );
  AND U12217 ( .A(n11527), .B(n11526), .Z(n11668) );
  NAND U12218 ( .A(n184), .B(n11528), .Z(n11530) );
  XOR U12219 ( .A(b[7]), .B(a[86]), .Z(n11681) );
  NAND U12220 ( .A(n36592), .B(n11681), .Z(n11529) );
  AND U12221 ( .A(n11530), .B(n11529), .Z(n11667) );
  NAND U12222 ( .A(n38289), .B(n11531), .Z(n11533) );
  XOR U12223 ( .A(b[25]), .B(a[68]), .Z(n11684) );
  NAND U12224 ( .A(n38247), .B(n11684), .Z(n11532) );
  NAND U12225 ( .A(n11533), .B(n11532), .Z(n11666) );
  XOR U12226 ( .A(n11667), .B(n11666), .Z(n11669) );
  XOR U12227 ( .A(n11668), .B(n11669), .Z(n11638) );
  XOR U12228 ( .A(n11639), .B(n11638), .Z(n11641) );
  NAND U12229 ( .A(n187), .B(n11534), .Z(n11536) );
  XOR U12230 ( .A(b[13]), .B(a[80]), .Z(n11687) );
  NAND U12231 ( .A(n37295), .B(n11687), .Z(n11535) );
  AND U12232 ( .A(n11536), .B(n11535), .Z(n11633) );
  NAND U12233 ( .A(n186), .B(n11537), .Z(n11539) );
  XOR U12234 ( .A(b[11]), .B(a[82]), .Z(n11690) );
  NAND U12235 ( .A(n37097), .B(n11690), .Z(n11538) );
  NAND U12236 ( .A(n11539), .B(n11538), .Z(n11632) );
  XNOR U12237 ( .A(n11633), .B(n11632), .Z(n11635) );
  NAND U12238 ( .A(n188), .B(n11540), .Z(n11542) );
  XOR U12239 ( .A(b[15]), .B(a[78]), .Z(n11693) );
  NAND U12240 ( .A(n37382), .B(n11693), .Z(n11541) );
  AND U12241 ( .A(n11542), .B(n11541), .Z(n11629) );
  NAND U12242 ( .A(n38064), .B(n11543), .Z(n11545) );
  XOR U12243 ( .A(b[21]), .B(a[72]), .Z(n11696) );
  NAND U12244 ( .A(n37993), .B(n11696), .Z(n11544) );
  AND U12245 ( .A(n11545), .B(n11544), .Z(n11627) );
  NAND U12246 ( .A(n185), .B(n11546), .Z(n11548) );
  XOR U12247 ( .A(b[9]), .B(a[84]), .Z(n11699) );
  NAND U12248 ( .A(n36805), .B(n11699), .Z(n11547) );
  NAND U12249 ( .A(n11548), .B(n11547), .Z(n11626) );
  XNOR U12250 ( .A(n11627), .B(n11626), .Z(n11628) );
  XNOR U12251 ( .A(n11629), .B(n11628), .Z(n11634) );
  XOR U12252 ( .A(n11635), .B(n11634), .Z(n11640) );
  XNOR U12253 ( .A(n11641), .B(n11640), .Z(n11652) );
  XNOR U12254 ( .A(n11653), .B(n11652), .Z(n11708) );
  XNOR U12255 ( .A(n11709), .B(n11708), .Z(n11710) );
  XOR U12256 ( .A(n11711), .B(n11710), .Z(n11715) );
  XOR U12257 ( .A(n11714), .B(n11715), .Z(n11717) );
  XOR U12258 ( .A(n11716), .B(n11717), .Z(n11593) );
  NANDN U12259 ( .A(n11550), .B(n11549), .Z(n11554) );
  NAND U12260 ( .A(n11552), .B(n11551), .Z(n11553) );
  AND U12261 ( .A(n11554), .B(n11553), .Z(n11591) );
  NANDN U12262 ( .A(n11556), .B(n11555), .Z(n11560) );
  NANDN U12263 ( .A(n11558), .B(n11557), .Z(n11559) );
  AND U12264 ( .A(n11560), .B(n11559), .Z(n11590) );
  XNOR U12265 ( .A(n11591), .B(n11590), .Z(n11592) );
  XNOR U12266 ( .A(n11593), .B(n11592), .Z(n11584) );
  NANDN U12267 ( .A(n11562), .B(n11561), .Z(n11566) );
  NANDN U12268 ( .A(n11564), .B(n11563), .Z(n11565) );
  NAND U12269 ( .A(n11566), .B(n11565), .Z(n11585) );
  XNOR U12270 ( .A(n11584), .B(n11585), .Z(n11586) );
  NANDN U12271 ( .A(n11568), .B(n11567), .Z(n11572) );
  NAND U12272 ( .A(n11570), .B(n11569), .Z(n11571) );
  NAND U12273 ( .A(n11572), .B(n11571), .Z(n11587) );
  XNOR U12274 ( .A(n11586), .B(n11587), .Z(n11578) );
  XNOR U12275 ( .A(n11579), .B(n11578), .Z(n11580) );
  XNOR U12276 ( .A(n11581), .B(n11580), .Z(n11720) );
  XNOR U12277 ( .A(sreg[316]), .B(n11720), .Z(n11722) );
  NANDN U12278 ( .A(sreg[315]), .B(n11573), .Z(n11577) );
  NAND U12279 ( .A(n11575), .B(n11574), .Z(n11576) );
  NAND U12280 ( .A(n11577), .B(n11576), .Z(n11721) );
  XNOR U12281 ( .A(n11722), .B(n11721), .Z(c[316]) );
  NANDN U12282 ( .A(n11579), .B(n11578), .Z(n11583) );
  NANDN U12283 ( .A(n11581), .B(n11580), .Z(n11582) );
  AND U12284 ( .A(n11583), .B(n11582), .Z(n11728) );
  NANDN U12285 ( .A(n11585), .B(n11584), .Z(n11589) );
  NANDN U12286 ( .A(n11587), .B(n11586), .Z(n11588) );
  AND U12287 ( .A(n11589), .B(n11588), .Z(n11726) );
  NANDN U12288 ( .A(n11591), .B(n11590), .Z(n11595) );
  NANDN U12289 ( .A(n11593), .B(n11592), .Z(n11594) );
  AND U12290 ( .A(n11595), .B(n11594), .Z(n11734) );
  NANDN U12291 ( .A(n11597), .B(n11596), .Z(n11601) );
  NANDN U12292 ( .A(n11599), .B(n11598), .Z(n11600) );
  AND U12293 ( .A(n11601), .B(n11600), .Z(n11805) );
  NAND U12294 ( .A(n38385), .B(n11602), .Z(n11604) );
  XOR U12295 ( .A(b[27]), .B(a[67]), .Z(n11749) );
  NAND U12296 ( .A(n38343), .B(n11749), .Z(n11603) );
  AND U12297 ( .A(n11604), .B(n11603), .Z(n11812) );
  NAND U12298 ( .A(n183), .B(n11605), .Z(n11607) );
  XOR U12299 ( .A(b[5]), .B(a[89]), .Z(n11752) );
  NAND U12300 ( .A(n36296), .B(n11752), .Z(n11606) );
  AND U12301 ( .A(n11607), .B(n11606), .Z(n11810) );
  NAND U12302 ( .A(n190), .B(n11608), .Z(n11610) );
  XOR U12303 ( .A(b[19]), .B(a[75]), .Z(n11755) );
  NAND U12304 ( .A(n37821), .B(n11755), .Z(n11609) );
  NAND U12305 ( .A(n11610), .B(n11609), .Z(n11809) );
  XNOR U12306 ( .A(n11810), .B(n11809), .Z(n11811) );
  XNOR U12307 ( .A(n11812), .B(n11811), .Z(n11803) );
  NAND U12308 ( .A(n38470), .B(n11611), .Z(n11613) );
  XOR U12309 ( .A(b[31]), .B(a[63]), .Z(n11758) );
  NAND U12310 ( .A(n38453), .B(n11758), .Z(n11612) );
  AND U12311 ( .A(n11613), .B(n11612), .Z(n11770) );
  NAND U12312 ( .A(n181), .B(n11614), .Z(n11616) );
  XOR U12313 ( .A(b[3]), .B(a[91]), .Z(n11761) );
  NAND U12314 ( .A(n182), .B(n11761), .Z(n11615) );
  AND U12315 ( .A(n11616), .B(n11615), .Z(n11768) );
  NAND U12316 ( .A(n189), .B(n11617), .Z(n11619) );
  XOR U12317 ( .A(b[17]), .B(a[77]), .Z(n11764) );
  NAND U12318 ( .A(n37652), .B(n11764), .Z(n11618) );
  NAND U12319 ( .A(n11619), .B(n11618), .Z(n11767) );
  XNOR U12320 ( .A(n11768), .B(n11767), .Z(n11769) );
  XOR U12321 ( .A(n11770), .B(n11769), .Z(n11804) );
  XOR U12322 ( .A(n11803), .B(n11804), .Z(n11806) );
  XOR U12323 ( .A(n11805), .B(n11806), .Z(n11852) );
  NANDN U12324 ( .A(n11621), .B(n11620), .Z(n11625) );
  NANDN U12325 ( .A(n11623), .B(n11622), .Z(n11624) );
  AND U12326 ( .A(n11625), .B(n11624), .Z(n11791) );
  NANDN U12327 ( .A(n11627), .B(n11626), .Z(n11631) );
  NANDN U12328 ( .A(n11629), .B(n11628), .Z(n11630) );
  NAND U12329 ( .A(n11631), .B(n11630), .Z(n11792) );
  XNOR U12330 ( .A(n11791), .B(n11792), .Z(n11793) );
  NANDN U12331 ( .A(n11633), .B(n11632), .Z(n11637) );
  NAND U12332 ( .A(n11635), .B(n11634), .Z(n11636) );
  NAND U12333 ( .A(n11637), .B(n11636), .Z(n11794) );
  XNOR U12334 ( .A(n11793), .B(n11794), .Z(n11851) );
  XNOR U12335 ( .A(n11852), .B(n11851), .Z(n11854) );
  NAND U12336 ( .A(n11639), .B(n11638), .Z(n11643) );
  NAND U12337 ( .A(n11641), .B(n11640), .Z(n11642) );
  AND U12338 ( .A(n11643), .B(n11642), .Z(n11853) );
  XOR U12339 ( .A(n11854), .B(n11853), .Z(n11865) );
  NANDN U12340 ( .A(n11645), .B(n11644), .Z(n11649) );
  NANDN U12341 ( .A(n11647), .B(n11646), .Z(n11648) );
  AND U12342 ( .A(n11649), .B(n11648), .Z(n11863) );
  NANDN U12343 ( .A(n11655), .B(n11654), .Z(n11659) );
  OR U12344 ( .A(n11657), .B(n11656), .Z(n11658) );
  AND U12345 ( .A(n11659), .B(n11658), .Z(n11858) );
  NANDN U12346 ( .A(n11661), .B(n11660), .Z(n11665) );
  NANDN U12347 ( .A(n11663), .B(n11662), .Z(n11664) );
  AND U12348 ( .A(n11665), .B(n11664), .Z(n11798) );
  NANDN U12349 ( .A(n11667), .B(n11666), .Z(n11671) );
  OR U12350 ( .A(n11669), .B(n11668), .Z(n11670) );
  NAND U12351 ( .A(n11671), .B(n11670), .Z(n11797) );
  XNOR U12352 ( .A(n11798), .B(n11797), .Z(n11799) );
  NAND U12353 ( .A(b[0]), .B(a[93]), .Z(n11672) );
  XNOR U12354 ( .A(b[1]), .B(n11672), .Z(n11674) );
  NANDN U12355 ( .A(b[0]), .B(a[92]), .Z(n11673) );
  NAND U12356 ( .A(n11674), .B(n11673), .Z(n11746) );
  NAND U12357 ( .A(n194), .B(n11675), .Z(n11677) );
  XOR U12358 ( .A(b[29]), .B(a[65]), .Z(n11824) );
  NAND U12359 ( .A(n38456), .B(n11824), .Z(n11676) );
  AND U12360 ( .A(n11677), .B(n11676), .Z(n11744) );
  AND U12361 ( .A(b[31]), .B(a[61]), .Z(n11743) );
  XNOR U12362 ( .A(n11744), .B(n11743), .Z(n11745) );
  XNOR U12363 ( .A(n11746), .B(n11745), .Z(n11785) );
  NAND U12364 ( .A(n38185), .B(n11678), .Z(n11680) );
  XOR U12365 ( .A(b[23]), .B(a[71]), .Z(n11827) );
  NAND U12366 ( .A(n38132), .B(n11827), .Z(n11679) );
  AND U12367 ( .A(n11680), .B(n11679), .Z(n11818) );
  NAND U12368 ( .A(n184), .B(n11681), .Z(n11683) );
  XOR U12369 ( .A(b[7]), .B(a[87]), .Z(n11830) );
  NAND U12370 ( .A(n36592), .B(n11830), .Z(n11682) );
  AND U12371 ( .A(n11683), .B(n11682), .Z(n11816) );
  NAND U12372 ( .A(n38289), .B(n11684), .Z(n11686) );
  XOR U12373 ( .A(b[25]), .B(a[69]), .Z(n11833) );
  NAND U12374 ( .A(n38247), .B(n11833), .Z(n11685) );
  NAND U12375 ( .A(n11686), .B(n11685), .Z(n11815) );
  XNOR U12376 ( .A(n11816), .B(n11815), .Z(n11817) );
  XOR U12377 ( .A(n11818), .B(n11817), .Z(n11786) );
  XNOR U12378 ( .A(n11785), .B(n11786), .Z(n11787) );
  NAND U12379 ( .A(n187), .B(n11687), .Z(n11689) );
  XOR U12380 ( .A(b[13]), .B(a[81]), .Z(n11836) );
  NAND U12381 ( .A(n37295), .B(n11836), .Z(n11688) );
  AND U12382 ( .A(n11689), .B(n11688), .Z(n11780) );
  NAND U12383 ( .A(n186), .B(n11690), .Z(n11692) );
  XOR U12384 ( .A(b[11]), .B(a[83]), .Z(n11839) );
  NAND U12385 ( .A(n37097), .B(n11839), .Z(n11691) );
  NAND U12386 ( .A(n11692), .B(n11691), .Z(n11779) );
  XNOR U12387 ( .A(n11780), .B(n11779), .Z(n11781) );
  NAND U12388 ( .A(n188), .B(n11693), .Z(n11695) );
  XOR U12389 ( .A(b[15]), .B(a[79]), .Z(n11842) );
  NAND U12390 ( .A(n37382), .B(n11842), .Z(n11694) );
  AND U12391 ( .A(n11695), .B(n11694), .Z(n11776) );
  NAND U12392 ( .A(n38064), .B(n11696), .Z(n11698) );
  XOR U12393 ( .A(b[21]), .B(a[73]), .Z(n11845) );
  NAND U12394 ( .A(n37993), .B(n11845), .Z(n11697) );
  AND U12395 ( .A(n11698), .B(n11697), .Z(n11774) );
  NAND U12396 ( .A(n185), .B(n11699), .Z(n11701) );
  XOR U12397 ( .A(b[9]), .B(a[85]), .Z(n11848) );
  NAND U12398 ( .A(n36805), .B(n11848), .Z(n11700) );
  NAND U12399 ( .A(n11701), .B(n11700), .Z(n11773) );
  XNOR U12400 ( .A(n11774), .B(n11773), .Z(n11775) );
  XOR U12401 ( .A(n11776), .B(n11775), .Z(n11782) );
  XOR U12402 ( .A(n11781), .B(n11782), .Z(n11788) );
  XOR U12403 ( .A(n11787), .B(n11788), .Z(n11800) );
  XNOR U12404 ( .A(n11799), .B(n11800), .Z(n11857) );
  XNOR U12405 ( .A(n11858), .B(n11857), .Z(n11859) );
  XOR U12406 ( .A(n11860), .B(n11859), .Z(n11864) );
  XOR U12407 ( .A(n11863), .B(n11864), .Z(n11866) );
  XOR U12408 ( .A(n11865), .B(n11866), .Z(n11740) );
  NANDN U12409 ( .A(n11703), .B(n11702), .Z(n11707) );
  NAND U12410 ( .A(n11705), .B(n11704), .Z(n11706) );
  AND U12411 ( .A(n11707), .B(n11706), .Z(n11738) );
  NANDN U12412 ( .A(n11709), .B(n11708), .Z(n11713) );
  NANDN U12413 ( .A(n11711), .B(n11710), .Z(n11712) );
  AND U12414 ( .A(n11713), .B(n11712), .Z(n11737) );
  XNOR U12415 ( .A(n11738), .B(n11737), .Z(n11739) );
  XNOR U12416 ( .A(n11740), .B(n11739), .Z(n11731) );
  NANDN U12417 ( .A(n11715), .B(n11714), .Z(n11719) );
  OR U12418 ( .A(n11717), .B(n11716), .Z(n11718) );
  NAND U12419 ( .A(n11719), .B(n11718), .Z(n11732) );
  XNOR U12420 ( .A(n11731), .B(n11732), .Z(n11733) );
  XNOR U12421 ( .A(n11734), .B(n11733), .Z(n11725) );
  XNOR U12422 ( .A(n11726), .B(n11725), .Z(n11727) );
  XNOR U12423 ( .A(n11728), .B(n11727), .Z(n11869) );
  XNOR U12424 ( .A(sreg[317]), .B(n11869), .Z(n11871) );
  NANDN U12425 ( .A(sreg[316]), .B(n11720), .Z(n11724) );
  NAND U12426 ( .A(n11722), .B(n11721), .Z(n11723) );
  NAND U12427 ( .A(n11724), .B(n11723), .Z(n11870) );
  XNOR U12428 ( .A(n11871), .B(n11870), .Z(c[317]) );
  NANDN U12429 ( .A(n11726), .B(n11725), .Z(n11730) );
  NANDN U12430 ( .A(n11728), .B(n11727), .Z(n11729) );
  AND U12431 ( .A(n11730), .B(n11729), .Z(n11877) );
  NANDN U12432 ( .A(n11732), .B(n11731), .Z(n11736) );
  NANDN U12433 ( .A(n11734), .B(n11733), .Z(n11735) );
  AND U12434 ( .A(n11736), .B(n11735), .Z(n11875) );
  NANDN U12435 ( .A(n11738), .B(n11737), .Z(n11742) );
  NANDN U12436 ( .A(n11740), .B(n11739), .Z(n11741) );
  AND U12437 ( .A(n11742), .B(n11741), .Z(n11883) );
  NANDN U12438 ( .A(n11744), .B(n11743), .Z(n11748) );
  NANDN U12439 ( .A(n11746), .B(n11745), .Z(n11747) );
  AND U12440 ( .A(n11748), .B(n11747), .Z(n11964) );
  NAND U12441 ( .A(n38385), .B(n11749), .Z(n11751) );
  XOR U12442 ( .A(b[27]), .B(a[68]), .Z(n11910) );
  NAND U12443 ( .A(n38343), .B(n11910), .Z(n11750) );
  AND U12444 ( .A(n11751), .B(n11750), .Z(n11971) );
  NAND U12445 ( .A(n183), .B(n11752), .Z(n11754) );
  XOR U12446 ( .A(b[5]), .B(a[90]), .Z(n11913) );
  NAND U12447 ( .A(n36296), .B(n11913), .Z(n11753) );
  AND U12448 ( .A(n11754), .B(n11753), .Z(n11969) );
  NAND U12449 ( .A(n190), .B(n11755), .Z(n11757) );
  XOR U12450 ( .A(b[19]), .B(a[76]), .Z(n11916) );
  NAND U12451 ( .A(n37821), .B(n11916), .Z(n11756) );
  NAND U12452 ( .A(n11757), .B(n11756), .Z(n11968) );
  XNOR U12453 ( .A(n11969), .B(n11968), .Z(n11970) );
  XNOR U12454 ( .A(n11971), .B(n11970), .Z(n11962) );
  NAND U12455 ( .A(n38470), .B(n11758), .Z(n11760) );
  XOR U12456 ( .A(b[31]), .B(a[64]), .Z(n11919) );
  NAND U12457 ( .A(n38453), .B(n11919), .Z(n11759) );
  AND U12458 ( .A(n11760), .B(n11759), .Z(n11931) );
  NAND U12459 ( .A(n181), .B(n11761), .Z(n11763) );
  XOR U12460 ( .A(b[3]), .B(a[92]), .Z(n11922) );
  NAND U12461 ( .A(n182), .B(n11922), .Z(n11762) );
  AND U12462 ( .A(n11763), .B(n11762), .Z(n11929) );
  NAND U12463 ( .A(n189), .B(n11764), .Z(n11766) );
  XOR U12464 ( .A(b[17]), .B(a[78]), .Z(n11925) );
  NAND U12465 ( .A(n37652), .B(n11925), .Z(n11765) );
  NAND U12466 ( .A(n11766), .B(n11765), .Z(n11928) );
  XNOR U12467 ( .A(n11929), .B(n11928), .Z(n11930) );
  XOR U12468 ( .A(n11931), .B(n11930), .Z(n11963) );
  XOR U12469 ( .A(n11962), .B(n11963), .Z(n11965) );
  XOR U12470 ( .A(n11964), .B(n11965), .Z(n11899) );
  NANDN U12471 ( .A(n11768), .B(n11767), .Z(n11772) );
  NANDN U12472 ( .A(n11770), .B(n11769), .Z(n11771) );
  AND U12473 ( .A(n11772), .B(n11771), .Z(n11952) );
  NANDN U12474 ( .A(n11774), .B(n11773), .Z(n11778) );
  NANDN U12475 ( .A(n11776), .B(n11775), .Z(n11777) );
  NAND U12476 ( .A(n11778), .B(n11777), .Z(n11953) );
  XNOR U12477 ( .A(n11952), .B(n11953), .Z(n11954) );
  NANDN U12478 ( .A(n11780), .B(n11779), .Z(n11784) );
  NANDN U12479 ( .A(n11782), .B(n11781), .Z(n11783) );
  NAND U12480 ( .A(n11784), .B(n11783), .Z(n11955) );
  XNOR U12481 ( .A(n11954), .B(n11955), .Z(n11898) );
  XNOR U12482 ( .A(n11899), .B(n11898), .Z(n11901) );
  NANDN U12483 ( .A(n11786), .B(n11785), .Z(n11790) );
  NANDN U12484 ( .A(n11788), .B(n11787), .Z(n11789) );
  AND U12485 ( .A(n11790), .B(n11789), .Z(n11900) );
  XOR U12486 ( .A(n11901), .B(n11900), .Z(n12012) );
  NANDN U12487 ( .A(n11792), .B(n11791), .Z(n11796) );
  NANDN U12488 ( .A(n11794), .B(n11793), .Z(n11795) );
  AND U12489 ( .A(n11796), .B(n11795), .Z(n12010) );
  NANDN U12490 ( .A(n11798), .B(n11797), .Z(n11802) );
  NANDN U12491 ( .A(n11800), .B(n11799), .Z(n11801) );
  AND U12492 ( .A(n11802), .B(n11801), .Z(n11895) );
  NANDN U12493 ( .A(n11804), .B(n11803), .Z(n11808) );
  OR U12494 ( .A(n11806), .B(n11805), .Z(n11807) );
  AND U12495 ( .A(n11808), .B(n11807), .Z(n11893) );
  NANDN U12496 ( .A(n11810), .B(n11809), .Z(n11814) );
  NANDN U12497 ( .A(n11812), .B(n11811), .Z(n11813) );
  AND U12498 ( .A(n11814), .B(n11813), .Z(n11959) );
  NANDN U12499 ( .A(n11816), .B(n11815), .Z(n11820) );
  NANDN U12500 ( .A(n11818), .B(n11817), .Z(n11819) );
  NAND U12501 ( .A(n11820), .B(n11819), .Z(n11958) );
  XNOR U12502 ( .A(n11959), .B(n11958), .Z(n11961) );
  NAND U12503 ( .A(b[0]), .B(a[94]), .Z(n11821) );
  XNOR U12504 ( .A(b[1]), .B(n11821), .Z(n11823) );
  NANDN U12505 ( .A(b[0]), .B(a[93]), .Z(n11822) );
  NAND U12506 ( .A(n11823), .B(n11822), .Z(n11907) );
  NAND U12507 ( .A(n194), .B(n11824), .Z(n11826) );
  XOR U12508 ( .A(b[29]), .B(a[66]), .Z(n11980) );
  NAND U12509 ( .A(n38456), .B(n11980), .Z(n11825) );
  AND U12510 ( .A(n11826), .B(n11825), .Z(n11905) );
  AND U12511 ( .A(b[31]), .B(a[62]), .Z(n11904) );
  XNOR U12512 ( .A(n11905), .B(n11904), .Z(n11906) );
  XNOR U12513 ( .A(n11907), .B(n11906), .Z(n11947) );
  NAND U12514 ( .A(n38185), .B(n11827), .Z(n11829) );
  XOR U12515 ( .A(b[23]), .B(a[72]), .Z(n11986) );
  NAND U12516 ( .A(n38132), .B(n11986), .Z(n11828) );
  AND U12517 ( .A(n11829), .B(n11828), .Z(n11976) );
  NAND U12518 ( .A(n184), .B(n11830), .Z(n11832) );
  XOR U12519 ( .A(b[7]), .B(a[88]), .Z(n11989) );
  NAND U12520 ( .A(n36592), .B(n11989), .Z(n11831) );
  AND U12521 ( .A(n11832), .B(n11831), .Z(n11975) );
  NAND U12522 ( .A(n38289), .B(n11833), .Z(n11835) );
  XOR U12523 ( .A(b[25]), .B(a[70]), .Z(n11992) );
  NAND U12524 ( .A(n38247), .B(n11992), .Z(n11834) );
  NAND U12525 ( .A(n11835), .B(n11834), .Z(n11974) );
  XOR U12526 ( .A(n11975), .B(n11974), .Z(n11977) );
  XOR U12527 ( .A(n11976), .B(n11977), .Z(n11946) );
  XOR U12528 ( .A(n11947), .B(n11946), .Z(n11949) );
  NAND U12529 ( .A(n187), .B(n11836), .Z(n11838) );
  XOR U12530 ( .A(b[13]), .B(a[82]), .Z(n11995) );
  NAND U12531 ( .A(n37295), .B(n11995), .Z(n11837) );
  AND U12532 ( .A(n11838), .B(n11837), .Z(n11941) );
  NAND U12533 ( .A(n186), .B(n11839), .Z(n11841) );
  XOR U12534 ( .A(b[11]), .B(a[84]), .Z(n11998) );
  NAND U12535 ( .A(n37097), .B(n11998), .Z(n11840) );
  NAND U12536 ( .A(n11841), .B(n11840), .Z(n11940) );
  XNOR U12537 ( .A(n11941), .B(n11940), .Z(n11943) );
  NAND U12538 ( .A(n188), .B(n11842), .Z(n11844) );
  XOR U12539 ( .A(b[15]), .B(a[80]), .Z(n12001) );
  NAND U12540 ( .A(n37382), .B(n12001), .Z(n11843) );
  AND U12541 ( .A(n11844), .B(n11843), .Z(n11937) );
  NAND U12542 ( .A(n38064), .B(n11845), .Z(n11847) );
  XOR U12543 ( .A(b[21]), .B(a[74]), .Z(n12004) );
  NAND U12544 ( .A(n37993), .B(n12004), .Z(n11846) );
  AND U12545 ( .A(n11847), .B(n11846), .Z(n11935) );
  NAND U12546 ( .A(n185), .B(n11848), .Z(n11850) );
  XOR U12547 ( .A(b[9]), .B(a[86]), .Z(n12007) );
  NAND U12548 ( .A(n36805), .B(n12007), .Z(n11849) );
  NAND U12549 ( .A(n11850), .B(n11849), .Z(n11934) );
  XNOR U12550 ( .A(n11935), .B(n11934), .Z(n11936) );
  XNOR U12551 ( .A(n11937), .B(n11936), .Z(n11942) );
  XOR U12552 ( .A(n11943), .B(n11942), .Z(n11948) );
  XNOR U12553 ( .A(n11949), .B(n11948), .Z(n11960) );
  XNOR U12554 ( .A(n11961), .B(n11960), .Z(n11892) );
  XNOR U12555 ( .A(n11893), .B(n11892), .Z(n11894) );
  XOR U12556 ( .A(n11895), .B(n11894), .Z(n12011) );
  XOR U12557 ( .A(n12010), .B(n12011), .Z(n12013) );
  XOR U12558 ( .A(n12012), .B(n12013), .Z(n11889) );
  NANDN U12559 ( .A(n11852), .B(n11851), .Z(n11856) );
  NAND U12560 ( .A(n11854), .B(n11853), .Z(n11855) );
  AND U12561 ( .A(n11856), .B(n11855), .Z(n11887) );
  NANDN U12562 ( .A(n11858), .B(n11857), .Z(n11862) );
  NANDN U12563 ( .A(n11860), .B(n11859), .Z(n11861) );
  AND U12564 ( .A(n11862), .B(n11861), .Z(n11886) );
  XNOR U12565 ( .A(n11887), .B(n11886), .Z(n11888) );
  XNOR U12566 ( .A(n11889), .B(n11888), .Z(n11880) );
  NANDN U12567 ( .A(n11864), .B(n11863), .Z(n11868) );
  OR U12568 ( .A(n11866), .B(n11865), .Z(n11867) );
  NAND U12569 ( .A(n11868), .B(n11867), .Z(n11881) );
  XNOR U12570 ( .A(n11880), .B(n11881), .Z(n11882) );
  XNOR U12571 ( .A(n11883), .B(n11882), .Z(n11874) );
  XNOR U12572 ( .A(n11875), .B(n11874), .Z(n11876) );
  XNOR U12573 ( .A(n11877), .B(n11876), .Z(n12016) );
  XNOR U12574 ( .A(sreg[318]), .B(n12016), .Z(n12018) );
  NANDN U12575 ( .A(sreg[317]), .B(n11869), .Z(n11873) );
  NAND U12576 ( .A(n11871), .B(n11870), .Z(n11872) );
  NAND U12577 ( .A(n11873), .B(n11872), .Z(n12017) );
  XNOR U12578 ( .A(n12018), .B(n12017), .Z(c[318]) );
  NANDN U12579 ( .A(n11875), .B(n11874), .Z(n11879) );
  NANDN U12580 ( .A(n11877), .B(n11876), .Z(n11878) );
  AND U12581 ( .A(n11879), .B(n11878), .Z(n12024) );
  NANDN U12582 ( .A(n11881), .B(n11880), .Z(n11885) );
  NANDN U12583 ( .A(n11883), .B(n11882), .Z(n11884) );
  AND U12584 ( .A(n11885), .B(n11884), .Z(n12022) );
  NANDN U12585 ( .A(n11887), .B(n11886), .Z(n11891) );
  NANDN U12586 ( .A(n11889), .B(n11888), .Z(n11890) );
  AND U12587 ( .A(n11891), .B(n11890), .Z(n12030) );
  NANDN U12588 ( .A(n11893), .B(n11892), .Z(n11897) );
  NANDN U12589 ( .A(n11895), .B(n11894), .Z(n11896) );
  AND U12590 ( .A(n11897), .B(n11896), .Z(n12160) );
  NANDN U12591 ( .A(n11899), .B(n11898), .Z(n11903) );
  NAND U12592 ( .A(n11901), .B(n11900), .Z(n11902) );
  AND U12593 ( .A(n11903), .B(n11902), .Z(n12159) );
  XNOR U12594 ( .A(n12160), .B(n12159), .Z(n12162) );
  NANDN U12595 ( .A(n11905), .B(n11904), .Z(n11909) );
  NANDN U12596 ( .A(n11907), .B(n11906), .Z(n11908) );
  AND U12597 ( .A(n11909), .B(n11908), .Z(n12095) );
  NAND U12598 ( .A(n38385), .B(n11910), .Z(n11912) );
  XOR U12599 ( .A(b[27]), .B(a[69]), .Z(n12039) );
  NAND U12600 ( .A(n38343), .B(n12039), .Z(n11911) );
  AND U12601 ( .A(n11912), .B(n11911), .Z(n12102) );
  NAND U12602 ( .A(n183), .B(n11913), .Z(n11915) );
  XOR U12603 ( .A(b[5]), .B(a[91]), .Z(n12042) );
  NAND U12604 ( .A(n36296), .B(n12042), .Z(n11914) );
  AND U12605 ( .A(n11915), .B(n11914), .Z(n12100) );
  NAND U12606 ( .A(n190), .B(n11916), .Z(n11918) );
  XOR U12607 ( .A(b[19]), .B(a[77]), .Z(n12045) );
  NAND U12608 ( .A(n37821), .B(n12045), .Z(n11917) );
  NAND U12609 ( .A(n11918), .B(n11917), .Z(n12099) );
  XNOR U12610 ( .A(n12100), .B(n12099), .Z(n12101) );
  XNOR U12611 ( .A(n12102), .B(n12101), .Z(n12093) );
  NAND U12612 ( .A(n38470), .B(n11919), .Z(n11921) );
  XOR U12613 ( .A(b[31]), .B(a[65]), .Z(n12048) );
  NAND U12614 ( .A(n38453), .B(n12048), .Z(n11920) );
  AND U12615 ( .A(n11921), .B(n11920), .Z(n12060) );
  NAND U12616 ( .A(n181), .B(n11922), .Z(n11924) );
  XOR U12617 ( .A(b[3]), .B(a[93]), .Z(n12051) );
  NAND U12618 ( .A(n182), .B(n12051), .Z(n11923) );
  AND U12619 ( .A(n11924), .B(n11923), .Z(n12058) );
  NAND U12620 ( .A(n189), .B(n11925), .Z(n11927) );
  XOR U12621 ( .A(b[17]), .B(a[79]), .Z(n12054) );
  NAND U12622 ( .A(n37652), .B(n12054), .Z(n11926) );
  NAND U12623 ( .A(n11927), .B(n11926), .Z(n12057) );
  XNOR U12624 ( .A(n12058), .B(n12057), .Z(n12059) );
  XOR U12625 ( .A(n12060), .B(n12059), .Z(n12094) );
  XOR U12626 ( .A(n12093), .B(n12094), .Z(n12096) );
  XOR U12627 ( .A(n12095), .B(n12096), .Z(n12142) );
  NANDN U12628 ( .A(n11929), .B(n11928), .Z(n11933) );
  NANDN U12629 ( .A(n11931), .B(n11930), .Z(n11932) );
  AND U12630 ( .A(n11933), .B(n11932), .Z(n12081) );
  NANDN U12631 ( .A(n11935), .B(n11934), .Z(n11939) );
  NANDN U12632 ( .A(n11937), .B(n11936), .Z(n11938) );
  NAND U12633 ( .A(n11939), .B(n11938), .Z(n12082) );
  XNOR U12634 ( .A(n12081), .B(n12082), .Z(n12083) );
  NANDN U12635 ( .A(n11941), .B(n11940), .Z(n11945) );
  NAND U12636 ( .A(n11943), .B(n11942), .Z(n11944) );
  NAND U12637 ( .A(n11945), .B(n11944), .Z(n12084) );
  XNOR U12638 ( .A(n12083), .B(n12084), .Z(n12141) );
  XNOR U12639 ( .A(n12142), .B(n12141), .Z(n12144) );
  NAND U12640 ( .A(n11947), .B(n11946), .Z(n11951) );
  NAND U12641 ( .A(n11949), .B(n11948), .Z(n11950) );
  AND U12642 ( .A(n11951), .B(n11950), .Z(n12143) );
  XOR U12643 ( .A(n12144), .B(n12143), .Z(n12156) );
  NANDN U12644 ( .A(n11953), .B(n11952), .Z(n11957) );
  NANDN U12645 ( .A(n11955), .B(n11954), .Z(n11956) );
  AND U12646 ( .A(n11957), .B(n11956), .Z(n12153) );
  NANDN U12647 ( .A(n11963), .B(n11962), .Z(n11967) );
  OR U12648 ( .A(n11965), .B(n11964), .Z(n11966) );
  AND U12649 ( .A(n11967), .B(n11966), .Z(n12148) );
  NANDN U12650 ( .A(n11969), .B(n11968), .Z(n11973) );
  NANDN U12651 ( .A(n11971), .B(n11970), .Z(n11972) );
  AND U12652 ( .A(n11973), .B(n11972), .Z(n12088) );
  NANDN U12653 ( .A(n11975), .B(n11974), .Z(n11979) );
  OR U12654 ( .A(n11977), .B(n11976), .Z(n11978) );
  NAND U12655 ( .A(n11979), .B(n11978), .Z(n12087) );
  XNOR U12656 ( .A(n12088), .B(n12087), .Z(n12089) );
  NAND U12657 ( .A(n194), .B(n11980), .Z(n11982) );
  XOR U12658 ( .A(b[29]), .B(a[67]), .Z(n12114) );
  NAND U12659 ( .A(n38456), .B(n12114), .Z(n11981) );
  AND U12660 ( .A(n11982), .B(n11981), .Z(n12034) );
  AND U12661 ( .A(b[31]), .B(a[63]), .Z(n12033) );
  XNOR U12662 ( .A(n12034), .B(n12033), .Z(n12035) );
  NAND U12663 ( .A(b[0]), .B(a[95]), .Z(n11983) );
  XNOR U12664 ( .A(b[1]), .B(n11983), .Z(n11985) );
  NANDN U12665 ( .A(b[0]), .B(a[94]), .Z(n11984) );
  NAND U12666 ( .A(n11985), .B(n11984), .Z(n12036) );
  XNOR U12667 ( .A(n12035), .B(n12036), .Z(n12075) );
  NAND U12668 ( .A(n38185), .B(n11986), .Z(n11988) );
  XOR U12669 ( .A(b[23]), .B(a[73]), .Z(n12117) );
  NAND U12670 ( .A(n38132), .B(n12117), .Z(n11987) );
  AND U12671 ( .A(n11988), .B(n11987), .Z(n12108) );
  NAND U12672 ( .A(n184), .B(n11989), .Z(n11991) );
  XOR U12673 ( .A(b[7]), .B(a[89]), .Z(n12120) );
  NAND U12674 ( .A(n36592), .B(n12120), .Z(n11990) );
  AND U12675 ( .A(n11991), .B(n11990), .Z(n12106) );
  NAND U12676 ( .A(n38289), .B(n11992), .Z(n11994) );
  XOR U12677 ( .A(b[25]), .B(a[71]), .Z(n12123) );
  NAND U12678 ( .A(n38247), .B(n12123), .Z(n11993) );
  NAND U12679 ( .A(n11994), .B(n11993), .Z(n12105) );
  XNOR U12680 ( .A(n12106), .B(n12105), .Z(n12107) );
  XOR U12681 ( .A(n12108), .B(n12107), .Z(n12076) );
  XNOR U12682 ( .A(n12075), .B(n12076), .Z(n12077) );
  NAND U12683 ( .A(n187), .B(n11995), .Z(n11997) );
  XOR U12684 ( .A(b[13]), .B(a[83]), .Z(n12126) );
  NAND U12685 ( .A(n37295), .B(n12126), .Z(n11996) );
  AND U12686 ( .A(n11997), .B(n11996), .Z(n12070) );
  NAND U12687 ( .A(n186), .B(n11998), .Z(n12000) );
  XOR U12688 ( .A(b[11]), .B(a[85]), .Z(n12129) );
  NAND U12689 ( .A(n37097), .B(n12129), .Z(n11999) );
  NAND U12690 ( .A(n12000), .B(n11999), .Z(n12069) );
  XNOR U12691 ( .A(n12070), .B(n12069), .Z(n12071) );
  NAND U12692 ( .A(n188), .B(n12001), .Z(n12003) );
  XOR U12693 ( .A(b[15]), .B(a[81]), .Z(n12132) );
  NAND U12694 ( .A(n37382), .B(n12132), .Z(n12002) );
  AND U12695 ( .A(n12003), .B(n12002), .Z(n12066) );
  NAND U12696 ( .A(n38064), .B(n12004), .Z(n12006) );
  XOR U12697 ( .A(b[21]), .B(a[75]), .Z(n12135) );
  NAND U12698 ( .A(n37993), .B(n12135), .Z(n12005) );
  AND U12699 ( .A(n12006), .B(n12005), .Z(n12064) );
  NAND U12700 ( .A(n185), .B(n12007), .Z(n12009) );
  XOR U12701 ( .A(b[9]), .B(a[87]), .Z(n12138) );
  NAND U12702 ( .A(n36805), .B(n12138), .Z(n12008) );
  NAND U12703 ( .A(n12009), .B(n12008), .Z(n12063) );
  XNOR U12704 ( .A(n12064), .B(n12063), .Z(n12065) );
  XOR U12705 ( .A(n12066), .B(n12065), .Z(n12072) );
  XOR U12706 ( .A(n12071), .B(n12072), .Z(n12078) );
  XOR U12707 ( .A(n12077), .B(n12078), .Z(n12090) );
  XNOR U12708 ( .A(n12089), .B(n12090), .Z(n12147) );
  XNOR U12709 ( .A(n12148), .B(n12147), .Z(n12149) );
  XOR U12710 ( .A(n12150), .B(n12149), .Z(n12154) );
  XNOR U12711 ( .A(n12153), .B(n12154), .Z(n12155) );
  XNOR U12712 ( .A(n12156), .B(n12155), .Z(n12161) );
  XOR U12713 ( .A(n12162), .B(n12161), .Z(n12028) );
  NANDN U12714 ( .A(n12011), .B(n12010), .Z(n12015) );
  OR U12715 ( .A(n12013), .B(n12012), .Z(n12014) );
  AND U12716 ( .A(n12015), .B(n12014), .Z(n12027) );
  XNOR U12717 ( .A(n12028), .B(n12027), .Z(n12029) );
  XNOR U12718 ( .A(n12030), .B(n12029), .Z(n12021) );
  XNOR U12719 ( .A(n12022), .B(n12021), .Z(n12023) );
  XNOR U12720 ( .A(n12024), .B(n12023), .Z(n12165) );
  XNOR U12721 ( .A(sreg[319]), .B(n12165), .Z(n12167) );
  NANDN U12722 ( .A(sreg[318]), .B(n12016), .Z(n12020) );
  NAND U12723 ( .A(n12018), .B(n12017), .Z(n12019) );
  NAND U12724 ( .A(n12020), .B(n12019), .Z(n12166) );
  XNOR U12725 ( .A(n12167), .B(n12166), .Z(c[319]) );
  NANDN U12726 ( .A(n12022), .B(n12021), .Z(n12026) );
  NANDN U12727 ( .A(n12024), .B(n12023), .Z(n12025) );
  AND U12728 ( .A(n12026), .B(n12025), .Z(n12173) );
  NANDN U12729 ( .A(n12028), .B(n12027), .Z(n12032) );
  NANDN U12730 ( .A(n12030), .B(n12029), .Z(n12031) );
  AND U12731 ( .A(n12032), .B(n12031), .Z(n12171) );
  NANDN U12732 ( .A(n12034), .B(n12033), .Z(n12038) );
  NANDN U12733 ( .A(n12036), .B(n12035), .Z(n12037) );
  AND U12734 ( .A(n12038), .B(n12037), .Z(n12262) );
  NAND U12735 ( .A(n38385), .B(n12039), .Z(n12041) );
  XOR U12736 ( .A(b[27]), .B(a[70]), .Z(n12206) );
  NAND U12737 ( .A(n38343), .B(n12206), .Z(n12040) );
  AND U12738 ( .A(n12041), .B(n12040), .Z(n12269) );
  NAND U12739 ( .A(n183), .B(n12042), .Z(n12044) );
  XOR U12740 ( .A(b[5]), .B(a[92]), .Z(n12209) );
  NAND U12741 ( .A(n36296), .B(n12209), .Z(n12043) );
  AND U12742 ( .A(n12044), .B(n12043), .Z(n12267) );
  NAND U12743 ( .A(n190), .B(n12045), .Z(n12047) );
  XOR U12744 ( .A(b[19]), .B(a[78]), .Z(n12212) );
  NAND U12745 ( .A(n37821), .B(n12212), .Z(n12046) );
  NAND U12746 ( .A(n12047), .B(n12046), .Z(n12266) );
  XNOR U12747 ( .A(n12267), .B(n12266), .Z(n12268) );
  XNOR U12748 ( .A(n12269), .B(n12268), .Z(n12260) );
  NAND U12749 ( .A(n38470), .B(n12048), .Z(n12050) );
  XOR U12750 ( .A(b[31]), .B(a[66]), .Z(n12215) );
  NAND U12751 ( .A(n38453), .B(n12215), .Z(n12049) );
  AND U12752 ( .A(n12050), .B(n12049), .Z(n12227) );
  NAND U12753 ( .A(n181), .B(n12051), .Z(n12053) );
  XOR U12754 ( .A(b[3]), .B(a[94]), .Z(n12218) );
  NAND U12755 ( .A(n182), .B(n12218), .Z(n12052) );
  AND U12756 ( .A(n12053), .B(n12052), .Z(n12225) );
  NAND U12757 ( .A(n189), .B(n12054), .Z(n12056) );
  XOR U12758 ( .A(b[17]), .B(a[80]), .Z(n12221) );
  NAND U12759 ( .A(n37652), .B(n12221), .Z(n12055) );
  NAND U12760 ( .A(n12056), .B(n12055), .Z(n12224) );
  XNOR U12761 ( .A(n12225), .B(n12224), .Z(n12226) );
  XOR U12762 ( .A(n12227), .B(n12226), .Z(n12261) );
  XOR U12763 ( .A(n12260), .B(n12261), .Z(n12263) );
  XOR U12764 ( .A(n12262), .B(n12263), .Z(n12195) );
  NANDN U12765 ( .A(n12058), .B(n12057), .Z(n12062) );
  NANDN U12766 ( .A(n12060), .B(n12059), .Z(n12061) );
  AND U12767 ( .A(n12062), .B(n12061), .Z(n12248) );
  NANDN U12768 ( .A(n12064), .B(n12063), .Z(n12068) );
  NANDN U12769 ( .A(n12066), .B(n12065), .Z(n12067) );
  NAND U12770 ( .A(n12068), .B(n12067), .Z(n12249) );
  XNOR U12771 ( .A(n12248), .B(n12249), .Z(n12250) );
  NANDN U12772 ( .A(n12070), .B(n12069), .Z(n12074) );
  NANDN U12773 ( .A(n12072), .B(n12071), .Z(n12073) );
  NAND U12774 ( .A(n12074), .B(n12073), .Z(n12251) );
  XNOR U12775 ( .A(n12250), .B(n12251), .Z(n12194) );
  XNOR U12776 ( .A(n12195), .B(n12194), .Z(n12197) );
  NANDN U12777 ( .A(n12076), .B(n12075), .Z(n12080) );
  NANDN U12778 ( .A(n12078), .B(n12077), .Z(n12079) );
  AND U12779 ( .A(n12080), .B(n12079), .Z(n12196) );
  XOR U12780 ( .A(n12197), .B(n12196), .Z(n12310) );
  NANDN U12781 ( .A(n12082), .B(n12081), .Z(n12086) );
  NANDN U12782 ( .A(n12084), .B(n12083), .Z(n12085) );
  AND U12783 ( .A(n12086), .B(n12085), .Z(n12308) );
  NANDN U12784 ( .A(n12088), .B(n12087), .Z(n12092) );
  NANDN U12785 ( .A(n12090), .B(n12089), .Z(n12091) );
  AND U12786 ( .A(n12092), .B(n12091), .Z(n12191) );
  NANDN U12787 ( .A(n12094), .B(n12093), .Z(n12098) );
  OR U12788 ( .A(n12096), .B(n12095), .Z(n12097) );
  AND U12789 ( .A(n12098), .B(n12097), .Z(n12189) );
  NANDN U12790 ( .A(n12100), .B(n12099), .Z(n12104) );
  NANDN U12791 ( .A(n12102), .B(n12101), .Z(n12103) );
  AND U12792 ( .A(n12104), .B(n12103), .Z(n12255) );
  NANDN U12793 ( .A(n12106), .B(n12105), .Z(n12110) );
  NANDN U12794 ( .A(n12108), .B(n12107), .Z(n12109) );
  NAND U12795 ( .A(n12110), .B(n12109), .Z(n12254) );
  XNOR U12796 ( .A(n12255), .B(n12254), .Z(n12256) );
  NAND U12797 ( .A(b[0]), .B(a[96]), .Z(n12111) );
  XNOR U12798 ( .A(b[1]), .B(n12111), .Z(n12113) );
  NANDN U12799 ( .A(b[0]), .B(a[95]), .Z(n12112) );
  NAND U12800 ( .A(n12113), .B(n12112), .Z(n12203) );
  NAND U12801 ( .A(n194), .B(n12114), .Z(n12116) );
  XOR U12802 ( .A(b[29]), .B(a[68]), .Z(n12281) );
  NAND U12803 ( .A(n38456), .B(n12281), .Z(n12115) );
  AND U12804 ( .A(n12116), .B(n12115), .Z(n12201) );
  AND U12805 ( .A(b[31]), .B(a[64]), .Z(n12200) );
  XNOR U12806 ( .A(n12201), .B(n12200), .Z(n12202) );
  XNOR U12807 ( .A(n12203), .B(n12202), .Z(n12242) );
  NAND U12808 ( .A(n38185), .B(n12117), .Z(n12119) );
  XOR U12809 ( .A(b[23]), .B(a[74]), .Z(n12284) );
  NAND U12810 ( .A(n38132), .B(n12284), .Z(n12118) );
  AND U12811 ( .A(n12119), .B(n12118), .Z(n12275) );
  NAND U12812 ( .A(n184), .B(n12120), .Z(n12122) );
  XOR U12813 ( .A(b[7]), .B(a[90]), .Z(n12287) );
  NAND U12814 ( .A(n36592), .B(n12287), .Z(n12121) );
  AND U12815 ( .A(n12122), .B(n12121), .Z(n12273) );
  NAND U12816 ( .A(n38289), .B(n12123), .Z(n12125) );
  XOR U12817 ( .A(b[25]), .B(a[72]), .Z(n12290) );
  NAND U12818 ( .A(n38247), .B(n12290), .Z(n12124) );
  NAND U12819 ( .A(n12125), .B(n12124), .Z(n12272) );
  XNOR U12820 ( .A(n12273), .B(n12272), .Z(n12274) );
  XOR U12821 ( .A(n12275), .B(n12274), .Z(n12243) );
  XNOR U12822 ( .A(n12242), .B(n12243), .Z(n12244) );
  NAND U12823 ( .A(n187), .B(n12126), .Z(n12128) );
  XOR U12824 ( .A(b[13]), .B(a[84]), .Z(n12293) );
  NAND U12825 ( .A(n37295), .B(n12293), .Z(n12127) );
  AND U12826 ( .A(n12128), .B(n12127), .Z(n12237) );
  NAND U12827 ( .A(n186), .B(n12129), .Z(n12131) );
  XOR U12828 ( .A(b[11]), .B(a[86]), .Z(n12296) );
  NAND U12829 ( .A(n37097), .B(n12296), .Z(n12130) );
  NAND U12830 ( .A(n12131), .B(n12130), .Z(n12236) );
  XNOR U12831 ( .A(n12237), .B(n12236), .Z(n12238) );
  NAND U12832 ( .A(n188), .B(n12132), .Z(n12134) );
  XOR U12833 ( .A(b[15]), .B(a[82]), .Z(n12299) );
  NAND U12834 ( .A(n37382), .B(n12299), .Z(n12133) );
  AND U12835 ( .A(n12134), .B(n12133), .Z(n12233) );
  NAND U12836 ( .A(n38064), .B(n12135), .Z(n12137) );
  XOR U12837 ( .A(b[21]), .B(a[76]), .Z(n12302) );
  NAND U12838 ( .A(n37993), .B(n12302), .Z(n12136) );
  AND U12839 ( .A(n12137), .B(n12136), .Z(n12231) );
  NAND U12840 ( .A(n185), .B(n12138), .Z(n12140) );
  XOR U12841 ( .A(b[9]), .B(a[88]), .Z(n12305) );
  NAND U12842 ( .A(n36805), .B(n12305), .Z(n12139) );
  NAND U12843 ( .A(n12140), .B(n12139), .Z(n12230) );
  XNOR U12844 ( .A(n12231), .B(n12230), .Z(n12232) );
  XOR U12845 ( .A(n12233), .B(n12232), .Z(n12239) );
  XOR U12846 ( .A(n12238), .B(n12239), .Z(n12245) );
  XOR U12847 ( .A(n12244), .B(n12245), .Z(n12257) );
  XNOR U12848 ( .A(n12256), .B(n12257), .Z(n12188) );
  XNOR U12849 ( .A(n12189), .B(n12188), .Z(n12190) );
  XOR U12850 ( .A(n12191), .B(n12190), .Z(n12309) );
  XOR U12851 ( .A(n12308), .B(n12309), .Z(n12311) );
  XOR U12852 ( .A(n12310), .B(n12311), .Z(n12185) );
  NANDN U12853 ( .A(n12142), .B(n12141), .Z(n12146) );
  NAND U12854 ( .A(n12144), .B(n12143), .Z(n12145) );
  AND U12855 ( .A(n12146), .B(n12145), .Z(n12183) );
  NANDN U12856 ( .A(n12148), .B(n12147), .Z(n12152) );
  NANDN U12857 ( .A(n12150), .B(n12149), .Z(n12151) );
  AND U12858 ( .A(n12152), .B(n12151), .Z(n12182) );
  XNOR U12859 ( .A(n12183), .B(n12182), .Z(n12184) );
  XNOR U12860 ( .A(n12185), .B(n12184), .Z(n12176) );
  NANDN U12861 ( .A(n12154), .B(n12153), .Z(n12158) );
  NANDN U12862 ( .A(n12156), .B(n12155), .Z(n12157) );
  NAND U12863 ( .A(n12158), .B(n12157), .Z(n12177) );
  XNOR U12864 ( .A(n12176), .B(n12177), .Z(n12178) );
  NANDN U12865 ( .A(n12160), .B(n12159), .Z(n12164) );
  NAND U12866 ( .A(n12162), .B(n12161), .Z(n12163) );
  NAND U12867 ( .A(n12164), .B(n12163), .Z(n12179) );
  XNOR U12868 ( .A(n12178), .B(n12179), .Z(n12170) );
  XNOR U12869 ( .A(n12171), .B(n12170), .Z(n12172) );
  XNOR U12870 ( .A(n12173), .B(n12172), .Z(n12314) );
  XNOR U12871 ( .A(sreg[320]), .B(n12314), .Z(n12316) );
  NANDN U12872 ( .A(sreg[319]), .B(n12165), .Z(n12169) );
  NAND U12873 ( .A(n12167), .B(n12166), .Z(n12168) );
  NAND U12874 ( .A(n12169), .B(n12168), .Z(n12315) );
  XNOR U12875 ( .A(n12316), .B(n12315), .Z(c[320]) );
  NANDN U12876 ( .A(n12171), .B(n12170), .Z(n12175) );
  NANDN U12877 ( .A(n12173), .B(n12172), .Z(n12174) );
  AND U12878 ( .A(n12175), .B(n12174), .Z(n12322) );
  NANDN U12879 ( .A(n12177), .B(n12176), .Z(n12181) );
  NANDN U12880 ( .A(n12179), .B(n12178), .Z(n12180) );
  AND U12881 ( .A(n12181), .B(n12180), .Z(n12320) );
  NANDN U12882 ( .A(n12183), .B(n12182), .Z(n12187) );
  NANDN U12883 ( .A(n12185), .B(n12184), .Z(n12186) );
  AND U12884 ( .A(n12187), .B(n12186), .Z(n12328) );
  NANDN U12885 ( .A(n12189), .B(n12188), .Z(n12193) );
  NANDN U12886 ( .A(n12191), .B(n12190), .Z(n12192) );
  AND U12887 ( .A(n12193), .B(n12192), .Z(n12332) );
  NANDN U12888 ( .A(n12195), .B(n12194), .Z(n12199) );
  NAND U12889 ( .A(n12197), .B(n12196), .Z(n12198) );
  AND U12890 ( .A(n12199), .B(n12198), .Z(n12331) );
  XNOR U12891 ( .A(n12332), .B(n12331), .Z(n12334) );
  NANDN U12892 ( .A(n12201), .B(n12200), .Z(n12205) );
  NANDN U12893 ( .A(n12203), .B(n12202), .Z(n12204) );
  AND U12894 ( .A(n12205), .B(n12204), .Z(n12411) );
  NAND U12895 ( .A(n38385), .B(n12206), .Z(n12208) );
  XOR U12896 ( .A(b[27]), .B(a[71]), .Z(n12355) );
  NAND U12897 ( .A(n38343), .B(n12355), .Z(n12207) );
  AND U12898 ( .A(n12208), .B(n12207), .Z(n12418) );
  NAND U12899 ( .A(n183), .B(n12209), .Z(n12211) );
  XOR U12900 ( .A(b[5]), .B(a[93]), .Z(n12358) );
  NAND U12901 ( .A(n36296), .B(n12358), .Z(n12210) );
  AND U12902 ( .A(n12211), .B(n12210), .Z(n12416) );
  NAND U12903 ( .A(n190), .B(n12212), .Z(n12214) );
  XOR U12904 ( .A(b[19]), .B(a[79]), .Z(n12361) );
  NAND U12905 ( .A(n37821), .B(n12361), .Z(n12213) );
  NAND U12906 ( .A(n12214), .B(n12213), .Z(n12415) );
  XNOR U12907 ( .A(n12416), .B(n12415), .Z(n12417) );
  XNOR U12908 ( .A(n12418), .B(n12417), .Z(n12409) );
  NAND U12909 ( .A(n38470), .B(n12215), .Z(n12217) );
  XOR U12910 ( .A(b[31]), .B(a[67]), .Z(n12364) );
  NAND U12911 ( .A(n38453), .B(n12364), .Z(n12216) );
  AND U12912 ( .A(n12217), .B(n12216), .Z(n12376) );
  NAND U12913 ( .A(n181), .B(n12218), .Z(n12220) );
  XOR U12914 ( .A(b[3]), .B(a[95]), .Z(n12367) );
  NAND U12915 ( .A(n182), .B(n12367), .Z(n12219) );
  AND U12916 ( .A(n12220), .B(n12219), .Z(n12374) );
  NAND U12917 ( .A(n189), .B(n12221), .Z(n12223) );
  XOR U12918 ( .A(b[17]), .B(a[81]), .Z(n12370) );
  NAND U12919 ( .A(n37652), .B(n12370), .Z(n12222) );
  NAND U12920 ( .A(n12223), .B(n12222), .Z(n12373) );
  XNOR U12921 ( .A(n12374), .B(n12373), .Z(n12375) );
  XOR U12922 ( .A(n12376), .B(n12375), .Z(n12410) );
  XOR U12923 ( .A(n12409), .B(n12410), .Z(n12412) );
  XOR U12924 ( .A(n12411), .B(n12412), .Z(n12344) );
  NANDN U12925 ( .A(n12225), .B(n12224), .Z(n12229) );
  NANDN U12926 ( .A(n12227), .B(n12226), .Z(n12228) );
  AND U12927 ( .A(n12229), .B(n12228), .Z(n12397) );
  NANDN U12928 ( .A(n12231), .B(n12230), .Z(n12235) );
  NANDN U12929 ( .A(n12233), .B(n12232), .Z(n12234) );
  NAND U12930 ( .A(n12235), .B(n12234), .Z(n12398) );
  XNOR U12931 ( .A(n12397), .B(n12398), .Z(n12399) );
  NANDN U12932 ( .A(n12237), .B(n12236), .Z(n12241) );
  NANDN U12933 ( .A(n12239), .B(n12238), .Z(n12240) );
  NAND U12934 ( .A(n12241), .B(n12240), .Z(n12400) );
  XNOR U12935 ( .A(n12399), .B(n12400), .Z(n12343) );
  XNOR U12936 ( .A(n12344), .B(n12343), .Z(n12346) );
  NANDN U12937 ( .A(n12243), .B(n12242), .Z(n12247) );
  NANDN U12938 ( .A(n12245), .B(n12244), .Z(n12246) );
  AND U12939 ( .A(n12247), .B(n12246), .Z(n12345) );
  XOR U12940 ( .A(n12346), .B(n12345), .Z(n12460) );
  NANDN U12941 ( .A(n12249), .B(n12248), .Z(n12253) );
  NANDN U12942 ( .A(n12251), .B(n12250), .Z(n12252) );
  AND U12943 ( .A(n12253), .B(n12252), .Z(n12457) );
  NANDN U12944 ( .A(n12255), .B(n12254), .Z(n12259) );
  NANDN U12945 ( .A(n12257), .B(n12256), .Z(n12258) );
  AND U12946 ( .A(n12259), .B(n12258), .Z(n12340) );
  NANDN U12947 ( .A(n12261), .B(n12260), .Z(n12265) );
  OR U12948 ( .A(n12263), .B(n12262), .Z(n12264) );
  AND U12949 ( .A(n12265), .B(n12264), .Z(n12338) );
  NANDN U12950 ( .A(n12267), .B(n12266), .Z(n12271) );
  NANDN U12951 ( .A(n12269), .B(n12268), .Z(n12270) );
  AND U12952 ( .A(n12271), .B(n12270), .Z(n12404) );
  NANDN U12953 ( .A(n12273), .B(n12272), .Z(n12277) );
  NANDN U12954 ( .A(n12275), .B(n12274), .Z(n12276) );
  NAND U12955 ( .A(n12277), .B(n12276), .Z(n12403) );
  XNOR U12956 ( .A(n12404), .B(n12403), .Z(n12405) );
  NAND U12957 ( .A(b[0]), .B(a[97]), .Z(n12278) );
  XNOR U12958 ( .A(b[1]), .B(n12278), .Z(n12280) );
  NANDN U12959 ( .A(b[0]), .B(a[96]), .Z(n12279) );
  NAND U12960 ( .A(n12280), .B(n12279), .Z(n12352) );
  NAND U12961 ( .A(n194), .B(n12281), .Z(n12283) );
  XOR U12962 ( .A(b[29]), .B(a[69]), .Z(n12430) );
  NAND U12963 ( .A(n38456), .B(n12430), .Z(n12282) );
  AND U12964 ( .A(n12283), .B(n12282), .Z(n12350) );
  AND U12965 ( .A(b[31]), .B(a[65]), .Z(n12349) );
  XNOR U12966 ( .A(n12350), .B(n12349), .Z(n12351) );
  XNOR U12967 ( .A(n12352), .B(n12351), .Z(n12391) );
  NAND U12968 ( .A(n38185), .B(n12284), .Z(n12286) );
  XOR U12969 ( .A(b[23]), .B(a[75]), .Z(n12433) );
  NAND U12970 ( .A(n38132), .B(n12433), .Z(n12285) );
  AND U12971 ( .A(n12286), .B(n12285), .Z(n12424) );
  NAND U12972 ( .A(n184), .B(n12287), .Z(n12289) );
  XOR U12973 ( .A(b[7]), .B(a[91]), .Z(n12436) );
  NAND U12974 ( .A(n36592), .B(n12436), .Z(n12288) );
  AND U12975 ( .A(n12289), .B(n12288), .Z(n12422) );
  NAND U12976 ( .A(n38289), .B(n12290), .Z(n12292) );
  XOR U12977 ( .A(b[25]), .B(a[73]), .Z(n12439) );
  NAND U12978 ( .A(n38247), .B(n12439), .Z(n12291) );
  NAND U12979 ( .A(n12292), .B(n12291), .Z(n12421) );
  XNOR U12980 ( .A(n12422), .B(n12421), .Z(n12423) );
  XOR U12981 ( .A(n12424), .B(n12423), .Z(n12392) );
  XNOR U12982 ( .A(n12391), .B(n12392), .Z(n12393) );
  NAND U12983 ( .A(n187), .B(n12293), .Z(n12295) );
  XOR U12984 ( .A(b[13]), .B(a[85]), .Z(n12442) );
  NAND U12985 ( .A(n37295), .B(n12442), .Z(n12294) );
  AND U12986 ( .A(n12295), .B(n12294), .Z(n12386) );
  NAND U12987 ( .A(n186), .B(n12296), .Z(n12298) );
  XOR U12988 ( .A(b[11]), .B(a[87]), .Z(n12445) );
  NAND U12989 ( .A(n37097), .B(n12445), .Z(n12297) );
  NAND U12990 ( .A(n12298), .B(n12297), .Z(n12385) );
  XNOR U12991 ( .A(n12386), .B(n12385), .Z(n12387) );
  NAND U12992 ( .A(n188), .B(n12299), .Z(n12301) );
  XOR U12993 ( .A(b[15]), .B(a[83]), .Z(n12448) );
  NAND U12994 ( .A(n37382), .B(n12448), .Z(n12300) );
  AND U12995 ( .A(n12301), .B(n12300), .Z(n12382) );
  NAND U12996 ( .A(n38064), .B(n12302), .Z(n12304) );
  XOR U12997 ( .A(b[21]), .B(a[77]), .Z(n12451) );
  NAND U12998 ( .A(n37993), .B(n12451), .Z(n12303) );
  AND U12999 ( .A(n12304), .B(n12303), .Z(n12380) );
  NAND U13000 ( .A(n185), .B(n12305), .Z(n12307) );
  XOR U13001 ( .A(b[9]), .B(a[89]), .Z(n12454) );
  NAND U13002 ( .A(n36805), .B(n12454), .Z(n12306) );
  NAND U13003 ( .A(n12307), .B(n12306), .Z(n12379) );
  XNOR U13004 ( .A(n12380), .B(n12379), .Z(n12381) );
  XOR U13005 ( .A(n12382), .B(n12381), .Z(n12388) );
  XOR U13006 ( .A(n12387), .B(n12388), .Z(n12394) );
  XOR U13007 ( .A(n12393), .B(n12394), .Z(n12406) );
  XNOR U13008 ( .A(n12405), .B(n12406), .Z(n12337) );
  XNOR U13009 ( .A(n12338), .B(n12337), .Z(n12339) );
  XOR U13010 ( .A(n12340), .B(n12339), .Z(n12458) );
  XNOR U13011 ( .A(n12457), .B(n12458), .Z(n12459) );
  XNOR U13012 ( .A(n12460), .B(n12459), .Z(n12333) );
  XOR U13013 ( .A(n12334), .B(n12333), .Z(n12326) );
  NANDN U13014 ( .A(n12309), .B(n12308), .Z(n12313) );
  OR U13015 ( .A(n12311), .B(n12310), .Z(n12312) );
  AND U13016 ( .A(n12313), .B(n12312), .Z(n12325) );
  XNOR U13017 ( .A(n12326), .B(n12325), .Z(n12327) );
  XNOR U13018 ( .A(n12328), .B(n12327), .Z(n12319) );
  XNOR U13019 ( .A(n12320), .B(n12319), .Z(n12321) );
  XNOR U13020 ( .A(n12322), .B(n12321), .Z(n12463) );
  XNOR U13021 ( .A(sreg[321]), .B(n12463), .Z(n12465) );
  NANDN U13022 ( .A(sreg[320]), .B(n12314), .Z(n12318) );
  NAND U13023 ( .A(n12316), .B(n12315), .Z(n12317) );
  NAND U13024 ( .A(n12318), .B(n12317), .Z(n12464) );
  XNOR U13025 ( .A(n12465), .B(n12464), .Z(c[321]) );
  NANDN U13026 ( .A(n12320), .B(n12319), .Z(n12324) );
  NANDN U13027 ( .A(n12322), .B(n12321), .Z(n12323) );
  AND U13028 ( .A(n12324), .B(n12323), .Z(n12471) );
  NANDN U13029 ( .A(n12326), .B(n12325), .Z(n12330) );
  NANDN U13030 ( .A(n12328), .B(n12327), .Z(n12329) );
  AND U13031 ( .A(n12330), .B(n12329), .Z(n12469) );
  NANDN U13032 ( .A(n12332), .B(n12331), .Z(n12336) );
  NAND U13033 ( .A(n12334), .B(n12333), .Z(n12335) );
  AND U13034 ( .A(n12336), .B(n12335), .Z(n12476) );
  NANDN U13035 ( .A(n12338), .B(n12337), .Z(n12342) );
  NANDN U13036 ( .A(n12340), .B(n12339), .Z(n12341) );
  AND U13037 ( .A(n12342), .B(n12341), .Z(n12607) );
  NANDN U13038 ( .A(n12344), .B(n12343), .Z(n12348) );
  NAND U13039 ( .A(n12346), .B(n12345), .Z(n12347) );
  AND U13040 ( .A(n12348), .B(n12347), .Z(n12606) );
  XNOR U13041 ( .A(n12607), .B(n12606), .Z(n12609) );
  NANDN U13042 ( .A(n12350), .B(n12349), .Z(n12354) );
  NANDN U13043 ( .A(n12352), .B(n12351), .Z(n12353) );
  AND U13044 ( .A(n12354), .B(n12353), .Z(n12554) );
  NAND U13045 ( .A(n38385), .B(n12355), .Z(n12357) );
  XOR U13046 ( .A(b[27]), .B(a[72]), .Z(n12498) );
  NAND U13047 ( .A(n38343), .B(n12498), .Z(n12356) );
  AND U13048 ( .A(n12357), .B(n12356), .Z(n12561) );
  NAND U13049 ( .A(n183), .B(n12358), .Z(n12360) );
  XOR U13050 ( .A(b[5]), .B(a[94]), .Z(n12501) );
  NAND U13051 ( .A(n36296), .B(n12501), .Z(n12359) );
  AND U13052 ( .A(n12360), .B(n12359), .Z(n12559) );
  NAND U13053 ( .A(n190), .B(n12361), .Z(n12363) );
  XOR U13054 ( .A(b[19]), .B(a[80]), .Z(n12504) );
  NAND U13055 ( .A(n37821), .B(n12504), .Z(n12362) );
  NAND U13056 ( .A(n12363), .B(n12362), .Z(n12558) );
  XNOR U13057 ( .A(n12559), .B(n12558), .Z(n12560) );
  XNOR U13058 ( .A(n12561), .B(n12560), .Z(n12552) );
  NAND U13059 ( .A(n38470), .B(n12364), .Z(n12366) );
  XOR U13060 ( .A(b[31]), .B(a[68]), .Z(n12507) );
  NAND U13061 ( .A(n38453), .B(n12507), .Z(n12365) );
  AND U13062 ( .A(n12366), .B(n12365), .Z(n12519) );
  NAND U13063 ( .A(n181), .B(n12367), .Z(n12369) );
  XOR U13064 ( .A(b[3]), .B(a[96]), .Z(n12510) );
  NAND U13065 ( .A(n182), .B(n12510), .Z(n12368) );
  AND U13066 ( .A(n12369), .B(n12368), .Z(n12517) );
  NAND U13067 ( .A(n189), .B(n12370), .Z(n12372) );
  XOR U13068 ( .A(b[17]), .B(a[82]), .Z(n12513) );
  NAND U13069 ( .A(n37652), .B(n12513), .Z(n12371) );
  NAND U13070 ( .A(n12372), .B(n12371), .Z(n12516) );
  XNOR U13071 ( .A(n12517), .B(n12516), .Z(n12518) );
  XOR U13072 ( .A(n12519), .B(n12518), .Z(n12553) );
  XOR U13073 ( .A(n12552), .B(n12553), .Z(n12555) );
  XOR U13074 ( .A(n12554), .B(n12555), .Z(n12487) );
  NANDN U13075 ( .A(n12374), .B(n12373), .Z(n12378) );
  NANDN U13076 ( .A(n12376), .B(n12375), .Z(n12377) );
  AND U13077 ( .A(n12378), .B(n12377), .Z(n12540) );
  NANDN U13078 ( .A(n12380), .B(n12379), .Z(n12384) );
  NANDN U13079 ( .A(n12382), .B(n12381), .Z(n12383) );
  NAND U13080 ( .A(n12384), .B(n12383), .Z(n12541) );
  XNOR U13081 ( .A(n12540), .B(n12541), .Z(n12542) );
  NANDN U13082 ( .A(n12386), .B(n12385), .Z(n12390) );
  NANDN U13083 ( .A(n12388), .B(n12387), .Z(n12389) );
  NAND U13084 ( .A(n12390), .B(n12389), .Z(n12543) );
  XNOR U13085 ( .A(n12542), .B(n12543), .Z(n12486) );
  XNOR U13086 ( .A(n12487), .B(n12486), .Z(n12489) );
  NANDN U13087 ( .A(n12392), .B(n12391), .Z(n12396) );
  NANDN U13088 ( .A(n12394), .B(n12393), .Z(n12395) );
  AND U13089 ( .A(n12396), .B(n12395), .Z(n12488) );
  XOR U13090 ( .A(n12489), .B(n12488), .Z(n12603) );
  NANDN U13091 ( .A(n12398), .B(n12397), .Z(n12402) );
  NANDN U13092 ( .A(n12400), .B(n12399), .Z(n12401) );
  AND U13093 ( .A(n12402), .B(n12401), .Z(n12600) );
  NANDN U13094 ( .A(n12404), .B(n12403), .Z(n12408) );
  NANDN U13095 ( .A(n12406), .B(n12405), .Z(n12407) );
  AND U13096 ( .A(n12408), .B(n12407), .Z(n12483) );
  NANDN U13097 ( .A(n12410), .B(n12409), .Z(n12414) );
  OR U13098 ( .A(n12412), .B(n12411), .Z(n12413) );
  AND U13099 ( .A(n12414), .B(n12413), .Z(n12481) );
  NANDN U13100 ( .A(n12416), .B(n12415), .Z(n12420) );
  NANDN U13101 ( .A(n12418), .B(n12417), .Z(n12419) );
  AND U13102 ( .A(n12420), .B(n12419), .Z(n12547) );
  NANDN U13103 ( .A(n12422), .B(n12421), .Z(n12426) );
  NANDN U13104 ( .A(n12424), .B(n12423), .Z(n12425) );
  NAND U13105 ( .A(n12426), .B(n12425), .Z(n12546) );
  XNOR U13106 ( .A(n12547), .B(n12546), .Z(n12548) );
  NAND U13107 ( .A(b[0]), .B(a[98]), .Z(n12427) );
  XNOR U13108 ( .A(b[1]), .B(n12427), .Z(n12429) );
  NANDN U13109 ( .A(b[0]), .B(a[97]), .Z(n12428) );
  NAND U13110 ( .A(n12429), .B(n12428), .Z(n12495) );
  NAND U13111 ( .A(n194), .B(n12430), .Z(n12432) );
  XOR U13112 ( .A(b[29]), .B(a[70]), .Z(n12573) );
  NAND U13113 ( .A(n38456), .B(n12573), .Z(n12431) );
  AND U13114 ( .A(n12432), .B(n12431), .Z(n12493) );
  AND U13115 ( .A(b[31]), .B(a[66]), .Z(n12492) );
  XNOR U13116 ( .A(n12493), .B(n12492), .Z(n12494) );
  XNOR U13117 ( .A(n12495), .B(n12494), .Z(n12534) );
  NAND U13118 ( .A(n38185), .B(n12433), .Z(n12435) );
  XOR U13119 ( .A(b[23]), .B(a[76]), .Z(n12576) );
  NAND U13120 ( .A(n38132), .B(n12576), .Z(n12434) );
  AND U13121 ( .A(n12435), .B(n12434), .Z(n12567) );
  NAND U13122 ( .A(n184), .B(n12436), .Z(n12438) );
  XOR U13123 ( .A(b[7]), .B(a[92]), .Z(n12579) );
  NAND U13124 ( .A(n36592), .B(n12579), .Z(n12437) );
  AND U13125 ( .A(n12438), .B(n12437), .Z(n12565) );
  NAND U13126 ( .A(n38289), .B(n12439), .Z(n12441) );
  XOR U13127 ( .A(b[25]), .B(a[74]), .Z(n12582) );
  NAND U13128 ( .A(n38247), .B(n12582), .Z(n12440) );
  NAND U13129 ( .A(n12441), .B(n12440), .Z(n12564) );
  XNOR U13130 ( .A(n12565), .B(n12564), .Z(n12566) );
  XOR U13131 ( .A(n12567), .B(n12566), .Z(n12535) );
  XNOR U13132 ( .A(n12534), .B(n12535), .Z(n12536) );
  NAND U13133 ( .A(n187), .B(n12442), .Z(n12444) );
  XOR U13134 ( .A(b[13]), .B(a[86]), .Z(n12585) );
  NAND U13135 ( .A(n37295), .B(n12585), .Z(n12443) );
  AND U13136 ( .A(n12444), .B(n12443), .Z(n12529) );
  NAND U13137 ( .A(n186), .B(n12445), .Z(n12447) );
  XOR U13138 ( .A(b[11]), .B(a[88]), .Z(n12588) );
  NAND U13139 ( .A(n37097), .B(n12588), .Z(n12446) );
  NAND U13140 ( .A(n12447), .B(n12446), .Z(n12528) );
  XNOR U13141 ( .A(n12529), .B(n12528), .Z(n12530) );
  NAND U13142 ( .A(n188), .B(n12448), .Z(n12450) );
  XOR U13143 ( .A(b[15]), .B(a[84]), .Z(n12591) );
  NAND U13144 ( .A(n37382), .B(n12591), .Z(n12449) );
  AND U13145 ( .A(n12450), .B(n12449), .Z(n12525) );
  NAND U13146 ( .A(n38064), .B(n12451), .Z(n12453) );
  XOR U13147 ( .A(b[21]), .B(a[78]), .Z(n12594) );
  NAND U13148 ( .A(n37993), .B(n12594), .Z(n12452) );
  AND U13149 ( .A(n12453), .B(n12452), .Z(n12523) );
  NAND U13150 ( .A(n185), .B(n12454), .Z(n12456) );
  XOR U13151 ( .A(b[9]), .B(a[90]), .Z(n12597) );
  NAND U13152 ( .A(n36805), .B(n12597), .Z(n12455) );
  NAND U13153 ( .A(n12456), .B(n12455), .Z(n12522) );
  XNOR U13154 ( .A(n12523), .B(n12522), .Z(n12524) );
  XOR U13155 ( .A(n12525), .B(n12524), .Z(n12531) );
  XOR U13156 ( .A(n12530), .B(n12531), .Z(n12537) );
  XOR U13157 ( .A(n12536), .B(n12537), .Z(n12549) );
  XNOR U13158 ( .A(n12548), .B(n12549), .Z(n12480) );
  XNOR U13159 ( .A(n12481), .B(n12480), .Z(n12482) );
  XOR U13160 ( .A(n12483), .B(n12482), .Z(n12601) );
  XNOR U13161 ( .A(n12600), .B(n12601), .Z(n12602) );
  XNOR U13162 ( .A(n12603), .B(n12602), .Z(n12608) );
  XOR U13163 ( .A(n12609), .B(n12608), .Z(n12475) );
  NANDN U13164 ( .A(n12458), .B(n12457), .Z(n12462) );
  NANDN U13165 ( .A(n12460), .B(n12459), .Z(n12461) );
  AND U13166 ( .A(n12462), .B(n12461), .Z(n12474) );
  XOR U13167 ( .A(n12475), .B(n12474), .Z(n12477) );
  XNOR U13168 ( .A(n12476), .B(n12477), .Z(n12468) );
  XNOR U13169 ( .A(n12469), .B(n12468), .Z(n12470) );
  XNOR U13170 ( .A(n12471), .B(n12470), .Z(n12612) );
  XNOR U13171 ( .A(sreg[322]), .B(n12612), .Z(n12614) );
  NANDN U13172 ( .A(sreg[321]), .B(n12463), .Z(n12467) );
  NAND U13173 ( .A(n12465), .B(n12464), .Z(n12466) );
  NAND U13174 ( .A(n12467), .B(n12466), .Z(n12613) );
  XNOR U13175 ( .A(n12614), .B(n12613), .Z(c[322]) );
  NANDN U13176 ( .A(n12469), .B(n12468), .Z(n12473) );
  NANDN U13177 ( .A(n12471), .B(n12470), .Z(n12472) );
  AND U13178 ( .A(n12473), .B(n12472), .Z(n12620) );
  NANDN U13179 ( .A(n12475), .B(n12474), .Z(n12479) );
  NANDN U13180 ( .A(n12477), .B(n12476), .Z(n12478) );
  AND U13181 ( .A(n12479), .B(n12478), .Z(n12618) );
  NANDN U13182 ( .A(n12481), .B(n12480), .Z(n12485) );
  NANDN U13183 ( .A(n12483), .B(n12482), .Z(n12484) );
  AND U13184 ( .A(n12485), .B(n12484), .Z(n12630) );
  NANDN U13185 ( .A(n12487), .B(n12486), .Z(n12491) );
  NAND U13186 ( .A(n12489), .B(n12488), .Z(n12490) );
  AND U13187 ( .A(n12491), .B(n12490), .Z(n12629) );
  XNOR U13188 ( .A(n12630), .B(n12629), .Z(n12632) );
  NANDN U13189 ( .A(n12493), .B(n12492), .Z(n12497) );
  NANDN U13190 ( .A(n12495), .B(n12494), .Z(n12496) );
  AND U13191 ( .A(n12497), .B(n12496), .Z(n12707) );
  NAND U13192 ( .A(n38385), .B(n12498), .Z(n12500) );
  XOR U13193 ( .A(b[27]), .B(a[73]), .Z(n12653) );
  NAND U13194 ( .A(n38343), .B(n12653), .Z(n12499) );
  AND U13195 ( .A(n12500), .B(n12499), .Z(n12714) );
  NAND U13196 ( .A(n183), .B(n12501), .Z(n12503) );
  XOR U13197 ( .A(b[5]), .B(a[95]), .Z(n12656) );
  NAND U13198 ( .A(n36296), .B(n12656), .Z(n12502) );
  AND U13199 ( .A(n12503), .B(n12502), .Z(n12712) );
  NAND U13200 ( .A(n190), .B(n12504), .Z(n12506) );
  XOR U13201 ( .A(b[19]), .B(a[81]), .Z(n12659) );
  NAND U13202 ( .A(n37821), .B(n12659), .Z(n12505) );
  NAND U13203 ( .A(n12506), .B(n12505), .Z(n12711) );
  XNOR U13204 ( .A(n12712), .B(n12711), .Z(n12713) );
  XNOR U13205 ( .A(n12714), .B(n12713), .Z(n12705) );
  NAND U13206 ( .A(n38470), .B(n12507), .Z(n12509) );
  XOR U13207 ( .A(b[31]), .B(a[69]), .Z(n12662) );
  NAND U13208 ( .A(n38453), .B(n12662), .Z(n12508) );
  AND U13209 ( .A(n12509), .B(n12508), .Z(n12674) );
  NAND U13210 ( .A(n181), .B(n12510), .Z(n12512) );
  XOR U13211 ( .A(b[3]), .B(a[97]), .Z(n12665) );
  NAND U13212 ( .A(n182), .B(n12665), .Z(n12511) );
  AND U13213 ( .A(n12512), .B(n12511), .Z(n12672) );
  NAND U13214 ( .A(n189), .B(n12513), .Z(n12515) );
  XOR U13215 ( .A(b[17]), .B(a[83]), .Z(n12668) );
  NAND U13216 ( .A(n37652), .B(n12668), .Z(n12514) );
  NAND U13217 ( .A(n12515), .B(n12514), .Z(n12671) );
  XNOR U13218 ( .A(n12672), .B(n12671), .Z(n12673) );
  XOR U13219 ( .A(n12674), .B(n12673), .Z(n12706) );
  XOR U13220 ( .A(n12705), .B(n12706), .Z(n12708) );
  XOR U13221 ( .A(n12707), .B(n12708), .Z(n12642) );
  NANDN U13222 ( .A(n12517), .B(n12516), .Z(n12521) );
  NANDN U13223 ( .A(n12519), .B(n12518), .Z(n12520) );
  AND U13224 ( .A(n12521), .B(n12520), .Z(n12695) );
  NANDN U13225 ( .A(n12523), .B(n12522), .Z(n12527) );
  NANDN U13226 ( .A(n12525), .B(n12524), .Z(n12526) );
  NAND U13227 ( .A(n12527), .B(n12526), .Z(n12696) );
  XNOR U13228 ( .A(n12695), .B(n12696), .Z(n12697) );
  NANDN U13229 ( .A(n12529), .B(n12528), .Z(n12533) );
  NANDN U13230 ( .A(n12531), .B(n12530), .Z(n12532) );
  NAND U13231 ( .A(n12533), .B(n12532), .Z(n12698) );
  XNOR U13232 ( .A(n12697), .B(n12698), .Z(n12641) );
  XNOR U13233 ( .A(n12642), .B(n12641), .Z(n12644) );
  NANDN U13234 ( .A(n12535), .B(n12534), .Z(n12539) );
  NANDN U13235 ( .A(n12537), .B(n12536), .Z(n12538) );
  AND U13236 ( .A(n12539), .B(n12538), .Z(n12643) );
  XOR U13237 ( .A(n12644), .B(n12643), .Z(n12756) );
  NANDN U13238 ( .A(n12541), .B(n12540), .Z(n12545) );
  NANDN U13239 ( .A(n12543), .B(n12542), .Z(n12544) );
  AND U13240 ( .A(n12545), .B(n12544), .Z(n12753) );
  NANDN U13241 ( .A(n12547), .B(n12546), .Z(n12551) );
  NANDN U13242 ( .A(n12549), .B(n12548), .Z(n12550) );
  AND U13243 ( .A(n12551), .B(n12550), .Z(n12638) );
  NANDN U13244 ( .A(n12553), .B(n12552), .Z(n12557) );
  OR U13245 ( .A(n12555), .B(n12554), .Z(n12556) );
  AND U13246 ( .A(n12557), .B(n12556), .Z(n12636) );
  NANDN U13247 ( .A(n12559), .B(n12558), .Z(n12563) );
  NANDN U13248 ( .A(n12561), .B(n12560), .Z(n12562) );
  AND U13249 ( .A(n12563), .B(n12562), .Z(n12702) );
  NANDN U13250 ( .A(n12565), .B(n12564), .Z(n12569) );
  NANDN U13251 ( .A(n12567), .B(n12566), .Z(n12568) );
  NAND U13252 ( .A(n12569), .B(n12568), .Z(n12701) );
  XNOR U13253 ( .A(n12702), .B(n12701), .Z(n12704) );
  NAND U13254 ( .A(b[0]), .B(a[99]), .Z(n12570) );
  XNOR U13255 ( .A(b[1]), .B(n12570), .Z(n12572) );
  NANDN U13256 ( .A(b[0]), .B(a[98]), .Z(n12571) );
  NAND U13257 ( .A(n12572), .B(n12571), .Z(n12650) );
  NAND U13258 ( .A(n194), .B(n12573), .Z(n12575) );
  XOR U13259 ( .A(b[29]), .B(a[71]), .Z(n12726) );
  NAND U13260 ( .A(n38456), .B(n12726), .Z(n12574) );
  AND U13261 ( .A(n12575), .B(n12574), .Z(n12648) );
  AND U13262 ( .A(b[31]), .B(a[67]), .Z(n12647) );
  XNOR U13263 ( .A(n12648), .B(n12647), .Z(n12649) );
  XNOR U13264 ( .A(n12650), .B(n12649), .Z(n12690) );
  NAND U13265 ( .A(n38185), .B(n12576), .Z(n12578) );
  XOR U13266 ( .A(b[23]), .B(a[77]), .Z(n12729) );
  NAND U13267 ( .A(n38132), .B(n12729), .Z(n12577) );
  AND U13268 ( .A(n12578), .B(n12577), .Z(n12719) );
  NAND U13269 ( .A(n184), .B(n12579), .Z(n12581) );
  XOR U13270 ( .A(b[7]), .B(a[93]), .Z(n12732) );
  NAND U13271 ( .A(n36592), .B(n12732), .Z(n12580) );
  AND U13272 ( .A(n12581), .B(n12580), .Z(n12718) );
  NAND U13273 ( .A(n38289), .B(n12582), .Z(n12584) );
  XOR U13274 ( .A(b[25]), .B(a[75]), .Z(n12735) );
  NAND U13275 ( .A(n38247), .B(n12735), .Z(n12583) );
  NAND U13276 ( .A(n12584), .B(n12583), .Z(n12717) );
  XOR U13277 ( .A(n12718), .B(n12717), .Z(n12720) );
  XOR U13278 ( .A(n12719), .B(n12720), .Z(n12689) );
  XOR U13279 ( .A(n12690), .B(n12689), .Z(n12692) );
  NAND U13280 ( .A(n187), .B(n12585), .Z(n12587) );
  XOR U13281 ( .A(b[13]), .B(a[87]), .Z(n12738) );
  NAND U13282 ( .A(n37295), .B(n12738), .Z(n12586) );
  AND U13283 ( .A(n12587), .B(n12586), .Z(n12684) );
  NAND U13284 ( .A(n186), .B(n12588), .Z(n12590) );
  XOR U13285 ( .A(b[11]), .B(a[89]), .Z(n12741) );
  NAND U13286 ( .A(n37097), .B(n12741), .Z(n12589) );
  NAND U13287 ( .A(n12590), .B(n12589), .Z(n12683) );
  XNOR U13288 ( .A(n12684), .B(n12683), .Z(n12686) );
  NAND U13289 ( .A(n188), .B(n12591), .Z(n12593) );
  XOR U13290 ( .A(b[15]), .B(a[85]), .Z(n12744) );
  NAND U13291 ( .A(n37382), .B(n12744), .Z(n12592) );
  AND U13292 ( .A(n12593), .B(n12592), .Z(n12680) );
  NAND U13293 ( .A(n38064), .B(n12594), .Z(n12596) );
  XOR U13294 ( .A(b[21]), .B(a[79]), .Z(n12747) );
  NAND U13295 ( .A(n37993), .B(n12747), .Z(n12595) );
  AND U13296 ( .A(n12596), .B(n12595), .Z(n12678) );
  NAND U13297 ( .A(n185), .B(n12597), .Z(n12599) );
  XOR U13298 ( .A(b[9]), .B(a[91]), .Z(n12750) );
  NAND U13299 ( .A(n36805), .B(n12750), .Z(n12598) );
  NAND U13300 ( .A(n12599), .B(n12598), .Z(n12677) );
  XNOR U13301 ( .A(n12678), .B(n12677), .Z(n12679) );
  XNOR U13302 ( .A(n12680), .B(n12679), .Z(n12685) );
  XOR U13303 ( .A(n12686), .B(n12685), .Z(n12691) );
  XNOR U13304 ( .A(n12692), .B(n12691), .Z(n12703) );
  XNOR U13305 ( .A(n12704), .B(n12703), .Z(n12635) );
  XNOR U13306 ( .A(n12636), .B(n12635), .Z(n12637) );
  XOR U13307 ( .A(n12638), .B(n12637), .Z(n12754) );
  XNOR U13308 ( .A(n12753), .B(n12754), .Z(n12755) );
  XNOR U13309 ( .A(n12756), .B(n12755), .Z(n12631) );
  XOR U13310 ( .A(n12632), .B(n12631), .Z(n12624) );
  NANDN U13311 ( .A(n12601), .B(n12600), .Z(n12605) );
  NANDN U13312 ( .A(n12603), .B(n12602), .Z(n12604) );
  AND U13313 ( .A(n12605), .B(n12604), .Z(n12623) );
  XNOR U13314 ( .A(n12624), .B(n12623), .Z(n12625) );
  NANDN U13315 ( .A(n12607), .B(n12606), .Z(n12611) );
  NAND U13316 ( .A(n12609), .B(n12608), .Z(n12610) );
  NAND U13317 ( .A(n12611), .B(n12610), .Z(n12626) );
  XNOR U13318 ( .A(n12625), .B(n12626), .Z(n12617) );
  XNOR U13319 ( .A(n12618), .B(n12617), .Z(n12619) );
  XNOR U13320 ( .A(n12620), .B(n12619), .Z(n12759) );
  XNOR U13321 ( .A(sreg[323]), .B(n12759), .Z(n12761) );
  NANDN U13322 ( .A(sreg[322]), .B(n12612), .Z(n12616) );
  NAND U13323 ( .A(n12614), .B(n12613), .Z(n12615) );
  NAND U13324 ( .A(n12616), .B(n12615), .Z(n12760) );
  XNOR U13325 ( .A(n12761), .B(n12760), .Z(c[323]) );
  NANDN U13326 ( .A(n12618), .B(n12617), .Z(n12622) );
  NANDN U13327 ( .A(n12620), .B(n12619), .Z(n12621) );
  AND U13328 ( .A(n12622), .B(n12621), .Z(n12767) );
  NANDN U13329 ( .A(n12624), .B(n12623), .Z(n12628) );
  NANDN U13330 ( .A(n12626), .B(n12625), .Z(n12627) );
  AND U13331 ( .A(n12628), .B(n12627), .Z(n12765) );
  NANDN U13332 ( .A(n12630), .B(n12629), .Z(n12634) );
  NAND U13333 ( .A(n12632), .B(n12631), .Z(n12633) );
  AND U13334 ( .A(n12634), .B(n12633), .Z(n12772) );
  NANDN U13335 ( .A(n12636), .B(n12635), .Z(n12640) );
  NANDN U13336 ( .A(n12638), .B(n12637), .Z(n12639) );
  AND U13337 ( .A(n12640), .B(n12639), .Z(n12903) );
  NANDN U13338 ( .A(n12642), .B(n12641), .Z(n12646) );
  NAND U13339 ( .A(n12644), .B(n12643), .Z(n12645) );
  AND U13340 ( .A(n12646), .B(n12645), .Z(n12902) );
  XNOR U13341 ( .A(n12903), .B(n12902), .Z(n12905) );
  NANDN U13342 ( .A(n12648), .B(n12647), .Z(n12652) );
  NANDN U13343 ( .A(n12650), .B(n12649), .Z(n12651) );
  AND U13344 ( .A(n12652), .B(n12651), .Z(n12838) );
  NAND U13345 ( .A(n38385), .B(n12653), .Z(n12655) );
  XOR U13346 ( .A(b[27]), .B(a[74]), .Z(n12782) );
  NAND U13347 ( .A(n38343), .B(n12782), .Z(n12654) );
  AND U13348 ( .A(n12655), .B(n12654), .Z(n12845) );
  NAND U13349 ( .A(n183), .B(n12656), .Z(n12658) );
  XOR U13350 ( .A(b[5]), .B(a[96]), .Z(n12785) );
  NAND U13351 ( .A(n36296), .B(n12785), .Z(n12657) );
  AND U13352 ( .A(n12658), .B(n12657), .Z(n12843) );
  NAND U13353 ( .A(n190), .B(n12659), .Z(n12661) );
  XOR U13354 ( .A(b[19]), .B(a[82]), .Z(n12788) );
  NAND U13355 ( .A(n37821), .B(n12788), .Z(n12660) );
  NAND U13356 ( .A(n12661), .B(n12660), .Z(n12842) );
  XNOR U13357 ( .A(n12843), .B(n12842), .Z(n12844) );
  XNOR U13358 ( .A(n12845), .B(n12844), .Z(n12836) );
  NAND U13359 ( .A(n38470), .B(n12662), .Z(n12664) );
  XOR U13360 ( .A(b[31]), .B(a[70]), .Z(n12791) );
  NAND U13361 ( .A(n38453), .B(n12791), .Z(n12663) );
  AND U13362 ( .A(n12664), .B(n12663), .Z(n12803) );
  NAND U13363 ( .A(n181), .B(n12665), .Z(n12667) );
  XOR U13364 ( .A(b[3]), .B(a[98]), .Z(n12794) );
  NAND U13365 ( .A(n182), .B(n12794), .Z(n12666) );
  AND U13366 ( .A(n12667), .B(n12666), .Z(n12801) );
  NAND U13367 ( .A(n189), .B(n12668), .Z(n12670) );
  XOR U13368 ( .A(b[17]), .B(a[84]), .Z(n12797) );
  NAND U13369 ( .A(n37652), .B(n12797), .Z(n12669) );
  NAND U13370 ( .A(n12670), .B(n12669), .Z(n12800) );
  XNOR U13371 ( .A(n12801), .B(n12800), .Z(n12802) );
  XOR U13372 ( .A(n12803), .B(n12802), .Z(n12837) );
  XOR U13373 ( .A(n12836), .B(n12837), .Z(n12839) );
  XOR U13374 ( .A(n12838), .B(n12839), .Z(n12885) );
  NANDN U13375 ( .A(n12672), .B(n12671), .Z(n12676) );
  NANDN U13376 ( .A(n12674), .B(n12673), .Z(n12675) );
  AND U13377 ( .A(n12676), .B(n12675), .Z(n12824) );
  NANDN U13378 ( .A(n12678), .B(n12677), .Z(n12682) );
  NANDN U13379 ( .A(n12680), .B(n12679), .Z(n12681) );
  NAND U13380 ( .A(n12682), .B(n12681), .Z(n12825) );
  XNOR U13381 ( .A(n12824), .B(n12825), .Z(n12826) );
  NANDN U13382 ( .A(n12684), .B(n12683), .Z(n12688) );
  NAND U13383 ( .A(n12686), .B(n12685), .Z(n12687) );
  NAND U13384 ( .A(n12688), .B(n12687), .Z(n12827) );
  XNOR U13385 ( .A(n12826), .B(n12827), .Z(n12884) );
  XNOR U13386 ( .A(n12885), .B(n12884), .Z(n12887) );
  NAND U13387 ( .A(n12690), .B(n12689), .Z(n12694) );
  NAND U13388 ( .A(n12692), .B(n12691), .Z(n12693) );
  AND U13389 ( .A(n12694), .B(n12693), .Z(n12886) );
  XOR U13390 ( .A(n12887), .B(n12886), .Z(n12899) );
  NANDN U13391 ( .A(n12696), .B(n12695), .Z(n12700) );
  NANDN U13392 ( .A(n12698), .B(n12697), .Z(n12699) );
  AND U13393 ( .A(n12700), .B(n12699), .Z(n12896) );
  NANDN U13394 ( .A(n12706), .B(n12705), .Z(n12710) );
  OR U13395 ( .A(n12708), .B(n12707), .Z(n12709) );
  AND U13396 ( .A(n12710), .B(n12709), .Z(n12891) );
  NANDN U13397 ( .A(n12712), .B(n12711), .Z(n12716) );
  NANDN U13398 ( .A(n12714), .B(n12713), .Z(n12715) );
  AND U13399 ( .A(n12716), .B(n12715), .Z(n12831) );
  NANDN U13400 ( .A(n12718), .B(n12717), .Z(n12722) );
  OR U13401 ( .A(n12720), .B(n12719), .Z(n12721) );
  NAND U13402 ( .A(n12722), .B(n12721), .Z(n12830) );
  XNOR U13403 ( .A(n12831), .B(n12830), .Z(n12832) );
  NAND U13404 ( .A(b[0]), .B(a[100]), .Z(n12723) );
  XNOR U13405 ( .A(b[1]), .B(n12723), .Z(n12725) );
  NANDN U13406 ( .A(b[0]), .B(a[99]), .Z(n12724) );
  NAND U13407 ( .A(n12725), .B(n12724), .Z(n12779) );
  NAND U13408 ( .A(n194), .B(n12726), .Z(n12728) );
  XOR U13409 ( .A(b[29]), .B(a[72]), .Z(n12857) );
  NAND U13410 ( .A(n38456), .B(n12857), .Z(n12727) );
  AND U13411 ( .A(n12728), .B(n12727), .Z(n12777) );
  AND U13412 ( .A(b[31]), .B(a[68]), .Z(n12776) );
  XNOR U13413 ( .A(n12777), .B(n12776), .Z(n12778) );
  XNOR U13414 ( .A(n12779), .B(n12778), .Z(n12818) );
  NAND U13415 ( .A(n38185), .B(n12729), .Z(n12731) );
  XOR U13416 ( .A(b[23]), .B(a[78]), .Z(n12860) );
  NAND U13417 ( .A(n38132), .B(n12860), .Z(n12730) );
  AND U13418 ( .A(n12731), .B(n12730), .Z(n12851) );
  NAND U13419 ( .A(n184), .B(n12732), .Z(n12734) );
  XOR U13420 ( .A(b[7]), .B(a[94]), .Z(n12863) );
  NAND U13421 ( .A(n36592), .B(n12863), .Z(n12733) );
  AND U13422 ( .A(n12734), .B(n12733), .Z(n12849) );
  NAND U13423 ( .A(n38289), .B(n12735), .Z(n12737) );
  XOR U13424 ( .A(b[25]), .B(a[76]), .Z(n12866) );
  NAND U13425 ( .A(n38247), .B(n12866), .Z(n12736) );
  NAND U13426 ( .A(n12737), .B(n12736), .Z(n12848) );
  XNOR U13427 ( .A(n12849), .B(n12848), .Z(n12850) );
  XOR U13428 ( .A(n12851), .B(n12850), .Z(n12819) );
  XNOR U13429 ( .A(n12818), .B(n12819), .Z(n12820) );
  NAND U13430 ( .A(n187), .B(n12738), .Z(n12740) );
  XOR U13431 ( .A(b[13]), .B(a[88]), .Z(n12869) );
  NAND U13432 ( .A(n37295), .B(n12869), .Z(n12739) );
  AND U13433 ( .A(n12740), .B(n12739), .Z(n12813) );
  NAND U13434 ( .A(n186), .B(n12741), .Z(n12743) );
  XOR U13435 ( .A(b[11]), .B(a[90]), .Z(n12872) );
  NAND U13436 ( .A(n37097), .B(n12872), .Z(n12742) );
  NAND U13437 ( .A(n12743), .B(n12742), .Z(n12812) );
  XNOR U13438 ( .A(n12813), .B(n12812), .Z(n12814) );
  NAND U13439 ( .A(n188), .B(n12744), .Z(n12746) );
  XOR U13440 ( .A(b[15]), .B(a[86]), .Z(n12875) );
  NAND U13441 ( .A(n37382), .B(n12875), .Z(n12745) );
  AND U13442 ( .A(n12746), .B(n12745), .Z(n12809) );
  NAND U13443 ( .A(n38064), .B(n12747), .Z(n12749) );
  XOR U13444 ( .A(b[21]), .B(a[80]), .Z(n12878) );
  NAND U13445 ( .A(n37993), .B(n12878), .Z(n12748) );
  AND U13446 ( .A(n12749), .B(n12748), .Z(n12807) );
  NAND U13447 ( .A(n185), .B(n12750), .Z(n12752) );
  XOR U13448 ( .A(b[9]), .B(a[92]), .Z(n12881) );
  NAND U13449 ( .A(n36805), .B(n12881), .Z(n12751) );
  NAND U13450 ( .A(n12752), .B(n12751), .Z(n12806) );
  XNOR U13451 ( .A(n12807), .B(n12806), .Z(n12808) );
  XOR U13452 ( .A(n12809), .B(n12808), .Z(n12815) );
  XOR U13453 ( .A(n12814), .B(n12815), .Z(n12821) );
  XOR U13454 ( .A(n12820), .B(n12821), .Z(n12833) );
  XNOR U13455 ( .A(n12832), .B(n12833), .Z(n12890) );
  XNOR U13456 ( .A(n12891), .B(n12890), .Z(n12892) );
  XOR U13457 ( .A(n12893), .B(n12892), .Z(n12897) );
  XNOR U13458 ( .A(n12896), .B(n12897), .Z(n12898) );
  XNOR U13459 ( .A(n12899), .B(n12898), .Z(n12904) );
  XOR U13460 ( .A(n12905), .B(n12904), .Z(n12771) );
  NANDN U13461 ( .A(n12754), .B(n12753), .Z(n12758) );
  NANDN U13462 ( .A(n12756), .B(n12755), .Z(n12757) );
  AND U13463 ( .A(n12758), .B(n12757), .Z(n12770) );
  XOR U13464 ( .A(n12771), .B(n12770), .Z(n12773) );
  XNOR U13465 ( .A(n12772), .B(n12773), .Z(n12764) );
  XNOR U13466 ( .A(n12765), .B(n12764), .Z(n12766) );
  XNOR U13467 ( .A(n12767), .B(n12766), .Z(n12908) );
  XNOR U13468 ( .A(sreg[324]), .B(n12908), .Z(n12910) );
  NANDN U13469 ( .A(sreg[323]), .B(n12759), .Z(n12763) );
  NAND U13470 ( .A(n12761), .B(n12760), .Z(n12762) );
  NAND U13471 ( .A(n12763), .B(n12762), .Z(n12909) );
  XNOR U13472 ( .A(n12910), .B(n12909), .Z(c[324]) );
  NANDN U13473 ( .A(n12765), .B(n12764), .Z(n12769) );
  NANDN U13474 ( .A(n12767), .B(n12766), .Z(n12768) );
  AND U13475 ( .A(n12769), .B(n12768), .Z(n12916) );
  NANDN U13476 ( .A(n12771), .B(n12770), .Z(n12775) );
  NANDN U13477 ( .A(n12773), .B(n12772), .Z(n12774) );
  AND U13478 ( .A(n12775), .B(n12774), .Z(n12914) );
  NANDN U13479 ( .A(n12777), .B(n12776), .Z(n12781) );
  NANDN U13480 ( .A(n12779), .B(n12778), .Z(n12780) );
  AND U13481 ( .A(n12781), .B(n12780), .Z(n13005) );
  NAND U13482 ( .A(n38385), .B(n12782), .Z(n12784) );
  XOR U13483 ( .A(b[27]), .B(a[75]), .Z(n12949) );
  NAND U13484 ( .A(n38343), .B(n12949), .Z(n12783) );
  AND U13485 ( .A(n12784), .B(n12783), .Z(n13012) );
  NAND U13486 ( .A(n183), .B(n12785), .Z(n12787) );
  XOR U13487 ( .A(b[5]), .B(a[97]), .Z(n12952) );
  NAND U13488 ( .A(n36296), .B(n12952), .Z(n12786) );
  AND U13489 ( .A(n12787), .B(n12786), .Z(n13010) );
  NAND U13490 ( .A(n190), .B(n12788), .Z(n12790) );
  XOR U13491 ( .A(b[19]), .B(a[83]), .Z(n12955) );
  NAND U13492 ( .A(n37821), .B(n12955), .Z(n12789) );
  NAND U13493 ( .A(n12790), .B(n12789), .Z(n13009) );
  XNOR U13494 ( .A(n13010), .B(n13009), .Z(n13011) );
  XNOR U13495 ( .A(n13012), .B(n13011), .Z(n13003) );
  NAND U13496 ( .A(n38470), .B(n12791), .Z(n12793) );
  XOR U13497 ( .A(b[31]), .B(a[71]), .Z(n12958) );
  NAND U13498 ( .A(n38453), .B(n12958), .Z(n12792) );
  AND U13499 ( .A(n12793), .B(n12792), .Z(n12970) );
  NAND U13500 ( .A(n181), .B(n12794), .Z(n12796) );
  XOR U13501 ( .A(b[3]), .B(a[99]), .Z(n12961) );
  NAND U13502 ( .A(n182), .B(n12961), .Z(n12795) );
  AND U13503 ( .A(n12796), .B(n12795), .Z(n12968) );
  NAND U13504 ( .A(n189), .B(n12797), .Z(n12799) );
  XOR U13505 ( .A(b[17]), .B(a[85]), .Z(n12964) );
  NAND U13506 ( .A(n37652), .B(n12964), .Z(n12798) );
  NAND U13507 ( .A(n12799), .B(n12798), .Z(n12967) );
  XNOR U13508 ( .A(n12968), .B(n12967), .Z(n12969) );
  XOR U13509 ( .A(n12970), .B(n12969), .Z(n13004) );
  XOR U13510 ( .A(n13003), .B(n13004), .Z(n13006) );
  XOR U13511 ( .A(n13005), .B(n13006), .Z(n12938) );
  NANDN U13512 ( .A(n12801), .B(n12800), .Z(n12805) );
  NANDN U13513 ( .A(n12803), .B(n12802), .Z(n12804) );
  AND U13514 ( .A(n12805), .B(n12804), .Z(n12991) );
  NANDN U13515 ( .A(n12807), .B(n12806), .Z(n12811) );
  NANDN U13516 ( .A(n12809), .B(n12808), .Z(n12810) );
  NAND U13517 ( .A(n12811), .B(n12810), .Z(n12992) );
  XNOR U13518 ( .A(n12991), .B(n12992), .Z(n12993) );
  NANDN U13519 ( .A(n12813), .B(n12812), .Z(n12817) );
  NANDN U13520 ( .A(n12815), .B(n12814), .Z(n12816) );
  NAND U13521 ( .A(n12817), .B(n12816), .Z(n12994) );
  XNOR U13522 ( .A(n12993), .B(n12994), .Z(n12937) );
  XNOR U13523 ( .A(n12938), .B(n12937), .Z(n12940) );
  NANDN U13524 ( .A(n12819), .B(n12818), .Z(n12823) );
  NANDN U13525 ( .A(n12821), .B(n12820), .Z(n12822) );
  AND U13526 ( .A(n12823), .B(n12822), .Z(n12939) );
  XOR U13527 ( .A(n12940), .B(n12939), .Z(n13053) );
  NANDN U13528 ( .A(n12825), .B(n12824), .Z(n12829) );
  NANDN U13529 ( .A(n12827), .B(n12826), .Z(n12828) );
  AND U13530 ( .A(n12829), .B(n12828), .Z(n13051) );
  NANDN U13531 ( .A(n12831), .B(n12830), .Z(n12835) );
  NANDN U13532 ( .A(n12833), .B(n12832), .Z(n12834) );
  AND U13533 ( .A(n12835), .B(n12834), .Z(n12934) );
  NANDN U13534 ( .A(n12837), .B(n12836), .Z(n12841) );
  OR U13535 ( .A(n12839), .B(n12838), .Z(n12840) );
  AND U13536 ( .A(n12841), .B(n12840), .Z(n12932) );
  NANDN U13537 ( .A(n12843), .B(n12842), .Z(n12847) );
  NANDN U13538 ( .A(n12845), .B(n12844), .Z(n12846) );
  AND U13539 ( .A(n12847), .B(n12846), .Z(n12998) );
  NANDN U13540 ( .A(n12849), .B(n12848), .Z(n12853) );
  NANDN U13541 ( .A(n12851), .B(n12850), .Z(n12852) );
  NAND U13542 ( .A(n12853), .B(n12852), .Z(n12997) );
  XNOR U13543 ( .A(n12998), .B(n12997), .Z(n12999) );
  NAND U13544 ( .A(b[0]), .B(a[101]), .Z(n12854) );
  XNOR U13545 ( .A(b[1]), .B(n12854), .Z(n12856) );
  NANDN U13546 ( .A(b[0]), .B(a[100]), .Z(n12855) );
  NAND U13547 ( .A(n12856), .B(n12855), .Z(n12946) );
  NAND U13548 ( .A(n194), .B(n12857), .Z(n12859) );
  XOR U13549 ( .A(b[29]), .B(a[73]), .Z(n13021) );
  NAND U13550 ( .A(n38456), .B(n13021), .Z(n12858) );
  AND U13551 ( .A(n12859), .B(n12858), .Z(n12944) );
  AND U13552 ( .A(b[31]), .B(a[69]), .Z(n12943) );
  XNOR U13553 ( .A(n12944), .B(n12943), .Z(n12945) );
  XNOR U13554 ( .A(n12946), .B(n12945), .Z(n12985) );
  NAND U13555 ( .A(n38185), .B(n12860), .Z(n12862) );
  XOR U13556 ( .A(b[23]), .B(a[79]), .Z(n13027) );
  NAND U13557 ( .A(n38132), .B(n13027), .Z(n12861) );
  AND U13558 ( .A(n12862), .B(n12861), .Z(n13018) );
  NAND U13559 ( .A(n184), .B(n12863), .Z(n12865) );
  XOR U13560 ( .A(b[7]), .B(a[95]), .Z(n13030) );
  NAND U13561 ( .A(n36592), .B(n13030), .Z(n12864) );
  AND U13562 ( .A(n12865), .B(n12864), .Z(n13016) );
  NAND U13563 ( .A(n38289), .B(n12866), .Z(n12868) );
  XOR U13564 ( .A(b[25]), .B(a[77]), .Z(n13033) );
  NAND U13565 ( .A(n38247), .B(n13033), .Z(n12867) );
  NAND U13566 ( .A(n12868), .B(n12867), .Z(n13015) );
  XNOR U13567 ( .A(n13016), .B(n13015), .Z(n13017) );
  XOR U13568 ( .A(n13018), .B(n13017), .Z(n12986) );
  XNOR U13569 ( .A(n12985), .B(n12986), .Z(n12987) );
  NAND U13570 ( .A(n187), .B(n12869), .Z(n12871) );
  XOR U13571 ( .A(b[13]), .B(a[89]), .Z(n13036) );
  NAND U13572 ( .A(n37295), .B(n13036), .Z(n12870) );
  AND U13573 ( .A(n12871), .B(n12870), .Z(n12980) );
  NAND U13574 ( .A(n186), .B(n12872), .Z(n12874) );
  XOR U13575 ( .A(b[11]), .B(a[91]), .Z(n13039) );
  NAND U13576 ( .A(n37097), .B(n13039), .Z(n12873) );
  NAND U13577 ( .A(n12874), .B(n12873), .Z(n12979) );
  XNOR U13578 ( .A(n12980), .B(n12979), .Z(n12981) );
  NAND U13579 ( .A(n188), .B(n12875), .Z(n12877) );
  XOR U13580 ( .A(b[15]), .B(a[87]), .Z(n13042) );
  NAND U13581 ( .A(n37382), .B(n13042), .Z(n12876) );
  AND U13582 ( .A(n12877), .B(n12876), .Z(n12976) );
  NAND U13583 ( .A(n38064), .B(n12878), .Z(n12880) );
  XOR U13584 ( .A(b[21]), .B(a[81]), .Z(n13045) );
  NAND U13585 ( .A(n37993), .B(n13045), .Z(n12879) );
  AND U13586 ( .A(n12880), .B(n12879), .Z(n12974) );
  NAND U13587 ( .A(n185), .B(n12881), .Z(n12883) );
  XOR U13588 ( .A(b[9]), .B(a[93]), .Z(n13048) );
  NAND U13589 ( .A(n36805), .B(n13048), .Z(n12882) );
  NAND U13590 ( .A(n12883), .B(n12882), .Z(n12973) );
  XNOR U13591 ( .A(n12974), .B(n12973), .Z(n12975) );
  XOR U13592 ( .A(n12976), .B(n12975), .Z(n12982) );
  XOR U13593 ( .A(n12981), .B(n12982), .Z(n12988) );
  XOR U13594 ( .A(n12987), .B(n12988), .Z(n13000) );
  XNOR U13595 ( .A(n12999), .B(n13000), .Z(n12931) );
  XNOR U13596 ( .A(n12932), .B(n12931), .Z(n12933) );
  XOR U13597 ( .A(n12934), .B(n12933), .Z(n13052) );
  XOR U13598 ( .A(n13051), .B(n13052), .Z(n13054) );
  XOR U13599 ( .A(n13053), .B(n13054), .Z(n12928) );
  NANDN U13600 ( .A(n12885), .B(n12884), .Z(n12889) );
  NAND U13601 ( .A(n12887), .B(n12886), .Z(n12888) );
  AND U13602 ( .A(n12889), .B(n12888), .Z(n12926) );
  NANDN U13603 ( .A(n12891), .B(n12890), .Z(n12895) );
  NANDN U13604 ( .A(n12893), .B(n12892), .Z(n12894) );
  AND U13605 ( .A(n12895), .B(n12894), .Z(n12925) );
  XNOR U13606 ( .A(n12926), .B(n12925), .Z(n12927) );
  XNOR U13607 ( .A(n12928), .B(n12927), .Z(n12919) );
  NANDN U13608 ( .A(n12897), .B(n12896), .Z(n12901) );
  NANDN U13609 ( .A(n12899), .B(n12898), .Z(n12900) );
  NAND U13610 ( .A(n12901), .B(n12900), .Z(n12920) );
  XNOR U13611 ( .A(n12919), .B(n12920), .Z(n12921) );
  NANDN U13612 ( .A(n12903), .B(n12902), .Z(n12907) );
  NAND U13613 ( .A(n12905), .B(n12904), .Z(n12906) );
  NAND U13614 ( .A(n12907), .B(n12906), .Z(n12922) );
  XNOR U13615 ( .A(n12921), .B(n12922), .Z(n12913) );
  XNOR U13616 ( .A(n12914), .B(n12913), .Z(n12915) );
  XNOR U13617 ( .A(n12916), .B(n12915), .Z(n13057) );
  XNOR U13618 ( .A(sreg[325]), .B(n13057), .Z(n13059) );
  NANDN U13619 ( .A(sreg[324]), .B(n12908), .Z(n12912) );
  NAND U13620 ( .A(n12910), .B(n12909), .Z(n12911) );
  NAND U13621 ( .A(n12912), .B(n12911), .Z(n13058) );
  XNOR U13622 ( .A(n13059), .B(n13058), .Z(c[325]) );
  NANDN U13623 ( .A(n12914), .B(n12913), .Z(n12918) );
  NANDN U13624 ( .A(n12916), .B(n12915), .Z(n12917) );
  AND U13625 ( .A(n12918), .B(n12917), .Z(n13065) );
  NANDN U13626 ( .A(n12920), .B(n12919), .Z(n12924) );
  NANDN U13627 ( .A(n12922), .B(n12921), .Z(n12923) );
  AND U13628 ( .A(n12924), .B(n12923), .Z(n13063) );
  NANDN U13629 ( .A(n12926), .B(n12925), .Z(n12930) );
  NANDN U13630 ( .A(n12928), .B(n12927), .Z(n12929) );
  AND U13631 ( .A(n12930), .B(n12929), .Z(n13071) );
  NANDN U13632 ( .A(n12932), .B(n12931), .Z(n12936) );
  NANDN U13633 ( .A(n12934), .B(n12933), .Z(n12935) );
  AND U13634 ( .A(n12936), .B(n12935), .Z(n13075) );
  NANDN U13635 ( .A(n12938), .B(n12937), .Z(n12942) );
  NAND U13636 ( .A(n12940), .B(n12939), .Z(n12941) );
  AND U13637 ( .A(n12942), .B(n12941), .Z(n13074) );
  XNOR U13638 ( .A(n13075), .B(n13074), .Z(n13077) );
  NANDN U13639 ( .A(n12944), .B(n12943), .Z(n12948) );
  NANDN U13640 ( .A(n12946), .B(n12945), .Z(n12947) );
  AND U13641 ( .A(n12948), .B(n12947), .Z(n13154) );
  NAND U13642 ( .A(n38385), .B(n12949), .Z(n12951) );
  XOR U13643 ( .A(b[27]), .B(a[76]), .Z(n13098) );
  NAND U13644 ( .A(n38343), .B(n13098), .Z(n12950) );
  AND U13645 ( .A(n12951), .B(n12950), .Z(n13161) );
  NAND U13646 ( .A(n183), .B(n12952), .Z(n12954) );
  XOR U13647 ( .A(b[5]), .B(a[98]), .Z(n13101) );
  NAND U13648 ( .A(n36296), .B(n13101), .Z(n12953) );
  AND U13649 ( .A(n12954), .B(n12953), .Z(n13159) );
  NAND U13650 ( .A(n190), .B(n12955), .Z(n12957) );
  XOR U13651 ( .A(b[19]), .B(a[84]), .Z(n13104) );
  NAND U13652 ( .A(n37821), .B(n13104), .Z(n12956) );
  NAND U13653 ( .A(n12957), .B(n12956), .Z(n13158) );
  XNOR U13654 ( .A(n13159), .B(n13158), .Z(n13160) );
  XNOR U13655 ( .A(n13161), .B(n13160), .Z(n13152) );
  NAND U13656 ( .A(n38470), .B(n12958), .Z(n12960) );
  XOR U13657 ( .A(b[31]), .B(a[72]), .Z(n13107) );
  NAND U13658 ( .A(n38453), .B(n13107), .Z(n12959) );
  AND U13659 ( .A(n12960), .B(n12959), .Z(n13119) );
  NAND U13660 ( .A(n181), .B(n12961), .Z(n12963) );
  XOR U13661 ( .A(b[3]), .B(a[100]), .Z(n13110) );
  NAND U13662 ( .A(n182), .B(n13110), .Z(n12962) );
  AND U13663 ( .A(n12963), .B(n12962), .Z(n13117) );
  NAND U13664 ( .A(n189), .B(n12964), .Z(n12966) );
  XOR U13665 ( .A(b[17]), .B(a[86]), .Z(n13113) );
  NAND U13666 ( .A(n37652), .B(n13113), .Z(n12965) );
  NAND U13667 ( .A(n12966), .B(n12965), .Z(n13116) );
  XNOR U13668 ( .A(n13117), .B(n13116), .Z(n13118) );
  XOR U13669 ( .A(n13119), .B(n13118), .Z(n13153) );
  XOR U13670 ( .A(n13152), .B(n13153), .Z(n13155) );
  XOR U13671 ( .A(n13154), .B(n13155), .Z(n13087) );
  NANDN U13672 ( .A(n12968), .B(n12967), .Z(n12972) );
  NANDN U13673 ( .A(n12970), .B(n12969), .Z(n12971) );
  AND U13674 ( .A(n12972), .B(n12971), .Z(n13140) );
  NANDN U13675 ( .A(n12974), .B(n12973), .Z(n12978) );
  NANDN U13676 ( .A(n12976), .B(n12975), .Z(n12977) );
  NAND U13677 ( .A(n12978), .B(n12977), .Z(n13141) );
  XNOR U13678 ( .A(n13140), .B(n13141), .Z(n13142) );
  NANDN U13679 ( .A(n12980), .B(n12979), .Z(n12984) );
  NANDN U13680 ( .A(n12982), .B(n12981), .Z(n12983) );
  NAND U13681 ( .A(n12984), .B(n12983), .Z(n13143) );
  XNOR U13682 ( .A(n13142), .B(n13143), .Z(n13086) );
  XNOR U13683 ( .A(n13087), .B(n13086), .Z(n13089) );
  NANDN U13684 ( .A(n12986), .B(n12985), .Z(n12990) );
  NANDN U13685 ( .A(n12988), .B(n12987), .Z(n12989) );
  AND U13686 ( .A(n12990), .B(n12989), .Z(n13088) );
  XOR U13687 ( .A(n13089), .B(n13088), .Z(n13203) );
  NANDN U13688 ( .A(n12992), .B(n12991), .Z(n12996) );
  NANDN U13689 ( .A(n12994), .B(n12993), .Z(n12995) );
  AND U13690 ( .A(n12996), .B(n12995), .Z(n13200) );
  NANDN U13691 ( .A(n12998), .B(n12997), .Z(n13002) );
  NANDN U13692 ( .A(n13000), .B(n12999), .Z(n13001) );
  AND U13693 ( .A(n13002), .B(n13001), .Z(n13083) );
  NANDN U13694 ( .A(n13004), .B(n13003), .Z(n13008) );
  OR U13695 ( .A(n13006), .B(n13005), .Z(n13007) );
  AND U13696 ( .A(n13008), .B(n13007), .Z(n13081) );
  NANDN U13697 ( .A(n13010), .B(n13009), .Z(n13014) );
  NANDN U13698 ( .A(n13012), .B(n13011), .Z(n13013) );
  AND U13699 ( .A(n13014), .B(n13013), .Z(n13147) );
  NANDN U13700 ( .A(n13016), .B(n13015), .Z(n13020) );
  NANDN U13701 ( .A(n13018), .B(n13017), .Z(n13019) );
  NAND U13702 ( .A(n13020), .B(n13019), .Z(n13146) );
  XNOR U13703 ( .A(n13147), .B(n13146), .Z(n13148) );
  NAND U13704 ( .A(n194), .B(n13021), .Z(n13023) );
  XOR U13705 ( .A(b[29]), .B(a[74]), .Z(n13173) );
  NAND U13706 ( .A(n38456), .B(n13173), .Z(n13022) );
  AND U13707 ( .A(n13023), .B(n13022), .Z(n13093) );
  AND U13708 ( .A(b[31]), .B(a[70]), .Z(n13092) );
  XNOR U13709 ( .A(n13093), .B(n13092), .Z(n13094) );
  NAND U13710 ( .A(b[0]), .B(a[102]), .Z(n13024) );
  XNOR U13711 ( .A(b[1]), .B(n13024), .Z(n13026) );
  NANDN U13712 ( .A(b[0]), .B(a[101]), .Z(n13025) );
  NAND U13713 ( .A(n13026), .B(n13025), .Z(n13095) );
  XNOR U13714 ( .A(n13094), .B(n13095), .Z(n13134) );
  NAND U13715 ( .A(n38185), .B(n13027), .Z(n13029) );
  XOR U13716 ( .A(b[23]), .B(a[80]), .Z(n13176) );
  NAND U13717 ( .A(n38132), .B(n13176), .Z(n13028) );
  AND U13718 ( .A(n13029), .B(n13028), .Z(n13167) );
  NAND U13719 ( .A(n184), .B(n13030), .Z(n13032) );
  XOR U13720 ( .A(b[7]), .B(a[96]), .Z(n13179) );
  NAND U13721 ( .A(n36592), .B(n13179), .Z(n13031) );
  AND U13722 ( .A(n13032), .B(n13031), .Z(n13165) );
  NAND U13723 ( .A(n38289), .B(n13033), .Z(n13035) );
  XOR U13724 ( .A(b[25]), .B(a[78]), .Z(n13182) );
  NAND U13725 ( .A(n38247), .B(n13182), .Z(n13034) );
  NAND U13726 ( .A(n13035), .B(n13034), .Z(n13164) );
  XNOR U13727 ( .A(n13165), .B(n13164), .Z(n13166) );
  XOR U13728 ( .A(n13167), .B(n13166), .Z(n13135) );
  XNOR U13729 ( .A(n13134), .B(n13135), .Z(n13136) );
  NAND U13730 ( .A(n187), .B(n13036), .Z(n13038) );
  XOR U13731 ( .A(b[13]), .B(a[90]), .Z(n13185) );
  NAND U13732 ( .A(n37295), .B(n13185), .Z(n13037) );
  AND U13733 ( .A(n13038), .B(n13037), .Z(n13129) );
  NAND U13734 ( .A(n186), .B(n13039), .Z(n13041) );
  XOR U13735 ( .A(b[11]), .B(a[92]), .Z(n13188) );
  NAND U13736 ( .A(n37097), .B(n13188), .Z(n13040) );
  NAND U13737 ( .A(n13041), .B(n13040), .Z(n13128) );
  XNOR U13738 ( .A(n13129), .B(n13128), .Z(n13130) );
  NAND U13739 ( .A(n188), .B(n13042), .Z(n13044) );
  XOR U13740 ( .A(b[15]), .B(a[88]), .Z(n13191) );
  NAND U13741 ( .A(n37382), .B(n13191), .Z(n13043) );
  AND U13742 ( .A(n13044), .B(n13043), .Z(n13125) );
  NAND U13743 ( .A(n38064), .B(n13045), .Z(n13047) );
  XOR U13744 ( .A(b[21]), .B(a[82]), .Z(n13194) );
  NAND U13745 ( .A(n37993), .B(n13194), .Z(n13046) );
  AND U13746 ( .A(n13047), .B(n13046), .Z(n13123) );
  NAND U13747 ( .A(n185), .B(n13048), .Z(n13050) );
  XOR U13748 ( .A(b[9]), .B(a[94]), .Z(n13197) );
  NAND U13749 ( .A(n36805), .B(n13197), .Z(n13049) );
  NAND U13750 ( .A(n13050), .B(n13049), .Z(n13122) );
  XNOR U13751 ( .A(n13123), .B(n13122), .Z(n13124) );
  XOR U13752 ( .A(n13125), .B(n13124), .Z(n13131) );
  XOR U13753 ( .A(n13130), .B(n13131), .Z(n13137) );
  XOR U13754 ( .A(n13136), .B(n13137), .Z(n13149) );
  XNOR U13755 ( .A(n13148), .B(n13149), .Z(n13080) );
  XNOR U13756 ( .A(n13081), .B(n13080), .Z(n13082) );
  XOR U13757 ( .A(n13083), .B(n13082), .Z(n13201) );
  XNOR U13758 ( .A(n13200), .B(n13201), .Z(n13202) );
  XNOR U13759 ( .A(n13203), .B(n13202), .Z(n13076) );
  XOR U13760 ( .A(n13077), .B(n13076), .Z(n13069) );
  NANDN U13761 ( .A(n13052), .B(n13051), .Z(n13056) );
  OR U13762 ( .A(n13054), .B(n13053), .Z(n13055) );
  AND U13763 ( .A(n13056), .B(n13055), .Z(n13068) );
  XNOR U13764 ( .A(n13069), .B(n13068), .Z(n13070) );
  XNOR U13765 ( .A(n13071), .B(n13070), .Z(n13062) );
  XNOR U13766 ( .A(n13063), .B(n13062), .Z(n13064) );
  XNOR U13767 ( .A(n13065), .B(n13064), .Z(n13206) );
  XNOR U13768 ( .A(sreg[326]), .B(n13206), .Z(n13208) );
  NANDN U13769 ( .A(sreg[325]), .B(n13057), .Z(n13061) );
  NAND U13770 ( .A(n13059), .B(n13058), .Z(n13060) );
  NAND U13771 ( .A(n13061), .B(n13060), .Z(n13207) );
  XNOR U13772 ( .A(n13208), .B(n13207), .Z(c[326]) );
  NANDN U13773 ( .A(n13063), .B(n13062), .Z(n13067) );
  NANDN U13774 ( .A(n13065), .B(n13064), .Z(n13066) );
  AND U13775 ( .A(n13067), .B(n13066), .Z(n13214) );
  NANDN U13776 ( .A(n13069), .B(n13068), .Z(n13073) );
  NANDN U13777 ( .A(n13071), .B(n13070), .Z(n13072) );
  AND U13778 ( .A(n13073), .B(n13072), .Z(n13212) );
  NANDN U13779 ( .A(n13075), .B(n13074), .Z(n13079) );
  NAND U13780 ( .A(n13077), .B(n13076), .Z(n13078) );
  AND U13781 ( .A(n13079), .B(n13078), .Z(n13219) );
  NANDN U13782 ( .A(n13081), .B(n13080), .Z(n13085) );
  NANDN U13783 ( .A(n13083), .B(n13082), .Z(n13084) );
  AND U13784 ( .A(n13085), .B(n13084), .Z(n13350) );
  NANDN U13785 ( .A(n13087), .B(n13086), .Z(n13091) );
  NAND U13786 ( .A(n13089), .B(n13088), .Z(n13090) );
  AND U13787 ( .A(n13091), .B(n13090), .Z(n13349) );
  XNOR U13788 ( .A(n13350), .B(n13349), .Z(n13352) );
  NANDN U13789 ( .A(n13093), .B(n13092), .Z(n13097) );
  NANDN U13790 ( .A(n13095), .B(n13094), .Z(n13096) );
  AND U13791 ( .A(n13097), .B(n13096), .Z(n13297) );
  NAND U13792 ( .A(n38385), .B(n13098), .Z(n13100) );
  XOR U13793 ( .A(b[27]), .B(a[77]), .Z(n13241) );
  NAND U13794 ( .A(n38343), .B(n13241), .Z(n13099) );
  AND U13795 ( .A(n13100), .B(n13099), .Z(n13304) );
  NAND U13796 ( .A(n183), .B(n13101), .Z(n13103) );
  XOR U13797 ( .A(b[5]), .B(a[99]), .Z(n13244) );
  NAND U13798 ( .A(n36296), .B(n13244), .Z(n13102) );
  AND U13799 ( .A(n13103), .B(n13102), .Z(n13302) );
  NAND U13800 ( .A(n190), .B(n13104), .Z(n13106) );
  XOR U13801 ( .A(b[19]), .B(a[85]), .Z(n13247) );
  NAND U13802 ( .A(n37821), .B(n13247), .Z(n13105) );
  NAND U13803 ( .A(n13106), .B(n13105), .Z(n13301) );
  XNOR U13804 ( .A(n13302), .B(n13301), .Z(n13303) );
  XNOR U13805 ( .A(n13304), .B(n13303), .Z(n13295) );
  NAND U13806 ( .A(n38470), .B(n13107), .Z(n13109) );
  XOR U13807 ( .A(b[31]), .B(a[73]), .Z(n13250) );
  NAND U13808 ( .A(n38453), .B(n13250), .Z(n13108) );
  AND U13809 ( .A(n13109), .B(n13108), .Z(n13262) );
  NAND U13810 ( .A(n181), .B(n13110), .Z(n13112) );
  XOR U13811 ( .A(b[3]), .B(a[101]), .Z(n13253) );
  NAND U13812 ( .A(n182), .B(n13253), .Z(n13111) );
  AND U13813 ( .A(n13112), .B(n13111), .Z(n13260) );
  NAND U13814 ( .A(n189), .B(n13113), .Z(n13115) );
  XOR U13815 ( .A(b[17]), .B(a[87]), .Z(n13256) );
  NAND U13816 ( .A(n37652), .B(n13256), .Z(n13114) );
  NAND U13817 ( .A(n13115), .B(n13114), .Z(n13259) );
  XNOR U13818 ( .A(n13260), .B(n13259), .Z(n13261) );
  XOR U13819 ( .A(n13262), .B(n13261), .Z(n13296) );
  XOR U13820 ( .A(n13295), .B(n13296), .Z(n13298) );
  XOR U13821 ( .A(n13297), .B(n13298), .Z(n13230) );
  NANDN U13822 ( .A(n13117), .B(n13116), .Z(n13121) );
  NANDN U13823 ( .A(n13119), .B(n13118), .Z(n13120) );
  AND U13824 ( .A(n13121), .B(n13120), .Z(n13283) );
  NANDN U13825 ( .A(n13123), .B(n13122), .Z(n13127) );
  NANDN U13826 ( .A(n13125), .B(n13124), .Z(n13126) );
  NAND U13827 ( .A(n13127), .B(n13126), .Z(n13284) );
  XNOR U13828 ( .A(n13283), .B(n13284), .Z(n13285) );
  NANDN U13829 ( .A(n13129), .B(n13128), .Z(n13133) );
  NANDN U13830 ( .A(n13131), .B(n13130), .Z(n13132) );
  NAND U13831 ( .A(n13133), .B(n13132), .Z(n13286) );
  XNOR U13832 ( .A(n13285), .B(n13286), .Z(n13229) );
  XNOR U13833 ( .A(n13230), .B(n13229), .Z(n13232) );
  NANDN U13834 ( .A(n13135), .B(n13134), .Z(n13139) );
  NANDN U13835 ( .A(n13137), .B(n13136), .Z(n13138) );
  AND U13836 ( .A(n13139), .B(n13138), .Z(n13231) );
  XOR U13837 ( .A(n13232), .B(n13231), .Z(n13346) );
  NANDN U13838 ( .A(n13141), .B(n13140), .Z(n13145) );
  NANDN U13839 ( .A(n13143), .B(n13142), .Z(n13144) );
  AND U13840 ( .A(n13145), .B(n13144), .Z(n13343) );
  NANDN U13841 ( .A(n13147), .B(n13146), .Z(n13151) );
  NANDN U13842 ( .A(n13149), .B(n13148), .Z(n13150) );
  AND U13843 ( .A(n13151), .B(n13150), .Z(n13226) );
  NANDN U13844 ( .A(n13153), .B(n13152), .Z(n13157) );
  OR U13845 ( .A(n13155), .B(n13154), .Z(n13156) );
  AND U13846 ( .A(n13157), .B(n13156), .Z(n13224) );
  NANDN U13847 ( .A(n13159), .B(n13158), .Z(n13163) );
  NANDN U13848 ( .A(n13161), .B(n13160), .Z(n13162) );
  AND U13849 ( .A(n13163), .B(n13162), .Z(n13290) );
  NANDN U13850 ( .A(n13165), .B(n13164), .Z(n13169) );
  NANDN U13851 ( .A(n13167), .B(n13166), .Z(n13168) );
  NAND U13852 ( .A(n13169), .B(n13168), .Z(n13289) );
  XNOR U13853 ( .A(n13290), .B(n13289), .Z(n13291) );
  NAND U13854 ( .A(b[0]), .B(a[103]), .Z(n13170) );
  XNOR U13855 ( .A(b[1]), .B(n13170), .Z(n13172) );
  NANDN U13856 ( .A(b[0]), .B(a[102]), .Z(n13171) );
  NAND U13857 ( .A(n13172), .B(n13171), .Z(n13238) );
  NAND U13858 ( .A(n194), .B(n13173), .Z(n13175) );
  XOR U13859 ( .A(b[29]), .B(a[75]), .Z(n13313) );
  NAND U13860 ( .A(n38456), .B(n13313), .Z(n13174) );
  AND U13861 ( .A(n13175), .B(n13174), .Z(n13236) );
  AND U13862 ( .A(b[31]), .B(a[71]), .Z(n13235) );
  XNOR U13863 ( .A(n13236), .B(n13235), .Z(n13237) );
  XNOR U13864 ( .A(n13238), .B(n13237), .Z(n13277) );
  NAND U13865 ( .A(n38185), .B(n13176), .Z(n13178) );
  XOR U13866 ( .A(b[23]), .B(a[81]), .Z(n13319) );
  NAND U13867 ( .A(n38132), .B(n13319), .Z(n13177) );
  AND U13868 ( .A(n13178), .B(n13177), .Z(n13310) );
  NAND U13869 ( .A(n184), .B(n13179), .Z(n13181) );
  XOR U13870 ( .A(b[7]), .B(a[97]), .Z(n13322) );
  NAND U13871 ( .A(n36592), .B(n13322), .Z(n13180) );
  AND U13872 ( .A(n13181), .B(n13180), .Z(n13308) );
  NAND U13873 ( .A(n38289), .B(n13182), .Z(n13184) );
  XOR U13874 ( .A(b[25]), .B(a[79]), .Z(n13325) );
  NAND U13875 ( .A(n38247), .B(n13325), .Z(n13183) );
  NAND U13876 ( .A(n13184), .B(n13183), .Z(n13307) );
  XNOR U13877 ( .A(n13308), .B(n13307), .Z(n13309) );
  XOR U13878 ( .A(n13310), .B(n13309), .Z(n13278) );
  XNOR U13879 ( .A(n13277), .B(n13278), .Z(n13279) );
  NAND U13880 ( .A(n187), .B(n13185), .Z(n13187) );
  XOR U13881 ( .A(b[13]), .B(a[91]), .Z(n13328) );
  NAND U13882 ( .A(n37295), .B(n13328), .Z(n13186) );
  AND U13883 ( .A(n13187), .B(n13186), .Z(n13272) );
  NAND U13884 ( .A(n186), .B(n13188), .Z(n13190) );
  XOR U13885 ( .A(b[11]), .B(a[93]), .Z(n13331) );
  NAND U13886 ( .A(n37097), .B(n13331), .Z(n13189) );
  NAND U13887 ( .A(n13190), .B(n13189), .Z(n13271) );
  XNOR U13888 ( .A(n13272), .B(n13271), .Z(n13273) );
  NAND U13889 ( .A(n188), .B(n13191), .Z(n13193) );
  XOR U13890 ( .A(b[15]), .B(a[89]), .Z(n13334) );
  NAND U13891 ( .A(n37382), .B(n13334), .Z(n13192) );
  AND U13892 ( .A(n13193), .B(n13192), .Z(n13268) );
  NAND U13893 ( .A(n38064), .B(n13194), .Z(n13196) );
  XOR U13894 ( .A(b[21]), .B(a[83]), .Z(n13337) );
  NAND U13895 ( .A(n37993), .B(n13337), .Z(n13195) );
  AND U13896 ( .A(n13196), .B(n13195), .Z(n13266) );
  NAND U13897 ( .A(n185), .B(n13197), .Z(n13199) );
  XOR U13898 ( .A(b[9]), .B(a[95]), .Z(n13340) );
  NAND U13899 ( .A(n36805), .B(n13340), .Z(n13198) );
  NAND U13900 ( .A(n13199), .B(n13198), .Z(n13265) );
  XNOR U13901 ( .A(n13266), .B(n13265), .Z(n13267) );
  XOR U13902 ( .A(n13268), .B(n13267), .Z(n13274) );
  XOR U13903 ( .A(n13273), .B(n13274), .Z(n13280) );
  XOR U13904 ( .A(n13279), .B(n13280), .Z(n13292) );
  XNOR U13905 ( .A(n13291), .B(n13292), .Z(n13223) );
  XNOR U13906 ( .A(n13224), .B(n13223), .Z(n13225) );
  XOR U13907 ( .A(n13226), .B(n13225), .Z(n13344) );
  XNOR U13908 ( .A(n13343), .B(n13344), .Z(n13345) );
  XNOR U13909 ( .A(n13346), .B(n13345), .Z(n13351) );
  XOR U13910 ( .A(n13352), .B(n13351), .Z(n13218) );
  NANDN U13911 ( .A(n13201), .B(n13200), .Z(n13205) );
  NANDN U13912 ( .A(n13203), .B(n13202), .Z(n13204) );
  AND U13913 ( .A(n13205), .B(n13204), .Z(n13217) );
  XOR U13914 ( .A(n13218), .B(n13217), .Z(n13220) );
  XNOR U13915 ( .A(n13219), .B(n13220), .Z(n13211) );
  XNOR U13916 ( .A(n13212), .B(n13211), .Z(n13213) );
  XNOR U13917 ( .A(n13214), .B(n13213), .Z(n13355) );
  XNOR U13918 ( .A(sreg[327]), .B(n13355), .Z(n13357) );
  NANDN U13919 ( .A(sreg[326]), .B(n13206), .Z(n13210) );
  NAND U13920 ( .A(n13208), .B(n13207), .Z(n13209) );
  NAND U13921 ( .A(n13210), .B(n13209), .Z(n13356) );
  XNOR U13922 ( .A(n13357), .B(n13356), .Z(c[327]) );
  NANDN U13923 ( .A(n13212), .B(n13211), .Z(n13216) );
  NANDN U13924 ( .A(n13214), .B(n13213), .Z(n13215) );
  AND U13925 ( .A(n13216), .B(n13215), .Z(n13363) );
  NANDN U13926 ( .A(n13218), .B(n13217), .Z(n13222) );
  NANDN U13927 ( .A(n13220), .B(n13219), .Z(n13221) );
  AND U13928 ( .A(n13222), .B(n13221), .Z(n13361) );
  NANDN U13929 ( .A(n13224), .B(n13223), .Z(n13228) );
  NANDN U13930 ( .A(n13226), .B(n13225), .Z(n13227) );
  AND U13931 ( .A(n13228), .B(n13227), .Z(n13499) );
  NANDN U13932 ( .A(n13230), .B(n13229), .Z(n13234) );
  NAND U13933 ( .A(n13232), .B(n13231), .Z(n13233) );
  AND U13934 ( .A(n13234), .B(n13233), .Z(n13498) );
  XNOR U13935 ( .A(n13499), .B(n13498), .Z(n13501) );
  NANDN U13936 ( .A(n13236), .B(n13235), .Z(n13240) );
  NANDN U13937 ( .A(n13238), .B(n13237), .Z(n13239) );
  AND U13938 ( .A(n13240), .B(n13239), .Z(n13446) );
  NAND U13939 ( .A(n38385), .B(n13241), .Z(n13243) );
  XOR U13940 ( .A(b[27]), .B(a[78]), .Z(n13390) );
  NAND U13941 ( .A(n38343), .B(n13390), .Z(n13242) );
  AND U13942 ( .A(n13243), .B(n13242), .Z(n13453) );
  NAND U13943 ( .A(n183), .B(n13244), .Z(n13246) );
  XOR U13944 ( .A(b[5]), .B(a[100]), .Z(n13393) );
  NAND U13945 ( .A(n36296), .B(n13393), .Z(n13245) );
  AND U13946 ( .A(n13246), .B(n13245), .Z(n13451) );
  NAND U13947 ( .A(n190), .B(n13247), .Z(n13249) );
  XOR U13948 ( .A(b[19]), .B(a[86]), .Z(n13396) );
  NAND U13949 ( .A(n37821), .B(n13396), .Z(n13248) );
  NAND U13950 ( .A(n13249), .B(n13248), .Z(n13450) );
  XNOR U13951 ( .A(n13451), .B(n13450), .Z(n13452) );
  XNOR U13952 ( .A(n13453), .B(n13452), .Z(n13444) );
  NAND U13953 ( .A(n38470), .B(n13250), .Z(n13252) );
  XOR U13954 ( .A(b[31]), .B(a[74]), .Z(n13399) );
  NAND U13955 ( .A(n38453), .B(n13399), .Z(n13251) );
  AND U13956 ( .A(n13252), .B(n13251), .Z(n13411) );
  NAND U13957 ( .A(n181), .B(n13253), .Z(n13255) );
  XOR U13958 ( .A(b[3]), .B(a[102]), .Z(n13402) );
  NAND U13959 ( .A(n182), .B(n13402), .Z(n13254) );
  AND U13960 ( .A(n13255), .B(n13254), .Z(n13409) );
  NAND U13961 ( .A(n189), .B(n13256), .Z(n13258) );
  XOR U13962 ( .A(b[17]), .B(a[88]), .Z(n13405) );
  NAND U13963 ( .A(n37652), .B(n13405), .Z(n13257) );
  NAND U13964 ( .A(n13258), .B(n13257), .Z(n13408) );
  XNOR U13965 ( .A(n13409), .B(n13408), .Z(n13410) );
  XOR U13966 ( .A(n13411), .B(n13410), .Z(n13445) );
  XOR U13967 ( .A(n13444), .B(n13445), .Z(n13447) );
  XOR U13968 ( .A(n13446), .B(n13447), .Z(n13379) );
  NANDN U13969 ( .A(n13260), .B(n13259), .Z(n13264) );
  NANDN U13970 ( .A(n13262), .B(n13261), .Z(n13263) );
  AND U13971 ( .A(n13264), .B(n13263), .Z(n13432) );
  NANDN U13972 ( .A(n13266), .B(n13265), .Z(n13270) );
  NANDN U13973 ( .A(n13268), .B(n13267), .Z(n13269) );
  NAND U13974 ( .A(n13270), .B(n13269), .Z(n13433) );
  XNOR U13975 ( .A(n13432), .B(n13433), .Z(n13434) );
  NANDN U13976 ( .A(n13272), .B(n13271), .Z(n13276) );
  NANDN U13977 ( .A(n13274), .B(n13273), .Z(n13275) );
  NAND U13978 ( .A(n13276), .B(n13275), .Z(n13435) );
  XNOR U13979 ( .A(n13434), .B(n13435), .Z(n13378) );
  XNOR U13980 ( .A(n13379), .B(n13378), .Z(n13381) );
  NANDN U13981 ( .A(n13278), .B(n13277), .Z(n13282) );
  NANDN U13982 ( .A(n13280), .B(n13279), .Z(n13281) );
  AND U13983 ( .A(n13282), .B(n13281), .Z(n13380) );
  XOR U13984 ( .A(n13381), .B(n13380), .Z(n13495) );
  NANDN U13985 ( .A(n13284), .B(n13283), .Z(n13288) );
  NANDN U13986 ( .A(n13286), .B(n13285), .Z(n13287) );
  AND U13987 ( .A(n13288), .B(n13287), .Z(n13492) );
  NANDN U13988 ( .A(n13290), .B(n13289), .Z(n13294) );
  NANDN U13989 ( .A(n13292), .B(n13291), .Z(n13293) );
  AND U13990 ( .A(n13294), .B(n13293), .Z(n13375) );
  NANDN U13991 ( .A(n13296), .B(n13295), .Z(n13300) );
  OR U13992 ( .A(n13298), .B(n13297), .Z(n13299) );
  AND U13993 ( .A(n13300), .B(n13299), .Z(n13373) );
  NANDN U13994 ( .A(n13302), .B(n13301), .Z(n13306) );
  NANDN U13995 ( .A(n13304), .B(n13303), .Z(n13305) );
  AND U13996 ( .A(n13306), .B(n13305), .Z(n13439) );
  NANDN U13997 ( .A(n13308), .B(n13307), .Z(n13312) );
  NANDN U13998 ( .A(n13310), .B(n13309), .Z(n13311) );
  NAND U13999 ( .A(n13312), .B(n13311), .Z(n13438) );
  XNOR U14000 ( .A(n13439), .B(n13438), .Z(n13440) );
  NAND U14001 ( .A(n194), .B(n13313), .Z(n13315) );
  XOR U14002 ( .A(b[29]), .B(a[76]), .Z(n13465) );
  NAND U14003 ( .A(n38456), .B(n13465), .Z(n13314) );
  AND U14004 ( .A(n13315), .B(n13314), .Z(n13385) );
  AND U14005 ( .A(b[31]), .B(a[72]), .Z(n13384) );
  XNOR U14006 ( .A(n13385), .B(n13384), .Z(n13386) );
  NAND U14007 ( .A(b[0]), .B(a[104]), .Z(n13316) );
  XNOR U14008 ( .A(b[1]), .B(n13316), .Z(n13318) );
  NANDN U14009 ( .A(b[0]), .B(a[103]), .Z(n13317) );
  NAND U14010 ( .A(n13318), .B(n13317), .Z(n13387) );
  XNOR U14011 ( .A(n13386), .B(n13387), .Z(n13426) );
  NAND U14012 ( .A(n38185), .B(n13319), .Z(n13321) );
  XOR U14013 ( .A(b[23]), .B(a[82]), .Z(n13468) );
  NAND U14014 ( .A(n38132), .B(n13468), .Z(n13320) );
  AND U14015 ( .A(n13321), .B(n13320), .Z(n13459) );
  NAND U14016 ( .A(n184), .B(n13322), .Z(n13324) );
  XOR U14017 ( .A(b[7]), .B(a[98]), .Z(n13471) );
  NAND U14018 ( .A(n36592), .B(n13471), .Z(n13323) );
  AND U14019 ( .A(n13324), .B(n13323), .Z(n13457) );
  NAND U14020 ( .A(n38289), .B(n13325), .Z(n13327) );
  XOR U14021 ( .A(b[25]), .B(a[80]), .Z(n13474) );
  NAND U14022 ( .A(n38247), .B(n13474), .Z(n13326) );
  NAND U14023 ( .A(n13327), .B(n13326), .Z(n13456) );
  XNOR U14024 ( .A(n13457), .B(n13456), .Z(n13458) );
  XOR U14025 ( .A(n13459), .B(n13458), .Z(n13427) );
  XNOR U14026 ( .A(n13426), .B(n13427), .Z(n13428) );
  NAND U14027 ( .A(n187), .B(n13328), .Z(n13330) );
  XOR U14028 ( .A(b[13]), .B(a[92]), .Z(n13477) );
  NAND U14029 ( .A(n37295), .B(n13477), .Z(n13329) );
  AND U14030 ( .A(n13330), .B(n13329), .Z(n13421) );
  NAND U14031 ( .A(n186), .B(n13331), .Z(n13333) );
  XOR U14032 ( .A(b[11]), .B(a[94]), .Z(n13480) );
  NAND U14033 ( .A(n37097), .B(n13480), .Z(n13332) );
  NAND U14034 ( .A(n13333), .B(n13332), .Z(n13420) );
  XNOR U14035 ( .A(n13421), .B(n13420), .Z(n13422) );
  NAND U14036 ( .A(n188), .B(n13334), .Z(n13336) );
  XOR U14037 ( .A(b[15]), .B(a[90]), .Z(n13483) );
  NAND U14038 ( .A(n37382), .B(n13483), .Z(n13335) );
  AND U14039 ( .A(n13336), .B(n13335), .Z(n13417) );
  NAND U14040 ( .A(n38064), .B(n13337), .Z(n13339) );
  XOR U14041 ( .A(b[21]), .B(a[84]), .Z(n13486) );
  NAND U14042 ( .A(n37993), .B(n13486), .Z(n13338) );
  AND U14043 ( .A(n13339), .B(n13338), .Z(n13415) );
  NAND U14044 ( .A(n185), .B(n13340), .Z(n13342) );
  XOR U14045 ( .A(b[9]), .B(a[96]), .Z(n13489) );
  NAND U14046 ( .A(n36805), .B(n13489), .Z(n13341) );
  NAND U14047 ( .A(n13342), .B(n13341), .Z(n13414) );
  XNOR U14048 ( .A(n13415), .B(n13414), .Z(n13416) );
  XOR U14049 ( .A(n13417), .B(n13416), .Z(n13423) );
  XOR U14050 ( .A(n13422), .B(n13423), .Z(n13429) );
  XOR U14051 ( .A(n13428), .B(n13429), .Z(n13441) );
  XNOR U14052 ( .A(n13440), .B(n13441), .Z(n13372) );
  XNOR U14053 ( .A(n13373), .B(n13372), .Z(n13374) );
  XOR U14054 ( .A(n13375), .B(n13374), .Z(n13493) );
  XNOR U14055 ( .A(n13492), .B(n13493), .Z(n13494) );
  XNOR U14056 ( .A(n13495), .B(n13494), .Z(n13500) );
  XOR U14057 ( .A(n13501), .B(n13500), .Z(n13367) );
  NANDN U14058 ( .A(n13344), .B(n13343), .Z(n13348) );
  NANDN U14059 ( .A(n13346), .B(n13345), .Z(n13347) );
  AND U14060 ( .A(n13348), .B(n13347), .Z(n13366) );
  XNOR U14061 ( .A(n13367), .B(n13366), .Z(n13368) );
  NANDN U14062 ( .A(n13350), .B(n13349), .Z(n13354) );
  NAND U14063 ( .A(n13352), .B(n13351), .Z(n13353) );
  NAND U14064 ( .A(n13354), .B(n13353), .Z(n13369) );
  XNOR U14065 ( .A(n13368), .B(n13369), .Z(n13360) );
  XNOR U14066 ( .A(n13361), .B(n13360), .Z(n13362) );
  XNOR U14067 ( .A(n13363), .B(n13362), .Z(n13504) );
  XNOR U14068 ( .A(sreg[328]), .B(n13504), .Z(n13506) );
  NANDN U14069 ( .A(sreg[327]), .B(n13355), .Z(n13359) );
  NAND U14070 ( .A(n13357), .B(n13356), .Z(n13358) );
  NAND U14071 ( .A(n13359), .B(n13358), .Z(n13505) );
  XNOR U14072 ( .A(n13506), .B(n13505), .Z(c[328]) );
  NANDN U14073 ( .A(n13361), .B(n13360), .Z(n13365) );
  NANDN U14074 ( .A(n13363), .B(n13362), .Z(n13364) );
  AND U14075 ( .A(n13365), .B(n13364), .Z(n13512) );
  NANDN U14076 ( .A(n13367), .B(n13366), .Z(n13371) );
  NANDN U14077 ( .A(n13369), .B(n13368), .Z(n13370) );
  AND U14078 ( .A(n13371), .B(n13370), .Z(n13510) );
  NANDN U14079 ( .A(n13373), .B(n13372), .Z(n13377) );
  NANDN U14080 ( .A(n13375), .B(n13374), .Z(n13376) );
  AND U14081 ( .A(n13377), .B(n13376), .Z(n13522) );
  NANDN U14082 ( .A(n13379), .B(n13378), .Z(n13383) );
  NAND U14083 ( .A(n13381), .B(n13380), .Z(n13382) );
  AND U14084 ( .A(n13383), .B(n13382), .Z(n13521) );
  XNOR U14085 ( .A(n13522), .B(n13521), .Z(n13524) );
  NANDN U14086 ( .A(n13385), .B(n13384), .Z(n13389) );
  NANDN U14087 ( .A(n13387), .B(n13386), .Z(n13388) );
  AND U14088 ( .A(n13389), .B(n13388), .Z(n13601) );
  NAND U14089 ( .A(n38385), .B(n13390), .Z(n13392) );
  XOR U14090 ( .A(b[27]), .B(a[79]), .Z(n13545) );
  NAND U14091 ( .A(n38343), .B(n13545), .Z(n13391) );
  AND U14092 ( .A(n13392), .B(n13391), .Z(n13608) );
  NAND U14093 ( .A(n183), .B(n13393), .Z(n13395) );
  XOR U14094 ( .A(b[5]), .B(a[101]), .Z(n13548) );
  NAND U14095 ( .A(n36296), .B(n13548), .Z(n13394) );
  AND U14096 ( .A(n13395), .B(n13394), .Z(n13606) );
  NAND U14097 ( .A(n190), .B(n13396), .Z(n13398) );
  XOR U14098 ( .A(b[19]), .B(a[87]), .Z(n13551) );
  NAND U14099 ( .A(n37821), .B(n13551), .Z(n13397) );
  NAND U14100 ( .A(n13398), .B(n13397), .Z(n13605) );
  XNOR U14101 ( .A(n13606), .B(n13605), .Z(n13607) );
  XNOR U14102 ( .A(n13608), .B(n13607), .Z(n13599) );
  NAND U14103 ( .A(n38470), .B(n13399), .Z(n13401) );
  XOR U14104 ( .A(b[31]), .B(a[75]), .Z(n13554) );
  NAND U14105 ( .A(n38453), .B(n13554), .Z(n13400) );
  AND U14106 ( .A(n13401), .B(n13400), .Z(n13566) );
  NAND U14107 ( .A(n181), .B(n13402), .Z(n13404) );
  XOR U14108 ( .A(b[3]), .B(a[103]), .Z(n13557) );
  NAND U14109 ( .A(n182), .B(n13557), .Z(n13403) );
  AND U14110 ( .A(n13404), .B(n13403), .Z(n13564) );
  NAND U14111 ( .A(n189), .B(n13405), .Z(n13407) );
  XOR U14112 ( .A(b[17]), .B(a[89]), .Z(n13560) );
  NAND U14113 ( .A(n37652), .B(n13560), .Z(n13406) );
  NAND U14114 ( .A(n13407), .B(n13406), .Z(n13563) );
  XNOR U14115 ( .A(n13564), .B(n13563), .Z(n13565) );
  XOR U14116 ( .A(n13566), .B(n13565), .Z(n13600) );
  XOR U14117 ( .A(n13599), .B(n13600), .Z(n13602) );
  XOR U14118 ( .A(n13601), .B(n13602), .Z(n13534) );
  NANDN U14119 ( .A(n13409), .B(n13408), .Z(n13413) );
  NANDN U14120 ( .A(n13411), .B(n13410), .Z(n13412) );
  AND U14121 ( .A(n13413), .B(n13412), .Z(n13587) );
  NANDN U14122 ( .A(n13415), .B(n13414), .Z(n13419) );
  NANDN U14123 ( .A(n13417), .B(n13416), .Z(n13418) );
  NAND U14124 ( .A(n13419), .B(n13418), .Z(n13588) );
  XNOR U14125 ( .A(n13587), .B(n13588), .Z(n13589) );
  NANDN U14126 ( .A(n13421), .B(n13420), .Z(n13425) );
  NANDN U14127 ( .A(n13423), .B(n13422), .Z(n13424) );
  NAND U14128 ( .A(n13425), .B(n13424), .Z(n13590) );
  XNOR U14129 ( .A(n13589), .B(n13590), .Z(n13533) );
  XNOR U14130 ( .A(n13534), .B(n13533), .Z(n13536) );
  NANDN U14131 ( .A(n13427), .B(n13426), .Z(n13431) );
  NANDN U14132 ( .A(n13429), .B(n13428), .Z(n13430) );
  AND U14133 ( .A(n13431), .B(n13430), .Z(n13535) );
  XOR U14134 ( .A(n13536), .B(n13535), .Z(n13650) );
  NANDN U14135 ( .A(n13433), .B(n13432), .Z(n13437) );
  NANDN U14136 ( .A(n13435), .B(n13434), .Z(n13436) );
  AND U14137 ( .A(n13437), .B(n13436), .Z(n13647) );
  NANDN U14138 ( .A(n13439), .B(n13438), .Z(n13443) );
  NANDN U14139 ( .A(n13441), .B(n13440), .Z(n13442) );
  AND U14140 ( .A(n13443), .B(n13442), .Z(n13530) );
  NANDN U14141 ( .A(n13445), .B(n13444), .Z(n13449) );
  OR U14142 ( .A(n13447), .B(n13446), .Z(n13448) );
  AND U14143 ( .A(n13449), .B(n13448), .Z(n13528) );
  NANDN U14144 ( .A(n13451), .B(n13450), .Z(n13455) );
  NANDN U14145 ( .A(n13453), .B(n13452), .Z(n13454) );
  AND U14146 ( .A(n13455), .B(n13454), .Z(n13594) );
  NANDN U14147 ( .A(n13457), .B(n13456), .Z(n13461) );
  NANDN U14148 ( .A(n13459), .B(n13458), .Z(n13460) );
  NAND U14149 ( .A(n13461), .B(n13460), .Z(n13593) );
  XNOR U14150 ( .A(n13594), .B(n13593), .Z(n13595) );
  NAND U14151 ( .A(b[0]), .B(a[105]), .Z(n13462) );
  XNOR U14152 ( .A(b[1]), .B(n13462), .Z(n13464) );
  NANDN U14153 ( .A(b[0]), .B(a[104]), .Z(n13463) );
  NAND U14154 ( .A(n13464), .B(n13463), .Z(n13542) );
  NAND U14155 ( .A(n194), .B(n13465), .Z(n13467) );
  XOR U14156 ( .A(b[29]), .B(a[77]), .Z(n13620) );
  NAND U14157 ( .A(n38456), .B(n13620), .Z(n13466) );
  AND U14158 ( .A(n13467), .B(n13466), .Z(n13540) );
  AND U14159 ( .A(b[31]), .B(a[73]), .Z(n13539) );
  XNOR U14160 ( .A(n13540), .B(n13539), .Z(n13541) );
  XNOR U14161 ( .A(n13542), .B(n13541), .Z(n13581) );
  NAND U14162 ( .A(n38185), .B(n13468), .Z(n13470) );
  XOR U14163 ( .A(b[23]), .B(a[83]), .Z(n13623) );
  NAND U14164 ( .A(n38132), .B(n13623), .Z(n13469) );
  AND U14165 ( .A(n13470), .B(n13469), .Z(n13614) );
  NAND U14166 ( .A(n184), .B(n13471), .Z(n13473) );
  XOR U14167 ( .A(b[7]), .B(a[99]), .Z(n13626) );
  NAND U14168 ( .A(n36592), .B(n13626), .Z(n13472) );
  AND U14169 ( .A(n13473), .B(n13472), .Z(n13612) );
  NAND U14170 ( .A(n38289), .B(n13474), .Z(n13476) );
  XOR U14171 ( .A(b[25]), .B(a[81]), .Z(n13629) );
  NAND U14172 ( .A(n38247), .B(n13629), .Z(n13475) );
  NAND U14173 ( .A(n13476), .B(n13475), .Z(n13611) );
  XNOR U14174 ( .A(n13612), .B(n13611), .Z(n13613) );
  XOR U14175 ( .A(n13614), .B(n13613), .Z(n13582) );
  XNOR U14176 ( .A(n13581), .B(n13582), .Z(n13583) );
  NAND U14177 ( .A(n187), .B(n13477), .Z(n13479) );
  XOR U14178 ( .A(b[13]), .B(a[93]), .Z(n13632) );
  NAND U14179 ( .A(n37295), .B(n13632), .Z(n13478) );
  AND U14180 ( .A(n13479), .B(n13478), .Z(n13576) );
  NAND U14181 ( .A(n186), .B(n13480), .Z(n13482) );
  XOR U14182 ( .A(b[11]), .B(a[95]), .Z(n13635) );
  NAND U14183 ( .A(n37097), .B(n13635), .Z(n13481) );
  NAND U14184 ( .A(n13482), .B(n13481), .Z(n13575) );
  XNOR U14185 ( .A(n13576), .B(n13575), .Z(n13577) );
  NAND U14186 ( .A(n188), .B(n13483), .Z(n13485) );
  XOR U14187 ( .A(b[15]), .B(a[91]), .Z(n13638) );
  NAND U14188 ( .A(n37382), .B(n13638), .Z(n13484) );
  AND U14189 ( .A(n13485), .B(n13484), .Z(n13572) );
  NAND U14190 ( .A(n38064), .B(n13486), .Z(n13488) );
  XOR U14191 ( .A(b[21]), .B(a[85]), .Z(n13641) );
  NAND U14192 ( .A(n37993), .B(n13641), .Z(n13487) );
  AND U14193 ( .A(n13488), .B(n13487), .Z(n13570) );
  NAND U14194 ( .A(n185), .B(n13489), .Z(n13491) );
  XOR U14195 ( .A(b[9]), .B(a[97]), .Z(n13644) );
  NAND U14196 ( .A(n36805), .B(n13644), .Z(n13490) );
  NAND U14197 ( .A(n13491), .B(n13490), .Z(n13569) );
  XNOR U14198 ( .A(n13570), .B(n13569), .Z(n13571) );
  XOR U14199 ( .A(n13572), .B(n13571), .Z(n13578) );
  XOR U14200 ( .A(n13577), .B(n13578), .Z(n13584) );
  XOR U14201 ( .A(n13583), .B(n13584), .Z(n13596) );
  XNOR U14202 ( .A(n13595), .B(n13596), .Z(n13527) );
  XNOR U14203 ( .A(n13528), .B(n13527), .Z(n13529) );
  XOR U14204 ( .A(n13530), .B(n13529), .Z(n13648) );
  XNOR U14205 ( .A(n13647), .B(n13648), .Z(n13649) );
  XNOR U14206 ( .A(n13650), .B(n13649), .Z(n13523) );
  XOR U14207 ( .A(n13524), .B(n13523), .Z(n13516) );
  NANDN U14208 ( .A(n13493), .B(n13492), .Z(n13497) );
  NANDN U14209 ( .A(n13495), .B(n13494), .Z(n13496) );
  AND U14210 ( .A(n13497), .B(n13496), .Z(n13515) );
  XNOR U14211 ( .A(n13516), .B(n13515), .Z(n13517) );
  NANDN U14212 ( .A(n13499), .B(n13498), .Z(n13503) );
  NAND U14213 ( .A(n13501), .B(n13500), .Z(n13502) );
  NAND U14214 ( .A(n13503), .B(n13502), .Z(n13518) );
  XNOR U14215 ( .A(n13517), .B(n13518), .Z(n13509) );
  XNOR U14216 ( .A(n13510), .B(n13509), .Z(n13511) );
  XNOR U14217 ( .A(n13512), .B(n13511), .Z(n13653) );
  XNOR U14218 ( .A(sreg[329]), .B(n13653), .Z(n13655) );
  NANDN U14219 ( .A(sreg[328]), .B(n13504), .Z(n13508) );
  NAND U14220 ( .A(n13506), .B(n13505), .Z(n13507) );
  NAND U14221 ( .A(n13508), .B(n13507), .Z(n13654) );
  XNOR U14222 ( .A(n13655), .B(n13654), .Z(c[329]) );
  NANDN U14223 ( .A(n13510), .B(n13509), .Z(n13514) );
  NANDN U14224 ( .A(n13512), .B(n13511), .Z(n13513) );
  AND U14225 ( .A(n13514), .B(n13513), .Z(n13661) );
  NANDN U14226 ( .A(n13516), .B(n13515), .Z(n13520) );
  NANDN U14227 ( .A(n13518), .B(n13517), .Z(n13519) );
  AND U14228 ( .A(n13520), .B(n13519), .Z(n13659) );
  NANDN U14229 ( .A(n13522), .B(n13521), .Z(n13526) );
  NAND U14230 ( .A(n13524), .B(n13523), .Z(n13525) );
  AND U14231 ( .A(n13526), .B(n13525), .Z(n13666) );
  NANDN U14232 ( .A(n13528), .B(n13527), .Z(n13532) );
  NANDN U14233 ( .A(n13530), .B(n13529), .Z(n13531) );
  AND U14234 ( .A(n13532), .B(n13531), .Z(n13797) );
  NANDN U14235 ( .A(n13534), .B(n13533), .Z(n13538) );
  NAND U14236 ( .A(n13536), .B(n13535), .Z(n13537) );
  AND U14237 ( .A(n13538), .B(n13537), .Z(n13796) );
  XNOR U14238 ( .A(n13797), .B(n13796), .Z(n13799) );
  NANDN U14239 ( .A(n13540), .B(n13539), .Z(n13544) );
  NANDN U14240 ( .A(n13542), .B(n13541), .Z(n13543) );
  AND U14241 ( .A(n13544), .B(n13543), .Z(n13744) );
  NAND U14242 ( .A(n38385), .B(n13545), .Z(n13547) );
  XOR U14243 ( .A(b[27]), .B(a[80]), .Z(n13688) );
  NAND U14244 ( .A(n38343), .B(n13688), .Z(n13546) );
  AND U14245 ( .A(n13547), .B(n13546), .Z(n13751) );
  NAND U14246 ( .A(n183), .B(n13548), .Z(n13550) );
  XOR U14247 ( .A(b[5]), .B(a[102]), .Z(n13691) );
  NAND U14248 ( .A(n36296), .B(n13691), .Z(n13549) );
  AND U14249 ( .A(n13550), .B(n13549), .Z(n13749) );
  NAND U14250 ( .A(n190), .B(n13551), .Z(n13553) );
  XOR U14251 ( .A(b[19]), .B(a[88]), .Z(n13694) );
  NAND U14252 ( .A(n37821), .B(n13694), .Z(n13552) );
  NAND U14253 ( .A(n13553), .B(n13552), .Z(n13748) );
  XNOR U14254 ( .A(n13749), .B(n13748), .Z(n13750) );
  XNOR U14255 ( .A(n13751), .B(n13750), .Z(n13742) );
  NAND U14256 ( .A(n38470), .B(n13554), .Z(n13556) );
  XOR U14257 ( .A(b[31]), .B(a[76]), .Z(n13697) );
  NAND U14258 ( .A(n38453), .B(n13697), .Z(n13555) );
  AND U14259 ( .A(n13556), .B(n13555), .Z(n13709) );
  NAND U14260 ( .A(n181), .B(n13557), .Z(n13559) );
  XOR U14261 ( .A(b[3]), .B(a[104]), .Z(n13700) );
  NAND U14262 ( .A(n182), .B(n13700), .Z(n13558) );
  AND U14263 ( .A(n13559), .B(n13558), .Z(n13707) );
  NAND U14264 ( .A(n189), .B(n13560), .Z(n13562) );
  XOR U14265 ( .A(b[17]), .B(a[90]), .Z(n13703) );
  NAND U14266 ( .A(n37652), .B(n13703), .Z(n13561) );
  NAND U14267 ( .A(n13562), .B(n13561), .Z(n13706) );
  XNOR U14268 ( .A(n13707), .B(n13706), .Z(n13708) );
  XOR U14269 ( .A(n13709), .B(n13708), .Z(n13743) );
  XOR U14270 ( .A(n13742), .B(n13743), .Z(n13745) );
  XOR U14271 ( .A(n13744), .B(n13745), .Z(n13677) );
  NANDN U14272 ( .A(n13564), .B(n13563), .Z(n13568) );
  NANDN U14273 ( .A(n13566), .B(n13565), .Z(n13567) );
  AND U14274 ( .A(n13568), .B(n13567), .Z(n13730) );
  NANDN U14275 ( .A(n13570), .B(n13569), .Z(n13574) );
  NANDN U14276 ( .A(n13572), .B(n13571), .Z(n13573) );
  NAND U14277 ( .A(n13574), .B(n13573), .Z(n13731) );
  XNOR U14278 ( .A(n13730), .B(n13731), .Z(n13732) );
  NANDN U14279 ( .A(n13576), .B(n13575), .Z(n13580) );
  NANDN U14280 ( .A(n13578), .B(n13577), .Z(n13579) );
  NAND U14281 ( .A(n13580), .B(n13579), .Z(n13733) );
  XNOR U14282 ( .A(n13732), .B(n13733), .Z(n13676) );
  XNOR U14283 ( .A(n13677), .B(n13676), .Z(n13679) );
  NANDN U14284 ( .A(n13582), .B(n13581), .Z(n13586) );
  NANDN U14285 ( .A(n13584), .B(n13583), .Z(n13585) );
  AND U14286 ( .A(n13586), .B(n13585), .Z(n13678) );
  XOR U14287 ( .A(n13679), .B(n13678), .Z(n13793) );
  NANDN U14288 ( .A(n13588), .B(n13587), .Z(n13592) );
  NANDN U14289 ( .A(n13590), .B(n13589), .Z(n13591) );
  AND U14290 ( .A(n13592), .B(n13591), .Z(n13790) );
  NANDN U14291 ( .A(n13594), .B(n13593), .Z(n13598) );
  NANDN U14292 ( .A(n13596), .B(n13595), .Z(n13597) );
  AND U14293 ( .A(n13598), .B(n13597), .Z(n13673) );
  NANDN U14294 ( .A(n13600), .B(n13599), .Z(n13604) );
  OR U14295 ( .A(n13602), .B(n13601), .Z(n13603) );
  AND U14296 ( .A(n13604), .B(n13603), .Z(n13671) );
  NANDN U14297 ( .A(n13606), .B(n13605), .Z(n13610) );
  NANDN U14298 ( .A(n13608), .B(n13607), .Z(n13609) );
  AND U14299 ( .A(n13610), .B(n13609), .Z(n13737) );
  NANDN U14300 ( .A(n13612), .B(n13611), .Z(n13616) );
  NANDN U14301 ( .A(n13614), .B(n13613), .Z(n13615) );
  NAND U14302 ( .A(n13616), .B(n13615), .Z(n13736) );
  XNOR U14303 ( .A(n13737), .B(n13736), .Z(n13738) );
  NAND U14304 ( .A(b[0]), .B(a[106]), .Z(n13617) );
  XNOR U14305 ( .A(b[1]), .B(n13617), .Z(n13619) );
  NANDN U14306 ( .A(b[0]), .B(a[105]), .Z(n13618) );
  NAND U14307 ( .A(n13619), .B(n13618), .Z(n13685) );
  NAND U14308 ( .A(n194), .B(n13620), .Z(n13622) );
  XOR U14309 ( .A(b[29]), .B(a[78]), .Z(n13760) );
  NAND U14310 ( .A(n38456), .B(n13760), .Z(n13621) );
  AND U14311 ( .A(n13622), .B(n13621), .Z(n13683) );
  AND U14312 ( .A(b[31]), .B(a[74]), .Z(n13682) );
  XNOR U14313 ( .A(n13683), .B(n13682), .Z(n13684) );
  XNOR U14314 ( .A(n13685), .B(n13684), .Z(n13724) );
  NAND U14315 ( .A(n38185), .B(n13623), .Z(n13625) );
  XOR U14316 ( .A(b[23]), .B(a[84]), .Z(n13766) );
  NAND U14317 ( .A(n38132), .B(n13766), .Z(n13624) );
  AND U14318 ( .A(n13625), .B(n13624), .Z(n13757) );
  NAND U14319 ( .A(n184), .B(n13626), .Z(n13628) );
  XOR U14320 ( .A(b[7]), .B(a[100]), .Z(n13769) );
  NAND U14321 ( .A(n36592), .B(n13769), .Z(n13627) );
  AND U14322 ( .A(n13628), .B(n13627), .Z(n13755) );
  NAND U14323 ( .A(n38289), .B(n13629), .Z(n13631) );
  XOR U14324 ( .A(b[25]), .B(a[82]), .Z(n13772) );
  NAND U14325 ( .A(n38247), .B(n13772), .Z(n13630) );
  NAND U14326 ( .A(n13631), .B(n13630), .Z(n13754) );
  XNOR U14327 ( .A(n13755), .B(n13754), .Z(n13756) );
  XOR U14328 ( .A(n13757), .B(n13756), .Z(n13725) );
  XNOR U14329 ( .A(n13724), .B(n13725), .Z(n13726) );
  NAND U14330 ( .A(n187), .B(n13632), .Z(n13634) );
  XOR U14331 ( .A(b[13]), .B(a[94]), .Z(n13775) );
  NAND U14332 ( .A(n37295), .B(n13775), .Z(n13633) );
  AND U14333 ( .A(n13634), .B(n13633), .Z(n13719) );
  NAND U14334 ( .A(n186), .B(n13635), .Z(n13637) );
  XOR U14335 ( .A(b[11]), .B(a[96]), .Z(n13778) );
  NAND U14336 ( .A(n37097), .B(n13778), .Z(n13636) );
  NAND U14337 ( .A(n13637), .B(n13636), .Z(n13718) );
  XNOR U14338 ( .A(n13719), .B(n13718), .Z(n13720) );
  NAND U14339 ( .A(n188), .B(n13638), .Z(n13640) );
  XOR U14340 ( .A(b[15]), .B(a[92]), .Z(n13781) );
  NAND U14341 ( .A(n37382), .B(n13781), .Z(n13639) );
  AND U14342 ( .A(n13640), .B(n13639), .Z(n13715) );
  NAND U14343 ( .A(n38064), .B(n13641), .Z(n13643) );
  XOR U14344 ( .A(b[21]), .B(a[86]), .Z(n13784) );
  NAND U14345 ( .A(n37993), .B(n13784), .Z(n13642) );
  AND U14346 ( .A(n13643), .B(n13642), .Z(n13713) );
  NAND U14347 ( .A(n185), .B(n13644), .Z(n13646) );
  XOR U14348 ( .A(b[9]), .B(a[98]), .Z(n13787) );
  NAND U14349 ( .A(n36805), .B(n13787), .Z(n13645) );
  NAND U14350 ( .A(n13646), .B(n13645), .Z(n13712) );
  XNOR U14351 ( .A(n13713), .B(n13712), .Z(n13714) );
  XOR U14352 ( .A(n13715), .B(n13714), .Z(n13721) );
  XOR U14353 ( .A(n13720), .B(n13721), .Z(n13727) );
  XOR U14354 ( .A(n13726), .B(n13727), .Z(n13739) );
  XNOR U14355 ( .A(n13738), .B(n13739), .Z(n13670) );
  XNOR U14356 ( .A(n13671), .B(n13670), .Z(n13672) );
  XOR U14357 ( .A(n13673), .B(n13672), .Z(n13791) );
  XNOR U14358 ( .A(n13790), .B(n13791), .Z(n13792) );
  XNOR U14359 ( .A(n13793), .B(n13792), .Z(n13798) );
  XOR U14360 ( .A(n13799), .B(n13798), .Z(n13665) );
  NANDN U14361 ( .A(n13648), .B(n13647), .Z(n13652) );
  NANDN U14362 ( .A(n13650), .B(n13649), .Z(n13651) );
  AND U14363 ( .A(n13652), .B(n13651), .Z(n13664) );
  XOR U14364 ( .A(n13665), .B(n13664), .Z(n13667) );
  XNOR U14365 ( .A(n13666), .B(n13667), .Z(n13658) );
  XNOR U14366 ( .A(n13659), .B(n13658), .Z(n13660) );
  XNOR U14367 ( .A(n13661), .B(n13660), .Z(n13802) );
  XNOR U14368 ( .A(sreg[330]), .B(n13802), .Z(n13804) );
  NANDN U14369 ( .A(sreg[329]), .B(n13653), .Z(n13657) );
  NAND U14370 ( .A(n13655), .B(n13654), .Z(n13656) );
  NAND U14371 ( .A(n13657), .B(n13656), .Z(n13803) );
  XNOR U14372 ( .A(n13804), .B(n13803), .Z(c[330]) );
  NANDN U14373 ( .A(n13659), .B(n13658), .Z(n13663) );
  NANDN U14374 ( .A(n13661), .B(n13660), .Z(n13662) );
  AND U14375 ( .A(n13663), .B(n13662), .Z(n13810) );
  NANDN U14376 ( .A(n13665), .B(n13664), .Z(n13669) );
  NANDN U14377 ( .A(n13667), .B(n13666), .Z(n13668) );
  AND U14378 ( .A(n13669), .B(n13668), .Z(n13808) );
  NANDN U14379 ( .A(n13671), .B(n13670), .Z(n13675) );
  NANDN U14380 ( .A(n13673), .B(n13672), .Z(n13674) );
  AND U14381 ( .A(n13675), .B(n13674), .Z(n13946) );
  NANDN U14382 ( .A(n13677), .B(n13676), .Z(n13681) );
  NAND U14383 ( .A(n13679), .B(n13678), .Z(n13680) );
  AND U14384 ( .A(n13681), .B(n13680), .Z(n13945) );
  XNOR U14385 ( .A(n13946), .B(n13945), .Z(n13948) );
  NANDN U14386 ( .A(n13683), .B(n13682), .Z(n13687) );
  NANDN U14387 ( .A(n13685), .B(n13684), .Z(n13686) );
  AND U14388 ( .A(n13687), .B(n13686), .Z(n13893) );
  NAND U14389 ( .A(n38385), .B(n13688), .Z(n13690) );
  XOR U14390 ( .A(b[27]), .B(a[81]), .Z(n13837) );
  NAND U14391 ( .A(n38343), .B(n13837), .Z(n13689) );
  AND U14392 ( .A(n13690), .B(n13689), .Z(n13900) );
  NAND U14393 ( .A(n183), .B(n13691), .Z(n13693) );
  XOR U14394 ( .A(b[5]), .B(a[103]), .Z(n13840) );
  NAND U14395 ( .A(n36296), .B(n13840), .Z(n13692) );
  AND U14396 ( .A(n13693), .B(n13692), .Z(n13898) );
  NAND U14397 ( .A(n190), .B(n13694), .Z(n13696) );
  XOR U14398 ( .A(b[19]), .B(a[89]), .Z(n13843) );
  NAND U14399 ( .A(n37821), .B(n13843), .Z(n13695) );
  NAND U14400 ( .A(n13696), .B(n13695), .Z(n13897) );
  XNOR U14401 ( .A(n13898), .B(n13897), .Z(n13899) );
  XNOR U14402 ( .A(n13900), .B(n13899), .Z(n13891) );
  NAND U14403 ( .A(n38470), .B(n13697), .Z(n13699) );
  XOR U14404 ( .A(b[31]), .B(a[77]), .Z(n13846) );
  NAND U14405 ( .A(n38453), .B(n13846), .Z(n13698) );
  AND U14406 ( .A(n13699), .B(n13698), .Z(n13858) );
  NAND U14407 ( .A(n181), .B(n13700), .Z(n13702) );
  XOR U14408 ( .A(b[3]), .B(a[105]), .Z(n13849) );
  NAND U14409 ( .A(n182), .B(n13849), .Z(n13701) );
  AND U14410 ( .A(n13702), .B(n13701), .Z(n13856) );
  NAND U14411 ( .A(n189), .B(n13703), .Z(n13705) );
  XOR U14412 ( .A(b[17]), .B(a[91]), .Z(n13852) );
  NAND U14413 ( .A(n37652), .B(n13852), .Z(n13704) );
  NAND U14414 ( .A(n13705), .B(n13704), .Z(n13855) );
  XNOR U14415 ( .A(n13856), .B(n13855), .Z(n13857) );
  XOR U14416 ( .A(n13858), .B(n13857), .Z(n13892) );
  XOR U14417 ( .A(n13891), .B(n13892), .Z(n13894) );
  XOR U14418 ( .A(n13893), .B(n13894), .Z(n13826) );
  NANDN U14419 ( .A(n13707), .B(n13706), .Z(n13711) );
  NANDN U14420 ( .A(n13709), .B(n13708), .Z(n13710) );
  AND U14421 ( .A(n13711), .B(n13710), .Z(n13879) );
  NANDN U14422 ( .A(n13713), .B(n13712), .Z(n13717) );
  NANDN U14423 ( .A(n13715), .B(n13714), .Z(n13716) );
  NAND U14424 ( .A(n13717), .B(n13716), .Z(n13880) );
  XNOR U14425 ( .A(n13879), .B(n13880), .Z(n13881) );
  NANDN U14426 ( .A(n13719), .B(n13718), .Z(n13723) );
  NANDN U14427 ( .A(n13721), .B(n13720), .Z(n13722) );
  NAND U14428 ( .A(n13723), .B(n13722), .Z(n13882) );
  XNOR U14429 ( .A(n13881), .B(n13882), .Z(n13825) );
  XNOR U14430 ( .A(n13826), .B(n13825), .Z(n13828) );
  NANDN U14431 ( .A(n13725), .B(n13724), .Z(n13729) );
  NANDN U14432 ( .A(n13727), .B(n13726), .Z(n13728) );
  AND U14433 ( .A(n13729), .B(n13728), .Z(n13827) );
  XOR U14434 ( .A(n13828), .B(n13827), .Z(n13942) );
  NANDN U14435 ( .A(n13731), .B(n13730), .Z(n13735) );
  NANDN U14436 ( .A(n13733), .B(n13732), .Z(n13734) );
  AND U14437 ( .A(n13735), .B(n13734), .Z(n13939) );
  NANDN U14438 ( .A(n13737), .B(n13736), .Z(n13741) );
  NANDN U14439 ( .A(n13739), .B(n13738), .Z(n13740) );
  AND U14440 ( .A(n13741), .B(n13740), .Z(n13822) );
  NANDN U14441 ( .A(n13743), .B(n13742), .Z(n13747) );
  OR U14442 ( .A(n13745), .B(n13744), .Z(n13746) );
  AND U14443 ( .A(n13747), .B(n13746), .Z(n13820) );
  NANDN U14444 ( .A(n13749), .B(n13748), .Z(n13753) );
  NANDN U14445 ( .A(n13751), .B(n13750), .Z(n13752) );
  AND U14446 ( .A(n13753), .B(n13752), .Z(n13886) );
  NANDN U14447 ( .A(n13755), .B(n13754), .Z(n13759) );
  NANDN U14448 ( .A(n13757), .B(n13756), .Z(n13758) );
  NAND U14449 ( .A(n13759), .B(n13758), .Z(n13885) );
  XNOR U14450 ( .A(n13886), .B(n13885), .Z(n13887) );
  NAND U14451 ( .A(n194), .B(n13760), .Z(n13762) );
  XOR U14452 ( .A(b[29]), .B(a[79]), .Z(n13909) );
  NAND U14453 ( .A(n38456), .B(n13909), .Z(n13761) );
  AND U14454 ( .A(n13762), .B(n13761), .Z(n13832) );
  AND U14455 ( .A(b[31]), .B(a[75]), .Z(n13831) );
  XNOR U14456 ( .A(n13832), .B(n13831), .Z(n13833) );
  NAND U14457 ( .A(b[0]), .B(a[107]), .Z(n13763) );
  XNOR U14458 ( .A(b[1]), .B(n13763), .Z(n13765) );
  NANDN U14459 ( .A(b[0]), .B(a[106]), .Z(n13764) );
  NAND U14460 ( .A(n13765), .B(n13764), .Z(n13834) );
  XNOR U14461 ( .A(n13833), .B(n13834), .Z(n13873) );
  NAND U14462 ( .A(n38185), .B(n13766), .Z(n13768) );
  XOR U14463 ( .A(b[23]), .B(a[85]), .Z(n13915) );
  NAND U14464 ( .A(n38132), .B(n13915), .Z(n13767) );
  AND U14465 ( .A(n13768), .B(n13767), .Z(n13906) );
  NAND U14466 ( .A(n184), .B(n13769), .Z(n13771) );
  XOR U14467 ( .A(b[7]), .B(a[101]), .Z(n13918) );
  NAND U14468 ( .A(n36592), .B(n13918), .Z(n13770) );
  AND U14469 ( .A(n13771), .B(n13770), .Z(n13904) );
  NAND U14470 ( .A(n38289), .B(n13772), .Z(n13774) );
  XOR U14471 ( .A(b[25]), .B(a[83]), .Z(n13921) );
  NAND U14472 ( .A(n38247), .B(n13921), .Z(n13773) );
  NAND U14473 ( .A(n13774), .B(n13773), .Z(n13903) );
  XNOR U14474 ( .A(n13904), .B(n13903), .Z(n13905) );
  XOR U14475 ( .A(n13906), .B(n13905), .Z(n13874) );
  XNOR U14476 ( .A(n13873), .B(n13874), .Z(n13875) );
  NAND U14477 ( .A(n187), .B(n13775), .Z(n13777) );
  XOR U14478 ( .A(b[13]), .B(a[95]), .Z(n13924) );
  NAND U14479 ( .A(n37295), .B(n13924), .Z(n13776) );
  AND U14480 ( .A(n13777), .B(n13776), .Z(n13868) );
  NAND U14481 ( .A(n186), .B(n13778), .Z(n13780) );
  XOR U14482 ( .A(b[11]), .B(a[97]), .Z(n13927) );
  NAND U14483 ( .A(n37097), .B(n13927), .Z(n13779) );
  NAND U14484 ( .A(n13780), .B(n13779), .Z(n13867) );
  XNOR U14485 ( .A(n13868), .B(n13867), .Z(n13869) );
  NAND U14486 ( .A(n188), .B(n13781), .Z(n13783) );
  XOR U14487 ( .A(b[15]), .B(a[93]), .Z(n13930) );
  NAND U14488 ( .A(n37382), .B(n13930), .Z(n13782) );
  AND U14489 ( .A(n13783), .B(n13782), .Z(n13864) );
  NAND U14490 ( .A(n38064), .B(n13784), .Z(n13786) );
  XOR U14491 ( .A(b[21]), .B(a[87]), .Z(n13933) );
  NAND U14492 ( .A(n37993), .B(n13933), .Z(n13785) );
  AND U14493 ( .A(n13786), .B(n13785), .Z(n13862) );
  NAND U14494 ( .A(n185), .B(n13787), .Z(n13789) );
  XOR U14495 ( .A(b[9]), .B(a[99]), .Z(n13936) );
  NAND U14496 ( .A(n36805), .B(n13936), .Z(n13788) );
  NAND U14497 ( .A(n13789), .B(n13788), .Z(n13861) );
  XNOR U14498 ( .A(n13862), .B(n13861), .Z(n13863) );
  XOR U14499 ( .A(n13864), .B(n13863), .Z(n13870) );
  XOR U14500 ( .A(n13869), .B(n13870), .Z(n13876) );
  XOR U14501 ( .A(n13875), .B(n13876), .Z(n13888) );
  XNOR U14502 ( .A(n13887), .B(n13888), .Z(n13819) );
  XNOR U14503 ( .A(n13820), .B(n13819), .Z(n13821) );
  XOR U14504 ( .A(n13822), .B(n13821), .Z(n13940) );
  XNOR U14505 ( .A(n13939), .B(n13940), .Z(n13941) );
  XNOR U14506 ( .A(n13942), .B(n13941), .Z(n13947) );
  XOR U14507 ( .A(n13948), .B(n13947), .Z(n13814) );
  NANDN U14508 ( .A(n13791), .B(n13790), .Z(n13795) );
  NANDN U14509 ( .A(n13793), .B(n13792), .Z(n13794) );
  AND U14510 ( .A(n13795), .B(n13794), .Z(n13813) );
  XNOR U14511 ( .A(n13814), .B(n13813), .Z(n13815) );
  NANDN U14512 ( .A(n13797), .B(n13796), .Z(n13801) );
  NAND U14513 ( .A(n13799), .B(n13798), .Z(n13800) );
  NAND U14514 ( .A(n13801), .B(n13800), .Z(n13816) );
  XNOR U14515 ( .A(n13815), .B(n13816), .Z(n13807) );
  XNOR U14516 ( .A(n13808), .B(n13807), .Z(n13809) );
  XNOR U14517 ( .A(n13810), .B(n13809), .Z(n13951) );
  XNOR U14518 ( .A(sreg[331]), .B(n13951), .Z(n13953) );
  NANDN U14519 ( .A(sreg[330]), .B(n13802), .Z(n13806) );
  NAND U14520 ( .A(n13804), .B(n13803), .Z(n13805) );
  NAND U14521 ( .A(n13806), .B(n13805), .Z(n13952) );
  XNOR U14522 ( .A(n13953), .B(n13952), .Z(c[331]) );
  NANDN U14523 ( .A(n13808), .B(n13807), .Z(n13812) );
  NANDN U14524 ( .A(n13810), .B(n13809), .Z(n13811) );
  AND U14525 ( .A(n13812), .B(n13811), .Z(n13959) );
  NANDN U14526 ( .A(n13814), .B(n13813), .Z(n13818) );
  NANDN U14527 ( .A(n13816), .B(n13815), .Z(n13817) );
  AND U14528 ( .A(n13818), .B(n13817), .Z(n13957) );
  NANDN U14529 ( .A(n13820), .B(n13819), .Z(n13824) );
  NANDN U14530 ( .A(n13822), .B(n13821), .Z(n13823) );
  AND U14531 ( .A(n13824), .B(n13823), .Z(n13969) );
  NANDN U14532 ( .A(n13826), .B(n13825), .Z(n13830) );
  NAND U14533 ( .A(n13828), .B(n13827), .Z(n13829) );
  AND U14534 ( .A(n13830), .B(n13829), .Z(n13968) );
  XNOR U14535 ( .A(n13969), .B(n13968), .Z(n13971) );
  NANDN U14536 ( .A(n13832), .B(n13831), .Z(n13836) );
  NANDN U14537 ( .A(n13834), .B(n13833), .Z(n13835) );
  AND U14538 ( .A(n13836), .B(n13835), .Z(n14048) );
  NAND U14539 ( .A(n38385), .B(n13837), .Z(n13839) );
  XOR U14540 ( .A(b[27]), .B(a[82]), .Z(n13992) );
  NAND U14541 ( .A(n38343), .B(n13992), .Z(n13838) );
  AND U14542 ( .A(n13839), .B(n13838), .Z(n14055) );
  NAND U14543 ( .A(n183), .B(n13840), .Z(n13842) );
  XOR U14544 ( .A(b[5]), .B(a[104]), .Z(n13995) );
  NAND U14545 ( .A(n36296), .B(n13995), .Z(n13841) );
  AND U14546 ( .A(n13842), .B(n13841), .Z(n14053) );
  NAND U14547 ( .A(n190), .B(n13843), .Z(n13845) );
  XOR U14548 ( .A(b[19]), .B(a[90]), .Z(n13998) );
  NAND U14549 ( .A(n37821), .B(n13998), .Z(n13844) );
  NAND U14550 ( .A(n13845), .B(n13844), .Z(n14052) );
  XNOR U14551 ( .A(n14053), .B(n14052), .Z(n14054) );
  XNOR U14552 ( .A(n14055), .B(n14054), .Z(n14046) );
  NAND U14553 ( .A(n38470), .B(n13846), .Z(n13848) );
  XOR U14554 ( .A(b[31]), .B(a[78]), .Z(n14001) );
  NAND U14555 ( .A(n38453), .B(n14001), .Z(n13847) );
  AND U14556 ( .A(n13848), .B(n13847), .Z(n14013) );
  NAND U14557 ( .A(n181), .B(n13849), .Z(n13851) );
  XOR U14558 ( .A(b[3]), .B(a[106]), .Z(n14004) );
  NAND U14559 ( .A(n182), .B(n14004), .Z(n13850) );
  AND U14560 ( .A(n13851), .B(n13850), .Z(n14011) );
  NAND U14561 ( .A(n189), .B(n13852), .Z(n13854) );
  XOR U14562 ( .A(b[17]), .B(a[92]), .Z(n14007) );
  NAND U14563 ( .A(n37652), .B(n14007), .Z(n13853) );
  NAND U14564 ( .A(n13854), .B(n13853), .Z(n14010) );
  XNOR U14565 ( .A(n14011), .B(n14010), .Z(n14012) );
  XOR U14566 ( .A(n14013), .B(n14012), .Z(n14047) );
  XOR U14567 ( .A(n14046), .B(n14047), .Z(n14049) );
  XOR U14568 ( .A(n14048), .B(n14049), .Z(n13981) );
  NANDN U14569 ( .A(n13856), .B(n13855), .Z(n13860) );
  NANDN U14570 ( .A(n13858), .B(n13857), .Z(n13859) );
  AND U14571 ( .A(n13860), .B(n13859), .Z(n14034) );
  NANDN U14572 ( .A(n13862), .B(n13861), .Z(n13866) );
  NANDN U14573 ( .A(n13864), .B(n13863), .Z(n13865) );
  NAND U14574 ( .A(n13866), .B(n13865), .Z(n14035) );
  XNOR U14575 ( .A(n14034), .B(n14035), .Z(n14036) );
  NANDN U14576 ( .A(n13868), .B(n13867), .Z(n13872) );
  NANDN U14577 ( .A(n13870), .B(n13869), .Z(n13871) );
  NAND U14578 ( .A(n13872), .B(n13871), .Z(n14037) );
  XNOR U14579 ( .A(n14036), .B(n14037), .Z(n13980) );
  XNOR U14580 ( .A(n13981), .B(n13980), .Z(n13983) );
  NANDN U14581 ( .A(n13874), .B(n13873), .Z(n13878) );
  NANDN U14582 ( .A(n13876), .B(n13875), .Z(n13877) );
  AND U14583 ( .A(n13878), .B(n13877), .Z(n13982) );
  XOR U14584 ( .A(n13983), .B(n13982), .Z(n14097) );
  NANDN U14585 ( .A(n13880), .B(n13879), .Z(n13884) );
  NANDN U14586 ( .A(n13882), .B(n13881), .Z(n13883) );
  AND U14587 ( .A(n13884), .B(n13883), .Z(n14094) );
  NANDN U14588 ( .A(n13886), .B(n13885), .Z(n13890) );
  NANDN U14589 ( .A(n13888), .B(n13887), .Z(n13889) );
  AND U14590 ( .A(n13890), .B(n13889), .Z(n13977) );
  NANDN U14591 ( .A(n13892), .B(n13891), .Z(n13896) );
  OR U14592 ( .A(n13894), .B(n13893), .Z(n13895) );
  AND U14593 ( .A(n13896), .B(n13895), .Z(n13975) );
  NANDN U14594 ( .A(n13898), .B(n13897), .Z(n13902) );
  NANDN U14595 ( .A(n13900), .B(n13899), .Z(n13901) );
  AND U14596 ( .A(n13902), .B(n13901), .Z(n14041) );
  NANDN U14597 ( .A(n13904), .B(n13903), .Z(n13908) );
  NANDN U14598 ( .A(n13906), .B(n13905), .Z(n13907) );
  NAND U14599 ( .A(n13908), .B(n13907), .Z(n14040) );
  XNOR U14600 ( .A(n14041), .B(n14040), .Z(n14042) );
  NAND U14601 ( .A(n194), .B(n13909), .Z(n13911) );
  XOR U14602 ( .A(b[29]), .B(a[80]), .Z(n14067) );
  NAND U14603 ( .A(n38456), .B(n14067), .Z(n13910) );
  AND U14604 ( .A(n13911), .B(n13910), .Z(n13987) );
  AND U14605 ( .A(b[31]), .B(a[76]), .Z(n13986) );
  XNOR U14606 ( .A(n13987), .B(n13986), .Z(n13988) );
  NAND U14607 ( .A(b[0]), .B(a[108]), .Z(n13912) );
  XNOR U14608 ( .A(b[1]), .B(n13912), .Z(n13914) );
  NANDN U14609 ( .A(b[0]), .B(a[107]), .Z(n13913) );
  NAND U14610 ( .A(n13914), .B(n13913), .Z(n13989) );
  XNOR U14611 ( .A(n13988), .B(n13989), .Z(n14028) );
  NAND U14612 ( .A(n38185), .B(n13915), .Z(n13917) );
  XOR U14613 ( .A(b[23]), .B(a[86]), .Z(n14070) );
  NAND U14614 ( .A(n38132), .B(n14070), .Z(n13916) );
  AND U14615 ( .A(n13917), .B(n13916), .Z(n14061) );
  NAND U14616 ( .A(n184), .B(n13918), .Z(n13920) );
  XOR U14617 ( .A(b[7]), .B(a[102]), .Z(n14073) );
  NAND U14618 ( .A(n36592), .B(n14073), .Z(n13919) );
  AND U14619 ( .A(n13920), .B(n13919), .Z(n14059) );
  NAND U14620 ( .A(n38289), .B(n13921), .Z(n13923) );
  XOR U14621 ( .A(b[25]), .B(a[84]), .Z(n14076) );
  NAND U14622 ( .A(n38247), .B(n14076), .Z(n13922) );
  NAND U14623 ( .A(n13923), .B(n13922), .Z(n14058) );
  XNOR U14624 ( .A(n14059), .B(n14058), .Z(n14060) );
  XOR U14625 ( .A(n14061), .B(n14060), .Z(n14029) );
  XNOR U14626 ( .A(n14028), .B(n14029), .Z(n14030) );
  NAND U14627 ( .A(n187), .B(n13924), .Z(n13926) );
  XOR U14628 ( .A(b[13]), .B(a[96]), .Z(n14079) );
  NAND U14629 ( .A(n37295), .B(n14079), .Z(n13925) );
  AND U14630 ( .A(n13926), .B(n13925), .Z(n14023) );
  NAND U14631 ( .A(n186), .B(n13927), .Z(n13929) );
  XOR U14632 ( .A(b[11]), .B(a[98]), .Z(n14082) );
  NAND U14633 ( .A(n37097), .B(n14082), .Z(n13928) );
  NAND U14634 ( .A(n13929), .B(n13928), .Z(n14022) );
  XNOR U14635 ( .A(n14023), .B(n14022), .Z(n14024) );
  NAND U14636 ( .A(n188), .B(n13930), .Z(n13932) );
  XOR U14637 ( .A(b[15]), .B(a[94]), .Z(n14085) );
  NAND U14638 ( .A(n37382), .B(n14085), .Z(n13931) );
  AND U14639 ( .A(n13932), .B(n13931), .Z(n14019) );
  NAND U14640 ( .A(n38064), .B(n13933), .Z(n13935) );
  XOR U14641 ( .A(b[21]), .B(a[88]), .Z(n14088) );
  NAND U14642 ( .A(n37993), .B(n14088), .Z(n13934) );
  AND U14643 ( .A(n13935), .B(n13934), .Z(n14017) );
  NAND U14644 ( .A(n185), .B(n13936), .Z(n13938) );
  XOR U14645 ( .A(b[9]), .B(a[100]), .Z(n14091) );
  NAND U14646 ( .A(n36805), .B(n14091), .Z(n13937) );
  NAND U14647 ( .A(n13938), .B(n13937), .Z(n14016) );
  XNOR U14648 ( .A(n14017), .B(n14016), .Z(n14018) );
  XOR U14649 ( .A(n14019), .B(n14018), .Z(n14025) );
  XOR U14650 ( .A(n14024), .B(n14025), .Z(n14031) );
  XOR U14651 ( .A(n14030), .B(n14031), .Z(n14043) );
  XNOR U14652 ( .A(n14042), .B(n14043), .Z(n13974) );
  XNOR U14653 ( .A(n13975), .B(n13974), .Z(n13976) );
  XOR U14654 ( .A(n13977), .B(n13976), .Z(n14095) );
  XNOR U14655 ( .A(n14094), .B(n14095), .Z(n14096) );
  XNOR U14656 ( .A(n14097), .B(n14096), .Z(n13970) );
  XOR U14657 ( .A(n13971), .B(n13970), .Z(n13963) );
  NANDN U14658 ( .A(n13940), .B(n13939), .Z(n13944) );
  NANDN U14659 ( .A(n13942), .B(n13941), .Z(n13943) );
  AND U14660 ( .A(n13944), .B(n13943), .Z(n13962) );
  XNOR U14661 ( .A(n13963), .B(n13962), .Z(n13964) );
  NANDN U14662 ( .A(n13946), .B(n13945), .Z(n13950) );
  NAND U14663 ( .A(n13948), .B(n13947), .Z(n13949) );
  NAND U14664 ( .A(n13950), .B(n13949), .Z(n13965) );
  XNOR U14665 ( .A(n13964), .B(n13965), .Z(n13956) );
  XNOR U14666 ( .A(n13957), .B(n13956), .Z(n13958) );
  XNOR U14667 ( .A(n13959), .B(n13958), .Z(n14100) );
  XNOR U14668 ( .A(sreg[332]), .B(n14100), .Z(n14102) );
  NANDN U14669 ( .A(sreg[331]), .B(n13951), .Z(n13955) );
  NAND U14670 ( .A(n13953), .B(n13952), .Z(n13954) );
  NAND U14671 ( .A(n13955), .B(n13954), .Z(n14101) );
  XNOR U14672 ( .A(n14102), .B(n14101), .Z(c[332]) );
  NANDN U14673 ( .A(n13957), .B(n13956), .Z(n13961) );
  NANDN U14674 ( .A(n13959), .B(n13958), .Z(n13960) );
  AND U14675 ( .A(n13961), .B(n13960), .Z(n14108) );
  NANDN U14676 ( .A(n13963), .B(n13962), .Z(n13967) );
  NANDN U14677 ( .A(n13965), .B(n13964), .Z(n13966) );
  AND U14678 ( .A(n13967), .B(n13966), .Z(n14106) );
  NANDN U14679 ( .A(n13969), .B(n13968), .Z(n13973) );
  NAND U14680 ( .A(n13971), .B(n13970), .Z(n13972) );
  AND U14681 ( .A(n13973), .B(n13972), .Z(n14113) );
  NANDN U14682 ( .A(n13975), .B(n13974), .Z(n13979) );
  NANDN U14683 ( .A(n13977), .B(n13976), .Z(n13978) );
  AND U14684 ( .A(n13979), .B(n13978), .Z(n14244) );
  NANDN U14685 ( .A(n13981), .B(n13980), .Z(n13985) );
  NAND U14686 ( .A(n13983), .B(n13982), .Z(n13984) );
  AND U14687 ( .A(n13985), .B(n13984), .Z(n14243) );
  XNOR U14688 ( .A(n14244), .B(n14243), .Z(n14246) );
  NANDN U14689 ( .A(n13987), .B(n13986), .Z(n13991) );
  NANDN U14690 ( .A(n13989), .B(n13988), .Z(n13990) );
  AND U14691 ( .A(n13991), .B(n13990), .Z(n14191) );
  NAND U14692 ( .A(n38385), .B(n13992), .Z(n13994) );
  XOR U14693 ( .A(b[27]), .B(a[83]), .Z(n14135) );
  NAND U14694 ( .A(n38343), .B(n14135), .Z(n13993) );
  AND U14695 ( .A(n13994), .B(n13993), .Z(n14198) );
  NAND U14696 ( .A(n183), .B(n13995), .Z(n13997) );
  XOR U14697 ( .A(b[5]), .B(a[105]), .Z(n14138) );
  NAND U14698 ( .A(n36296), .B(n14138), .Z(n13996) );
  AND U14699 ( .A(n13997), .B(n13996), .Z(n14196) );
  NAND U14700 ( .A(n190), .B(n13998), .Z(n14000) );
  XOR U14701 ( .A(b[19]), .B(a[91]), .Z(n14141) );
  NAND U14702 ( .A(n37821), .B(n14141), .Z(n13999) );
  NAND U14703 ( .A(n14000), .B(n13999), .Z(n14195) );
  XNOR U14704 ( .A(n14196), .B(n14195), .Z(n14197) );
  XNOR U14705 ( .A(n14198), .B(n14197), .Z(n14189) );
  NAND U14706 ( .A(n38470), .B(n14001), .Z(n14003) );
  XOR U14707 ( .A(b[31]), .B(a[79]), .Z(n14144) );
  NAND U14708 ( .A(n38453), .B(n14144), .Z(n14002) );
  AND U14709 ( .A(n14003), .B(n14002), .Z(n14156) );
  NAND U14710 ( .A(n181), .B(n14004), .Z(n14006) );
  XOR U14711 ( .A(b[3]), .B(a[107]), .Z(n14147) );
  NAND U14712 ( .A(n182), .B(n14147), .Z(n14005) );
  AND U14713 ( .A(n14006), .B(n14005), .Z(n14154) );
  NAND U14714 ( .A(n189), .B(n14007), .Z(n14009) );
  XOR U14715 ( .A(b[17]), .B(a[93]), .Z(n14150) );
  NAND U14716 ( .A(n37652), .B(n14150), .Z(n14008) );
  NAND U14717 ( .A(n14009), .B(n14008), .Z(n14153) );
  XNOR U14718 ( .A(n14154), .B(n14153), .Z(n14155) );
  XOR U14719 ( .A(n14156), .B(n14155), .Z(n14190) );
  XOR U14720 ( .A(n14189), .B(n14190), .Z(n14192) );
  XOR U14721 ( .A(n14191), .B(n14192), .Z(n14124) );
  NANDN U14722 ( .A(n14011), .B(n14010), .Z(n14015) );
  NANDN U14723 ( .A(n14013), .B(n14012), .Z(n14014) );
  AND U14724 ( .A(n14015), .B(n14014), .Z(n14177) );
  NANDN U14725 ( .A(n14017), .B(n14016), .Z(n14021) );
  NANDN U14726 ( .A(n14019), .B(n14018), .Z(n14020) );
  NAND U14727 ( .A(n14021), .B(n14020), .Z(n14178) );
  XNOR U14728 ( .A(n14177), .B(n14178), .Z(n14179) );
  NANDN U14729 ( .A(n14023), .B(n14022), .Z(n14027) );
  NANDN U14730 ( .A(n14025), .B(n14024), .Z(n14026) );
  NAND U14731 ( .A(n14027), .B(n14026), .Z(n14180) );
  XNOR U14732 ( .A(n14179), .B(n14180), .Z(n14123) );
  XNOR U14733 ( .A(n14124), .B(n14123), .Z(n14126) );
  NANDN U14734 ( .A(n14029), .B(n14028), .Z(n14033) );
  NANDN U14735 ( .A(n14031), .B(n14030), .Z(n14032) );
  AND U14736 ( .A(n14033), .B(n14032), .Z(n14125) );
  XOR U14737 ( .A(n14126), .B(n14125), .Z(n14240) );
  NANDN U14738 ( .A(n14035), .B(n14034), .Z(n14039) );
  NANDN U14739 ( .A(n14037), .B(n14036), .Z(n14038) );
  AND U14740 ( .A(n14039), .B(n14038), .Z(n14237) );
  NANDN U14741 ( .A(n14041), .B(n14040), .Z(n14045) );
  NANDN U14742 ( .A(n14043), .B(n14042), .Z(n14044) );
  AND U14743 ( .A(n14045), .B(n14044), .Z(n14120) );
  NANDN U14744 ( .A(n14047), .B(n14046), .Z(n14051) );
  OR U14745 ( .A(n14049), .B(n14048), .Z(n14050) );
  AND U14746 ( .A(n14051), .B(n14050), .Z(n14118) );
  NANDN U14747 ( .A(n14053), .B(n14052), .Z(n14057) );
  NANDN U14748 ( .A(n14055), .B(n14054), .Z(n14056) );
  AND U14749 ( .A(n14057), .B(n14056), .Z(n14184) );
  NANDN U14750 ( .A(n14059), .B(n14058), .Z(n14063) );
  NANDN U14751 ( .A(n14061), .B(n14060), .Z(n14062) );
  NAND U14752 ( .A(n14063), .B(n14062), .Z(n14183) );
  XNOR U14753 ( .A(n14184), .B(n14183), .Z(n14185) );
  NAND U14754 ( .A(b[0]), .B(a[109]), .Z(n14064) );
  XNOR U14755 ( .A(b[1]), .B(n14064), .Z(n14066) );
  NANDN U14756 ( .A(b[0]), .B(a[108]), .Z(n14065) );
  NAND U14757 ( .A(n14066), .B(n14065), .Z(n14132) );
  NAND U14758 ( .A(n194), .B(n14067), .Z(n14069) );
  XOR U14759 ( .A(b[29]), .B(a[81]), .Z(n14210) );
  NAND U14760 ( .A(n38456), .B(n14210), .Z(n14068) );
  AND U14761 ( .A(n14069), .B(n14068), .Z(n14130) );
  AND U14762 ( .A(b[31]), .B(a[77]), .Z(n14129) );
  XNOR U14763 ( .A(n14130), .B(n14129), .Z(n14131) );
  XNOR U14764 ( .A(n14132), .B(n14131), .Z(n14171) );
  NAND U14765 ( .A(n38185), .B(n14070), .Z(n14072) );
  XOR U14766 ( .A(b[23]), .B(a[87]), .Z(n14213) );
  NAND U14767 ( .A(n38132), .B(n14213), .Z(n14071) );
  AND U14768 ( .A(n14072), .B(n14071), .Z(n14204) );
  NAND U14769 ( .A(n184), .B(n14073), .Z(n14075) );
  XOR U14770 ( .A(b[7]), .B(a[103]), .Z(n14216) );
  NAND U14771 ( .A(n36592), .B(n14216), .Z(n14074) );
  AND U14772 ( .A(n14075), .B(n14074), .Z(n14202) );
  NAND U14773 ( .A(n38289), .B(n14076), .Z(n14078) );
  XOR U14774 ( .A(b[25]), .B(a[85]), .Z(n14219) );
  NAND U14775 ( .A(n38247), .B(n14219), .Z(n14077) );
  NAND U14776 ( .A(n14078), .B(n14077), .Z(n14201) );
  XNOR U14777 ( .A(n14202), .B(n14201), .Z(n14203) );
  XOR U14778 ( .A(n14204), .B(n14203), .Z(n14172) );
  XNOR U14779 ( .A(n14171), .B(n14172), .Z(n14173) );
  NAND U14780 ( .A(n187), .B(n14079), .Z(n14081) );
  XOR U14781 ( .A(b[13]), .B(a[97]), .Z(n14222) );
  NAND U14782 ( .A(n37295), .B(n14222), .Z(n14080) );
  AND U14783 ( .A(n14081), .B(n14080), .Z(n14166) );
  NAND U14784 ( .A(n186), .B(n14082), .Z(n14084) );
  XOR U14785 ( .A(b[11]), .B(a[99]), .Z(n14225) );
  NAND U14786 ( .A(n37097), .B(n14225), .Z(n14083) );
  NAND U14787 ( .A(n14084), .B(n14083), .Z(n14165) );
  XNOR U14788 ( .A(n14166), .B(n14165), .Z(n14167) );
  NAND U14789 ( .A(n188), .B(n14085), .Z(n14087) );
  XOR U14790 ( .A(b[15]), .B(a[95]), .Z(n14228) );
  NAND U14791 ( .A(n37382), .B(n14228), .Z(n14086) );
  AND U14792 ( .A(n14087), .B(n14086), .Z(n14162) );
  NAND U14793 ( .A(n38064), .B(n14088), .Z(n14090) );
  XOR U14794 ( .A(b[21]), .B(a[89]), .Z(n14231) );
  NAND U14795 ( .A(n37993), .B(n14231), .Z(n14089) );
  AND U14796 ( .A(n14090), .B(n14089), .Z(n14160) );
  NAND U14797 ( .A(n185), .B(n14091), .Z(n14093) );
  XOR U14798 ( .A(b[9]), .B(a[101]), .Z(n14234) );
  NAND U14799 ( .A(n36805), .B(n14234), .Z(n14092) );
  NAND U14800 ( .A(n14093), .B(n14092), .Z(n14159) );
  XNOR U14801 ( .A(n14160), .B(n14159), .Z(n14161) );
  XOR U14802 ( .A(n14162), .B(n14161), .Z(n14168) );
  XOR U14803 ( .A(n14167), .B(n14168), .Z(n14174) );
  XOR U14804 ( .A(n14173), .B(n14174), .Z(n14186) );
  XNOR U14805 ( .A(n14185), .B(n14186), .Z(n14117) );
  XNOR U14806 ( .A(n14118), .B(n14117), .Z(n14119) );
  XOR U14807 ( .A(n14120), .B(n14119), .Z(n14238) );
  XNOR U14808 ( .A(n14237), .B(n14238), .Z(n14239) );
  XNOR U14809 ( .A(n14240), .B(n14239), .Z(n14245) );
  XOR U14810 ( .A(n14246), .B(n14245), .Z(n14112) );
  NANDN U14811 ( .A(n14095), .B(n14094), .Z(n14099) );
  NANDN U14812 ( .A(n14097), .B(n14096), .Z(n14098) );
  AND U14813 ( .A(n14099), .B(n14098), .Z(n14111) );
  XOR U14814 ( .A(n14112), .B(n14111), .Z(n14114) );
  XNOR U14815 ( .A(n14113), .B(n14114), .Z(n14105) );
  XNOR U14816 ( .A(n14106), .B(n14105), .Z(n14107) );
  XNOR U14817 ( .A(n14108), .B(n14107), .Z(n14249) );
  XNOR U14818 ( .A(sreg[333]), .B(n14249), .Z(n14251) );
  NANDN U14819 ( .A(sreg[332]), .B(n14100), .Z(n14104) );
  NAND U14820 ( .A(n14102), .B(n14101), .Z(n14103) );
  NAND U14821 ( .A(n14104), .B(n14103), .Z(n14250) );
  XNOR U14822 ( .A(n14251), .B(n14250), .Z(c[333]) );
  NANDN U14823 ( .A(n14106), .B(n14105), .Z(n14110) );
  NANDN U14824 ( .A(n14108), .B(n14107), .Z(n14109) );
  AND U14825 ( .A(n14110), .B(n14109), .Z(n14257) );
  NANDN U14826 ( .A(n14112), .B(n14111), .Z(n14116) );
  NANDN U14827 ( .A(n14114), .B(n14113), .Z(n14115) );
  AND U14828 ( .A(n14116), .B(n14115), .Z(n14255) );
  NANDN U14829 ( .A(n14118), .B(n14117), .Z(n14122) );
  NANDN U14830 ( .A(n14120), .B(n14119), .Z(n14121) );
  AND U14831 ( .A(n14122), .B(n14121), .Z(n14267) );
  NANDN U14832 ( .A(n14124), .B(n14123), .Z(n14128) );
  NAND U14833 ( .A(n14126), .B(n14125), .Z(n14127) );
  AND U14834 ( .A(n14128), .B(n14127), .Z(n14266) );
  XNOR U14835 ( .A(n14267), .B(n14266), .Z(n14269) );
  NANDN U14836 ( .A(n14130), .B(n14129), .Z(n14134) );
  NANDN U14837 ( .A(n14132), .B(n14131), .Z(n14133) );
  AND U14838 ( .A(n14134), .B(n14133), .Z(n14346) );
  NAND U14839 ( .A(n38385), .B(n14135), .Z(n14137) );
  XOR U14840 ( .A(b[27]), .B(a[84]), .Z(n14290) );
  NAND U14841 ( .A(n38343), .B(n14290), .Z(n14136) );
  AND U14842 ( .A(n14137), .B(n14136), .Z(n14353) );
  NAND U14843 ( .A(n183), .B(n14138), .Z(n14140) );
  XOR U14844 ( .A(b[5]), .B(a[106]), .Z(n14293) );
  NAND U14845 ( .A(n36296), .B(n14293), .Z(n14139) );
  AND U14846 ( .A(n14140), .B(n14139), .Z(n14351) );
  NAND U14847 ( .A(n190), .B(n14141), .Z(n14143) );
  XOR U14848 ( .A(b[19]), .B(a[92]), .Z(n14296) );
  NAND U14849 ( .A(n37821), .B(n14296), .Z(n14142) );
  NAND U14850 ( .A(n14143), .B(n14142), .Z(n14350) );
  XNOR U14851 ( .A(n14351), .B(n14350), .Z(n14352) );
  XNOR U14852 ( .A(n14353), .B(n14352), .Z(n14344) );
  NAND U14853 ( .A(n38470), .B(n14144), .Z(n14146) );
  XOR U14854 ( .A(b[31]), .B(a[80]), .Z(n14299) );
  NAND U14855 ( .A(n38453), .B(n14299), .Z(n14145) );
  AND U14856 ( .A(n14146), .B(n14145), .Z(n14311) );
  NAND U14857 ( .A(n181), .B(n14147), .Z(n14149) );
  XOR U14858 ( .A(b[3]), .B(a[108]), .Z(n14302) );
  NAND U14859 ( .A(n182), .B(n14302), .Z(n14148) );
  AND U14860 ( .A(n14149), .B(n14148), .Z(n14309) );
  NAND U14861 ( .A(n189), .B(n14150), .Z(n14152) );
  XOR U14862 ( .A(b[17]), .B(a[94]), .Z(n14305) );
  NAND U14863 ( .A(n37652), .B(n14305), .Z(n14151) );
  NAND U14864 ( .A(n14152), .B(n14151), .Z(n14308) );
  XNOR U14865 ( .A(n14309), .B(n14308), .Z(n14310) );
  XOR U14866 ( .A(n14311), .B(n14310), .Z(n14345) );
  XOR U14867 ( .A(n14344), .B(n14345), .Z(n14347) );
  XOR U14868 ( .A(n14346), .B(n14347), .Z(n14279) );
  NANDN U14869 ( .A(n14154), .B(n14153), .Z(n14158) );
  NANDN U14870 ( .A(n14156), .B(n14155), .Z(n14157) );
  AND U14871 ( .A(n14158), .B(n14157), .Z(n14332) );
  NANDN U14872 ( .A(n14160), .B(n14159), .Z(n14164) );
  NANDN U14873 ( .A(n14162), .B(n14161), .Z(n14163) );
  NAND U14874 ( .A(n14164), .B(n14163), .Z(n14333) );
  XNOR U14875 ( .A(n14332), .B(n14333), .Z(n14334) );
  NANDN U14876 ( .A(n14166), .B(n14165), .Z(n14170) );
  NANDN U14877 ( .A(n14168), .B(n14167), .Z(n14169) );
  NAND U14878 ( .A(n14170), .B(n14169), .Z(n14335) );
  XNOR U14879 ( .A(n14334), .B(n14335), .Z(n14278) );
  XNOR U14880 ( .A(n14279), .B(n14278), .Z(n14281) );
  NANDN U14881 ( .A(n14172), .B(n14171), .Z(n14176) );
  NANDN U14882 ( .A(n14174), .B(n14173), .Z(n14175) );
  AND U14883 ( .A(n14176), .B(n14175), .Z(n14280) );
  XOR U14884 ( .A(n14281), .B(n14280), .Z(n14395) );
  NANDN U14885 ( .A(n14178), .B(n14177), .Z(n14182) );
  NANDN U14886 ( .A(n14180), .B(n14179), .Z(n14181) );
  AND U14887 ( .A(n14182), .B(n14181), .Z(n14392) );
  NANDN U14888 ( .A(n14184), .B(n14183), .Z(n14188) );
  NANDN U14889 ( .A(n14186), .B(n14185), .Z(n14187) );
  AND U14890 ( .A(n14188), .B(n14187), .Z(n14275) );
  NANDN U14891 ( .A(n14190), .B(n14189), .Z(n14194) );
  OR U14892 ( .A(n14192), .B(n14191), .Z(n14193) );
  AND U14893 ( .A(n14194), .B(n14193), .Z(n14273) );
  NANDN U14894 ( .A(n14196), .B(n14195), .Z(n14200) );
  NANDN U14895 ( .A(n14198), .B(n14197), .Z(n14199) );
  AND U14896 ( .A(n14200), .B(n14199), .Z(n14339) );
  NANDN U14897 ( .A(n14202), .B(n14201), .Z(n14206) );
  NANDN U14898 ( .A(n14204), .B(n14203), .Z(n14205) );
  NAND U14899 ( .A(n14206), .B(n14205), .Z(n14338) );
  XNOR U14900 ( .A(n14339), .B(n14338), .Z(n14340) );
  NAND U14901 ( .A(b[0]), .B(a[110]), .Z(n14207) );
  XNOR U14902 ( .A(b[1]), .B(n14207), .Z(n14209) );
  NANDN U14903 ( .A(b[0]), .B(a[109]), .Z(n14208) );
  NAND U14904 ( .A(n14209), .B(n14208), .Z(n14287) );
  NAND U14905 ( .A(n194), .B(n14210), .Z(n14212) );
  XOR U14906 ( .A(b[29]), .B(a[82]), .Z(n14362) );
  NAND U14907 ( .A(n38456), .B(n14362), .Z(n14211) );
  AND U14908 ( .A(n14212), .B(n14211), .Z(n14285) );
  AND U14909 ( .A(b[31]), .B(a[78]), .Z(n14284) );
  XNOR U14910 ( .A(n14285), .B(n14284), .Z(n14286) );
  XNOR U14911 ( .A(n14287), .B(n14286), .Z(n14326) );
  NAND U14912 ( .A(n38185), .B(n14213), .Z(n14215) );
  XOR U14913 ( .A(b[23]), .B(a[88]), .Z(n14368) );
  NAND U14914 ( .A(n38132), .B(n14368), .Z(n14214) );
  AND U14915 ( .A(n14215), .B(n14214), .Z(n14359) );
  NAND U14916 ( .A(n184), .B(n14216), .Z(n14218) );
  XOR U14917 ( .A(b[7]), .B(a[104]), .Z(n14371) );
  NAND U14918 ( .A(n36592), .B(n14371), .Z(n14217) );
  AND U14919 ( .A(n14218), .B(n14217), .Z(n14357) );
  NAND U14920 ( .A(n38289), .B(n14219), .Z(n14221) );
  XOR U14921 ( .A(b[25]), .B(a[86]), .Z(n14374) );
  NAND U14922 ( .A(n38247), .B(n14374), .Z(n14220) );
  NAND U14923 ( .A(n14221), .B(n14220), .Z(n14356) );
  XNOR U14924 ( .A(n14357), .B(n14356), .Z(n14358) );
  XOR U14925 ( .A(n14359), .B(n14358), .Z(n14327) );
  XNOR U14926 ( .A(n14326), .B(n14327), .Z(n14328) );
  NAND U14927 ( .A(n187), .B(n14222), .Z(n14224) );
  XOR U14928 ( .A(b[13]), .B(a[98]), .Z(n14377) );
  NAND U14929 ( .A(n37295), .B(n14377), .Z(n14223) );
  AND U14930 ( .A(n14224), .B(n14223), .Z(n14321) );
  NAND U14931 ( .A(n186), .B(n14225), .Z(n14227) );
  XOR U14932 ( .A(b[11]), .B(a[100]), .Z(n14380) );
  NAND U14933 ( .A(n37097), .B(n14380), .Z(n14226) );
  NAND U14934 ( .A(n14227), .B(n14226), .Z(n14320) );
  XNOR U14935 ( .A(n14321), .B(n14320), .Z(n14322) );
  NAND U14936 ( .A(n188), .B(n14228), .Z(n14230) );
  XOR U14937 ( .A(b[15]), .B(a[96]), .Z(n14383) );
  NAND U14938 ( .A(n37382), .B(n14383), .Z(n14229) );
  AND U14939 ( .A(n14230), .B(n14229), .Z(n14317) );
  NAND U14940 ( .A(n38064), .B(n14231), .Z(n14233) );
  XOR U14941 ( .A(b[21]), .B(a[90]), .Z(n14386) );
  NAND U14942 ( .A(n37993), .B(n14386), .Z(n14232) );
  AND U14943 ( .A(n14233), .B(n14232), .Z(n14315) );
  NAND U14944 ( .A(n185), .B(n14234), .Z(n14236) );
  XOR U14945 ( .A(b[9]), .B(a[102]), .Z(n14389) );
  NAND U14946 ( .A(n36805), .B(n14389), .Z(n14235) );
  NAND U14947 ( .A(n14236), .B(n14235), .Z(n14314) );
  XNOR U14948 ( .A(n14315), .B(n14314), .Z(n14316) );
  XOR U14949 ( .A(n14317), .B(n14316), .Z(n14323) );
  XOR U14950 ( .A(n14322), .B(n14323), .Z(n14329) );
  XOR U14951 ( .A(n14328), .B(n14329), .Z(n14341) );
  XNOR U14952 ( .A(n14340), .B(n14341), .Z(n14272) );
  XNOR U14953 ( .A(n14273), .B(n14272), .Z(n14274) );
  XOR U14954 ( .A(n14275), .B(n14274), .Z(n14393) );
  XNOR U14955 ( .A(n14392), .B(n14393), .Z(n14394) );
  XNOR U14956 ( .A(n14395), .B(n14394), .Z(n14268) );
  XOR U14957 ( .A(n14269), .B(n14268), .Z(n14261) );
  NANDN U14958 ( .A(n14238), .B(n14237), .Z(n14242) );
  NANDN U14959 ( .A(n14240), .B(n14239), .Z(n14241) );
  AND U14960 ( .A(n14242), .B(n14241), .Z(n14260) );
  XNOR U14961 ( .A(n14261), .B(n14260), .Z(n14262) );
  NANDN U14962 ( .A(n14244), .B(n14243), .Z(n14248) );
  NAND U14963 ( .A(n14246), .B(n14245), .Z(n14247) );
  NAND U14964 ( .A(n14248), .B(n14247), .Z(n14263) );
  XNOR U14965 ( .A(n14262), .B(n14263), .Z(n14254) );
  XNOR U14966 ( .A(n14255), .B(n14254), .Z(n14256) );
  XNOR U14967 ( .A(n14257), .B(n14256), .Z(n14398) );
  XNOR U14968 ( .A(sreg[334]), .B(n14398), .Z(n14400) );
  NANDN U14969 ( .A(sreg[333]), .B(n14249), .Z(n14253) );
  NAND U14970 ( .A(n14251), .B(n14250), .Z(n14252) );
  NAND U14971 ( .A(n14253), .B(n14252), .Z(n14399) );
  XNOR U14972 ( .A(n14400), .B(n14399), .Z(c[334]) );
  NANDN U14973 ( .A(n14255), .B(n14254), .Z(n14259) );
  NANDN U14974 ( .A(n14257), .B(n14256), .Z(n14258) );
  AND U14975 ( .A(n14259), .B(n14258), .Z(n14406) );
  NANDN U14976 ( .A(n14261), .B(n14260), .Z(n14265) );
  NANDN U14977 ( .A(n14263), .B(n14262), .Z(n14264) );
  AND U14978 ( .A(n14265), .B(n14264), .Z(n14404) );
  NANDN U14979 ( .A(n14267), .B(n14266), .Z(n14271) );
  NAND U14980 ( .A(n14269), .B(n14268), .Z(n14270) );
  AND U14981 ( .A(n14271), .B(n14270), .Z(n14411) );
  NANDN U14982 ( .A(n14273), .B(n14272), .Z(n14277) );
  NANDN U14983 ( .A(n14275), .B(n14274), .Z(n14276) );
  AND U14984 ( .A(n14277), .B(n14276), .Z(n14542) );
  NANDN U14985 ( .A(n14279), .B(n14278), .Z(n14283) );
  NAND U14986 ( .A(n14281), .B(n14280), .Z(n14282) );
  AND U14987 ( .A(n14283), .B(n14282), .Z(n14541) );
  XNOR U14988 ( .A(n14542), .B(n14541), .Z(n14544) );
  NANDN U14989 ( .A(n14285), .B(n14284), .Z(n14289) );
  NANDN U14990 ( .A(n14287), .B(n14286), .Z(n14288) );
  AND U14991 ( .A(n14289), .B(n14288), .Z(n14489) );
  NAND U14992 ( .A(n38385), .B(n14290), .Z(n14292) );
  XOR U14993 ( .A(b[27]), .B(a[85]), .Z(n14433) );
  NAND U14994 ( .A(n38343), .B(n14433), .Z(n14291) );
  AND U14995 ( .A(n14292), .B(n14291), .Z(n14496) );
  NAND U14996 ( .A(n183), .B(n14293), .Z(n14295) );
  XOR U14997 ( .A(b[5]), .B(a[107]), .Z(n14436) );
  NAND U14998 ( .A(n36296), .B(n14436), .Z(n14294) );
  AND U14999 ( .A(n14295), .B(n14294), .Z(n14494) );
  NAND U15000 ( .A(n190), .B(n14296), .Z(n14298) );
  XOR U15001 ( .A(b[19]), .B(a[93]), .Z(n14439) );
  NAND U15002 ( .A(n37821), .B(n14439), .Z(n14297) );
  NAND U15003 ( .A(n14298), .B(n14297), .Z(n14493) );
  XNOR U15004 ( .A(n14494), .B(n14493), .Z(n14495) );
  XNOR U15005 ( .A(n14496), .B(n14495), .Z(n14487) );
  NAND U15006 ( .A(n38470), .B(n14299), .Z(n14301) );
  XOR U15007 ( .A(b[31]), .B(a[81]), .Z(n14442) );
  NAND U15008 ( .A(n38453), .B(n14442), .Z(n14300) );
  AND U15009 ( .A(n14301), .B(n14300), .Z(n14454) );
  NAND U15010 ( .A(n181), .B(n14302), .Z(n14304) );
  XOR U15011 ( .A(b[3]), .B(a[109]), .Z(n14445) );
  NAND U15012 ( .A(n182), .B(n14445), .Z(n14303) );
  AND U15013 ( .A(n14304), .B(n14303), .Z(n14452) );
  NAND U15014 ( .A(n189), .B(n14305), .Z(n14307) );
  XOR U15015 ( .A(b[17]), .B(a[95]), .Z(n14448) );
  NAND U15016 ( .A(n37652), .B(n14448), .Z(n14306) );
  NAND U15017 ( .A(n14307), .B(n14306), .Z(n14451) );
  XNOR U15018 ( .A(n14452), .B(n14451), .Z(n14453) );
  XOR U15019 ( .A(n14454), .B(n14453), .Z(n14488) );
  XOR U15020 ( .A(n14487), .B(n14488), .Z(n14490) );
  XOR U15021 ( .A(n14489), .B(n14490), .Z(n14422) );
  NANDN U15022 ( .A(n14309), .B(n14308), .Z(n14313) );
  NANDN U15023 ( .A(n14311), .B(n14310), .Z(n14312) );
  AND U15024 ( .A(n14313), .B(n14312), .Z(n14475) );
  NANDN U15025 ( .A(n14315), .B(n14314), .Z(n14319) );
  NANDN U15026 ( .A(n14317), .B(n14316), .Z(n14318) );
  NAND U15027 ( .A(n14319), .B(n14318), .Z(n14476) );
  XNOR U15028 ( .A(n14475), .B(n14476), .Z(n14477) );
  NANDN U15029 ( .A(n14321), .B(n14320), .Z(n14325) );
  NANDN U15030 ( .A(n14323), .B(n14322), .Z(n14324) );
  NAND U15031 ( .A(n14325), .B(n14324), .Z(n14478) );
  XNOR U15032 ( .A(n14477), .B(n14478), .Z(n14421) );
  XNOR U15033 ( .A(n14422), .B(n14421), .Z(n14424) );
  NANDN U15034 ( .A(n14327), .B(n14326), .Z(n14331) );
  NANDN U15035 ( .A(n14329), .B(n14328), .Z(n14330) );
  AND U15036 ( .A(n14331), .B(n14330), .Z(n14423) );
  XOR U15037 ( .A(n14424), .B(n14423), .Z(n14538) );
  NANDN U15038 ( .A(n14333), .B(n14332), .Z(n14337) );
  NANDN U15039 ( .A(n14335), .B(n14334), .Z(n14336) );
  AND U15040 ( .A(n14337), .B(n14336), .Z(n14535) );
  NANDN U15041 ( .A(n14339), .B(n14338), .Z(n14343) );
  NANDN U15042 ( .A(n14341), .B(n14340), .Z(n14342) );
  AND U15043 ( .A(n14343), .B(n14342), .Z(n14418) );
  NANDN U15044 ( .A(n14345), .B(n14344), .Z(n14349) );
  OR U15045 ( .A(n14347), .B(n14346), .Z(n14348) );
  AND U15046 ( .A(n14349), .B(n14348), .Z(n14416) );
  NANDN U15047 ( .A(n14351), .B(n14350), .Z(n14355) );
  NANDN U15048 ( .A(n14353), .B(n14352), .Z(n14354) );
  AND U15049 ( .A(n14355), .B(n14354), .Z(n14482) );
  NANDN U15050 ( .A(n14357), .B(n14356), .Z(n14361) );
  NANDN U15051 ( .A(n14359), .B(n14358), .Z(n14360) );
  NAND U15052 ( .A(n14361), .B(n14360), .Z(n14481) );
  XNOR U15053 ( .A(n14482), .B(n14481), .Z(n14483) );
  NAND U15054 ( .A(n194), .B(n14362), .Z(n14364) );
  XOR U15055 ( .A(b[29]), .B(a[83]), .Z(n14508) );
  NAND U15056 ( .A(n38456), .B(n14508), .Z(n14363) );
  AND U15057 ( .A(n14364), .B(n14363), .Z(n14428) );
  AND U15058 ( .A(b[31]), .B(a[79]), .Z(n14427) );
  XNOR U15059 ( .A(n14428), .B(n14427), .Z(n14429) );
  NAND U15060 ( .A(b[0]), .B(a[111]), .Z(n14365) );
  XNOR U15061 ( .A(b[1]), .B(n14365), .Z(n14367) );
  NANDN U15062 ( .A(b[0]), .B(a[110]), .Z(n14366) );
  NAND U15063 ( .A(n14367), .B(n14366), .Z(n14430) );
  XNOR U15064 ( .A(n14429), .B(n14430), .Z(n14469) );
  NAND U15065 ( .A(n38185), .B(n14368), .Z(n14370) );
  XOR U15066 ( .A(b[23]), .B(a[89]), .Z(n14511) );
  NAND U15067 ( .A(n38132), .B(n14511), .Z(n14369) );
  AND U15068 ( .A(n14370), .B(n14369), .Z(n14502) );
  NAND U15069 ( .A(n184), .B(n14371), .Z(n14373) );
  XOR U15070 ( .A(b[7]), .B(a[105]), .Z(n14514) );
  NAND U15071 ( .A(n36592), .B(n14514), .Z(n14372) );
  AND U15072 ( .A(n14373), .B(n14372), .Z(n14500) );
  NAND U15073 ( .A(n38289), .B(n14374), .Z(n14376) );
  XOR U15074 ( .A(b[25]), .B(a[87]), .Z(n14517) );
  NAND U15075 ( .A(n38247), .B(n14517), .Z(n14375) );
  NAND U15076 ( .A(n14376), .B(n14375), .Z(n14499) );
  XNOR U15077 ( .A(n14500), .B(n14499), .Z(n14501) );
  XOR U15078 ( .A(n14502), .B(n14501), .Z(n14470) );
  XNOR U15079 ( .A(n14469), .B(n14470), .Z(n14471) );
  NAND U15080 ( .A(n187), .B(n14377), .Z(n14379) );
  XOR U15081 ( .A(b[13]), .B(a[99]), .Z(n14520) );
  NAND U15082 ( .A(n37295), .B(n14520), .Z(n14378) );
  AND U15083 ( .A(n14379), .B(n14378), .Z(n14464) );
  NAND U15084 ( .A(n186), .B(n14380), .Z(n14382) );
  XOR U15085 ( .A(b[11]), .B(a[101]), .Z(n14523) );
  NAND U15086 ( .A(n37097), .B(n14523), .Z(n14381) );
  NAND U15087 ( .A(n14382), .B(n14381), .Z(n14463) );
  XNOR U15088 ( .A(n14464), .B(n14463), .Z(n14465) );
  NAND U15089 ( .A(n188), .B(n14383), .Z(n14385) );
  XOR U15090 ( .A(b[15]), .B(a[97]), .Z(n14526) );
  NAND U15091 ( .A(n37382), .B(n14526), .Z(n14384) );
  AND U15092 ( .A(n14385), .B(n14384), .Z(n14460) );
  NAND U15093 ( .A(n38064), .B(n14386), .Z(n14388) );
  XOR U15094 ( .A(b[21]), .B(a[91]), .Z(n14529) );
  NAND U15095 ( .A(n37993), .B(n14529), .Z(n14387) );
  AND U15096 ( .A(n14388), .B(n14387), .Z(n14458) );
  NAND U15097 ( .A(n185), .B(n14389), .Z(n14391) );
  XOR U15098 ( .A(b[9]), .B(a[103]), .Z(n14532) );
  NAND U15099 ( .A(n36805), .B(n14532), .Z(n14390) );
  NAND U15100 ( .A(n14391), .B(n14390), .Z(n14457) );
  XNOR U15101 ( .A(n14458), .B(n14457), .Z(n14459) );
  XOR U15102 ( .A(n14460), .B(n14459), .Z(n14466) );
  XOR U15103 ( .A(n14465), .B(n14466), .Z(n14472) );
  XOR U15104 ( .A(n14471), .B(n14472), .Z(n14484) );
  XNOR U15105 ( .A(n14483), .B(n14484), .Z(n14415) );
  XNOR U15106 ( .A(n14416), .B(n14415), .Z(n14417) );
  XOR U15107 ( .A(n14418), .B(n14417), .Z(n14536) );
  XNOR U15108 ( .A(n14535), .B(n14536), .Z(n14537) );
  XNOR U15109 ( .A(n14538), .B(n14537), .Z(n14543) );
  XOR U15110 ( .A(n14544), .B(n14543), .Z(n14410) );
  NANDN U15111 ( .A(n14393), .B(n14392), .Z(n14397) );
  NANDN U15112 ( .A(n14395), .B(n14394), .Z(n14396) );
  AND U15113 ( .A(n14397), .B(n14396), .Z(n14409) );
  XOR U15114 ( .A(n14410), .B(n14409), .Z(n14412) );
  XNOR U15115 ( .A(n14411), .B(n14412), .Z(n14403) );
  XNOR U15116 ( .A(n14404), .B(n14403), .Z(n14405) );
  XNOR U15117 ( .A(n14406), .B(n14405), .Z(n14547) );
  XNOR U15118 ( .A(sreg[335]), .B(n14547), .Z(n14549) );
  NANDN U15119 ( .A(sreg[334]), .B(n14398), .Z(n14402) );
  NAND U15120 ( .A(n14400), .B(n14399), .Z(n14401) );
  NAND U15121 ( .A(n14402), .B(n14401), .Z(n14548) );
  XNOR U15122 ( .A(n14549), .B(n14548), .Z(c[335]) );
  NANDN U15123 ( .A(n14404), .B(n14403), .Z(n14408) );
  NANDN U15124 ( .A(n14406), .B(n14405), .Z(n14407) );
  AND U15125 ( .A(n14408), .B(n14407), .Z(n14555) );
  NANDN U15126 ( .A(n14410), .B(n14409), .Z(n14414) );
  NANDN U15127 ( .A(n14412), .B(n14411), .Z(n14413) );
  AND U15128 ( .A(n14414), .B(n14413), .Z(n14553) );
  NANDN U15129 ( .A(n14416), .B(n14415), .Z(n14420) );
  NANDN U15130 ( .A(n14418), .B(n14417), .Z(n14419) );
  AND U15131 ( .A(n14420), .B(n14419), .Z(n14565) );
  NANDN U15132 ( .A(n14422), .B(n14421), .Z(n14426) );
  NAND U15133 ( .A(n14424), .B(n14423), .Z(n14425) );
  AND U15134 ( .A(n14426), .B(n14425), .Z(n14564) );
  XNOR U15135 ( .A(n14565), .B(n14564), .Z(n14567) );
  NANDN U15136 ( .A(n14428), .B(n14427), .Z(n14432) );
  NANDN U15137 ( .A(n14430), .B(n14429), .Z(n14431) );
  AND U15138 ( .A(n14432), .B(n14431), .Z(n14644) );
  NAND U15139 ( .A(n38385), .B(n14433), .Z(n14435) );
  XOR U15140 ( .A(b[27]), .B(a[86]), .Z(n14588) );
  NAND U15141 ( .A(n38343), .B(n14588), .Z(n14434) );
  AND U15142 ( .A(n14435), .B(n14434), .Z(n14651) );
  NAND U15143 ( .A(n183), .B(n14436), .Z(n14438) );
  XOR U15144 ( .A(b[5]), .B(a[108]), .Z(n14591) );
  NAND U15145 ( .A(n36296), .B(n14591), .Z(n14437) );
  AND U15146 ( .A(n14438), .B(n14437), .Z(n14649) );
  NAND U15147 ( .A(n190), .B(n14439), .Z(n14441) );
  XOR U15148 ( .A(b[19]), .B(a[94]), .Z(n14594) );
  NAND U15149 ( .A(n37821), .B(n14594), .Z(n14440) );
  NAND U15150 ( .A(n14441), .B(n14440), .Z(n14648) );
  XNOR U15151 ( .A(n14649), .B(n14648), .Z(n14650) );
  XNOR U15152 ( .A(n14651), .B(n14650), .Z(n14642) );
  NAND U15153 ( .A(n38470), .B(n14442), .Z(n14444) );
  XOR U15154 ( .A(b[31]), .B(a[82]), .Z(n14597) );
  NAND U15155 ( .A(n38453), .B(n14597), .Z(n14443) );
  AND U15156 ( .A(n14444), .B(n14443), .Z(n14609) );
  NAND U15157 ( .A(n181), .B(n14445), .Z(n14447) );
  XOR U15158 ( .A(b[3]), .B(a[110]), .Z(n14600) );
  NAND U15159 ( .A(n182), .B(n14600), .Z(n14446) );
  AND U15160 ( .A(n14447), .B(n14446), .Z(n14607) );
  NAND U15161 ( .A(n189), .B(n14448), .Z(n14450) );
  XOR U15162 ( .A(b[17]), .B(a[96]), .Z(n14603) );
  NAND U15163 ( .A(n37652), .B(n14603), .Z(n14449) );
  NAND U15164 ( .A(n14450), .B(n14449), .Z(n14606) );
  XNOR U15165 ( .A(n14607), .B(n14606), .Z(n14608) );
  XOR U15166 ( .A(n14609), .B(n14608), .Z(n14643) );
  XOR U15167 ( .A(n14642), .B(n14643), .Z(n14645) );
  XOR U15168 ( .A(n14644), .B(n14645), .Z(n14577) );
  NANDN U15169 ( .A(n14452), .B(n14451), .Z(n14456) );
  NANDN U15170 ( .A(n14454), .B(n14453), .Z(n14455) );
  AND U15171 ( .A(n14456), .B(n14455), .Z(n14630) );
  NANDN U15172 ( .A(n14458), .B(n14457), .Z(n14462) );
  NANDN U15173 ( .A(n14460), .B(n14459), .Z(n14461) );
  NAND U15174 ( .A(n14462), .B(n14461), .Z(n14631) );
  XNOR U15175 ( .A(n14630), .B(n14631), .Z(n14632) );
  NANDN U15176 ( .A(n14464), .B(n14463), .Z(n14468) );
  NANDN U15177 ( .A(n14466), .B(n14465), .Z(n14467) );
  NAND U15178 ( .A(n14468), .B(n14467), .Z(n14633) );
  XNOR U15179 ( .A(n14632), .B(n14633), .Z(n14576) );
  XNOR U15180 ( .A(n14577), .B(n14576), .Z(n14579) );
  NANDN U15181 ( .A(n14470), .B(n14469), .Z(n14474) );
  NANDN U15182 ( .A(n14472), .B(n14471), .Z(n14473) );
  AND U15183 ( .A(n14474), .B(n14473), .Z(n14578) );
  XOR U15184 ( .A(n14579), .B(n14578), .Z(n14693) );
  NANDN U15185 ( .A(n14476), .B(n14475), .Z(n14480) );
  NANDN U15186 ( .A(n14478), .B(n14477), .Z(n14479) );
  AND U15187 ( .A(n14480), .B(n14479), .Z(n14690) );
  NANDN U15188 ( .A(n14482), .B(n14481), .Z(n14486) );
  NANDN U15189 ( .A(n14484), .B(n14483), .Z(n14485) );
  AND U15190 ( .A(n14486), .B(n14485), .Z(n14573) );
  NANDN U15191 ( .A(n14488), .B(n14487), .Z(n14492) );
  OR U15192 ( .A(n14490), .B(n14489), .Z(n14491) );
  AND U15193 ( .A(n14492), .B(n14491), .Z(n14571) );
  NANDN U15194 ( .A(n14494), .B(n14493), .Z(n14498) );
  NANDN U15195 ( .A(n14496), .B(n14495), .Z(n14497) );
  AND U15196 ( .A(n14498), .B(n14497), .Z(n14637) );
  NANDN U15197 ( .A(n14500), .B(n14499), .Z(n14504) );
  NANDN U15198 ( .A(n14502), .B(n14501), .Z(n14503) );
  NAND U15199 ( .A(n14504), .B(n14503), .Z(n14636) );
  XNOR U15200 ( .A(n14637), .B(n14636), .Z(n14638) );
  NAND U15201 ( .A(b[0]), .B(a[112]), .Z(n14505) );
  XNOR U15202 ( .A(b[1]), .B(n14505), .Z(n14507) );
  NANDN U15203 ( .A(b[0]), .B(a[111]), .Z(n14506) );
  NAND U15204 ( .A(n14507), .B(n14506), .Z(n14585) );
  NAND U15205 ( .A(n194), .B(n14508), .Z(n14510) );
  XOR U15206 ( .A(b[29]), .B(a[84]), .Z(n14663) );
  NAND U15207 ( .A(n38456), .B(n14663), .Z(n14509) );
  AND U15208 ( .A(n14510), .B(n14509), .Z(n14583) );
  AND U15209 ( .A(b[31]), .B(a[80]), .Z(n14582) );
  XNOR U15210 ( .A(n14583), .B(n14582), .Z(n14584) );
  XNOR U15211 ( .A(n14585), .B(n14584), .Z(n14624) );
  NAND U15212 ( .A(n38185), .B(n14511), .Z(n14513) );
  XOR U15213 ( .A(b[23]), .B(a[90]), .Z(n14666) );
  NAND U15214 ( .A(n38132), .B(n14666), .Z(n14512) );
  AND U15215 ( .A(n14513), .B(n14512), .Z(n14657) );
  NAND U15216 ( .A(n184), .B(n14514), .Z(n14516) );
  XOR U15217 ( .A(b[7]), .B(a[106]), .Z(n14669) );
  NAND U15218 ( .A(n36592), .B(n14669), .Z(n14515) );
  AND U15219 ( .A(n14516), .B(n14515), .Z(n14655) );
  NAND U15220 ( .A(n38289), .B(n14517), .Z(n14519) );
  XOR U15221 ( .A(b[25]), .B(a[88]), .Z(n14672) );
  NAND U15222 ( .A(n38247), .B(n14672), .Z(n14518) );
  NAND U15223 ( .A(n14519), .B(n14518), .Z(n14654) );
  XNOR U15224 ( .A(n14655), .B(n14654), .Z(n14656) );
  XOR U15225 ( .A(n14657), .B(n14656), .Z(n14625) );
  XNOR U15226 ( .A(n14624), .B(n14625), .Z(n14626) );
  NAND U15227 ( .A(n187), .B(n14520), .Z(n14522) );
  XOR U15228 ( .A(b[13]), .B(a[100]), .Z(n14675) );
  NAND U15229 ( .A(n37295), .B(n14675), .Z(n14521) );
  AND U15230 ( .A(n14522), .B(n14521), .Z(n14619) );
  NAND U15231 ( .A(n186), .B(n14523), .Z(n14525) );
  XOR U15232 ( .A(b[11]), .B(a[102]), .Z(n14678) );
  NAND U15233 ( .A(n37097), .B(n14678), .Z(n14524) );
  NAND U15234 ( .A(n14525), .B(n14524), .Z(n14618) );
  XNOR U15235 ( .A(n14619), .B(n14618), .Z(n14620) );
  NAND U15236 ( .A(n188), .B(n14526), .Z(n14528) );
  XOR U15237 ( .A(b[15]), .B(a[98]), .Z(n14681) );
  NAND U15238 ( .A(n37382), .B(n14681), .Z(n14527) );
  AND U15239 ( .A(n14528), .B(n14527), .Z(n14615) );
  NAND U15240 ( .A(n38064), .B(n14529), .Z(n14531) );
  XOR U15241 ( .A(b[21]), .B(a[92]), .Z(n14684) );
  NAND U15242 ( .A(n37993), .B(n14684), .Z(n14530) );
  AND U15243 ( .A(n14531), .B(n14530), .Z(n14613) );
  NAND U15244 ( .A(n185), .B(n14532), .Z(n14534) );
  XOR U15245 ( .A(b[9]), .B(a[104]), .Z(n14687) );
  NAND U15246 ( .A(n36805), .B(n14687), .Z(n14533) );
  NAND U15247 ( .A(n14534), .B(n14533), .Z(n14612) );
  XNOR U15248 ( .A(n14613), .B(n14612), .Z(n14614) );
  XOR U15249 ( .A(n14615), .B(n14614), .Z(n14621) );
  XOR U15250 ( .A(n14620), .B(n14621), .Z(n14627) );
  XOR U15251 ( .A(n14626), .B(n14627), .Z(n14639) );
  XNOR U15252 ( .A(n14638), .B(n14639), .Z(n14570) );
  XNOR U15253 ( .A(n14571), .B(n14570), .Z(n14572) );
  XOR U15254 ( .A(n14573), .B(n14572), .Z(n14691) );
  XNOR U15255 ( .A(n14690), .B(n14691), .Z(n14692) );
  XNOR U15256 ( .A(n14693), .B(n14692), .Z(n14566) );
  XOR U15257 ( .A(n14567), .B(n14566), .Z(n14559) );
  NANDN U15258 ( .A(n14536), .B(n14535), .Z(n14540) );
  NANDN U15259 ( .A(n14538), .B(n14537), .Z(n14539) );
  AND U15260 ( .A(n14540), .B(n14539), .Z(n14558) );
  XNOR U15261 ( .A(n14559), .B(n14558), .Z(n14560) );
  NANDN U15262 ( .A(n14542), .B(n14541), .Z(n14546) );
  NAND U15263 ( .A(n14544), .B(n14543), .Z(n14545) );
  NAND U15264 ( .A(n14546), .B(n14545), .Z(n14561) );
  XNOR U15265 ( .A(n14560), .B(n14561), .Z(n14552) );
  XNOR U15266 ( .A(n14553), .B(n14552), .Z(n14554) );
  XNOR U15267 ( .A(n14555), .B(n14554), .Z(n14696) );
  XNOR U15268 ( .A(sreg[336]), .B(n14696), .Z(n14698) );
  NANDN U15269 ( .A(sreg[335]), .B(n14547), .Z(n14551) );
  NAND U15270 ( .A(n14549), .B(n14548), .Z(n14550) );
  NAND U15271 ( .A(n14551), .B(n14550), .Z(n14697) );
  XNOR U15272 ( .A(n14698), .B(n14697), .Z(c[336]) );
  NANDN U15273 ( .A(n14553), .B(n14552), .Z(n14557) );
  NANDN U15274 ( .A(n14555), .B(n14554), .Z(n14556) );
  AND U15275 ( .A(n14557), .B(n14556), .Z(n14704) );
  NANDN U15276 ( .A(n14559), .B(n14558), .Z(n14563) );
  NANDN U15277 ( .A(n14561), .B(n14560), .Z(n14562) );
  AND U15278 ( .A(n14563), .B(n14562), .Z(n14702) );
  NANDN U15279 ( .A(n14565), .B(n14564), .Z(n14569) );
  NAND U15280 ( .A(n14567), .B(n14566), .Z(n14568) );
  AND U15281 ( .A(n14569), .B(n14568), .Z(n14709) );
  NANDN U15282 ( .A(n14571), .B(n14570), .Z(n14575) );
  NANDN U15283 ( .A(n14573), .B(n14572), .Z(n14574) );
  AND U15284 ( .A(n14575), .B(n14574), .Z(n14714) );
  NANDN U15285 ( .A(n14577), .B(n14576), .Z(n14581) );
  NAND U15286 ( .A(n14579), .B(n14578), .Z(n14580) );
  AND U15287 ( .A(n14581), .B(n14580), .Z(n14713) );
  XNOR U15288 ( .A(n14714), .B(n14713), .Z(n14716) );
  NANDN U15289 ( .A(n14583), .B(n14582), .Z(n14587) );
  NANDN U15290 ( .A(n14585), .B(n14584), .Z(n14586) );
  AND U15291 ( .A(n14587), .B(n14586), .Z(n14793) );
  NAND U15292 ( .A(n38385), .B(n14588), .Z(n14590) );
  XOR U15293 ( .A(b[27]), .B(a[87]), .Z(n14737) );
  NAND U15294 ( .A(n38343), .B(n14737), .Z(n14589) );
  AND U15295 ( .A(n14590), .B(n14589), .Z(n14800) );
  NAND U15296 ( .A(n183), .B(n14591), .Z(n14593) );
  XOR U15297 ( .A(b[5]), .B(a[109]), .Z(n14740) );
  NAND U15298 ( .A(n36296), .B(n14740), .Z(n14592) );
  AND U15299 ( .A(n14593), .B(n14592), .Z(n14798) );
  NAND U15300 ( .A(n190), .B(n14594), .Z(n14596) );
  XOR U15301 ( .A(b[19]), .B(a[95]), .Z(n14743) );
  NAND U15302 ( .A(n37821), .B(n14743), .Z(n14595) );
  NAND U15303 ( .A(n14596), .B(n14595), .Z(n14797) );
  XNOR U15304 ( .A(n14798), .B(n14797), .Z(n14799) );
  XNOR U15305 ( .A(n14800), .B(n14799), .Z(n14791) );
  NAND U15306 ( .A(n38470), .B(n14597), .Z(n14599) );
  XOR U15307 ( .A(b[31]), .B(a[83]), .Z(n14746) );
  NAND U15308 ( .A(n38453), .B(n14746), .Z(n14598) );
  AND U15309 ( .A(n14599), .B(n14598), .Z(n14758) );
  NAND U15310 ( .A(n181), .B(n14600), .Z(n14602) );
  XOR U15311 ( .A(b[3]), .B(a[111]), .Z(n14749) );
  NAND U15312 ( .A(n182), .B(n14749), .Z(n14601) );
  AND U15313 ( .A(n14602), .B(n14601), .Z(n14756) );
  NAND U15314 ( .A(n189), .B(n14603), .Z(n14605) );
  XOR U15315 ( .A(b[17]), .B(a[97]), .Z(n14752) );
  NAND U15316 ( .A(n37652), .B(n14752), .Z(n14604) );
  NAND U15317 ( .A(n14605), .B(n14604), .Z(n14755) );
  XNOR U15318 ( .A(n14756), .B(n14755), .Z(n14757) );
  XOR U15319 ( .A(n14758), .B(n14757), .Z(n14792) );
  XOR U15320 ( .A(n14791), .B(n14792), .Z(n14794) );
  XOR U15321 ( .A(n14793), .B(n14794), .Z(n14726) );
  NANDN U15322 ( .A(n14607), .B(n14606), .Z(n14611) );
  NANDN U15323 ( .A(n14609), .B(n14608), .Z(n14610) );
  AND U15324 ( .A(n14611), .B(n14610), .Z(n14779) );
  NANDN U15325 ( .A(n14613), .B(n14612), .Z(n14617) );
  NANDN U15326 ( .A(n14615), .B(n14614), .Z(n14616) );
  NAND U15327 ( .A(n14617), .B(n14616), .Z(n14780) );
  XNOR U15328 ( .A(n14779), .B(n14780), .Z(n14781) );
  NANDN U15329 ( .A(n14619), .B(n14618), .Z(n14623) );
  NANDN U15330 ( .A(n14621), .B(n14620), .Z(n14622) );
  NAND U15331 ( .A(n14623), .B(n14622), .Z(n14782) );
  XNOR U15332 ( .A(n14781), .B(n14782), .Z(n14725) );
  XNOR U15333 ( .A(n14726), .B(n14725), .Z(n14728) );
  NANDN U15334 ( .A(n14625), .B(n14624), .Z(n14629) );
  NANDN U15335 ( .A(n14627), .B(n14626), .Z(n14628) );
  AND U15336 ( .A(n14629), .B(n14628), .Z(n14727) );
  XOR U15337 ( .A(n14728), .B(n14727), .Z(n14842) );
  NANDN U15338 ( .A(n14631), .B(n14630), .Z(n14635) );
  NANDN U15339 ( .A(n14633), .B(n14632), .Z(n14634) );
  AND U15340 ( .A(n14635), .B(n14634), .Z(n14839) );
  NANDN U15341 ( .A(n14637), .B(n14636), .Z(n14641) );
  NANDN U15342 ( .A(n14639), .B(n14638), .Z(n14640) );
  AND U15343 ( .A(n14641), .B(n14640), .Z(n14722) );
  NANDN U15344 ( .A(n14643), .B(n14642), .Z(n14647) );
  OR U15345 ( .A(n14645), .B(n14644), .Z(n14646) );
  AND U15346 ( .A(n14647), .B(n14646), .Z(n14720) );
  NANDN U15347 ( .A(n14649), .B(n14648), .Z(n14653) );
  NANDN U15348 ( .A(n14651), .B(n14650), .Z(n14652) );
  AND U15349 ( .A(n14653), .B(n14652), .Z(n14786) );
  NANDN U15350 ( .A(n14655), .B(n14654), .Z(n14659) );
  NANDN U15351 ( .A(n14657), .B(n14656), .Z(n14658) );
  NAND U15352 ( .A(n14659), .B(n14658), .Z(n14785) );
  XNOR U15353 ( .A(n14786), .B(n14785), .Z(n14787) );
  NAND U15354 ( .A(b[0]), .B(a[113]), .Z(n14660) );
  XNOR U15355 ( .A(b[1]), .B(n14660), .Z(n14662) );
  NANDN U15356 ( .A(b[0]), .B(a[112]), .Z(n14661) );
  NAND U15357 ( .A(n14662), .B(n14661), .Z(n14734) );
  NAND U15358 ( .A(n194), .B(n14663), .Z(n14665) );
  XOR U15359 ( .A(b[29]), .B(a[85]), .Z(n14812) );
  NAND U15360 ( .A(n38456), .B(n14812), .Z(n14664) );
  AND U15361 ( .A(n14665), .B(n14664), .Z(n14732) );
  AND U15362 ( .A(b[31]), .B(a[81]), .Z(n14731) );
  XNOR U15363 ( .A(n14732), .B(n14731), .Z(n14733) );
  XNOR U15364 ( .A(n14734), .B(n14733), .Z(n14773) );
  NAND U15365 ( .A(n38185), .B(n14666), .Z(n14668) );
  XOR U15366 ( .A(b[23]), .B(a[91]), .Z(n14815) );
  NAND U15367 ( .A(n38132), .B(n14815), .Z(n14667) );
  AND U15368 ( .A(n14668), .B(n14667), .Z(n14806) );
  NAND U15369 ( .A(n184), .B(n14669), .Z(n14671) );
  XOR U15370 ( .A(b[7]), .B(a[107]), .Z(n14818) );
  NAND U15371 ( .A(n36592), .B(n14818), .Z(n14670) );
  AND U15372 ( .A(n14671), .B(n14670), .Z(n14804) );
  NAND U15373 ( .A(n38289), .B(n14672), .Z(n14674) );
  XOR U15374 ( .A(b[25]), .B(a[89]), .Z(n14821) );
  NAND U15375 ( .A(n38247), .B(n14821), .Z(n14673) );
  NAND U15376 ( .A(n14674), .B(n14673), .Z(n14803) );
  XNOR U15377 ( .A(n14804), .B(n14803), .Z(n14805) );
  XOR U15378 ( .A(n14806), .B(n14805), .Z(n14774) );
  XNOR U15379 ( .A(n14773), .B(n14774), .Z(n14775) );
  NAND U15380 ( .A(n187), .B(n14675), .Z(n14677) );
  XOR U15381 ( .A(b[13]), .B(a[101]), .Z(n14824) );
  NAND U15382 ( .A(n37295), .B(n14824), .Z(n14676) );
  AND U15383 ( .A(n14677), .B(n14676), .Z(n14768) );
  NAND U15384 ( .A(n186), .B(n14678), .Z(n14680) );
  XOR U15385 ( .A(b[11]), .B(a[103]), .Z(n14827) );
  NAND U15386 ( .A(n37097), .B(n14827), .Z(n14679) );
  NAND U15387 ( .A(n14680), .B(n14679), .Z(n14767) );
  XNOR U15388 ( .A(n14768), .B(n14767), .Z(n14769) );
  NAND U15389 ( .A(n188), .B(n14681), .Z(n14683) );
  XOR U15390 ( .A(b[15]), .B(a[99]), .Z(n14830) );
  NAND U15391 ( .A(n37382), .B(n14830), .Z(n14682) );
  AND U15392 ( .A(n14683), .B(n14682), .Z(n14764) );
  NAND U15393 ( .A(n38064), .B(n14684), .Z(n14686) );
  XOR U15394 ( .A(b[21]), .B(a[93]), .Z(n14833) );
  NAND U15395 ( .A(n37993), .B(n14833), .Z(n14685) );
  AND U15396 ( .A(n14686), .B(n14685), .Z(n14762) );
  NAND U15397 ( .A(n185), .B(n14687), .Z(n14689) );
  XOR U15398 ( .A(b[9]), .B(a[105]), .Z(n14836) );
  NAND U15399 ( .A(n36805), .B(n14836), .Z(n14688) );
  NAND U15400 ( .A(n14689), .B(n14688), .Z(n14761) );
  XNOR U15401 ( .A(n14762), .B(n14761), .Z(n14763) );
  XOR U15402 ( .A(n14764), .B(n14763), .Z(n14770) );
  XOR U15403 ( .A(n14769), .B(n14770), .Z(n14776) );
  XOR U15404 ( .A(n14775), .B(n14776), .Z(n14788) );
  XNOR U15405 ( .A(n14787), .B(n14788), .Z(n14719) );
  XNOR U15406 ( .A(n14720), .B(n14719), .Z(n14721) );
  XOR U15407 ( .A(n14722), .B(n14721), .Z(n14840) );
  XNOR U15408 ( .A(n14839), .B(n14840), .Z(n14841) );
  XNOR U15409 ( .A(n14842), .B(n14841), .Z(n14715) );
  XOR U15410 ( .A(n14716), .B(n14715), .Z(n14708) );
  NANDN U15411 ( .A(n14691), .B(n14690), .Z(n14695) );
  NANDN U15412 ( .A(n14693), .B(n14692), .Z(n14694) );
  AND U15413 ( .A(n14695), .B(n14694), .Z(n14707) );
  XOR U15414 ( .A(n14708), .B(n14707), .Z(n14710) );
  XNOR U15415 ( .A(n14709), .B(n14710), .Z(n14701) );
  XNOR U15416 ( .A(n14702), .B(n14701), .Z(n14703) );
  XNOR U15417 ( .A(n14704), .B(n14703), .Z(n14845) );
  XNOR U15418 ( .A(sreg[337]), .B(n14845), .Z(n14847) );
  NANDN U15419 ( .A(sreg[336]), .B(n14696), .Z(n14700) );
  NAND U15420 ( .A(n14698), .B(n14697), .Z(n14699) );
  NAND U15421 ( .A(n14700), .B(n14699), .Z(n14846) );
  XNOR U15422 ( .A(n14847), .B(n14846), .Z(c[337]) );
  NANDN U15423 ( .A(n14702), .B(n14701), .Z(n14706) );
  NANDN U15424 ( .A(n14704), .B(n14703), .Z(n14705) );
  AND U15425 ( .A(n14706), .B(n14705), .Z(n14853) );
  NANDN U15426 ( .A(n14708), .B(n14707), .Z(n14712) );
  NANDN U15427 ( .A(n14710), .B(n14709), .Z(n14711) );
  AND U15428 ( .A(n14712), .B(n14711), .Z(n14851) );
  NANDN U15429 ( .A(n14714), .B(n14713), .Z(n14718) );
  NAND U15430 ( .A(n14716), .B(n14715), .Z(n14717) );
  AND U15431 ( .A(n14718), .B(n14717), .Z(n14858) );
  NANDN U15432 ( .A(n14720), .B(n14719), .Z(n14724) );
  NANDN U15433 ( .A(n14722), .B(n14721), .Z(n14723) );
  AND U15434 ( .A(n14724), .B(n14723), .Z(n14989) );
  NANDN U15435 ( .A(n14726), .B(n14725), .Z(n14730) );
  NAND U15436 ( .A(n14728), .B(n14727), .Z(n14729) );
  AND U15437 ( .A(n14730), .B(n14729), .Z(n14988) );
  XNOR U15438 ( .A(n14989), .B(n14988), .Z(n14991) );
  NANDN U15439 ( .A(n14732), .B(n14731), .Z(n14736) );
  NANDN U15440 ( .A(n14734), .B(n14733), .Z(n14735) );
  AND U15441 ( .A(n14736), .B(n14735), .Z(n14936) );
  NAND U15442 ( .A(n38385), .B(n14737), .Z(n14739) );
  XOR U15443 ( .A(b[27]), .B(a[88]), .Z(n14880) );
  NAND U15444 ( .A(n38343), .B(n14880), .Z(n14738) );
  AND U15445 ( .A(n14739), .B(n14738), .Z(n14943) );
  NAND U15446 ( .A(n183), .B(n14740), .Z(n14742) );
  XOR U15447 ( .A(b[5]), .B(a[110]), .Z(n14883) );
  NAND U15448 ( .A(n36296), .B(n14883), .Z(n14741) );
  AND U15449 ( .A(n14742), .B(n14741), .Z(n14941) );
  NAND U15450 ( .A(n190), .B(n14743), .Z(n14745) );
  XOR U15451 ( .A(b[19]), .B(a[96]), .Z(n14886) );
  NAND U15452 ( .A(n37821), .B(n14886), .Z(n14744) );
  NAND U15453 ( .A(n14745), .B(n14744), .Z(n14940) );
  XNOR U15454 ( .A(n14941), .B(n14940), .Z(n14942) );
  XNOR U15455 ( .A(n14943), .B(n14942), .Z(n14934) );
  NAND U15456 ( .A(n38470), .B(n14746), .Z(n14748) );
  XOR U15457 ( .A(b[31]), .B(a[84]), .Z(n14889) );
  NAND U15458 ( .A(n38453), .B(n14889), .Z(n14747) );
  AND U15459 ( .A(n14748), .B(n14747), .Z(n14901) );
  NAND U15460 ( .A(n181), .B(n14749), .Z(n14751) );
  XOR U15461 ( .A(b[3]), .B(a[112]), .Z(n14892) );
  NAND U15462 ( .A(n182), .B(n14892), .Z(n14750) );
  AND U15463 ( .A(n14751), .B(n14750), .Z(n14899) );
  NAND U15464 ( .A(n189), .B(n14752), .Z(n14754) );
  XOR U15465 ( .A(b[17]), .B(a[98]), .Z(n14895) );
  NAND U15466 ( .A(n37652), .B(n14895), .Z(n14753) );
  NAND U15467 ( .A(n14754), .B(n14753), .Z(n14898) );
  XNOR U15468 ( .A(n14899), .B(n14898), .Z(n14900) );
  XOR U15469 ( .A(n14901), .B(n14900), .Z(n14935) );
  XOR U15470 ( .A(n14934), .B(n14935), .Z(n14937) );
  XOR U15471 ( .A(n14936), .B(n14937), .Z(n14869) );
  NANDN U15472 ( .A(n14756), .B(n14755), .Z(n14760) );
  NANDN U15473 ( .A(n14758), .B(n14757), .Z(n14759) );
  AND U15474 ( .A(n14760), .B(n14759), .Z(n14922) );
  NANDN U15475 ( .A(n14762), .B(n14761), .Z(n14766) );
  NANDN U15476 ( .A(n14764), .B(n14763), .Z(n14765) );
  NAND U15477 ( .A(n14766), .B(n14765), .Z(n14923) );
  XNOR U15478 ( .A(n14922), .B(n14923), .Z(n14924) );
  NANDN U15479 ( .A(n14768), .B(n14767), .Z(n14772) );
  NANDN U15480 ( .A(n14770), .B(n14769), .Z(n14771) );
  NAND U15481 ( .A(n14772), .B(n14771), .Z(n14925) );
  XNOR U15482 ( .A(n14924), .B(n14925), .Z(n14868) );
  XNOR U15483 ( .A(n14869), .B(n14868), .Z(n14871) );
  NANDN U15484 ( .A(n14774), .B(n14773), .Z(n14778) );
  NANDN U15485 ( .A(n14776), .B(n14775), .Z(n14777) );
  AND U15486 ( .A(n14778), .B(n14777), .Z(n14870) );
  XOR U15487 ( .A(n14871), .B(n14870), .Z(n14985) );
  NANDN U15488 ( .A(n14780), .B(n14779), .Z(n14784) );
  NANDN U15489 ( .A(n14782), .B(n14781), .Z(n14783) );
  AND U15490 ( .A(n14784), .B(n14783), .Z(n14982) );
  NANDN U15491 ( .A(n14786), .B(n14785), .Z(n14790) );
  NANDN U15492 ( .A(n14788), .B(n14787), .Z(n14789) );
  AND U15493 ( .A(n14790), .B(n14789), .Z(n14865) );
  NANDN U15494 ( .A(n14792), .B(n14791), .Z(n14796) );
  OR U15495 ( .A(n14794), .B(n14793), .Z(n14795) );
  AND U15496 ( .A(n14796), .B(n14795), .Z(n14863) );
  NANDN U15497 ( .A(n14798), .B(n14797), .Z(n14802) );
  NANDN U15498 ( .A(n14800), .B(n14799), .Z(n14801) );
  AND U15499 ( .A(n14802), .B(n14801), .Z(n14929) );
  NANDN U15500 ( .A(n14804), .B(n14803), .Z(n14808) );
  NANDN U15501 ( .A(n14806), .B(n14805), .Z(n14807) );
  NAND U15502 ( .A(n14808), .B(n14807), .Z(n14928) );
  XNOR U15503 ( .A(n14929), .B(n14928), .Z(n14930) );
  NAND U15504 ( .A(b[0]), .B(a[114]), .Z(n14809) );
  XNOR U15505 ( .A(b[1]), .B(n14809), .Z(n14811) );
  NANDN U15506 ( .A(b[0]), .B(a[113]), .Z(n14810) );
  NAND U15507 ( .A(n14811), .B(n14810), .Z(n14877) );
  NAND U15508 ( .A(n194), .B(n14812), .Z(n14814) );
  XOR U15509 ( .A(b[29]), .B(a[86]), .Z(n14955) );
  NAND U15510 ( .A(n38456), .B(n14955), .Z(n14813) );
  AND U15511 ( .A(n14814), .B(n14813), .Z(n14875) );
  AND U15512 ( .A(b[31]), .B(a[82]), .Z(n14874) );
  XNOR U15513 ( .A(n14875), .B(n14874), .Z(n14876) );
  XNOR U15514 ( .A(n14877), .B(n14876), .Z(n14916) );
  NAND U15515 ( .A(n38185), .B(n14815), .Z(n14817) );
  XOR U15516 ( .A(b[23]), .B(a[92]), .Z(n14958) );
  NAND U15517 ( .A(n38132), .B(n14958), .Z(n14816) );
  AND U15518 ( .A(n14817), .B(n14816), .Z(n14949) );
  NAND U15519 ( .A(n184), .B(n14818), .Z(n14820) );
  XOR U15520 ( .A(b[7]), .B(a[108]), .Z(n14961) );
  NAND U15521 ( .A(n36592), .B(n14961), .Z(n14819) );
  AND U15522 ( .A(n14820), .B(n14819), .Z(n14947) );
  NAND U15523 ( .A(n38289), .B(n14821), .Z(n14823) );
  XOR U15524 ( .A(b[25]), .B(a[90]), .Z(n14964) );
  NAND U15525 ( .A(n38247), .B(n14964), .Z(n14822) );
  NAND U15526 ( .A(n14823), .B(n14822), .Z(n14946) );
  XNOR U15527 ( .A(n14947), .B(n14946), .Z(n14948) );
  XOR U15528 ( .A(n14949), .B(n14948), .Z(n14917) );
  XNOR U15529 ( .A(n14916), .B(n14917), .Z(n14918) );
  NAND U15530 ( .A(n187), .B(n14824), .Z(n14826) );
  XOR U15531 ( .A(b[13]), .B(a[102]), .Z(n14967) );
  NAND U15532 ( .A(n37295), .B(n14967), .Z(n14825) );
  AND U15533 ( .A(n14826), .B(n14825), .Z(n14911) );
  NAND U15534 ( .A(n186), .B(n14827), .Z(n14829) );
  XOR U15535 ( .A(b[11]), .B(a[104]), .Z(n14970) );
  NAND U15536 ( .A(n37097), .B(n14970), .Z(n14828) );
  NAND U15537 ( .A(n14829), .B(n14828), .Z(n14910) );
  XNOR U15538 ( .A(n14911), .B(n14910), .Z(n14912) );
  NAND U15539 ( .A(n188), .B(n14830), .Z(n14832) );
  XOR U15540 ( .A(b[15]), .B(a[100]), .Z(n14973) );
  NAND U15541 ( .A(n37382), .B(n14973), .Z(n14831) );
  AND U15542 ( .A(n14832), .B(n14831), .Z(n14907) );
  NAND U15543 ( .A(n38064), .B(n14833), .Z(n14835) );
  XOR U15544 ( .A(b[21]), .B(a[94]), .Z(n14976) );
  NAND U15545 ( .A(n37993), .B(n14976), .Z(n14834) );
  AND U15546 ( .A(n14835), .B(n14834), .Z(n14905) );
  NAND U15547 ( .A(n185), .B(n14836), .Z(n14838) );
  XOR U15548 ( .A(b[9]), .B(a[106]), .Z(n14979) );
  NAND U15549 ( .A(n36805), .B(n14979), .Z(n14837) );
  NAND U15550 ( .A(n14838), .B(n14837), .Z(n14904) );
  XNOR U15551 ( .A(n14905), .B(n14904), .Z(n14906) );
  XOR U15552 ( .A(n14907), .B(n14906), .Z(n14913) );
  XOR U15553 ( .A(n14912), .B(n14913), .Z(n14919) );
  XOR U15554 ( .A(n14918), .B(n14919), .Z(n14931) );
  XNOR U15555 ( .A(n14930), .B(n14931), .Z(n14862) );
  XNOR U15556 ( .A(n14863), .B(n14862), .Z(n14864) );
  XOR U15557 ( .A(n14865), .B(n14864), .Z(n14983) );
  XNOR U15558 ( .A(n14982), .B(n14983), .Z(n14984) );
  XNOR U15559 ( .A(n14985), .B(n14984), .Z(n14990) );
  XOR U15560 ( .A(n14991), .B(n14990), .Z(n14857) );
  NANDN U15561 ( .A(n14840), .B(n14839), .Z(n14844) );
  NANDN U15562 ( .A(n14842), .B(n14841), .Z(n14843) );
  AND U15563 ( .A(n14844), .B(n14843), .Z(n14856) );
  XOR U15564 ( .A(n14857), .B(n14856), .Z(n14859) );
  XNOR U15565 ( .A(n14858), .B(n14859), .Z(n14850) );
  XNOR U15566 ( .A(n14851), .B(n14850), .Z(n14852) );
  XNOR U15567 ( .A(n14853), .B(n14852), .Z(n14994) );
  XNOR U15568 ( .A(sreg[338]), .B(n14994), .Z(n14996) );
  NANDN U15569 ( .A(sreg[337]), .B(n14845), .Z(n14849) );
  NAND U15570 ( .A(n14847), .B(n14846), .Z(n14848) );
  NAND U15571 ( .A(n14849), .B(n14848), .Z(n14995) );
  XNOR U15572 ( .A(n14996), .B(n14995), .Z(c[338]) );
  NANDN U15573 ( .A(n14851), .B(n14850), .Z(n14855) );
  NANDN U15574 ( .A(n14853), .B(n14852), .Z(n14854) );
  AND U15575 ( .A(n14855), .B(n14854), .Z(n15002) );
  NANDN U15576 ( .A(n14857), .B(n14856), .Z(n14861) );
  NANDN U15577 ( .A(n14859), .B(n14858), .Z(n14860) );
  AND U15578 ( .A(n14861), .B(n14860), .Z(n15000) );
  NANDN U15579 ( .A(n14863), .B(n14862), .Z(n14867) );
  NANDN U15580 ( .A(n14865), .B(n14864), .Z(n14866) );
  AND U15581 ( .A(n14867), .B(n14866), .Z(n15138) );
  NANDN U15582 ( .A(n14869), .B(n14868), .Z(n14873) );
  NAND U15583 ( .A(n14871), .B(n14870), .Z(n14872) );
  AND U15584 ( .A(n14873), .B(n14872), .Z(n15137) );
  XNOR U15585 ( .A(n15138), .B(n15137), .Z(n15140) );
  NANDN U15586 ( .A(n14875), .B(n14874), .Z(n14879) );
  NANDN U15587 ( .A(n14877), .B(n14876), .Z(n14878) );
  AND U15588 ( .A(n14879), .B(n14878), .Z(n15085) );
  NAND U15589 ( .A(n38385), .B(n14880), .Z(n14882) );
  XOR U15590 ( .A(b[27]), .B(a[89]), .Z(n15029) );
  NAND U15591 ( .A(n38343), .B(n15029), .Z(n14881) );
  AND U15592 ( .A(n14882), .B(n14881), .Z(n15092) );
  NAND U15593 ( .A(n183), .B(n14883), .Z(n14885) );
  XOR U15594 ( .A(b[5]), .B(a[111]), .Z(n15032) );
  NAND U15595 ( .A(n36296), .B(n15032), .Z(n14884) );
  AND U15596 ( .A(n14885), .B(n14884), .Z(n15090) );
  NAND U15597 ( .A(n190), .B(n14886), .Z(n14888) );
  XOR U15598 ( .A(b[19]), .B(a[97]), .Z(n15035) );
  NAND U15599 ( .A(n37821), .B(n15035), .Z(n14887) );
  NAND U15600 ( .A(n14888), .B(n14887), .Z(n15089) );
  XNOR U15601 ( .A(n15090), .B(n15089), .Z(n15091) );
  XNOR U15602 ( .A(n15092), .B(n15091), .Z(n15083) );
  NAND U15603 ( .A(n38470), .B(n14889), .Z(n14891) );
  XOR U15604 ( .A(b[31]), .B(a[85]), .Z(n15038) );
  NAND U15605 ( .A(n38453), .B(n15038), .Z(n14890) );
  AND U15606 ( .A(n14891), .B(n14890), .Z(n15050) );
  NAND U15607 ( .A(n181), .B(n14892), .Z(n14894) );
  XOR U15608 ( .A(b[3]), .B(a[113]), .Z(n15041) );
  NAND U15609 ( .A(n182), .B(n15041), .Z(n14893) );
  AND U15610 ( .A(n14894), .B(n14893), .Z(n15048) );
  NAND U15611 ( .A(n189), .B(n14895), .Z(n14897) );
  XOR U15612 ( .A(b[17]), .B(a[99]), .Z(n15044) );
  NAND U15613 ( .A(n37652), .B(n15044), .Z(n14896) );
  NAND U15614 ( .A(n14897), .B(n14896), .Z(n15047) );
  XNOR U15615 ( .A(n15048), .B(n15047), .Z(n15049) );
  XOR U15616 ( .A(n15050), .B(n15049), .Z(n15084) );
  XOR U15617 ( .A(n15083), .B(n15084), .Z(n15086) );
  XOR U15618 ( .A(n15085), .B(n15086), .Z(n15018) );
  NANDN U15619 ( .A(n14899), .B(n14898), .Z(n14903) );
  NANDN U15620 ( .A(n14901), .B(n14900), .Z(n14902) );
  AND U15621 ( .A(n14903), .B(n14902), .Z(n15071) );
  NANDN U15622 ( .A(n14905), .B(n14904), .Z(n14909) );
  NANDN U15623 ( .A(n14907), .B(n14906), .Z(n14908) );
  NAND U15624 ( .A(n14909), .B(n14908), .Z(n15072) );
  XNOR U15625 ( .A(n15071), .B(n15072), .Z(n15073) );
  NANDN U15626 ( .A(n14911), .B(n14910), .Z(n14915) );
  NANDN U15627 ( .A(n14913), .B(n14912), .Z(n14914) );
  NAND U15628 ( .A(n14915), .B(n14914), .Z(n15074) );
  XNOR U15629 ( .A(n15073), .B(n15074), .Z(n15017) );
  XNOR U15630 ( .A(n15018), .B(n15017), .Z(n15020) );
  NANDN U15631 ( .A(n14917), .B(n14916), .Z(n14921) );
  NANDN U15632 ( .A(n14919), .B(n14918), .Z(n14920) );
  AND U15633 ( .A(n14921), .B(n14920), .Z(n15019) );
  XOR U15634 ( .A(n15020), .B(n15019), .Z(n15134) );
  NANDN U15635 ( .A(n14923), .B(n14922), .Z(n14927) );
  NANDN U15636 ( .A(n14925), .B(n14924), .Z(n14926) );
  AND U15637 ( .A(n14927), .B(n14926), .Z(n15131) );
  NANDN U15638 ( .A(n14929), .B(n14928), .Z(n14933) );
  NANDN U15639 ( .A(n14931), .B(n14930), .Z(n14932) );
  AND U15640 ( .A(n14933), .B(n14932), .Z(n15014) );
  NANDN U15641 ( .A(n14935), .B(n14934), .Z(n14939) );
  OR U15642 ( .A(n14937), .B(n14936), .Z(n14938) );
  AND U15643 ( .A(n14939), .B(n14938), .Z(n15012) );
  NANDN U15644 ( .A(n14941), .B(n14940), .Z(n14945) );
  NANDN U15645 ( .A(n14943), .B(n14942), .Z(n14944) );
  AND U15646 ( .A(n14945), .B(n14944), .Z(n15078) );
  NANDN U15647 ( .A(n14947), .B(n14946), .Z(n14951) );
  NANDN U15648 ( .A(n14949), .B(n14948), .Z(n14950) );
  NAND U15649 ( .A(n14951), .B(n14950), .Z(n15077) );
  XNOR U15650 ( .A(n15078), .B(n15077), .Z(n15079) );
  NAND U15651 ( .A(b[0]), .B(a[115]), .Z(n14952) );
  XNOR U15652 ( .A(b[1]), .B(n14952), .Z(n14954) );
  NANDN U15653 ( .A(b[0]), .B(a[114]), .Z(n14953) );
  NAND U15654 ( .A(n14954), .B(n14953), .Z(n15026) );
  NAND U15655 ( .A(n194), .B(n14955), .Z(n14957) );
  XOR U15656 ( .A(b[29]), .B(a[87]), .Z(n15104) );
  NAND U15657 ( .A(n38456), .B(n15104), .Z(n14956) );
  AND U15658 ( .A(n14957), .B(n14956), .Z(n15024) );
  AND U15659 ( .A(b[31]), .B(a[83]), .Z(n15023) );
  XNOR U15660 ( .A(n15024), .B(n15023), .Z(n15025) );
  XNOR U15661 ( .A(n15026), .B(n15025), .Z(n15065) );
  NAND U15662 ( .A(n38185), .B(n14958), .Z(n14960) );
  XOR U15663 ( .A(b[23]), .B(a[93]), .Z(n15107) );
  NAND U15664 ( .A(n38132), .B(n15107), .Z(n14959) );
  AND U15665 ( .A(n14960), .B(n14959), .Z(n15098) );
  NAND U15666 ( .A(n184), .B(n14961), .Z(n14963) );
  XOR U15667 ( .A(b[7]), .B(a[109]), .Z(n15110) );
  NAND U15668 ( .A(n36592), .B(n15110), .Z(n14962) );
  AND U15669 ( .A(n14963), .B(n14962), .Z(n15096) );
  NAND U15670 ( .A(n38289), .B(n14964), .Z(n14966) );
  XOR U15671 ( .A(b[25]), .B(a[91]), .Z(n15113) );
  NAND U15672 ( .A(n38247), .B(n15113), .Z(n14965) );
  NAND U15673 ( .A(n14966), .B(n14965), .Z(n15095) );
  XNOR U15674 ( .A(n15096), .B(n15095), .Z(n15097) );
  XOR U15675 ( .A(n15098), .B(n15097), .Z(n15066) );
  XNOR U15676 ( .A(n15065), .B(n15066), .Z(n15067) );
  NAND U15677 ( .A(n187), .B(n14967), .Z(n14969) );
  XOR U15678 ( .A(b[13]), .B(a[103]), .Z(n15116) );
  NAND U15679 ( .A(n37295), .B(n15116), .Z(n14968) );
  AND U15680 ( .A(n14969), .B(n14968), .Z(n15060) );
  NAND U15681 ( .A(n186), .B(n14970), .Z(n14972) );
  XOR U15682 ( .A(b[11]), .B(a[105]), .Z(n15119) );
  NAND U15683 ( .A(n37097), .B(n15119), .Z(n14971) );
  NAND U15684 ( .A(n14972), .B(n14971), .Z(n15059) );
  XNOR U15685 ( .A(n15060), .B(n15059), .Z(n15061) );
  NAND U15686 ( .A(n188), .B(n14973), .Z(n14975) );
  XOR U15687 ( .A(b[15]), .B(a[101]), .Z(n15122) );
  NAND U15688 ( .A(n37382), .B(n15122), .Z(n14974) );
  AND U15689 ( .A(n14975), .B(n14974), .Z(n15056) );
  NAND U15690 ( .A(n38064), .B(n14976), .Z(n14978) );
  XOR U15691 ( .A(b[21]), .B(a[95]), .Z(n15125) );
  NAND U15692 ( .A(n37993), .B(n15125), .Z(n14977) );
  AND U15693 ( .A(n14978), .B(n14977), .Z(n15054) );
  NAND U15694 ( .A(n185), .B(n14979), .Z(n14981) );
  XOR U15695 ( .A(b[9]), .B(a[107]), .Z(n15128) );
  NAND U15696 ( .A(n36805), .B(n15128), .Z(n14980) );
  NAND U15697 ( .A(n14981), .B(n14980), .Z(n15053) );
  XNOR U15698 ( .A(n15054), .B(n15053), .Z(n15055) );
  XOR U15699 ( .A(n15056), .B(n15055), .Z(n15062) );
  XOR U15700 ( .A(n15061), .B(n15062), .Z(n15068) );
  XOR U15701 ( .A(n15067), .B(n15068), .Z(n15080) );
  XNOR U15702 ( .A(n15079), .B(n15080), .Z(n15011) );
  XNOR U15703 ( .A(n15012), .B(n15011), .Z(n15013) );
  XOR U15704 ( .A(n15014), .B(n15013), .Z(n15132) );
  XNOR U15705 ( .A(n15131), .B(n15132), .Z(n15133) );
  XNOR U15706 ( .A(n15134), .B(n15133), .Z(n15139) );
  XOR U15707 ( .A(n15140), .B(n15139), .Z(n15006) );
  NANDN U15708 ( .A(n14983), .B(n14982), .Z(n14987) );
  NANDN U15709 ( .A(n14985), .B(n14984), .Z(n14986) );
  AND U15710 ( .A(n14987), .B(n14986), .Z(n15005) );
  XNOR U15711 ( .A(n15006), .B(n15005), .Z(n15007) );
  NANDN U15712 ( .A(n14989), .B(n14988), .Z(n14993) );
  NAND U15713 ( .A(n14991), .B(n14990), .Z(n14992) );
  NAND U15714 ( .A(n14993), .B(n14992), .Z(n15008) );
  XNOR U15715 ( .A(n15007), .B(n15008), .Z(n14999) );
  XNOR U15716 ( .A(n15000), .B(n14999), .Z(n15001) );
  XNOR U15717 ( .A(n15002), .B(n15001), .Z(n15143) );
  XNOR U15718 ( .A(sreg[339]), .B(n15143), .Z(n15145) );
  NANDN U15719 ( .A(sreg[338]), .B(n14994), .Z(n14998) );
  NAND U15720 ( .A(n14996), .B(n14995), .Z(n14997) );
  NAND U15721 ( .A(n14998), .B(n14997), .Z(n15144) );
  XNOR U15722 ( .A(n15145), .B(n15144), .Z(c[339]) );
  NANDN U15723 ( .A(n15000), .B(n14999), .Z(n15004) );
  NANDN U15724 ( .A(n15002), .B(n15001), .Z(n15003) );
  AND U15725 ( .A(n15004), .B(n15003), .Z(n15151) );
  NANDN U15726 ( .A(n15006), .B(n15005), .Z(n15010) );
  NANDN U15727 ( .A(n15008), .B(n15007), .Z(n15009) );
  AND U15728 ( .A(n15010), .B(n15009), .Z(n15149) );
  NANDN U15729 ( .A(n15012), .B(n15011), .Z(n15016) );
  NANDN U15730 ( .A(n15014), .B(n15013), .Z(n15015) );
  AND U15731 ( .A(n15016), .B(n15015), .Z(n15287) );
  NANDN U15732 ( .A(n15018), .B(n15017), .Z(n15022) );
  NAND U15733 ( .A(n15020), .B(n15019), .Z(n15021) );
  AND U15734 ( .A(n15022), .B(n15021), .Z(n15286) );
  XNOR U15735 ( .A(n15287), .B(n15286), .Z(n15289) );
  NANDN U15736 ( .A(n15024), .B(n15023), .Z(n15028) );
  NANDN U15737 ( .A(n15026), .B(n15025), .Z(n15027) );
  AND U15738 ( .A(n15028), .B(n15027), .Z(n15234) );
  NAND U15739 ( .A(n38385), .B(n15029), .Z(n15031) );
  XOR U15740 ( .A(b[27]), .B(a[90]), .Z(n15178) );
  NAND U15741 ( .A(n38343), .B(n15178), .Z(n15030) );
  AND U15742 ( .A(n15031), .B(n15030), .Z(n15241) );
  NAND U15743 ( .A(n183), .B(n15032), .Z(n15034) );
  XOR U15744 ( .A(b[5]), .B(a[112]), .Z(n15181) );
  NAND U15745 ( .A(n36296), .B(n15181), .Z(n15033) );
  AND U15746 ( .A(n15034), .B(n15033), .Z(n15239) );
  NAND U15747 ( .A(n190), .B(n15035), .Z(n15037) );
  XOR U15748 ( .A(b[19]), .B(a[98]), .Z(n15184) );
  NAND U15749 ( .A(n37821), .B(n15184), .Z(n15036) );
  NAND U15750 ( .A(n15037), .B(n15036), .Z(n15238) );
  XNOR U15751 ( .A(n15239), .B(n15238), .Z(n15240) );
  XNOR U15752 ( .A(n15241), .B(n15240), .Z(n15232) );
  NAND U15753 ( .A(n38470), .B(n15038), .Z(n15040) );
  XOR U15754 ( .A(b[31]), .B(a[86]), .Z(n15187) );
  NAND U15755 ( .A(n38453), .B(n15187), .Z(n15039) );
  AND U15756 ( .A(n15040), .B(n15039), .Z(n15199) );
  NAND U15757 ( .A(n181), .B(n15041), .Z(n15043) );
  XOR U15758 ( .A(b[3]), .B(a[114]), .Z(n15190) );
  NAND U15759 ( .A(n182), .B(n15190), .Z(n15042) );
  AND U15760 ( .A(n15043), .B(n15042), .Z(n15197) );
  NAND U15761 ( .A(n189), .B(n15044), .Z(n15046) );
  XOR U15762 ( .A(b[17]), .B(a[100]), .Z(n15193) );
  NAND U15763 ( .A(n37652), .B(n15193), .Z(n15045) );
  NAND U15764 ( .A(n15046), .B(n15045), .Z(n15196) );
  XNOR U15765 ( .A(n15197), .B(n15196), .Z(n15198) );
  XOR U15766 ( .A(n15199), .B(n15198), .Z(n15233) );
  XOR U15767 ( .A(n15232), .B(n15233), .Z(n15235) );
  XOR U15768 ( .A(n15234), .B(n15235), .Z(n15167) );
  NANDN U15769 ( .A(n15048), .B(n15047), .Z(n15052) );
  NANDN U15770 ( .A(n15050), .B(n15049), .Z(n15051) );
  AND U15771 ( .A(n15052), .B(n15051), .Z(n15220) );
  NANDN U15772 ( .A(n15054), .B(n15053), .Z(n15058) );
  NANDN U15773 ( .A(n15056), .B(n15055), .Z(n15057) );
  NAND U15774 ( .A(n15058), .B(n15057), .Z(n15221) );
  XNOR U15775 ( .A(n15220), .B(n15221), .Z(n15222) );
  NANDN U15776 ( .A(n15060), .B(n15059), .Z(n15064) );
  NANDN U15777 ( .A(n15062), .B(n15061), .Z(n15063) );
  NAND U15778 ( .A(n15064), .B(n15063), .Z(n15223) );
  XNOR U15779 ( .A(n15222), .B(n15223), .Z(n15166) );
  XNOR U15780 ( .A(n15167), .B(n15166), .Z(n15169) );
  NANDN U15781 ( .A(n15066), .B(n15065), .Z(n15070) );
  NANDN U15782 ( .A(n15068), .B(n15067), .Z(n15069) );
  AND U15783 ( .A(n15070), .B(n15069), .Z(n15168) );
  XOR U15784 ( .A(n15169), .B(n15168), .Z(n15283) );
  NANDN U15785 ( .A(n15072), .B(n15071), .Z(n15076) );
  NANDN U15786 ( .A(n15074), .B(n15073), .Z(n15075) );
  AND U15787 ( .A(n15076), .B(n15075), .Z(n15280) );
  NANDN U15788 ( .A(n15078), .B(n15077), .Z(n15082) );
  NANDN U15789 ( .A(n15080), .B(n15079), .Z(n15081) );
  AND U15790 ( .A(n15082), .B(n15081), .Z(n15163) );
  NANDN U15791 ( .A(n15084), .B(n15083), .Z(n15088) );
  OR U15792 ( .A(n15086), .B(n15085), .Z(n15087) );
  AND U15793 ( .A(n15088), .B(n15087), .Z(n15161) );
  NANDN U15794 ( .A(n15090), .B(n15089), .Z(n15094) );
  NANDN U15795 ( .A(n15092), .B(n15091), .Z(n15093) );
  AND U15796 ( .A(n15094), .B(n15093), .Z(n15227) );
  NANDN U15797 ( .A(n15096), .B(n15095), .Z(n15100) );
  NANDN U15798 ( .A(n15098), .B(n15097), .Z(n15099) );
  NAND U15799 ( .A(n15100), .B(n15099), .Z(n15226) );
  XNOR U15800 ( .A(n15227), .B(n15226), .Z(n15228) );
  NAND U15801 ( .A(b[0]), .B(a[116]), .Z(n15101) );
  XNOR U15802 ( .A(b[1]), .B(n15101), .Z(n15103) );
  NANDN U15803 ( .A(b[0]), .B(a[115]), .Z(n15102) );
  NAND U15804 ( .A(n15103), .B(n15102), .Z(n15175) );
  NAND U15805 ( .A(n194), .B(n15104), .Z(n15106) );
  XOR U15806 ( .A(b[29]), .B(a[88]), .Z(n15253) );
  NAND U15807 ( .A(n38456), .B(n15253), .Z(n15105) );
  AND U15808 ( .A(n15106), .B(n15105), .Z(n15173) );
  AND U15809 ( .A(b[31]), .B(a[84]), .Z(n15172) );
  XNOR U15810 ( .A(n15173), .B(n15172), .Z(n15174) );
  XNOR U15811 ( .A(n15175), .B(n15174), .Z(n15214) );
  NAND U15812 ( .A(n38185), .B(n15107), .Z(n15109) );
  XOR U15813 ( .A(b[23]), .B(a[94]), .Z(n15256) );
  NAND U15814 ( .A(n38132), .B(n15256), .Z(n15108) );
  AND U15815 ( .A(n15109), .B(n15108), .Z(n15247) );
  NAND U15816 ( .A(n184), .B(n15110), .Z(n15112) );
  XOR U15817 ( .A(b[7]), .B(a[110]), .Z(n15259) );
  NAND U15818 ( .A(n36592), .B(n15259), .Z(n15111) );
  AND U15819 ( .A(n15112), .B(n15111), .Z(n15245) );
  NAND U15820 ( .A(n38289), .B(n15113), .Z(n15115) );
  XOR U15821 ( .A(b[25]), .B(a[92]), .Z(n15262) );
  NAND U15822 ( .A(n38247), .B(n15262), .Z(n15114) );
  NAND U15823 ( .A(n15115), .B(n15114), .Z(n15244) );
  XNOR U15824 ( .A(n15245), .B(n15244), .Z(n15246) );
  XOR U15825 ( .A(n15247), .B(n15246), .Z(n15215) );
  XNOR U15826 ( .A(n15214), .B(n15215), .Z(n15216) );
  NAND U15827 ( .A(n187), .B(n15116), .Z(n15118) );
  XOR U15828 ( .A(b[13]), .B(a[104]), .Z(n15265) );
  NAND U15829 ( .A(n37295), .B(n15265), .Z(n15117) );
  AND U15830 ( .A(n15118), .B(n15117), .Z(n15209) );
  NAND U15831 ( .A(n186), .B(n15119), .Z(n15121) );
  XOR U15832 ( .A(b[11]), .B(a[106]), .Z(n15268) );
  NAND U15833 ( .A(n37097), .B(n15268), .Z(n15120) );
  NAND U15834 ( .A(n15121), .B(n15120), .Z(n15208) );
  XNOR U15835 ( .A(n15209), .B(n15208), .Z(n15210) );
  NAND U15836 ( .A(n188), .B(n15122), .Z(n15124) );
  XOR U15837 ( .A(b[15]), .B(a[102]), .Z(n15271) );
  NAND U15838 ( .A(n37382), .B(n15271), .Z(n15123) );
  AND U15839 ( .A(n15124), .B(n15123), .Z(n15205) );
  NAND U15840 ( .A(n38064), .B(n15125), .Z(n15127) );
  XOR U15841 ( .A(b[21]), .B(a[96]), .Z(n15274) );
  NAND U15842 ( .A(n37993), .B(n15274), .Z(n15126) );
  AND U15843 ( .A(n15127), .B(n15126), .Z(n15203) );
  NAND U15844 ( .A(n185), .B(n15128), .Z(n15130) );
  XOR U15845 ( .A(b[9]), .B(a[108]), .Z(n15277) );
  NAND U15846 ( .A(n36805), .B(n15277), .Z(n15129) );
  NAND U15847 ( .A(n15130), .B(n15129), .Z(n15202) );
  XNOR U15848 ( .A(n15203), .B(n15202), .Z(n15204) );
  XOR U15849 ( .A(n15205), .B(n15204), .Z(n15211) );
  XOR U15850 ( .A(n15210), .B(n15211), .Z(n15217) );
  XOR U15851 ( .A(n15216), .B(n15217), .Z(n15229) );
  XNOR U15852 ( .A(n15228), .B(n15229), .Z(n15160) );
  XNOR U15853 ( .A(n15161), .B(n15160), .Z(n15162) );
  XOR U15854 ( .A(n15163), .B(n15162), .Z(n15281) );
  XNOR U15855 ( .A(n15280), .B(n15281), .Z(n15282) );
  XNOR U15856 ( .A(n15283), .B(n15282), .Z(n15288) );
  XOR U15857 ( .A(n15289), .B(n15288), .Z(n15155) );
  NANDN U15858 ( .A(n15132), .B(n15131), .Z(n15136) );
  NANDN U15859 ( .A(n15134), .B(n15133), .Z(n15135) );
  AND U15860 ( .A(n15136), .B(n15135), .Z(n15154) );
  XNOR U15861 ( .A(n15155), .B(n15154), .Z(n15156) );
  NANDN U15862 ( .A(n15138), .B(n15137), .Z(n15142) );
  NAND U15863 ( .A(n15140), .B(n15139), .Z(n15141) );
  NAND U15864 ( .A(n15142), .B(n15141), .Z(n15157) );
  XNOR U15865 ( .A(n15156), .B(n15157), .Z(n15148) );
  XNOR U15866 ( .A(n15149), .B(n15148), .Z(n15150) );
  XNOR U15867 ( .A(n15151), .B(n15150), .Z(n15292) );
  XNOR U15868 ( .A(sreg[340]), .B(n15292), .Z(n15294) );
  NANDN U15869 ( .A(sreg[339]), .B(n15143), .Z(n15147) );
  NAND U15870 ( .A(n15145), .B(n15144), .Z(n15146) );
  NAND U15871 ( .A(n15147), .B(n15146), .Z(n15293) );
  XNOR U15872 ( .A(n15294), .B(n15293), .Z(c[340]) );
  NANDN U15873 ( .A(n15149), .B(n15148), .Z(n15153) );
  NANDN U15874 ( .A(n15151), .B(n15150), .Z(n15152) );
  AND U15875 ( .A(n15153), .B(n15152), .Z(n15300) );
  NANDN U15876 ( .A(n15155), .B(n15154), .Z(n15159) );
  NANDN U15877 ( .A(n15157), .B(n15156), .Z(n15158) );
  AND U15878 ( .A(n15159), .B(n15158), .Z(n15298) );
  NANDN U15879 ( .A(n15161), .B(n15160), .Z(n15165) );
  NANDN U15880 ( .A(n15163), .B(n15162), .Z(n15164) );
  AND U15881 ( .A(n15165), .B(n15164), .Z(n15310) );
  NANDN U15882 ( .A(n15167), .B(n15166), .Z(n15171) );
  NAND U15883 ( .A(n15169), .B(n15168), .Z(n15170) );
  AND U15884 ( .A(n15171), .B(n15170), .Z(n15309) );
  XNOR U15885 ( .A(n15310), .B(n15309), .Z(n15312) );
  NANDN U15886 ( .A(n15173), .B(n15172), .Z(n15177) );
  NANDN U15887 ( .A(n15175), .B(n15174), .Z(n15176) );
  AND U15888 ( .A(n15177), .B(n15176), .Z(n15389) );
  NAND U15889 ( .A(n38385), .B(n15178), .Z(n15180) );
  XOR U15890 ( .A(b[27]), .B(a[91]), .Z(n15333) );
  NAND U15891 ( .A(n38343), .B(n15333), .Z(n15179) );
  AND U15892 ( .A(n15180), .B(n15179), .Z(n15396) );
  NAND U15893 ( .A(n183), .B(n15181), .Z(n15183) );
  XOR U15894 ( .A(b[5]), .B(a[113]), .Z(n15336) );
  NAND U15895 ( .A(n36296), .B(n15336), .Z(n15182) );
  AND U15896 ( .A(n15183), .B(n15182), .Z(n15394) );
  NAND U15897 ( .A(n190), .B(n15184), .Z(n15186) );
  XOR U15898 ( .A(b[19]), .B(a[99]), .Z(n15339) );
  NAND U15899 ( .A(n37821), .B(n15339), .Z(n15185) );
  NAND U15900 ( .A(n15186), .B(n15185), .Z(n15393) );
  XNOR U15901 ( .A(n15394), .B(n15393), .Z(n15395) );
  XNOR U15902 ( .A(n15396), .B(n15395), .Z(n15387) );
  NAND U15903 ( .A(n38470), .B(n15187), .Z(n15189) );
  XOR U15904 ( .A(b[31]), .B(a[87]), .Z(n15342) );
  NAND U15905 ( .A(n38453), .B(n15342), .Z(n15188) );
  AND U15906 ( .A(n15189), .B(n15188), .Z(n15354) );
  NAND U15907 ( .A(n181), .B(n15190), .Z(n15192) );
  XOR U15908 ( .A(b[3]), .B(a[115]), .Z(n15345) );
  NAND U15909 ( .A(n182), .B(n15345), .Z(n15191) );
  AND U15910 ( .A(n15192), .B(n15191), .Z(n15352) );
  NAND U15911 ( .A(n189), .B(n15193), .Z(n15195) );
  XOR U15912 ( .A(b[17]), .B(a[101]), .Z(n15348) );
  NAND U15913 ( .A(n37652), .B(n15348), .Z(n15194) );
  NAND U15914 ( .A(n15195), .B(n15194), .Z(n15351) );
  XNOR U15915 ( .A(n15352), .B(n15351), .Z(n15353) );
  XOR U15916 ( .A(n15354), .B(n15353), .Z(n15388) );
  XOR U15917 ( .A(n15387), .B(n15388), .Z(n15390) );
  XOR U15918 ( .A(n15389), .B(n15390), .Z(n15322) );
  NANDN U15919 ( .A(n15197), .B(n15196), .Z(n15201) );
  NANDN U15920 ( .A(n15199), .B(n15198), .Z(n15200) );
  AND U15921 ( .A(n15201), .B(n15200), .Z(n15375) );
  NANDN U15922 ( .A(n15203), .B(n15202), .Z(n15207) );
  NANDN U15923 ( .A(n15205), .B(n15204), .Z(n15206) );
  NAND U15924 ( .A(n15207), .B(n15206), .Z(n15376) );
  XNOR U15925 ( .A(n15375), .B(n15376), .Z(n15377) );
  NANDN U15926 ( .A(n15209), .B(n15208), .Z(n15213) );
  NANDN U15927 ( .A(n15211), .B(n15210), .Z(n15212) );
  NAND U15928 ( .A(n15213), .B(n15212), .Z(n15378) );
  XNOR U15929 ( .A(n15377), .B(n15378), .Z(n15321) );
  XNOR U15930 ( .A(n15322), .B(n15321), .Z(n15324) );
  NANDN U15931 ( .A(n15215), .B(n15214), .Z(n15219) );
  NANDN U15932 ( .A(n15217), .B(n15216), .Z(n15218) );
  AND U15933 ( .A(n15219), .B(n15218), .Z(n15323) );
  XOR U15934 ( .A(n15324), .B(n15323), .Z(n15438) );
  NANDN U15935 ( .A(n15221), .B(n15220), .Z(n15225) );
  NANDN U15936 ( .A(n15223), .B(n15222), .Z(n15224) );
  AND U15937 ( .A(n15225), .B(n15224), .Z(n15435) );
  NANDN U15938 ( .A(n15227), .B(n15226), .Z(n15231) );
  NANDN U15939 ( .A(n15229), .B(n15228), .Z(n15230) );
  AND U15940 ( .A(n15231), .B(n15230), .Z(n15318) );
  NANDN U15941 ( .A(n15233), .B(n15232), .Z(n15237) );
  OR U15942 ( .A(n15235), .B(n15234), .Z(n15236) );
  AND U15943 ( .A(n15237), .B(n15236), .Z(n15316) );
  NANDN U15944 ( .A(n15239), .B(n15238), .Z(n15243) );
  NANDN U15945 ( .A(n15241), .B(n15240), .Z(n15242) );
  AND U15946 ( .A(n15243), .B(n15242), .Z(n15382) );
  NANDN U15947 ( .A(n15245), .B(n15244), .Z(n15249) );
  NANDN U15948 ( .A(n15247), .B(n15246), .Z(n15248) );
  NAND U15949 ( .A(n15249), .B(n15248), .Z(n15381) );
  XNOR U15950 ( .A(n15382), .B(n15381), .Z(n15383) );
  NAND U15951 ( .A(b[0]), .B(a[117]), .Z(n15250) );
  XNOR U15952 ( .A(b[1]), .B(n15250), .Z(n15252) );
  NANDN U15953 ( .A(b[0]), .B(a[116]), .Z(n15251) );
  NAND U15954 ( .A(n15252), .B(n15251), .Z(n15330) );
  NAND U15955 ( .A(n194), .B(n15253), .Z(n15255) );
  XOR U15956 ( .A(b[29]), .B(a[89]), .Z(n15408) );
  NAND U15957 ( .A(n38456), .B(n15408), .Z(n15254) );
  AND U15958 ( .A(n15255), .B(n15254), .Z(n15328) );
  AND U15959 ( .A(b[31]), .B(a[85]), .Z(n15327) );
  XNOR U15960 ( .A(n15328), .B(n15327), .Z(n15329) );
  XNOR U15961 ( .A(n15330), .B(n15329), .Z(n15369) );
  NAND U15962 ( .A(n38185), .B(n15256), .Z(n15258) );
  XOR U15963 ( .A(b[23]), .B(a[95]), .Z(n15411) );
  NAND U15964 ( .A(n38132), .B(n15411), .Z(n15257) );
  AND U15965 ( .A(n15258), .B(n15257), .Z(n15402) );
  NAND U15966 ( .A(n184), .B(n15259), .Z(n15261) );
  XOR U15967 ( .A(b[7]), .B(a[111]), .Z(n15414) );
  NAND U15968 ( .A(n36592), .B(n15414), .Z(n15260) );
  AND U15969 ( .A(n15261), .B(n15260), .Z(n15400) );
  NAND U15970 ( .A(n38289), .B(n15262), .Z(n15264) );
  XOR U15971 ( .A(b[25]), .B(a[93]), .Z(n15417) );
  NAND U15972 ( .A(n38247), .B(n15417), .Z(n15263) );
  NAND U15973 ( .A(n15264), .B(n15263), .Z(n15399) );
  XNOR U15974 ( .A(n15400), .B(n15399), .Z(n15401) );
  XOR U15975 ( .A(n15402), .B(n15401), .Z(n15370) );
  XNOR U15976 ( .A(n15369), .B(n15370), .Z(n15371) );
  NAND U15977 ( .A(n187), .B(n15265), .Z(n15267) );
  XOR U15978 ( .A(b[13]), .B(a[105]), .Z(n15420) );
  NAND U15979 ( .A(n37295), .B(n15420), .Z(n15266) );
  AND U15980 ( .A(n15267), .B(n15266), .Z(n15364) );
  NAND U15981 ( .A(n186), .B(n15268), .Z(n15270) );
  XOR U15982 ( .A(b[11]), .B(a[107]), .Z(n15423) );
  NAND U15983 ( .A(n37097), .B(n15423), .Z(n15269) );
  NAND U15984 ( .A(n15270), .B(n15269), .Z(n15363) );
  XNOR U15985 ( .A(n15364), .B(n15363), .Z(n15365) );
  NAND U15986 ( .A(n188), .B(n15271), .Z(n15273) );
  XOR U15987 ( .A(b[15]), .B(a[103]), .Z(n15426) );
  NAND U15988 ( .A(n37382), .B(n15426), .Z(n15272) );
  AND U15989 ( .A(n15273), .B(n15272), .Z(n15360) );
  NAND U15990 ( .A(n38064), .B(n15274), .Z(n15276) );
  XOR U15991 ( .A(b[21]), .B(a[97]), .Z(n15429) );
  NAND U15992 ( .A(n37993), .B(n15429), .Z(n15275) );
  AND U15993 ( .A(n15276), .B(n15275), .Z(n15358) );
  NAND U15994 ( .A(n185), .B(n15277), .Z(n15279) );
  XOR U15995 ( .A(b[9]), .B(a[109]), .Z(n15432) );
  NAND U15996 ( .A(n36805), .B(n15432), .Z(n15278) );
  NAND U15997 ( .A(n15279), .B(n15278), .Z(n15357) );
  XNOR U15998 ( .A(n15358), .B(n15357), .Z(n15359) );
  XOR U15999 ( .A(n15360), .B(n15359), .Z(n15366) );
  XOR U16000 ( .A(n15365), .B(n15366), .Z(n15372) );
  XOR U16001 ( .A(n15371), .B(n15372), .Z(n15384) );
  XNOR U16002 ( .A(n15383), .B(n15384), .Z(n15315) );
  XNOR U16003 ( .A(n15316), .B(n15315), .Z(n15317) );
  XOR U16004 ( .A(n15318), .B(n15317), .Z(n15436) );
  XNOR U16005 ( .A(n15435), .B(n15436), .Z(n15437) );
  XNOR U16006 ( .A(n15438), .B(n15437), .Z(n15311) );
  XOR U16007 ( .A(n15312), .B(n15311), .Z(n15304) );
  NANDN U16008 ( .A(n15281), .B(n15280), .Z(n15285) );
  NANDN U16009 ( .A(n15283), .B(n15282), .Z(n15284) );
  AND U16010 ( .A(n15285), .B(n15284), .Z(n15303) );
  XNOR U16011 ( .A(n15304), .B(n15303), .Z(n15305) );
  NANDN U16012 ( .A(n15287), .B(n15286), .Z(n15291) );
  NAND U16013 ( .A(n15289), .B(n15288), .Z(n15290) );
  NAND U16014 ( .A(n15291), .B(n15290), .Z(n15306) );
  XNOR U16015 ( .A(n15305), .B(n15306), .Z(n15297) );
  XNOR U16016 ( .A(n15298), .B(n15297), .Z(n15299) );
  XNOR U16017 ( .A(n15300), .B(n15299), .Z(n15441) );
  XNOR U16018 ( .A(sreg[341]), .B(n15441), .Z(n15443) );
  NANDN U16019 ( .A(sreg[340]), .B(n15292), .Z(n15296) );
  NAND U16020 ( .A(n15294), .B(n15293), .Z(n15295) );
  NAND U16021 ( .A(n15296), .B(n15295), .Z(n15442) );
  XNOR U16022 ( .A(n15443), .B(n15442), .Z(c[341]) );
  NANDN U16023 ( .A(n15298), .B(n15297), .Z(n15302) );
  NANDN U16024 ( .A(n15300), .B(n15299), .Z(n15301) );
  AND U16025 ( .A(n15302), .B(n15301), .Z(n15449) );
  NANDN U16026 ( .A(n15304), .B(n15303), .Z(n15308) );
  NANDN U16027 ( .A(n15306), .B(n15305), .Z(n15307) );
  AND U16028 ( .A(n15308), .B(n15307), .Z(n15447) );
  NANDN U16029 ( .A(n15310), .B(n15309), .Z(n15314) );
  NAND U16030 ( .A(n15312), .B(n15311), .Z(n15313) );
  AND U16031 ( .A(n15314), .B(n15313), .Z(n15454) );
  NANDN U16032 ( .A(n15316), .B(n15315), .Z(n15320) );
  NANDN U16033 ( .A(n15318), .B(n15317), .Z(n15319) );
  AND U16034 ( .A(n15320), .B(n15319), .Z(n15459) );
  NANDN U16035 ( .A(n15322), .B(n15321), .Z(n15326) );
  NAND U16036 ( .A(n15324), .B(n15323), .Z(n15325) );
  AND U16037 ( .A(n15326), .B(n15325), .Z(n15458) );
  XNOR U16038 ( .A(n15459), .B(n15458), .Z(n15461) );
  NANDN U16039 ( .A(n15328), .B(n15327), .Z(n15332) );
  NANDN U16040 ( .A(n15330), .B(n15329), .Z(n15331) );
  AND U16041 ( .A(n15332), .B(n15331), .Z(n15538) );
  NAND U16042 ( .A(n38385), .B(n15333), .Z(n15335) );
  XOR U16043 ( .A(b[27]), .B(a[92]), .Z(n15482) );
  NAND U16044 ( .A(n38343), .B(n15482), .Z(n15334) );
  AND U16045 ( .A(n15335), .B(n15334), .Z(n15545) );
  NAND U16046 ( .A(n183), .B(n15336), .Z(n15338) );
  XOR U16047 ( .A(b[5]), .B(a[114]), .Z(n15485) );
  NAND U16048 ( .A(n36296), .B(n15485), .Z(n15337) );
  AND U16049 ( .A(n15338), .B(n15337), .Z(n15543) );
  NAND U16050 ( .A(n190), .B(n15339), .Z(n15341) );
  XOR U16051 ( .A(b[19]), .B(a[100]), .Z(n15488) );
  NAND U16052 ( .A(n37821), .B(n15488), .Z(n15340) );
  NAND U16053 ( .A(n15341), .B(n15340), .Z(n15542) );
  XNOR U16054 ( .A(n15543), .B(n15542), .Z(n15544) );
  XNOR U16055 ( .A(n15545), .B(n15544), .Z(n15536) );
  NAND U16056 ( .A(n38470), .B(n15342), .Z(n15344) );
  XOR U16057 ( .A(b[31]), .B(a[88]), .Z(n15491) );
  NAND U16058 ( .A(n38453), .B(n15491), .Z(n15343) );
  AND U16059 ( .A(n15344), .B(n15343), .Z(n15503) );
  NAND U16060 ( .A(n181), .B(n15345), .Z(n15347) );
  XOR U16061 ( .A(b[3]), .B(a[116]), .Z(n15494) );
  NAND U16062 ( .A(n182), .B(n15494), .Z(n15346) );
  AND U16063 ( .A(n15347), .B(n15346), .Z(n15501) );
  NAND U16064 ( .A(n189), .B(n15348), .Z(n15350) );
  XOR U16065 ( .A(b[17]), .B(a[102]), .Z(n15497) );
  NAND U16066 ( .A(n37652), .B(n15497), .Z(n15349) );
  NAND U16067 ( .A(n15350), .B(n15349), .Z(n15500) );
  XNOR U16068 ( .A(n15501), .B(n15500), .Z(n15502) );
  XOR U16069 ( .A(n15503), .B(n15502), .Z(n15537) );
  XOR U16070 ( .A(n15536), .B(n15537), .Z(n15539) );
  XOR U16071 ( .A(n15538), .B(n15539), .Z(n15471) );
  NANDN U16072 ( .A(n15352), .B(n15351), .Z(n15356) );
  NANDN U16073 ( .A(n15354), .B(n15353), .Z(n15355) );
  AND U16074 ( .A(n15356), .B(n15355), .Z(n15524) );
  NANDN U16075 ( .A(n15358), .B(n15357), .Z(n15362) );
  NANDN U16076 ( .A(n15360), .B(n15359), .Z(n15361) );
  NAND U16077 ( .A(n15362), .B(n15361), .Z(n15525) );
  XNOR U16078 ( .A(n15524), .B(n15525), .Z(n15526) );
  NANDN U16079 ( .A(n15364), .B(n15363), .Z(n15368) );
  NANDN U16080 ( .A(n15366), .B(n15365), .Z(n15367) );
  NAND U16081 ( .A(n15368), .B(n15367), .Z(n15527) );
  XNOR U16082 ( .A(n15526), .B(n15527), .Z(n15470) );
  XNOR U16083 ( .A(n15471), .B(n15470), .Z(n15473) );
  NANDN U16084 ( .A(n15370), .B(n15369), .Z(n15374) );
  NANDN U16085 ( .A(n15372), .B(n15371), .Z(n15373) );
  AND U16086 ( .A(n15374), .B(n15373), .Z(n15472) );
  XOR U16087 ( .A(n15473), .B(n15472), .Z(n15587) );
  NANDN U16088 ( .A(n15376), .B(n15375), .Z(n15380) );
  NANDN U16089 ( .A(n15378), .B(n15377), .Z(n15379) );
  AND U16090 ( .A(n15380), .B(n15379), .Z(n15584) );
  NANDN U16091 ( .A(n15382), .B(n15381), .Z(n15386) );
  NANDN U16092 ( .A(n15384), .B(n15383), .Z(n15385) );
  AND U16093 ( .A(n15386), .B(n15385), .Z(n15467) );
  NANDN U16094 ( .A(n15388), .B(n15387), .Z(n15392) );
  OR U16095 ( .A(n15390), .B(n15389), .Z(n15391) );
  AND U16096 ( .A(n15392), .B(n15391), .Z(n15465) );
  NANDN U16097 ( .A(n15394), .B(n15393), .Z(n15398) );
  NANDN U16098 ( .A(n15396), .B(n15395), .Z(n15397) );
  AND U16099 ( .A(n15398), .B(n15397), .Z(n15531) );
  NANDN U16100 ( .A(n15400), .B(n15399), .Z(n15404) );
  NANDN U16101 ( .A(n15402), .B(n15401), .Z(n15403) );
  NAND U16102 ( .A(n15404), .B(n15403), .Z(n15530) );
  XNOR U16103 ( .A(n15531), .B(n15530), .Z(n15532) );
  NAND U16104 ( .A(b[0]), .B(a[118]), .Z(n15405) );
  XNOR U16105 ( .A(b[1]), .B(n15405), .Z(n15407) );
  NANDN U16106 ( .A(b[0]), .B(a[117]), .Z(n15406) );
  NAND U16107 ( .A(n15407), .B(n15406), .Z(n15479) );
  NAND U16108 ( .A(n194), .B(n15408), .Z(n15410) );
  XOR U16109 ( .A(b[29]), .B(a[90]), .Z(n15557) );
  NAND U16110 ( .A(n38456), .B(n15557), .Z(n15409) );
  AND U16111 ( .A(n15410), .B(n15409), .Z(n15477) );
  AND U16112 ( .A(b[31]), .B(a[86]), .Z(n15476) );
  XNOR U16113 ( .A(n15477), .B(n15476), .Z(n15478) );
  XNOR U16114 ( .A(n15479), .B(n15478), .Z(n15518) );
  NAND U16115 ( .A(n38185), .B(n15411), .Z(n15413) );
  XOR U16116 ( .A(b[23]), .B(a[96]), .Z(n15560) );
  NAND U16117 ( .A(n38132), .B(n15560), .Z(n15412) );
  AND U16118 ( .A(n15413), .B(n15412), .Z(n15551) );
  NAND U16119 ( .A(n184), .B(n15414), .Z(n15416) );
  XOR U16120 ( .A(b[7]), .B(a[112]), .Z(n15563) );
  NAND U16121 ( .A(n36592), .B(n15563), .Z(n15415) );
  AND U16122 ( .A(n15416), .B(n15415), .Z(n15549) );
  NAND U16123 ( .A(n38289), .B(n15417), .Z(n15419) );
  XOR U16124 ( .A(b[25]), .B(a[94]), .Z(n15566) );
  NAND U16125 ( .A(n38247), .B(n15566), .Z(n15418) );
  NAND U16126 ( .A(n15419), .B(n15418), .Z(n15548) );
  XNOR U16127 ( .A(n15549), .B(n15548), .Z(n15550) );
  XOR U16128 ( .A(n15551), .B(n15550), .Z(n15519) );
  XNOR U16129 ( .A(n15518), .B(n15519), .Z(n15520) );
  NAND U16130 ( .A(n187), .B(n15420), .Z(n15422) );
  XOR U16131 ( .A(b[13]), .B(a[106]), .Z(n15569) );
  NAND U16132 ( .A(n37295), .B(n15569), .Z(n15421) );
  AND U16133 ( .A(n15422), .B(n15421), .Z(n15513) );
  NAND U16134 ( .A(n186), .B(n15423), .Z(n15425) );
  XOR U16135 ( .A(b[11]), .B(a[108]), .Z(n15572) );
  NAND U16136 ( .A(n37097), .B(n15572), .Z(n15424) );
  NAND U16137 ( .A(n15425), .B(n15424), .Z(n15512) );
  XNOR U16138 ( .A(n15513), .B(n15512), .Z(n15514) );
  NAND U16139 ( .A(n188), .B(n15426), .Z(n15428) );
  XOR U16140 ( .A(b[15]), .B(a[104]), .Z(n15575) );
  NAND U16141 ( .A(n37382), .B(n15575), .Z(n15427) );
  AND U16142 ( .A(n15428), .B(n15427), .Z(n15509) );
  NAND U16143 ( .A(n38064), .B(n15429), .Z(n15431) );
  XOR U16144 ( .A(b[21]), .B(a[98]), .Z(n15578) );
  NAND U16145 ( .A(n37993), .B(n15578), .Z(n15430) );
  AND U16146 ( .A(n15431), .B(n15430), .Z(n15507) );
  NAND U16147 ( .A(n185), .B(n15432), .Z(n15434) );
  XOR U16148 ( .A(b[9]), .B(a[110]), .Z(n15581) );
  NAND U16149 ( .A(n36805), .B(n15581), .Z(n15433) );
  NAND U16150 ( .A(n15434), .B(n15433), .Z(n15506) );
  XNOR U16151 ( .A(n15507), .B(n15506), .Z(n15508) );
  XOR U16152 ( .A(n15509), .B(n15508), .Z(n15515) );
  XOR U16153 ( .A(n15514), .B(n15515), .Z(n15521) );
  XOR U16154 ( .A(n15520), .B(n15521), .Z(n15533) );
  XNOR U16155 ( .A(n15532), .B(n15533), .Z(n15464) );
  XNOR U16156 ( .A(n15465), .B(n15464), .Z(n15466) );
  XOR U16157 ( .A(n15467), .B(n15466), .Z(n15585) );
  XNOR U16158 ( .A(n15584), .B(n15585), .Z(n15586) );
  XNOR U16159 ( .A(n15587), .B(n15586), .Z(n15460) );
  XOR U16160 ( .A(n15461), .B(n15460), .Z(n15453) );
  NANDN U16161 ( .A(n15436), .B(n15435), .Z(n15440) );
  NANDN U16162 ( .A(n15438), .B(n15437), .Z(n15439) );
  AND U16163 ( .A(n15440), .B(n15439), .Z(n15452) );
  XOR U16164 ( .A(n15453), .B(n15452), .Z(n15455) );
  XNOR U16165 ( .A(n15454), .B(n15455), .Z(n15446) );
  XNOR U16166 ( .A(n15447), .B(n15446), .Z(n15448) );
  XNOR U16167 ( .A(n15449), .B(n15448), .Z(n15590) );
  XNOR U16168 ( .A(sreg[342]), .B(n15590), .Z(n15592) );
  NANDN U16169 ( .A(sreg[341]), .B(n15441), .Z(n15445) );
  NAND U16170 ( .A(n15443), .B(n15442), .Z(n15444) );
  NAND U16171 ( .A(n15445), .B(n15444), .Z(n15591) );
  XNOR U16172 ( .A(n15592), .B(n15591), .Z(c[342]) );
  NANDN U16173 ( .A(n15447), .B(n15446), .Z(n15451) );
  NANDN U16174 ( .A(n15449), .B(n15448), .Z(n15450) );
  AND U16175 ( .A(n15451), .B(n15450), .Z(n15602) );
  NANDN U16176 ( .A(n15453), .B(n15452), .Z(n15457) );
  NANDN U16177 ( .A(n15455), .B(n15454), .Z(n15456) );
  AND U16178 ( .A(n15457), .B(n15456), .Z(n15601) );
  NANDN U16179 ( .A(n15459), .B(n15458), .Z(n15463) );
  NAND U16180 ( .A(n15461), .B(n15460), .Z(n15462) );
  AND U16181 ( .A(n15463), .B(n15462), .Z(n15608) );
  NANDN U16182 ( .A(n15465), .B(n15464), .Z(n15469) );
  NANDN U16183 ( .A(n15467), .B(n15466), .Z(n15468) );
  AND U16184 ( .A(n15469), .B(n15468), .Z(n15739) );
  NANDN U16185 ( .A(n15471), .B(n15470), .Z(n15475) );
  NAND U16186 ( .A(n15473), .B(n15472), .Z(n15474) );
  AND U16187 ( .A(n15475), .B(n15474), .Z(n15738) );
  XNOR U16188 ( .A(n15739), .B(n15738), .Z(n15741) );
  NANDN U16189 ( .A(n15477), .B(n15476), .Z(n15481) );
  NANDN U16190 ( .A(n15479), .B(n15478), .Z(n15480) );
  AND U16191 ( .A(n15481), .B(n15480), .Z(n15686) );
  NAND U16192 ( .A(n38385), .B(n15482), .Z(n15484) );
  XOR U16193 ( .A(b[27]), .B(a[93]), .Z(n15630) );
  NAND U16194 ( .A(n38343), .B(n15630), .Z(n15483) );
  AND U16195 ( .A(n15484), .B(n15483), .Z(n15693) );
  NAND U16196 ( .A(n183), .B(n15485), .Z(n15487) );
  XOR U16197 ( .A(b[5]), .B(a[115]), .Z(n15633) );
  NAND U16198 ( .A(n36296), .B(n15633), .Z(n15486) );
  AND U16199 ( .A(n15487), .B(n15486), .Z(n15691) );
  NAND U16200 ( .A(n190), .B(n15488), .Z(n15490) );
  XOR U16201 ( .A(b[19]), .B(a[101]), .Z(n15636) );
  NAND U16202 ( .A(n37821), .B(n15636), .Z(n15489) );
  NAND U16203 ( .A(n15490), .B(n15489), .Z(n15690) );
  XNOR U16204 ( .A(n15691), .B(n15690), .Z(n15692) );
  XNOR U16205 ( .A(n15693), .B(n15692), .Z(n15684) );
  NAND U16206 ( .A(n38470), .B(n15491), .Z(n15493) );
  XOR U16207 ( .A(b[31]), .B(a[89]), .Z(n15639) );
  NAND U16208 ( .A(n38453), .B(n15639), .Z(n15492) );
  AND U16209 ( .A(n15493), .B(n15492), .Z(n15651) );
  NAND U16210 ( .A(n181), .B(n15494), .Z(n15496) );
  XOR U16211 ( .A(b[3]), .B(a[117]), .Z(n15642) );
  NAND U16212 ( .A(n182), .B(n15642), .Z(n15495) );
  AND U16213 ( .A(n15496), .B(n15495), .Z(n15649) );
  NAND U16214 ( .A(n189), .B(n15497), .Z(n15499) );
  XOR U16215 ( .A(b[17]), .B(a[103]), .Z(n15645) );
  NAND U16216 ( .A(n37652), .B(n15645), .Z(n15498) );
  NAND U16217 ( .A(n15499), .B(n15498), .Z(n15648) );
  XNOR U16218 ( .A(n15649), .B(n15648), .Z(n15650) );
  XOR U16219 ( .A(n15651), .B(n15650), .Z(n15685) );
  XOR U16220 ( .A(n15684), .B(n15685), .Z(n15687) );
  XOR U16221 ( .A(n15686), .B(n15687), .Z(n15619) );
  NANDN U16222 ( .A(n15501), .B(n15500), .Z(n15505) );
  NANDN U16223 ( .A(n15503), .B(n15502), .Z(n15504) );
  AND U16224 ( .A(n15505), .B(n15504), .Z(n15672) );
  NANDN U16225 ( .A(n15507), .B(n15506), .Z(n15511) );
  NANDN U16226 ( .A(n15509), .B(n15508), .Z(n15510) );
  NAND U16227 ( .A(n15511), .B(n15510), .Z(n15673) );
  XNOR U16228 ( .A(n15672), .B(n15673), .Z(n15674) );
  NANDN U16229 ( .A(n15513), .B(n15512), .Z(n15517) );
  NANDN U16230 ( .A(n15515), .B(n15514), .Z(n15516) );
  NAND U16231 ( .A(n15517), .B(n15516), .Z(n15675) );
  XNOR U16232 ( .A(n15674), .B(n15675), .Z(n15618) );
  XNOR U16233 ( .A(n15619), .B(n15618), .Z(n15621) );
  NANDN U16234 ( .A(n15519), .B(n15518), .Z(n15523) );
  NANDN U16235 ( .A(n15521), .B(n15520), .Z(n15522) );
  AND U16236 ( .A(n15523), .B(n15522), .Z(n15620) );
  XOR U16237 ( .A(n15621), .B(n15620), .Z(n15735) );
  NANDN U16238 ( .A(n15525), .B(n15524), .Z(n15529) );
  NANDN U16239 ( .A(n15527), .B(n15526), .Z(n15528) );
  AND U16240 ( .A(n15529), .B(n15528), .Z(n15732) );
  NANDN U16241 ( .A(n15531), .B(n15530), .Z(n15535) );
  NANDN U16242 ( .A(n15533), .B(n15532), .Z(n15534) );
  AND U16243 ( .A(n15535), .B(n15534), .Z(n15615) );
  NANDN U16244 ( .A(n15537), .B(n15536), .Z(n15541) );
  OR U16245 ( .A(n15539), .B(n15538), .Z(n15540) );
  AND U16246 ( .A(n15541), .B(n15540), .Z(n15613) );
  NANDN U16247 ( .A(n15543), .B(n15542), .Z(n15547) );
  NANDN U16248 ( .A(n15545), .B(n15544), .Z(n15546) );
  AND U16249 ( .A(n15547), .B(n15546), .Z(n15679) );
  NANDN U16250 ( .A(n15549), .B(n15548), .Z(n15553) );
  NANDN U16251 ( .A(n15551), .B(n15550), .Z(n15552) );
  NAND U16252 ( .A(n15553), .B(n15552), .Z(n15678) );
  XNOR U16253 ( .A(n15679), .B(n15678), .Z(n15680) );
  NAND U16254 ( .A(b[0]), .B(a[119]), .Z(n15554) );
  XNOR U16255 ( .A(b[1]), .B(n15554), .Z(n15556) );
  NANDN U16256 ( .A(b[0]), .B(a[118]), .Z(n15555) );
  NAND U16257 ( .A(n15556), .B(n15555), .Z(n15627) );
  NAND U16258 ( .A(n194), .B(n15557), .Z(n15559) );
  XOR U16259 ( .A(b[29]), .B(a[91]), .Z(n15705) );
  NAND U16260 ( .A(n38456), .B(n15705), .Z(n15558) );
  AND U16261 ( .A(n15559), .B(n15558), .Z(n15625) );
  AND U16262 ( .A(b[31]), .B(a[87]), .Z(n15624) );
  XNOR U16263 ( .A(n15625), .B(n15624), .Z(n15626) );
  XNOR U16264 ( .A(n15627), .B(n15626), .Z(n15666) );
  NAND U16265 ( .A(n38185), .B(n15560), .Z(n15562) );
  XOR U16266 ( .A(b[23]), .B(a[97]), .Z(n15708) );
  NAND U16267 ( .A(n38132), .B(n15708), .Z(n15561) );
  AND U16268 ( .A(n15562), .B(n15561), .Z(n15699) );
  NAND U16269 ( .A(n184), .B(n15563), .Z(n15565) );
  XOR U16270 ( .A(b[7]), .B(a[113]), .Z(n15711) );
  NAND U16271 ( .A(n36592), .B(n15711), .Z(n15564) );
  AND U16272 ( .A(n15565), .B(n15564), .Z(n15697) );
  NAND U16273 ( .A(n38289), .B(n15566), .Z(n15568) );
  XOR U16274 ( .A(b[25]), .B(a[95]), .Z(n15714) );
  NAND U16275 ( .A(n38247), .B(n15714), .Z(n15567) );
  NAND U16276 ( .A(n15568), .B(n15567), .Z(n15696) );
  XNOR U16277 ( .A(n15697), .B(n15696), .Z(n15698) );
  XOR U16278 ( .A(n15699), .B(n15698), .Z(n15667) );
  XNOR U16279 ( .A(n15666), .B(n15667), .Z(n15668) );
  NAND U16280 ( .A(n187), .B(n15569), .Z(n15571) );
  XOR U16281 ( .A(b[13]), .B(a[107]), .Z(n15717) );
  NAND U16282 ( .A(n37295), .B(n15717), .Z(n15570) );
  AND U16283 ( .A(n15571), .B(n15570), .Z(n15661) );
  NAND U16284 ( .A(n186), .B(n15572), .Z(n15574) );
  XOR U16285 ( .A(b[11]), .B(a[109]), .Z(n15720) );
  NAND U16286 ( .A(n37097), .B(n15720), .Z(n15573) );
  NAND U16287 ( .A(n15574), .B(n15573), .Z(n15660) );
  XNOR U16288 ( .A(n15661), .B(n15660), .Z(n15662) );
  NAND U16289 ( .A(n188), .B(n15575), .Z(n15577) );
  XOR U16290 ( .A(b[15]), .B(a[105]), .Z(n15723) );
  NAND U16291 ( .A(n37382), .B(n15723), .Z(n15576) );
  AND U16292 ( .A(n15577), .B(n15576), .Z(n15657) );
  NAND U16293 ( .A(n38064), .B(n15578), .Z(n15580) );
  XOR U16294 ( .A(b[21]), .B(a[99]), .Z(n15726) );
  NAND U16295 ( .A(n37993), .B(n15726), .Z(n15579) );
  AND U16296 ( .A(n15580), .B(n15579), .Z(n15655) );
  NAND U16297 ( .A(n185), .B(n15581), .Z(n15583) );
  XOR U16298 ( .A(b[9]), .B(a[111]), .Z(n15729) );
  NAND U16299 ( .A(n36805), .B(n15729), .Z(n15582) );
  NAND U16300 ( .A(n15583), .B(n15582), .Z(n15654) );
  XNOR U16301 ( .A(n15655), .B(n15654), .Z(n15656) );
  XOR U16302 ( .A(n15657), .B(n15656), .Z(n15663) );
  XOR U16303 ( .A(n15662), .B(n15663), .Z(n15669) );
  XOR U16304 ( .A(n15668), .B(n15669), .Z(n15681) );
  XNOR U16305 ( .A(n15680), .B(n15681), .Z(n15612) );
  XNOR U16306 ( .A(n15613), .B(n15612), .Z(n15614) );
  XOR U16307 ( .A(n15615), .B(n15614), .Z(n15733) );
  XNOR U16308 ( .A(n15732), .B(n15733), .Z(n15734) );
  XNOR U16309 ( .A(n15735), .B(n15734), .Z(n15740) );
  XOR U16310 ( .A(n15741), .B(n15740), .Z(n15607) );
  NANDN U16311 ( .A(n15585), .B(n15584), .Z(n15589) );
  NANDN U16312 ( .A(n15587), .B(n15586), .Z(n15588) );
  AND U16313 ( .A(n15589), .B(n15588), .Z(n15606) );
  XOR U16314 ( .A(n15607), .B(n15606), .Z(n15609) );
  XNOR U16315 ( .A(n15608), .B(n15609), .Z(n15600) );
  XOR U16316 ( .A(n15601), .B(n15600), .Z(n15603) );
  XOR U16317 ( .A(n15602), .B(n15603), .Z(n15595) );
  XNOR U16318 ( .A(n15595), .B(sreg[343]), .Z(n15597) );
  NANDN U16319 ( .A(sreg[342]), .B(n15590), .Z(n15594) );
  NAND U16320 ( .A(n15592), .B(n15591), .Z(n15593) );
  AND U16321 ( .A(n15594), .B(n15593), .Z(n15596) );
  XOR U16322 ( .A(n15597), .B(n15596), .Z(c[343]) );
  NANDN U16323 ( .A(n15595), .B(sreg[343]), .Z(n15599) );
  NAND U16324 ( .A(n15597), .B(n15596), .Z(n15598) );
  AND U16325 ( .A(n15599), .B(n15598), .Z(n15888) );
  NANDN U16326 ( .A(n15601), .B(n15600), .Z(n15605) );
  OR U16327 ( .A(n15603), .B(n15602), .Z(n15604) );
  AND U16328 ( .A(n15605), .B(n15604), .Z(n15747) );
  NANDN U16329 ( .A(n15607), .B(n15606), .Z(n15611) );
  NANDN U16330 ( .A(n15609), .B(n15608), .Z(n15610) );
  AND U16331 ( .A(n15611), .B(n15610), .Z(n15745) );
  NANDN U16332 ( .A(n15613), .B(n15612), .Z(n15617) );
  NANDN U16333 ( .A(n15615), .B(n15614), .Z(n15616) );
  AND U16334 ( .A(n15617), .B(n15616), .Z(n15757) );
  NANDN U16335 ( .A(n15619), .B(n15618), .Z(n15623) );
  NAND U16336 ( .A(n15621), .B(n15620), .Z(n15622) );
  AND U16337 ( .A(n15623), .B(n15622), .Z(n15756) );
  XNOR U16338 ( .A(n15757), .B(n15756), .Z(n15759) );
  NANDN U16339 ( .A(n15625), .B(n15624), .Z(n15629) );
  NANDN U16340 ( .A(n15627), .B(n15626), .Z(n15628) );
  AND U16341 ( .A(n15629), .B(n15628), .Z(n15834) );
  NAND U16342 ( .A(n38385), .B(n15630), .Z(n15632) );
  XOR U16343 ( .A(b[27]), .B(a[94]), .Z(n15780) );
  NAND U16344 ( .A(n38343), .B(n15780), .Z(n15631) );
  AND U16345 ( .A(n15632), .B(n15631), .Z(n15841) );
  NAND U16346 ( .A(n183), .B(n15633), .Z(n15635) );
  XOR U16347 ( .A(b[5]), .B(a[116]), .Z(n15783) );
  NAND U16348 ( .A(n36296), .B(n15783), .Z(n15634) );
  AND U16349 ( .A(n15635), .B(n15634), .Z(n15839) );
  NAND U16350 ( .A(n190), .B(n15636), .Z(n15638) );
  XOR U16351 ( .A(b[19]), .B(a[102]), .Z(n15786) );
  NAND U16352 ( .A(n37821), .B(n15786), .Z(n15637) );
  NAND U16353 ( .A(n15638), .B(n15637), .Z(n15838) );
  XNOR U16354 ( .A(n15839), .B(n15838), .Z(n15840) );
  XNOR U16355 ( .A(n15841), .B(n15840), .Z(n15832) );
  NAND U16356 ( .A(n38470), .B(n15639), .Z(n15641) );
  XOR U16357 ( .A(b[31]), .B(a[90]), .Z(n15789) );
  NAND U16358 ( .A(n38453), .B(n15789), .Z(n15640) );
  AND U16359 ( .A(n15641), .B(n15640), .Z(n15801) );
  NAND U16360 ( .A(n181), .B(n15642), .Z(n15644) );
  XOR U16361 ( .A(b[3]), .B(a[118]), .Z(n15792) );
  NAND U16362 ( .A(n182), .B(n15792), .Z(n15643) );
  AND U16363 ( .A(n15644), .B(n15643), .Z(n15799) );
  NAND U16364 ( .A(n189), .B(n15645), .Z(n15647) );
  XOR U16365 ( .A(b[17]), .B(a[104]), .Z(n15795) );
  NAND U16366 ( .A(n37652), .B(n15795), .Z(n15646) );
  NAND U16367 ( .A(n15647), .B(n15646), .Z(n15798) );
  XNOR U16368 ( .A(n15799), .B(n15798), .Z(n15800) );
  XOR U16369 ( .A(n15801), .B(n15800), .Z(n15833) );
  XOR U16370 ( .A(n15832), .B(n15833), .Z(n15835) );
  XOR U16371 ( .A(n15834), .B(n15835), .Z(n15769) );
  NANDN U16372 ( .A(n15649), .B(n15648), .Z(n15653) );
  NANDN U16373 ( .A(n15651), .B(n15650), .Z(n15652) );
  AND U16374 ( .A(n15653), .B(n15652), .Z(n15822) );
  NANDN U16375 ( .A(n15655), .B(n15654), .Z(n15659) );
  NANDN U16376 ( .A(n15657), .B(n15656), .Z(n15658) );
  NAND U16377 ( .A(n15659), .B(n15658), .Z(n15823) );
  XNOR U16378 ( .A(n15822), .B(n15823), .Z(n15824) );
  NANDN U16379 ( .A(n15661), .B(n15660), .Z(n15665) );
  NANDN U16380 ( .A(n15663), .B(n15662), .Z(n15664) );
  NAND U16381 ( .A(n15665), .B(n15664), .Z(n15825) );
  XNOR U16382 ( .A(n15824), .B(n15825), .Z(n15768) );
  XNOR U16383 ( .A(n15769), .B(n15768), .Z(n15771) );
  NANDN U16384 ( .A(n15667), .B(n15666), .Z(n15671) );
  NANDN U16385 ( .A(n15669), .B(n15668), .Z(n15670) );
  AND U16386 ( .A(n15671), .B(n15670), .Z(n15770) );
  XOR U16387 ( .A(n15771), .B(n15770), .Z(n15883) );
  NANDN U16388 ( .A(n15673), .B(n15672), .Z(n15677) );
  NANDN U16389 ( .A(n15675), .B(n15674), .Z(n15676) );
  AND U16390 ( .A(n15677), .B(n15676), .Z(n15880) );
  NANDN U16391 ( .A(n15679), .B(n15678), .Z(n15683) );
  NANDN U16392 ( .A(n15681), .B(n15680), .Z(n15682) );
  AND U16393 ( .A(n15683), .B(n15682), .Z(n15765) );
  NANDN U16394 ( .A(n15685), .B(n15684), .Z(n15689) );
  OR U16395 ( .A(n15687), .B(n15686), .Z(n15688) );
  AND U16396 ( .A(n15689), .B(n15688), .Z(n15763) );
  NANDN U16397 ( .A(n15691), .B(n15690), .Z(n15695) );
  NANDN U16398 ( .A(n15693), .B(n15692), .Z(n15694) );
  AND U16399 ( .A(n15695), .B(n15694), .Z(n15829) );
  NANDN U16400 ( .A(n15697), .B(n15696), .Z(n15701) );
  NANDN U16401 ( .A(n15699), .B(n15698), .Z(n15700) );
  NAND U16402 ( .A(n15701), .B(n15700), .Z(n15828) );
  XNOR U16403 ( .A(n15829), .B(n15828), .Z(n15831) );
  NAND U16404 ( .A(b[0]), .B(a[120]), .Z(n15702) );
  XNOR U16405 ( .A(b[1]), .B(n15702), .Z(n15704) );
  NANDN U16406 ( .A(b[0]), .B(a[119]), .Z(n15703) );
  NAND U16407 ( .A(n15704), .B(n15703), .Z(n15777) );
  NAND U16408 ( .A(n194), .B(n15705), .Z(n15707) );
  XOR U16409 ( .A(b[29]), .B(a[92]), .Z(n15853) );
  NAND U16410 ( .A(n38456), .B(n15853), .Z(n15706) );
  AND U16411 ( .A(n15707), .B(n15706), .Z(n15775) );
  AND U16412 ( .A(b[31]), .B(a[88]), .Z(n15774) );
  XNOR U16413 ( .A(n15775), .B(n15774), .Z(n15776) );
  XNOR U16414 ( .A(n15777), .B(n15776), .Z(n15817) );
  NAND U16415 ( .A(n38185), .B(n15708), .Z(n15710) );
  XOR U16416 ( .A(b[23]), .B(a[98]), .Z(n15856) );
  NAND U16417 ( .A(n38132), .B(n15856), .Z(n15709) );
  AND U16418 ( .A(n15710), .B(n15709), .Z(n15846) );
  NAND U16419 ( .A(n184), .B(n15711), .Z(n15713) );
  XOR U16420 ( .A(b[7]), .B(a[114]), .Z(n15859) );
  NAND U16421 ( .A(n36592), .B(n15859), .Z(n15712) );
  AND U16422 ( .A(n15713), .B(n15712), .Z(n15845) );
  NAND U16423 ( .A(n38289), .B(n15714), .Z(n15716) );
  XOR U16424 ( .A(b[25]), .B(a[96]), .Z(n15862) );
  NAND U16425 ( .A(n38247), .B(n15862), .Z(n15715) );
  NAND U16426 ( .A(n15716), .B(n15715), .Z(n15844) );
  XOR U16427 ( .A(n15845), .B(n15844), .Z(n15847) );
  XOR U16428 ( .A(n15846), .B(n15847), .Z(n15816) );
  XOR U16429 ( .A(n15817), .B(n15816), .Z(n15819) );
  NAND U16430 ( .A(n187), .B(n15717), .Z(n15719) );
  XOR U16431 ( .A(b[13]), .B(a[108]), .Z(n15865) );
  NAND U16432 ( .A(n37295), .B(n15865), .Z(n15718) );
  AND U16433 ( .A(n15719), .B(n15718), .Z(n15811) );
  NAND U16434 ( .A(n186), .B(n15720), .Z(n15722) );
  XOR U16435 ( .A(b[11]), .B(a[110]), .Z(n15868) );
  NAND U16436 ( .A(n37097), .B(n15868), .Z(n15721) );
  NAND U16437 ( .A(n15722), .B(n15721), .Z(n15810) );
  XNOR U16438 ( .A(n15811), .B(n15810), .Z(n15813) );
  NAND U16439 ( .A(n188), .B(n15723), .Z(n15725) );
  XOR U16440 ( .A(b[15]), .B(a[106]), .Z(n15871) );
  NAND U16441 ( .A(n37382), .B(n15871), .Z(n15724) );
  AND U16442 ( .A(n15725), .B(n15724), .Z(n15807) );
  NAND U16443 ( .A(n38064), .B(n15726), .Z(n15728) );
  XOR U16444 ( .A(b[21]), .B(a[100]), .Z(n15874) );
  NAND U16445 ( .A(n37993), .B(n15874), .Z(n15727) );
  AND U16446 ( .A(n15728), .B(n15727), .Z(n15805) );
  NAND U16447 ( .A(n185), .B(n15729), .Z(n15731) );
  XOR U16448 ( .A(b[9]), .B(a[112]), .Z(n15877) );
  NAND U16449 ( .A(n36805), .B(n15877), .Z(n15730) );
  NAND U16450 ( .A(n15731), .B(n15730), .Z(n15804) );
  XNOR U16451 ( .A(n15805), .B(n15804), .Z(n15806) );
  XNOR U16452 ( .A(n15807), .B(n15806), .Z(n15812) );
  XOR U16453 ( .A(n15813), .B(n15812), .Z(n15818) );
  XNOR U16454 ( .A(n15819), .B(n15818), .Z(n15830) );
  XNOR U16455 ( .A(n15831), .B(n15830), .Z(n15762) );
  XNOR U16456 ( .A(n15763), .B(n15762), .Z(n15764) );
  XOR U16457 ( .A(n15765), .B(n15764), .Z(n15881) );
  XNOR U16458 ( .A(n15880), .B(n15881), .Z(n15882) );
  XNOR U16459 ( .A(n15883), .B(n15882), .Z(n15758) );
  XOR U16460 ( .A(n15759), .B(n15758), .Z(n15751) );
  NANDN U16461 ( .A(n15733), .B(n15732), .Z(n15737) );
  NANDN U16462 ( .A(n15735), .B(n15734), .Z(n15736) );
  AND U16463 ( .A(n15737), .B(n15736), .Z(n15750) );
  XNOR U16464 ( .A(n15751), .B(n15750), .Z(n15752) );
  NANDN U16465 ( .A(n15739), .B(n15738), .Z(n15743) );
  NAND U16466 ( .A(n15741), .B(n15740), .Z(n15742) );
  NAND U16467 ( .A(n15743), .B(n15742), .Z(n15753) );
  XNOR U16468 ( .A(n15752), .B(n15753), .Z(n15744) );
  XNOR U16469 ( .A(n15745), .B(n15744), .Z(n15746) );
  XNOR U16470 ( .A(n15747), .B(n15746), .Z(n15886) );
  XNOR U16471 ( .A(sreg[344]), .B(n15886), .Z(n15887) );
  XNOR U16472 ( .A(n15888), .B(n15887), .Z(c[344]) );
  NANDN U16473 ( .A(n15745), .B(n15744), .Z(n15749) );
  NANDN U16474 ( .A(n15747), .B(n15746), .Z(n15748) );
  AND U16475 ( .A(n15749), .B(n15748), .Z(n15894) );
  NANDN U16476 ( .A(n15751), .B(n15750), .Z(n15755) );
  NANDN U16477 ( .A(n15753), .B(n15752), .Z(n15754) );
  AND U16478 ( .A(n15755), .B(n15754), .Z(n15892) );
  NANDN U16479 ( .A(n15757), .B(n15756), .Z(n15761) );
  NAND U16480 ( .A(n15759), .B(n15758), .Z(n15760) );
  AND U16481 ( .A(n15761), .B(n15760), .Z(n15899) );
  NANDN U16482 ( .A(n15763), .B(n15762), .Z(n15767) );
  NANDN U16483 ( .A(n15765), .B(n15764), .Z(n15766) );
  AND U16484 ( .A(n15767), .B(n15766), .Z(n16030) );
  NANDN U16485 ( .A(n15769), .B(n15768), .Z(n15773) );
  NAND U16486 ( .A(n15771), .B(n15770), .Z(n15772) );
  AND U16487 ( .A(n15773), .B(n15772), .Z(n16029) );
  XNOR U16488 ( .A(n16030), .B(n16029), .Z(n16032) );
  NANDN U16489 ( .A(n15775), .B(n15774), .Z(n15779) );
  NANDN U16490 ( .A(n15777), .B(n15776), .Z(n15778) );
  AND U16491 ( .A(n15779), .B(n15778), .Z(n15965) );
  NAND U16492 ( .A(n38385), .B(n15780), .Z(n15782) );
  XOR U16493 ( .A(b[27]), .B(a[95]), .Z(n15909) );
  NAND U16494 ( .A(n38343), .B(n15909), .Z(n15781) );
  AND U16495 ( .A(n15782), .B(n15781), .Z(n15972) );
  NAND U16496 ( .A(n183), .B(n15783), .Z(n15785) );
  XOR U16497 ( .A(b[5]), .B(a[117]), .Z(n15912) );
  NAND U16498 ( .A(n36296), .B(n15912), .Z(n15784) );
  AND U16499 ( .A(n15785), .B(n15784), .Z(n15970) );
  NAND U16500 ( .A(n190), .B(n15786), .Z(n15788) );
  XOR U16501 ( .A(b[19]), .B(a[103]), .Z(n15915) );
  NAND U16502 ( .A(n37821), .B(n15915), .Z(n15787) );
  NAND U16503 ( .A(n15788), .B(n15787), .Z(n15969) );
  XNOR U16504 ( .A(n15970), .B(n15969), .Z(n15971) );
  XNOR U16505 ( .A(n15972), .B(n15971), .Z(n15963) );
  NAND U16506 ( .A(n38470), .B(n15789), .Z(n15791) );
  XOR U16507 ( .A(b[31]), .B(a[91]), .Z(n15918) );
  NAND U16508 ( .A(n38453), .B(n15918), .Z(n15790) );
  AND U16509 ( .A(n15791), .B(n15790), .Z(n15930) );
  NAND U16510 ( .A(n181), .B(n15792), .Z(n15794) );
  XOR U16511 ( .A(b[3]), .B(a[119]), .Z(n15921) );
  NAND U16512 ( .A(n182), .B(n15921), .Z(n15793) );
  AND U16513 ( .A(n15794), .B(n15793), .Z(n15928) );
  NAND U16514 ( .A(n189), .B(n15795), .Z(n15797) );
  XOR U16515 ( .A(b[17]), .B(a[105]), .Z(n15924) );
  NAND U16516 ( .A(n37652), .B(n15924), .Z(n15796) );
  NAND U16517 ( .A(n15797), .B(n15796), .Z(n15927) );
  XNOR U16518 ( .A(n15928), .B(n15927), .Z(n15929) );
  XOR U16519 ( .A(n15930), .B(n15929), .Z(n15964) );
  XOR U16520 ( .A(n15963), .B(n15964), .Z(n15966) );
  XOR U16521 ( .A(n15965), .B(n15966), .Z(n16012) );
  NANDN U16522 ( .A(n15799), .B(n15798), .Z(n15803) );
  NANDN U16523 ( .A(n15801), .B(n15800), .Z(n15802) );
  AND U16524 ( .A(n15803), .B(n15802), .Z(n15951) );
  NANDN U16525 ( .A(n15805), .B(n15804), .Z(n15809) );
  NANDN U16526 ( .A(n15807), .B(n15806), .Z(n15808) );
  NAND U16527 ( .A(n15809), .B(n15808), .Z(n15952) );
  XNOR U16528 ( .A(n15951), .B(n15952), .Z(n15953) );
  NANDN U16529 ( .A(n15811), .B(n15810), .Z(n15815) );
  NAND U16530 ( .A(n15813), .B(n15812), .Z(n15814) );
  NAND U16531 ( .A(n15815), .B(n15814), .Z(n15954) );
  XNOR U16532 ( .A(n15953), .B(n15954), .Z(n16011) );
  XNOR U16533 ( .A(n16012), .B(n16011), .Z(n16014) );
  NAND U16534 ( .A(n15817), .B(n15816), .Z(n15821) );
  NAND U16535 ( .A(n15819), .B(n15818), .Z(n15820) );
  AND U16536 ( .A(n15821), .B(n15820), .Z(n16013) );
  XOR U16537 ( .A(n16014), .B(n16013), .Z(n16026) );
  NANDN U16538 ( .A(n15823), .B(n15822), .Z(n15827) );
  NANDN U16539 ( .A(n15825), .B(n15824), .Z(n15826) );
  AND U16540 ( .A(n15827), .B(n15826), .Z(n16023) );
  NANDN U16541 ( .A(n15833), .B(n15832), .Z(n15837) );
  OR U16542 ( .A(n15835), .B(n15834), .Z(n15836) );
  AND U16543 ( .A(n15837), .B(n15836), .Z(n16018) );
  NANDN U16544 ( .A(n15839), .B(n15838), .Z(n15843) );
  NANDN U16545 ( .A(n15841), .B(n15840), .Z(n15842) );
  AND U16546 ( .A(n15843), .B(n15842), .Z(n15958) );
  NANDN U16547 ( .A(n15845), .B(n15844), .Z(n15849) );
  OR U16548 ( .A(n15847), .B(n15846), .Z(n15848) );
  NAND U16549 ( .A(n15849), .B(n15848), .Z(n15957) );
  XNOR U16550 ( .A(n15958), .B(n15957), .Z(n15959) );
  NAND U16551 ( .A(b[0]), .B(a[121]), .Z(n15850) );
  XNOR U16552 ( .A(b[1]), .B(n15850), .Z(n15852) );
  NANDN U16553 ( .A(b[0]), .B(a[120]), .Z(n15851) );
  NAND U16554 ( .A(n15852), .B(n15851), .Z(n15906) );
  NAND U16555 ( .A(n194), .B(n15853), .Z(n15855) );
  XOR U16556 ( .A(b[29]), .B(a[93]), .Z(n15984) );
  NAND U16557 ( .A(n38456), .B(n15984), .Z(n15854) );
  AND U16558 ( .A(n15855), .B(n15854), .Z(n15904) );
  AND U16559 ( .A(b[31]), .B(a[89]), .Z(n15903) );
  XNOR U16560 ( .A(n15904), .B(n15903), .Z(n15905) );
  XNOR U16561 ( .A(n15906), .B(n15905), .Z(n15945) );
  NAND U16562 ( .A(n38185), .B(n15856), .Z(n15858) );
  XOR U16563 ( .A(b[23]), .B(a[99]), .Z(n15987) );
  NAND U16564 ( .A(n38132), .B(n15987), .Z(n15857) );
  AND U16565 ( .A(n15858), .B(n15857), .Z(n15978) );
  NAND U16566 ( .A(n184), .B(n15859), .Z(n15861) );
  XOR U16567 ( .A(b[7]), .B(a[115]), .Z(n15990) );
  NAND U16568 ( .A(n36592), .B(n15990), .Z(n15860) );
  AND U16569 ( .A(n15861), .B(n15860), .Z(n15976) );
  NAND U16570 ( .A(n38289), .B(n15862), .Z(n15864) );
  XOR U16571 ( .A(b[25]), .B(a[97]), .Z(n15993) );
  NAND U16572 ( .A(n38247), .B(n15993), .Z(n15863) );
  NAND U16573 ( .A(n15864), .B(n15863), .Z(n15975) );
  XNOR U16574 ( .A(n15976), .B(n15975), .Z(n15977) );
  XOR U16575 ( .A(n15978), .B(n15977), .Z(n15946) );
  XNOR U16576 ( .A(n15945), .B(n15946), .Z(n15947) );
  NAND U16577 ( .A(n187), .B(n15865), .Z(n15867) );
  XOR U16578 ( .A(b[13]), .B(a[109]), .Z(n15996) );
  NAND U16579 ( .A(n37295), .B(n15996), .Z(n15866) );
  AND U16580 ( .A(n15867), .B(n15866), .Z(n15940) );
  NAND U16581 ( .A(n186), .B(n15868), .Z(n15870) );
  XOR U16582 ( .A(b[11]), .B(a[111]), .Z(n15999) );
  NAND U16583 ( .A(n37097), .B(n15999), .Z(n15869) );
  NAND U16584 ( .A(n15870), .B(n15869), .Z(n15939) );
  XNOR U16585 ( .A(n15940), .B(n15939), .Z(n15941) );
  NAND U16586 ( .A(n188), .B(n15871), .Z(n15873) );
  XOR U16587 ( .A(b[15]), .B(a[107]), .Z(n16002) );
  NAND U16588 ( .A(n37382), .B(n16002), .Z(n15872) );
  AND U16589 ( .A(n15873), .B(n15872), .Z(n15936) );
  NAND U16590 ( .A(n38064), .B(n15874), .Z(n15876) );
  XOR U16591 ( .A(b[21]), .B(a[101]), .Z(n16005) );
  NAND U16592 ( .A(n37993), .B(n16005), .Z(n15875) );
  AND U16593 ( .A(n15876), .B(n15875), .Z(n15934) );
  NAND U16594 ( .A(n185), .B(n15877), .Z(n15879) );
  XOR U16595 ( .A(b[9]), .B(a[113]), .Z(n16008) );
  NAND U16596 ( .A(n36805), .B(n16008), .Z(n15878) );
  NAND U16597 ( .A(n15879), .B(n15878), .Z(n15933) );
  XNOR U16598 ( .A(n15934), .B(n15933), .Z(n15935) );
  XOR U16599 ( .A(n15936), .B(n15935), .Z(n15942) );
  XOR U16600 ( .A(n15941), .B(n15942), .Z(n15948) );
  XOR U16601 ( .A(n15947), .B(n15948), .Z(n15960) );
  XNOR U16602 ( .A(n15959), .B(n15960), .Z(n16017) );
  XNOR U16603 ( .A(n16018), .B(n16017), .Z(n16019) );
  XOR U16604 ( .A(n16020), .B(n16019), .Z(n16024) );
  XNOR U16605 ( .A(n16023), .B(n16024), .Z(n16025) );
  XNOR U16606 ( .A(n16026), .B(n16025), .Z(n16031) );
  XOR U16607 ( .A(n16032), .B(n16031), .Z(n15898) );
  NANDN U16608 ( .A(n15881), .B(n15880), .Z(n15885) );
  NANDN U16609 ( .A(n15883), .B(n15882), .Z(n15884) );
  AND U16610 ( .A(n15885), .B(n15884), .Z(n15897) );
  XOR U16611 ( .A(n15898), .B(n15897), .Z(n15900) );
  XNOR U16612 ( .A(n15899), .B(n15900), .Z(n15891) );
  XNOR U16613 ( .A(n15892), .B(n15891), .Z(n15893) );
  XNOR U16614 ( .A(n15894), .B(n15893), .Z(n16035) );
  XNOR U16615 ( .A(sreg[345]), .B(n16035), .Z(n16037) );
  NANDN U16616 ( .A(sreg[344]), .B(n15886), .Z(n15890) );
  NAND U16617 ( .A(n15888), .B(n15887), .Z(n15889) );
  NAND U16618 ( .A(n15890), .B(n15889), .Z(n16036) );
  XNOR U16619 ( .A(n16037), .B(n16036), .Z(c[345]) );
  NANDN U16620 ( .A(n15892), .B(n15891), .Z(n15896) );
  NANDN U16621 ( .A(n15894), .B(n15893), .Z(n15895) );
  AND U16622 ( .A(n15896), .B(n15895), .Z(n16043) );
  NANDN U16623 ( .A(n15898), .B(n15897), .Z(n15902) );
  NANDN U16624 ( .A(n15900), .B(n15899), .Z(n15901) );
  AND U16625 ( .A(n15902), .B(n15901), .Z(n16041) );
  NANDN U16626 ( .A(n15904), .B(n15903), .Z(n15908) );
  NANDN U16627 ( .A(n15906), .B(n15905), .Z(n15907) );
  AND U16628 ( .A(n15908), .B(n15907), .Z(n16130) );
  NAND U16629 ( .A(n38385), .B(n15909), .Z(n15911) );
  XOR U16630 ( .A(b[27]), .B(a[96]), .Z(n16076) );
  NAND U16631 ( .A(n38343), .B(n16076), .Z(n15910) );
  AND U16632 ( .A(n15911), .B(n15910), .Z(n16137) );
  NAND U16633 ( .A(n183), .B(n15912), .Z(n15914) );
  XOR U16634 ( .A(b[5]), .B(a[118]), .Z(n16079) );
  NAND U16635 ( .A(n36296), .B(n16079), .Z(n15913) );
  AND U16636 ( .A(n15914), .B(n15913), .Z(n16135) );
  NAND U16637 ( .A(n190), .B(n15915), .Z(n15917) );
  XOR U16638 ( .A(b[19]), .B(a[104]), .Z(n16082) );
  NAND U16639 ( .A(n37821), .B(n16082), .Z(n15916) );
  NAND U16640 ( .A(n15917), .B(n15916), .Z(n16134) );
  XNOR U16641 ( .A(n16135), .B(n16134), .Z(n16136) );
  XNOR U16642 ( .A(n16137), .B(n16136), .Z(n16128) );
  NAND U16643 ( .A(n38470), .B(n15918), .Z(n15920) );
  XOR U16644 ( .A(b[31]), .B(a[92]), .Z(n16085) );
  NAND U16645 ( .A(n38453), .B(n16085), .Z(n15919) );
  AND U16646 ( .A(n15920), .B(n15919), .Z(n16097) );
  NAND U16647 ( .A(n181), .B(n15921), .Z(n15923) );
  XOR U16648 ( .A(b[3]), .B(a[120]), .Z(n16088) );
  NAND U16649 ( .A(n182), .B(n16088), .Z(n15922) );
  AND U16650 ( .A(n15923), .B(n15922), .Z(n16095) );
  NAND U16651 ( .A(n189), .B(n15924), .Z(n15926) );
  XOR U16652 ( .A(b[17]), .B(a[106]), .Z(n16091) );
  NAND U16653 ( .A(n37652), .B(n16091), .Z(n15925) );
  NAND U16654 ( .A(n15926), .B(n15925), .Z(n16094) );
  XNOR U16655 ( .A(n16095), .B(n16094), .Z(n16096) );
  XOR U16656 ( .A(n16097), .B(n16096), .Z(n16129) );
  XOR U16657 ( .A(n16128), .B(n16129), .Z(n16131) );
  XOR U16658 ( .A(n16130), .B(n16131), .Z(n16065) );
  NANDN U16659 ( .A(n15928), .B(n15927), .Z(n15932) );
  NANDN U16660 ( .A(n15930), .B(n15929), .Z(n15931) );
  AND U16661 ( .A(n15932), .B(n15931), .Z(n16118) );
  NANDN U16662 ( .A(n15934), .B(n15933), .Z(n15938) );
  NANDN U16663 ( .A(n15936), .B(n15935), .Z(n15937) );
  NAND U16664 ( .A(n15938), .B(n15937), .Z(n16119) );
  XNOR U16665 ( .A(n16118), .B(n16119), .Z(n16120) );
  NANDN U16666 ( .A(n15940), .B(n15939), .Z(n15944) );
  NANDN U16667 ( .A(n15942), .B(n15941), .Z(n15943) );
  NAND U16668 ( .A(n15944), .B(n15943), .Z(n16121) );
  XNOR U16669 ( .A(n16120), .B(n16121), .Z(n16064) );
  XNOR U16670 ( .A(n16065), .B(n16064), .Z(n16067) );
  NANDN U16671 ( .A(n15946), .B(n15945), .Z(n15950) );
  NANDN U16672 ( .A(n15948), .B(n15947), .Z(n15949) );
  AND U16673 ( .A(n15950), .B(n15949), .Z(n16066) );
  XOR U16674 ( .A(n16067), .B(n16066), .Z(n16178) );
  NANDN U16675 ( .A(n15952), .B(n15951), .Z(n15956) );
  NANDN U16676 ( .A(n15954), .B(n15953), .Z(n15955) );
  AND U16677 ( .A(n15956), .B(n15955), .Z(n16176) );
  NANDN U16678 ( .A(n15958), .B(n15957), .Z(n15962) );
  NANDN U16679 ( .A(n15960), .B(n15959), .Z(n15961) );
  AND U16680 ( .A(n15962), .B(n15961), .Z(n16061) );
  NANDN U16681 ( .A(n15964), .B(n15963), .Z(n15968) );
  OR U16682 ( .A(n15966), .B(n15965), .Z(n15967) );
  AND U16683 ( .A(n15968), .B(n15967), .Z(n16059) );
  NANDN U16684 ( .A(n15970), .B(n15969), .Z(n15974) );
  NANDN U16685 ( .A(n15972), .B(n15971), .Z(n15973) );
  AND U16686 ( .A(n15974), .B(n15973), .Z(n16125) );
  NANDN U16687 ( .A(n15976), .B(n15975), .Z(n15980) );
  NANDN U16688 ( .A(n15978), .B(n15977), .Z(n15979) );
  NAND U16689 ( .A(n15980), .B(n15979), .Z(n16124) );
  XNOR U16690 ( .A(n16125), .B(n16124), .Z(n16127) );
  NAND U16691 ( .A(b[0]), .B(a[122]), .Z(n15981) );
  XNOR U16692 ( .A(b[1]), .B(n15981), .Z(n15983) );
  NANDN U16693 ( .A(b[0]), .B(a[121]), .Z(n15982) );
  NAND U16694 ( .A(n15983), .B(n15982), .Z(n16073) );
  NAND U16695 ( .A(n194), .B(n15984), .Z(n15986) );
  XOR U16696 ( .A(b[29]), .B(a[94]), .Z(n16149) );
  NAND U16697 ( .A(n38456), .B(n16149), .Z(n15985) );
  AND U16698 ( .A(n15986), .B(n15985), .Z(n16071) );
  AND U16699 ( .A(b[31]), .B(a[90]), .Z(n16070) );
  XNOR U16700 ( .A(n16071), .B(n16070), .Z(n16072) );
  XNOR U16701 ( .A(n16073), .B(n16072), .Z(n16113) );
  NAND U16702 ( .A(n38185), .B(n15987), .Z(n15989) );
  XOR U16703 ( .A(b[23]), .B(a[100]), .Z(n16152) );
  NAND U16704 ( .A(n38132), .B(n16152), .Z(n15988) );
  AND U16705 ( .A(n15989), .B(n15988), .Z(n16142) );
  NAND U16706 ( .A(n184), .B(n15990), .Z(n15992) );
  XOR U16707 ( .A(b[7]), .B(a[116]), .Z(n16155) );
  NAND U16708 ( .A(n36592), .B(n16155), .Z(n15991) );
  AND U16709 ( .A(n15992), .B(n15991), .Z(n16141) );
  NAND U16710 ( .A(n38289), .B(n15993), .Z(n15995) );
  XOR U16711 ( .A(b[25]), .B(a[98]), .Z(n16158) );
  NAND U16712 ( .A(n38247), .B(n16158), .Z(n15994) );
  NAND U16713 ( .A(n15995), .B(n15994), .Z(n16140) );
  XOR U16714 ( .A(n16141), .B(n16140), .Z(n16143) );
  XOR U16715 ( .A(n16142), .B(n16143), .Z(n16112) );
  XOR U16716 ( .A(n16113), .B(n16112), .Z(n16115) );
  NAND U16717 ( .A(n187), .B(n15996), .Z(n15998) );
  XOR U16718 ( .A(b[13]), .B(a[110]), .Z(n16161) );
  NAND U16719 ( .A(n37295), .B(n16161), .Z(n15997) );
  AND U16720 ( .A(n15998), .B(n15997), .Z(n16107) );
  NAND U16721 ( .A(n186), .B(n15999), .Z(n16001) );
  XOR U16722 ( .A(b[11]), .B(a[112]), .Z(n16164) );
  NAND U16723 ( .A(n37097), .B(n16164), .Z(n16000) );
  NAND U16724 ( .A(n16001), .B(n16000), .Z(n16106) );
  XNOR U16725 ( .A(n16107), .B(n16106), .Z(n16109) );
  NAND U16726 ( .A(n188), .B(n16002), .Z(n16004) );
  XOR U16727 ( .A(b[15]), .B(a[108]), .Z(n16167) );
  NAND U16728 ( .A(n37382), .B(n16167), .Z(n16003) );
  AND U16729 ( .A(n16004), .B(n16003), .Z(n16103) );
  NAND U16730 ( .A(n38064), .B(n16005), .Z(n16007) );
  XOR U16731 ( .A(b[21]), .B(a[102]), .Z(n16170) );
  NAND U16732 ( .A(n37993), .B(n16170), .Z(n16006) );
  AND U16733 ( .A(n16007), .B(n16006), .Z(n16101) );
  NAND U16734 ( .A(n185), .B(n16008), .Z(n16010) );
  XOR U16735 ( .A(b[9]), .B(a[114]), .Z(n16173) );
  NAND U16736 ( .A(n36805), .B(n16173), .Z(n16009) );
  NAND U16737 ( .A(n16010), .B(n16009), .Z(n16100) );
  XNOR U16738 ( .A(n16101), .B(n16100), .Z(n16102) );
  XNOR U16739 ( .A(n16103), .B(n16102), .Z(n16108) );
  XOR U16740 ( .A(n16109), .B(n16108), .Z(n16114) );
  XNOR U16741 ( .A(n16115), .B(n16114), .Z(n16126) );
  XNOR U16742 ( .A(n16127), .B(n16126), .Z(n16058) );
  XNOR U16743 ( .A(n16059), .B(n16058), .Z(n16060) );
  XOR U16744 ( .A(n16061), .B(n16060), .Z(n16177) );
  XOR U16745 ( .A(n16176), .B(n16177), .Z(n16179) );
  XOR U16746 ( .A(n16178), .B(n16179), .Z(n16055) );
  NANDN U16747 ( .A(n16012), .B(n16011), .Z(n16016) );
  NAND U16748 ( .A(n16014), .B(n16013), .Z(n16015) );
  AND U16749 ( .A(n16016), .B(n16015), .Z(n16053) );
  NANDN U16750 ( .A(n16018), .B(n16017), .Z(n16022) );
  NANDN U16751 ( .A(n16020), .B(n16019), .Z(n16021) );
  AND U16752 ( .A(n16022), .B(n16021), .Z(n16052) );
  XNOR U16753 ( .A(n16053), .B(n16052), .Z(n16054) );
  XNOR U16754 ( .A(n16055), .B(n16054), .Z(n16046) );
  NANDN U16755 ( .A(n16024), .B(n16023), .Z(n16028) );
  NANDN U16756 ( .A(n16026), .B(n16025), .Z(n16027) );
  NAND U16757 ( .A(n16028), .B(n16027), .Z(n16047) );
  XNOR U16758 ( .A(n16046), .B(n16047), .Z(n16048) );
  NANDN U16759 ( .A(n16030), .B(n16029), .Z(n16034) );
  NAND U16760 ( .A(n16032), .B(n16031), .Z(n16033) );
  NAND U16761 ( .A(n16034), .B(n16033), .Z(n16049) );
  XNOR U16762 ( .A(n16048), .B(n16049), .Z(n16040) );
  XNOR U16763 ( .A(n16041), .B(n16040), .Z(n16042) );
  XNOR U16764 ( .A(n16043), .B(n16042), .Z(n16182) );
  XNOR U16765 ( .A(sreg[346]), .B(n16182), .Z(n16184) );
  NANDN U16766 ( .A(sreg[345]), .B(n16035), .Z(n16039) );
  NAND U16767 ( .A(n16037), .B(n16036), .Z(n16038) );
  NAND U16768 ( .A(n16039), .B(n16038), .Z(n16183) );
  XNOR U16769 ( .A(n16184), .B(n16183), .Z(c[346]) );
  NANDN U16770 ( .A(n16041), .B(n16040), .Z(n16045) );
  NANDN U16771 ( .A(n16043), .B(n16042), .Z(n16044) );
  AND U16772 ( .A(n16045), .B(n16044), .Z(n16190) );
  NANDN U16773 ( .A(n16047), .B(n16046), .Z(n16051) );
  NANDN U16774 ( .A(n16049), .B(n16048), .Z(n16050) );
  AND U16775 ( .A(n16051), .B(n16050), .Z(n16188) );
  NANDN U16776 ( .A(n16053), .B(n16052), .Z(n16057) );
  NANDN U16777 ( .A(n16055), .B(n16054), .Z(n16056) );
  AND U16778 ( .A(n16057), .B(n16056), .Z(n16196) );
  NANDN U16779 ( .A(n16059), .B(n16058), .Z(n16063) );
  NANDN U16780 ( .A(n16061), .B(n16060), .Z(n16062) );
  AND U16781 ( .A(n16063), .B(n16062), .Z(n16326) );
  NANDN U16782 ( .A(n16065), .B(n16064), .Z(n16069) );
  NAND U16783 ( .A(n16067), .B(n16066), .Z(n16068) );
  AND U16784 ( .A(n16069), .B(n16068), .Z(n16325) );
  XNOR U16785 ( .A(n16326), .B(n16325), .Z(n16328) );
  NANDN U16786 ( .A(n16071), .B(n16070), .Z(n16075) );
  NANDN U16787 ( .A(n16073), .B(n16072), .Z(n16074) );
  AND U16788 ( .A(n16075), .B(n16074), .Z(n16261) );
  NAND U16789 ( .A(n38385), .B(n16076), .Z(n16078) );
  XOR U16790 ( .A(b[27]), .B(a[97]), .Z(n16205) );
  NAND U16791 ( .A(n38343), .B(n16205), .Z(n16077) );
  AND U16792 ( .A(n16078), .B(n16077), .Z(n16268) );
  NAND U16793 ( .A(n183), .B(n16079), .Z(n16081) );
  XOR U16794 ( .A(b[5]), .B(a[119]), .Z(n16208) );
  NAND U16795 ( .A(n36296), .B(n16208), .Z(n16080) );
  AND U16796 ( .A(n16081), .B(n16080), .Z(n16266) );
  NAND U16797 ( .A(n190), .B(n16082), .Z(n16084) );
  XOR U16798 ( .A(b[19]), .B(a[105]), .Z(n16211) );
  NAND U16799 ( .A(n37821), .B(n16211), .Z(n16083) );
  NAND U16800 ( .A(n16084), .B(n16083), .Z(n16265) );
  XNOR U16801 ( .A(n16266), .B(n16265), .Z(n16267) );
  XNOR U16802 ( .A(n16268), .B(n16267), .Z(n16259) );
  NAND U16803 ( .A(n38470), .B(n16085), .Z(n16087) );
  XOR U16804 ( .A(b[31]), .B(a[93]), .Z(n16214) );
  NAND U16805 ( .A(n38453), .B(n16214), .Z(n16086) );
  AND U16806 ( .A(n16087), .B(n16086), .Z(n16226) );
  NAND U16807 ( .A(n181), .B(n16088), .Z(n16090) );
  XOR U16808 ( .A(b[3]), .B(a[121]), .Z(n16217) );
  NAND U16809 ( .A(n182), .B(n16217), .Z(n16089) );
  AND U16810 ( .A(n16090), .B(n16089), .Z(n16224) );
  NAND U16811 ( .A(n189), .B(n16091), .Z(n16093) );
  XOR U16812 ( .A(b[17]), .B(a[107]), .Z(n16220) );
  NAND U16813 ( .A(n37652), .B(n16220), .Z(n16092) );
  NAND U16814 ( .A(n16093), .B(n16092), .Z(n16223) );
  XNOR U16815 ( .A(n16224), .B(n16223), .Z(n16225) );
  XOR U16816 ( .A(n16226), .B(n16225), .Z(n16260) );
  XOR U16817 ( .A(n16259), .B(n16260), .Z(n16262) );
  XOR U16818 ( .A(n16261), .B(n16262), .Z(n16308) );
  NANDN U16819 ( .A(n16095), .B(n16094), .Z(n16099) );
  NANDN U16820 ( .A(n16097), .B(n16096), .Z(n16098) );
  AND U16821 ( .A(n16099), .B(n16098), .Z(n16247) );
  NANDN U16822 ( .A(n16101), .B(n16100), .Z(n16105) );
  NANDN U16823 ( .A(n16103), .B(n16102), .Z(n16104) );
  NAND U16824 ( .A(n16105), .B(n16104), .Z(n16248) );
  XNOR U16825 ( .A(n16247), .B(n16248), .Z(n16249) );
  NANDN U16826 ( .A(n16107), .B(n16106), .Z(n16111) );
  NAND U16827 ( .A(n16109), .B(n16108), .Z(n16110) );
  NAND U16828 ( .A(n16111), .B(n16110), .Z(n16250) );
  XNOR U16829 ( .A(n16249), .B(n16250), .Z(n16307) );
  XNOR U16830 ( .A(n16308), .B(n16307), .Z(n16310) );
  NAND U16831 ( .A(n16113), .B(n16112), .Z(n16117) );
  NAND U16832 ( .A(n16115), .B(n16114), .Z(n16116) );
  AND U16833 ( .A(n16117), .B(n16116), .Z(n16309) );
  XOR U16834 ( .A(n16310), .B(n16309), .Z(n16322) );
  NANDN U16835 ( .A(n16119), .B(n16118), .Z(n16123) );
  NANDN U16836 ( .A(n16121), .B(n16120), .Z(n16122) );
  AND U16837 ( .A(n16123), .B(n16122), .Z(n16319) );
  NANDN U16838 ( .A(n16129), .B(n16128), .Z(n16133) );
  OR U16839 ( .A(n16131), .B(n16130), .Z(n16132) );
  AND U16840 ( .A(n16133), .B(n16132), .Z(n16314) );
  NANDN U16841 ( .A(n16135), .B(n16134), .Z(n16139) );
  NANDN U16842 ( .A(n16137), .B(n16136), .Z(n16138) );
  AND U16843 ( .A(n16139), .B(n16138), .Z(n16254) );
  NANDN U16844 ( .A(n16141), .B(n16140), .Z(n16145) );
  OR U16845 ( .A(n16143), .B(n16142), .Z(n16144) );
  NAND U16846 ( .A(n16145), .B(n16144), .Z(n16253) );
  XNOR U16847 ( .A(n16254), .B(n16253), .Z(n16255) );
  NAND U16848 ( .A(b[0]), .B(a[123]), .Z(n16146) );
  XNOR U16849 ( .A(b[1]), .B(n16146), .Z(n16148) );
  NANDN U16850 ( .A(b[0]), .B(a[122]), .Z(n16147) );
  NAND U16851 ( .A(n16148), .B(n16147), .Z(n16202) );
  NAND U16852 ( .A(n194), .B(n16149), .Z(n16151) );
  XOR U16853 ( .A(b[29]), .B(a[95]), .Z(n16280) );
  NAND U16854 ( .A(n38456), .B(n16280), .Z(n16150) );
  AND U16855 ( .A(n16151), .B(n16150), .Z(n16200) );
  AND U16856 ( .A(b[31]), .B(a[91]), .Z(n16199) );
  XNOR U16857 ( .A(n16200), .B(n16199), .Z(n16201) );
  XNOR U16858 ( .A(n16202), .B(n16201), .Z(n16241) );
  NAND U16859 ( .A(n38185), .B(n16152), .Z(n16154) );
  XOR U16860 ( .A(b[23]), .B(a[101]), .Z(n16283) );
  NAND U16861 ( .A(n38132), .B(n16283), .Z(n16153) );
  AND U16862 ( .A(n16154), .B(n16153), .Z(n16274) );
  NAND U16863 ( .A(n184), .B(n16155), .Z(n16157) );
  XOR U16864 ( .A(b[7]), .B(a[117]), .Z(n16286) );
  NAND U16865 ( .A(n36592), .B(n16286), .Z(n16156) );
  AND U16866 ( .A(n16157), .B(n16156), .Z(n16272) );
  NAND U16867 ( .A(n38289), .B(n16158), .Z(n16160) );
  XOR U16868 ( .A(b[25]), .B(a[99]), .Z(n16289) );
  NAND U16869 ( .A(n38247), .B(n16289), .Z(n16159) );
  NAND U16870 ( .A(n16160), .B(n16159), .Z(n16271) );
  XNOR U16871 ( .A(n16272), .B(n16271), .Z(n16273) );
  XOR U16872 ( .A(n16274), .B(n16273), .Z(n16242) );
  XNOR U16873 ( .A(n16241), .B(n16242), .Z(n16243) );
  NAND U16874 ( .A(n187), .B(n16161), .Z(n16163) );
  XOR U16875 ( .A(b[13]), .B(a[111]), .Z(n16292) );
  NAND U16876 ( .A(n37295), .B(n16292), .Z(n16162) );
  AND U16877 ( .A(n16163), .B(n16162), .Z(n16236) );
  NAND U16878 ( .A(n186), .B(n16164), .Z(n16166) );
  XOR U16879 ( .A(b[11]), .B(a[113]), .Z(n16295) );
  NAND U16880 ( .A(n37097), .B(n16295), .Z(n16165) );
  NAND U16881 ( .A(n16166), .B(n16165), .Z(n16235) );
  XNOR U16882 ( .A(n16236), .B(n16235), .Z(n16237) );
  NAND U16883 ( .A(n188), .B(n16167), .Z(n16169) );
  XOR U16884 ( .A(b[15]), .B(a[109]), .Z(n16298) );
  NAND U16885 ( .A(n37382), .B(n16298), .Z(n16168) );
  AND U16886 ( .A(n16169), .B(n16168), .Z(n16232) );
  NAND U16887 ( .A(n38064), .B(n16170), .Z(n16172) );
  XOR U16888 ( .A(b[21]), .B(a[103]), .Z(n16301) );
  NAND U16889 ( .A(n37993), .B(n16301), .Z(n16171) );
  AND U16890 ( .A(n16172), .B(n16171), .Z(n16230) );
  NAND U16891 ( .A(n185), .B(n16173), .Z(n16175) );
  XOR U16892 ( .A(b[9]), .B(a[115]), .Z(n16304) );
  NAND U16893 ( .A(n36805), .B(n16304), .Z(n16174) );
  NAND U16894 ( .A(n16175), .B(n16174), .Z(n16229) );
  XNOR U16895 ( .A(n16230), .B(n16229), .Z(n16231) );
  XOR U16896 ( .A(n16232), .B(n16231), .Z(n16238) );
  XOR U16897 ( .A(n16237), .B(n16238), .Z(n16244) );
  XOR U16898 ( .A(n16243), .B(n16244), .Z(n16256) );
  XNOR U16899 ( .A(n16255), .B(n16256), .Z(n16313) );
  XNOR U16900 ( .A(n16314), .B(n16313), .Z(n16315) );
  XOR U16901 ( .A(n16316), .B(n16315), .Z(n16320) );
  XNOR U16902 ( .A(n16319), .B(n16320), .Z(n16321) );
  XNOR U16903 ( .A(n16322), .B(n16321), .Z(n16327) );
  XOR U16904 ( .A(n16328), .B(n16327), .Z(n16194) );
  NANDN U16905 ( .A(n16177), .B(n16176), .Z(n16181) );
  OR U16906 ( .A(n16179), .B(n16178), .Z(n16180) );
  AND U16907 ( .A(n16181), .B(n16180), .Z(n16193) );
  XNOR U16908 ( .A(n16194), .B(n16193), .Z(n16195) );
  XNOR U16909 ( .A(n16196), .B(n16195), .Z(n16187) );
  XNOR U16910 ( .A(n16188), .B(n16187), .Z(n16189) );
  XNOR U16911 ( .A(n16190), .B(n16189), .Z(n16331) );
  XNOR U16912 ( .A(sreg[347]), .B(n16331), .Z(n16333) );
  NANDN U16913 ( .A(sreg[346]), .B(n16182), .Z(n16186) );
  NAND U16914 ( .A(n16184), .B(n16183), .Z(n16185) );
  NAND U16915 ( .A(n16186), .B(n16185), .Z(n16332) );
  XNOR U16916 ( .A(n16333), .B(n16332), .Z(c[347]) );
  NANDN U16917 ( .A(n16188), .B(n16187), .Z(n16192) );
  NANDN U16918 ( .A(n16190), .B(n16189), .Z(n16191) );
  AND U16919 ( .A(n16192), .B(n16191), .Z(n16339) );
  NANDN U16920 ( .A(n16194), .B(n16193), .Z(n16198) );
  NANDN U16921 ( .A(n16196), .B(n16195), .Z(n16197) );
  AND U16922 ( .A(n16198), .B(n16197), .Z(n16337) );
  NANDN U16923 ( .A(n16200), .B(n16199), .Z(n16204) );
  NANDN U16924 ( .A(n16202), .B(n16201), .Z(n16203) );
  AND U16925 ( .A(n16204), .B(n16203), .Z(n16428) );
  NAND U16926 ( .A(n38385), .B(n16205), .Z(n16207) );
  XOR U16927 ( .A(b[27]), .B(a[98]), .Z(n16372) );
  NAND U16928 ( .A(n38343), .B(n16372), .Z(n16206) );
  AND U16929 ( .A(n16207), .B(n16206), .Z(n16435) );
  NAND U16930 ( .A(n183), .B(n16208), .Z(n16210) );
  XOR U16931 ( .A(b[5]), .B(a[120]), .Z(n16375) );
  NAND U16932 ( .A(n36296), .B(n16375), .Z(n16209) );
  AND U16933 ( .A(n16210), .B(n16209), .Z(n16433) );
  NAND U16934 ( .A(n190), .B(n16211), .Z(n16213) );
  XOR U16935 ( .A(b[19]), .B(a[106]), .Z(n16378) );
  NAND U16936 ( .A(n37821), .B(n16378), .Z(n16212) );
  NAND U16937 ( .A(n16213), .B(n16212), .Z(n16432) );
  XNOR U16938 ( .A(n16433), .B(n16432), .Z(n16434) );
  XNOR U16939 ( .A(n16435), .B(n16434), .Z(n16426) );
  NAND U16940 ( .A(n38470), .B(n16214), .Z(n16216) );
  XOR U16941 ( .A(b[31]), .B(a[94]), .Z(n16381) );
  NAND U16942 ( .A(n38453), .B(n16381), .Z(n16215) );
  AND U16943 ( .A(n16216), .B(n16215), .Z(n16393) );
  NAND U16944 ( .A(n181), .B(n16217), .Z(n16219) );
  XOR U16945 ( .A(b[3]), .B(a[122]), .Z(n16384) );
  NAND U16946 ( .A(n182), .B(n16384), .Z(n16218) );
  AND U16947 ( .A(n16219), .B(n16218), .Z(n16391) );
  NAND U16948 ( .A(n189), .B(n16220), .Z(n16222) );
  XOR U16949 ( .A(b[17]), .B(a[108]), .Z(n16387) );
  NAND U16950 ( .A(n37652), .B(n16387), .Z(n16221) );
  NAND U16951 ( .A(n16222), .B(n16221), .Z(n16390) );
  XNOR U16952 ( .A(n16391), .B(n16390), .Z(n16392) );
  XOR U16953 ( .A(n16393), .B(n16392), .Z(n16427) );
  XOR U16954 ( .A(n16426), .B(n16427), .Z(n16429) );
  XOR U16955 ( .A(n16428), .B(n16429), .Z(n16361) );
  NANDN U16956 ( .A(n16224), .B(n16223), .Z(n16228) );
  NANDN U16957 ( .A(n16226), .B(n16225), .Z(n16227) );
  AND U16958 ( .A(n16228), .B(n16227), .Z(n16414) );
  NANDN U16959 ( .A(n16230), .B(n16229), .Z(n16234) );
  NANDN U16960 ( .A(n16232), .B(n16231), .Z(n16233) );
  NAND U16961 ( .A(n16234), .B(n16233), .Z(n16415) );
  XNOR U16962 ( .A(n16414), .B(n16415), .Z(n16416) );
  NANDN U16963 ( .A(n16236), .B(n16235), .Z(n16240) );
  NANDN U16964 ( .A(n16238), .B(n16237), .Z(n16239) );
  NAND U16965 ( .A(n16240), .B(n16239), .Z(n16417) );
  XNOR U16966 ( .A(n16416), .B(n16417), .Z(n16360) );
  XNOR U16967 ( .A(n16361), .B(n16360), .Z(n16363) );
  NANDN U16968 ( .A(n16242), .B(n16241), .Z(n16246) );
  NANDN U16969 ( .A(n16244), .B(n16243), .Z(n16245) );
  AND U16970 ( .A(n16246), .B(n16245), .Z(n16362) );
  XOR U16971 ( .A(n16363), .B(n16362), .Z(n16476) );
  NANDN U16972 ( .A(n16248), .B(n16247), .Z(n16252) );
  NANDN U16973 ( .A(n16250), .B(n16249), .Z(n16251) );
  AND U16974 ( .A(n16252), .B(n16251), .Z(n16474) );
  NANDN U16975 ( .A(n16254), .B(n16253), .Z(n16258) );
  NANDN U16976 ( .A(n16256), .B(n16255), .Z(n16257) );
  AND U16977 ( .A(n16258), .B(n16257), .Z(n16357) );
  NANDN U16978 ( .A(n16260), .B(n16259), .Z(n16264) );
  OR U16979 ( .A(n16262), .B(n16261), .Z(n16263) );
  AND U16980 ( .A(n16264), .B(n16263), .Z(n16355) );
  NANDN U16981 ( .A(n16266), .B(n16265), .Z(n16270) );
  NANDN U16982 ( .A(n16268), .B(n16267), .Z(n16269) );
  AND U16983 ( .A(n16270), .B(n16269), .Z(n16421) );
  NANDN U16984 ( .A(n16272), .B(n16271), .Z(n16276) );
  NANDN U16985 ( .A(n16274), .B(n16273), .Z(n16275) );
  NAND U16986 ( .A(n16276), .B(n16275), .Z(n16420) );
  XNOR U16987 ( .A(n16421), .B(n16420), .Z(n16422) );
  NAND U16988 ( .A(b[0]), .B(a[124]), .Z(n16277) );
  XNOR U16989 ( .A(b[1]), .B(n16277), .Z(n16279) );
  NANDN U16990 ( .A(b[0]), .B(a[123]), .Z(n16278) );
  NAND U16991 ( .A(n16279), .B(n16278), .Z(n16369) );
  NAND U16992 ( .A(n194), .B(n16280), .Z(n16282) );
  XOR U16993 ( .A(b[29]), .B(a[96]), .Z(n16444) );
  NAND U16994 ( .A(n38456), .B(n16444), .Z(n16281) );
  AND U16995 ( .A(n16282), .B(n16281), .Z(n16367) );
  AND U16996 ( .A(b[31]), .B(a[92]), .Z(n16366) );
  XNOR U16997 ( .A(n16367), .B(n16366), .Z(n16368) );
  XNOR U16998 ( .A(n16369), .B(n16368), .Z(n16408) );
  NAND U16999 ( .A(n38185), .B(n16283), .Z(n16285) );
  XOR U17000 ( .A(b[23]), .B(a[102]), .Z(n16450) );
  NAND U17001 ( .A(n38132), .B(n16450), .Z(n16284) );
  AND U17002 ( .A(n16285), .B(n16284), .Z(n16441) );
  NAND U17003 ( .A(n184), .B(n16286), .Z(n16288) );
  XOR U17004 ( .A(b[7]), .B(a[118]), .Z(n16453) );
  NAND U17005 ( .A(n36592), .B(n16453), .Z(n16287) );
  AND U17006 ( .A(n16288), .B(n16287), .Z(n16439) );
  NAND U17007 ( .A(n38289), .B(n16289), .Z(n16291) );
  XOR U17008 ( .A(b[25]), .B(a[100]), .Z(n16456) );
  NAND U17009 ( .A(n38247), .B(n16456), .Z(n16290) );
  NAND U17010 ( .A(n16291), .B(n16290), .Z(n16438) );
  XNOR U17011 ( .A(n16439), .B(n16438), .Z(n16440) );
  XOR U17012 ( .A(n16441), .B(n16440), .Z(n16409) );
  XNOR U17013 ( .A(n16408), .B(n16409), .Z(n16410) );
  NAND U17014 ( .A(n187), .B(n16292), .Z(n16294) );
  XOR U17015 ( .A(b[13]), .B(a[112]), .Z(n16459) );
  NAND U17016 ( .A(n37295), .B(n16459), .Z(n16293) );
  AND U17017 ( .A(n16294), .B(n16293), .Z(n16403) );
  NAND U17018 ( .A(n186), .B(n16295), .Z(n16297) );
  XOR U17019 ( .A(b[11]), .B(a[114]), .Z(n16462) );
  NAND U17020 ( .A(n37097), .B(n16462), .Z(n16296) );
  NAND U17021 ( .A(n16297), .B(n16296), .Z(n16402) );
  XNOR U17022 ( .A(n16403), .B(n16402), .Z(n16404) );
  NAND U17023 ( .A(n188), .B(n16298), .Z(n16300) );
  XOR U17024 ( .A(b[15]), .B(a[110]), .Z(n16465) );
  NAND U17025 ( .A(n37382), .B(n16465), .Z(n16299) );
  AND U17026 ( .A(n16300), .B(n16299), .Z(n16399) );
  NAND U17027 ( .A(n38064), .B(n16301), .Z(n16303) );
  XOR U17028 ( .A(b[21]), .B(a[104]), .Z(n16468) );
  NAND U17029 ( .A(n37993), .B(n16468), .Z(n16302) );
  AND U17030 ( .A(n16303), .B(n16302), .Z(n16397) );
  NAND U17031 ( .A(n185), .B(n16304), .Z(n16306) );
  XOR U17032 ( .A(b[9]), .B(a[116]), .Z(n16471) );
  NAND U17033 ( .A(n36805), .B(n16471), .Z(n16305) );
  NAND U17034 ( .A(n16306), .B(n16305), .Z(n16396) );
  XNOR U17035 ( .A(n16397), .B(n16396), .Z(n16398) );
  XOR U17036 ( .A(n16399), .B(n16398), .Z(n16405) );
  XOR U17037 ( .A(n16404), .B(n16405), .Z(n16411) );
  XOR U17038 ( .A(n16410), .B(n16411), .Z(n16423) );
  XNOR U17039 ( .A(n16422), .B(n16423), .Z(n16354) );
  XNOR U17040 ( .A(n16355), .B(n16354), .Z(n16356) );
  XOR U17041 ( .A(n16357), .B(n16356), .Z(n16475) );
  XOR U17042 ( .A(n16474), .B(n16475), .Z(n16477) );
  XOR U17043 ( .A(n16476), .B(n16477), .Z(n16351) );
  NANDN U17044 ( .A(n16308), .B(n16307), .Z(n16312) );
  NAND U17045 ( .A(n16310), .B(n16309), .Z(n16311) );
  AND U17046 ( .A(n16312), .B(n16311), .Z(n16349) );
  NANDN U17047 ( .A(n16314), .B(n16313), .Z(n16318) );
  NANDN U17048 ( .A(n16316), .B(n16315), .Z(n16317) );
  AND U17049 ( .A(n16318), .B(n16317), .Z(n16348) );
  XNOR U17050 ( .A(n16349), .B(n16348), .Z(n16350) );
  XNOR U17051 ( .A(n16351), .B(n16350), .Z(n16342) );
  NANDN U17052 ( .A(n16320), .B(n16319), .Z(n16324) );
  NANDN U17053 ( .A(n16322), .B(n16321), .Z(n16323) );
  NAND U17054 ( .A(n16324), .B(n16323), .Z(n16343) );
  XNOR U17055 ( .A(n16342), .B(n16343), .Z(n16344) );
  NANDN U17056 ( .A(n16326), .B(n16325), .Z(n16330) );
  NAND U17057 ( .A(n16328), .B(n16327), .Z(n16329) );
  NAND U17058 ( .A(n16330), .B(n16329), .Z(n16345) );
  XNOR U17059 ( .A(n16344), .B(n16345), .Z(n16336) );
  XNOR U17060 ( .A(n16337), .B(n16336), .Z(n16338) );
  XNOR U17061 ( .A(n16339), .B(n16338), .Z(n16480) );
  XNOR U17062 ( .A(sreg[348]), .B(n16480), .Z(n16482) );
  NANDN U17063 ( .A(sreg[347]), .B(n16331), .Z(n16335) );
  NAND U17064 ( .A(n16333), .B(n16332), .Z(n16334) );
  NAND U17065 ( .A(n16335), .B(n16334), .Z(n16481) );
  XNOR U17066 ( .A(n16482), .B(n16481), .Z(c[348]) );
  NANDN U17067 ( .A(n16337), .B(n16336), .Z(n16341) );
  NANDN U17068 ( .A(n16339), .B(n16338), .Z(n16340) );
  AND U17069 ( .A(n16341), .B(n16340), .Z(n16488) );
  NANDN U17070 ( .A(n16343), .B(n16342), .Z(n16347) );
  NANDN U17071 ( .A(n16345), .B(n16344), .Z(n16346) );
  AND U17072 ( .A(n16347), .B(n16346), .Z(n16486) );
  NANDN U17073 ( .A(n16349), .B(n16348), .Z(n16353) );
  NANDN U17074 ( .A(n16351), .B(n16350), .Z(n16352) );
  AND U17075 ( .A(n16353), .B(n16352), .Z(n16494) );
  NANDN U17076 ( .A(n16355), .B(n16354), .Z(n16359) );
  NANDN U17077 ( .A(n16357), .B(n16356), .Z(n16358) );
  AND U17078 ( .A(n16359), .B(n16358), .Z(n16498) );
  NANDN U17079 ( .A(n16361), .B(n16360), .Z(n16365) );
  NAND U17080 ( .A(n16363), .B(n16362), .Z(n16364) );
  AND U17081 ( .A(n16365), .B(n16364), .Z(n16497) );
  XNOR U17082 ( .A(n16498), .B(n16497), .Z(n16500) );
  NANDN U17083 ( .A(n16367), .B(n16366), .Z(n16371) );
  NANDN U17084 ( .A(n16369), .B(n16368), .Z(n16370) );
  AND U17085 ( .A(n16371), .B(n16370), .Z(n16577) );
  NAND U17086 ( .A(n38385), .B(n16372), .Z(n16374) );
  XOR U17087 ( .A(b[27]), .B(a[99]), .Z(n16521) );
  NAND U17088 ( .A(n38343), .B(n16521), .Z(n16373) );
  AND U17089 ( .A(n16374), .B(n16373), .Z(n16584) );
  NAND U17090 ( .A(n183), .B(n16375), .Z(n16377) );
  XOR U17091 ( .A(b[5]), .B(a[121]), .Z(n16524) );
  NAND U17092 ( .A(n36296), .B(n16524), .Z(n16376) );
  AND U17093 ( .A(n16377), .B(n16376), .Z(n16582) );
  NAND U17094 ( .A(n190), .B(n16378), .Z(n16380) );
  XOR U17095 ( .A(b[19]), .B(a[107]), .Z(n16527) );
  NAND U17096 ( .A(n37821), .B(n16527), .Z(n16379) );
  NAND U17097 ( .A(n16380), .B(n16379), .Z(n16581) );
  XNOR U17098 ( .A(n16582), .B(n16581), .Z(n16583) );
  XNOR U17099 ( .A(n16584), .B(n16583), .Z(n16575) );
  NAND U17100 ( .A(n38470), .B(n16381), .Z(n16383) );
  XOR U17101 ( .A(b[31]), .B(a[95]), .Z(n16530) );
  NAND U17102 ( .A(n38453), .B(n16530), .Z(n16382) );
  AND U17103 ( .A(n16383), .B(n16382), .Z(n16542) );
  NAND U17104 ( .A(n181), .B(n16384), .Z(n16386) );
  XOR U17105 ( .A(b[3]), .B(a[123]), .Z(n16533) );
  NAND U17106 ( .A(n182), .B(n16533), .Z(n16385) );
  AND U17107 ( .A(n16386), .B(n16385), .Z(n16540) );
  NAND U17108 ( .A(n189), .B(n16387), .Z(n16389) );
  XOR U17109 ( .A(b[17]), .B(a[109]), .Z(n16536) );
  NAND U17110 ( .A(n37652), .B(n16536), .Z(n16388) );
  NAND U17111 ( .A(n16389), .B(n16388), .Z(n16539) );
  XNOR U17112 ( .A(n16540), .B(n16539), .Z(n16541) );
  XOR U17113 ( .A(n16542), .B(n16541), .Z(n16576) );
  XOR U17114 ( .A(n16575), .B(n16576), .Z(n16578) );
  XOR U17115 ( .A(n16577), .B(n16578), .Z(n16510) );
  NANDN U17116 ( .A(n16391), .B(n16390), .Z(n16395) );
  NANDN U17117 ( .A(n16393), .B(n16392), .Z(n16394) );
  AND U17118 ( .A(n16395), .B(n16394), .Z(n16563) );
  NANDN U17119 ( .A(n16397), .B(n16396), .Z(n16401) );
  NANDN U17120 ( .A(n16399), .B(n16398), .Z(n16400) );
  NAND U17121 ( .A(n16401), .B(n16400), .Z(n16564) );
  XNOR U17122 ( .A(n16563), .B(n16564), .Z(n16565) );
  NANDN U17123 ( .A(n16403), .B(n16402), .Z(n16407) );
  NANDN U17124 ( .A(n16405), .B(n16404), .Z(n16406) );
  NAND U17125 ( .A(n16407), .B(n16406), .Z(n16566) );
  XNOR U17126 ( .A(n16565), .B(n16566), .Z(n16509) );
  XNOR U17127 ( .A(n16510), .B(n16509), .Z(n16512) );
  NANDN U17128 ( .A(n16409), .B(n16408), .Z(n16413) );
  NANDN U17129 ( .A(n16411), .B(n16410), .Z(n16412) );
  AND U17130 ( .A(n16413), .B(n16412), .Z(n16511) );
  XOR U17131 ( .A(n16512), .B(n16511), .Z(n16626) );
  NANDN U17132 ( .A(n16415), .B(n16414), .Z(n16419) );
  NANDN U17133 ( .A(n16417), .B(n16416), .Z(n16418) );
  AND U17134 ( .A(n16419), .B(n16418), .Z(n16623) );
  NANDN U17135 ( .A(n16421), .B(n16420), .Z(n16425) );
  NANDN U17136 ( .A(n16423), .B(n16422), .Z(n16424) );
  AND U17137 ( .A(n16425), .B(n16424), .Z(n16506) );
  NANDN U17138 ( .A(n16427), .B(n16426), .Z(n16431) );
  OR U17139 ( .A(n16429), .B(n16428), .Z(n16430) );
  AND U17140 ( .A(n16431), .B(n16430), .Z(n16504) );
  NANDN U17141 ( .A(n16433), .B(n16432), .Z(n16437) );
  NANDN U17142 ( .A(n16435), .B(n16434), .Z(n16436) );
  AND U17143 ( .A(n16437), .B(n16436), .Z(n16570) );
  NANDN U17144 ( .A(n16439), .B(n16438), .Z(n16443) );
  NANDN U17145 ( .A(n16441), .B(n16440), .Z(n16442) );
  NAND U17146 ( .A(n16443), .B(n16442), .Z(n16569) );
  XNOR U17147 ( .A(n16570), .B(n16569), .Z(n16571) );
  NAND U17148 ( .A(n194), .B(n16444), .Z(n16446) );
  XOR U17149 ( .A(b[29]), .B(a[97]), .Z(n16596) );
  NAND U17150 ( .A(n38456), .B(n16596), .Z(n16445) );
  AND U17151 ( .A(n16446), .B(n16445), .Z(n16516) );
  AND U17152 ( .A(b[31]), .B(a[93]), .Z(n16515) );
  XNOR U17153 ( .A(n16516), .B(n16515), .Z(n16517) );
  NAND U17154 ( .A(b[0]), .B(a[125]), .Z(n16447) );
  XNOR U17155 ( .A(b[1]), .B(n16447), .Z(n16449) );
  NANDN U17156 ( .A(b[0]), .B(a[124]), .Z(n16448) );
  NAND U17157 ( .A(n16449), .B(n16448), .Z(n16518) );
  XNOR U17158 ( .A(n16517), .B(n16518), .Z(n16557) );
  NAND U17159 ( .A(n38185), .B(n16450), .Z(n16452) );
  XOR U17160 ( .A(b[23]), .B(a[103]), .Z(n16599) );
  NAND U17161 ( .A(n38132), .B(n16599), .Z(n16451) );
  AND U17162 ( .A(n16452), .B(n16451), .Z(n16590) );
  NAND U17163 ( .A(n184), .B(n16453), .Z(n16455) );
  XOR U17164 ( .A(b[7]), .B(a[119]), .Z(n16602) );
  NAND U17165 ( .A(n36592), .B(n16602), .Z(n16454) );
  AND U17166 ( .A(n16455), .B(n16454), .Z(n16588) );
  NAND U17167 ( .A(n38289), .B(n16456), .Z(n16458) );
  XOR U17168 ( .A(b[25]), .B(a[101]), .Z(n16605) );
  NAND U17169 ( .A(n38247), .B(n16605), .Z(n16457) );
  NAND U17170 ( .A(n16458), .B(n16457), .Z(n16587) );
  XNOR U17171 ( .A(n16588), .B(n16587), .Z(n16589) );
  XOR U17172 ( .A(n16590), .B(n16589), .Z(n16558) );
  XNOR U17173 ( .A(n16557), .B(n16558), .Z(n16559) );
  NAND U17174 ( .A(n187), .B(n16459), .Z(n16461) );
  XOR U17175 ( .A(b[13]), .B(a[113]), .Z(n16608) );
  NAND U17176 ( .A(n37295), .B(n16608), .Z(n16460) );
  AND U17177 ( .A(n16461), .B(n16460), .Z(n16552) );
  NAND U17178 ( .A(n186), .B(n16462), .Z(n16464) );
  XOR U17179 ( .A(b[11]), .B(a[115]), .Z(n16611) );
  NAND U17180 ( .A(n37097), .B(n16611), .Z(n16463) );
  NAND U17181 ( .A(n16464), .B(n16463), .Z(n16551) );
  XNOR U17182 ( .A(n16552), .B(n16551), .Z(n16553) );
  NAND U17183 ( .A(n188), .B(n16465), .Z(n16467) );
  XOR U17184 ( .A(b[15]), .B(a[111]), .Z(n16614) );
  NAND U17185 ( .A(n37382), .B(n16614), .Z(n16466) );
  AND U17186 ( .A(n16467), .B(n16466), .Z(n16548) );
  NAND U17187 ( .A(n38064), .B(n16468), .Z(n16470) );
  XOR U17188 ( .A(b[21]), .B(a[105]), .Z(n16617) );
  NAND U17189 ( .A(n37993), .B(n16617), .Z(n16469) );
  AND U17190 ( .A(n16470), .B(n16469), .Z(n16546) );
  NAND U17191 ( .A(n185), .B(n16471), .Z(n16473) );
  XOR U17192 ( .A(b[9]), .B(a[117]), .Z(n16620) );
  NAND U17193 ( .A(n36805), .B(n16620), .Z(n16472) );
  NAND U17194 ( .A(n16473), .B(n16472), .Z(n16545) );
  XNOR U17195 ( .A(n16546), .B(n16545), .Z(n16547) );
  XOR U17196 ( .A(n16548), .B(n16547), .Z(n16554) );
  XOR U17197 ( .A(n16553), .B(n16554), .Z(n16560) );
  XOR U17198 ( .A(n16559), .B(n16560), .Z(n16572) );
  XNOR U17199 ( .A(n16571), .B(n16572), .Z(n16503) );
  XNOR U17200 ( .A(n16504), .B(n16503), .Z(n16505) );
  XOR U17201 ( .A(n16506), .B(n16505), .Z(n16624) );
  XNOR U17202 ( .A(n16623), .B(n16624), .Z(n16625) );
  XNOR U17203 ( .A(n16626), .B(n16625), .Z(n16499) );
  XOR U17204 ( .A(n16500), .B(n16499), .Z(n16492) );
  NANDN U17205 ( .A(n16475), .B(n16474), .Z(n16479) );
  OR U17206 ( .A(n16477), .B(n16476), .Z(n16478) );
  AND U17207 ( .A(n16479), .B(n16478), .Z(n16491) );
  XNOR U17208 ( .A(n16492), .B(n16491), .Z(n16493) );
  XNOR U17209 ( .A(n16494), .B(n16493), .Z(n16485) );
  XNOR U17210 ( .A(n16486), .B(n16485), .Z(n16487) );
  XNOR U17211 ( .A(n16488), .B(n16487), .Z(n16629) );
  XNOR U17212 ( .A(sreg[349]), .B(n16629), .Z(n16631) );
  NANDN U17213 ( .A(sreg[348]), .B(n16480), .Z(n16484) );
  NAND U17214 ( .A(n16482), .B(n16481), .Z(n16483) );
  NAND U17215 ( .A(n16484), .B(n16483), .Z(n16630) );
  XNOR U17216 ( .A(n16631), .B(n16630), .Z(c[349]) );
  NANDN U17217 ( .A(n16486), .B(n16485), .Z(n16490) );
  NANDN U17218 ( .A(n16488), .B(n16487), .Z(n16489) );
  AND U17219 ( .A(n16490), .B(n16489), .Z(n16637) );
  NANDN U17220 ( .A(n16492), .B(n16491), .Z(n16496) );
  NANDN U17221 ( .A(n16494), .B(n16493), .Z(n16495) );
  AND U17222 ( .A(n16496), .B(n16495), .Z(n16635) );
  NANDN U17223 ( .A(n16498), .B(n16497), .Z(n16502) );
  NAND U17224 ( .A(n16500), .B(n16499), .Z(n16501) );
  AND U17225 ( .A(n16502), .B(n16501), .Z(n16642) );
  NANDN U17226 ( .A(n16504), .B(n16503), .Z(n16508) );
  NANDN U17227 ( .A(n16506), .B(n16505), .Z(n16507) );
  AND U17228 ( .A(n16508), .B(n16507), .Z(n16647) );
  NANDN U17229 ( .A(n16510), .B(n16509), .Z(n16514) );
  NAND U17230 ( .A(n16512), .B(n16511), .Z(n16513) );
  AND U17231 ( .A(n16514), .B(n16513), .Z(n16646) );
  XNOR U17232 ( .A(n16647), .B(n16646), .Z(n16649) );
  NANDN U17233 ( .A(n16516), .B(n16515), .Z(n16520) );
  NANDN U17234 ( .A(n16518), .B(n16517), .Z(n16519) );
  AND U17235 ( .A(n16520), .B(n16519), .Z(n16726) );
  NAND U17236 ( .A(n38385), .B(n16521), .Z(n16523) );
  XOR U17237 ( .A(b[27]), .B(a[100]), .Z(n16670) );
  NAND U17238 ( .A(n38343), .B(n16670), .Z(n16522) );
  AND U17239 ( .A(n16523), .B(n16522), .Z(n16733) );
  NAND U17240 ( .A(n183), .B(n16524), .Z(n16526) );
  XOR U17241 ( .A(b[5]), .B(a[122]), .Z(n16673) );
  NAND U17242 ( .A(n36296), .B(n16673), .Z(n16525) );
  AND U17243 ( .A(n16526), .B(n16525), .Z(n16731) );
  NAND U17244 ( .A(n190), .B(n16527), .Z(n16529) );
  XOR U17245 ( .A(b[19]), .B(a[108]), .Z(n16676) );
  NAND U17246 ( .A(n37821), .B(n16676), .Z(n16528) );
  NAND U17247 ( .A(n16529), .B(n16528), .Z(n16730) );
  XNOR U17248 ( .A(n16731), .B(n16730), .Z(n16732) );
  XNOR U17249 ( .A(n16733), .B(n16732), .Z(n16724) );
  NAND U17250 ( .A(n38470), .B(n16530), .Z(n16532) );
  XOR U17251 ( .A(b[31]), .B(a[96]), .Z(n16679) );
  NAND U17252 ( .A(n38453), .B(n16679), .Z(n16531) );
  AND U17253 ( .A(n16532), .B(n16531), .Z(n16691) );
  NAND U17254 ( .A(n181), .B(n16533), .Z(n16535) );
  XOR U17255 ( .A(b[3]), .B(a[124]), .Z(n16682) );
  NAND U17256 ( .A(n182), .B(n16682), .Z(n16534) );
  AND U17257 ( .A(n16535), .B(n16534), .Z(n16689) );
  NAND U17258 ( .A(n189), .B(n16536), .Z(n16538) );
  XOR U17259 ( .A(b[17]), .B(a[110]), .Z(n16685) );
  NAND U17260 ( .A(n37652), .B(n16685), .Z(n16537) );
  NAND U17261 ( .A(n16538), .B(n16537), .Z(n16688) );
  XNOR U17262 ( .A(n16689), .B(n16688), .Z(n16690) );
  XOR U17263 ( .A(n16691), .B(n16690), .Z(n16725) );
  XOR U17264 ( .A(n16724), .B(n16725), .Z(n16727) );
  XOR U17265 ( .A(n16726), .B(n16727), .Z(n16659) );
  NANDN U17266 ( .A(n16540), .B(n16539), .Z(n16544) );
  NANDN U17267 ( .A(n16542), .B(n16541), .Z(n16543) );
  AND U17268 ( .A(n16544), .B(n16543), .Z(n16712) );
  NANDN U17269 ( .A(n16546), .B(n16545), .Z(n16550) );
  NANDN U17270 ( .A(n16548), .B(n16547), .Z(n16549) );
  NAND U17271 ( .A(n16550), .B(n16549), .Z(n16713) );
  XNOR U17272 ( .A(n16712), .B(n16713), .Z(n16714) );
  NANDN U17273 ( .A(n16552), .B(n16551), .Z(n16556) );
  NANDN U17274 ( .A(n16554), .B(n16553), .Z(n16555) );
  NAND U17275 ( .A(n16556), .B(n16555), .Z(n16715) );
  XNOR U17276 ( .A(n16714), .B(n16715), .Z(n16658) );
  XNOR U17277 ( .A(n16659), .B(n16658), .Z(n16661) );
  NANDN U17278 ( .A(n16558), .B(n16557), .Z(n16562) );
  NANDN U17279 ( .A(n16560), .B(n16559), .Z(n16561) );
  AND U17280 ( .A(n16562), .B(n16561), .Z(n16660) );
  XOR U17281 ( .A(n16661), .B(n16660), .Z(n16775) );
  NANDN U17282 ( .A(n16564), .B(n16563), .Z(n16568) );
  NANDN U17283 ( .A(n16566), .B(n16565), .Z(n16567) );
  AND U17284 ( .A(n16568), .B(n16567), .Z(n16772) );
  NANDN U17285 ( .A(n16570), .B(n16569), .Z(n16574) );
  NANDN U17286 ( .A(n16572), .B(n16571), .Z(n16573) );
  AND U17287 ( .A(n16574), .B(n16573), .Z(n16655) );
  NANDN U17288 ( .A(n16576), .B(n16575), .Z(n16580) );
  OR U17289 ( .A(n16578), .B(n16577), .Z(n16579) );
  AND U17290 ( .A(n16580), .B(n16579), .Z(n16653) );
  NANDN U17291 ( .A(n16582), .B(n16581), .Z(n16586) );
  NANDN U17292 ( .A(n16584), .B(n16583), .Z(n16585) );
  AND U17293 ( .A(n16586), .B(n16585), .Z(n16719) );
  NANDN U17294 ( .A(n16588), .B(n16587), .Z(n16592) );
  NANDN U17295 ( .A(n16590), .B(n16589), .Z(n16591) );
  NAND U17296 ( .A(n16592), .B(n16591), .Z(n16718) );
  XNOR U17297 ( .A(n16719), .B(n16718), .Z(n16720) );
  NAND U17298 ( .A(b[0]), .B(a[126]), .Z(n16593) );
  XNOR U17299 ( .A(b[1]), .B(n16593), .Z(n16595) );
  NANDN U17300 ( .A(b[0]), .B(a[125]), .Z(n16594) );
  NAND U17301 ( .A(n16595), .B(n16594), .Z(n16667) );
  NAND U17302 ( .A(n194), .B(n16596), .Z(n16598) );
  XOR U17303 ( .A(b[29]), .B(a[98]), .Z(n16745) );
  NAND U17304 ( .A(n38456), .B(n16745), .Z(n16597) );
  AND U17305 ( .A(n16598), .B(n16597), .Z(n16665) );
  AND U17306 ( .A(b[31]), .B(a[94]), .Z(n16664) );
  XNOR U17307 ( .A(n16665), .B(n16664), .Z(n16666) );
  XNOR U17308 ( .A(n16667), .B(n16666), .Z(n16706) );
  NAND U17309 ( .A(n38185), .B(n16599), .Z(n16601) );
  XOR U17310 ( .A(b[23]), .B(a[104]), .Z(n16748) );
  NAND U17311 ( .A(n38132), .B(n16748), .Z(n16600) );
  AND U17312 ( .A(n16601), .B(n16600), .Z(n16739) );
  NAND U17313 ( .A(n184), .B(n16602), .Z(n16604) );
  XOR U17314 ( .A(b[7]), .B(a[120]), .Z(n16751) );
  NAND U17315 ( .A(n36592), .B(n16751), .Z(n16603) );
  AND U17316 ( .A(n16604), .B(n16603), .Z(n16737) );
  NAND U17317 ( .A(n38289), .B(n16605), .Z(n16607) );
  XOR U17318 ( .A(b[25]), .B(a[102]), .Z(n16754) );
  NAND U17319 ( .A(n38247), .B(n16754), .Z(n16606) );
  NAND U17320 ( .A(n16607), .B(n16606), .Z(n16736) );
  XNOR U17321 ( .A(n16737), .B(n16736), .Z(n16738) );
  XOR U17322 ( .A(n16739), .B(n16738), .Z(n16707) );
  XNOR U17323 ( .A(n16706), .B(n16707), .Z(n16708) );
  NAND U17324 ( .A(n187), .B(n16608), .Z(n16610) );
  XOR U17325 ( .A(b[13]), .B(a[114]), .Z(n16757) );
  NAND U17326 ( .A(n37295), .B(n16757), .Z(n16609) );
  AND U17327 ( .A(n16610), .B(n16609), .Z(n16701) );
  NAND U17328 ( .A(n186), .B(n16611), .Z(n16613) );
  XOR U17329 ( .A(b[11]), .B(a[116]), .Z(n16760) );
  NAND U17330 ( .A(n37097), .B(n16760), .Z(n16612) );
  NAND U17331 ( .A(n16613), .B(n16612), .Z(n16700) );
  XNOR U17332 ( .A(n16701), .B(n16700), .Z(n16702) );
  NAND U17333 ( .A(n188), .B(n16614), .Z(n16616) );
  XOR U17334 ( .A(b[15]), .B(a[112]), .Z(n16763) );
  NAND U17335 ( .A(n37382), .B(n16763), .Z(n16615) );
  AND U17336 ( .A(n16616), .B(n16615), .Z(n16697) );
  NAND U17337 ( .A(n38064), .B(n16617), .Z(n16619) );
  XOR U17338 ( .A(b[21]), .B(a[106]), .Z(n16766) );
  NAND U17339 ( .A(n37993), .B(n16766), .Z(n16618) );
  AND U17340 ( .A(n16619), .B(n16618), .Z(n16695) );
  NAND U17341 ( .A(n185), .B(n16620), .Z(n16622) );
  XOR U17342 ( .A(b[9]), .B(a[118]), .Z(n16769) );
  NAND U17343 ( .A(n36805), .B(n16769), .Z(n16621) );
  NAND U17344 ( .A(n16622), .B(n16621), .Z(n16694) );
  XNOR U17345 ( .A(n16695), .B(n16694), .Z(n16696) );
  XOR U17346 ( .A(n16697), .B(n16696), .Z(n16703) );
  XOR U17347 ( .A(n16702), .B(n16703), .Z(n16709) );
  XOR U17348 ( .A(n16708), .B(n16709), .Z(n16721) );
  XNOR U17349 ( .A(n16720), .B(n16721), .Z(n16652) );
  XNOR U17350 ( .A(n16653), .B(n16652), .Z(n16654) );
  XOR U17351 ( .A(n16655), .B(n16654), .Z(n16773) );
  XNOR U17352 ( .A(n16772), .B(n16773), .Z(n16774) );
  XNOR U17353 ( .A(n16775), .B(n16774), .Z(n16648) );
  XOR U17354 ( .A(n16649), .B(n16648), .Z(n16641) );
  NANDN U17355 ( .A(n16624), .B(n16623), .Z(n16628) );
  NANDN U17356 ( .A(n16626), .B(n16625), .Z(n16627) );
  AND U17357 ( .A(n16628), .B(n16627), .Z(n16640) );
  XOR U17358 ( .A(n16641), .B(n16640), .Z(n16643) );
  XNOR U17359 ( .A(n16642), .B(n16643), .Z(n16634) );
  XNOR U17360 ( .A(n16635), .B(n16634), .Z(n16636) );
  XNOR U17361 ( .A(n16637), .B(n16636), .Z(n16778) );
  XNOR U17362 ( .A(sreg[350]), .B(n16778), .Z(n16780) );
  NANDN U17363 ( .A(sreg[349]), .B(n16629), .Z(n16633) );
  NAND U17364 ( .A(n16631), .B(n16630), .Z(n16632) );
  NAND U17365 ( .A(n16633), .B(n16632), .Z(n16779) );
  XNOR U17366 ( .A(n16780), .B(n16779), .Z(c[350]) );
  NANDN U17367 ( .A(n16635), .B(n16634), .Z(n16639) );
  NANDN U17368 ( .A(n16637), .B(n16636), .Z(n16638) );
  AND U17369 ( .A(n16639), .B(n16638), .Z(n16786) );
  NANDN U17370 ( .A(n16641), .B(n16640), .Z(n16645) );
  NANDN U17371 ( .A(n16643), .B(n16642), .Z(n16644) );
  AND U17372 ( .A(n16645), .B(n16644), .Z(n16784) );
  NANDN U17373 ( .A(n16647), .B(n16646), .Z(n16651) );
  NAND U17374 ( .A(n16649), .B(n16648), .Z(n16650) );
  AND U17375 ( .A(n16651), .B(n16650), .Z(n16791) );
  NANDN U17376 ( .A(n16653), .B(n16652), .Z(n16657) );
  NANDN U17377 ( .A(n16655), .B(n16654), .Z(n16656) );
  AND U17378 ( .A(n16657), .B(n16656), .Z(n16796) );
  NANDN U17379 ( .A(n16659), .B(n16658), .Z(n16663) );
  NAND U17380 ( .A(n16661), .B(n16660), .Z(n16662) );
  AND U17381 ( .A(n16663), .B(n16662), .Z(n16795) );
  XNOR U17382 ( .A(n16796), .B(n16795), .Z(n16798) );
  NANDN U17383 ( .A(n16665), .B(n16664), .Z(n16669) );
  NANDN U17384 ( .A(n16667), .B(n16666), .Z(n16668) );
  AND U17385 ( .A(n16669), .B(n16668), .Z(n16875) );
  NAND U17386 ( .A(n38385), .B(n16670), .Z(n16672) );
  XOR U17387 ( .A(b[27]), .B(a[101]), .Z(n16819) );
  NAND U17388 ( .A(n38343), .B(n16819), .Z(n16671) );
  AND U17389 ( .A(n16672), .B(n16671), .Z(n16882) );
  NAND U17390 ( .A(n183), .B(n16673), .Z(n16675) );
  XOR U17391 ( .A(b[5]), .B(a[123]), .Z(n16822) );
  NAND U17392 ( .A(n36296), .B(n16822), .Z(n16674) );
  AND U17393 ( .A(n16675), .B(n16674), .Z(n16880) );
  NAND U17394 ( .A(n190), .B(n16676), .Z(n16678) );
  XOR U17395 ( .A(b[19]), .B(a[109]), .Z(n16825) );
  NAND U17396 ( .A(n37821), .B(n16825), .Z(n16677) );
  NAND U17397 ( .A(n16678), .B(n16677), .Z(n16879) );
  XNOR U17398 ( .A(n16880), .B(n16879), .Z(n16881) );
  XNOR U17399 ( .A(n16882), .B(n16881), .Z(n16873) );
  NAND U17400 ( .A(n38470), .B(n16679), .Z(n16681) );
  XOR U17401 ( .A(b[31]), .B(a[97]), .Z(n16828) );
  NAND U17402 ( .A(n38453), .B(n16828), .Z(n16680) );
  AND U17403 ( .A(n16681), .B(n16680), .Z(n16840) );
  NAND U17404 ( .A(n181), .B(n16682), .Z(n16684) );
  XOR U17405 ( .A(b[3]), .B(a[125]), .Z(n16831) );
  NAND U17406 ( .A(n182), .B(n16831), .Z(n16683) );
  AND U17407 ( .A(n16684), .B(n16683), .Z(n16838) );
  NAND U17408 ( .A(n189), .B(n16685), .Z(n16687) );
  XOR U17409 ( .A(b[17]), .B(a[111]), .Z(n16834) );
  NAND U17410 ( .A(n37652), .B(n16834), .Z(n16686) );
  NAND U17411 ( .A(n16687), .B(n16686), .Z(n16837) );
  XNOR U17412 ( .A(n16838), .B(n16837), .Z(n16839) );
  XOR U17413 ( .A(n16840), .B(n16839), .Z(n16874) );
  XOR U17414 ( .A(n16873), .B(n16874), .Z(n16876) );
  XOR U17415 ( .A(n16875), .B(n16876), .Z(n16808) );
  NANDN U17416 ( .A(n16689), .B(n16688), .Z(n16693) );
  NANDN U17417 ( .A(n16691), .B(n16690), .Z(n16692) );
  AND U17418 ( .A(n16693), .B(n16692), .Z(n16861) );
  NANDN U17419 ( .A(n16695), .B(n16694), .Z(n16699) );
  NANDN U17420 ( .A(n16697), .B(n16696), .Z(n16698) );
  NAND U17421 ( .A(n16699), .B(n16698), .Z(n16862) );
  XNOR U17422 ( .A(n16861), .B(n16862), .Z(n16863) );
  NANDN U17423 ( .A(n16701), .B(n16700), .Z(n16705) );
  NANDN U17424 ( .A(n16703), .B(n16702), .Z(n16704) );
  NAND U17425 ( .A(n16705), .B(n16704), .Z(n16864) );
  XNOR U17426 ( .A(n16863), .B(n16864), .Z(n16807) );
  XNOR U17427 ( .A(n16808), .B(n16807), .Z(n16810) );
  NANDN U17428 ( .A(n16707), .B(n16706), .Z(n16711) );
  NANDN U17429 ( .A(n16709), .B(n16708), .Z(n16710) );
  AND U17430 ( .A(n16711), .B(n16710), .Z(n16809) );
  XOR U17431 ( .A(n16810), .B(n16809), .Z(n16924) );
  NANDN U17432 ( .A(n16713), .B(n16712), .Z(n16717) );
  NANDN U17433 ( .A(n16715), .B(n16714), .Z(n16716) );
  AND U17434 ( .A(n16717), .B(n16716), .Z(n16921) );
  NANDN U17435 ( .A(n16719), .B(n16718), .Z(n16723) );
  NANDN U17436 ( .A(n16721), .B(n16720), .Z(n16722) );
  AND U17437 ( .A(n16723), .B(n16722), .Z(n16804) );
  NANDN U17438 ( .A(n16725), .B(n16724), .Z(n16729) );
  OR U17439 ( .A(n16727), .B(n16726), .Z(n16728) );
  AND U17440 ( .A(n16729), .B(n16728), .Z(n16802) );
  NANDN U17441 ( .A(n16731), .B(n16730), .Z(n16735) );
  NANDN U17442 ( .A(n16733), .B(n16732), .Z(n16734) );
  AND U17443 ( .A(n16735), .B(n16734), .Z(n16868) );
  NANDN U17444 ( .A(n16737), .B(n16736), .Z(n16741) );
  NANDN U17445 ( .A(n16739), .B(n16738), .Z(n16740) );
  NAND U17446 ( .A(n16741), .B(n16740), .Z(n16867) );
  XNOR U17447 ( .A(n16868), .B(n16867), .Z(n16869) );
  NAND U17448 ( .A(b[0]), .B(a[127]), .Z(n16742) );
  XNOR U17449 ( .A(b[1]), .B(n16742), .Z(n16744) );
  NANDN U17450 ( .A(b[0]), .B(a[126]), .Z(n16743) );
  NAND U17451 ( .A(n16744), .B(n16743), .Z(n16816) );
  NAND U17452 ( .A(n194), .B(n16745), .Z(n16747) );
  XOR U17453 ( .A(b[29]), .B(a[99]), .Z(n16894) );
  NAND U17454 ( .A(n38456), .B(n16894), .Z(n16746) );
  AND U17455 ( .A(n16747), .B(n16746), .Z(n16814) );
  AND U17456 ( .A(b[31]), .B(a[95]), .Z(n16813) );
  XNOR U17457 ( .A(n16814), .B(n16813), .Z(n16815) );
  XNOR U17458 ( .A(n16816), .B(n16815), .Z(n16855) );
  NAND U17459 ( .A(n38185), .B(n16748), .Z(n16750) );
  XOR U17460 ( .A(b[23]), .B(a[105]), .Z(n16897) );
  NAND U17461 ( .A(n38132), .B(n16897), .Z(n16749) );
  AND U17462 ( .A(n16750), .B(n16749), .Z(n16888) );
  NAND U17463 ( .A(n184), .B(n16751), .Z(n16753) );
  XOR U17464 ( .A(b[7]), .B(a[121]), .Z(n16900) );
  NAND U17465 ( .A(n36592), .B(n16900), .Z(n16752) );
  AND U17466 ( .A(n16753), .B(n16752), .Z(n16886) );
  NAND U17467 ( .A(n38289), .B(n16754), .Z(n16756) );
  XOR U17468 ( .A(b[25]), .B(a[103]), .Z(n16903) );
  NAND U17469 ( .A(n38247), .B(n16903), .Z(n16755) );
  NAND U17470 ( .A(n16756), .B(n16755), .Z(n16885) );
  XNOR U17471 ( .A(n16886), .B(n16885), .Z(n16887) );
  XOR U17472 ( .A(n16888), .B(n16887), .Z(n16856) );
  XNOR U17473 ( .A(n16855), .B(n16856), .Z(n16857) );
  NAND U17474 ( .A(n187), .B(n16757), .Z(n16759) );
  XOR U17475 ( .A(b[13]), .B(a[115]), .Z(n16906) );
  NAND U17476 ( .A(n37295), .B(n16906), .Z(n16758) );
  AND U17477 ( .A(n16759), .B(n16758), .Z(n16850) );
  NAND U17478 ( .A(n186), .B(n16760), .Z(n16762) );
  XOR U17479 ( .A(b[11]), .B(a[117]), .Z(n16909) );
  NAND U17480 ( .A(n37097), .B(n16909), .Z(n16761) );
  NAND U17481 ( .A(n16762), .B(n16761), .Z(n16849) );
  XNOR U17482 ( .A(n16850), .B(n16849), .Z(n16851) );
  NAND U17483 ( .A(n188), .B(n16763), .Z(n16765) );
  XOR U17484 ( .A(b[15]), .B(a[113]), .Z(n16912) );
  NAND U17485 ( .A(n37382), .B(n16912), .Z(n16764) );
  AND U17486 ( .A(n16765), .B(n16764), .Z(n16846) );
  NAND U17487 ( .A(n38064), .B(n16766), .Z(n16768) );
  XOR U17488 ( .A(b[21]), .B(a[107]), .Z(n16915) );
  NAND U17489 ( .A(n37993), .B(n16915), .Z(n16767) );
  AND U17490 ( .A(n16768), .B(n16767), .Z(n16844) );
  NAND U17491 ( .A(n185), .B(n16769), .Z(n16771) );
  XOR U17492 ( .A(b[9]), .B(a[119]), .Z(n16918) );
  NAND U17493 ( .A(n36805), .B(n16918), .Z(n16770) );
  NAND U17494 ( .A(n16771), .B(n16770), .Z(n16843) );
  XNOR U17495 ( .A(n16844), .B(n16843), .Z(n16845) );
  XOR U17496 ( .A(n16846), .B(n16845), .Z(n16852) );
  XOR U17497 ( .A(n16851), .B(n16852), .Z(n16858) );
  XOR U17498 ( .A(n16857), .B(n16858), .Z(n16870) );
  XNOR U17499 ( .A(n16869), .B(n16870), .Z(n16801) );
  XNOR U17500 ( .A(n16802), .B(n16801), .Z(n16803) );
  XOR U17501 ( .A(n16804), .B(n16803), .Z(n16922) );
  XNOR U17502 ( .A(n16921), .B(n16922), .Z(n16923) );
  XNOR U17503 ( .A(n16924), .B(n16923), .Z(n16797) );
  XOR U17504 ( .A(n16798), .B(n16797), .Z(n16790) );
  NANDN U17505 ( .A(n16773), .B(n16772), .Z(n16777) );
  NANDN U17506 ( .A(n16775), .B(n16774), .Z(n16776) );
  AND U17507 ( .A(n16777), .B(n16776), .Z(n16789) );
  XOR U17508 ( .A(n16790), .B(n16789), .Z(n16792) );
  XNOR U17509 ( .A(n16791), .B(n16792), .Z(n16783) );
  XNOR U17510 ( .A(n16784), .B(n16783), .Z(n16785) );
  XNOR U17511 ( .A(n16786), .B(n16785), .Z(n16927) );
  XNOR U17512 ( .A(sreg[351]), .B(n16927), .Z(n16929) );
  NANDN U17513 ( .A(sreg[350]), .B(n16778), .Z(n16782) );
  NAND U17514 ( .A(n16780), .B(n16779), .Z(n16781) );
  NAND U17515 ( .A(n16782), .B(n16781), .Z(n16928) );
  XNOR U17516 ( .A(n16929), .B(n16928), .Z(c[351]) );
  NANDN U17517 ( .A(n16784), .B(n16783), .Z(n16788) );
  NANDN U17518 ( .A(n16786), .B(n16785), .Z(n16787) );
  AND U17519 ( .A(n16788), .B(n16787), .Z(n16935) );
  NANDN U17520 ( .A(n16790), .B(n16789), .Z(n16794) );
  NANDN U17521 ( .A(n16792), .B(n16791), .Z(n16793) );
  AND U17522 ( .A(n16794), .B(n16793), .Z(n16933) );
  NANDN U17523 ( .A(n16796), .B(n16795), .Z(n16800) );
  NAND U17524 ( .A(n16798), .B(n16797), .Z(n16799) );
  AND U17525 ( .A(n16800), .B(n16799), .Z(n16940) );
  NANDN U17526 ( .A(n16802), .B(n16801), .Z(n16806) );
  NANDN U17527 ( .A(n16804), .B(n16803), .Z(n16805) );
  AND U17528 ( .A(n16806), .B(n16805), .Z(n16945) );
  NANDN U17529 ( .A(n16808), .B(n16807), .Z(n16812) );
  NAND U17530 ( .A(n16810), .B(n16809), .Z(n16811) );
  AND U17531 ( .A(n16812), .B(n16811), .Z(n16944) );
  XNOR U17532 ( .A(n16945), .B(n16944), .Z(n16947) );
  NANDN U17533 ( .A(n16814), .B(n16813), .Z(n16818) );
  NANDN U17534 ( .A(n16816), .B(n16815), .Z(n16817) );
  AND U17535 ( .A(n16818), .B(n16817), .Z(n17024) );
  NAND U17536 ( .A(n38385), .B(n16819), .Z(n16821) );
  XOR U17537 ( .A(b[27]), .B(a[102]), .Z(n16968) );
  NAND U17538 ( .A(n38343), .B(n16968), .Z(n16820) );
  AND U17539 ( .A(n16821), .B(n16820), .Z(n17031) );
  NAND U17540 ( .A(n183), .B(n16822), .Z(n16824) );
  XOR U17541 ( .A(b[5]), .B(a[124]), .Z(n16971) );
  NAND U17542 ( .A(n36296), .B(n16971), .Z(n16823) );
  AND U17543 ( .A(n16824), .B(n16823), .Z(n17029) );
  NAND U17544 ( .A(n190), .B(n16825), .Z(n16827) );
  XOR U17545 ( .A(b[19]), .B(a[110]), .Z(n16974) );
  NAND U17546 ( .A(n37821), .B(n16974), .Z(n16826) );
  NAND U17547 ( .A(n16827), .B(n16826), .Z(n17028) );
  XNOR U17548 ( .A(n17029), .B(n17028), .Z(n17030) );
  XNOR U17549 ( .A(n17031), .B(n17030), .Z(n17022) );
  NAND U17550 ( .A(n38470), .B(n16828), .Z(n16830) );
  XOR U17551 ( .A(b[31]), .B(a[98]), .Z(n16977) );
  NAND U17552 ( .A(n38453), .B(n16977), .Z(n16829) );
  AND U17553 ( .A(n16830), .B(n16829), .Z(n16989) );
  NAND U17554 ( .A(n181), .B(n16831), .Z(n16833) );
  XOR U17555 ( .A(b[3]), .B(a[126]), .Z(n16980) );
  NAND U17556 ( .A(n182), .B(n16980), .Z(n16832) );
  AND U17557 ( .A(n16833), .B(n16832), .Z(n16987) );
  NAND U17558 ( .A(n189), .B(n16834), .Z(n16836) );
  XOR U17559 ( .A(b[17]), .B(a[112]), .Z(n16983) );
  NAND U17560 ( .A(n37652), .B(n16983), .Z(n16835) );
  NAND U17561 ( .A(n16836), .B(n16835), .Z(n16986) );
  XNOR U17562 ( .A(n16987), .B(n16986), .Z(n16988) );
  XOR U17563 ( .A(n16989), .B(n16988), .Z(n17023) );
  XOR U17564 ( .A(n17022), .B(n17023), .Z(n17025) );
  XOR U17565 ( .A(n17024), .B(n17025), .Z(n16957) );
  NANDN U17566 ( .A(n16838), .B(n16837), .Z(n16842) );
  NANDN U17567 ( .A(n16840), .B(n16839), .Z(n16841) );
  AND U17568 ( .A(n16842), .B(n16841), .Z(n17010) );
  NANDN U17569 ( .A(n16844), .B(n16843), .Z(n16848) );
  NANDN U17570 ( .A(n16846), .B(n16845), .Z(n16847) );
  NAND U17571 ( .A(n16848), .B(n16847), .Z(n17011) );
  XNOR U17572 ( .A(n17010), .B(n17011), .Z(n17012) );
  NANDN U17573 ( .A(n16850), .B(n16849), .Z(n16854) );
  NANDN U17574 ( .A(n16852), .B(n16851), .Z(n16853) );
  NAND U17575 ( .A(n16854), .B(n16853), .Z(n17013) );
  XNOR U17576 ( .A(n17012), .B(n17013), .Z(n16956) );
  XNOR U17577 ( .A(n16957), .B(n16956), .Z(n16959) );
  NANDN U17578 ( .A(n16856), .B(n16855), .Z(n16860) );
  NANDN U17579 ( .A(n16858), .B(n16857), .Z(n16859) );
  AND U17580 ( .A(n16860), .B(n16859), .Z(n16958) );
  XOR U17581 ( .A(n16959), .B(n16958), .Z(n17073) );
  NANDN U17582 ( .A(n16862), .B(n16861), .Z(n16866) );
  NANDN U17583 ( .A(n16864), .B(n16863), .Z(n16865) );
  AND U17584 ( .A(n16866), .B(n16865), .Z(n17070) );
  NANDN U17585 ( .A(n16868), .B(n16867), .Z(n16872) );
  NANDN U17586 ( .A(n16870), .B(n16869), .Z(n16871) );
  AND U17587 ( .A(n16872), .B(n16871), .Z(n16953) );
  NANDN U17588 ( .A(n16874), .B(n16873), .Z(n16878) );
  OR U17589 ( .A(n16876), .B(n16875), .Z(n16877) );
  AND U17590 ( .A(n16878), .B(n16877), .Z(n16951) );
  NANDN U17591 ( .A(n16880), .B(n16879), .Z(n16884) );
  NANDN U17592 ( .A(n16882), .B(n16881), .Z(n16883) );
  AND U17593 ( .A(n16884), .B(n16883), .Z(n17017) );
  NANDN U17594 ( .A(n16886), .B(n16885), .Z(n16890) );
  NANDN U17595 ( .A(n16888), .B(n16887), .Z(n16889) );
  NAND U17596 ( .A(n16890), .B(n16889), .Z(n17016) );
  XNOR U17597 ( .A(n17017), .B(n17016), .Z(n17018) );
  NAND U17598 ( .A(b[0]), .B(a[128]), .Z(n16891) );
  XNOR U17599 ( .A(b[1]), .B(n16891), .Z(n16893) );
  NANDN U17600 ( .A(b[0]), .B(a[127]), .Z(n16892) );
  NAND U17601 ( .A(n16893), .B(n16892), .Z(n16965) );
  NAND U17602 ( .A(n194), .B(n16894), .Z(n16896) );
  XOR U17603 ( .A(b[29]), .B(a[100]), .Z(n17043) );
  NAND U17604 ( .A(n38456), .B(n17043), .Z(n16895) );
  AND U17605 ( .A(n16896), .B(n16895), .Z(n16963) );
  AND U17606 ( .A(b[31]), .B(a[96]), .Z(n16962) );
  XNOR U17607 ( .A(n16963), .B(n16962), .Z(n16964) );
  XNOR U17608 ( .A(n16965), .B(n16964), .Z(n17004) );
  NAND U17609 ( .A(n38185), .B(n16897), .Z(n16899) );
  XOR U17610 ( .A(b[23]), .B(a[106]), .Z(n17046) );
  NAND U17611 ( .A(n38132), .B(n17046), .Z(n16898) );
  AND U17612 ( .A(n16899), .B(n16898), .Z(n17037) );
  NAND U17613 ( .A(n184), .B(n16900), .Z(n16902) );
  XOR U17614 ( .A(b[7]), .B(a[122]), .Z(n17049) );
  NAND U17615 ( .A(n36592), .B(n17049), .Z(n16901) );
  AND U17616 ( .A(n16902), .B(n16901), .Z(n17035) );
  NAND U17617 ( .A(n38289), .B(n16903), .Z(n16905) );
  XOR U17618 ( .A(b[25]), .B(a[104]), .Z(n17052) );
  NAND U17619 ( .A(n38247), .B(n17052), .Z(n16904) );
  NAND U17620 ( .A(n16905), .B(n16904), .Z(n17034) );
  XNOR U17621 ( .A(n17035), .B(n17034), .Z(n17036) );
  XOR U17622 ( .A(n17037), .B(n17036), .Z(n17005) );
  XNOR U17623 ( .A(n17004), .B(n17005), .Z(n17006) );
  NAND U17624 ( .A(n187), .B(n16906), .Z(n16908) );
  XOR U17625 ( .A(b[13]), .B(a[116]), .Z(n17055) );
  NAND U17626 ( .A(n37295), .B(n17055), .Z(n16907) );
  AND U17627 ( .A(n16908), .B(n16907), .Z(n16999) );
  NAND U17628 ( .A(n186), .B(n16909), .Z(n16911) );
  XOR U17629 ( .A(b[11]), .B(a[118]), .Z(n17058) );
  NAND U17630 ( .A(n37097), .B(n17058), .Z(n16910) );
  NAND U17631 ( .A(n16911), .B(n16910), .Z(n16998) );
  XNOR U17632 ( .A(n16999), .B(n16998), .Z(n17000) );
  NAND U17633 ( .A(n188), .B(n16912), .Z(n16914) );
  XOR U17634 ( .A(b[15]), .B(a[114]), .Z(n17061) );
  NAND U17635 ( .A(n37382), .B(n17061), .Z(n16913) );
  AND U17636 ( .A(n16914), .B(n16913), .Z(n16995) );
  NAND U17637 ( .A(n38064), .B(n16915), .Z(n16917) );
  XOR U17638 ( .A(b[21]), .B(a[108]), .Z(n17064) );
  NAND U17639 ( .A(n37993), .B(n17064), .Z(n16916) );
  AND U17640 ( .A(n16917), .B(n16916), .Z(n16993) );
  NAND U17641 ( .A(n185), .B(n16918), .Z(n16920) );
  XOR U17642 ( .A(b[9]), .B(a[120]), .Z(n17067) );
  NAND U17643 ( .A(n36805), .B(n17067), .Z(n16919) );
  NAND U17644 ( .A(n16920), .B(n16919), .Z(n16992) );
  XNOR U17645 ( .A(n16993), .B(n16992), .Z(n16994) );
  XOR U17646 ( .A(n16995), .B(n16994), .Z(n17001) );
  XOR U17647 ( .A(n17000), .B(n17001), .Z(n17007) );
  XOR U17648 ( .A(n17006), .B(n17007), .Z(n17019) );
  XNOR U17649 ( .A(n17018), .B(n17019), .Z(n16950) );
  XNOR U17650 ( .A(n16951), .B(n16950), .Z(n16952) );
  XOR U17651 ( .A(n16953), .B(n16952), .Z(n17071) );
  XNOR U17652 ( .A(n17070), .B(n17071), .Z(n17072) );
  XNOR U17653 ( .A(n17073), .B(n17072), .Z(n16946) );
  XOR U17654 ( .A(n16947), .B(n16946), .Z(n16939) );
  NANDN U17655 ( .A(n16922), .B(n16921), .Z(n16926) );
  NANDN U17656 ( .A(n16924), .B(n16923), .Z(n16925) );
  AND U17657 ( .A(n16926), .B(n16925), .Z(n16938) );
  XOR U17658 ( .A(n16939), .B(n16938), .Z(n16941) );
  XNOR U17659 ( .A(n16940), .B(n16941), .Z(n16932) );
  XNOR U17660 ( .A(n16933), .B(n16932), .Z(n16934) );
  XNOR U17661 ( .A(n16935), .B(n16934), .Z(n17076) );
  XNOR U17662 ( .A(sreg[352]), .B(n17076), .Z(n17078) );
  NANDN U17663 ( .A(sreg[351]), .B(n16927), .Z(n16931) );
  NAND U17664 ( .A(n16929), .B(n16928), .Z(n16930) );
  NAND U17665 ( .A(n16931), .B(n16930), .Z(n17077) );
  XNOR U17666 ( .A(n17078), .B(n17077), .Z(c[352]) );
  NANDN U17667 ( .A(n16933), .B(n16932), .Z(n16937) );
  NANDN U17668 ( .A(n16935), .B(n16934), .Z(n16936) );
  AND U17669 ( .A(n16937), .B(n16936), .Z(n17084) );
  NANDN U17670 ( .A(n16939), .B(n16938), .Z(n16943) );
  NANDN U17671 ( .A(n16941), .B(n16940), .Z(n16942) );
  AND U17672 ( .A(n16943), .B(n16942), .Z(n17082) );
  NANDN U17673 ( .A(n16945), .B(n16944), .Z(n16949) );
  NAND U17674 ( .A(n16947), .B(n16946), .Z(n16948) );
  AND U17675 ( .A(n16949), .B(n16948), .Z(n17089) );
  NANDN U17676 ( .A(n16951), .B(n16950), .Z(n16955) );
  NANDN U17677 ( .A(n16953), .B(n16952), .Z(n16954) );
  AND U17678 ( .A(n16955), .B(n16954), .Z(n17218) );
  NANDN U17679 ( .A(n16957), .B(n16956), .Z(n16961) );
  NAND U17680 ( .A(n16959), .B(n16958), .Z(n16960) );
  AND U17681 ( .A(n16961), .B(n16960), .Z(n17217) );
  XNOR U17682 ( .A(n17218), .B(n17217), .Z(n17220) );
  NANDN U17683 ( .A(n16963), .B(n16962), .Z(n16967) );
  NANDN U17684 ( .A(n16965), .B(n16964), .Z(n16966) );
  AND U17685 ( .A(n16967), .B(n16966), .Z(n17165) );
  NAND U17686 ( .A(n38385), .B(n16968), .Z(n16970) );
  XOR U17687 ( .A(b[27]), .B(a[103]), .Z(n17111) );
  NAND U17688 ( .A(n38343), .B(n17111), .Z(n16969) );
  AND U17689 ( .A(n16970), .B(n16969), .Z(n17172) );
  NAND U17690 ( .A(n183), .B(n16971), .Z(n16973) );
  XOR U17691 ( .A(b[5]), .B(a[125]), .Z(n17114) );
  NAND U17692 ( .A(n36296), .B(n17114), .Z(n16972) );
  AND U17693 ( .A(n16973), .B(n16972), .Z(n17170) );
  NAND U17694 ( .A(n190), .B(n16974), .Z(n16976) );
  XOR U17695 ( .A(b[19]), .B(a[111]), .Z(n17117) );
  NAND U17696 ( .A(n37821), .B(n17117), .Z(n16975) );
  NAND U17697 ( .A(n16976), .B(n16975), .Z(n17169) );
  XNOR U17698 ( .A(n17170), .B(n17169), .Z(n17171) );
  XNOR U17699 ( .A(n17172), .B(n17171), .Z(n17163) );
  NAND U17700 ( .A(n38470), .B(n16977), .Z(n16979) );
  XOR U17701 ( .A(b[31]), .B(a[99]), .Z(n17120) );
  NAND U17702 ( .A(n38453), .B(n17120), .Z(n16978) );
  AND U17703 ( .A(n16979), .B(n16978), .Z(n17132) );
  NAND U17704 ( .A(n181), .B(n16980), .Z(n16982) );
  XOR U17705 ( .A(b[3]), .B(a[127]), .Z(n17123) );
  NAND U17706 ( .A(n182), .B(n17123), .Z(n16981) );
  AND U17707 ( .A(n16982), .B(n16981), .Z(n17130) );
  NAND U17708 ( .A(n189), .B(n16983), .Z(n16985) );
  XOR U17709 ( .A(b[17]), .B(a[113]), .Z(n17126) );
  NAND U17710 ( .A(n37652), .B(n17126), .Z(n16984) );
  NAND U17711 ( .A(n16985), .B(n16984), .Z(n17129) );
  XNOR U17712 ( .A(n17130), .B(n17129), .Z(n17131) );
  XOR U17713 ( .A(n17132), .B(n17131), .Z(n17164) );
  XOR U17714 ( .A(n17163), .B(n17164), .Z(n17166) );
  XOR U17715 ( .A(n17165), .B(n17166), .Z(n17100) );
  NANDN U17716 ( .A(n16987), .B(n16986), .Z(n16991) );
  NANDN U17717 ( .A(n16989), .B(n16988), .Z(n16990) );
  AND U17718 ( .A(n16991), .B(n16990), .Z(n17153) );
  NANDN U17719 ( .A(n16993), .B(n16992), .Z(n16997) );
  NANDN U17720 ( .A(n16995), .B(n16994), .Z(n16996) );
  NAND U17721 ( .A(n16997), .B(n16996), .Z(n17154) );
  XNOR U17722 ( .A(n17153), .B(n17154), .Z(n17155) );
  NANDN U17723 ( .A(n16999), .B(n16998), .Z(n17003) );
  NANDN U17724 ( .A(n17001), .B(n17000), .Z(n17002) );
  NAND U17725 ( .A(n17003), .B(n17002), .Z(n17156) );
  XNOR U17726 ( .A(n17155), .B(n17156), .Z(n17099) );
  XNOR U17727 ( .A(n17100), .B(n17099), .Z(n17102) );
  NANDN U17728 ( .A(n17005), .B(n17004), .Z(n17009) );
  NANDN U17729 ( .A(n17007), .B(n17006), .Z(n17008) );
  AND U17730 ( .A(n17009), .B(n17008), .Z(n17101) );
  XOR U17731 ( .A(n17102), .B(n17101), .Z(n17214) );
  NANDN U17732 ( .A(n17011), .B(n17010), .Z(n17015) );
  NANDN U17733 ( .A(n17013), .B(n17012), .Z(n17014) );
  AND U17734 ( .A(n17015), .B(n17014), .Z(n17211) );
  NANDN U17735 ( .A(n17017), .B(n17016), .Z(n17021) );
  NANDN U17736 ( .A(n17019), .B(n17018), .Z(n17020) );
  AND U17737 ( .A(n17021), .B(n17020), .Z(n17096) );
  NANDN U17738 ( .A(n17023), .B(n17022), .Z(n17027) );
  OR U17739 ( .A(n17025), .B(n17024), .Z(n17026) );
  AND U17740 ( .A(n17027), .B(n17026), .Z(n17094) );
  NANDN U17741 ( .A(n17029), .B(n17028), .Z(n17033) );
  NANDN U17742 ( .A(n17031), .B(n17030), .Z(n17032) );
  AND U17743 ( .A(n17033), .B(n17032), .Z(n17160) );
  NANDN U17744 ( .A(n17035), .B(n17034), .Z(n17039) );
  NANDN U17745 ( .A(n17037), .B(n17036), .Z(n17038) );
  NAND U17746 ( .A(n17039), .B(n17038), .Z(n17159) );
  XNOR U17747 ( .A(n17160), .B(n17159), .Z(n17162) );
  NAND U17748 ( .A(b[0]), .B(a[129]), .Z(n17040) );
  XNOR U17749 ( .A(b[1]), .B(n17040), .Z(n17042) );
  NANDN U17750 ( .A(b[0]), .B(a[128]), .Z(n17041) );
  NAND U17751 ( .A(n17042), .B(n17041), .Z(n17108) );
  NAND U17752 ( .A(n194), .B(n17043), .Z(n17045) );
  XOR U17753 ( .A(b[29]), .B(a[101]), .Z(n17181) );
  NAND U17754 ( .A(n38456), .B(n17181), .Z(n17044) );
  AND U17755 ( .A(n17045), .B(n17044), .Z(n17106) );
  AND U17756 ( .A(b[31]), .B(a[97]), .Z(n17105) );
  XNOR U17757 ( .A(n17106), .B(n17105), .Z(n17107) );
  XNOR U17758 ( .A(n17108), .B(n17107), .Z(n17148) );
  NAND U17759 ( .A(n38185), .B(n17046), .Z(n17048) );
  XOR U17760 ( .A(b[23]), .B(a[107]), .Z(n17187) );
  NAND U17761 ( .A(n38132), .B(n17187), .Z(n17047) );
  AND U17762 ( .A(n17048), .B(n17047), .Z(n17177) );
  NAND U17763 ( .A(n184), .B(n17049), .Z(n17051) );
  XOR U17764 ( .A(b[7]), .B(a[123]), .Z(n17190) );
  NAND U17765 ( .A(n36592), .B(n17190), .Z(n17050) );
  AND U17766 ( .A(n17051), .B(n17050), .Z(n17176) );
  NAND U17767 ( .A(n38289), .B(n17052), .Z(n17054) );
  XOR U17768 ( .A(b[25]), .B(a[105]), .Z(n17193) );
  NAND U17769 ( .A(n38247), .B(n17193), .Z(n17053) );
  NAND U17770 ( .A(n17054), .B(n17053), .Z(n17175) );
  XOR U17771 ( .A(n17176), .B(n17175), .Z(n17178) );
  XOR U17772 ( .A(n17177), .B(n17178), .Z(n17147) );
  XOR U17773 ( .A(n17148), .B(n17147), .Z(n17150) );
  NAND U17774 ( .A(n187), .B(n17055), .Z(n17057) );
  XOR U17775 ( .A(b[13]), .B(a[117]), .Z(n17196) );
  NAND U17776 ( .A(n37295), .B(n17196), .Z(n17056) );
  AND U17777 ( .A(n17057), .B(n17056), .Z(n17142) );
  NAND U17778 ( .A(n186), .B(n17058), .Z(n17060) );
  XOR U17779 ( .A(b[11]), .B(a[119]), .Z(n17199) );
  NAND U17780 ( .A(n37097), .B(n17199), .Z(n17059) );
  NAND U17781 ( .A(n17060), .B(n17059), .Z(n17141) );
  XNOR U17782 ( .A(n17142), .B(n17141), .Z(n17144) );
  NAND U17783 ( .A(n188), .B(n17061), .Z(n17063) );
  XOR U17784 ( .A(b[15]), .B(a[115]), .Z(n17202) );
  NAND U17785 ( .A(n37382), .B(n17202), .Z(n17062) );
  AND U17786 ( .A(n17063), .B(n17062), .Z(n17138) );
  NAND U17787 ( .A(n38064), .B(n17064), .Z(n17066) );
  XOR U17788 ( .A(b[21]), .B(a[109]), .Z(n17205) );
  NAND U17789 ( .A(n37993), .B(n17205), .Z(n17065) );
  AND U17790 ( .A(n17066), .B(n17065), .Z(n17136) );
  NAND U17791 ( .A(n185), .B(n17067), .Z(n17069) );
  XOR U17792 ( .A(b[9]), .B(a[121]), .Z(n17208) );
  NAND U17793 ( .A(n36805), .B(n17208), .Z(n17068) );
  NAND U17794 ( .A(n17069), .B(n17068), .Z(n17135) );
  XNOR U17795 ( .A(n17136), .B(n17135), .Z(n17137) );
  XNOR U17796 ( .A(n17138), .B(n17137), .Z(n17143) );
  XOR U17797 ( .A(n17144), .B(n17143), .Z(n17149) );
  XNOR U17798 ( .A(n17150), .B(n17149), .Z(n17161) );
  XNOR U17799 ( .A(n17162), .B(n17161), .Z(n17093) );
  XNOR U17800 ( .A(n17094), .B(n17093), .Z(n17095) );
  XOR U17801 ( .A(n17096), .B(n17095), .Z(n17212) );
  XNOR U17802 ( .A(n17211), .B(n17212), .Z(n17213) );
  XNOR U17803 ( .A(n17214), .B(n17213), .Z(n17219) );
  XOR U17804 ( .A(n17220), .B(n17219), .Z(n17088) );
  NANDN U17805 ( .A(n17071), .B(n17070), .Z(n17075) );
  NANDN U17806 ( .A(n17073), .B(n17072), .Z(n17074) );
  AND U17807 ( .A(n17075), .B(n17074), .Z(n17087) );
  XOR U17808 ( .A(n17088), .B(n17087), .Z(n17090) );
  XNOR U17809 ( .A(n17089), .B(n17090), .Z(n17081) );
  XNOR U17810 ( .A(n17082), .B(n17081), .Z(n17083) );
  XNOR U17811 ( .A(n17084), .B(n17083), .Z(n17223) );
  XNOR U17812 ( .A(sreg[353]), .B(n17223), .Z(n17225) );
  NANDN U17813 ( .A(sreg[352]), .B(n17076), .Z(n17080) );
  NAND U17814 ( .A(n17078), .B(n17077), .Z(n17079) );
  NAND U17815 ( .A(n17080), .B(n17079), .Z(n17224) );
  XNOR U17816 ( .A(n17225), .B(n17224), .Z(c[353]) );
  NANDN U17817 ( .A(n17082), .B(n17081), .Z(n17086) );
  NANDN U17818 ( .A(n17084), .B(n17083), .Z(n17085) );
  AND U17819 ( .A(n17086), .B(n17085), .Z(n17231) );
  NANDN U17820 ( .A(n17088), .B(n17087), .Z(n17092) );
  NANDN U17821 ( .A(n17090), .B(n17089), .Z(n17091) );
  AND U17822 ( .A(n17092), .B(n17091), .Z(n17229) );
  NANDN U17823 ( .A(n17094), .B(n17093), .Z(n17098) );
  NANDN U17824 ( .A(n17096), .B(n17095), .Z(n17097) );
  AND U17825 ( .A(n17098), .B(n17097), .Z(n17367) );
  NANDN U17826 ( .A(n17100), .B(n17099), .Z(n17104) );
  NAND U17827 ( .A(n17102), .B(n17101), .Z(n17103) );
  AND U17828 ( .A(n17104), .B(n17103), .Z(n17366) );
  XNOR U17829 ( .A(n17367), .B(n17366), .Z(n17369) );
  NANDN U17830 ( .A(n17106), .B(n17105), .Z(n17110) );
  NANDN U17831 ( .A(n17108), .B(n17107), .Z(n17109) );
  AND U17832 ( .A(n17110), .B(n17109), .Z(n17302) );
  NAND U17833 ( .A(n38385), .B(n17111), .Z(n17113) );
  XOR U17834 ( .A(b[27]), .B(a[104]), .Z(n17246) );
  NAND U17835 ( .A(n38343), .B(n17246), .Z(n17112) );
  AND U17836 ( .A(n17113), .B(n17112), .Z(n17309) );
  NAND U17837 ( .A(n183), .B(n17114), .Z(n17116) );
  XOR U17838 ( .A(b[5]), .B(a[126]), .Z(n17249) );
  NAND U17839 ( .A(n36296), .B(n17249), .Z(n17115) );
  AND U17840 ( .A(n17116), .B(n17115), .Z(n17307) );
  NAND U17841 ( .A(n190), .B(n17117), .Z(n17119) );
  XOR U17842 ( .A(b[19]), .B(a[112]), .Z(n17252) );
  NAND U17843 ( .A(n37821), .B(n17252), .Z(n17118) );
  NAND U17844 ( .A(n17119), .B(n17118), .Z(n17306) );
  XNOR U17845 ( .A(n17307), .B(n17306), .Z(n17308) );
  XNOR U17846 ( .A(n17309), .B(n17308), .Z(n17300) );
  NAND U17847 ( .A(n38470), .B(n17120), .Z(n17122) );
  XOR U17848 ( .A(b[31]), .B(a[100]), .Z(n17255) );
  NAND U17849 ( .A(n38453), .B(n17255), .Z(n17121) );
  AND U17850 ( .A(n17122), .B(n17121), .Z(n17267) );
  NAND U17851 ( .A(n181), .B(n17123), .Z(n17125) );
  XOR U17852 ( .A(b[3]), .B(a[128]), .Z(n17258) );
  NAND U17853 ( .A(n182), .B(n17258), .Z(n17124) );
  AND U17854 ( .A(n17125), .B(n17124), .Z(n17265) );
  NAND U17855 ( .A(n189), .B(n17126), .Z(n17128) );
  XOR U17856 ( .A(b[17]), .B(a[114]), .Z(n17261) );
  NAND U17857 ( .A(n37652), .B(n17261), .Z(n17127) );
  NAND U17858 ( .A(n17128), .B(n17127), .Z(n17264) );
  XNOR U17859 ( .A(n17265), .B(n17264), .Z(n17266) );
  XOR U17860 ( .A(n17267), .B(n17266), .Z(n17301) );
  XOR U17861 ( .A(n17300), .B(n17301), .Z(n17303) );
  XOR U17862 ( .A(n17302), .B(n17303), .Z(n17349) );
  NANDN U17863 ( .A(n17130), .B(n17129), .Z(n17134) );
  NANDN U17864 ( .A(n17132), .B(n17131), .Z(n17133) );
  AND U17865 ( .A(n17134), .B(n17133), .Z(n17288) );
  NANDN U17866 ( .A(n17136), .B(n17135), .Z(n17140) );
  NANDN U17867 ( .A(n17138), .B(n17137), .Z(n17139) );
  NAND U17868 ( .A(n17140), .B(n17139), .Z(n17289) );
  XNOR U17869 ( .A(n17288), .B(n17289), .Z(n17290) );
  NANDN U17870 ( .A(n17142), .B(n17141), .Z(n17146) );
  NAND U17871 ( .A(n17144), .B(n17143), .Z(n17145) );
  NAND U17872 ( .A(n17146), .B(n17145), .Z(n17291) );
  XNOR U17873 ( .A(n17290), .B(n17291), .Z(n17348) );
  XNOR U17874 ( .A(n17349), .B(n17348), .Z(n17351) );
  NAND U17875 ( .A(n17148), .B(n17147), .Z(n17152) );
  NAND U17876 ( .A(n17150), .B(n17149), .Z(n17151) );
  AND U17877 ( .A(n17152), .B(n17151), .Z(n17350) );
  XOR U17878 ( .A(n17351), .B(n17350), .Z(n17363) );
  NANDN U17879 ( .A(n17154), .B(n17153), .Z(n17158) );
  NANDN U17880 ( .A(n17156), .B(n17155), .Z(n17157) );
  AND U17881 ( .A(n17158), .B(n17157), .Z(n17360) );
  NANDN U17882 ( .A(n17164), .B(n17163), .Z(n17168) );
  OR U17883 ( .A(n17166), .B(n17165), .Z(n17167) );
  AND U17884 ( .A(n17168), .B(n17167), .Z(n17355) );
  NANDN U17885 ( .A(n17170), .B(n17169), .Z(n17174) );
  NANDN U17886 ( .A(n17172), .B(n17171), .Z(n17173) );
  AND U17887 ( .A(n17174), .B(n17173), .Z(n17295) );
  NANDN U17888 ( .A(n17176), .B(n17175), .Z(n17180) );
  OR U17889 ( .A(n17178), .B(n17177), .Z(n17179) );
  NAND U17890 ( .A(n17180), .B(n17179), .Z(n17294) );
  XNOR U17891 ( .A(n17295), .B(n17294), .Z(n17296) );
  NAND U17892 ( .A(n194), .B(n17181), .Z(n17183) );
  XOR U17893 ( .A(b[29]), .B(a[102]), .Z(n17321) );
  NAND U17894 ( .A(n38456), .B(n17321), .Z(n17182) );
  AND U17895 ( .A(n17183), .B(n17182), .Z(n17241) );
  AND U17896 ( .A(b[31]), .B(a[98]), .Z(n17240) );
  XNOR U17897 ( .A(n17241), .B(n17240), .Z(n17242) );
  NAND U17898 ( .A(b[0]), .B(a[130]), .Z(n17184) );
  XNOR U17899 ( .A(b[1]), .B(n17184), .Z(n17186) );
  NANDN U17900 ( .A(b[0]), .B(a[129]), .Z(n17185) );
  NAND U17901 ( .A(n17186), .B(n17185), .Z(n17243) );
  XNOR U17902 ( .A(n17242), .B(n17243), .Z(n17282) );
  NAND U17903 ( .A(n38185), .B(n17187), .Z(n17189) );
  XOR U17904 ( .A(b[23]), .B(a[108]), .Z(n17324) );
  NAND U17905 ( .A(n38132), .B(n17324), .Z(n17188) );
  AND U17906 ( .A(n17189), .B(n17188), .Z(n17315) );
  NAND U17907 ( .A(n184), .B(n17190), .Z(n17192) );
  XOR U17908 ( .A(b[7]), .B(a[124]), .Z(n17327) );
  NAND U17909 ( .A(n36592), .B(n17327), .Z(n17191) );
  AND U17910 ( .A(n17192), .B(n17191), .Z(n17313) );
  NAND U17911 ( .A(n38289), .B(n17193), .Z(n17195) );
  XOR U17912 ( .A(b[25]), .B(a[106]), .Z(n17330) );
  NAND U17913 ( .A(n38247), .B(n17330), .Z(n17194) );
  NAND U17914 ( .A(n17195), .B(n17194), .Z(n17312) );
  XNOR U17915 ( .A(n17313), .B(n17312), .Z(n17314) );
  XOR U17916 ( .A(n17315), .B(n17314), .Z(n17283) );
  XNOR U17917 ( .A(n17282), .B(n17283), .Z(n17284) );
  NAND U17918 ( .A(n187), .B(n17196), .Z(n17198) );
  XOR U17919 ( .A(b[13]), .B(a[118]), .Z(n17333) );
  NAND U17920 ( .A(n37295), .B(n17333), .Z(n17197) );
  AND U17921 ( .A(n17198), .B(n17197), .Z(n17277) );
  NAND U17922 ( .A(n186), .B(n17199), .Z(n17201) );
  XOR U17923 ( .A(b[11]), .B(a[120]), .Z(n17336) );
  NAND U17924 ( .A(n37097), .B(n17336), .Z(n17200) );
  NAND U17925 ( .A(n17201), .B(n17200), .Z(n17276) );
  XNOR U17926 ( .A(n17277), .B(n17276), .Z(n17278) );
  NAND U17927 ( .A(n188), .B(n17202), .Z(n17204) );
  XOR U17928 ( .A(b[15]), .B(a[116]), .Z(n17339) );
  NAND U17929 ( .A(n37382), .B(n17339), .Z(n17203) );
  AND U17930 ( .A(n17204), .B(n17203), .Z(n17273) );
  NAND U17931 ( .A(n38064), .B(n17205), .Z(n17207) );
  XOR U17932 ( .A(b[21]), .B(a[110]), .Z(n17342) );
  NAND U17933 ( .A(n37993), .B(n17342), .Z(n17206) );
  AND U17934 ( .A(n17207), .B(n17206), .Z(n17271) );
  NAND U17935 ( .A(n185), .B(n17208), .Z(n17210) );
  XOR U17936 ( .A(b[9]), .B(a[122]), .Z(n17345) );
  NAND U17937 ( .A(n36805), .B(n17345), .Z(n17209) );
  NAND U17938 ( .A(n17210), .B(n17209), .Z(n17270) );
  XNOR U17939 ( .A(n17271), .B(n17270), .Z(n17272) );
  XOR U17940 ( .A(n17273), .B(n17272), .Z(n17279) );
  XOR U17941 ( .A(n17278), .B(n17279), .Z(n17285) );
  XOR U17942 ( .A(n17284), .B(n17285), .Z(n17297) );
  XNOR U17943 ( .A(n17296), .B(n17297), .Z(n17354) );
  XNOR U17944 ( .A(n17355), .B(n17354), .Z(n17356) );
  XOR U17945 ( .A(n17357), .B(n17356), .Z(n17361) );
  XNOR U17946 ( .A(n17360), .B(n17361), .Z(n17362) );
  XNOR U17947 ( .A(n17363), .B(n17362), .Z(n17368) );
  XOR U17948 ( .A(n17369), .B(n17368), .Z(n17235) );
  NANDN U17949 ( .A(n17212), .B(n17211), .Z(n17216) );
  NANDN U17950 ( .A(n17214), .B(n17213), .Z(n17215) );
  AND U17951 ( .A(n17216), .B(n17215), .Z(n17234) );
  XNOR U17952 ( .A(n17235), .B(n17234), .Z(n17236) );
  NANDN U17953 ( .A(n17218), .B(n17217), .Z(n17222) );
  NAND U17954 ( .A(n17220), .B(n17219), .Z(n17221) );
  NAND U17955 ( .A(n17222), .B(n17221), .Z(n17237) );
  XNOR U17956 ( .A(n17236), .B(n17237), .Z(n17228) );
  XNOR U17957 ( .A(n17229), .B(n17228), .Z(n17230) );
  XNOR U17958 ( .A(n17231), .B(n17230), .Z(n17372) );
  XNOR U17959 ( .A(sreg[354]), .B(n17372), .Z(n17374) );
  NANDN U17960 ( .A(sreg[353]), .B(n17223), .Z(n17227) );
  NAND U17961 ( .A(n17225), .B(n17224), .Z(n17226) );
  NAND U17962 ( .A(n17227), .B(n17226), .Z(n17373) );
  XNOR U17963 ( .A(n17374), .B(n17373), .Z(c[354]) );
  NANDN U17964 ( .A(n17229), .B(n17228), .Z(n17233) );
  NANDN U17965 ( .A(n17231), .B(n17230), .Z(n17232) );
  AND U17966 ( .A(n17233), .B(n17232), .Z(n17380) );
  NANDN U17967 ( .A(n17235), .B(n17234), .Z(n17239) );
  NANDN U17968 ( .A(n17237), .B(n17236), .Z(n17238) );
  AND U17969 ( .A(n17239), .B(n17238), .Z(n17378) );
  NANDN U17970 ( .A(n17241), .B(n17240), .Z(n17245) );
  NANDN U17971 ( .A(n17243), .B(n17242), .Z(n17244) );
  AND U17972 ( .A(n17245), .B(n17244), .Z(n17469) );
  NAND U17973 ( .A(n38385), .B(n17246), .Z(n17248) );
  XOR U17974 ( .A(b[27]), .B(a[105]), .Z(n17413) );
  NAND U17975 ( .A(n38343), .B(n17413), .Z(n17247) );
  AND U17976 ( .A(n17248), .B(n17247), .Z(n17476) );
  NAND U17977 ( .A(n183), .B(n17249), .Z(n17251) );
  XOR U17978 ( .A(b[5]), .B(a[127]), .Z(n17416) );
  NAND U17979 ( .A(n36296), .B(n17416), .Z(n17250) );
  AND U17980 ( .A(n17251), .B(n17250), .Z(n17474) );
  NAND U17981 ( .A(n190), .B(n17252), .Z(n17254) );
  XOR U17982 ( .A(b[19]), .B(a[113]), .Z(n17419) );
  NAND U17983 ( .A(n37821), .B(n17419), .Z(n17253) );
  NAND U17984 ( .A(n17254), .B(n17253), .Z(n17473) );
  XNOR U17985 ( .A(n17474), .B(n17473), .Z(n17475) );
  XNOR U17986 ( .A(n17476), .B(n17475), .Z(n17467) );
  NAND U17987 ( .A(n38470), .B(n17255), .Z(n17257) );
  XOR U17988 ( .A(b[31]), .B(a[101]), .Z(n17422) );
  NAND U17989 ( .A(n38453), .B(n17422), .Z(n17256) );
  AND U17990 ( .A(n17257), .B(n17256), .Z(n17434) );
  NAND U17991 ( .A(n181), .B(n17258), .Z(n17260) );
  XOR U17992 ( .A(b[3]), .B(a[129]), .Z(n17425) );
  NAND U17993 ( .A(n182), .B(n17425), .Z(n17259) );
  AND U17994 ( .A(n17260), .B(n17259), .Z(n17432) );
  NAND U17995 ( .A(n189), .B(n17261), .Z(n17263) );
  XOR U17996 ( .A(b[17]), .B(a[115]), .Z(n17428) );
  NAND U17997 ( .A(n37652), .B(n17428), .Z(n17262) );
  NAND U17998 ( .A(n17263), .B(n17262), .Z(n17431) );
  XNOR U17999 ( .A(n17432), .B(n17431), .Z(n17433) );
  XOR U18000 ( .A(n17434), .B(n17433), .Z(n17468) );
  XOR U18001 ( .A(n17467), .B(n17468), .Z(n17470) );
  XOR U18002 ( .A(n17469), .B(n17470), .Z(n17402) );
  NANDN U18003 ( .A(n17265), .B(n17264), .Z(n17269) );
  NANDN U18004 ( .A(n17267), .B(n17266), .Z(n17268) );
  AND U18005 ( .A(n17269), .B(n17268), .Z(n17455) );
  NANDN U18006 ( .A(n17271), .B(n17270), .Z(n17275) );
  NANDN U18007 ( .A(n17273), .B(n17272), .Z(n17274) );
  NAND U18008 ( .A(n17275), .B(n17274), .Z(n17456) );
  XNOR U18009 ( .A(n17455), .B(n17456), .Z(n17457) );
  NANDN U18010 ( .A(n17277), .B(n17276), .Z(n17281) );
  NANDN U18011 ( .A(n17279), .B(n17278), .Z(n17280) );
  NAND U18012 ( .A(n17281), .B(n17280), .Z(n17458) );
  XNOR U18013 ( .A(n17457), .B(n17458), .Z(n17401) );
  XNOR U18014 ( .A(n17402), .B(n17401), .Z(n17404) );
  NANDN U18015 ( .A(n17283), .B(n17282), .Z(n17287) );
  NANDN U18016 ( .A(n17285), .B(n17284), .Z(n17286) );
  AND U18017 ( .A(n17287), .B(n17286), .Z(n17403) );
  XOR U18018 ( .A(n17404), .B(n17403), .Z(n17517) );
  NANDN U18019 ( .A(n17289), .B(n17288), .Z(n17293) );
  NANDN U18020 ( .A(n17291), .B(n17290), .Z(n17292) );
  AND U18021 ( .A(n17293), .B(n17292), .Z(n17515) );
  NANDN U18022 ( .A(n17295), .B(n17294), .Z(n17299) );
  NANDN U18023 ( .A(n17297), .B(n17296), .Z(n17298) );
  AND U18024 ( .A(n17299), .B(n17298), .Z(n17398) );
  NANDN U18025 ( .A(n17301), .B(n17300), .Z(n17305) );
  OR U18026 ( .A(n17303), .B(n17302), .Z(n17304) );
  AND U18027 ( .A(n17305), .B(n17304), .Z(n17396) );
  NANDN U18028 ( .A(n17307), .B(n17306), .Z(n17311) );
  NANDN U18029 ( .A(n17309), .B(n17308), .Z(n17310) );
  AND U18030 ( .A(n17311), .B(n17310), .Z(n17462) );
  NANDN U18031 ( .A(n17313), .B(n17312), .Z(n17317) );
  NANDN U18032 ( .A(n17315), .B(n17314), .Z(n17316) );
  NAND U18033 ( .A(n17317), .B(n17316), .Z(n17461) );
  XNOR U18034 ( .A(n17462), .B(n17461), .Z(n17463) );
  NAND U18035 ( .A(b[0]), .B(a[131]), .Z(n17318) );
  XNOR U18036 ( .A(b[1]), .B(n17318), .Z(n17320) );
  NANDN U18037 ( .A(b[0]), .B(a[130]), .Z(n17319) );
  NAND U18038 ( .A(n17320), .B(n17319), .Z(n17410) );
  NAND U18039 ( .A(n194), .B(n17321), .Z(n17323) );
  XOR U18040 ( .A(b[29]), .B(a[103]), .Z(n17485) );
  NAND U18041 ( .A(n38456), .B(n17485), .Z(n17322) );
  AND U18042 ( .A(n17323), .B(n17322), .Z(n17408) );
  AND U18043 ( .A(b[31]), .B(a[99]), .Z(n17407) );
  XNOR U18044 ( .A(n17408), .B(n17407), .Z(n17409) );
  XNOR U18045 ( .A(n17410), .B(n17409), .Z(n17449) );
  NAND U18046 ( .A(n38185), .B(n17324), .Z(n17326) );
  XOR U18047 ( .A(b[23]), .B(a[109]), .Z(n17491) );
  NAND U18048 ( .A(n38132), .B(n17491), .Z(n17325) );
  AND U18049 ( .A(n17326), .B(n17325), .Z(n17482) );
  NAND U18050 ( .A(n184), .B(n17327), .Z(n17329) );
  XOR U18051 ( .A(b[7]), .B(a[125]), .Z(n17494) );
  NAND U18052 ( .A(n36592), .B(n17494), .Z(n17328) );
  AND U18053 ( .A(n17329), .B(n17328), .Z(n17480) );
  NAND U18054 ( .A(n38289), .B(n17330), .Z(n17332) );
  XOR U18055 ( .A(b[25]), .B(a[107]), .Z(n17497) );
  NAND U18056 ( .A(n38247), .B(n17497), .Z(n17331) );
  NAND U18057 ( .A(n17332), .B(n17331), .Z(n17479) );
  XNOR U18058 ( .A(n17480), .B(n17479), .Z(n17481) );
  XOR U18059 ( .A(n17482), .B(n17481), .Z(n17450) );
  XNOR U18060 ( .A(n17449), .B(n17450), .Z(n17451) );
  NAND U18061 ( .A(n187), .B(n17333), .Z(n17335) );
  XOR U18062 ( .A(b[13]), .B(a[119]), .Z(n17500) );
  NAND U18063 ( .A(n37295), .B(n17500), .Z(n17334) );
  AND U18064 ( .A(n17335), .B(n17334), .Z(n17444) );
  NAND U18065 ( .A(n186), .B(n17336), .Z(n17338) );
  XOR U18066 ( .A(b[11]), .B(a[121]), .Z(n17503) );
  NAND U18067 ( .A(n37097), .B(n17503), .Z(n17337) );
  NAND U18068 ( .A(n17338), .B(n17337), .Z(n17443) );
  XNOR U18069 ( .A(n17444), .B(n17443), .Z(n17445) );
  NAND U18070 ( .A(n188), .B(n17339), .Z(n17341) );
  XOR U18071 ( .A(b[15]), .B(a[117]), .Z(n17506) );
  NAND U18072 ( .A(n37382), .B(n17506), .Z(n17340) );
  AND U18073 ( .A(n17341), .B(n17340), .Z(n17440) );
  NAND U18074 ( .A(n38064), .B(n17342), .Z(n17344) );
  XOR U18075 ( .A(b[21]), .B(a[111]), .Z(n17509) );
  NAND U18076 ( .A(n37993), .B(n17509), .Z(n17343) );
  AND U18077 ( .A(n17344), .B(n17343), .Z(n17438) );
  NAND U18078 ( .A(n185), .B(n17345), .Z(n17347) );
  XOR U18079 ( .A(b[9]), .B(a[123]), .Z(n17512) );
  NAND U18080 ( .A(n36805), .B(n17512), .Z(n17346) );
  NAND U18081 ( .A(n17347), .B(n17346), .Z(n17437) );
  XNOR U18082 ( .A(n17438), .B(n17437), .Z(n17439) );
  XOR U18083 ( .A(n17440), .B(n17439), .Z(n17446) );
  XOR U18084 ( .A(n17445), .B(n17446), .Z(n17452) );
  XOR U18085 ( .A(n17451), .B(n17452), .Z(n17464) );
  XNOR U18086 ( .A(n17463), .B(n17464), .Z(n17395) );
  XNOR U18087 ( .A(n17396), .B(n17395), .Z(n17397) );
  XOR U18088 ( .A(n17398), .B(n17397), .Z(n17516) );
  XOR U18089 ( .A(n17515), .B(n17516), .Z(n17518) );
  XOR U18090 ( .A(n17517), .B(n17518), .Z(n17392) );
  NANDN U18091 ( .A(n17349), .B(n17348), .Z(n17353) );
  NAND U18092 ( .A(n17351), .B(n17350), .Z(n17352) );
  AND U18093 ( .A(n17353), .B(n17352), .Z(n17390) );
  NANDN U18094 ( .A(n17355), .B(n17354), .Z(n17359) );
  NANDN U18095 ( .A(n17357), .B(n17356), .Z(n17358) );
  AND U18096 ( .A(n17359), .B(n17358), .Z(n17389) );
  XNOR U18097 ( .A(n17390), .B(n17389), .Z(n17391) );
  XNOR U18098 ( .A(n17392), .B(n17391), .Z(n17383) );
  NANDN U18099 ( .A(n17361), .B(n17360), .Z(n17365) );
  NANDN U18100 ( .A(n17363), .B(n17362), .Z(n17364) );
  NAND U18101 ( .A(n17365), .B(n17364), .Z(n17384) );
  XNOR U18102 ( .A(n17383), .B(n17384), .Z(n17385) );
  NANDN U18103 ( .A(n17367), .B(n17366), .Z(n17371) );
  NAND U18104 ( .A(n17369), .B(n17368), .Z(n17370) );
  NAND U18105 ( .A(n17371), .B(n17370), .Z(n17386) );
  XNOR U18106 ( .A(n17385), .B(n17386), .Z(n17377) );
  XNOR U18107 ( .A(n17378), .B(n17377), .Z(n17379) );
  XNOR U18108 ( .A(n17380), .B(n17379), .Z(n17521) );
  XNOR U18109 ( .A(sreg[355]), .B(n17521), .Z(n17523) );
  NANDN U18110 ( .A(sreg[354]), .B(n17372), .Z(n17376) );
  NAND U18111 ( .A(n17374), .B(n17373), .Z(n17375) );
  NAND U18112 ( .A(n17376), .B(n17375), .Z(n17522) );
  XNOR U18113 ( .A(n17523), .B(n17522), .Z(c[355]) );
  NANDN U18114 ( .A(n17378), .B(n17377), .Z(n17382) );
  NANDN U18115 ( .A(n17380), .B(n17379), .Z(n17381) );
  AND U18116 ( .A(n17382), .B(n17381), .Z(n17529) );
  NANDN U18117 ( .A(n17384), .B(n17383), .Z(n17388) );
  NANDN U18118 ( .A(n17386), .B(n17385), .Z(n17387) );
  AND U18119 ( .A(n17388), .B(n17387), .Z(n17527) );
  NANDN U18120 ( .A(n17390), .B(n17389), .Z(n17394) );
  NANDN U18121 ( .A(n17392), .B(n17391), .Z(n17393) );
  AND U18122 ( .A(n17394), .B(n17393), .Z(n17535) );
  NANDN U18123 ( .A(n17396), .B(n17395), .Z(n17400) );
  NANDN U18124 ( .A(n17398), .B(n17397), .Z(n17399) );
  AND U18125 ( .A(n17400), .B(n17399), .Z(n17539) );
  NANDN U18126 ( .A(n17402), .B(n17401), .Z(n17406) );
  NAND U18127 ( .A(n17404), .B(n17403), .Z(n17405) );
  AND U18128 ( .A(n17406), .B(n17405), .Z(n17538) );
  XNOR U18129 ( .A(n17539), .B(n17538), .Z(n17541) );
  NANDN U18130 ( .A(n17408), .B(n17407), .Z(n17412) );
  NANDN U18131 ( .A(n17410), .B(n17409), .Z(n17411) );
  AND U18132 ( .A(n17412), .B(n17411), .Z(n17616) );
  NAND U18133 ( .A(n38385), .B(n17413), .Z(n17415) );
  XOR U18134 ( .A(b[27]), .B(a[106]), .Z(n17562) );
  NAND U18135 ( .A(n38343), .B(n17562), .Z(n17414) );
  AND U18136 ( .A(n17415), .B(n17414), .Z(n17623) );
  NAND U18137 ( .A(n183), .B(n17416), .Z(n17418) );
  XOR U18138 ( .A(b[5]), .B(a[128]), .Z(n17565) );
  NAND U18139 ( .A(n36296), .B(n17565), .Z(n17417) );
  AND U18140 ( .A(n17418), .B(n17417), .Z(n17621) );
  NAND U18141 ( .A(n190), .B(n17419), .Z(n17421) );
  XOR U18142 ( .A(b[19]), .B(a[114]), .Z(n17568) );
  NAND U18143 ( .A(n37821), .B(n17568), .Z(n17420) );
  NAND U18144 ( .A(n17421), .B(n17420), .Z(n17620) );
  XNOR U18145 ( .A(n17621), .B(n17620), .Z(n17622) );
  XNOR U18146 ( .A(n17623), .B(n17622), .Z(n17614) );
  NAND U18147 ( .A(n38470), .B(n17422), .Z(n17424) );
  XOR U18148 ( .A(b[31]), .B(a[102]), .Z(n17571) );
  NAND U18149 ( .A(n38453), .B(n17571), .Z(n17423) );
  AND U18150 ( .A(n17424), .B(n17423), .Z(n17583) );
  NAND U18151 ( .A(n181), .B(n17425), .Z(n17427) );
  XOR U18152 ( .A(b[3]), .B(a[130]), .Z(n17574) );
  NAND U18153 ( .A(n182), .B(n17574), .Z(n17426) );
  AND U18154 ( .A(n17427), .B(n17426), .Z(n17581) );
  NAND U18155 ( .A(n189), .B(n17428), .Z(n17430) );
  XOR U18156 ( .A(b[17]), .B(a[116]), .Z(n17577) );
  NAND U18157 ( .A(n37652), .B(n17577), .Z(n17429) );
  NAND U18158 ( .A(n17430), .B(n17429), .Z(n17580) );
  XNOR U18159 ( .A(n17581), .B(n17580), .Z(n17582) );
  XOR U18160 ( .A(n17583), .B(n17582), .Z(n17615) );
  XOR U18161 ( .A(n17614), .B(n17615), .Z(n17617) );
  XOR U18162 ( .A(n17616), .B(n17617), .Z(n17551) );
  NANDN U18163 ( .A(n17432), .B(n17431), .Z(n17436) );
  NANDN U18164 ( .A(n17434), .B(n17433), .Z(n17435) );
  AND U18165 ( .A(n17436), .B(n17435), .Z(n17604) );
  NANDN U18166 ( .A(n17438), .B(n17437), .Z(n17442) );
  NANDN U18167 ( .A(n17440), .B(n17439), .Z(n17441) );
  NAND U18168 ( .A(n17442), .B(n17441), .Z(n17605) );
  XNOR U18169 ( .A(n17604), .B(n17605), .Z(n17606) );
  NANDN U18170 ( .A(n17444), .B(n17443), .Z(n17448) );
  NANDN U18171 ( .A(n17446), .B(n17445), .Z(n17447) );
  NAND U18172 ( .A(n17448), .B(n17447), .Z(n17607) );
  XNOR U18173 ( .A(n17606), .B(n17607), .Z(n17550) );
  XNOR U18174 ( .A(n17551), .B(n17550), .Z(n17553) );
  NANDN U18175 ( .A(n17450), .B(n17449), .Z(n17454) );
  NANDN U18176 ( .A(n17452), .B(n17451), .Z(n17453) );
  AND U18177 ( .A(n17454), .B(n17453), .Z(n17552) );
  XOR U18178 ( .A(n17553), .B(n17552), .Z(n17665) );
  NANDN U18179 ( .A(n17456), .B(n17455), .Z(n17460) );
  NANDN U18180 ( .A(n17458), .B(n17457), .Z(n17459) );
  AND U18181 ( .A(n17460), .B(n17459), .Z(n17662) );
  NANDN U18182 ( .A(n17462), .B(n17461), .Z(n17466) );
  NANDN U18183 ( .A(n17464), .B(n17463), .Z(n17465) );
  AND U18184 ( .A(n17466), .B(n17465), .Z(n17547) );
  NANDN U18185 ( .A(n17468), .B(n17467), .Z(n17472) );
  OR U18186 ( .A(n17470), .B(n17469), .Z(n17471) );
  AND U18187 ( .A(n17472), .B(n17471), .Z(n17545) );
  NANDN U18188 ( .A(n17474), .B(n17473), .Z(n17478) );
  NANDN U18189 ( .A(n17476), .B(n17475), .Z(n17477) );
  AND U18190 ( .A(n17478), .B(n17477), .Z(n17611) );
  NANDN U18191 ( .A(n17480), .B(n17479), .Z(n17484) );
  NANDN U18192 ( .A(n17482), .B(n17481), .Z(n17483) );
  NAND U18193 ( .A(n17484), .B(n17483), .Z(n17610) );
  XNOR U18194 ( .A(n17611), .B(n17610), .Z(n17613) );
  NAND U18195 ( .A(n194), .B(n17485), .Z(n17487) );
  XOR U18196 ( .A(b[29]), .B(a[104]), .Z(n17635) );
  NAND U18197 ( .A(n38456), .B(n17635), .Z(n17486) );
  AND U18198 ( .A(n17487), .B(n17486), .Z(n17557) );
  AND U18199 ( .A(b[31]), .B(a[100]), .Z(n17556) );
  XNOR U18200 ( .A(n17557), .B(n17556), .Z(n17558) );
  NAND U18201 ( .A(b[0]), .B(a[132]), .Z(n17488) );
  XNOR U18202 ( .A(b[1]), .B(n17488), .Z(n17490) );
  NANDN U18203 ( .A(b[0]), .B(a[131]), .Z(n17489) );
  NAND U18204 ( .A(n17490), .B(n17489), .Z(n17559) );
  XNOR U18205 ( .A(n17558), .B(n17559), .Z(n17599) );
  NAND U18206 ( .A(n38185), .B(n17491), .Z(n17493) );
  XOR U18207 ( .A(b[23]), .B(a[110]), .Z(n17638) );
  NAND U18208 ( .A(n38132), .B(n17638), .Z(n17492) );
  AND U18209 ( .A(n17493), .B(n17492), .Z(n17628) );
  NAND U18210 ( .A(n184), .B(n17494), .Z(n17496) );
  XOR U18211 ( .A(b[7]), .B(a[126]), .Z(n17641) );
  NAND U18212 ( .A(n36592), .B(n17641), .Z(n17495) );
  AND U18213 ( .A(n17496), .B(n17495), .Z(n17627) );
  NAND U18214 ( .A(n38289), .B(n17497), .Z(n17499) );
  XOR U18215 ( .A(b[25]), .B(a[108]), .Z(n17644) );
  NAND U18216 ( .A(n38247), .B(n17644), .Z(n17498) );
  NAND U18217 ( .A(n17499), .B(n17498), .Z(n17626) );
  XOR U18218 ( .A(n17627), .B(n17626), .Z(n17629) );
  XOR U18219 ( .A(n17628), .B(n17629), .Z(n17598) );
  XOR U18220 ( .A(n17599), .B(n17598), .Z(n17601) );
  NAND U18221 ( .A(n187), .B(n17500), .Z(n17502) );
  XOR U18222 ( .A(b[13]), .B(a[120]), .Z(n17647) );
  NAND U18223 ( .A(n37295), .B(n17647), .Z(n17501) );
  AND U18224 ( .A(n17502), .B(n17501), .Z(n17593) );
  NAND U18225 ( .A(n186), .B(n17503), .Z(n17505) );
  XOR U18226 ( .A(b[11]), .B(a[122]), .Z(n17650) );
  NAND U18227 ( .A(n37097), .B(n17650), .Z(n17504) );
  NAND U18228 ( .A(n17505), .B(n17504), .Z(n17592) );
  XNOR U18229 ( .A(n17593), .B(n17592), .Z(n17595) );
  NAND U18230 ( .A(n188), .B(n17506), .Z(n17508) );
  XOR U18231 ( .A(b[15]), .B(a[118]), .Z(n17653) );
  NAND U18232 ( .A(n37382), .B(n17653), .Z(n17507) );
  AND U18233 ( .A(n17508), .B(n17507), .Z(n17589) );
  NAND U18234 ( .A(n38064), .B(n17509), .Z(n17511) );
  XOR U18235 ( .A(b[21]), .B(a[112]), .Z(n17656) );
  NAND U18236 ( .A(n37993), .B(n17656), .Z(n17510) );
  AND U18237 ( .A(n17511), .B(n17510), .Z(n17587) );
  NAND U18238 ( .A(n185), .B(n17512), .Z(n17514) );
  XOR U18239 ( .A(b[9]), .B(a[124]), .Z(n17659) );
  NAND U18240 ( .A(n36805), .B(n17659), .Z(n17513) );
  NAND U18241 ( .A(n17514), .B(n17513), .Z(n17586) );
  XNOR U18242 ( .A(n17587), .B(n17586), .Z(n17588) );
  XNOR U18243 ( .A(n17589), .B(n17588), .Z(n17594) );
  XOR U18244 ( .A(n17595), .B(n17594), .Z(n17600) );
  XNOR U18245 ( .A(n17601), .B(n17600), .Z(n17612) );
  XNOR U18246 ( .A(n17613), .B(n17612), .Z(n17544) );
  XNOR U18247 ( .A(n17545), .B(n17544), .Z(n17546) );
  XOR U18248 ( .A(n17547), .B(n17546), .Z(n17663) );
  XNOR U18249 ( .A(n17662), .B(n17663), .Z(n17664) );
  XNOR U18250 ( .A(n17665), .B(n17664), .Z(n17540) );
  XOR U18251 ( .A(n17541), .B(n17540), .Z(n17533) );
  NANDN U18252 ( .A(n17516), .B(n17515), .Z(n17520) );
  OR U18253 ( .A(n17518), .B(n17517), .Z(n17519) );
  AND U18254 ( .A(n17520), .B(n17519), .Z(n17532) );
  XNOR U18255 ( .A(n17533), .B(n17532), .Z(n17534) );
  XNOR U18256 ( .A(n17535), .B(n17534), .Z(n17526) );
  XNOR U18257 ( .A(n17527), .B(n17526), .Z(n17528) );
  XNOR U18258 ( .A(n17529), .B(n17528), .Z(n17668) );
  XNOR U18259 ( .A(sreg[356]), .B(n17668), .Z(n17670) );
  NANDN U18260 ( .A(sreg[355]), .B(n17521), .Z(n17525) );
  NAND U18261 ( .A(n17523), .B(n17522), .Z(n17524) );
  NAND U18262 ( .A(n17525), .B(n17524), .Z(n17669) );
  XNOR U18263 ( .A(n17670), .B(n17669), .Z(c[356]) );
  NANDN U18264 ( .A(n17527), .B(n17526), .Z(n17531) );
  NANDN U18265 ( .A(n17529), .B(n17528), .Z(n17530) );
  AND U18266 ( .A(n17531), .B(n17530), .Z(n17676) );
  NANDN U18267 ( .A(n17533), .B(n17532), .Z(n17537) );
  NANDN U18268 ( .A(n17535), .B(n17534), .Z(n17536) );
  AND U18269 ( .A(n17537), .B(n17536), .Z(n17674) );
  NANDN U18270 ( .A(n17539), .B(n17538), .Z(n17543) );
  NAND U18271 ( .A(n17541), .B(n17540), .Z(n17542) );
  AND U18272 ( .A(n17543), .B(n17542), .Z(n17681) );
  NANDN U18273 ( .A(n17545), .B(n17544), .Z(n17549) );
  NANDN U18274 ( .A(n17547), .B(n17546), .Z(n17548) );
  AND U18275 ( .A(n17549), .B(n17548), .Z(n17810) );
  NANDN U18276 ( .A(n17551), .B(n17550), .Z(n17555) );
  NAND U18277 ( .A(n17553), .B(n17552), .Z(n17554) );
  AND U18278 ( .A(n17555), .B(n17554), .Z(n17809) );
  XNOR U18279 ( .A(n17810), .B(n17809), .Z(n17812) );
  NANDN U18280 ( .A(n17557), .B(n17556), .Z(n17561) );
  NANDN U18281 ( .A(n17559), .B(n17558), .Z(n17560) );
  AND U18282 ( .A(n17561), .B(n17560), .Z(n17745) );
  NAND U18283 ( .A(n38385), .B(n17562), .Z(n17564) );
  XOR U18284 ( .A(b[27]), .B(a[107]), .Z(n17691) );
  NAND U18285 ( .A(n38343), .B(n17691), .Z(n17563) );
  AND U18286 ( .A(n17564), .B(n17563), .Z(n17752) );
  NAND U18287 ( .A(n183), .B(n17565), .Z(n17567) );
  XOR U18288 ( .A(b[5]), .B(a[129]), .Z(n17694) );
  NAND U18289 ( .A(n36296), .B(n17694), .Z(n17566) );
  AND U18290 ( .A(n17567), .B(n17566), .Z(n17750) );
  NAND U18291 ( .A(n190), .B(n17568), .Z(n17570) );
  XOR U18292 ( .A(b[19]), .B(a[115]), .Z(n17697) );
  NAND U18293 ( .A(n37821), .B(n17697), .Z(n17569) );
  NAND U18294 ( .A(n17570), .B(n17569), .Z(n17749) );
  XNOR U18295 ( .A(n17750), .B(n17749), .Z(n17751) );
  XNOR U18296 ( .A(n17752), .B(n17751), .Z(n17743) );
  NAND U18297 ( .A(n38470), .B(n17571), .Z(n17573) );
  XOR U18298 ( .A(b[31]), .B(a[103]), .Z(n17700) );
  NAND U18299 ( .A(n38453), .B(n17700), .Z(n17572) );
  AND U18300 ( .A(n17573), .B(n17572), .Z(n17712) );
  NAND U18301 ( .A(n181), .B(n17574), .Z(n17576) );
  XOR U18302 ( .A(b[3]), .B(a[131]), .Z(n17703) );
  NAND U18303 ( .A(n182), .B(n17703), .Z(n17575) );
  AND U18304 ( .A(n17576), .B(n17575), .Z(n17710) );
  NAND U18305 ( .A(n189), .B(n17577), .Z(n17579) );
  XOR U18306 ( .A(b[17]), .B(a[117]), .Z(n17706) );
  NAND U18307 ( .A(n37652), .B(n17706), .Z(n17578) );
  NAND U18308 ( .A(n17579), .B(n17578), .Z(n17709) );
  XNOR U18309 ( .A(n17710), .B(n17709), .Z(n17711) );
  XOR U18310 ( .A(n17712), .B(n17711), .Z(n17744) );
  XOR U18311 ( .A(n17743), .B(n17744), .Z(n17746) );
  XOR U18312 ( .A(n17745), .B(n17746), .Z(n17792) );
  NANDN U18313 ( .A(n17581), .B(n17580), .Z(n17585) );
  NANDN U18314 ( .A(n17583), .B(n17582), .Z(n17584) );
  AND U18315 ( .A(n17585), .B(n17584), .Z(n17733) );
  NANDN U18316 ( .A(n17587), .B(n17586), .Z(n17591) );
  NANDN U18317 ( .A(n17589), .B(n17588), .Z(n17590) );
  NAND U18318 ( .A(n17591), .B(n17590), .Z(n17734) );
  XNOR U18319 ( .A(n17733), .B(n17734), .Z(n17735) );
  NANDN U18320 ( .A(n17593), .B(n17592), .Z(n17597) );
  NAND U18321 ( .A(n17595), .B(n17594), .Z(n17596) );
  NAND U18322 ( .A(n17597), .B(n17596), .Z(n17736) );
  XNOR U18323 ( .A(n17735), .B(n17736), .Z(n17791) );
  XNOR U18324 ( .A(n17792), .B(n17791), .Z(n17794) );
  NAND U18325 ( .A(n17599), .B(n17598), .Z(n17603) );
  NAND U18326 ( .A(n17601), .B(n17600), .Z(n17602) );
  AND U18327 ( .A(n17603), .B(n17602), .Z(n17793) );
  XOR U18328 ( .A(n17794), .B(n17793), .Z(n17806) );
  NANDN U18329 ( .A(n17605), .B(n17604), .Z(n17609) );
  NANDN U18330 ( .A(n17607), .B(n17606), .Z(n17608) );
  AND U18331 ( .A(n17609), .B(n17608), .Z(n17803) );
  NANDN U18332 ( .A(n17615), .B(n17614), .Z(n17619) );
  OR U18333 ( .A(n17617), .B(n17616), .Z(n17618) );
  AND U18334 ( .A(n17619), .B(n17618), .Z(n17798) );
  NANDN U18335 ( .A(n17621), .B(n17620), .Z(n17625) );
  NANDN U18336 ( .A(n17623), .B(n17622), .Z(n17624) );
  AND U18337 ( .A(n17625), .B(n17624), .Z(n17740) );
  NANDN U18338 ( .A(n17627), .B(n17626), .Z(n17631) );
  OR U18339 ( .A(n17629), .B(n17628), .Z(n17630) );
  NAND U18340 ( .A(n17631), .B(n17630), .Z(n17739) );
  XNOR U18341 ( .A(n17740), .B(n17739), .Z(n17742) );
  NAND U18342 ( .A(b[0]), .B(a[133]), .Z(n17632) );
  XNOR U18343 ( .A(b[1]), .B(n17632), .Z(n17634) );
  NANDN U18344 ( .A(b[0]), .B(a[132]), .Z(n17633) );
  NAND U18345 ( .A(n17634), .B(n17633), .Z(n17688) );
  NAND U18346 ( .A(n194), .B(n17635), .Z(n17637) );
  XOR U18347 ( .A(b[29]), .B(a[105]), .Z(n17764) );
  NAND U18348 ( .A(n38456), .B(n17764), .Z(n17636) );
  AND U18349 ( .A(n17637), .B(n17636), .Z(n17686) );
  AND U18350 ( .A(b[31]), .B(a[101]), .Z(n17685) );
  XNOR U18351 ( .A(n17686), .B(n17685), .Z(n17687) );
  XNOR U18352 ( .A(n17688), .B(n17687), .Z(n17728) );
  NAND U18353 ( .A(n38185), .B(n17638), .Z(n17640) );
  XOR U18354 ( .A(b[23]), .B(a[111]), .Z(n17767) );
  NAND U18355 ( .A(n38132), .B(n17767), .Z(n17639) );
  AND U18356 ( .A(n17640), .B(n17639), .Z(n17757) );
  NAND U18357 ( .A(n184), .B(n17641), .Z(n17643) );
  XOR U18358 ( .A(b[7]), .B(a[127]), .Z(n17770) );
  NAND U18359 ( .A(n36592), .B(n17770), .Z(n17642) );
  AND U18360 ( .A(n17643), .B(n17642), .Z(n17756) );
  NAND U18361 ( .A(n38289), .B(n17644), .Z(n17646) );
  XOR U18362 ( .A(b[25]), .B(a[109]), .Z(n17773) );
  NAND U18363 ( .A(n38247), .B(n17773), .Z(n17645) );
  NAND U18364 ( .A(n17646), .B(n17645), .Z(n17755) );
  XOR U18365 ( .A(n17756), .B(n17755), .Z(n17758) );
  XOR U18366 ( .A(n17757), .B(n17758), .Z(n17727) );
  XOR U18367 ( .A(n17728), .B(n17727), .Z(n17730) );
  NAND U18368 ( .A(n187), .B(n17647), .Z(n17649) );
  XOR U18369 ( .A(b[13]), .B(a[121]), .Z(n17776) );
  NAND U18370 ( .A(n37295), .B(n17776), .Z(n17648) );
  AND U18371 ( .A(n17649), .B(n17648), .Z(n17722) );
  NAND U18372 ( .A(n186), .B(n17650), .Z(n17652) );
  XOR U18373 ( .A(b[11]), .B(a[123]), .Z(n17779) );
  NAND U18374 ( .A(n37097), .B(n17779), .Z(n17651) );
  NAND U18375 ( .A(n17652), .B(n17651), .Z(n17721) );
  XNOR U18376 ( .A(n17722), .B(n17721), .Z(n17724) );
  NAND U18377 ( .A(n188), .B(n17653), .Z(n17655) );
  XOR U18378 ( .A(b[15]), .B(a[119]), .Z(n17782) );
  NAND U18379 ( .A(n37382), .B(n17782), .Z(n17654) );
  AND U18380 ( .A(n17655), .B(n17654), .Z(n17718) );
  NAND U18381 ( .A(n38064), .B(n17656), .Z(n17658) );
  XOR U18382 ( .A(b[21]), .B(a[113]), .Z(n17785) );
  NAND U18383 ( .A(n37993), .B(n17785), .Z(n17657) );
  AND U18384 ( .A(n17658), .B(n17657), .Z(n17716) );
  NAND U18385 ( .A(n185), .B(n17659), .Z(n17661) );
  XOR U18386 ( .A(b[9]), .B(a[125]), .Z(n17788) );
  NAND U18387 ( .A(n36805), .B(n17788), .Z(n17660) );
  NAND U18388 ( .A(n17661), .B(n17660), .Z(n17715) );
  XNOR U18389 ( .A(n17716), .B(n17715), .Z(n17717) );
  XNOR U18390 ( .A(n17718), .B(n17717), .Z(n17723) );
  XOR U18391 ( .A(n17724), .B(n17723), .Z(n17729) );
  XNOR U18392 ( .A(n17730), .B(n17729), .Z(n17741) );
  XNOR U18393 ( .A(n17742), .B(n17741), .Z(n17797) );
  XNOR U18394 ( .A(n17798), .B(n17797), .Z(n17799) );
  XOR U18395 ( .A(n17800), .B(n17799), .Z(n17804) );
  XNOR U18396 ( .A(n17803), .B(n17804), .Z(n17805) );
  XNOR U18397 ( .A(n17806), .B(n17805), .Z(n17811) );
  XOR U18398 ( .A(n17812), .B(n17811), .Z(n17680) );
  NANDN U18399 ( .A(n17663), .B(n17662), .Z(n17667) );
  NANDN U18400 ( .A(n17665), .B(n17664), .Z(n17666) );
  AND U18401 ( .A(n17667), .B(n17666), .Z(n17679) );
  XOR U18402 ( .A(n17680), .B(n17679), .Z(n17682) );
  XNOR U18403 ( .A(n17681), .B(n17682), .Z(n17673) );
  XNOR U18404 ( .A(n17674), .B(n17673), .Z(n17675) );
  XNOR U18405 ( .A(n17676), .B(n17675), .Z(n17815) );
  XNOR U18406 ( .A(sreg[357]), .B(n17815), .Z(n17817) );
  NANDN U18407 ( .A(sreg[356]), .B(n17668), .Z(n17672) );
  NAND U18408 ( .A(n17670), .B(n17669), .Z(n17671) );
  NAND U18409 ( .A(n17672), .B(n17671), .Z(n17816) );
  XNOR U18410 ( .A(n17817), .B(n17816), .Z(c[357]) );
  NANDN U18411 ( .A(n17674), .B(n17673), .Z(n17678) );
  NANDN U18412 ( .A(n17676), .B(n17675), .Z(n17677) );
  AND U18413 ( .A(n17678), .B(n17677), .Z(n17823) );
  NANDN U18414 ( .A(n17680), .B(n17679), .Z(n17684) );
  NANDN U18415 ( .A(n17682), .B(n17681), .Z(n17683) );
  AND U18416 ( .A(n17684), .B(n17683), .Z(n17821) );
  NANDN U18417 ( .A(n17686), .B(n17685), .Z(n17690) );
  NANDN U18418 ( .A(n17688), .B(n17687), .Z(n17689) );
  AND U18419 ( .A(n17690), .B(n17689), .Z(n17900) );
  NAND U18420 ( .A(n38385), .B(n17691), .Z(n17693) );
  XOR U18421 ( .A(b[27]), .B(a[108]), .Z(n17844) );
  NAND U18422 ( .A(n38343), .B(n17844), .Z(n17692) );
  AND U18423 ( .A(n17693), .B(n17692), .Z(n17907) );
  NAND U18424 ( .A(n183), .B(n17694), .Z(n17696) );
  XOR U18425 ( .A(b[5]), .B(a[130]), .Z(n17847) );
  NAND U18426 ( .A(n36296), .B(n17847), .Z(n17695) );
  AND U18427 ( .A(n17696), .B(n17695), .Z(n17905) );
  NAND U18428 ( .A(n190), .B(n17697), .Z(n17699) );
  XOR U18429 ( .A(b[19]), .B(a[116]), .Z(n17850) );
  NAND U18430 ( .A(n37821), .B(n17850), .Z(n17698) );
  NAND U18431 ( .A(n17699), .B(n17698), .Z(n17904) );
  XNOR U18432 ( .A(n17905), .B(n17904), .Z(n17906) );
  XNOR U18433 ( .A(n17907), .B(n17906), .Z(n17898) );
  NAND U18434 ( .A(n38470), .B(n17700), .Z(n17702) );
  XOR U18435 ( .A(b[31]), .B(a[104]), .Z(n17853) );
  NAND U18436 ( .A(n38453), .B(n17853), .Z(n17701) );
  AND U18437 ( .A(n17702), .B(n17701), .Z(n17865) );
  NAND U18438 ( .A(n181), .B(n17703), .Z(n17705) );
  XOR U18439 ( .A(b[3]), .B(a[132]), .Z(n17856) );
  NAND U18440 ( .A(n182), .B(n17856), .Z(n17704) );
  AND U18441 ( .A(n17705), .B(n17704), .Z(n17863) );
  NAND U18442 ( .A(n189), .B(n17706), .Z(n17708) );
  XOR U18443 ( .A(b[17]), .B(a[118]), .Z(n17859) );
  NAND U18444 ( .A(n37652), .B(n17859), .Z(n17707) );
  NAND U18445 ( .A(n17708), .B(n17707), .Z(n17862) );
  XNOR U18446 ( .A(n17863), .B(n17862), .Z(n17864) );
  XOR U18447 ( .A(n17865), .B(n17864), .Z(n17899) );
  XOR U18448 ( .A(n17898), .B(n17899), .Z(n17901) );
  XOR U18449 ( .A(n17900), .B(n17901), .Z(n17947) );
  NANDN U18450 ( .A(n17710), .B(n17709), .Z(n17714) );
  NANDN U18451 ( .A(n17712), .B(n17711), .Z(n17713) );
  AND U18452 ( .A(n17714), .B(n17713), .Z(n17886) );
  NANDN U18453 ( .A(n17716), .B(n17715), .Z(n17720) );
  NANDN U18454 ( .A(n17718), .B(n17717), .Z(n17719) );
  NAND U18455 ( .A(n17720), .B(n17719), .Z(n17887) );
  XNOR U18456 ( .A(n17886), .B(n17887), .Z(n17888) );
  NANDN U18457 ( .A(n17722), .B(n17721), .Z(n17726) );
  NAND U18458 ( .A(n17724), .B(n17723), .Z(n17725) );
  NAND U18459 ( .A(n17726), .B(n17725), .Z(n17889) );
  XNOR U18460 ( .A(n17888), .B(n17889), .Z(n17946) );
  XNOR U18461 ( .A(n17947), .B(n17946), .Z(n17949) );
  NAND U18462 ( .A(n17728), .B(n17727), .Z(n17732) );
  NAND U18463 ( .A(n17730), .B(n17729), .Z(n17731) );
  AND U18464 ( .A(n17732), .B(n17731), .Z(n17948) );
  XOR U18465 ( .A(n17949), .B(n17948), .Z(n17960) );
  NANDN U18466 ( .A(n17734), .B(n17733), .Z(n17738) );
  NANDN U18467 ( .A(n17736), .B(n17735), .Z(n17737) );
  AND U18468 ( .A(n17738), .B(n17737), .Z(n17958) );
  NANDN U18469 ( .A(n17744), .B(n17743), .Z(n17748) );
  OR U18470 ( .A(n17746), .B(n17745), .Z(n17747) );
  AND U18471 ( .A(n17748), .B(n17747), .Z(n17953) );
  NANDN U18472 ( .A(n17750), .B(n17749), .Z(n17754) );
  NANDN U18473 ( .A(n17752), .B(n17751), .Z(n17753) );
  AND U18474 ( .A(n17754), .B(n17753), .Z(n17893) );
  NANDN U18475 ( .A(n17756), .B(n17755), .Z(n17760) );
  OR U18476 ( .A(n17758), .B(n17757), .Z(n17759) );
  NAND U18477 ( .A(n17760), .B(n17759), .Z(n17892) );
  XNOR U18478 ( .A(n17893), .B(n17892), .Z(n17894) );
  NAND U18479 ( .A(b[0]), .B(a[134]), .Z(n17761) );
  XNOR U18480 ( .A(b[1]), .B(n17761), .Z(n17763) );
  NANDN U18481 ( .A(b[0]), .B(a[133]), .Z(n17762) );
  NAND U18482 ( .A(n17763), .B(n17762), .Z(n17841) );
  NAND U18483 ( .A(n194), .B(n17764), .Z(n17766) );
  XOR U18484 ( .A(b[29]), .B(a[106]), .Z(n17919) );
  NAND U18485 ( .A(n38456), .B(n17919), .Z(n17765) );
  AND U18486 ( .A(n17766), .B(n17765), .Z(n17839) );
  AND U18487 ( .A(b[31]), .B(a[102]), .Z(n17838) );
  XNOR U18488 ( .A(n17839), .B(n17838), .Z(n17840) );
  XNOR U18489 ( .A(n17841), .B(n17840), .Z(n17880) );
  NAND U18490 ( .A(n38185), .B(n17767), .Z(n17769) );
  XOR U18491 ( .A(b[23]), .B(a[112]), .Z(n17922) );
  NAND U18492 ( .A(n38132), .B(n17922), .Z(n17768) );
  AND U18493 ( .A(n17769), .B(n17768), .Z(n17913) );
  NAND U18494 ( .A(n184), .B(n17770), .Z(n17772) );
  XOR U18495 ( .A(b[7]), .B(a[128]), .Z(n17925) );
  NAND U18496 ( .A(n36592), .B(n17925), .Z(n17771) );
  AND U18497 ( .A(n17772), .B(n17771), .Z(n17911) );
  NAND U18498 ( .A(n38289), .B(n17773), .Z(n17775) );
  XOR U18499 ( .A(b[25]), .B(a[110]), .Z(n17928) );
  NAND U18500 ( .A(n38247), .B(n17928), .Z(n17774) );
  NAND U18501 ( .A(n17775), .B(n17774), .Z(n17910) );
  XNOR U18502 ( .A(n17911), .B(n17910), .Z(n17912) );
  XOR U18503 ( .A(n17913), .B(n17912), .Z(n17881) );
  XNOR U18504 ( .A(n17880), .B(n17881), .Z(n17882) );
  NAND U18505 ( .A(n187), .B(n17776), .Z(n17778) );
  XOR U18506 ( .A(b[13]), .B(a[122]), .Z(n17931) );
  NAND U18507 ( .A(n37295), .B(n17931), .Z(n17777) );
  AND U18508 ( .A(n17778), .B(n17777), .Z(n17875) );
  NAND U18509 ( .A(n186), .B(n17779), .Z(n17781) );
  XOR U18510 ( .A(b[11]), .B(a[124]), .Z(n17934) );
  NAND U18511 ( .A(n37097), .B(n17934), .Z(n17780) );
  NAND U18512 ( .A(n17781), .B(n17780), .Z(n17874) );
  XNOR U18513 ( .A(n17875), .B(n17874), .Z(n17876) );
  NAND U18514 ( .A(n188), .B(n17782), .Z(n17784) );
  XOR U18515 ( .A(b[15]), .B(a[120]), .Z(n17937) );
  NAND U18516 ( .A(n37382), .B(n17937), .Z(n17783) );
  AND U18517 ( .A(n17784), .B(n17783), .Z(n17871) );
  NAND U18518 ( .A(n38064), .B(n17785), .Z(n17787) );
  XOR U18519 ( .A(b[21]), .B(a[114]), .Z(n17940) );
  NAND U18520 ( .A(n37993), .B(n17940), .Z(n17786) );
  AND U18521 ( .A(n17787), .B(n17786), .Z(n17869) );
  NAND U18522 ( .A(n185), .B(n17788), .Z(n17790) );
  XOR U18523 ( .A(b[9]), .B(a[126]), .Z(n17943) );
  NAND U18524 ( .A(n36805), .B(n17943), .Z(n17789) );
  NAND U18525 ( .A(n17790), .B(n17789), .Z(n17868) );
  XNOR U18526 ( .A(n17869), .B(n17868), .Z(n17870) );
  XOR U18527 ( .A(n17871), .B(n17870), .Z(n17877) );
  XOR U18528 ( .A(n17876), .B(n17877), .Z(n17883) );
  XOR U18529 ( .A(n17882), .B(n17883), .Z(n17895) );
  XNOR U18530 ( .A(n17894), .B(n17895), .Z(n17952) );
  XNOR U18531 ( .A(n17953), .B(n17952), .Z(n17954) );
  XOR U18532 ( .A(n17955), .B(n17954), .Z(n17959) );
  XOR U18533 ( .A(n17958), .B(n17959), .Z(n17961) );
  XOR U18534 ( .A(n17960), .B(n17961), .Z(n17835) );
  NANDN U18535 ( .A(n17792), .B(n17791), .Z(n17796) );
  NAND U18536 ( .A(n17794), .B(n17793), .Z(n17795) );
  AND U18537 ( .A(n17796), .B(n17795), .Z(n17833) );
  NANDN U18538 ( .A(n17798), .B(n17797), .Z(n17802) );
  NANDN U18539 ( .A(n17800), .B(n17799), .Z(n17801) );
  AND U18540 ( .A(n17802), .B(n17801), .Z(n17832) );
  XNOR U18541 ( .A(n17833), .B(n17832), .Z(n17834) );
  XNOR U18542 ( .A(n17835), .B(n17834), .Z(n17826) );
  NANDN U18543 ( .A(n17804), .B(n17803), .Z(n17808) );
  NANDN U18544 ( .A(n17806), .B(n17805), .Z(n17807) );
  NAND U18545 ( .A(n17808), .B(n17807), .Z(n17827) );
  XNOR U18546 ( .A(n17826), .B(n17827), .Z(n17828) );
  NANDN U18547 ( .A(n17810), .B(n17809), .Z(n17814) );
  NAND U18548 ( .A(n17812), .B(n17811), .Z(n17813) );
  NAND U18549 ( .A(n17814), .B(n17813), .Z(n17829) );
  XNOR U18550 ( .A(n17828), .B(n17829), .Z(n17820) );
  XNOR U18551 ( .A(n17821), .B(n17820), .Z(n17822) );
  XNOR U18552 ( .A(n17823), .B(n17822), .Z(n17964) );
  XNOR U18553 ( .A(sreg[358]), .B(n17964), .Z(n17966) );
  NANDN U18554 ( .A(sreg[357]), .B(n17815), .Z(n17819) );
  NAND U18555 ( .A(n17817), .B(n17816), .Z(n17818) );
  NAND U18556 ( .A(n17819), .B(n17818), .Z(n17965) );
  XNOR U18557 ( .A(n17966), .B(n17965), .Z(c[358]) );
  NANDN U18558 ( .A(n17821), .B(n17820), .Z(n17825) );
  NANDN U18559 ( .A(n17823), .B(n17822), .Z(n17824) );
  AND U18560 ( .A(n17825), .B(n17824), .Z(n17972) );
  NANDN U18561 ( .A(n17827), .B(n17826), .Z(n17831) );
  NANDN U18562 ( .A(n17829), .B(n17828), .Z(n17830) );
  AND U18563 ( .A(n17831), .B(n17830), .Z(n17970) );
  NANDN U18564 ( .A(n17833), .B(n17832), .Z(n17837) );
  NANDN U18565 ( .A(n17835), .B(n17834), .Z(n17836) );
  AND U18566 ( .A(n17837), .B(n17836), .Z(n17978) );
  NANDN U18567 ( .A(n17839), .B(n17838), .Z(n17843) );
  NANDN U18568 ( .A(n17841), .B(n17840), .Z(n17842) );
  AND U18569 ( .A(n17843), .B(n17842), .Z(n18061) );
  NAND U18570 ( .A(n38385), .B(n17844), .Z(n17846) );
  XOR U18571 ( .A(b[27]), .B(a[109]), .Z(n18005) );
  NAND U18572 ( .A(n38343), .B(n18005), .Z(n17845) );
  AND U18573 ( .A(n17846), .B(n17845), .Z(n18068) );
  NAND U18574 ( .A(n183), .B(n17847), .Z(n17849) );
  XOR U18575 ( .A(b[5]), .B(a[131]), .Z(n18008) );
  NAND U18576 ( .A(n36296), .B(n18008), .Z(n17848) );
  AND U18577 ( .A(n17849), .B(n17848), .Z(n18066) );
  NAND U18578 ( .A(n190), .B(n17850), .Z(n17852) );
  XOR U18579 ( .A(b[19]), .B(a[117]), .Z(n18011) );
  NAND U18580 ( .A(n37821), .B(n18011), .Z(n17851) );
  NAND U18581 ( .A(n17852), .B(n17851), .Z(n18065) );
  XNOR U18582 ( .A(n18066), .B(n18065), .Z(n18067) );
  XNOR U18583 ( .A(n18068), .B(n18067), .Z(n18059) );
  NAND U18584 ( .A(n38470), .B(n17853), .Z(n17855) );
  XOR U18585 ( .A(b[31]), .B(a[105]), .Z(n18014) );
  NAND U18586 ( .A(n38453), .B(n18014), .Z(n17854) );
  AND U18587 ( .A(n17855), .B(n17854), .Z(n18026) );
  NAND U18588 ( .A(n181), .B(n17856), .Z(n17858) );
  XOR U18589 ( .A(b[3]), .B(a[133]), .Z(n18017) );
  NAND U18590 ( .A(n182), .B(n18017), .Z(n17857) );
  AND U18591 ( .A(n17858), .B(n17857), .Z(n18024) );
  NAND U18592 ( .A(n189), .B(n17859), .Z(n17861) );
  XOR U18593 ( .A(b[17]), .B(a[119]), .Z(n18020) );
  NAND U18594 ( .A(n37652), .B(n18020), .Z(n17860) );
  NAND U18595 ( .A(n17861), .B(n17860), .Z(n18023) );
  XNOR U18596 ( .A(n18024), .B(n18023), .Z(n18025) );
  XOR U18597 ( .A(n18026), .B(n18025), .Z(n18060) );
  XOR U18598 ( .A(n18059), .B(n18060), .Z(n18062) );
  XOR U18599 ( .A(n18061), .B(n18062), .Z(n17994) );
  NANDN U18600 ( .A(n17863), .B(n17862), .Z(n17867) );
  NANDN U18601 ( .A(n17865), .B(n17864), .Z(n17866) );
  AND U18602 ( .A(n17867), .B(n17866), .Z(n18047) );
  NANDN U18603 ( .A(n17869), .B(n17868), .Z(n17873) );
  NANDN U18604 ( .A(n17871), .B(n17870), .Z(n17872) );
  NAND U18605 ( .A(n17873), .B(n17872), .Z(n18048) );
  XNOR U18606 ( .A(n18047), .B(n18048), .Z(n18049) );
  NANDN U18607 ( .A(n17875), .B(n17874), .Z(n17879) );
  NANDN U18608 ( .A(n17877), .B(n17876), .Z(n17878) );
  NAND U18609 ( .A(n17879), .B(n17878), .Z(n18050) );
  XNOR U18610 ( .A(n18049), .B(n18050), .Z(n17993) );
  XNOR U18611 ( .A(n17994), .B(n17993), .Z(n17996) );
  NANDN U18612 ( .A(n17881), .B(n17880), .Z(n17885) );
  NANDN U18613 ( .A(n17883), .B(n17882), .Z(n17884) );
  AND U18614 ( .A(n17885), .B(n17884), .Z(n17995) );
  XOR U18615 ( .A(n17996), .B(n17995), .Z(n18109) );
  NANDN U18616 ( .A(n17887), .B(n17886), .Z(n17891) );
  NANDN U18617 ( .A(n17889), .B(n17888), .Z(n17890) );
  AND U18618 ( .A(n17891), .B(n17890), .Z(n18107) );
  NANDN U18619 ( .A(n17893), .B(n17892), .Z(n17897) );
  NANDN U18620 ( .A(n17895), .B(n17894), .Z(n17896) );
  AND U18621 ( .A(n17897), .B(n17896), .Z(n17990) );
  NANDN U18622 ( .A(n17899), .B(n17898), .Z(n17903) );
  OR U18623 ( .A(n17901), .B(n17900), .Z(n17902) );
  AND U18624 ( .A(n17903), .B(n17902), .Z(n17988) );
  NANDN U18625 ( .A(n17905), .B(n17904), .Z(n17909) );
  NANDN U18626 ( .A(n17907), .B(n17906), .Z(n17908) );
  AND U18627 ( .A(n17909), .B(n17908), .Z(n18054) );
  NANDN U18628 ( .A(n17911), .B(n17910), .Z(n17915) );
  NANDN U18629 ( .A(n17913), .B(n17912), .Z(n17914) );
  NAND U18630 ( .A(n17915), .B(n17914), .Z(n18053) );
  XNOR U18631 ( .A(n18054), .B(n18053), .Z(n18055) );
  NAND U18632 ( .A(b[0]), .B(a[135]), .Z(n17916) );
  XNOR U18633 ( .A(b[1]), .B(n17916), .Z(n17918) );
  NANDN U18634 ( .A(b[0]), .B(a[134]), .Z(n17917) );
  NAND U18635 ( .A(n17918), .B(n17917), .Z(n18002) );
  NAND U18636 ( .A(n194), .B(n17919), .Z(n17921) );
  XOR U18637 ( .A(b[29]), .B(a[107]), .Z(n18077) );
  NAND U18638 ( .A(n38456), .B(n18077), .Z(n17920) );
  AND U18639 ( .A(n17921), .B(n17920), .Z(n18000) );
  AND U18640 ( .A(b[31]), .B(a[103]), .Z(n17999) );
  XNOR U18641 ( .A(n18000), .B(n17999), .Z(n18001) );
  XNOR U18642 ( .A(n18002), .B(n18001), .Z(n18041) );
  NAND U18643 ( .A(n38185), .B(n17922), .Z(n17924) );
  XOR U18644 ( .A(b[23]), .B(a[113]), .Z(n18083) );
  NAND U18645 ( .A(n38132), .B(n18083), .Z(n17923) );
  AND U18646 ( .A(n17924), .B(n17923), .Z(n18074) );
  NAND U18647 ( .A(n184), .B(n17925), .Z(n17927) );
  XOR U18648 ( .A(b[7]), .B(a[129]), .Z(n18086) );
  NAND U18649 ( .A(n36592), .B(n18086), .Z(n17926) );
  AND U18650 ( .A(n17927), .B(n17926), .Z(n18072) );
  NAND U18651 ( .A(n38289), .B(n17928), .Z(n17930) );
  XOR U18652 ( .A(b[25]), .B(a[111]), .Z(n18089) );
  NAND U18653 ( .A(n38247), .B(n18089), .Z(n17929) );
  NAND U18654 ( .A(n17930), .B(n17929), .Z(n18071) );
  XNOR U18655 ( .A(n18072), .B(n18071), .Z(n18073) );
  XOR U18656 ( .A(n18074), .B(n18073), .Z(n18042) );
  XNOR U18657 ( .A(n18041), .B(n18042), .Z(n18043) );
  NAND U18658 ( .A(n187), .B(n17931), .Z(n17933) );
  XOR U18659 ( .A(b[13]), .B(a[123]), .Z(n18092) );
  NAND U18660 ( .A(n37295), .B(n18092), .Z(n17932) );
  AND U18661 ( .A(n17933), .B(n17932), .Z(n18036) );
  NAND U18662 ( .A(n186), .B(n17934), .Z(n17936) );
  XOR U18663 ( .A(b[11]), .B(a[125]), .Z(n18095) );
  NAND U18664 ( .A(n37097), .B(n18095), .Z(n17935) );
  NAND U18665 ( .A(n17936), .B(n17935), .Z(n18035) );
  XNOR U18666 ( .A(n18036), .B(n18035), .Z(n18037) );
  NAND U18667 ( .A(n188), .B(n17937), .Z(n17939) );
  XOR U18668 ( .A(b[15]), .B(a[121]), .Z(n18098) );
  NAND U18669 ( .A(n37382), .B(n18098), .Z(n17938) );
  AND U18670 ( .A(n17939), .B(n17938), .Z(n18032) );
  NAND U18671 ( .A(n38064), .B(n17940), .Z(n17942) );
  XOR U18672 ( .A(b[21]), .B(a[115]), .Z(n18101) );
  NAND U18673 ( .A(n37993), .B(n18101), .Z(n17941) );
  AND U18674 ( .A(n17942), .B(n17941), .Z(n18030) );
  NAND U18675 ( .A(n185), .B(n17943), .Z(n17945) );
  XOR U18676 ( .A(b[9]), .B(a[127]), .Z(n18104) );
  NAND U18677 ( .A(n36805), .B(n18104), .Z(n17944) );
  NAND U18678 ( .A(n17945), .B(n17944), .Z(n18029) );
  XNOR U18679 ( .A(n18030), .B(n18029), .Z(n18031) );
  XOR U18680 ( .A(n18032), .B(n18031), .Z(n18038) );
  XOR U18681 ( .A(n18037), .B(n18038), .Z(n18044) );
  XOR U18682 ( .A(n18043), .B(n18044), .Z(n18056) );
  XNOR U18683 ( .A(n18055), .B(n18056), .Z(n17987) );
  XNOR U18684 ( .A(n17988), .B(n17987), .Z(n17989) );
  XOR U18685 ( .A(n17990), .B(n17989), .Z(n18108) );
  XOR U18686 ( .A(n18107), .B(n18108), .Z(n18110) );
  XOR U18687 ( .A(n18109), .B(n18110), .Z(n17984) );
  NANDN U18688 ( .A(n17947), .B(n17946), .Z(n17951) );
  NAND U18689 ( .A(n17949), .B(n17948), .Z(n17950) );
  AND U18690 ( .A(n17951), .B(n17950), .Z(n17982) );
  NANDN U18691 ( .A(n17953), .B(n17952), .Z(n17957) );
  NANDN U18692 ( .A(n17955), .B(n17954), .Z(n17956) );
  AND U18693 ( .A(n17957), .B(n17956), .Z(n17981) );
  XNOR U18694 ( .A(n17982), .B(n17981), .Z(n17983) );
  XNOR U18695 ( .A(n17984), .B(n17983), .Z(n17975) );
  NANDN U18696 ( .A(n17959), .B(n17958), .Z(n17963) );
  OR U18697 ( .A(n17961), .B(n17960), .Z(n17962) );
  NAND U18698 ( .A(n17963), .B(n17962), .Z(n17976) );
  XNOR U18699 ( .A(n17975), .B(n17976), .Z(n17977) );
  XNOR U18700 ( .A(n17978), .B(n17977), .Z(n17969) );
  XNOR U18701 ( .A(n17970), .B(n17969), .Z(n17971) );
  XNOR U18702 ( .A(n17972), .B(n17971), .Z(n18113) );
  XNOR U18703 ( .A(sreg[359]), .B(n18113), .Z(n18115) );
  NANDN U18704 ( .A(sreg[358]), .B(n17964), .Z(n17968) );
  NAND U18705 ( .A(n17966), .B(n17965), .Z(n17967) );
  NAND U18706 ( .A(n17968), .B(n17967), .Z(n18114) );
  XNOR U18707 ( .A(n18115), .B(n18114), .Z(c[359]) );
  NANDN U18708 ( .A(n17970), .B(n17969), .Z(n17974) );
  NANDN U18709 ( .A(n17972), .B(n17971), .Z(n17973) );
  AND U18710 ( .A(n17974), .B(n17973), .Z(n18121) );
  NANDN U18711 ( .A(n17976), .B(n17975), .Z(n17980) );
  NANDN U18712 ( .A(n17978), .B(n17977), .Z(n17979) );
  AND U18713 ( .A(n17980), .B(n17979), .Z(n18119) );
  NANDN U18714 ( .A(n17982), .B(n17981), .Z(n17986) );
  NANDN U18715 ( .A(n17984), .B(n17983), .Z(n17985) );
  AND U18716 ( .A(n17986), .B(n17985), .Z(n18127) );
  NANDN U18717 ( .A(n17988), .B(n17987), .Z(n17992) );
  NANDN U18718 ( .A(n17990), .B(n17989), .Z(n17991) );
  AND U18719 ( .A(n17992), .B(n17991), .Z(n18255) );
  NANDN U18720 ( .A(n17994), .B(n17993), .Z(n17998) );
  NAND U18721 ( .A(n17996), .B(n17995), .Z(n17997) );
  AND U18722 ( .A(n17998), .B(n17997), .Z(n18254) );
  XNOR U18723 ( .A(n18255), .B(n18254), .Z(n18257) );
  NANDN U18724 ( .A(n18000), .B(n17999), .Z(n18004) );
  NANDN U18725 ( .A(n18002), .B(n18001), .Z(n18003) );
  AND U18726 ( .A(n18004), .B(n18003), .Z(n18202) );
  NAND U18727 ( .A(n38385), .B(n18005), .Z(n18007) );
  XOR U18728 ( .A(b[27]), .B(a[110]), .Z(n18148) );
  NAND U18729 ( .A(n38343), .B(n18148), .Z(n18006) );
  AND U18730 ( .A(n18007), .B(n18006), .Z(n18209) );
  NAND U18731 ( .A(n183), .B(n18008), .Z(n18010) );
  XOR U18732 ( .A(b[5]), .B(a[132]), .Z(n18151) );
  NAND U18733 ( .A(n36296), .B(n18151), .Z(n18009) );
  AND U18734 ( .A(n18010), .B(n18009), .Z(n18207) );
  NAND U18735 ( .A(n190), .B(n18011), .Z(n18013) );
  XOR U18736 ( .A(b[19]), .B(a[118]), .Z(n18154) );
  NAND U18737 ( .A(n37821), .B(n18154), .Z(n18012) );
  NAND U18738 ( .A(n18013), .B(n18012), .Z(n18206) );
  XNOR U18739 ( .A(n18207), .B(n18206), .Z(n18208) );
  XNOR U18740 ( .A(n18209), .B(n18208), .Z(n18200) );
  NAND U18741 ( .A(n38470), .B(n18014), .Z(n18016) );
  XOR U18742 ( .A(b[31]), .B(a[106]), .Z(n18157) );
  NAND U18743 ( .A(n38453), .B(n18157), .Z(n18015) );
  AND U18744 ( .A(n18016), .B(n18015), .Z(n18169) );
  NAND U18745 ( .A(n181), .B(n18017), .Z(n18019) );
  XOR U18746 ( .A(b[3]), .B(a[134]), .Z(n18160) );
  NAND U18747 ( .A(n182), .B(n18160), .Z(n18018) );
  AND U18748 ( .A(n18019), .B(n18018), .Z(n18167) );
  NAND U18749 ( .A(n189), .B(n18020), .Z(n18022) );
  XOR U18750 ( .A(b[17]), .B(a[120]), .Z(n18163) );
  NAND U18751 ( .A(n37652), .B(n18163), .Z(n18021) );
  NAND U18752 ( .A(n18022), .B(n18021), .Z(n18166) );
  XNOR U18753 ( .A(n18167), .B(n18166), .Z(n18168) );
  XOR U18754 ( .A(n18169), .B(n18168), .Z(n18201) );
  XOR U18755 ( .A(n18200), .B(n18201), .Z(n18203) );
  XOR U18756 ( .A(n18202), .B(n18203), .Z(n18137) );
  NANDN U18757 ( .A(n18024), .B(n18023), .Z(n18028) );
  NANDN U18758 ( .A(n18026), .B(n18025), .Z(n18027) );
  AND U18759 ( .A(n18028), .B(n18027), .Z(n18190) );
  NANDN U18760 ( .A(n18030), .B(n18029), .Z(n18034) );
  NANDN U18761 ( .A(n18032), .B(n18031), .Z(n18033) );
  NAND U18762 ( .A(n18034), .B(n18033), .Z(n18191) );
  XNOR U18763 ( .A(n18190), .B(n18191), .Z(n18192) );
  NANDN U18764 ( .A(n18036), .B(n18035), .Z(n18040) );
  NANDN U18765 ( .A(n18038), .B(n18037), .Z(n18039) );
  NAND U18766 ( .A(n18040), .B(n18039), .Z(n18193) );
  XNOR U18767 ( .A(n18192), .B(n18193), .Z(n18136) );
  XNOR U18768 ( .A(n18137), .B(n18136), .Z(n18139) );
  NANDN U18769 ( .A(n18042), .B(n18041), .Z(n18046) );
  NANDN U18770 ( .A(n18044), .B(n18043), .Z(n18045) );
  AND U18771 ( .A(n18046), .B(n18045), .Z(n18138) );
  XOR U18772 ( .A(n18139), .B(n18138), .Z(n18251) );
  NANDN U18773 ( .A(n18048), .B(n18047), .Z(n18052) );
  NANDN U18774 ( .A(n18050), .B(n18049), .Z(n18051) );
  AND U18775 ( .A(n18052), .B(n18051), .Z(n18248) );
  NANDN U18776 ( .A(n18054), .B(n18053), .Z(n18058) );
  NANDN U18777 ( .A(n18056), .B(n18055), .Z(n18057) );
  AND U18778 ( .A(n18058), .B(n18057), .Z(n18133) );
  NANDN U18779 ( .A(n18060), .B(n18059), .Z(n18064) );
  OR U18780 ( .A(n18062), .B(n18061), .Z(n18063) );
  AND U18781 ( .A(n18064), .B(n18063), .Z(n18131) );
  NANDN U18782 ( .A(n18066), .B(n18065), .Z(n18070) );
  NANDN U18783 ( .A(n18068), .B(n18067), .Z(n18069) );
  AND U18784 ( .A(n18070), .B(n18069), .Z(n18197) );
  NANDN U18785 ( .A(n18072), .B(n18071), .Z(n18076) );
  NANDN U18786 ( .A(n18074), .B(n18073), .Z(n18075) );
  NAND U18787 ( .A(n18076), .B(n18075), .Z(n18196) );
  XNOR U18788 ( .A(n18197), .B(n18196), .Z(n18199) );
  NAND U18789 ( .A(n194), .B(n18077), .Z(n18079) );
  XOR U18790 ( .A(b[29]), .B(a[108]), .Z(n18221) );
  NAND U18791 ( .A(n38456), .B(n18221), .Z(n18078) );
  AND U18792 ( .A(n18079), .B(n18078), .Z(n18143) );
  AND U18793 ( .A(b[31]), .B(a[104]), .Z(n18142) );
  XNOR U18794 ( .A(n18143), .B(n18142), .Z(n18144) );
  NAND U18795 ( .A(b[0]), .B(a[136]), .Z(n18080) );
  XNOR U18796 ( .A(b[1]), .B(n18080), .Z(n18082) );
  NANDN U18797 ( .A(b[0]), .B(a[135]), .Z(n18081) );
  NAND U18798 ( .A(n18082), .B(n18081), .Z(n18145) );
  XNOR U18799 ( .A(n18144), .B(n18145), .Z(n18185) );
  NAND U18800 ( .A(n38185), .B(n18083), .Z(n18085) );
  XOR U18801 ( .A(b[23]), .B(a[114]), .Z(n18224) );
  NAND U18802 ( .A(n38132), .B(n18224), .Z(n18084) );
  AND U18803 ( .A(n18085), .B(n18084), .Z(n18214) );
  NAND U18804 ( .A(n184), .B(n18086), .Z(n18088) );
  XOR U18805 ( .A(b[7]), .B(a[130]), .Z(n18227) );
  NAND U18806 ( .A(n36592), .B(n18227), .Z(n18087) );
  AND U18807 ( .A(n18088), .B(n18087), .Z(n18213) );
  NAND U18808 ( .A(n38289), .B(n18089), .Z(n18091) );
  XOR U18809 ( .A(b[25]), .B(a[112]), .Z(n18230) );
  NAND U18810 ( .A(n38247), .B(n18230), .Z(n18090) );
  NAND U18811 ( .A(n18091), .B(n18090), .Z(n18212) );
  XOR U18812 ( .A(n18213), .B(n18212), .Z(n18215) );
  XOR U18813 ( .A(n18214), .B(n18215), .Z(n18184) );
  XOR U18814 ( .A(n18185), .B(n18184), .Z(n18187) );
  NAND U18815 ( .A(n187), .B(n18092), .Z(n18094) );
  XOR U18816 ( .A(b[13]), .B(a[124]), .Z(n18233) );
  NAND U18817 ( .A(n37295), .B(n18233), .Z(n18093) );
  AND U18818 ( .A(n18094), .B(n18093), .Z(n18179) );
  NAND U18819 ( .A(n186), .B(n18095), .Z(n18097) );
  XOR U18820 ( .A(b[11]), .B(a[126]), .Z(n18236) );
  NAND U18821 ( .A(n37097), .B(n18236), .Z(n18096) );
  NAND U18822 ( .A(n18097), .B(n18096), .Z(n18178) );
  XNOR U18823 ( .A(n18179), .B(n18178), .Z(n18181) );
  NAND U18824 ( .A(n188), .B(n18098), .Z(n18100) );
  XOR U18825 ( .A(b[15]), .B(a[122]), .Z(n18239) );
  NAND U18826 ( .A(n37382), .B(n18239), .Z(n18099) );
  AND U18827 ( .A(n18100), .B(n18099), .Z(n18175) );
  NAND U18828 ( .A(n38064), .B(n18101), .Z(n18103) );
  XOR U18829 ( .A(b[21]), .B(a[116]), .Z(n18242) );
  NAND U18830 ( .A(n37993), .B(n18242), .Z(n18102) );
  AND U18831 ( .A(n18103), .B(n18102), .Z(n18173) );
  NAND U18832 ( .A(n185), .B(n18104), .Z(n18106) );
  XOR U18833 ( .A(b[9]), .B(a[128]), .Z(n18245) );
  NAND U18834 ( .A(n36805), .B(n18245), .Z(n18105) );
  NAND U18835 ( .A(n18106), .B(n18105), .Z(n18172) );
  XNOR U18836 ( .A(n18173), .B(n18172), .Z(n18174) );
  XNOR U18837 ( .A(n18175), .B(n18174), .Z(n18180) );
  XOR U18838 ( .A(n18181), .B(n18180), .Z(n18186) );
  XNOR U18839 ( .A(n18187), .B(n18186), .Z(n18198) );
  XNOR U18840 ( .A(n18199), .B(n18198), .Z(n18130) );
  XNOR U18841 ( .A(n18131), .B(n18130), .Z(n18132) );
  XOR U18842 ( .A(n18133), .B(n18132), .Z(n18249) );
  XNOR U18843 ( .A(n18248), .B(n18249), .Z(n18250) );
  XNOR U18844 ( .A(n18251), .B(n18250), .Z(n18256) );
  XOR U18845 ( .A(n18257), .B(n18256), .Z(n18125) );
  NANDN U18846 ( .A(n18108), .B(n18107), .Z(n18112) );
  OR U18847 ( .A(n18110), .B(n18109), .Z(n18111) );
  AND U18848 ( .A(n18112), .B(n18111), .Z(n18124) );
  XNOR U18849 ( .A(n18125), .B(n18124), .Z(n18126) );
  XNOR U18850 ( .A(n18127), .B(n18126), .Z(n18118) );
  XNOR U18851 ( .A(n18119), .B(n18118), .Z(n18120) );
  XNOR U18852 ( .A(n18121), .B(n18120), .Z(n18260) );
  XNOR U18853 ( .A(sreg[360]), .B(n18260), .Z(n18262) );
  NANDN U18854 ( .A(sreg[359]), .B(n18113), .Z(n18117) );
  NAND U18855 ( .A(n18115), .B(n18114), .Z(n18116) );
  NAND U18856 ( .A(n18117), .B(n18116), .Z(n18261) );
  XNOR U18857 ( .A(n18262), .B(n18261), .Z(c[360]) );
  NANDN U18858 ( .A(n18119), .B(n18118), .Z(n18123) );
  NANDN U18859 ( .A(n18121), .B(n18120), .Z(n18122) );
  AND U18860 ( .A(n18123), .B(n18122), .Z(n18268) );
  NANDN U18861 ( .A(n18125), .B(n18124), .Z(n18129) );
  NANDN U18862 ( .A(n18127), .B(n18126), .Z(n18128) );
  AND U18863 ( .A(n18129), .B(n18128), .Z(n18266) );
  NANDN U18864 ( .A(n18131), .B(n18130), .Z(n18135) );
  NANDN U18865 ( .A(n18133), .B(n18132), .Z(n18134) );
  AND U18866 ( .A(n18135), .B(n18134), .Z(n18278) );
  NANDN U18867 ( .A(n18137), .B(n18136), .Z(n18141) );
  NAND U18868 ( .A(n18139), .B(n18138), .Z(n18140) );
  AND U18869 ( .A(n18141), .B(n18140), .Z(n18277) );
  XNOR U18870 ( .A(n18278), .B(n18277), .Z(n18280) );
  NANDN U18871 ( .A(n18143), .B(n18142), .Z(n18147) );
  NANDN U18872 ( .A(n18145), .B(n18144), .Z(n18146) );
  AND U18873 ( .A(n18147), .B(n18146), .Z(n18345) );
  NAND U18874 ( .A(n38385), .B(n18148), .Z(n18150) );
  XOR U18875 ( .A(b[27]), .B(a[111]), .Z(n18289) );
  NAND U18876 ( .A(n38343), .B(n18289), .Z(n18149) );
  AND U18877 ( .A(n18150), .B(n18149), .Z(n18352) );
  NAND U18878 ( .A(n183), .B(n18151), .Z(n18153) );
  XOR U18879 ( .A(b[5]), .B(a[133]), .Z(n18292) );
  NAND U18880 ( .A(n36296), .B(n18292), .Z(n18152) );
  AND U18881 ( .A(n18153), .B(n18152), .Z(n18350) );
  NAND U18882 ( .A(n190), .B(n18154), .Z(n18156) );
  XOR U18883 ( .A(b[19]), .B(a[119]), .Z(n18295) );
  NAND U18884 ( .A(n37821), .B(n18295), .Z(n18155) );
  NAND U18885 ( .A(n18156), .B(n18155), .Z(n18349) );
  XNOR U18886 ( .A(n18350), .B(n18349), .Z(n18351) );
  XNOR U18887 ( .A(n18352), .B(n18351), .Z(n18343) );
  NAND U18888 ( .A(n38470), .B(n18157), .Z(n18159) );
  XOR U18889 ( .A(b[31]), .B(a[107]), .Z(n18298) );
  NAND U18890 ( .A(n38453), .B(n18298), .Z(n18158) );
  AND U18891 ( .A(n18159), .B(n18158), .Z(n18310) );
  NAND U18892 ( .A(n181), .B(n18160), .Z(n18162) );
  XOR U18893 ( .A(b[3]), .B(a[135]), .Z(n18301) );
  NAND U18894 ( .A(n182), .B(n18301), .Z(n18161) );
  AND U18895 ( .A(n18162), .B(n18161), .Z(n18308) );
  NAND U18896 ( .A(n189), .B(n18163), .Z(n18165) );
  XOR U18897 ( .A(b[17]), .B(a[121]), .Z(n18304) );
  NAND U18898 ( .A(n37652), .B(n18304), .Z(n18164) );
  NAND U18899 ( .A(n18165), .B(n18164), .Z(n18307) );
  XNOR U18900 ( .A(n18308), .B(n18307), .Z(n18309) );
  XOR U18901 ( .A(n18310), .B(n18309), .Z(n18344) );
  XOR U18902 ( .A(n18343), .B(n18344), .Z(n18346) );
  XOR U18903 ( .A(n18345), .B(n18346), .Z(n18392) );
  NANDN U18904 ( .A(n18167), .B(n18166), .Z(n18171) );
  NANDN U18905 ( .A(n18169), .B(n18168), .Z(n18170) );
  AND U18906 ( .A(n18171), .B(n18170), .Z(n18331) );
  NANDN U18907 ( .A(n18173), .B(n18172), .Z(n18177) );
  NANDN U18908 ( .A(n18175), .B(n18174), .Z(n18176) );
  NAND U18909 ( .A(n18177), .B(n18176), .Z(n18332) );
  XNOR U18910 ( .A(n18331), .B(n18332), .Z(n18333) );
  NANDN U18911 ( .A(n18179), .B(n18178), .Z(n18183) );
  NAND U18912 ( .A(n18181), .B(n18180), .Z(n18182) );
  NAND U18913 ( .A(n18183), .B(n18182), .Z(n18334) );
  XNOR U18914 ( .A(n18333), .B(n18334), .Z(n18391) );
  XNOR U18915 ( .A(n18392), .B(n18391), .Z(n18394) );
  NAND U18916 ( .A(n18185), .B(n18184), .Z(n18189) );
  NAND U18917 ( .A(n18187), .B(n18186), .Z(n18188) );
  AND U18918 ( .A(n18189), .B(n18188), .Z(n18393) );
  XOR U18919 ( .A(n18394), .B(n18393), .Z(n18406) );
  NANDN U18920 ( .A(n18191), .B(n18190), .Z(n18195) );
  NANDN U18921 ( .A(n18193), .B(n18192), .Z(n18194) );
  AND U18922 ( .A(n18195), .B(n18194), .Z(n18403) );
  NANDN U18923 ( .A(n18201), .B(n18200), .Z(n18205) );
  OR U18924 ( .A(n18203), .B(n18202), .Z(n18204) );
  AND U18925 ( .A(n18205), .B(n18204), .Z(n18398) );
  NANDN U18926 ( .A(n18207), .B(n18206), .Z(n18211) );
  NANDN U18927 ( .A(n18209), .B(n18208), .Z(n18210) );
  AND U18928 ( .A(n18211), .B(n18210), .Z(n18338) );
  NANDN U18929 ( .A(n18213), .B(n18212), .Z(n18217) );
  OR U18930 ( .A(n18215), .B(n18214), .Z(n18216) );
  NAND U18931 ( .A(n18217), .B(n18216), .Z(n18337) );
  XNOR U18932 ( .A(n18338), .B(n18337), .Z(n18339) );
  NAND U18933 ( .A(b[0]), .B(a[137]), .Z(n18218) );
  XNOR U18934 ( .A(b[1]), .B(n18218), .Z(n18220) );
  NANDN U18935 ( .A(b[0]), .B(a[136]), .Z(n18219) );
  NAND U18936 ( .A(n18220), .B(n18219), .Z(n18286) );
  NAND U18937 ( .A(n194), .B(n18221), .Z(n18223) );
  XOR U18938 ( .A(b[29]), .B(a[109]), .Z(n18364) );
  NAND U18939 ( .A(n38456), .B(n18364), .Z(n18222) );
  AND U18940 ( .A(n18223), .B(n18222), .Z(n18284) );
  AND U18941 ( .A(b[31]), .B(a[105]), .Z(n18283) );
  XNOR U18942 ( .A(n18284), .B(n18283), .Z(n18285) );
  XNOR U18943 ( .A(n18286), .B(n18285), .Z(n18325) );
  NAND U18944 ( .A(n38185), .B(n18224), .Z(n18226) );
  XOR U18945 ( .A(b[23]), .B(a[115]), .Z(n18367) );
  NAND U18946 ( .A(n38132), .B(n18367), .Z(n18225) );
  AND U18947 ( .A(n18226), .B(n18225), .Z(n18358) );
  NAND U18948 ( .A(n184), .B(n18227), .Z(n18229) );
  XOR U18949 ( .A(b[7]), .B(a[131]), .Z(n18370) );
  NAND U18950 ( .A(n36592), .B(n18370), .Z(n18228) );
  AND U18951 ( .A(n18229), .B(n18228), .Z(n18356) );
  NAND U18952 ( .A(n38289), .B(n18230), .Z(n18232) );
  XOR U18953 ( .A(b[25]), .B(a[113]), .Z(n18373) );
  NAND U18954 ( .A(n38247), .B(n18373), .Z(n18231) );
  NAND U18955 ( .A(n18232), .B(n18231), .Z(n18355) );
  XNOR U18956 ( .A(n18356), .B(n18355), .Z(n18357) );
  XOR U18957 ( .A(n18358), .B(n18357), .Z(n18326) );
  XNOR U18958 ( .A(n18325), .B(n18326), .Z(n18327) );
  NAND U18959 ( .A(n187), .B(n18233), .Z(n18235) );
  XOR U18960 ( .A(b[13]), .B(a[125]), .Z(n18376) );
  NAND U18961 ( .A(n37295), .B(n18376), .Z(n18234) );
  AND U18962 ( .A(n18235), .B(n18234), .Z(n18320) );
  NAND U18963 ( .A(n186), .B(n18236), .Z(n18238) );
  XOR U18964 ( .A(b[11]), .B(a[127]), .Z(n18379) );
  NAND U18965 ( .A(n37097), .B(n18379), .Z(n18237) );
  NAND U18966 ( .A(n18238), .B(n18237), .Z(n18319) );
  XNOR U18967 ( .A(n18320), .B(n18319), .Z(n18321) );
  NAND U18968 ( .A(n188), .B(n18239), .Z(n18241) );
  XOR U18969 ( .A(b[15]), .B(a[123]), .Z(n18382) );
  NAND U18970 ( .A(n37382), .B(n18382), .Z(n18240) );
  AND U18971 ( .A(n18241), .B(n18240), .Z(n18316) );
  NAND U18972 ( .A(n38064), .B(n18242), .Z(n18244) );
  XOR U18973 ( .A(b[21]), .B(a[117]), .Z(n18385) );
  NAND U18974 ( .A(n37993), .B(n18385), .Z(n18243) );
  AND U18975 ( .A(n18244), .B(n18243), .Z(n18314) );
  NAND U18976 ( .A(n185), .B(n18245), .Z(n18247) );
  XOR U18977 ( .A(b[9]), .B(a[129]), .Z(n18388) );
  NAND U18978 ( .A(n36805), .B(n18388), .Z(n18246) );
  NAND U18979 ( .A(n18247), .B(n18246), .Z(n18313) );
  XNOR U18980 ( .A(n18314), .B(n18313), .Z(n18315) );
  XOR U18981 ( .A(n18316), .B(n18315), .Z(n18322) );
  XOR U18982 ( .A(n18321), .B(n18322), .Z(n18328) );
  XOR U18983 ( .A(n18327), .B(n18328), .Z(n18340) );
  XNOR U18984 ( .A(n18339), .B(n18340), .Z(n18397) );
  XNOR U18985 ( .A(n18398), .B(n18397), .Z(n18399) );
  XOR U18986 ( .A(n18400), .B(n18399), .Z(n18404) );
  XNOR U18987 ( .A(n18403), .B(n18404), .Z(n18405) );
  XNOR U18988 ( .A(n18406), .B(n18405), .Z(n18279) );
  XOR U18989 ( .A(n18280), .B(n18279), .Z(n18272) );
  NANDN U18990 ( .A(n18249), .B(n18248), .Z(n18253) );
  NANDN U18991 ( .A(n18251), .B(n18250), .Z(n18252) );
  AND U18992 ( .A(n18253), .B(n18252), .Z(n18271) );
  XNOR U18993 ( .A(n18272), .B(n18271), .Z(n18273) );
  NANDN U18994 ( .A(n18255), .B(n18254), .Z(n18259) );
  NAND U18995 ( .A(n18257), .B(n18256), .Z(n18258) );
  NAND U18996 ( .A(n18259), .B(n18258), .Z(n18274) );
  XNOR U18997 ( .A(n18273), .B(n18274), .Z(n18265) );
  XNOR U18998 ( .A(n18266), .B(n18265), .Z(n18267) );
  XNOR U18999 ( .A(n18268), .B(n18267), .Z(n18409) );
  XNOR U19000 ( .A(sreg[361]), .B(n18409), .Z(n18411) );
  NANDN U19001 ( .A(sreg[360]), .B(n18260), .Z(n18264) );
  NAND U19002 ( .A(n18262), .B(n18261), .Z(n18263) );
  NAND U19003 ( .A(n18264), .B(n18263), .Z(n18410) );
  XNOR U19004 ( .A(n18411), .B(n18410), .Z(c[361]) );
  NANDN U19005 ( .A(n18266), .B(n18265), .Z(n18270) );
  NANDN U19006 ( .A(n18268), .B(n18267), .Z(n18269) );
  AND U19007 ( .A(n18270), .B(n18269), .Z(n18417) );
  NANDN U19008 ( .A(n18272), .B(n18271), .Z(n18276) );
  NANDN U19009 ( .A(n18274), .B(n18273), .Z(n18275) );
  AND U19010 ( .A(n18276), .B(n18275), .Z(n18415) );
  NANDN U19011 ( .A(n18278), .B(n18277), .Z(n18282) );
  NAND U19012 ( .A(n18280), .B(n18279), .Z(n18281) );
  AND U19013 ( .A(n18282), .B(n18281), .Z(n18422) );
  NANDN U19014 ( .A(n18284), .B(n18283), .Z(n18288) );
  NANDN U19015 ( .A(n18286), .B(n18285), .Z(n18287) );
  AND U19016 ( .A(n18288), .B(n18287), .Z(n18506) );
  NAND U19017 ( .A(n38385), .B(n18289), .Z(n18291) );
  XOR U19018 ( .A(b[27]), .B(a[112]), .Z(n18450) );
  NAND U19019 ( .A(n38343), .B(n18450), .Z(n18290) );
  AND U19020 ( .A(n18291), .B(n18290), .Z(n18513) );
  NAND U19021 ( .A(n183), .B(n18292), .Z(n18294) );
  XOR U19022 ( .A(b[5]), .B(a[134]), .Z(n18453) );
  NAND U19023 ( .A(n36296), .B(n18453), .Z(n18293) );
  AND U19024 ( .A(n18294), .B(n18293), .Z(n18511) );
  NAND U19025 ( .A(n190), .B(n18295), .Z(n18297) );
  XOR U19026 ( .A(b[19]), .B(a[120]), .Z(n18456) );
  NAND U19027 ( .A(n37821), .B(n18456), .Z(n18296) );
  NAND U19028 ( .A(n18297), .B(n18296), .Z(n18510) );
  XNOR U19029 ( .A(n18511), .B(n18510), .Z(n18512) );
  XNOR U19030 ( .A(n18513), .B(n18512), .Z(n18504) );
  NAND U19031 ( .A(n38470), .B(n18298), .Z(n18300) );
  XOR U19032 ( .A(b[31]), .B(a[108]), .Z(n18459) );
  NAND U19033 ( .A(n38453), .B(n18459), .Z(n18299) );
  AND U19034 ( .A(n18300), .B(n18299), .Z(n18471) );
  NAND U19035 ( .A(n181), .B(n18301), .Z(n18303) );
  XOR U19036 ( .A(b[3]), .B(a[136]), .Z(n18462) );
  NAND U19037 ( .A(n182), .B(n18462), .Z(n18302) );
  AND U19038 ( .A(n18303), .B(n18302), .Z(n18469) );
  NAND U19039 ( .A(n189), .B(n18304), .Z(n18306) );
  XOR U19040 ( .A(b[17]), .B(a[122]), .Z(n18465) );
  NAND U19041 ( .A(n37652), .B(n18465), .Z(n18305) );
  NAND U19042 ( .A(n18306), .B(n18305), .Z(n18468) );
  XNOR U19043 ( .A(n18469), .B(n18468), .Z(n18470) );
  XOR U19044 ( .A(n18471), .B(n18470), .Z(n18505) );
  XOR U19045 ( .A(n18504), .B(n18505), .Z(n18507) );
  XOR U19046 ( .A(n18506), .B(n18507), .Z(n18439) );
  NANDN U19047 ( .A(n18308), .B(n18307), .Z(n18312) );
  NANDN U19048 ( .A(n18310), .B(n18309), .Z(n18311) );
  AND U19049 ( .A(n18312), .B(n18311), .Z(n18492) );
  NANDN U19050 ( .A(n18314), .B(n18313), .Z(n18318) );
  NANDN U19051 ( .A(n18316), .B(n18315), .Z(n18317) );
  NAND U19052 ( .A(n18318), .B(n18317), .Z(n18493) );
  XNOR U19053 ( .A(n18492), .B(n18493), .Z(n18494) );
  NANDN U19054 ( .A(n18320), .B(n18319), .Z(n18324) );
  NANDN U19055 ( .A(n18322), .B(n18321), .Z(n18323) );
  NAND U19056 ( .A(n18324), .B(n18323), .Z(n18495) );
  XNOR U19057 ( .A(n18494), .B(n18495), .Z(n18438) );
  XNOR U19058 ( .A(n18439), .B(n18438), .Z(n18441) );
  NANDN U19059 ( .A(n18326), .B(n18325), .Z(n18330) );
  NANDN U19060 ( .A(n18328), .B(n18327), .Z(n18329) );
  AND U19061 ( .A(n18330), .B(n18329), .Z(n18440) );
  XOR U19062 ( .A(n18441), .B(n18440), .Z(n18554) );
  NANDN U19063 ( .A(n18332), .B(n18331), .Z(n18336) );
  NANDN U19064 ( .A(n18334), .B(n18333), .Z(n18335) );
  AND U19065 ( .A(n18336), .B(n18335), .Z(n18552) );
  NANDN U19066 ( .A(n18338), .B(n18337), .Z(n18342) );
  NANDN U19067 ( .A(n18340), .B(n18339), .Z(n18341) );
  AND U19068 ( .A(n18342), .B(n18341), .Z(n18435) );
  NANDN U19069 ( .A(n18344), .B(n18343), .Z(n18348) );
  OR U19070 ( .A(n18346), .B(n18345), .Z(n18347) );
  AND U19071 ( .A(n18348), .B(n18347), .Z(n18433) );
  NANDN U19072 ( .A(n18350), .B(n18349), .Z(n18354) );
  NANDN U19073 ( .A(n18352), .B(n18351), .Z(n18353) );
  AND U19074 ( .A(n18354), .B(n18353), .Z(n18499) );
  NANDN U19075 ( .A(n18356), .B(n18355), .Z(n18360) );
  NANDN U19076 ( .A(n18358), .B(n18357), .Z(n18359) );
  NAND U19077 ( .A(n18360), .B(n18359), .Z(n18498) );
  XNOR U19078 ( .A(n18499), .B(n18498), .Z(n18500) );
  NAND U19079 ( .A(b[0]), .B(a[138]), .Z(n18361) );
  XNOR U19080 ( .A(b[1]), .B(n18361), .Z(n18363) );
  NANDN U19081 ( .A(b[0]), .B(a[137]), .Z(n18362) );
  NAND U19082 ( .A(n18363), .B(n18362), .Z(n18447) );
  NAND U19083 ( .A(n194), .B(n18364), .Z(n18366) );
  XOR U19084 ( .A(b[29]), .B(a[110]), .Z(n18522) );
  NAND U19085 ( .A(n38456), .B(n18522), .Z(n18365) );
  AND U19086 ( .A(n18366), .B(n18365), .Z(n18445) );
  AND U19087 ( .A(b[31]), .B(a[106]), .Z(n18444) );
  XNOR U19088 ( .A(n18445), .B(n18444), .Z(n18446) );
  XNOR U19089 ( .A(n18447), .B(n18446), .Z(n18486) );
  NAND U19090 ( .A(n38185), .B(n18367), .Z(n18369) );
  XOR U19091 ( .A(b[23]), .B(a[116]), .Z(n18528) );
  NAND U19092 ( .A(n38132), .B(n18528), .Z(n18368) );
  AND U19093 ( .A(n18369), .B(n18368), .Z(n18519) );
  NAND U19094 ( .A(n184), .B(n18370), .Z(n18372) );
  XOR U19095 ( .A(b[7]), .B(a[132]), .Z(n18531) );
  NAND U19096 ( .A(n36592), .B(n18531), .Z(n18371) );
  AND U19097 ( .A(n18372), .B(n18371), .Z(n18517) );
  NAND U19098 ( .A(n38289), .B(n18373), .Z(n18375) );
  XOR U19099 ( .A(b[25]), .B(a[114]), .Z(n18534) );
  NAND U19100 ( .A(n38247), .B(n18534), .Z(n18374) );
  NAND U19101 ( .A(n18375), .B(n18374), .Z(n18516) );
  XNOR U19102 ( .A(n18517), .B(n18516), .Z(n18518) );
  XOR U19103 ( .A(n18519), .B(n18518), .Z(n18487) );
  XNOR U19104 ( .A(n18486), .B(n18487), .Z(n18488) );
  NAND U19105 ( .A(n187), .B(n18376), .Z(n18378) );
  XOR U19106 ( .A(b[13]), .B(a[126]), .Z(n18537) );
  NAND U19107 ( .A(n37295), .B(n18537), .Z(n18377) );
  AND U19108 ( .A(n18378), .B(n18377), .Z(n18481) );
  NAND U19109 ( .A(n186), .B(n18379), .Z(n18381) );
  XOR U19110 ( .A(b[11]), .B(a[128]), .Z(n18540) );
  NAND U19111 ( .A(n37097), .B(n18540), .Z(n18380) );
  NAND U19112 ( .A(n18381), .B(n18380), .Z(n18480) );
  XNOR U19113 ( .A(n18481), .B(n18480), .Z(n18482) );
  NAND U19114 ( .A(n188), .B(n18382), .Z(n18384) );
  XOR U19115 ( .A(b[15]), .B(a[124]), .Z(n18543) );
  NAND U19116 ( .A(n37382), .B(n18543), .Z(n18383) );
  AND U19117 ( .A(n18384), .B(n18383), .Z(n18477) );
  NAND U19118 ( .A(n38064), .B(n18385), .Z(n18387) );
  XOR U19119 ( .A(b[21]), .B(a[118]), .Z(n18546) );
  NAND U19120 ( .A(n37993), .B(n18546), .Z(n18386) );
  AND U19121 ( .A(n18387), .B(n18386), .Z(n18475) );
  NAND U19122 ( .A(n185), .B(n18388), .Z(n18390) );
  XOR U19123 ( .A(b[9]), .B(a[130]), .Z(n18549) );
  NAND U19124 ( .A(n36805), .B(n18549), .Z(n18389) );
  NAND U19125 ( .A(n18390), .B(n18389), .Z(n18474) );
  XNOR U19126 ( .A(n18475), .B(n18474), .Z(n18476) );
  XOR U19127 ( .A(n18477), .B(n18476), .Z(n18483) );
  XOR U19128 ( .A(n18482), .B(n18483), .Z(n18489) );
  XOR U19129 ( .A(n18488), .B(n18489), .Z(n18501) );
  XNOR U19130 ( .A(n18500), .B(n18501), .Z(n18432) );
  XNOR U19131 ( .A(n18433), .B(n18432), .Z(n18434) );
  XOR U19132 ( .A(n18435), .B(n18434), .Z(n18553) );
  XOR U19133 ( .A(n18552), .B(n18553), .Z(n18555) );
  XOR U19134 ( .A(n18554), .B(n18555), .Z(n18429) );
  NANDN U19135 ( .A(n18392), .B(n18391), .Z(n18396) );
  NAND U19136 ( .A(n18394), .B(n18393), .Z(n18395) );
  AND U19137 ( .A(n18396), .B(n18395), .Z(n18427) );
  NANDN U19138 ( .A(n18398), .B(n18397), .Z(n18402) );
  NANDN U19139 ( .A(n18400), .B(n18399), .Z(n18401) );
  AND U19140 ( .A(n18402), .B(n18401), .Z(n18426) );
  XNOR U19141 ( .A(n18427), .B(n18426), .Z(n18428) );
  XNOR U19142 ( .A(n18429), .B(n18428), .Z(n18420) );
  NANDN U19143 ( .A(n18404), .B(n18403), .Z(n18408) );
  NANDN U19144 ( .A(n18406), .B(n18405), .Z(n18407) );
  NAND U19145 ( .A(n18408), .B(n18407), .Z(n18421) );
  XOR U19146 ( .A(n18420), .B(n18421), .Z(n18423) );
  XNOR U19147 ( .A(n18422), .B(n18423), .Z(n18414) );
  XNOR U19148 ( .A(n18415), .B(n18414), .Z(n18416) );
  XNOR U19149 ( .A(n18417), .B(n18416), .Z(n18558) );
  XNOR U19150 ( .A(sreg[362]), .B(n18558), .Z(n18560) );
  NANDN U19151 ( .A(sreg[361]), .B(n18409), .Z(n18413) );
  NAND U19152 ( .A(n18411), .B(n18410), .Z(n18412) );
  NAND U19153 ( .A(n18413), .B(n18412), .Z(n18559) );
  XNOR U19154 ( .A(n18560), .B(n18559), .Z(c[362]) );
  NANDN U19155 ( .A(n18415), .B(n18414), .Z(n18419) );
  NANDN U19156 ( .A(n18417), .B(n18416), .Z(n18418) );
  AND U19157 ( .A(n18419), .B(n18418), .Z(n18566) );
  NANDN U19158 ( .A(n18421), .B(n18420), .Z(n18425) );
  NANDN U19159 ( .A(n18423), .B(n18422), .Z(n18424) );
  AND U19160 ( .A(n18425), .B(n18424), .Z(n18564) );
  NANDN U19161 ( .A(n18427), .B(n18426), .Z(n18431) );
  NANDN U19162 ( .A(n18429), .B(n18428), .Z(n18430) );
  AND U19163 ( .A(n18431), .B(n18430), .Z(n18572) );
  NANDN U19164 ( .A(n18433), .B(n18432), .Z(n18437) );
  NANDN U19165 ( .A(n18435), .B(n18434), .Z(n18436) );
  AND U19166 ( .A(n18437), .B(n18436), .Z(n18576) );
  NANDN U19167 ( .A(n18439), .B(n18438), .Z(n18443) );
  NAND U19168 ( .A(n18441), .B(n18440), .Z(n18442) );
  AND U19169 ( .A(n18443), .B(n18442), .Z(n18575) );
  XNOR U19170 ( .A(n18576), .B(n18575), .Z(n18578) );
  NANDN U19171 ( .A(n18445), .B(n18444), .Z(n18449) );
  NANDN U19172 ( .A(n18447), .B(n18446), .Z(n18448) );
  AND U19173 ( .A(n18449), .B(n18448), .Z(n18655) );
  NAND U19174 ( .A(n38385), .B(n18450), .Z(n18452) );
  XOR U19175 ( .A(b[27]), .B(a[113]), .Z(n18599) );
  NAND U19176 ( .A(n38343), .B(n18599), .Z(n18451) );
  AND U19177 ( .A(n18452), .B(n18451), .Z(n18662) );
  NAND U19178 ( .A(n183), .B(n18453), .Z(n18455) );
  XOR U19179 ( .A(b[5]), .B(a[135]), .Z(n18602) );
  NAND U19180 ( .A(n36296), .B(n18602), .Z(n18454) );
  AND U19181 ( .A(n18455), .B(n18454), .Z(n18660) );
  NAND U19182 ( .A(n190), .B(n18456), .Z(n18458) );
  XOR U19183 ( .A(b[19]), .B(a[121]), .Z(n18605) );
  NAND U19184 ( .A(n37821), .B(n18605), .Z(n18457) );
  NAND U19185 ( .A(n18458), .B(n18457), .Z(n18659) );
  XNOR U19186 ( .A(n18660), .B(n18659), .Z(n18661) );
  XNOR U19187 ( .A(n18662), .B(n18661), .Z(n18653) );
  NAND U19188 ( .A(n38470), .B(n18459), .Z(n18461) );
  XOR U19189 ( .A(b[31]), .B(a[109]), .Z(n18608) );
  NAND U19190 ( .A(n38453), .B(n18608), .Z(n18460) );
  AND U19191 ( .A(n18461), .B(n18460), .Z(n18620) );
  NAND U19192 ( .A(n181), .B(n18462), .Z(n18464) );
  XOR U19193 ( .A(b[3]), .B(a[137]), .Z(n18611) );
  NAND U19194 ( .A(n182), .B(n18611), .Z(n18463) );
  AND U19195 ( .A(n18464), .B(n18463), .Z(n18618) );
  NAND U19196 ( .A(n189), .B(n18465), .Z(n18467) );
  XOR U19197 ( .A(b[17]), .B(a[123]), .Z(n18614) );
  NAND U19198 ( .A(n37652), .B(n18614), .Z(n18466) );
  NAND U19199 ( .A(n18467), .B(n18466), .Z(n18617) );
  XNOR U19200 ( .A(n18618), .B(n18617), .Z(n18619) );
  XOR U19201 ( .A(n18620), .B(n18619), .Z(n18654) );
  XOR U19202 ( .A(n18653), .B(n18654), .Z(n18656) );
  XOR U19203 ( .A(n18655), .B(n18656), .Z(n18588) );
  NANDN U19204 ( .A(n18469), .B(n18468), .Z(n18473) );
  NANDN U19205 ( .A(n18471), .B(n18470), .Z(n18472) );
  AND U19206 ( .A(n18473), .B(n18472), .Z(n18641) );
  NANDN U19207 ( .A(n18475), .B(n18474), .Z(n18479) );
  NANDN U19208 ( .A(n18477), .B(n18476), .Z(n18478) );
  NAND U19209 ( .A(n18479), .B(n18478), .Z(n18642) );
  XNOR U19210 ( .A(n18641), .B(n18642), .Z(n18643) );
  NANDN U19211 ( .A(n18481), .B(n18480), .Z(n18485) );
  NANDN U19212 ( .A(n18483), .B(n18482), .Z(n18484) );
  NAND U19213 ( .A(n18485), .B(n18484), .Z(n18644) );
  XNOR U19214 ( .A(n18643), .B(n18644), .Z(n18587) );
  XNOR U19215 ( .A(n18588), .B(n18587), .Z(n18590) );
  NANDN U19216 ( .A(n18487), .B(n18486), .Z(n18491) );
  NANDN U19217 ( .A(n18489), .B(n18488), .Z(n18490) );
  AND U19218 ( .A(n18491), .B(n18490), .Z(n18589) );
  XOR U19219 ( .A(n18590), .B(n18589), .Z(n18704) );
  NANDN U19220 ( .A(n18493), .B(n18492), .Z(n18497) );
  NANDN U19221 ( .A(n18495), .B(n18494), .Z(n18496) );
  AND U19222 ( .A(n18497), .B(n18496), .Z(n18701) );
  NANDN U19223 ( .A(n18499), .B(n18498), .Z(n18503) );
  NANDN U19224 ( .A(n18501), .B(n18500), .Z(n18502) );
  AND U19225 ( .A(n18503), .B(n18502), .Z(n18584) );
  NANDN U19226 ( .A(n18505), .B(n18504), .Z(n18509) );
  OR U19227 ( .A(n18507), .B(n18506), .Z(n18508) );
  AND U19228 ( .A(n18509), .B(n18508), .Z(n18582) );
  NANDN U19229 ( .A(n18511), .B(n18510), .Z(n18515) );
  NANDN U19230 ( .A(n18513), .B(n18512), .Z(n18514) );
  AND U19231 ( .A(n18515), .B(n18514), .Z(n18648) );
  NANDN U19232 ( .A(n18517), .B(n18516), .Z(n18521) );
  NANDN U19233 ( .A(n18519), .B(n18518), .Z(n18520) );
  NAND U19234 ( .A(n18521), .B(n18520), .Z(n18647) );
  XNOR U19235 ( .A(n18648), .B(n18647), .Z(n18649) );
  NAND U19236 ( .A(n194), .B(n18522), .Z(n18524) );
  XOR U19237 ( .A(b[29]), .B(a[111]), .Z(n18674) );
  NAND U19238 ( .A(n38456), .B(n18674), .Z(n18523) );
  AND U19239 ( .A(n18524), .B(n18523), .Z(n18594) );
  AND U19240 ( .A(b[31]), .B(a[107]), .Z(n18593) );
  XNOR U19241 ( .A(n18594), .B(n18593), .Z(n18595) );
  NAND U19242 ( .A(b[0]), .B(a[139]), .Z(n18525) );
  XNOR U19243 ( .A(b[1]), .B(n18525), .Z(n18527) );
  NANDN U19244 ( .A(b[0]), .B(a[138]), .Z(n18526) );
  NAND U19245 ( .A(n18527), .B(n18526), .Z(n18596) );
  XNOR U19246 ( .A(n18595), .B(n18596), .Z(n18635) );
  NAND U19247 ( .A(n38185), .B(n18528), .Z(n18530) );
  XOR U19248 ( .A(b[23]), .B(a[117]), .Z(n18677) );
  NAND U19249 ( .A(n38132), .B(n18677), .Z(n18529) );
  AND U19250 ( .A(n18530), .B(n18529), .Z(n18668) );
  NAND U19251 ( .A(n184), .B(n18531), .Z(n18533) );
  XOR U19252 ( .A(b[7]), .B(a[133]), .Z(n18680) );
  NAND U19253 ( .A(n36592), .B(n18680), .Z(n18532) );
  AND U19254 ( .A(n18533), .B(n18532), .Z(n18666) );
  NAND U19255 ( .A(n38289), .B(n18534), .Z(n18536) );
  XOR U19256 ( .A(b[25]), .B(a[115]), .Z(n18683) );
  NAND U19257 ( .A(n38247), .B(n18683), .Z(n18535) );
  NAND U19258 ( .A(n18536), .B(n18535), .Z(n18665) );
  XNOR U19259 ( .A(n18666), .B(n18665), .Z(n18667) );
  XOR U19260 ( .A(n18668), .B(n18667), .Z(n18636) );
  XNOR U19261 ( .A(n18635), .B(n18636), .Z(n18637) );
  NAND U19262 ( .A(n187), .B(n18537), .Z(n18539) );
  XOR U19263 ( .A(b[13]), .B(a[127]), .Z(n18686) );
  NAND U19264 ( .A(n37295), .B(n18686), .Z(n18538) );
  AND U19265 ( .A(n18539), .B(n18538), .Z(n18630) );
  NAND U19266 ( .A(n186), .B(n18540), .Z(n18542) );
  XOR U19267 ( .A(b[11]), .B(a[129]), .Z(n18689) );
  NAND U19268 ( .A(n37097), .B(n18689), .Z(n18541) );
  NAND U19269 ( .A(n18542), .B(n18541), .Z(n18629) );
  XNOR U19270 ( .A(n18630), .B(n18629), .Z(n18631) );
  NAND U19271 ( .A(n188), .B(n18543), .Z(n18545) );
  XOR U19272 ( .A(b[15]), .B(a[125]), .Z(n18692) );
  NAND U19273 ( .A(n37382), .B(n18692), .Z(n18544) );
  AND U19274 ( .A(n18545), .B(n18544), .Z(n18626) );
  NAND U19275 ( .A(n38064), .B(n18546), .Z(n18548) );
  XOR U19276 ( .A(b[21]), .B(a[119]), .Z(n18695) );
  NAND U19277 ( .A(n37993), .B(n18695), .Z(n18547) );
  AND U19278 ( .A(n18548), .B(n18547), .Z(n18624) );
  NAND U19279 ( .A(n185), .B(n18549), .Z(n18551) );
  XOR U19280 ( .A(b[9]), .B(a[131]), .Z(n18698) );
  NAND U19281 ( .A(n36805), .B(n18698), .Z(n18550) );
  NAND U19282 ( .A(n18551), .B(n18550), .Z(n18623) );
  XNOR U19283 ( .A(n18624), .B(n18623), .Z(n18625) );
  XOR U19284 ( .A(n18626), .B(n18625), .Z(n18632) );
  XOR U19285 ( .A(n18631), .B(n18632), .Z(n18638) );
  XOR U19286 ( .A(n18637), .B(n18638), .Z(n18650) );
  XNOR U19287 ( .A(n18649), .B(n18650), .Z(n18581) );
  XNOR U19288 ( .A(n18582), .B(n18581), .Z(n18583) );
  XOR U19289 ( .A(n18584), .B(n18583), .Z(n18702) );
  XNOR U19290 ( .A(n18701), .B(n18702), .Z(n18703) );
  XNOR U19291 ( .A(n18704), .B(n18703), .Z(n18577) );
  XOR U19292 ( .A(n18578), .B(n18577), .Z(n18570) );
  NANDN U19293 ( .A(n18553), .B(n18552), .Z(n18557) );
  OR U19294 ( .A(n18555), .B(n18554), .Z(n18556) );
  AND U19295 ( .A(n18557), .B(n18556), .Z(n18569) );
  XNOR U19296 ( .A(n18570), .B(n18569), .Z(n18571) );
  XNOR U19297 ( .A(n18572), .B(n18571), .Z(n18563) );
  XNOR U19298 ( .A(n18564), .B(n18563), .Z(n18565) );
  XNOR U19299 ( .A(n18566), .B(n18565), .Z(n18707) );
  XNOR U19300 ( .A(sreg[363]), .B(n18707), .Z(n18709) );
  NANDN U19301 ( .A(sreg[362]), .B(n18558), .Z(n18562) );
  NAND U19302 ( .A(n18560), .B(n18559), .Z(n18561) );
  NAND U19303 ( .A(n18562), .B(n18561), .Z(n18708) );
  XNOR U19304 ( .A(n18709), .B(n18708), .Z(c[363]) );
  NANDN U19305 ( .A(n18564), .B(n18563), .Z(n18568) );
  NANDN U19306 ( .A(n18566), .B(n18565), .Z(n18567) );
  AND U19307 ( .A(n18568), .B(n18567), .Z(n18715) );
  NANDN U19308 ( .A(n18570), .B(n18569), .Z(n18574) );
  NANDN U19309 ( .A(n18572), .B(n18571), .Z(n18573) );
  AND U19310 ( .A(n18574), .B(n18573), .Z(n18713) );
  NANDN U19311 ( .A(n18576), .B(n18575), .Z(n18580) );
  NAND U19312 ( .A(n18578), .B(n18577), .Z(n18579) );
  AND U19313 ( .A(n18580), .B(n18579), .Z(n18720) );
  NANDN U19314 ( .A(n18582), .B(n18581), .Z(n18586) );
  NANDN U19315 ( .A(n18584), .B(n18583), .Z(n18585) );
  AND U19316 ( .A(n18586), .B(n18585), .Z(n18851) );
  NANDN U19317 ( .A(n18588), .B(n18587), .Z(n18592) );
  NAND U19318 ( .A(n18590), .B(n18589), .Z(n18591) );
  AND U19319 ( .A(n18592), .B(n18591), .Z(n18850) );
  XNOR U19320 ( .A(n18851), .B(n18850), .Z(n18853) );
  NANDN U19321 ( .A(n18594), .B(n18593), .Z(n18598) );
  NANDN U19322 ( .A(n18596), .B(n18595), .Z(n18597) );
  AND U19323 ( .A(n18598), .B(n18597), .Z(n18798) );
  NAND U19324 ( .A(n38385), .B(n18599), .Z(n18601) );
  XOR U19325 ( .A(b[27]), .B(a[114]), .Z(n18742) );
  NAND U19326 ( .A(n38343), .B(n18742), .Z(n18600) );
  AND U19327 ( .A(n18601), .B(n18600), .Z(n18805) );
  NAND U19328 ( .A(n183), .B(n18602), .Z(n18604) );
  XOR U19329 ( .A(b[5]), .B(a[136]), .Z(n18745) );
  NAND U19330 ( .A(n36296), .B(n18745), .Z(n18603) );
  AND U19331 ( .A(n18604), .B(n18603), .Z(n18803) );
  NAND U19332 ( .A(n190), .B(n18605), .Z(n18607) );
  XOR U19333 ( .A(b[19]), .B(a[122]), .Z(n18748) );
  NAND U19334 ( .A(n37821), .B(n18748), .Z(n18606) );
  NAND U19335 ( .A(n18607), .B(n18606), .Z(n18802) );
  XNOR U19336 ( .A(n18803), .B(n18802), .Z(n18804) );
  XNOR U19337 ( .A(n18805), .B(n18804), .Z(n18796) );
  NAND U19338 ( .A(n38470), .B(n18608), .Z(n18610) );
  XOR U19339 ( .A(b[31]), .B(a[110]), .Z(n18751) );
  NAND U19340 ( .A(n38453), .B(n18751), .Z(n18609) );
  AND U19341 ( .A(n18610), .B(n18609), .Z(n18763) );
  NAND U19342 ( .A(n181), .B(n18611), .Z(n18613) );
  XOR U19343 ( .A(b[3]), .B(a[138]), .Z(n18754) );
  NAND U19344 ( .A(n182), .B(n18754), .Z(n18612) );
  AND U19345 ( .A(n18613), .B(n18612), .Z(n18761) );
  NAND U19346 ( .A(n189), .B(n18614), .Z(n18616) );
  XOR U19347 ( .A(b[17]), .B(a[124]), .Z(n18757) );
  NAND U19348 ( .A(n37652), .B(n18757), .Z(n18615) );
  NAND U19349 ( .A(n18616), .B(n18615), .Z(n18760) );
  XNOR U19350 ( .A(n18761), .B(n18760), .Z(n18762) );
  XOR U19351 ( .A(n18763), .B(n18762), .Z(n18797) );
  XOR U19352 ( .A(n18796), .B(n18797), .Z(n18799) );
  XOR U19353 ( .A(n18798), .B(n18799), .Z(n18731) );
  NANDN U19354 ( .A(n18618), .B(n18617), .Z(n18622) );
  NANDN U19355 ( .A(n18620), .B(n18619), .Z(n18621) );
  AND U19356 ( .A(n18622), .B(n18621), .Z(n18784) );
  NANDN U19357 ( .A(n18624), .B(n18623), .Z(n18628) );
  NANDN U19358 ( .A(n18626), .B(n18625), .Z(n18627) );
  NAND U19359 ( .A(n18628), .B(n18627), .Z(n18785) );
  XNOR U19360 ( .A(n18784), .B(n18785), .Z(n18786) );
  NANDN U19361 ( .A(n18630), .B(n18629), .Z(n18634) );
  NANDN U19362 ( .A(n18632), .B(n18631), .Z(n18633) );
  NAND U19363 ( .A(n18634), .B(n18633), .Z(n18787) );
  XNOR U19364 ( .A(n18786), .B(n18787), .Z(n18730) );
  XNOR U19365 ( .A(n18731), .B(n18730), .Z(n18733) );
  NANDN U19366 ( .A(n18636), .B(n18635), .Z(n18640) );
  NANDN U19367 ( .A(n18638), .B(n18637), .Z(n18639) );
  AND U19368 ( .A(n18640), .B(n18639), .Z(n18732) );
  XOR U19369 ( .A(n18733), .B(n18732), .Z(n18847) );
  NANDN U19370 ( .A(n18642), .B(n18641), .Z(n18646) );
  NANDN U19371 ( .A(n18644), .B(n18643), .Z(n18645) );
  AND U19372 ( .A(n18646), .B(n18645), .Z(n18844) );
  NANDN U19373 ( .A(n18648), .B(n18647), .Z(n18652) );
  NANDN U19374 ( .A(n18650), .B(n18649), .Z(n18651) );
  AND U19375 ( .A(n18652), .B(n18651), .Z(n18727) );
  NANDN U19376 ( .A(n18654), .B(n18653), .Z(n18658) );
  OR U19377 ( .A(n18656), .B(n18655), .Z(n18657) );
  AND U19378 ( .A(n18658), .B(n18657), .Z(n18725) );
  NANDN U19379 ( .A(n18660), .B(n18659), .Z(n18664) );
  NANDN U19380 ( .A(n18662), .B(n18661), .Z(n18663) );
  AND U19381 ( .A(n18664), .B(n18663), .Z(n18791) );
  NANDN U19382 ( .A(n18666), .B(n18665), .Z(n18670) );
  NANDN U19383 ( .A(n18668), .B(n18667), .Z(n18669) );
  NAND U19384 ( .A(n18670), .B(n18669), .Z(n18790) );
  XNOR U19385 ( .A(n18791), .B(n18790), .Z(n18792) );
  NAND U19386 ( .A(b[0]), .B(a[140]), .Z(n18671) );
  XNOR U19387 ( .A(b[1]), .B(n18671), .Z(n18673) );
  NANDN U19388 ( .A(b[0]), .B(a[139]), .Z(n18672) );
  NAND U19389 ( .A(n18673), .B(n18672), .Z(n18739) );
  NAND U19390 ( .A(n194), .B(n18674), .Z(n18676) );
  XOR U19391 ( .A(b[29]), .B(a[112]), .Z(n18817) );
  NAND U19392 ( .A(n38456), .B(n18817), .Z(n18675) );
  AND U19393 ( .A(n18676), .B(n18675), .Z(n18737) );
  AND U19394 ( .A(b[31]), .B(a[108]), .Z(n18736) );
  XNOR U19395 ( .A(n18737), .B(n18736), .Z(n18738) );
  XNOR U19396 ( .A(n18739), .B(n18738), .Z(n18778) );
  NAND U19397 ( .A(n38185), .B(n18677), .Z(n18679) );
  XOR U19398 ( .A(b[23]), .B(a[118]), .Z(n18820) );
  NAND U19399 ( .A(n38132), .B(n18820), .Z(n18678) );
  AND U19400 ( .A(n18679), .B(n18678), .Z(n18811) );
  NAND U19401 ( .A(n184), .B(n18680), .Z(n18682) );
  XOR U19402 ( .A(b[7]), .B(a[134]), .Z(n18823) );
  NAND U19403 ( .A(n36592), .B(n18823), .Z(n18681) );
  AND U19404 ( .A(n18682), .B(n18681), .Z(n18809) );
  NAND U19405 ( .A(n38289), .B(n18683), .Z(n18685) );
  XOR U19406 ( .A(b[25]), .B(a[116]), .Z(n18826) );
  NAND U19407 ( .A(n38247), .B(n18826), .Z(n18684) );
  NAND U19408 ( .A(n18685), .B(n18684), .Z(n18808) );
  XNOR U19409 ( .A(n18809), .B(n18808), .Z(n18810) );
  XOR U19410 ( .A(n18811), .B(n18810), .Z(n18779) );
  XNOR U19411 ( .A(n18778), .B(n18779), .Z(n18780) );
  NAND U19412 ( .A(n187), .B(n18686), .Z(n18688) );
  XOR U19413 ( .A(b[13]), .B(a[128]), .Z(n18829) );
  NAND U19414 ( .A(n37295), .B(n18829), .Z(n18687) );
  AND U19415 ( .A(n18688), .B(n18687), .Z(n18773) );
  NAND U19416 ( .A(n186), .B(n18689), .Z(n18691) );
  XOR U19417 ( .A(b[11]), .B(a[130]), .Z(n18832) );
  NAND U19418 ( .A(n37097), .B(n18832), .Z(n18690) );
  NAND U19419 ( .A(n18691), .B(n18690), .Z(n18772) );
  XNOR U19420 ( .A(n18773), .B(n18772), .Z(n18774) );
  NAND U19421 ( .A(n188), .B(n18692), .Z(n18694) );
  XOR U19422 ( .A(b[15]), .B(a[126]), .Z(n18835) );
  NAND U19423 ( .A(n37382), .B(n18835), .Z(n18693) );
  AND U19424 ( .A(n18694), .B(n18693), .Z(n18769) );
  NAND U19425 ( .A(n38064), .B(n18695), .Z(n18697) );
  XOR U19426 ( .A(b[21]), .B(a[120]), .Z(n18838) );
  NAND U19427 ( .A(n37993), .B(n18838), .Z(n18696) );
  AND U19428 ( .A(n18697), .B(n18696), .Z(n18767) );
  NAND U19429 ( .A(n185), .B(n18698), .Z(n18700) );
  XOR U19430 ( .A(b[9]), .B(a[132]), .Z(n18841) );
  NAND U19431 ( .A(n36805), .B(n18841), .Z(n18699) );
  NAND U19432 ( .A(n18700), .B(n18699), .Z(n18766) );
  XNOR U19433 ( .A(n18767), .B(n18766), .Z(n18768) );
  XOR U19434 ( .A(n18769), .B(n18768), .Z(n18775) );
  XOR U19435 ( .A(n18774), .B(n18775), .Z(n18781) );
  XOR U19436 ( .A(n18780), .B(n18781), .Z(n18793) );
  XNOR U19437 ( .A(n18792), .B(n18793), .Z(n18724) );
  XNOR U19438 ( .A(n18725), .B(n18724), .Z(n18726) );
  XOR U19439 ( .A(n18727), .B(n18726), .Z(n18845) );
  XNOR U19440 ( .A(n18844), .B(n18845), .Z(n18846) );
  XNOR U19441 ( .A(n18847), .B(n18846), .Z(n18852) );
  XOR U19442 ( .A(n18853), .B(n18852), .Z(n18719) );
  NANDN U19443 ( .A(n18702), .B(n18701), .Z(n18706) );
  NANDN U19444 ( .A(n18704), .B(n18703), .Z(n18705) );
  AND U19445 ( .A(n18706), .B(n18705), .Z(n18718) );
  XOR U19446 ( .A(n18719), .B(n18718), .Z(n18721) );
  XNOR U19447 ( .A(n18720), .B(n18721), .Z(n18712) );
  XNOR U19448 ( .A(n18713), .B(n18712), .Z(n18714) );
  XNOR U19449 ( .A(n18715), .B(n18714), .Z(n18856) );
  XNOR U19450 ( .A(sreg[364]), .B(n18856), .Z(n18858) );
  NANDN U19451 ( .A(sreg[363]), .B(n18707), .Z(n18711) );
  NAND U19452 ( .A(n18709), .B(n18708), .Z(n18710) );
  NAND U19453 ( .A(n18711), .B(n18710), .Z(n18857) );
  XNOR U19454 ( .A(n18858), .B(n18857), .Z(c[364]) );
  NANDN U19455 ( .A(n18713), .B(n18712), .Z(n18717) );
  NANDN U19456 ( .A(n18715), .B(n18714), .Z(n18716) );
  AND U19457 ( .A(n18717), .B(n18716), .Z(n18864) );
  NANDN U19458 ( .A(n18719), .B(n18718), .Z(n18723) );
  NANDN U19459 ( .A(n18721), .B(n18720), .Z(n18722) );
  AND U19460 ( .A(n18723), .B(n18722), .Z(n18862) );
  NANDN U19461 ( .A(n18725), .B(n18724), .Z(n18729) );
  NANDN U19462 ( .A(n18727), .B(n18726), .Z(n18728) );
  AND U19463 ( .A(n18729), .B(n18728), .Z(n18874) );
  NANDN U19464 ( .A(n18731), .B(n18730), .Z(n18735) );
  NAND U19465 ( .A(n18733), .B(n18732), .Z(n18734) );
  AND U19466 ( .A(n18735), .B(n18734), .Z(n18873) );
  XNOR U19467 ( .A(n18874), .B(n18873), .Z(n18876) );
  NANDN U19468 ( .A(n18737), .B(n18736), .Z(n18741) );
  NANDN U19469 ( .A(n18739), .B(n18738), .Z(n18740) );
  AND U19470 ( .A(n18741), .B(n18740), .Z(n18953) );
  NAND U19471 ( .A(n38385), .B(n18742), .Z(n18744) );
  XOR U19472 ( .A(b[27]), .B(a[115]), .Z(n18897) );
  NAND U19473 ( .A(n38343), .B(n18897), .Z(n18743) );
  AND U19474 ( .A(n18744), .B(n18743), .Z(n18960) );
  NAND U19475 ( .A(n183), .B(n18745), .Z(n18747) );
  XOR U19476 ( .A(b[5]), .B(a[137]), .Z(n18900) );
  NAND U19477 ( .A(n36296), .B(n18900), .Z(n18746) );
  AND U19478 ( .A(n18747), .B(n18746), .Z(n18958) );
  NAND U19479 ( .A(n190), .B(n18748), .Z(n18750) );
  XOR U19480 ( .A(b[19]), .B(a[123]), .Z(n18903) );
  NAND U19481 ( .A(n37821), .B(n18903), .Z(n18749) );
  NAND U19482 ( .A(n18750), .B(n18749), .Z(n18957) );
  XNOR U19483 ( .A(n18958), .B(n18957), .Z(n18959) );
  XNOR U19484 ( .A(n18960), .B(n18959), .Z(n18951) );
  NAND U19485 ( .A(n38470), .B(n18751), .Z(n18753) );
  XOR U19486 ( .A(b[31]), .B(a[111]), .Z(n18906) );
  NAND U19487 ( .A(n38453), .B(n18906), .Z(n18752) );
  AND U19488 ( .A(n18753), .B(n18752), .Z(n18918) );
  NAND U19489 ( .A(n181), .B(n18754), .Z(n18756) );
  XOR U19490 ( .A(b[3]), .B(a[139]), .Z(n18909) );
  NAND U19491 ( .A(n182), .B(n18909), .Z(n18755) );
  AND U19492 ( .A(n18756), .B(n18755), .Z(n18916) );
  NAND U19493 ( .A(n189), .B(n18757), .Z(n18759) );
  XOR U19494 ( .A(b[17]), .B(a[125]), .Z(n18912) );
  NAND U19495 ( .A(n37652), .B(n18912), .Z(n18758) );
  NAND U19496 ( .A(n18759), .B(n18758), .Z(n18915) );
  XNOR U19497 ( .A(n18916), .B(n18915), .Z(n18917) );
  XOR U19498 ( .A(n18918), .B(n18917), .Z(n18952) );
  XOR U19499 ( .A(n18951), .B(n18952), .Z(n18954) );
  XOR U19500 ( .A(n18953), .B(n18954), .Z(n18886) );
  NANDN U19501 ( .A(n18761), .B(n18760), .Z(n18765) );
  NANDN U19502 ( .A(n18763), .B(n18762), .Z(n18764) );
  AND U19503 ( .A(n18765), .B(n18764), .Z(n18939) );
  NANDN U19504 ( .A(n18767), .B(n18766), .Z(n18771) );
  NANDN U19505 ( .A(n18769), .B(n18768), .Z(n18770) );
  NAND U19506 ( .A(n18771), .B(n18770), .Z(n18940) );
  XNOR U19507 ( .A(n18939), .B(n18940), .Z(n18941) );
  NANDN U19508 ( .A(n18773), .B(n18772), .Z(n18777) );
  NANDN U19509 ( .A(n18775), .B(n18774), .Z(n18776) );
  NAND U19510 ( .A(n18777), .B(n18776), .Z(n18942) );
  XNOR U19511 ( .A(n18941), .B(n18942), .Z(n18885) );
  XNOR U19512 ( .A(n18886), .B(n18885), .Z(n18888) );
  NANDN U19513 ( .A(n18779), .B(n18778), .Z(n18783) );
  NANDN U19514 ( .A(n18781), .B(n18780), .Z(n18782) );
  AND U19515 ( .A(n18783), .B(n18782), .Z(n18887) );
  XOR U19516 ( .A(n18888), .B(n18887), .Z(n19002) );
  NANDN U19517 ( .A(n18785), .B(n18784), .Z(n18789) );
  NANDN U19518 ( .A(n18787), .B(n18786), .Z(n18788) );
  AND U19519 ( .A(n18789), .B(n18788), .Z(n18999) );
  NANDN U19520 ( .A(n18791), .B(n18790), .Z(n18795) );
  NANDN U19521 ( .A(n18793), .B(n18792), .Z(n18794) );
  AND U19522 ( .A(n18795), .B(n18794), .Z(n18882) );
  NANDN U19523 ( .A(n18797), .B(n18796), .Z(n18801) );
  OR U19524 ( .A(n18799), .B(n18798), .Z(n18800) );
  AND U19525 ( .A(n18801), .B(n18800), .Z(n18880) );
  NANDN U19526 ( .A(n18803), .B(n18802), .Z(n18807) );
  NANDN U19527 ( .A(n18805), .B(n18804), .Z(n18806) );
  AND U19528 ( .A(n18807), .B(n18806), .Z(n18946) );
  NANDN U19529 ( .A(n18809), .B(n18808), .Z(n18813) );
  NANDN U19530 ( .A(n18811), .B(n18810), .Z(n18812) );
  NAND U19531 ( .A(n18813), .B(n18812), .Z(n18945) );
  XNOR U19532 ( .A(n18946), .B(n18945), .Z(n18947) );
  NAND U19533 ( .A(b[0]), .B(a[141]), .Z(n18814) );
  XNOR U19534 ( .A(b[1]), .B(n18814), .Z(n18816) );
  NANDN U19535 ( .A(b[0]), .B(a[140]), .Z(n18815) );
  NAND U19536 ( .A(n18816), .B(n18815), .Z(n18894) );
  NAND U19537 ( .A(n194), .B(n18817), .Z(n18819) );
  XOR U19538 ( .A(b[29]), .B(a[113]), .Z(n18972) );
  NAND U19539 ( .A(n38456), .B(n18972), .Z(n18818) );
  AND U19540 ( .A(n18819), .B(n18818), .Z(n18892) );
  AND U19541 ( .A(b[31]), .B(a[109]), .Z(n18891) );
  XNOR U19542 ( .A(n18892), .B(n18891), .Z(n18893) );
  XNOR U19543 ( .A(n18894), .B(n18893), .Z(n18933) );
  NAND U19544 ( .A(n38185), .B(n18820), .Z(n18822) );
  XOR U19545 ( .A(b[23]), .B(a[119]), .Z(n18975) );
  NAND U19546 ( .A(n38132), .B(n18975), .Z(n18821) );
  AND U19547 ( .A(n18822), .B(n18821), .Z(n18966) );
  NAND U19548 ( .A(n184), .B(n18823), .Z(n18825) );
  XOR U19549 ( .A(b[7]), .B(a[135]), .Z(n18978) );
  NAND U19550 ( .A(n36592), .B(n18978), .Z(n18824) );
  AND U19551 ( .A(n18825), .B(n18824), .Z(n18964) );
  NAND U19552 ( .A(n38289), .B(n18826), .Z(n18828) );
  XOR U19553 ( .A(b[25]), .B(a[117]), .Z(n18981) );
  NAND U19554 ( .A(n38247), .B(n18981), .Z(n18827) );
  NAND U19555 ( .A(n18828), .B(n18827), .Z(n18963) );
  XNOR U19556 ( .A(n18964), .B(n18963), .Z(n18965) );
  XOR U19557 ( .A(n18966), .B(n18965), .Z(n18934) );
  XNOR U19558 ( .A(n18933), .B(n18934), .Z(n18935) );
  NAND U19559 ( .A(n187), .B(n18829), .Z(n18831) );
  XOR U19560 ( .A(b[13]), .B(a[129]), .Z(n18984) );
  NAND U19561 ( .A(n37295), .B(n18984), .Z(n18830) );
  AND U19562 ( .A(n18831), .B(n18830), .Z(n18928) );
  NAND U19563 ( .A(n186), .B(n18832), .Z(n18834) );
  XOR U19564 ( .A(b[11]), .B(a[131]), .Z(n18987) );
  NAND U19565 ( .A(n37097), .B(n18987), .Z(n18833) );
  NAND U19566 ( .A(n18834), .B(n18833), .Z(n18927) );
  XNOR U19567 ( .A(n18928), .B(n18927), .Z(n18929) );
  NAND U19568 ( .A(n188), .B(n18835), .Z(n18837) );
  XOR U19569 ( .A(b[15]), .B(a[127]), .Z(n18990) );
  NAND U19570 ( .A(n37382), .B(n18990), .Z(n18836) );
  AND U19571 ( .A(n18837), .B(n18836), .Z(n18924) );
  NAND U19572 ( .A(n38064), .B(n18838), .Z(n18840) );
  XOR U19573 ( .A(b[21]), .B(a[121]), .Z(n18993) );
  NAND U19574 ( .A(n37993), .B(n18993), .Z(n18839) );
  AND U19575 ( .A(n18840), .B(n18839), .Z(n18922) );
  NAND U19576 ( .A(n185), .B(n18841), .Z(n18843) );
  XOR U19577 ( .A(b[9]), .B(a[133]), .Z(n18996) );
  NAND U19578 ( .A(n36805), .B(n18996), .Z(n18842) );
  NAND U19579 ( .A(n18843), .B(n18842), .Z(n18921) );
  XNOR U19580 ( .A(n18922), .B(n18921), .Z(n18923) );
  XOR U19581 ( .A(n18924), .B(n18923), .Z(n18930) );
  XOR U19582 ( .A(n18929), .B(n18930), .Z(n18936) );
  XOR U19583 ( .A(n18935), .B(n18936), .Z(n18948) );
  XNOR U19584 ( .A(n18947), .B(n18948), .Z(n18879) );
  XNOR U19585 ( .A(n18880), .B(n18879), .Z(n18881) );
  XOR U19586 ( .A(n18882), .B(n18881), .Z(n19000) );
  XNOR U19587 ( .A(n18999), .B(n19000), .Z(n19001) );
  XNOR U19588 ( .A(n19002), .B(n19001), .Z(n18875) );
  XOR U19589 ( .A(n18876), .B(n18875), .Z(n18868) );
  NANDN U19590 ( .A(n18845), .B(n18844), .Z(n18849) );
  NANDN U19591 ( .A(n18847), .B(n18846), .Z(n18848) );
  AND U19592 ( .A(n18849), .B(n18848), .Z(n18867) );
  XNOR U19593 ( .A(n18868), .B(n18867), .Z(n18869) );
  NANDN U19594 ( .A(n18851), .B(n18850), .Z(n18855) );
  NAND U19595 ( .A(n18853), .B(n18852), .Z(n18854) );
  NAND U19596 ( .A(n18855), .B(n18854), .Z(n18870) );
  XNOR U19597 ( .A(n18869), .B(n18870), .Z(n18861) );
  XNOR U19598 ( .A(n18862), .B(n18861), .Z(n18863) );
  XNOR U19599 ( .A(n18864), .B(n18863), .Z(n19005) );
  XNOR U19600 ( .A(sreg[365]), .B(n19005), .Z(n19007) );
  NANDN U19601 ( .A(sreg[364]), .B(n18856), .Z(n18860) );
  NAND U19602 ( .A(n18858), .B(n18857), .Z(n18859) );
  NAND U19603 ( .A(n18860), .B(n18859), .Z(n19006) );
  XNOR U19604 ( .A(n19007), .B(n19006), .Z(c[365]) );
  NANDN U19605 ( .A(n18862), .B(n18861), .Z(n18866) );
  NANDN U19606 ( .A(n18864), .B(n18863), .Z(n18865) );
  AND U19607 ( .A(n18866), .B(n18865), .Z(n19013) );
  NANDN U19608 ( .A(n18868), .B(n18867), .Z(n18872) );
  NANDN U19609 ( .A(n18870), .B(n18869), .Z(n18871) );
  AND U19610 ( .A(n18872), .B(n18871), .Z(n19011) );
  NANDN U19611 ( .A(n18874), .B(n18873), .Z(n18878) );
  NAND U19612 ( .A(n18876), .B(n18875), .Z(n18877) );
  AND U19613 ( .A(n18878), .B(n18877), .Z(n19018) );
  NANDN U19614 ( .A(n18880), .B(n18879), .Z(n18884) );
  NANDN U19615 ( .A(n18882), .B(n18881), .Z(n18883) );
  AND U19616 ( .A(n18884), .B(n18883), .Z(n19023) );
  NANDN U19617 ( .A(n18886), .B(n18885), .Z(n18890) );
  NAND U19618 ( .A(n18888), .B(n18887), .Z(n18889) );
  AND U19619 ( .A(n18890), .B(n18889), .Z(n19022) );
  XNOR U19620 ( .A(n19023), .B(n19022), .Z(n19025) );
  NANDN U19621 ( .A(n18892), .B(n18891), .Z(n18896) );
  NANDN U19622 ( .A(n18894), .B(n18893), .Z(n18895) );
  AND U19623 ( .A(n18896), .B(n18895), .Z(n19100) );
  NAND U19624 ( .A(n38385), .B(n18897), .Z(n18899) );
  XOR U19625 ( .A(b[27]), .B(a[116]), .Z(n19046) );
  NAND U19626 ( .A(n38343), .B(n19046), .Z(n18898) );
  AND U19627 ( .A(n18899), .B(n18898), .Z(n19107) );
  NAND U19628 ( .A(n183), .B(n18900), .Z(n18902) );
  XOR U19629 ( .A(b[5]), .B(a[138]), .Z(n19049) );
  NAND U19630 ( .A(n36296), .B(n19049), .Z(n18901) );
  AND U19631 ( .A(n18902), .B(n18901), .Z(n19105) );
  NAND U19632 ( .A(n190), .B(n18903), .Z(n18905) );
  XOR U19633 ( .A(b[19]), .B(a[124]), .Z(n19052) );
  NAND U19634 ( .A(n37821), .B(n19052), .Z(n18904) );
  NAND U19635 ( .A(n18905), .B(n18904), .Z(n19104) );
  XNOR U19636 ( .A(n19105), .B(n19104), .Z(n19106) );
  XNOR U19637 ( .A(n19107), .B(n19106), .Z(n19098) );
  NAND U19638 ( .A(n38470), .B(n18906), .Z(n18908) );
  XOR U19639 ( .A(b[31]), .B(a[112]), .Z(n19055) );
  NAND U19640 ( .A(n38453), .B(n19055), .Z(n18907) );
  AND U19641 ( .A(n18908), .B(n18907), .Z(n19067) );
  NAND U19642 ( .A(n181), .B(n18909), .Z(n18911) );
  XOR U19643 ( .A(b[3]), .B(a[140]), .Z(n19058) );
  NAND U19644 ( .A(n182), .B(n19058), .Z(n18910) );
  AND U19645 ( .A(n18911), .B(n18910), .Z(n19065) );
  NAND U19646 ( .A(n189), .B(n18912), .Z(n18914) );
  XOR U19647 ( .A(b[17]), .B(a[126]), .Z(n19061) );
  NAND U19648 ( .A(n37652), .B(n19061), .Z(n18913) );
  NAND U19649 ( .A(n18914), .B(n18913), .Z(n19064) );
  XNOR U19650 ( .A(n19065), .B(n19064), .Z(n19066) );
  XOR U19651 ( .A(n19067), .B(n19066), .Z(n19099) );
  XOR U19652 ( .A(n19098), .B(n19099), .Z(n19101) );
  XOR U19653 ( .A(n19100), .B(n19101), .Z(n19035) );
  NANDN U19654 ( .A(n18916), .B(n18915), .Z(n18920) );
  NANDN U19655 ( .A(n18918), .B(n18917), .Z(n18919) );
  AND U19656 ( .A(n18920), .B(n18919), .Z(n19088) );
  NANDN U19657 ( .A(n18922), .B(n18921), .Z(n18926) );
  NANDN U19658 ( .A(n18924), .B(n18923), .Z(n18925) );
  NAND U19659 ( .A(n18926), .B(n18925), .Z(n19089) );
  XNOR U19660 ( .A(n19088), .B(n19089), .Z(n19090) );
  NANDN U19661 ( .A(n18928), .B(n18927), .Z(n18932) );
  NANDN U19662 ( .A(n18930), .B(n18929), .Z(n18931) );
  NAND U19663 ( .A(n18932), .B(n18931), .Z(n19091) );
  XNOR U19664 ( .A(n19090), .B(n19091), .Z(n19034) );
  XNOR U19665 ( .A(n19035), .B(n19034), .Z(n19037) );
  NANDN U19666 ( .A(n18934), .B(n18933), .Z(n18938) );
  NANDN U19667 ( .A(n18936), .B(n18935), .Z(n18937) );
  AND U19668 ( .A(n18938), .B(n18937), .Z(n19036) );
  XOR U19669 ( .A(n19037), .B(n19036), .Z(n19149) );
  NANDN U19670 ( .A(n18940), .B(n18939), .Z(n18944) );
  NANDN U19671 ( .A(n18942), .B(n18941), .Z(n18943) );
  AND U19672 ( .A(n18944), .B(n18943), .Z(n19146) );
  NANDN U19673 ( .A(n18946), .B(n18945), .Z(n18950) );
  NANDN U19674 ( .A(n18948), .B(n18947), .Z(n18949) );
  AND U19675 ( .A(n18950), .B(n18949), .Z(n19031) );
  NANDN U19676 ( .A(n18952), .B(n18951), .Z(n18956) );
  OR U19677 ( .A(n18954), .B(n18953), .Z(n18955) );
  AND U19678 ( .A(n18956), .B(n18955), .Z(n19029) );
  NANDN U19679 ( .A(n18958), .B(n18957), .Z(n18962) );
  NANDN U19680 ( .A(n18960), .B(n18959), .Z(n18961) );
  AND U19681 ( .A(n18962), .B(n18961), .Z(n19095) );
  NANDN U19682 ( .A(n18964), .B(n18963), .Z(n18968) );
  NANDN U19683 ( .A(n18966), .B(n18965), .Z(n18967) );
  NAND U19684 ( .A(n18968), .B(n18967), .Z(n19094) );
  XNOR U19685 ( .A(n19095), .B(n19094), .Z(n19097) );
  NAND U19686 ( .A(b[0]), .B(a[142]), .Z(n18969) );
  XNOR U19687 ( .A(b[1]), .B(n18969), .Z(n18971) );
  NANDN U19688 ( .A(b[0]), .B(a[141]), .Z(n18970) );
  NAND U19689 ( .A(n18971), .B(n18970), .Z(n19043) );
  NAND U19690 ( .A(n194), .B(n18972), .Z(n18974) );
  XOR U19691 ( .A(b[29]), .B(a[114]), .Z(n19116) );
  NAND U19692 ( .A(n38456), .B(n19116), .Z(n18973) );
  AND U19693 ( .A(n18974), .B(n18973), .Z(n19041) );
  AND U19694 ( .A(b[31]), .B(a[110]), .Z(n19040) );
  XNOR U19695 ( .A(n19041), .B(n19040), .Z(n19042) );
  XNOR U19696 ( .A(n19043), .B(n19042), .Z(n19083) );
  NAND U19697 ( .A(n38185), .B(n18975), .Z(n18977) );
  XOR U19698 ( .A(b[23]), .B(a[120]), .Z(n19122) );
  NAND U19699 ( .A(n38132), .B(n19122), .Z(n18976) );
  AND U19700 ( .A(n18977), .B(n18976), .Z(n19112) );
  NAND U19701 ( .A(n184), .B(n18978), .Z(n18980) );
  XOR U19702 ( .A(b[7]), .B(a[136]), .Z(n19125) );
  NAND U19703 ( .A(n36592), .B(n19125), .Z(n18979) );
  AND U19704 ( .A(n18980), .B(n18979), .Z(n19111) );
  NAND U19705 ( .A(n38289), .B(n18981), .Z(n18983) );
  XOR U19706 ( .A(b[25]), .B(a[118]), .Z(n19128) );
  NAND U19707 ( .A(n38247), .B(n19128), .Z(n18982) );
  NAND U19708 ( .A(n18983), .B(n18982), .Z(n19110) );
  XOR U19709 ( .A(n19111), .B(n19110), .Z(n19113) );
  XOR U19710 ( .A(n19112), .B(n19113), .Z(n19082) );
  XOR U19711 ( .A(n19083), .B(n19082), .Z(n19085) );
  NAND U19712 ( .A(n187), .B(n18984), .Z(n18986) );
  XOR U19713 ( .A(b[13]), .B(a[130]), .Z(n19131) );
  NAND U19714 ( .A(n37295), .B(n19131), .Z(n18985) );
  AND U19715 ( .A(n18986), .B(n18985), .Z(n19077) );
  NAND U19716 ( .A(n186), .B(n18987), .Z(n18989) );
  XOR U19717 ( .A(b[11]), .B(a[132]), .Z(n19134) );
  NAND U19718 ( .A(n37097), .B(n19134), .Z(n18988) );
  NAND U19719 ( .A(n18989), .B(n18988), .Z(n19076) );
  XNOR U19720 ( .A(n19077), .B(n19076), .Z(n19079) );
  NAND U19721 ( .A(n188), .B(n18990), .Z(n18992) );
  XOR U19722 ( .A(b[15]), .B(a[128]), .Z(n19137) );
  NAND U19723 ( .A(n37382), .B(n19137), .Z(n18991) );
  AND U19724 ( .A(n18992), .B(n18991), .Z(n19073) );
  NAND U19725 ( .A(n38064), .B(n18993), .Z(n18995) );
  XOR U19726 ( .A(b[21]), .B(a[122]), .Z(n19140) );
  NAND U19727 ( .A(n37993), .B(n19140), .Z(n18994) );
  AND U19728 ( .A(n18995), .B(n18994), .Z(n19071) );
  NAND U19729 ( .A(n185), .B(n18996), .Z(n18998) );
  XOR U19730 ( .A(b[9]), .B(a[134]), .Z(n19143) );
  NAND U19731 ( .A(n36805), .B(n19143), .Z(n18997) );
  NAND U19732 ( .A(n18998), .B(n18997), .Z(n19070) );
  XNOR U19733 ( .A(n19071), .B(n19070), .Z(n19072) );
  XNOR U19734 ( .A(n19073), .B(n19072), .Z(n19078) );
  XOR U19735 ( .A(n19079), .B(n19078), .Z(n19084) );
  XNOR U19736 ( .A(n19085), .B(n19084), .Z(n19096) );
  XNOR U19737 ( .A(n19097), .B(n19096), .Z(n19028) );
  XNOR U19738 ( .A(n19029), .B(n19028), .Z(n19030) );
  XOR U19739 ( .A(n19031), .B(n19030), .Z(n19147) );
  XNOR U19740 ( .A(n19146), .B(n19147), .Z(n19148) );
  XNOR U19741 ( .A(n19149), .B(n19148), .Z(n19024) );
  XOR U19742 ( .A(n19025), .B(n19024), .Z(n19017) );
  NANDN U19743 ( .A(n19000), .B(n18999), .Z(n19004) );
  NANDN U19744 ( .A(n19002), .B(n19001), .Z(n19003) );
  AND U19745 ( .A(n19004), .B(n19003), .Z(n19016) );
  XOR U19746 ( .A(n19017), .B(n19016), .Z(n19019) );
  XNOR U19747 ( .A(n19018), .B(n19019), .Z(n19010) );
  XNOR U19748 ( .A(n19011), .B(n19010), .Z(n19012) );
  XNOR U19749 ( .A(n19013), .B(n19012), .Z(n19152) );
  XNOR U19750 ( .A(sreg[366]), .B(n19152), .Z(n19154) );
  NANDN U19751 ( .A(sreg[365]), .B(n19005), .Z(n19009) );
  NAND U19752 ( .A(n19007), .B(n19006), .Z(n19008) );
  NAND U19753 ( .A(n19009), .B(n19008), .Z(n19153) );
  XNOR U19754 ( .A(n19154), .B(n19153), .Z(c[366]) );
  NANDN U19755 ( .A(n19011), .B(n19010), .Z(n19015) );
  NANDN U19756 ( .A(n19013), .B(n19012), .Z(n19014) );
  AND U19757 ( .A(n19015), .B(n19014), .Z(n19160) );
  NANDN U19758 ( .A(n19017), .B(n19016), .Z(n19021) );
  NANDN U19759 ( .A(n19019), .B(n19018), .Z(n19020) );
  AND U19760 ( .A(n19021), .B(n19020), .Z(n19158) );
  NANDN U19761 ( .A(n19023), .B(n19022), .Z(n19027) );
  NAND U19762 ( .A(n19025), .B(n19024), .Z(n19026) );
  AND U19763 ( .A(n19027), .B(n19026), .Z(n19165) );
  NANDN U19764 ( .A(n19029), .B(n19028), .Z(n19033) );
  NANDN U19765 ( .A(n19031), .B(n19030), .Z(n19032) );
  AND U19766 ( .A(n19033), .B(n19032), .Z(n19170) );
  NANDN U19767 ( .A(n19035), .B(n19034), .Z(n19039) );
  NAND U19768 ( .A(n19037), .B(n19036), .Z(n19038) );
  AND U19769 ( .A(n19039), .B(n19038), .Z(n19169) );
  XNOR U19770 ( .A(n19170), .B(n19169), .Z(n19172) );
  NANDN U19771 ( .A(n19041), .B(n19040), .Z(n19045) );
  NANDN U19772 ( .A(n19043), .B(n19042), .Z(n19044) );
  AND U19773 ( .A(n19045), .B(n19044), .Z(n19237) );
  NAND U19774 ( .A(n38385), .B(n19046), .Z(n19048) );
  XOR U19775 ( .A(b[27]), .B(a[117]), .Z(n19181) );
  NAND U19776 ( .A(n38343), .B(n19181), .Z(n19047) );
  AND U19777 ( .A(n19048), .B(n19047), .Z(n19244) );
  NAND U19778 ( .A(n183), .B(n19049), .Z(n19051) );
  XOR U19779 ( .A(b[5]), .B(a[139]), .Z(n19184) );
  NAND U19780 ( .A(n36296), .B(n19184), .Z(n19050) );
  AND U19781 ( .A(n19051), .B(n19050), .Z(n19242) );
  NAND U19782 ( .A(n190), .B(n19052), .Z(n19054) );
  XOR U19783 ( .A(b[19]), .B(a[125]), .Z(n19187) );
  NAND U19784 ( .A(n37821), .B(n19187), .Z(n19053) );
  NAND U19785 ( .A(n19054), .B(n19053), .Z(n19241) );
  XNOR U19786 ( .A(n19242), .B(n19241), .Z(n19243) );
  XNOR U19787 ( .A(n19244), .B(n19243), .Z(n19235) );
  NAND U19788 ( .A(n38470), .B(n19055), .Z(n19057) );
  XOR U19789 ( .A(b[31]), .B(a[113]), .Z(n19190) );
  NAND U19790 ( .A(n38453), .B(n19190), .Z(n19056) );
  AND U19791 ( .A(n19057), .B(n19056), .Z(n19202) );
  NAND U19792 ( .A(n181), .B(n19058), .Z(n19060) );
  XOR U19793 ( .A(b[3]), .B(a[141]), .Z(n19193) );
  NAND U19794 ( .A(n182), .B(n19193), .Z(n19059) );
  AND U19795 ( .A(n19060), .B(n19059), .Z(n19200) );
  NAND U19796 ( .A(n189), .B(n19061), .Z(n19063) );
  XOR U19797 ( .A(b[17]), .B(a[127]), .Z(n19196) );
  NAND U19798 ( .A(n37652), .B(n19196), .Z(n19062) );
  NAND U19799 ( .A(n19063), .B(n19062), .Z(n19199) );
  XNOR U19800 ( .A(n19200), .B(n19199), .Z(n19201) );
  XOR U19801 ( .A(n19202), .B(n19201), .Z(n19236) );
  XOR U19802 ( .A(n19235), .B(n19236), .Z(n19238) );
  XOR U19803 ( .A(n19237), .B(n19238), .Z(n19284) );
  NANDN U19804 ( .A(n19065), .B(n19064), .Z(n19069) );
  NANDN U19805 ( .A(n19067), .B(n19066), .Z(n19068) );
  AND U19806 ( .A(n19069), .B(n19068), .Z(n19223) );
  NANDN U19807 ( .A(n19071), .B(n19070), .Z(n19075) );
  NANDN U19808 ( .A(n19073), .B(n19072), .Z(n19074) );
  NAND U19809 ( .A(n19075), .B(n19074), .Z(n19224) );
  XNOR U19810 ( .A(n19223), .B(n19224), .Z(n19225) );
  NANDN U19811 ( .A(n19077), .B(n19076), .Z(n19081) );
  NAND U19812 ( .A(n19079), .B(n19078), .Z(n19080) );
  NAND U19813 ( .A(n19081), .B(n19080), .Z(n19226) );
  XNOR U19814 ( .A(n19225), .B(n19226), .Z(n19283) );
  XNOR U19815 ( .A(n19284), .B(n19283), .Z(n19286) );
  NAND U19816 ( .A(n19083), .B(n19082), .Z(n19087) );
  NAND U19817 ( .A(n19085), .B(n19084), .Z(n19086) );
  AND U19818 ( .A(n19087), .B(n19086), .Z(n19285) );
  XOR U19819 ( .A(n19286), .B(n19285), .Z(n19298) );
  NANDN U19820 ( .A(n19089), .B(n19088), .Z(n19093) );
  NANDN U19821 ( .A(n19091), .B(n19090), .Z(n19092) );
  AND U19822 ( .A(n19093), .B(n19092), .Z(n19295) );
  NANDN U19823 ( .A(n19099), .B(n19098), .Z(n19103) );
  OR U19824 ( .A(n19101), .B(n19100), .Z(n19102) );
  AND U19825 ( .A(n19103), .B(n19102), .Z(n19290) );
  NANDN U19826 ( .A(n19105), .B(n19104), .Z(n19109) );
  NANDN U19827 ( .A(n19107), .B(n19106), .Z(n19108) );
  AND U19828 ( .A(n19109), .B(n19108), .Z(n19230) );
  NANDN U19829 ( .A(n19111), .B(n19110), .Z(n19115) );
  OR U19830 ( .A(n19113), .B(n19112), .Z(n19114) );
  NAND U19831 ( .A(n19115), .B(n19114), .Z(n19229) );
  XNOR U19832 ( .A(n19230), .B(n19229), .Z(n19231) );
  NAND U19833 ( .A(n194), .B(n19116), .Z(n19118) );
  XOR U19834 ( .A(b[29]), .B(a[115]), .Z(n19256) );
  NAND U19835 ( .A(n38456), .B(n19256), .Z(n19117) );
  AND U19836 ( .A(n19118), .B(n19117), .Z(n19176) );
  AND U19837 ( .A(b[31]), .B(a[111]), .Z(n19175) );
  XNOR U19838 ( .A(n19176), .B(n19175), .Z(n19177) );
  NAND U19839 ( .A(b[0]), .B(a[143]), .Z(n19119) );
  XNOR U19840 ( .A(b[1]), .B(n19119), .Z(n19121) );
  NANDN U19841 ( .A(b[0]), .B(a[142]), .Z(n19120) );
  NAND U19842 ( .A(n19121), .B(n19120), .Z(n19178) );
  XNOR U19843 ( .A(n19177), .B(n19178), .Z(n19217) );
  NAND U19844 ( .A(n38185), .B(n19122), .Z(n19124) );
  XOR U19845 ( .A(b[23]), .B(a[121]), .Z(n19259) );
  NAND U19846 ( .A(n38132), .B(n19259), .Z(n19123) );
  AND U19847 ( .A(n19124), .B(n19123), .Z(n19250) );
  NAND U19848 ( .A(n184), .B(n19125), .Z(n19127) );
  XOR U19849 ( .A(b[7]), .B(a[137]), .Z(n19262) );
  NAND U19850 ( .A(n36592), .B(n19262), .Z(n19126) );
  AND U19851 ( .A(n19127), .B(n19126), .Z(n19248) );
  NAND U19852 ( .A(n38289), .B(n19128), .Z(n19130) );
  XOR U19853 ( .A(b[25]), .B(a[119]), .Z(n19265) );
  NAND U19854 ( .A(n38247), .B(n19265), .Z(n19129) );
  NAND U19855 ( .A(n19130), .B(n19129), .Z(n19247) );
  XNOR U19856 ( .A(n19248), .B(n19247), .Z(n19249) );
  XOR U19857 ( .A(n19250), .B(n19249), .Z(n19218) );
  XNOR U19858 ( .A(n19217), .B(n19218), .Z(n19219) );
  NAND U19859 ( .A(n187), .B(n19131), .Z(n19133) );
  XOR U19860 ( .A(b[13]), .B(a[131]), .Z(n19268) );
  NAND U19861 ( .A(n37295), .B(n19268), .Z(n19132) );
  AND U19862 ( .A(n19133), .B(n19132), .Z(n19212) );
  NAND U19863 ( .A(n186), .B(n19134), .Z(n19136) );
  XOR U19864 ( .A(b[11]), .B(a[133]), .Z(n19271) );
  NAND U19865 ( .A(n37097), .B(n19271), .Z(n19135) );
  NAND U19866 ( .A(n19136), .B(n19135), .Z(n19211) );
  XNOR U19867 ( .A(n19212), .B(n19211), .Z(n19213) );
  NAND U19868 ( .A(n188), .B(n19137), .Z(n19139) );
  XOR U19869 ( .A(b[15]), .B(a[129]), .Z(n19274) );
  NAND U19870 ( .A(n37382), .B(n19274), .Z(n19138) );
  AND U19871 ( .A(n19139), .B(n19138), .Z(n19208) );
  NAND U19872 ( .A(n38064), .B(n19140), .Z(n19142) );
  XOR U19873 ( .A(b[21]), .B(a[123]), .Z(n19277) );
  NAND U19874 ( .A(n37993), .B(n19277), .Z(n19141) );
  AND U19875 ( .A(n19142), .B(n19141), .Z(n19206) );
  NAND U19876 ( .A(n185), .B(n19143), .Z(n19145) );
  XOR U19877 ( .A(b[9]), .B(a[135]), .Z(n19280) );
  NAND U19878 ( .A(n36805), .B(n19280), .Z(n19144) );
  NAND U19879 ( .A(n19145), .B(n19144), .Z(n19205) );
  XNOR U19880 ( .A(n19206), .B(n19205), .Z(n19207) );
  XOR U19881 ( .A(n19208), .B(n19207), .Z(n19214) );
  XOR U19882 ( .A(n19213), .B(n19214), .Z(n19220) );
  XOR U19883 ( .A(n19219), .B(n19220), .Z(n19232) );
  XNOR U19884 ( .A(n19231), .B(n19232), .Z(n19289) );
  XNOR U19885 ( .A(n19290), .B(n19289), .Z(n19291) );
  XOR U19886 ( .A(n19292), .B(n19291), .Z(n19296) );
  XNOR U19887 ( .A(n19295), .B(n19296), .Z(n19297) );
  XNOR U19888 ( .A(n19298), .B(n19297), .Z(n19171) );
  XOR U19889 ( .A(n19172), .B(n19171), .Z(n19164) );
  NANDN U19890 ( .A(n19147), .B(n19146), .Z(n19151) );
  NANDN U19891 ( .A(n19149), .B(n19148), .Z(n19150) );
  AND U19892 ( .A(n19151), .B(n19150), .Z(n19163) );
  XOR U19893 ( .A(n19164), .B(n19163), .Z(n19166) );
  XNOR U19894 ( .A(n19165), .B(n19166), .Z(n19157) );
  XNOR U19895 ( .A(n19158), .B(n19157), .Z(n19159) );
  XNOR U19896 ( .A(n19160), .B(n19159), .Z(n19301) );
  XNOR U19897 ( .A(sreg[367]), .B(n19301), .Z(n19303) );
  NANDN U19898 ( .A(sreg[366]), .B(n19152), .Z(n19156) );
  NAND U19899 ( .A(n19154), .B(n19153), .Z(n19155) );
  NAND U19900 ( .A(n19156), .B(n19155), .Z(n19302) );
  XNOR U19901 ( .A(n19303), .B(n19302), .Z(c[367]) );
  NANDN U19902 ( .A(n19158), .B(n19157), .Z(n19162) );
  NANDN U19903 ( .A(n19160), .B(n19159), .Z(n19161) );
  AND U19904 ( .A(n19162), .B(n19161), .Z(n19309) );
  NANDN U19905 ( .A(n19164), .B(n19163), .Z(n19168) );
  NANDN U19906 ( .A(n19166), .B(n19165), .Z(n19167) );
  AND U19907 ( .A(n19168), .B(n19167), .Z(n19307) );
  NANDN U19908 ( .A(n19170), .B(n19169), .Z(n19174) );
  NAND U19909 ( .A(n19172), .B(n19171), .Z(n19173) );
  AND U19910 ( .A(n19174), .B(n19173), .Z(n19314) );
  NANDN U19911 ( .A(n19176), .B(n19175), .Z(n19180) );
  NANDN U19912 ( .A(n19178), .B(n19177), .Z(n19179) );
  AND U19913 ( .A(n19180), .B(n19179), .Z(n19396) );
  NAND U19914 ( .A(n38385), .B(n19181), .Z(n19183) );
  XOR U19915 ( .A(b[27]), .B(a[118]), .Z(n19342) );
  NAND U19916 ( .A(n38343), .B(n19342), .Z(n19182) );
  AND U19917 ( .A(n19183), .B(n19182), .Z(n19403) );
  NAND U19918 ( .A(n183), .B(n19184), .Z(n19186) );
  XOR U19919 ( .A(b[5]), .B(a[140]), .Z(n19345) );
  NAND U19920 ( .A(n36296), .B(n19345), .Z(n19185) );
  AND U19921 ( .A(n19186), .B(n19185), .Z(n19401) );
  NAND U19922 ( .A(n190), .B(n19187), .Z(n19189) );
  XOR U19923 ( .A(b[19]), .B(a[126]), .Z(n19348) );
  NAND U19924 ( .A(n37821), .B(n19348), .Z(n19188) );
  NAND U19925 ( .A(n19189), .B(n19188), .Z(n19400) );
  XNOR U19926 ( .A(n19401), .B(n19400), .Z(n19402) );
  XNOR U19927 ( .A(n19403), .B(n19402), .Z(n19394) );
  NAND U19928 ( .A(n38470), .B(n19190), .Z(n19192) );
  XOR U19929 ( .A(b[31]), .B(a[114]), .Z(n19351) );
  NAND U19930 ( .A(n38453), .B(n19351), .Z(n19191) );
  AND U19931 ( .A(n19192), .B(n19191), .Z(n19363) );
  NAND U19932 ( .A(n181), .B(n19193), .Z(n19195) );
  XOR U19933 ( .A(b[3]), .B(a[142]), .Z(n19354) );
  NAND U19934 ( .A(n182), .B(n19354), .Z(n19194) );
  AND U19935 ( .A(n19195), .B(n19194), .Z(n19361) );
  NAND U19936 ( .A(n189), .B(n19196), .Z(n19198) );
  XOR U19937 ( .A(b[17]), .B(a[128]), .Z(n19357) );
  NAND U19938 ( .A(n37652), .B(n19357), .Z(n19197) );
  NAND U19939 ( .A(n19198), .B(n19197), .Z(n19360) );
  XNOR U19940 ( .A(n19361), .B(n19360), .Z(n19362) );
  XOR U19941 ( .A(n19363), .B(n19362), .Z(n19395) );
  XOR U19942 ( .A(n19394), .B(n19395), .Z(n19397) );
  XOR U19943 ( .A(n19396), .B(n19397), .Z(n19331) );
  NANDN U19944 ( .A(n19200), .B(n19199), .Z(n19204) );
  NANDN U19945 ( .A(n19202), .B(n19201), .Z(n19203) );
  AND U19946 ( .A(n19204), .B(n19203), .Z(n19384) );
  NANDN U19947 ( .A(n19206), .B(n19205), .Z(n19210) );
  NANDN U19948 ( .A(n19208), .B(n19207), .Z(n19209) );
  NAND U19949 ( .A(n19210), .B(n19209), .Z(n19385) );
  XNOR U19950 ( .A(n19384), .B(n19385), .Z(n19386) );
  NANDN U19951 ( .A(n19212), .B(n19211), .Z(n19216) );
  NANDN U19952 ( .A(n19214), .B(n19213), .Z(n19215) );
  NAND U19953 ( .A(n19216), .B(n19215), .Z(n19387) );
  XNOR U19954 ( .A(n19386), .B(n19387), .Z(n19330) );
  XNOR U19955 ( .A(n19331), .B(n19330), .Z(n19333) );
  NANDN U19956 ( .A(n19218), .B(n19217), .Z(n19222) );
  NANDN U19957 ( .A(n19220), .B(n19219), .Z(n19221) );
  AND U19958 ( .A(n19222), .B(n19221), .Z(n19332) );
  XOR U19959 ( .A(n19333), .B(n19332), .Z(n19444) );
  NANDN U19960 ( .A(n19224), .B(n19223), .Z(n19228) );
  NANDN U19961 ( .A(n19226), .B(n19225), .Z(n19227) );
  AND U19962 ( .A(n19228), .B(n19227), .Z(n19442) );
  NANDN U19963 ( .A(n19230), .B(n19229), .Z(n19234) );
  NANDN U19964 ( .A(n19232), .B(n19231), .Z(n19233) );
  AND U19965 ( .A(n19234), .B(n19233), .Z(n19327) );
  NANDN U19966 ( .A(n19236), .B(n19235), .Z(n19240) );
  OR U19967 ( .A(n19238), .B(n19237), .Z(n19239) );
  AND U19968 ( .A(n19240), .B(n19239), .Z(n19325) );
  NANDN U19969 ( .A(n19242), .B(n19241), .Z(n19246) );
  NANDN U19970 ( .A(n19244), .B(n19243), .Z(n19245) );
  AND U19971 ( .A(n19246), .B(n19245), .Z(n19391) );
  NANDN U19972 ( .A(n19248), .B(n19247), .Z(n19252) );
  NANDN U19973 ( .A(n19250), .B(n19249), .Z(n19251) );
  NAND U19974 ( .A(n19252), .B(n19251), .Z(n19390) );
  XNOR U19975 ( .A(n19391), .B(n19390), .Z(n19393) );
  NAND U19976 ( .A(b[0]), .B(a[144]), .Z(n19253) );
  XNOR U19977 ( .A(b[1]), .B(n19253), .Z(n19255) );
  NANDN U19978 ( .A(b[0]), .B(a[143]), .Z(n19254) );
  NAND U19979 ( .A(n19255), .B(n19254), .Z(n19339) );
  NAND U19980 ( .A(n194), .B(n19256), .Z(n19258) );
  XOR U19981 ( .A(b[29]), .B(a[116]), .Z(n19412) );
  NAND U19982 ( .A(n38456), .B(n19412), .Z(n19257) );
  AND U19983 ( .A(n19258), .B(n19257), .Z(n19337) );
  AND U19984 ( .A(b[31]), .B(a[112]), .Z(n19336) );
  XNOR U19985 ( .A(n19337), .B(n19336), .Z(n19338) );
  XNOR U19986 ( .A(n19339), .B(n19338), .Z(n19379) );
  NAND U19987 ( .A(n38185), .B(n19259), .Z(n19261) );
  XOR U19988 ( .A(b[23]), .B(a[122]), .Z(n19418) );
  NAND U19989 ( .A(n38132), .B(n19418), .Z(n19260) );
  AND U19990 ( .A(n19261), .B(n19260), .Z(n19408) );
  NAND U19991 ( .A(n184), .B(n19262), .Z(n19264) );
  XOR U19992 ( .A(b[7]), .B(a[138]), .Z(n19421) );
  NAND U19993 ( .A(n36592), .B(n19421), .Z(n19263) );
  AND U19994 ( .A(n19264), .B(n19263), .Z(n19407) );
  NAND U19995 ( .A(n38289), .B(n19265), .Z(n19267) );
  XOR U19996 ( .A(b[25]), .B(a[120]), .Z(n19424) );
  NAND U19997 ( .A(n38247), .B(n19424), .Z(n19266) );
  NAND U19998 ( .A(n19267), .B(n19266), .Z(n19406) );
  XOR U19999 ( .A(n19407), .B(n19406), .Z(n19409) );
  XOR U20000 ( .A(n19408), .B(n19409), .Z(n19378) );
  XOR U20001 ( .A(n19379), .B(n19378), .Z(n19381) );
  NAND U20002 ( .A(n187), .B(n19268), .Z(n19270) );
  XOR U20003 ( .A(b[13]), .B(a[132]), .Z(n19427) );
  NAND U20004 ( .A(n37295), .B(n19427), .Z(n19269) );
  AND U20005 ( .A(n19270), .B(n19269), .Z(n19373) );
  NAND U20006 ( .A(n186), .B(n19271), .Z(n19273) );
  XOR U20007 ( .A(b[11]), .B(a[134]), .Z(n19430) );
  NAND U20008 ( .A(n37097), .B(n19430), .Z(n19272) );
  NAND U20009 ( .A(n19273), .B(n19272), .Z(n19372) );
  XNOR U20010 ( .A(n19373), .B(n19372), .Z(n19375) );
  NAND U20011 ( .A(n188), .B(n19274), .Z(n19276) );
  XOR U20012 ( .A(b[15]), .B(a[130]), .Z(n19433) );
  NAND U20013 ( .A(n37382), .B(n19433), .Z(n19275) );
  AND U20014 ( .A(n19276), .B(n19275), .Z(n19369) );
  NAND U20015 ( .A(n38064), .B(n19277), .Z(n19279) );
  XOR U20016 ( .A(b[21]), .B(a[124]), .Z(n19436) );
  NAND U20017 ( .A(n37993), .B(n19436), .Z(n19278) );
  AND U20018 ( .A(n19279), .B(n19278), .Z(n19367) );
  NAND U20019 ( .A(n185), .B(n19280), .Z(n19282) );
  XOR U20020 ( .A(b[9]), .B(a[136]), .Z(n19439) );
  NAND U20021 ( .A(n36805), .B(n19439), .Z(n19281) );
  NAND U20022 ( .A(n19282), .B(n19281), .Z(n19366) );
  XNOR U20023 ( .A(n19367), .B(n19366), .Z(n19368) );
  XNOR U20024 ( .A(n19369), .B(n19368), .Z(n19374) );
  XOR U20025 ( .A(n19375), .B(n19374), .Z(n19380) );
  XNOR U20026 ( .A(n19381), .B(n19380), .Z(n19392) );
  XNOR U20027 ( .A(n19393), .B(n19392), .Z(n19324) );
  XNOR U20028 ( .A(n19325), .B(n19324), .Z(n19326) );
  XOR U20029 ( .A(n19327), .B(n19326), .Z(n19443) );
  XOR U20030 ( .A(n19442), .B(n19443), .Z(n19445) );
  XOR U20031 ( .A(n19444), .B(n19445), .Z(n19321) );
  NANDN U20032 ( .A(n19284), .B(n19283), .Z(n19288) );
  NAND U20033 ( .A(n19286), .B(n19285), .Z(n19287) );
  AND U20034 ( .A(n19288), .B(n19287), .Z(n19319) );
  NANDN U20035 ( .A(n19290), .B(n19289), .Z(n19294) );
  NANDN U20036 ( .A(n19292), .B(n19291), .Z(n19293) );
  AND U20037 ( .A(n19294), .B(n19293), .Z(n19318) );
  XNOR U20038 ( .A(n19319), .B(n19318), .Z(n19320) );
  XNOR U20039 ( .A(n19321), .B(n19320), .Z(n19312) );
  NANDN U20040 ( .A(n19296), .B(n19295), .Z(n19300) );
  NANDN U20041 ( .A(n19298), .B(n19297), .Z(n19299) );
  NAND U20042 ( .A(n19300), .B(n19299), .Z(n19313) );
  XOR U20043 ( .A(n19312), .B(n19313), .Z(n19315) );
  XNOR U20044 ( .A(n19314), .B(n19315), .Z(n19306) );
  XNOR U20045 ( .A(n19307), .B(n19306), .Z(n19308) );
  XNOR U20046 ( .A(n19309), .B(n19308), .Z(n19448) );
  XNOR U20047 ( .A(sreg[368]), .B(n19448), .Z(n19450) );
  NANDN U20048 ( .A(sreg[367]), .B(n19301), .Z(n19305) );
  NAND U20049 ( .A(n19303), .B(n19302), .Z(n19304) );
  NAND U20050 ( .A(n19305), .B(n19304), .Z(n19449) );
  XNOR U20051 ( .A(n19450), .B(n19449), .Z(c[368]) );
  NANDN U20052 ( .A(n19307), .B(n19306), .Z(n19311) );
  NANDN U20053 ( .A(n19309), .B(n19308), .Z(n19310) );
  AND U20054 ( .A(n19311), .B(n19310), .Z(n19456) );
  NANDN U20055 ( .A(n19313), .B(n19312), .Z(n19317) );
  NANDN U20056 ( .A(n19315), .B(n19314), .Z(n19316) );
  AND U20057 ( .A(n19317), .B(n19316), .Z(n19454) );
  NANDN U20058 ( .A(n19319), .B(n19318), .Z(n19323) );
  NANDN U20059 ( .A(n19321), .B(n19320), .Z(n19322) );
  AND U20060 ( .A(n19323), .B(n19322), .Z(n19462) );
  NANDN U20061 ( .A(n19325), .B(n19324), .Z(n19329) );
  NANDN U20062 ( .A(n19327), .B(n19326), .Z(n19328) );
  AND U20063 ( .A(n19329), .B(n19328), .Z(n19466) );
  NANDN U20064 ( .A(n19331), .B(n19330), .Z(n19335) );
  NAND U20065 ( .A(n19333), .B(n19332), .Z(n19334) );
  AND U20066 ( .A(n19335), .B(n19334), .Z(n19465) );
  XNOR U20067 ( .A(n19466), .B(n19465), .Z(n19468) );
  NANDN U20068 ( .A(n19337), .B(n19336), .Z(n19341) );
  NANDN U20069 ( .A(n19339), .B(n19338), .Z(n19340) );
  AND U20070 ( .A(n19341), .B(n19340), .Z(n19533) );
  NAND U20071 ( .A(n38385), .B(n19342), .Z(n19344) );
  XOR U20072 ( .A(b[27]), .B(a[119]), .Z(n19477) );
  NAND U20073 ( .A(n38343), .B(n19477), .Z(n19343) );
  AND U20074 ( .A(n19344), .B(n19343), .Z(n19540) );
  NAND U20075 ( .A(n183), .B(n19345), .Z(n19347) );
  XOR U20076 ( .A(b[5]), .B(a[141]), .Z(n19480) );
  NAND U20077 ( .A(n36296), .B(n19480), .Z(n19346) );
  AND U20078 ( .A(n19347), .B(n19346), .Z(n19538) );
  NAND U20079 ( .A(n190), .B(n19348), .Z(n19350) );
  XOR U20080 ( .A(b[19]), .B(a[127]), .Z(n19483) );
  NAND U20081 ( .A(n37821), .B(n19483), .Z(n19349) );
  NAND U20082 ( .A(n19350), .B(n19349), .Z(n19537) );
  XNOR U20083 ( .A(n19538), .B(n19537), .Z(n19539) );
  XNOR U20084 ( .A(n19540), .B(n19539), .Z(n19531) );
  NAND U20085 ( .A(n38470), .B(n19351), .Z(n19353) );
  XOR U20086 ( .A(b[31]), .B(a[115]), .Z(n19486) );
  NAND U20087 ( .A(n38453), .B(n19486), .Z(n19352) );
  AND U20088 ( .A(n19353), .B(n19352), .Z(n19498) );
  NAND U20089 ( .A(n181), .B(n19354), .Z(n19356) );
  XOR U20090 ( .A(b[3]), .B(a[143]), .Z(n19489) );
  NAND U20091 ( .A(n182), .B(n19489), .Z(n19355) );
  AND U20092 ( .A(n19356), .B(n19355), .Z(n19496) );
  NAND U20093 ( .A(n189), .B(n19357), .Z(n19359) );
  XOR U20094 ( .A(b[17]), .B(a[129]), .Z(n19492) );
  NAND U20095 ( .A(n37652), .B(n19492), .Z(n19358) );
  NAND U20096 ( .A(n19359), .B(n19358), .Z(n19495) );
  XNOR U20097 ( .A(n19496), .B(n19495), .Z(n19497) );
  XOR U20098 ( .A(n19498), .B(n19497), .Z(n19532) );
  XOR U20099 ( .A(n19531), .B(n19532), .Z(n19534) );
  XOR U20100 ( .A(n19533), .B(n19534), .Z(n19580) );
  NANDN U20101 ( .A(n19361), .B(n19360), .Z(n19365) );
  NANDN U20102 ( .A(n19363), .B(n19362), .Z(n19364) );
  AND U20103 ( .A(n19365), .B(n19364), .Z(n19519) );
  NANDN U20104 ( .A(n19367), .B(n19366), .Z(n19371) );
  NANDN U20105 ( .A(n19369), .B(n19368), .Z(n19370) );
  NAND U20106 ( .A(n19371), .B(n19370), .Z(n19520) );
  XNOR U20107 ( .A(n19519), .B(n19520), .Z(n19521) );
  NANDN U20108 ( .A(n19373), .B(n19372), .Z(n19377) );
  NAND U20109 ( .A(n19375), .B(n19374), .Z(n19376) );
  NAND U20110 ( .A(n19377), .B(n19376), .Z(n19522) );
  XNOR U20111 ( .A(n19521), .B(n19522), .Z(n19579) );
  XNOR U20112 ( .A(n19580), .B(n19579), .Z(n19582) );
  NAND U20113 ( .A(n19379), .B(n19378), .Z(n19383) );
  NAND U20114 ( .A(n19381), .B(n19380), .Z(n19382) );
  AND U20115 ( .A(n19383), .B(n19382), .Z(n19581) );
  XOR U20116 ( .A(n19582), .B(n19581), .Z(n19594) );
  NANDN U20117 ( .A(n19385), .B(n19384), .Z(n19389) );
  NANDN U20118 ( .A(n19387), .B(n19386), .Z(n19388) );
  AND U20119 ( .A(n19389), .B(n19388), .Z(n19591) );
  NANDN U20120 ( .A(n19395), .B(n19394), .Z(n19399) );
  OR U20121 ( .A(n19397), .B(n19396), .Z(n19398) );
  AND U20122 ( .A(n19399), .B(n19398), .Z(n19586) );
  NANDN U20123 ( .A(n19401), .B(n19400), .Z(n19405) );
  NANDN U20124 ( .A(n19403), .B(n19402), .Z(n19404) );
  AND U20125 ( .A(n19405), .B(n19404), .Z(n19526) );
  NANDN U20126 ( .A(n19407), .B(n19406), .Z(n19411) );
  OR U20127 ( .A(n19409), .B(n19408), .Z(n19410) );
  NAND U20128 ( .A(n19411), .B(n19410), .Z(n19525) );
  XNOR U20129 ( .A(n19526), .B(n19525), .Z(n19527) );
  NAND U20130 ( .A(n194), .B(n19412), .Z(n19414) );
  XOR U20131 ( .A(b[29]), .B(a[117]), .Z(n19552) );
  NAND U20132 ( .A(n38456), .B(n19552), .Z(n19413) );
  AND U20133 ( .A(n19414), .B(n19413), .Z(n19472) );
  AND U20134 ( .A(b[31]), .B(a[113]), .Z(n19471) );
  XNOR U20135 ( .A(n19472), .B(n19471), .Z(n19473) );
  NAND U20136 ( .A(b[0]), .B(a[145]), .Z(n19415) );
  XNOR U20137 ( .A(b[1]), .B(n19415), .Z(n19417) );
  NANDN U20138 ( .A(b[0]), .B(a[144]), .Z(n19416) );
  NAND U20139 ( .A(n19417), .B(n19416), .Z(n19474) );
  XNOR U20140 ( .A(n19473), .B(n19474), .Z(n19513) );
  NAND U20141 ( .A(n38185), .B(n19418), .Z(n19420) );
  XOR U20142 ( .A(b[23]), .B(a[123]), .Z(n19555) );
  NAND U20143 ( .A(n38132), .B(n19555), .Z(n19419) );
  AND U20144 ( .A(n19420), .B(n19419), .Z(n19546) );
  NAND U20145 ( .A(n184), .B(n19421), .Z(n19423) );
  XOR U20146 ( .A(b[7]), .B(a[139]), .Z(n19558) );
  NAND U20147 ( .A(n36592), .B(n19558), .Z(n19422) );
  AND U20148 ( .A(n19423), .B(n19422), .Z(n19544) );
  NAND U20149 ( .A(n38289), .B(n19424), .Z(n19426) );
  XOR U20150 ( .A(b[25]), .B(a[121]), .Z(n19561) );
  NAND U20151 ( .A(n38247), .B(n19561), .Z(n19425) );
  NAND U20152 ( .A(n19426), .B(n19425), .Z(n19543) );
  XNOR U20153 ( .A(n19544), .B(n19543), .Z(n19545) );
  XOR U20154 ( .A(n19546), .B(n19545), .Z(n19514) );
  XNOR U20155 ( .A(n19513), .B(n19514), .Z(n19515) );
  NAND U20156 ( .A(n187), .B(n19427), .Z(n19429) );
  XOR U20157 ( .A(b[13]), .B(a[133]), .Z(n19564) );
  NAND U20158 ( .A(n37295), .B(n19564), .Z(n19428) );
  AND U20159 ( .A(n19429), .B(n19428), .Z(n19508) );
  NAND U20160 ( .A(n186), .B(n19430), .Z(n19432) );
  XOR U20161 ( .A(b[11]), .B(a[135]), .Z(n19567) );
  NAND U20162 ( .A(n37097), .B(n19567), .Z(n19431) );
  NAND U20163 ( .A(n19432), .B(n19431), .Z(n19507) );
  XNOR U20164 ( .A(n19508), .B(n19507), .Z(n19509) );
  NAND U20165 ( .A(n188), .B(n19433), .Z(n19435) );
  XOR U20166 ( .A(b[15]), .B(a[131]), .Z(n19570) );
  NAND U20167 ( .A(n37382), .B(n19570), .Z(n19434) );
  AND U20168 ( .A(n19435), .B(n19434), .Z(n19504) );
  NAND U20169 ( .A(n38064), .B(n19436), .Z(n19438) );
  XOR U20170 ( .A(b[21]), .B(a[125]), .Z(n19573) );
  NAND U20171 ( .A(n37993), .B(n19573), .Z(n19437) );
  AND U20172 ( .A(n19438), .B(n19437), .Z(n19502) );
  NAND U20173 ( .A(n185), .B(n19439), .Z(n19441) );
  XOR U20174 ( .A(b[9]), .B(a[137]), .Z(n19576) );
  NAND U20175 ( .A(n36805), .B(n19576), .Z(n19440) );
  NAND U20176 ( .A(n19441), .B(n19440), .Z(n19501) );
  XNOR U20177 ( .A(n19502), .B(n19501), .Z(n19503) );
  XOR U20178 ( .A(n19504), .B(n19503), .Z(n19510) );
  XOR U20179 ( .A(n19509), .B(n19510), .Z(n19516) );
  XOR U20180 ( .A(n19515), .B(n19516), .Z(n19528) );
  XNOR U20181 ( .A(n19527), .B(n19528), .Z(n19585) );
  XNOR U20182 ( .A(n19586), .B(n19585), .Z(n19587) );
  XOR U20183 ( .A(n19588), .B(n19587), .Z(n19592) );
  XNOR U20184 ( .A(n19591), .B(n19592), .Z(n19593) );
  XNOR U20185 ( .A(n19594), .B(n19593), .Z(n19467) );
  XOR U20186 ( .A(n19468), .B(n19467), .Z(n19460) );
  NANDN U20187 ( .A(n19443), .B(n19442), .Z(n19447) );
  OR U20188 ( .A(n19445), .B(n19444), .Z(n19446) );
  AND U20189 ( .A(n19447), .B(n19446), .Z(n19459) );
  XNOR U20190 ( .A(n19460), .B(n19459), .Z(n19461) );
  XNOR U20191 ( .A(n19462), .B(n19461), .Z(n19453) );
  XNOR U20192 ( .A(n19454), .B(n19453), .Z(n19455) );
  XNOR U20193 ( .A(n19456), .B(n19455), .Z(n19597) );
  XNOR U20194 ( .A(sreg[369]), .B(n19597), .Z(n19599) );
  NANDN U20195 ( .A(sreg[368]), .B(n19448), .Z(n19452) );
  NAND U20196 ( .A(n19450), .B(n19449), .Z(n19451) );
  NAND U20197 ( .A(n19452), .B(n19451), .Z(n19598) );
  XNOR U20198 ( .A(n19599), .B(n19598), .Z(c[369]) );
  NANDN U20199 ( .A(n19454), .B(n19453), .Z(n19458) );
  NANDN U20200 ( .A(n19456), .B(n19455), .Z(n19457) );
  AND U20201 ( .A(n19458), .B(n19457), .Z(n19605) );
  NANDN U20202 ( .A(n19460), .B(n19459), .Z(n19464) );
  NANDN U20203 ( .A(n19462), .B(n19461), .Z(n19463) );
  AND U20204 ( .A(n19464), .B(n19463), .Z(n19603) );
  NANDN U20205 ( .A(n19466), .B(n19465), .Z(n19470) );
  NAND U20206 ( .A(n19468), .B(n19467), .Z(n19469) );
  AND U20207 ( .A(n19470), .B(n19469), .Z(n19610) );
  NANDN U20208 ( .A(n19472), .B(n19471), .Z(n19476) );
  NANDN U20209 ( .A(n19474), .B(n19473), .Z(n19475) );
  AND U20210 ( .A(n19476), .B(n19475), .Z(n19694) );
  NAND U20211 ( .A(n38385), .B(n19477), .Z(n19479) );
  XOR U20212 ( .A(b[27]), .B(a[120]), .Z(n19638) );
  NAND U20213 ( .A(n38343), .B(n19638), .Z(n19478) );
  AND U20214 ( .A(n19479), .B(n19478), .Z(n19701) );
  NAND U20215 ( .A(n183), .B(n19480), .Z(n19482) );
  XOR U20216 ( .A(b[5]), .B(a[142]), .Z(n19641) );
  NAND U20217 ( .A(n36296), .B(n19641), .Z(n19481) );
  AND U20218 ( .A(n19482), .B(n19481), .Z(n19699) );
  NAND U20219 ( .A(n190), .B(n19483), .Z(n19485) );
  XOR U20220 ( .A(b[19]), .B(a[128]), .Z(n19644) );
  NAND U20221 ( .A(n37821), .B(n19644), .Z(n19484) );
  NAND U20222 ( .A(n19485), .B(n19484), .Z(n19698) );
  XNOR U20223 ( .A(n19699), .B(n19698), .Z(n19700) );
  XNOR U20224 ( .A(n19701), .B(n19700), .Z(n19692) );
  NAND U20225 ( .A(n38470), .B(n19486), .Z(n19488) );
  XOR U20226 ( .A(b[31]), .B(a[116]), .Z(n19647) );
  NAND U20227 ( .A(n38453), .B(n19647), .Z(n19487) );
  AND U20228 ( .A(n19488), .B(n19487), .Z(n19659) );
  NAND U20229 ( .A(n181), .B(n19489), .Z(n19491) );
  XOR U20230 ( .A(b[3]), .B(a[144]), .Z(n19650) );
  NAND U20231 ( .A(n182), .B(n19650), .Z(n19490) );
  AND U20232 ( .A(n19491), .B(n19490), .Z(n19657) );
  NAND U20233 ( .A(n189), .B(n19492), .Z(n19494) );
  XOR U20234 ( .A(b[17]), .B(a[130]), .Z(n19653) );
  NAND U20235 ( .A(n37652), .B(n19653), .Z(n19493) );
  NAND U20236 ( .A(n19494), .B(n19493), .Z(n19656) );
  XNOR U20237 ( .A(n19657), .B(n19656), .Z(n19658) );
  XOR U20238 ( .A(n19659), .B(n19658), .Z(n19693) );
  XOR U20239 ( .A(n19692), .B(n19693), .Z(n19695) );
  XOR U20240 ( .A(n19694), .B(n19695), .Z(n19627) );
  NANDN U20241 ( .A(n19496), .B(n19495), .Z(n19500) );
  NANDN U20242 ( .A(n19498), .B(n19497), .Z(n19499) );
  AND U20243 ( .A(n19500), .B(n19499), .Z(n19680) );
  NANDN U20244 ( .A(n19502), .B(n19501), .Z(n19506) );
  NANDN U20245 ( .A(n19504), .B(n19503), .Z(n19505) );
  NAND U20246 ( .A(n19506), .B(n19505), .Z(n19681) );
  XNOR U20247 ( .A(n19680), .B(n19681), .Z(n19682) );
  NANDN U20248 ( .A(n19508), .B(n19507), .Z(n19512) );
  NANDN U20249 ( .A(n19510), .B(n19509), .Z(n19511) );
  NAND U20250 ( .A(n19512), .B(n19511), .Z(n19683) );
  XNOR U20251 ( .A(n19682), .B(n19683), .Z(n19626) );
  XNOR U20252 ( .A(n19627), .B(n19626), .Z(n19629) );
  NANDN U20253 ( .A(n19514), .B(n19513), .Z(n19518) );
  NANDN U20254 ( .A(n19516), .B(n19515), .Z(n19517) );
  AND U20255 ( .A(n19518), .B(n19517), .Z(n19628) );
  XOR U20256 ( .A(n19629), .B(n19628), .Z(n19742) );
  NANDN U20257 ( .A(n19520), .B(n19519), .Z(n19524) );
  NANDN U20258 ( .A(n19522), .B(n19521), .Z(n19523) );
  AND U20259 ( .A(n19524), .B(n19523), .Z(n19740) );
  NANDN U20260 ( .A(n19526), .B(n19525), .Z(n19530) );
  NANDN U20261 ( .A(n19528), .B(n19527), .Z(n19529) );
  AND U20262 ( .A(n19530), .B(n19529), .Z(n19623) );
  NANDN U20263 ( .A(n19532), .B(n19531), .Z(n19536) );
  OR U20264 ( .A(n19534), .B(n19533), .Z(n19535) );
  AND U20265 ( .A(n19536), .B(n19535), .Z(n19621) );
  NANDN U20266 ( .A(n19538), .B(n19537), .Z(n19542) );
  NANDN U20267 ( .A(n19540), .B(n19539), .Z(n19541) );
  AND U20268 ( .A(n19542), .B(n19541), .Z(n19687) );
  NANDN U20269 ( .A(n19544), .B(n19543), .Z(n19548) );
  NANDN U20270 ( .A(n19546), .B(n19545), .Z(n19547) );
  NAND U20271 ( .A(n19548), .B(n19547), .Z(n19686) );
  XNOR U20272 ( .A(n19687), .B(n19686), .Z(n19688) );
  NAND U20273 ( .A(b[0]), .B(a[146]), .Z(n19549) );
  XNOR U20274 ( .A(b[1]), .B(n19549), .Z(n19551) );
  NANDN U20275 ( .A(b[0]), .B(a[145]), .Z(n19550) );
  NAND U20276 ( .A(n19551), .B(n19550), .Z(n19635) );
  NAND U20277 ( .A(n194), .B(n19552), .Z(n19554) );
  XOR U20278 ( .A(b[29]), .B(a[118]), .Z(n19713) );
  NAND U20279 ( .A(n38456), .B(n19713), .Z(n19553) );
  AND U20280 ( .A(n19554), .B(n19553), .Z(n19633) );
  AND U20281 ( .A(b[31]), .B(a[114]), .Z(n19632) );
  XNOR U20282 ( .A(n19633), .B(n19632), .Z(n19634) );
  XNOR U20283 ( .A(n19635), .B(n19634), .Z(n19674) );
  NAND U20284 ( .A(n38185), .B(n19555), .Z(n19557) );
  XOR U20285 ( .A(b[23]), .B(a[124]), .Z(n19716) );
  NAND U20286 ( .A(n38132), .B(n19716), .Z(n19556) );
  AND U20287 ( .A(n19557), .B(n19556), .Z(n19707) );
  NAND U20288 ( .A(n184), .B(n19558), .Z(n19560) );
  XOR U20289 ( .A(b[7]), .B(a[140]), .Z(n19719) );
  NAND U20290 ( .A(n36592), .B(n19719), .Z(n19559) );
  AND U20291 ( .A(n19560), .B(n19559), .Z(n19705) );
  NAND U20292 ( .A(n38289), .B(n19561), .Z(n19563) );
  XOR U20293 ( .A(b[25]), .B(a[122]), .Z(n19722) );
  NAND U20294 ( .A(n38247), .B(n19722), .Z(n19562) );
  NAND U20295 ( .A(n19563), .B(n19562), .Z(n19704) );
  XNOR U20296 ( .A(n19705), .B(n19704), .Z(n19706) );
  XOR U20297 ( .A(n19707), .B(n19706), .Z(n19675) );
  XNOR U20298 ( .A(n19674), .B(n19675), .Z(n19676) );
  NAND U20299 ( .A(n187), .B(n19564), .Z(n19566) );
  XOR U20300 ( .A(b[13]), .B(a[134]), .Z(n19725) );
  NAND U20301 ( .A(n37295), .B(n19725), .Z(n19565) );
  AND U20302 ( .A(n19566), .B(n19565), .Z(n19669) );
  NAND U20303 ( .A(n186), .B(n19567), .Z(n19569) );
  XOR U20304 ( .A(b[11]), .B(a[136]), .Z(n19728) );
  NAND U20305 ( .A(n37097), .B(n19728), .Z(n19568) );
  NAND U20306 ( .A(n19569), .B(n19568), .Z(n19668) );
  XNOR U20307 ( .A(n19669), .B(n19668), .Z(n19670) );
  NAND U20308 ( .A(n188), .B(n19570), .Z(n19572) );
  XOR U20309 ( .A(b[15]), .B(a[132]), .Z(n19731) );
  NAND U20310 ( .A(n37382), .B(n19731), .Z(n19571) );
  AND U20311 ( .A(n19572), .B(n19571), .Z(n19665) );
  NAND U20312 ( .A(n38064), .B(n19573), .Z(n19575) );
  XOR U20313 ( .A(b[21]), .B(a[126]), .Z(n19734) );
  NAND U20314 ( .A(n37993), .B(n19734), .Z(n19574) );
  AND U20315 ( .A(n19575), .B(n19574), .Z(n19663) );
  NAND U20316 ( .A(n185), .B(n19576), .Z(n19578) );
  XOR U20317 ( .A(b[9]), .B(a[138]), .Z(n19737) );
  NAND U20318 ( .A(n36805), .B(n19737), .Z(n19577) );
  NAND U20319 ( .A(n19578), .B(n19577), .Z(n19662) );
  XNOR U20320 ( .A(n19663), .B(n19662), .Z(n19664) );
  XOR U20321 ( .A(n19665), .B(n19664), .Z(n19671) );
  XOR U20322 ( .A(n19670), .B(n19671), .Z(n19677) );
  XOR U20323 ( .A(n19676), .B(n19677), .Z(n19689) );
  XNOR U20324 ( .A(n19688), .B(n19689), .Z(n19620) );
  XNOR U20325 ( .A(n19621), .B(n19620), .Z(n19622) );
  XOR U20326 ( .A(n19623), .B(n19622), .Z(n19741) );
  XOR U20327 ( .A(n19740), .B(n19741), .Z(n19743) );
  XOR U20328 ( .A(n19742), .B(n19743), .Z(n19617) );
  NANDN U20329 ( .A(n19580), .B(n19579), .Z(n19584) );
  NAND U20330 ( .A(n19582), .B(n19581), .Z(n19583) );
  AND U20331 ( .A(n19584), .B(n19583), .Z(n19615) );
  NANDN U20332 ( .A(n19586), .B(n19585), .Z(n19590) );
  NANDN U20333 ( .A(n19588), .B(n19587), .Z(n19589) );
  AND U20334 ( .A(n19590), .B(n19589), .Z(n19614) );
  XNOR U20335 ( .A(n19615), .B(n19614), .Z(n19616) );
  XNOR U20336 ( .A(n19617), .B(n19616), .Z(n19608) );
  NANDN U20337 ( .A(n19592), .B(n19591), .Z(n19596) );
  NANDN U20338 ( .A(n19594), .B(n19593), .Z(n19595) );
  NAND U20339 ( .A(n19596), .B(n19595), .Z(n19609) );
  XOR U20340 ( .A(n19608), .B(n19609), .Z(n19611) );
  XNOR U20341 ( .A(n19610), .B(n19611), .Z(n19602) );
  XNOR U20342 ( .A(n19603), .B(n19602), .Z(n19604) );
  XNOR U20343 ( .A(n19605), .B(n19604), .Z(n19746) );
  XNOR U20344 ( .A(sreg[370]), .B(n19746), .Z(n19748) );
  NANDN U20345 ( .A(sreg[369]), .B(n19597), .Z(n19601) );
  NAND U20346 ( .A(n19599), .B(n19598), .Z(n19600) );
  NAND U20347 ( .A(n19601), .B(n19600), .Z(n19747) );
  XNOR U20348 ( .A(n19748), .B(n19747), .Z(c[370]) );
  NANDN U20349 ( .A(n19603), .B(n19602), .Z(n19607) );
  NANDN U20350 ( .A(n19605), .B(n19604), .Z(n19606) );
  AND U20351 ( .A(n19607), .B(n19606), .Z(n19754) );
  NANDN U20352 ( .A(n19609), .B(n19608), .Z(n19613) );
  NANDN U20353 ( .A(n19611), .B(n19610), .Z(n19612) );
  AND U20354 ( .A(n19613), .B(n19612), .Z(n19752) );
  NANDN U20355 ( .A(n19615), .B(n19614), .Z(n19619) );
  NANDN U20356 ( .A(n19617), .B(n19616), .Z(n19618) );
  AND U20357 ( .A(n19619), .B(n19618), .Z(n19760) );
  NANDN U20358 ( .A(n19621), .B(n19620), .Z(n19625) );
  NANDN U20359 ( .A(n19623), .B(n19622), .Z(n19624) );
  AND U20360 ( .A(n19625), .B(n19624), .Z(n19764) );
  NANDN U20361 ( .A(n19627), .B(n19626), .Z(n19631) );
  NAND U20362 ( .A(n19629), .B(n19628), .Z(n19630) );
  AND U20363 ( .A(n19631), .B(n19630), .Z(n19763) );
  XNOR U20364 ( .A(n19764), .B(n19763), .Z(n19766) );
  NANDN U20365 ( .A(n19633), .B(n19632), .Z(n19637) );
  NANDN U20366 ( .A(n19635), .B(n19634), .Z(n19636) );
  AND U20367 ( .A(n19637), .B(n19636), .Z(n19843) );
  NAND U20368 ( .A(n38385), .B(n19638), .Z(n19640) );
  XOR U20369 ( .A(b[27]), .B(a[121]), .Z(n19787) );
  NAND U20370 ( .A(n38343), .B(n19787), .Z(n19639) );
  AND U20371 ( .A(n19640), .B(n19639), .Z(n19850) );
  NAND U20372 ( .A(n183), .B(n19641), .Z(n19643) );
  XOR U20373 ( .A(b[5]), .B(a[143]), .Z(n19790) );
  NAND U20374 ( .A(n36296), .B(n19790), .Z(n19642) );
  AND U20375 ( .A(n19643), .B(n19642), .Z(n19848) );
  NAND U20376 ( .A(n190), .B(n19644), .Z(n19646) );
  XOR U20377 ( .A(b[19]), .B(a[129]), .Z(n19793) );
  NAND U20378 ( .A(n37821), .B(n19793), .Z(n19645) );
  NAND U20379 ( .A(n19646), .B(n19645), .Z(n19847) );
  XNOR U20380 ( .A(n19848), .B(n19847), .Z(n19849) );
  XNOR U20381 ( .A(n19850), .B(n19849), .Z(n19841) );
  NAND U20382 ( .A(n38470), .B(n19647), .Z(n19649) );
  XOR U20383 ( .A(b[31]), .B(a[117]), .Z(n19796) );
  NAND U20384 ( .A(n38453), .B(n19796), .Z(n19648) );
  AND U20385 ( .A(n19649), .B(n19648), .Z(n19808) );
  NAND U20386 ( .A(n181), .B(n19650), .Z(n19652) );
  XOR U20387 ( .A(b[3]), .B(a[145]), .Z(n19799) );
  NAND U20388 ( .A(n182), .B(n19799), .Z(n19651) );
  AND U20389 ( .A(n19652), .B(n19651), .Z(n19806) );
  NAND U20390 ( .A(n189), .B(n19653), .Z(n19655) );
  XOR U20391 ( .A(b[17]), .B(a[131]), .Z(n19802) );
  NAND U20392 ( .A(n37652), .B(n19802), .Z(n19654) );
  NAND U20393 ( .A(n19655), .B(n19654), .Z(n19805) );
  XNOR U20394 ( .A(n19806), .B(n19805), .Z(n19807) );
  XOR U20395 ( .A(n19808), .B(n19807), .Z(n19842) );
  XOR U20396 ( .A(n19841), .B(n19842), .Z(n19844) );
  XOR U20397 ( .A(n19843), .B(n19844), .Z(n19776) );
  NANDN U20398 ( .A(n19657), .B(n19656), .Z(n19661) );
  NANDN U20399 ( .A(n19659), .B(n19658), .Z(n19660) );
  AND U20400 ( .A(n19661), .B(n19660), .Z(n19829) );
  NANDN U20401 ( .A(n19663), .B(n19662), .Z(n19667) );
  NANDN U20402 ( .A(n19665), .B(n19664), .Z(n19666) );
  NAND U20403 ( .A(n19667), .B(n19666), .Z(n19830) );
  XNOR U20404 ( .A(n19829), .B(n19830), .Z(n19831) );
  NANDN U20405 ( .A(n19669), .B(n19668), .Z(n19673) );
  NANDN U20406 ( .A(n19671), .B(n19670), .Z(n19672) );
  NAND U20407 ( .A(n19673), .B(n19672), .Z(n19832) );
  XNOR U20408 ( .A(n19831), .B(n19832), .Z(n19775) );
  XNOR U20409 ( .A(n19776), .B(n19775), .Z(n19778) );
  NANDN U20410 ( .A(n19675), .B(n19674), .Z(n19679) );
  NANDN U20411 ( .A(n19677), .B(n19676), .Z(n19678) );
  AND U20412 ( .A(n19679), .B(n19678), .Z(n19777) );
  XOR U20413 ( .A(n19778), .B(n19777), .Z(n19892) );
  NANDN U20414 ( .A(n19681), .B(n19680), .Z(n19685) );
  NANDN U20415 ( .A(n19683), .B(n19682), .Z(n19684) );
  AND U20416 ( .A(n19685), .B(n19684), .Z(n19889) );
  NANDN U20417 ( .A(n19687), .B(n19686), .Z(n19691) );
  NANDN U20418 ( .A(n19689), .B(n19688), .Z(n19690) );
  AND U20419 ( .A(n19691), .B(n19690), .Z(n19772) );
  NANDN U20420 ( .A(n19693), .B(n19692), .Z(n19697) );
  OR U20421 ( .A(n19695), .B(n19694), .Z(n19696) );
  AND U20422 ( .A(n19697), .B(n19696), .Z(n19770) );
  NANDN U20423 ( .A(n19699), .B(n19698), .Z(n19703) );
  NANDN U20424 ( .A(n19701), .B(n19700), .Z(n19702) );
  AND U20425 ( .A(n19703), .B(n19702), .Z(n19836) );
  NANDN U20426 ( .A(n19705), .B(n19704), .Z(n19709) );
  NANDN U20427 ( .A(n19707), .B(n19706), .Z(n19708) );
  NAND U20428 ( .A(n19709), .B(n19708), .Z(n19835) );
  XNOR U20429 ( .A(n19836), .B(n19835), .Z(n19837) );
  NAND U20430 ( .A(b[0]), .B(a[147]), .Z(n19710) );
  XNOR U20431 ( .A(b[1]), .B(n19710), .Z(n19712) );
  NANDN U20432 ( .A(b[0]), .B(a[146]), .Z(n19711) );
  NAND U20433 ( .A(n19712), .B(n19711), .Z(n19784) );
  NAND U20434 ( .A(n194), .B(n19713), .Z(n19715) );
  XOR U20435 ( .A(b[29]), .B(a[119]), .Z(n19862) );
  NAND U20436 ( .A(n38456), .B(n19862), .Z(n19714) );
  AND U20437 ( .A(n19715), .B(n19714), .Z(n19782) );
  AND U20438 ( .A(b[31]), .B(a[115]), .Z(n19781) );
  XNOR U20439 ( .A(n19782), .B(n19781), .Z(n19783) );
  XNOR U20440 ( .A(n19784), .B(n19783), .Z(n19823) );
  NAND U20441 ( .A(n38185), .B(n19716), .Z(n19718) );
  XOR U20442 ( .A(b[23]), .B(a[125]), .Z(n19865) );
  NAND U20443 ( .A(n38132), .B(n19865), .Z(n19717) );
  AND U20444 ( .A(n19718), .B(n19717), .Z(n19856) );
  NAND U20445 ( .A(n184), .B(n19719), .Z(n19721) );
  XOR U20446 ( .A(b[7]), .B(a[141]), .Z(n19868) );
  NAND U20447 ( .A(n36592), .B(n19868), .Z(n19720) );
  AND U20448 ( .A(n19721), .B(n19720), .Z(n19854) );
  NAND U20449 ( .A(n38289), .B(n19722), .Z(n19724) );
  XOR U20450 ( .A(b[25]), .B(a[123]), .Z(n19871) );
  NAND U20451 ( .A(n38247), .B(n19871), .Z(n19723) );
  NAND U20452 ( .A(n19724), .B(n19723), .Z(n19853) );
  XNOR U20453 ( .A(n19854), .B(n19853), .Z(n19855) );
  XOR U20454 ( .A(n19856), .B(n19855), .Z(n19824) );
  XNOR U20455 ( .A(n19823), .B(n19824), .Z(n19825) );
  NAND U20456 ( .A(n187), .B(n19725), .Z(n19727) );
  XOR U20457 ( .A(b[13]), .B(a[135]), .Z(n19874) );
  NAND U20458 ( .A(n37295), .B(n19874), .Z(n19726) );
  AND U20459 ( .A(n19727), .B(n19726), .Z(n19818) );
  NAND U20460 ( .A(n186), .B(n19728), .Z(n19730) );
  XOR U20461 ( .A(b[11]), .B(a[137]), .Z(n19877) );
  NAND U20462 ( .A(n37097), .B(n19877), .Z(n19729) );
  NAND U20463 ( .A(n19730), .B(n19729), .Z(n19817) );
  XNOR U20464 ( .A(n19818), .B(n19817), .Z(n19819) );
  NAND U20465 ( .A(n188), .B(n19731), .Z(n19733) );
  XOR U20466 ( .A(b[15]), .B(a[133]), .Z(n19880) );
  NAND U20467 ( .A(n37382), .B(n19880), .Z(n19732) );
  AND U20468 ( .A(n19733), .B(n19732), .Z(n19814) );
  NAND U20469 ( .A(n38064), .B(n19734), .Z(n19736) );
  XOR U20470 ( .A(b[21]), .B(a[127]), .Z(n19883) );
  NAND U20471 ( .A(n37993), .B(n19883), .Z(n19735) );
  AND U20472 ( .A(n19736), .B(n19735), .Z(n19812) );
  NAND U20473 ( .A(n185), .B(n19737), .Z(n19739) );
  XOR U20474 ( .A(b[9]), .B(a[139]), .Z(n19886) );
  NAND U20475 ( .A(n36805), .B(n19886), .Z(n19738) );
  NAND U20476 ( .A(n19739), .B(n19738), .Z(n19811) );
  XNOR U20477 ( .A(n19812), .B(n19811), .Z(n19813) );
  XOR U20478 ( .A(n19814), .B(n19813), .Z(n19820) );
  XOR U20479 ( .A(n19819), .B(n19820), .Z(n19826) );
  XOR U20480 ( .A(n19825), .B(n19826), .Z(n19838) );
  XNOR U20481 ( .A(n19837), .B(n19838), .Z(n19769) );
  XNOR U20482 ( .A(n19770), .B(n19769), .Z(n19771) );
  XOR U20483 ( .A(n19772), .B(n19771), .Z(n19890) );
  XNOR U20484 ( .A(n19889), .B(n19890), .Z(n19891) );
  XNOR U20485 ( .A(n19892), .B(n19891), .Z(n19765) );
  XOR U20486 ( .A(n19766), .B(n19765), .Z(n19758) );
  NANDN U20487 ( .A(n19741), .B(n19740), .Z(n19745) );
  OR U20488 ( .A(n19743), .B(n19742), .Z(n19744) );
  AND U20489 ( .A(n19745), .B(n19744), .Z(n19757) );
  XNOR U20490 ( .A(n19758), .B(n19757), .Z(n19759) );
  XNOR U20491 ( .A(n19760), .B(n19759), .Z(n19751) );
  XNOR U20492 ( .A(n19752), .B(n19751), .Z(n19753) );
  XNOR U20493 ( .A(n19754), .B(n19753), .Z(n19895) );
  XNOR U20494 ( .A(sreg[371]), .B(n19895), .Z(n19897) );
  NANDN U20495 ( .A(sreg[370]), .B(n19746), .Z(n19750) );
  NAND U20496 ( .A(n19748), .B(n19747), .Z(n19749) );
  NAND U20497 ( .A(n19750), .B(n19749), .Z(n19896) );
  XNOR U20498 ( .A(n19897), .B(n19896), .Z(c[371]) );
  NANDN U20499 ( .A(n19752), .B(n19751), .Z(n19756) );
  NANDN U20500 ( .A(n19754), .B(n19753), .Z(n19755) );
  AND U20501 ( .A(n19756), .B(n19755), .Z(n19903) );
  NANDN U20502 ( .A(n19758), .B(n19757), .Z(n19762) );
  NANDN U20503 ( .A(n19760), .B(n19759), .Z(n19761) );
  AND U20504 ( .A(n19762), .B(n19761), .Z(n19901) );
  NANDN U20505 ( .A(n19764), .B(n19763), .Z(n19768) );
  NAND U20506 ( .A(n19766), .B(n19765), .Z(n19767) );
  AND U20507 ( .A(n19768), .B(n19767), .Z(n19908) );
  NANDN U20508 ( .A(n19770), .B(n19769), .Z(n19774) );
  NANDN U20509 ( .A(n19772), .B(n19771), .Z(n19773) );
  AND U20510 ( .A(n19774), .B(n19773), .Z(n19913) );
  NANDN U20511 ( .A(n19776), .B(n19775), .Z(n19780) );
  NAND U20512 ( .A(n19778), .B(n19777), .Z(n19779) );
  AND U20513 ( .A(n19780), .B(n19779), .Z(n19912) );
  XNOR U20514 ( .A(n19913), .B(n19912), .Z(n19915) );
  NANDN U20515 ( .A(n19782), .B(n19781), .Z(n19786) );
  NANDN U20516 ( .A(n19784), .B(n19783), .Z(n19785) );
  AND U20517 ( .A(n19786), .B(n19785), .Z(n19990) );
  NAND U20518 ( .A(n38385), .B(n19787), .Z(n19789) );
  XOR U20519 ( .A(b[27]), .B(a[122]), .Z(n19936) );
  NAND U20520 ( .A(n38343), .B(n19936), .Z(n19788) );
  AND U20521 ( .A(n19789), .B(n19788), .Z(n19997) );
  NAND U20522 ( .A(n183), .B(n19790), .Z(n19792) );
  XOR U20523 ( .A(b[5]), .B(a[144]), .Z(n19939) );
  NAND U20524 ( .A(n36296), .B(n19939), .Z(n19791) );
  AND U20525 ( .A(n19792), .B(n19791), .Z(n19995) );
  NAND U20526 ( .A(n190), .B(n19793), .Z(n19795) );
  XOR U20527 ( .A(b[19]), .B(a[130]), .Z(n19942) );
  NAND U20528 ( .A(n37821), .B(n19942), .Z(n19794) );
  NAND U20529 ( .A(n19795), .B(n19794), .Z(n19994) );
  XNOR U20530 ( .A(n19995), .B(n19994), .Z(n19996) );
  XNOR U20531 ( .A(n19997), .B(n19996), .Z(n19988) );
  NAND U20532 ( .A(n38470), .B(n19796), .Z(n19798) );
  XOR U20533 ( .A(b[31]), .B(a[118]), .Z(n19945) );
  NAND U20534 ( .A(n38453), .B(n19945), .Z(n19797) );
  AND U20535 ( .A(n19798), .B(n19797), .Z(n19957) );
  NAND U20536 ( .A(n181), .B(n19799), .Z(n19801) );
  XOR U20537 ( .A(b[3]), .B(a[146]), .Z(n19948) );
  NAND U20538 ( .A(n182), .B(n19948), .Z(n19800) );
  AND U20539 ( .A(n19801), .B(n19800), .Z(n19955) );
  NAND U20540 ( .A(n189), .B(n19802), .Z(n19804) );
  XOR U20541 ( .A(b[17]), .B(a[132]), .Z(n19951) );
  NAND U20542 ( .A(n37652), .B(n19951), .Z(n19803) );
  NAND U20543 ( .A(n19804), .B(n19803), .Z(n19954) );
  XNOR U20544 ( .A(n19955), .B(n19954), .Z(n19956) );
  XOR U20545 ( .A(n19957), .B(n19956), .Z(n19989) );
  XOR U20546 ( .A(n19988), .B(n19989), .Z(n19991) );
  XOR U20547 ( .A(n19990), .B(n19991), .Z(n19925) );
  NANDN U20548 ( .A(n19806), .B(n19805), .Z(n19810) );
  NANDN U20549 ( .A(n19808), .B(n19807), .Z(n19809) );
  AND U20550 ( .A(n19810), .B(n19809), .Z(n19978) );
  NANDN U20551 ( .A(n19812), .B(n19811), .Z(n19816) );
  NANDN U20552 ( .A(n19814), .B(n19813), .Z(n19815) );
  NAND U20553 ( .A(n19816), .B(n19815), .Z(n19979) );
  XNOR U20554 ( .A(n19978), .B(n19979), .Z(n19980) );
  NANDN U20555 ( .A(n19818), .B(n19817), .Z(n19822) );
  NANDN U20556 ( .A(n19820), .B(n19819), .Z(n19821) );
  NAND U20557 ( .A(n19822), .B(n19821), .Z(n19981) );
  XNOR U20558 ( .A(n19980), .B(n19981), .Z(n19924) );
  XNOR U20559 ( .A(n19925), .B(n19924), .Z(n19927) );
  NANDN U20560 ( .A(n19824), .B(n19823), .Z(n19828) );
  NANDN U20561 ( .A(n19826), .B(n19825), .Z(n19827) );
  AND U20562 ( .A(n19828), .B(n19827), .Z(n19926) );
  XOR U20563 ( .A(n19927), .B(n19926), .Z(n20039) );
  NANDN U20564 ( .A(n19830), .B(n19829), .Z(n19834) );
  NANDN U20565 ( .A(n19832), .B(n19831), .Z(n19833) );
  AND U20566 ( .A(n19834), .B(n19833), .Z(n20036) );
  NANDN U20567 ( .A(n19836), .B(n19835), .Z(n19840) );
  NANDN U20568 ( .A(n19838), .B(n19837), .Z(n19839) );
  AND U20569 ( .A(n19840), .B(n19839), .Z(n19921) );
  NANDN U20570 ( .A(n19842), .B(n19841), .Z(n19846) );
  OR U20571 ( .A(n19844), .B(n19843), .Z(n19845) );
  AND U20572 ( .A(n19846), .B(n19845), .Z(n19919) );
  NANDN U20573 ( .A(n19848), .B(n19847), .Z(n19852) );
  NANDN U20574 ( .A(n19850), .B(n19849), .Z(n19851) );
  AND U20575 ( .A(n19852), .B(n19851), .Z(n19985) );
  NANDN U20576 ( .A(n19854), .B(n19853), .Z(n19858) );
  NANDN U20577 ( .A(n19856), .B(n19855), .Z(n19857) );
  NAND U20578 ( .A(n19858), .B(n19857), .Z(n19984) );
  XNOR U20579 ( .A(n19985), .B(n19984), .Z(n19987) );
  NAND U20580 ( .A(b[0]), .B(a[148]), .Z(n19859) );
  XNOR U20581 ( .A(b[1]), .B(n19859), .Z(n19861) );
  NANDN U20582 ( .A(b[0]), .B(a[147]), .Z(n19860) );
  NAND U20583 ( .A(n19861), .B(n19860), .Z(n19933) );
  NAND U20584 ( .A(n194), .B(n19862), .Z(n19864) );
  XOR U20585 ( .A(b[29]), .B(a[120]), .Z(n20009) );
  NAND U20586 ( .A(n38456), .B(n20009), .Z(n19863) );
  AND U20587 ( .A(n19864), .B(n19863), .Z(n19931) );
  AND U20588 ( .A(b[31]), .B(a[116]), .Z(n19930) );
  XNOR U20589 ( .A(n19931), .B(n19930), .Z(n19932) );
  XNOR U20590 ( .A(n19933), .B(n19932), .Z(n19973) );
  NAND U20591 ( .A(n38185), .B(n19865), .Z(n19867) );
  XOR U20592 ( .A(b[23]), .B(a[126]), .Z(n20012) );
  NAND U20593 ( .A(n38132), .B(n20012), .Z(n19866) );
  AND U20594 ( .A(n19867), .B(n19866), .Z(n20002) );
  NAND U20595 ( .A(n184), .B(n19868), .Z(n19870) );
  XOR U20596 ( .A(b[7]), .B(a[142]), .Z(n20015) );
  NAND U20597 ( .A(n36592), .B(n20015), .Z(n19869) );
  AND U20598 ( .A(n19870), .B(n19869), .Z(n20001) );
  NAND U20599 ( .A(n38289), .B(n19871), .Z(n19873) );
  XOR U20600 ( .A(b[25]), .B(a[124]), .Z(n20018) );
  NAND U20601 ( .A(n38247), .B(n20018), .Z(n19872) );
  NAND U20602 ( .A(n19873), .B(n19872), .Z(n20000) );
  XOR U20603 ( .A(n20001), .B(n20000), .Z(n20003) );
  XOR U20604 ( .A(n20002), .B(n20003), .Z(n19972) );
  XOR U20605 ( .A(n19973), .B(n19972), .Z(n19975) );
  NAND U20606 ( .A(n187), .B(n19874), .Z(n19876) );
  XOR U20607 ( .A(b[13]), .B(a[136]), .Z(n20021) );
  NAND U20608 ( .A(n37295), .B(n20021), .Z(n19875) );
  AND U20609 ( .A(n19876), .B(n19875), .Z(n19967) );
  NAND U20610 ( .A(n186), .B(n19877), .Z(n19879) );
  XOR U20611 ( .A(b[11]), .B(a[138]), .Z(n20024) );
  NAND U20612 ( .A(n37097), .B(n20024), .Z(n19878) );
  NAND U20613 ( .A(n19879), .B(n19878), .Z(n19966) );
  XNOR U20614 ( .A(n19967), .B(n19966), .Z(n19969) );
  NAND U20615 ( .A(n188), .B(n19880), .Z(n19882) );
  XOR U20616 ( .A(b[15]), .B(a[134]), .Z(n20027) );
  NAND U20617 ( .A(n37382), .B(n20027), .Z(n19881) );
  AND U20618 ( .A(n19882), .B(n19881), .Z(n19963) );
  NAND U20619 ( .A(n38064), .B(n19883), .Z(n19885) );
  XOR U20620 ( .A(b[21]), .B(a[128]), .Z(n20030) );
  NAND U20621 ( .A(n37993), .B(n20030), .Z(n19884) );
  AND U20622 ( .A(n19885), .B(n19884), .Z(n19961) );
  NAND U20623 ( .A(n185), .B(n19886), .Z(n19888) );
  XOR U20624 ( .A(b[9]), .B(a[140]), .Z(n20033) );
  NAND U20625 ( .A(n36805), .B(n20033), .Z(n19887) );
  NAND U20626 ( .A(n19888), .B(n19887), .Z(n19960) );
  XNOR U20627 ( .A(n19961), .B(n19960), .Z(n19962) );
  XNOR U20628 ( .A(n19963), .B(n19962), .Z(n19968) );
  XOR U20629 ( .A(n19969), .B(n19968), .Z(n19974) );
  XNOR U20630 ( .A(n19975), .B(n19974), .Z(n19986) );
  XNOR U20631 ( .A(n19987), .B(n19986), .Z(n19918) );
  XNOR U20632 ( .A(n19919), .B(n19918), .Z(n19920) );
  XOR U20633 ( .A(n19921), .B(n19920), .Z(n20037) );
  XNOR U20634 ( .A(n20036), .B(n20037), .Z(n20038) );
  XNOR U20635 ( .A(n20039), .B(n20038), .Z(n19914) );
  XOR U20636 ( .A(n19915), .B(n19914), .Z(n19907) );
  NANDN U20637 ( .A(n19890), .B(n19889), .Z(n19894) );
  NANDN U20638 ( .A(n19892), .B(n19891), .Z(n19893) );
  AND U20639 ( .A(n19894), .B(n19893), .Z(n19906) );
  XOR U20640 ( .A(n19907), .B(n19906), .Z(n19909) );
  XNOR U20641 ( .A(n19908), .B(n19909), .Z(n19900) );
  XNOR U20642 ( .A(n19901), .B(n19900), .Z(n19902) );
  XNOR U20643 ( .A(n19903), .B(n19902), .Z(n20042) );
  XNOR U20644 ( .A(sreg[372]), .B(n20042), .Z(n20044) );
  NANDN U20645 ( .A(sreg[371]), .B(n19895), .Z(n19899) );
  NAND U20646 ( .A(n19897), .B(n19896), .Z(n19898) );
  NAND U20647 ( .A(n19899), .B(n19898), .Z(n20043) );
  XNOR U20648 ( .A(n20044), .B(n20043), .Z(c[372]) );
  NANDN U20649 ( .A(n19901), .B(n19900), .Z(n19905) );
  NANDN U20650 ( .A(n19903), .B(n19902), .Z(n19904) );
  AND U20651 ( .A(n19905), .B(n19904), .Z(n20050) );
  NANDN U20652 ( .A(n19907), .B(n19906), .Z(n19911) );
  NANDN U20653 ( .A(n19909), .B(n19908), .Z(n19910) );
  AND U20654 ( .A(n19911), .B(n19910), .Z(n20048) );
  NANDN U20655 ( .A(n19913), .B(n19912), .Z(n19917) );
  NAND U20656 ( .A(n19915), .B(n19914), .Z(n19916) );
  AND U20657 ( .A(n19917), .B(n19916), .Z(n20055) );
  NANDN U20658 ( .A(n19919), .B(n19918), .Z(n19923) );
  NANDN U20659 ( .A(n19921), .B(n19920), .Z(n19922) );
  AND U20660 ( .A(n19923), .B(n19922), .Z(n20060) );
  NANDN U20661 ( .A(n19925), .B(n19924), .Z(n19929) );
  NAND U20662 ( .A(n19927), .B(n19926), .Z(n19928) );
  AND U20663 ( .A(n19929), .B(n19928), .Z(n20059) );
  XNOR U20664 ( .A(n20060), .B(n20059), .Z(n20062) );
  NANDN U20665 ( .A(n19931), .B(n19930), .Z(n19935) );
  NANDN U20666 ( .A(n19933), .B(n19932), .Z(n19934) );
  AND U20667 ( .A(n19935), .B(n19934), .Z(n20127) );
  NAND U20668 ( .A(n38385), .B(n19936), .Z(n19938) );
  XOR U20669 ( .A(b[27]), .B(a[123]), .Z(n20071) );
  NAND U20670 ( .A(n38343), .B(n20071), .Z(n19937) );
  AND U20671 ( .A(n19938), .B(n19937), .Z(n20134) );
  NAND U20672 ( .A(n183), .B(n19939), .Z(n19941) );
  XOR U20673 ( .A(b[5]), .B(a[145]), .Z(n20074) );
  NAND U20674 ( .A(n36296), .B(n20074), .Z(n19940) );
  AND U20675 ( .A(n19941), .B(n19940), .Z(n20132) );
  NAND U20676 ( .A(n190), .B(n19942), .Z(n19944) );
  XOR U20677 ( .A(b[19]), .B(a[131]), .Z(n20077) );
  NAND U20678 ( .A(n37821), .B(n20077), .Z(n19943) );
  NAND U20679 ( .A(n19944), .B(n19943), .Z(n20131) );
  XNOR U20680 ( .A(n20132), .B(n20131), .Z(n20133) );
  XNOR U20681 ( .A(n20134), .B(n20133), .Z(n20125) );
  NAND U20682 ( .A(n38470), .B(n19945), .Z(n19947) );
  XOR U20683 ( .A(b[31]), .B(a[119]), .Z(n20080) );
  NAND U20684 ( .A(n38453), .B(n20080), .Z(n19946) );
  AND U20685 ( .A(n19947), .B(n19946), .Z(n20092) );
  NAND U20686 ( .A(n181), .B(n19948), .Z(n19950) );
  XOR U20687 ( .A(b[3]), .B(a[147]), .Z(n20083) );
  NAND U20688 ( .A(n182), .B(n20083), .Z(n19949) );
  AND U20689 ( .A(n19950), .B(n19949), .Z(n20090) );
  NAND U20690 ( .A(n189), .B(n19951), .Z(n19953) );
  XOR U20691 ( .A(b[17]), .B(a[133]), .Z(n20086) );
  NAND U20692 ( .A(n37652), .B(n20086), .Z(n19952) );
  NAND U20693 ( .A(n19953), .B(n19952), .Z(n20089) );
  XNOR U20694 ( .A(n20090), .B(n20089), .Z(n20091) );
  XOR U20695 ( .A(n20092), .B(n20091), .Z(n20126) );
  XOR U20696 ( .A(n20125), .B(n20126), .Z(n20128) );
  XOR U20697 ( .A(n20127), .B(n20128), .Z(n20174) );
  NANDN U20698 ( .A(n19955), .B(n19954), .Z(n19959) );
  NANDN U20699 ( .A(n19957), .B(n19956), .Z(n19958) );
  AND U20700 ( .A(n19959), .B(n19958), .Z(n20113) );
  NANDN U20701 ( .A(n19961), .B(n19960), .Z(n19965) );
  NANDN U20702 ( .A(n19963), .B(n19962), .Z(n19964) );
  NAND U20703 ( .A(n19965), .B(n19964), .Z(n20114) );
  XNOR U20704 ( .A(n20113), .B(n20114), .Z(n20115) );
  NANDN U20705 ( .A(n19967), .B(n19966), .Z(n19971) );
  NAND U20706 ( .A(n19969), .B(n19968), .Z(n19970) );
  NAND U20707 ( .A(n19971), .B(n19970), .Z(n20116) );
  XNOR U20708 ( .A(n20115), .B(n20116), .Z(n20173) );
  XNOR U20709 ( .A(n20174), .B(n20173), .Z(n20176) );
  NAND U20710 ( .A(n19973), .B(n19972), .Z(n19977) );
  NAND U20711 ( .A(n19975), .B(n19974), .Z(n19976) );
  AND U20712 ( .A(n19977), .B(n19976), .Z(n20175) );
  XOR U20713 ( .A(n20176), .B(n20175), .Z(n20188) );
  NANDN U20714 ( .A(n19979), .B(n19978), .Z(n19983) );
  NANDN U20715 ( .A(n19981), .B(n19980), .Z(n19982) );
  AND U20716 ( .A(n19983), .B(n19982), .Z(n20185) );
  NANDN U20717 ( .A(n19989), .B(n19988), .Z(n19993) );
  OR U20718 ( .A(n19991), .B(n19990), .Z(n19992) );
  AND U20719 ( .A(n19993), .B(n19992), .Z(n20180) );
  NANDN U20720 ( .A(n19995), .B(n19994), .Z(n19999) );
  NANDN U20721 ( .A(n19997), .B(n19996), .Z(n19998) );
  AND U20722 ( .A(n19999), .B(n19998), .Z(n20120) );
  NANDN U20723 ( .A(n20001), .B(n20000), .Z(n20005) );
  OR U20724 ( .A(n20003), .B(n20002), .Z(n20004) );
  NAND U20725 ( .A(n20005), .B(n20004), .Z(n20119) );
  XNOR U20726 ( .A(n20120), .B(n20119), .Z(n20121) );
  NAND U20727 ( .A(b[0]), .B(a[149]), .Z(n20006) );
  XNOR U20728 ( .A(b[1]), .B(n20006), .Z(n20008) );
  NANDN U20729 ( .A(b[0]), .B(a[148]), .Z(n20007) );
  NAND U20730 ( .A(n20008), .B(n20007), .Z(n20068) );
  NAND U20731 ( .A(n194), .B(n20009), .Z(n20011) );
  XOR U20732 ( .A(b[29]), .B(a[121]), .Z(n20146) );
  NAND U20733 ( .A(n38456), .B(n20146), .Z(n20010) );
  AND U20734 ( .A(n20011), .B(n20010), .Z(n20066) );
  AND U20735 ( .A(b[31]), .B(a[117]), .Z(n20065) );
  XNOR U20736 ( .A(n20066), .B(n20065), .Z(n20067) );
  XNOR U20737 ( .A(n20068), .B(n20067), .Z(n20107) );
  NAND U20738 ( .A(n38185), .B(n20012), .Z(n20014) );
  XOR U20739 ( .A(b[23]), .B(a[127]), .Z(n20149) );
  NAND U20740 ( .A(n38132), .B(n20149), .Z(n20013) );
  AND U20741 ( .A(n20014), .B(n20013), .Z(n20140) );
  NAND U20742 ( .A(n184), .B(n20015), .Z(n20017) );
  XOR U20743 ( .A(b[7]), .B(a[143]), .Z(n20152) );
  NAND U20744 ( .A(n36592), .B(n20152), .Z(n20016) );
  AND U20745 ( .A(n20017), .B(n20016), .Z(n20138) );
  NAND U20746 ( .A(n38289), .B(n20018), .Z(n20020) );
  XOR U20747 ( .A(b[25]), .B(a[125]), .Z(n20155) );
  NAND U20748 ( .A(n38247), .B(n20155), .Z(n20019) );
  NAND U20749 ( .A(n20020), .B(n20019), .Z(n20137) );
  XNOR U20750 ( .A(n20138), .B(n20137), .Z(n20139) );
  XOR U20751 ( .A(n20140), .B(n20139), .Z(n20108) );
  XNOR U20752 ( .A(n20107), .B(n20108), .Z(n20109) );
  NAND U20753 ( .A(n187), .B(n20021), .Z(n20023) );
  XOR U20754 ( .A(b[13]), .B(a[137]), .Z(n20158) );
  NAND U20755 ( .A(n37295), .B(n20158), .Z(n20022) );
  AND U20756 ( .A(n20023), .B(n20022), .Z(n20102) );
  NAND U20757 ( .A(n186), .B(n20024), .Z(n20026) );
  XOR U20758 ( .A(b[11]), .B(a[139]), .Z(n20161) );
  NAND U20759 ( .A(n37097), .B(n20161), .Z(n20025) );
  NAND U20760 ( .A(n20026), .B(n20025), .Z(n20101) );
  XNOR U20761 ( .A(n20102), .B(n20101), .Z(n20103) );
  NAND U20762 ( .A(n188), .B(n20027), .Z(n20029) );
  XOR U20763 ( .A(b[15]), .B(a[135]), .Z(n20164) );
  NAND U20764 ( .A(n37382), .B(n20164), .Z(n20028) );
  AND U20765 ( .A(n20029), .B(n20028), .Z(n20098) );
  NAND U20766 ( .A(n38064), .B(n20030), .Z(n20032) );
  XOR U20767 ( .A(b[21]), .B(a[129]), .Z(n20167) );
  NAND U20768 ( .A(n37993), .B(n20167), .Z(n20031) );
  AND U20769 ( .A(n20032), .B(n20031), .Z(n20096) );
  NAND U20770 ( .A(n185), .B(n20033), .Z(n20035) );
  XOR U20771 ( .A(b[9]), .B(a[141]), .Z(n20170) );
  NAND U20772 ( .A(n36805), .B(n20170), .Z(n20034) );
  NAND U20773 ( .A(n20035), .B(n20034), .Z(n20095) );
  XNOR U20774 ( .A(n20096), .B(n20095), .Z(n20097) );
  XOR U20775 ( .A(n20098), .B(n20097), .Z(n20104) );
  XOR U20776 ( .A(n20103), .B(n20104), .Z(n20110) );
  XOR U20777 ( .A(n20109), .B(n20110), .Z(n20122) );
  XNOR U20778 ( .A(n20121), .B(n20122), .Z(n20179) );
  XNOR U20779 ( .A(n20180), .B(n20179), .Z(n20181) );
  XOR U20780 ( .A(n20182), .B(n20181), .Z(n20186) );
  XNOR U20781 ( .A(n20185), .B(n20186), .Z(n20187) );
  XNOR U20782 ( .A(n20188), .B(n20187), .Z(n20061) );
  XOR U20783 ( .A(n20062), .B(n20061), .Z(n20054) );
  NANDN U20784 ( .A(n20037), .B(n20036), .Z(n20041) );
  NANDN U20785 ( .A(n20039), .B(n20038), .Z(n20040) );
  AND U20786 ( .A(n20041), .B(n20040), .Z(n20053) );
  XOR U20787 ( .A(n20054), .B(n20053), .Z(n20056) );
  XNOR U20788 ( .A(n20055), .B(n20056), .Z(n20047) );
  XNOR U20789 ( .A(n20048), .B(n20047), .Z(n20049) );
  XNOR U20790 ( .A(n20050), .B(n20049), .Z(n20191) );
  XNOR U20791 ( .A(sreg[373]), .B(n20191), .Z(n20193) );
  NANDN U20792 ( .A(sreg[372]), .B(n20042), .Z(n20046) );
  NAND U20793 ( .A(n20044), .B(n20043), .Z(n20045) );
  NAND U20794 ( .A(n20046), .B(n20045), .Z(n20192) );
  XNOR U20795 ( .A(n20193), .B(n20192), .Z(c[373]) );
  NANDN U20796 ( .A(n20048), .B(n20047), .Z(n20052) );
  NANDN U20797 ( .A(n20050), .B(n20049), .Z(n20051) );
  AND U20798 ( .A(n20052), .B(n20051), .Z(n20199) );
  NANDN U20799 ( .A(n20054), .B(n20053), .Z(n20058) );
  NANDN U20800 ( .A(n20056), .B(n20055), .Z(n20057) );
  AND U20801 ( .A(n20058), .B(n20057), .Z(n20197) );
  NANDN U20802 ( .A(n20060), .B(n20059), .Z(n20064) );
  NAND U20803 ( .A(n20062), .B(n20061), .Z(n20063) );
  AND U20804 ( .A(n20064), .B(n20063), .Z(n20204) );
  NANDN U20805 ( .A(n20066), .B(n20065), .Z(n20070) );
  NANDN U20806 ( .A(n20068), .B(n20067), .Z(n20069) );
  AND U20807 ( .A(n20070), .B(n20069), .Z(n20288) );
  NAND U20808 ( .A(n38385), .B(n20071), .Z(n20073) );
  XOR U20809 ( .A(b[27]), .B(a[124]), .Z(n20232) );
  NAND U20810 ( .A(n38343), .B(n20232), .Z(n20072) );
  AND U20811 ( .A(n20073), .B(n20072), .Z(n20295) );
  NAND U20812 ( .A(n183), .B(n20074), .Z(n20076) );
  XOR U20813 ( .A(b[5]), .B(a[146]), .Z(n20235) );
  NAND U20814 ( .A(n36296), .B(n20235), .Z(n20075) );
  AND U20815 ( .A(n20076), .B(n20075), .Z(n20293) );
  NAND U20816 ( .A(n190), .B(n20077), .Z(n20079) );
  XOR U20817 ( .A(b[19]), .B(a[132]), .Z(n20238) );
  NAND U20818 ( .A(n37821), .B(n20238), .Z(n20078) );
  NAND U20819 ( .A(n20079), .B(n20078), .Z(n20292) );
  XNOR U20820 ( .A(n20293), .B(n20292), .Z(n20294) );
  XNOR U20821 ( .A(n20295), .B(n20294), .Z(n20286) );
  NAND U20822 ( .A(n38470), .B(n20080), .Z(n20082) );
  XOR U20823 ( .A(b[31]), .B(a[120]), .Z(n20241) );
  NAND U20824 ( .A(n38453), .B(n20241), .Z(n20081) );
  AND U20825 ( .A(n20082), .B(n20081), .Z(n20253) );
  NAND U20826 ( .A(n181), .B(n20083), .Z(n20085) );
  XOR U20827 ( .A(b[3]), .B(a[148]), .Z(n20244) );
  NAND U20828 ( .A(n182), .B(n20244), .Z(n20084) );
  AND U20829 ( .A(n20085), .B(n20084), .Z(n20251) );
  NAND U20830 ( .A(n189), .B(n20086), .Z(n20088) );
  XOR U20831 ( .A(b[17]), .B(a[134]), .Z(n20247) );
  NAND U20832 ( .A(n37652), .B(n20247), .Z(n20087) );
  NAND U20833 ( .A(n20088), .B(n20087), .Z(n20250) );
  XNOR U20834 ( .A(n20251), .B(n20250), .Z(n20252) );
  XOR U20835 ( .A(n20253), .B(n20252), .Z(n20287) );
  XOR U20836 ( .A(n20286), .B(n20287), .Z(n20289) );
  XOR U20837 ( .A(n20288), .B(n20289), .Z(n20221) );
  NANDN U20838 ( .A(n20090), .B(n20089), .Z(n20094) );
  NANDN U20839 ( .A(n20092), .B(n20091), .Z(n20093) );
  AND U20840 ( .A(n20094), .B(n20093), .Z(n20274) );
  NANDN U20841 ( .A(n20096), .B(n20095), .Z(n20100) );
  NANDN U20842 ( .A(n20098), .B(n20097), .Z(n20099) );
  NAND U20843 ( .A(n20100), .B(n20099), .Z(n20275) );
  XNOR U20844 ( .A(n20274), .B(n20275), .Z(n20276) );
  NANDN U20845 ( .A(n20102), .B(n20101), .Z(n20106) );
  NANDN U20846 ( .A(n20104), .B(n20103), .Z(n20105) );
  NAND U20847 ( .A(n20106), .B(n20105), .Z(n20277) );
  XNOR U20848 ( .A(n20276), .B(n20277), .Z(n20220) );
  XNOR U20849 ( .A(n20221), .B(n20220), .Z(n20223) );
  NANDN U20850 ( .A(n20108), .B(n20107), .Z(n20112) );
  NANDN U20851 ( .A(n20110), .B(n20109), .Z(n20111) );
  AND U20852 ( .A(n20112), .B(n20111), .Z(n20222) );
  XOR U20853 ( .A(n20223), .B(n20222), .Z(n20336) );
  NANDN U20854 ( .A(n20114), .B(n20113), .Z(n20118) );
  NANDN U20855 ( .A(n20116), .B(n20115), .Z(n20117) );
  AND U20856 ( .A(n20118), .B(n20117), .Z(n20334) );
  NANDN U20857 ( .A(n20120), .B(n20119), .Z(n20124) );
  NANDN U20858 ( .A(n20122), .B(n20121), .Z(n20123) );
  AND U20859 ( .A(n20124), .B(n20123), .Z(n20217) );
  NANDN U20860 ( .A(n20126), .B(n20125), .Z(n20130) );
  OR U20861 ( .A(n20128), .B(n20127), .Z(n20129) );
  AND U20862 ( .A(n20130), .B(n20129), .Z(n20215) );
  NANDN U20863 ( .A(n20132), .B(n20131), .Z(n20136) );
  NANDN U20864 ( .A(n20134), .B(n20133), .Z(n20135) );
  AND U20865 ( .A(n20136), .B(n20135), .Z(n20281) );
  NANDN U20866 ( .A(n20138), .B(n20137), .Z(n20142) );
  NANDN U20867 ( .A(n20140), .B(n20139), .Z(n20141) );
  NAND U20868 ( .A(n20142), .B(n20141), .Z(n20280) );
  XNOR U20869 ( .A(n20281), .B(n20280), .Z(n20282) );
  NAND U20870 ( .A(b[0]), .B(a[150]), .Z(n20143) );
  XNOR U20871 ( .A(b[1]), .B(n20143), .Z(n20145) );
  NANDN U20872 ( .A(b[0]), .B(a[149]), .Z(n20144) );
  NAND U20873 ( .A(n20145), .B(n20144), .Z(n20229) );
  NAND U20874 ( .A(n194), .B(n20146), .Z(n20148) );
  XOR U20875 ( .A(b[29]), .B(a[122]), .Z(n20304) );
  NAND U20876 ( .A(n38456), .B(n20304), .Z(n20147) );
  AND U20877 ( .A(n20148), .B(n20147), .Z(n20227) );
  AND U20878 ( .A(b[31]), .B(a[118]), .Z(n20226) );
  XNOR U20879 ( .A(n20227), .B(n20226), .Z(n20228) );
  XNOR U20880 ( .A(n20229), .B(n20228), .Z(n20268) );
  NAND U20881 ( .A(n38185), .B(n20149), .Z(n20151) );
  XOR U20882 ( .A(b[23]), .B(a[128]), .Z(n20310) );
  NAND U20883 ( .A(n38132), .B(n20310), .Z(n20150) );
  AND U20884 ( .A(n20151), .B(n20150), .Z(n20301) );
  NAND U20885 ( .A(n184), .B(n20152), .Z(n20154) );
  XOR U20886 ( .A(b[7]), .B(a[144]), .Z(n20313) );
  NAND U20887 ( .A(n36592), .B(n20313), .Z(n20153) );
  AND U20888 ( .A(n20154), .B(n20153), .Z(n20299) );
  NAND U20889 ( .A(n38289), .B(n20155), .Z(n20157) );
  XOR U20890 ( .A(b[25]), .B(a[126]), .Z(n20316) );
  NAND U20891 ( .A(n38247), .B(n20316), .Z(n20156) );
  NAND U20892 ( .A(n20157), .B(n20156), .Z(n20298) );
  XNOR U20893 ( .A(n20299), .B(n20298), .Z(n20300) );
  XOR U20894 ( .A(n20301), .B(n20300), .Z(n20269) );
  XNOR U20895 ( .A(n20268), .B(n20269), .Z(n20270) );
  NAND U20896 ( .A(n187), .B(n20158), .Z(n20160) );
  XOR U20897 ( .A(b[13]), .B(a[138]), .Z(n20319) );
  NAND U20898 ( .A(n37295), .B(n20319), .Z(n20159) );
  AND U20899 ( .A(n20160), .B(n20159), .Z(n20263) );
  NAND U20900 ( .A(n186), .B(n20161), .Z(n20163) );
  XOR U20901 ( .A(b[11]), .B(a[140]), .Z(n20322) );
  NAND U20902 ( .A(n37097), .B(n20322), .Z(n20162) );
  NAND U20903 ( .A(n20163), .B(n20162), .Z(n20262) );
  XNOR U20904 ( .A(n20263), .B(n20262), .Z(n20264) );
  NAND U20905 ( .A(n188), .B(n20164), .Z(n20166) );
  XOR U20906 ( .A(b[15]), .B(a[136]), .Z(n20325) );
  NAND U20907 ( .A(n37382), .B(n20325), .Z(n20165) );
  AND U20908 ( .A(n20166), .B(n20165), .Z(n20259) );
  NAND U20909 ( .A(n38064), .B(n20167), .Z(n20169) );
  XOR U20910 ( .A(b[21]), .B(a[130]), .Z(n20328) );
  NAND U20911 ( .A(n37993), .B(n20328), .Z(n20168) );
  AND U20912 ( .A(n20169), .B(n20168), .Z(n20257) );
  NAND U20913 ( .A(n185), .B(n20170), .Z(n20172) );
  XOR U20914 ( .A(b[9]), .B(a[142]), .Z(n20331) );
  NAND U20915 ( .A(n36805), .B(n20331), .Z(n20171) );
  NAND U20916 ( .A(n20172), .B(n20171), .Z(n20256) );
  XNOR U20917 ( .A(n20257), .B(n20256), .Z(n20258) );
  XOR U20918 ( .A(n20259), .B(n20258), .Z(n20265) );
  XOR U20919 ( .A(n20264), .B(n20265), .Z(n20271) );
  XOR U20920 ( .A(n20270), .B(n20271), .Z(n20283) );
  XNOR U20921 ( .A(n20282), .B(n20283), .Z(n20214) );
  XNOR U20922 ( .A(n20215), .B(n20214), .Z(n20216) );
  XOR U20923 ( .A(n20217), .B(n20216), .Z(n20335) );
  XOR U20924 ( .A(n20334), .B(n20335), .Z(n20337) );
  XOR U20925 ( .A(n20336), .B(n20337), .Z(n20211) );
  NANDN U20926 ( .A(n20174), .B(n20173), .Z(n20178) );
  NAND U20927 ( .A(n20176), .B(n20175), .Z(n20177) );
  AND U20928 ( .A(n20178), .B(n20177), .Z(n20209) );
  NANDN U20929 ( .A(n20180), .B(n20179), .Z(n20184) );
  NANDN U20930 ( .A(n20182), .B(n20181), .Z(n20183) );
  AND U20931 ( .A(n20184), .B(n20183), .Z(n20208) );
  XNOR U20932 ( .A(n20209), .B(n20208), .Z(n20210) );
  XNOR U20933 ( .A(n20211), .B(n20210), .Z(n20202) );
  NANDN U20934 ( .A(n20186), .B(n20185), .Z(n20190) );
  NANDN U20935 ( .A(n20188), .B(n20187), .Z(n20189) );
  NAND U20936 ( .A(n20190), .B(n20189), .Z(n20203) );
  XOR U20937 ( .A(n20202), .B(n20203), .Z(n20205) );
  XNOR U20938 ( .A(n20204), .B(n20205), .Z(n20196) );
  XNOR U20939 ( .A(n20197), .B(n20196), .Z(n20198) );
  XNOR U20940 ( .A(n20199), .B(n20198), .Z(n20340) );
  XNOR U20941 ( .A(sreg[374]), .B(n20340), .Z(n20342) );
  NANDN U20942 ( .A(sreg[373]), .B(n20191), .Z(n20195) );
  NAND U20943 ( .A(n20193), .B(n20192), .Z(n20194) );
  NAND U20944 ( .A(n20195), .B(n20194), .Z(n20341) );
  XNOR U20945 ( .A(n20342), .B(n20341), .Z(c[374]) );
  NANDN U20946 ( .A(n20197), .B(n20196), .Z(n20201) );
  NANDN U20947 ( .A(n20199), .B(n20198), .Z(n20200) );
  AND U20948 ( .A(n20201), .B(n20200), .Z(n20348) );
  NANDN U20949 ( .A(n20203), .B(n20202), .Z(n20207) );
  NANDN U20950 ( .A(n20205), .B(n20204), .Z(n20206) );
  AND U20951 ( .A(n20207), .B(n20206), .Z(n20346) );
  NANDN U20952 ( .A(n20209), .B(n20208), .Z(n20213) );
  NANDN U20953 ( .A(n20211), .B(n20210), .Z(n20212) );
  AND U20954 ( .A(n20213), .B(n20212), .Z(n20354) );
  NANDN U20955 ( .A(n20215), .B(n20214), .Z(n20219) );
  NANDN U20956 ( .A(n20217), .B(n20216), .Z(n20218) );
  AND U20957 ( .A(n20219), .B(n20218), .Z(n20358) );
  NANDN U20958 ( .A(n20221), .B(n20220), .Z(n20225) );
  NAND U20959 ( .A(n20223), .B(n20222), .Z(n20224) );
  AND U20960 ( .A(n20225), .B(n20224), .Z(n20357) );
  XNOR U20961 ( .A(n20358), .B(n20357), .Z(n20360) );
  NANDN U20962 ( .A(n20227), .B(n20226), .Z(n20231) );
  NANDN U20963 ( .A(n20229), .B(n20228), .Z(n20230) );
  AND U20964 ( .A(n20231), .B(n20230), .Z(n20437) );
  NAND U20965 ( .A(n38385), .B(n20232), .Z(n20234) );
  XOR U20966 ( .A(b[27]), .B(a[125]), .Z(n20381) );
  NAND U20967 ( .A(n38343), .B(n20381), .Z(n20233) );
  AND U20968 ( .A(n20234), .B(n20233), .Z(n20444) );
  NAND U20969 ( .A(n183), .B(n20235), .Z(n20237) );
  XOR U20970 ( .A(b[5]), .B(a[147]), .Z(n20384) );
  NAND U20971 ( .A(n36296), .B(n20384), .Z(n20236) );
  AND U20972 ( .A(n20237), .B(n20236), .Z(n20442) );
  NAND U20973 ( .A(n190), .B(n20238), .Z(n20240) );
  XOR U20974 ( .A(b[19]), .B(a[133]), .Z(n20387) );
  NAND U20975 ( .A(n37821), .B(n20387), .Z(n20239) );
  NAND U20976 ( .A(n20240), .B(n20239), .Z(n20441) );
  XNOR U20977 ( .A(n20442), .B(n20441), .Z(n20443) );
  XNOR U20978 ( .A(n20444), .B(n20443), .Z(n20435) );
  NAND U20979 ( .A(n38470), .B(n20241), .Z(n20243) );
  XOR U20980 ( .A(b[31]), .B(a[121]), .Z(n20390) );
  NAND U20981 ( .A(n38453), .B(n20390), .Z(n20242) );
  AND U20982 ( .A(n20243), .B(n20242), .Z(n20402) );
  NAND U20983 ( .A(n181), .B(n20244), .Z(n20246) );
  XOR U20984 ( .A(b[3]), .B(a[149]), .Z(n20393) );
  NAND U20985 ( .A(n182), .B(n20393), .Z(n20245) );
  AND U20986 ( .A(n20246), .B(n20245), .Z(n20400) );
  NAND U20987 ( .A(n189), .B(n20247), .Z(n20249) );
  XOR U20988 ( .A(b[17]), .B(a[135]), .Z(n20396) );
  NAND U20989 ( .A(n37652), .B(n20396), .Z(n20248) );
  NAND U20990 ( .A(n20249), .B(n20248), .Z(n20399) );
  XNOR U20991 ( .A(n20400), .B(n20399), .Z(n20401) );
  XOR U20992 ( .A(n20402), .B(n20401), .Z(n20436) );
  XOR U20993 ( .A(n20435), .B(n20436), .Z(n20438) );
  XOR U20994 ( .A(n20437), .B(n20438), .Z(n20370) );
  NANDN U20995 ( .A(n20251), .B(n20250), .Z(n20255) );
  NANDN U20996 ( .A(n20253), .B(n20252), .Z(n20254) );
  AND U20997 ( .A(n20255), .B(n20254), .Z(n20423) );
  NANDN U20998 ( .A(n20257), .B(n20256), .Z(n20261) );
  NANDN U20999 ( .A(n20259), .B(n20258), .Z(n20260) );
  NAND U21000 ( .A(n20261), .B(n20260), .Z(n20424) );
  XNOR U21001 ( .A(n20423), .B(n20424), .Z(n20425) );
  NANDN U21002 ( .A(n20263), .B(n20262), .Z(n20267) );
  NANDN U21003 ( .A(n20265), .B(n20264), .Z(n20266) );
  NAND U21004 ( .A(n20267), .B(n20266), .Z(n20426) );
  XNOR U21005 ( .A(n20425), .B(n20426), .Z(n20369) );
  XNOR U21006 ( .A(n20370), .B(n20369), .Z(n20372) );
  NANDN U21007 ( .A(n20269), .B(n20268), .Z(n20273) );
  NANDN U21008 ( .A(n20271), .B(n20270), .Z(n20272) );
  AND U21009 ( .A(n20273), .B(n20272), .Z(n20371) );
  XOR U21010 ( .A(n20372), .B(n20371), .Z(n20486) );
  NANDN U21011 ( .A(n20275), .B(n20274), .Z(n20279) );
  NANDN U21012 ( .A(n20277), .B(n20276), .Z(n20278) );
  AND U21013 ( .A(n20279), .B(n20278), .Z(n20483) );
  NANDN U21014 ( .A(n20281), .B(n20280), .Z(n20285) );
  NANDN U21015 ( .A(n20283), .B(n20282), .Z(n20284) );
  AND U21016 ( .A(n20285), .B(n20284), .Z(n20366) );
  NANDN U21017 ( .A(n20287), .B(n20286), .Z(n20291) );
  OR U21018 ( .A(n20289), .B(n20288), .Z(n20290) );
  AND U21019 ( .A(n20291), .B(n20290), .Z(n20364) );
  NANDN U21020 ( .A(n20293), .B(n20292), .Z(n20297) );
  NANDN U21021 ( .A(n20295), .B(n20294), .Z(n20296) );
  AND U21022 ( .A(n20297), .B(n20296), .Z(n20430) );
  NANDN U21023 ( .A(n20299), .B(n20298), .Z(n20303) );
  NANDN U21024 ( .A(n20301), .B(n20300), .Z(n20302) );
  NAND U21025 ( .A(n20303), .B(n20302), .Z(n20429) );
  XNOR U21026 ( .A(n20430), .B(n20429), .Z(n20431) );
  NAND U21027 ( .A(n194), .B(n20304), .Z(n20306) );
  XOR U21028 ( .A(b[29]), .B(a[123]), .Z(n20456) );
  NAND U21029 ( .A(n38456), .B(n20456), .Z(n20305) );
  AND U21030 ( .A(n20306), .B(n20305), .Z(n20376) );
  AND U21031 ( .A(b[31]), .B(a[119]), .Z(n20375) );
  XNOR U21032 ( .A(n20376), .B(n20375), .Z(n20377) );
  NAND U21033 ( .A(b[0]), .B(a[151]), .Z(n20307) );
  XNOR U21034 ( .A(b[1]), .B(n20307), .Z(n20309) );
  NANDN U21035 ( .A(b[0]), .B(a[150]), .Z(n20308) );
  NAND U21036 ( .A(n20309), .B(n20308), .Z(n20378) );
  XNOR U21037 ( .A(n20377), .B(n20378), .Z(n20417) );
  NAND U21038 ( .A(n38185), .B(n20310), .Z(n20312) );
  XOR U21039 ( .A(b[23]), .B(a[129]), .Z(n20459) );
  NAND U21040 ( .A(n38132), .B(n20459), .Z(n20311) );
  AND U21041 ( .A(n20312), .B(n20311), .Z(n20450) );
  NAND U21042 ( .A(n184), .B(n20313), .Z(n20315) );
  XOR U21043 ( .A(b[7]), .B(a[145]), .Z(n20462) );
  NAND U21044 ( .A(n36592), .B(n20462), .Z(n20314) );
  AND U21045 ( .A(n20315), .B(n20314), .Z(n20448) );
  NAND U21046 ( .A(n38289), .B(n20316), .Z(n20318) );
  XOR U21047 ( .A(b[25]), .B(a[127]), .Z(n20465) );
  NAND U21048 ( .A(n38247), .B(n20465), .Z(n20317) );
  NAND U21049 ( .A(n20318), .B(n20317), .Z(n20447) );
  XNOR U21050 ( .A(n20448), .B(n20447), .Z(n20449) );
  XOR U21051 ( .A(n20450), .B(n20449), .Z(n20418) );
  XNOR U21052 ( .A(n20417), .B(n20418), .Z(n20419) );
  NAND U21053 ( .A(n187), .B(n20319), .Z(n20321) );
  XOR U21054 ( .A(b[13]), .B(a[139]), .Z(n20468) );
  NAND U21055 ( .A(n37295), .B(n20468), .Z(n20320) );
  AND U21056 ( .A(n20321), .B(n20320), .Z(n20412) );
  NAND U21057 ( .A(n186), .B(n20322), .Z(n20324) );
  XOR U21058 ( .A(b[11]), .B(a[141]), .Z(n20471) );
  NAND U21059 ( .A(n37097), .B(n20471), .Z(n20323) );
  NAND U21060 ( .A(n20324), .B(n20323), .Z(n20411) );
  XNOR U21061 ( .A(n20412), .B(n20411), .Z(n20413) );
  NAND U21062 ( .A(n188), .B(n20325), .Z(n20327) );
  XOR U21063 ( .A(b[15]), .B(a[137]), .Z(n20474) );
  NAND U21064 ( .A(n37382), .B(n20474), .Z(n20326) );
  AND U21065 ( .A(n20327), .B(n20326), .Z(n20408) );
  NAND U21066 ( .A(n38064), .B(n20328), .Z(n20330) );
  XOR U21067 ( .A(b[21]), .B(a[131]), .Z(n20477) );
  NAND U21068 ( .A(n37993), .B(n20477), .Z(n20329) );
  AND U21069 ( .A(n20330), .B(n20329), .Z(n20406) );
  NAND U21070 ( .A(n185), .B(n20331), .Z(n20333) );
  XOR U21071 ( .A(b[9]), .B(a[143]), .Z(n20480) );
  NAND U21072 ( .A(n36805), .B(n20480), .Z(n20332) );
  NAND U21073 ( .A(n20333), .B(n20332), .Z(n20405) );
  XNOR U21074 ( .A(n20406), .B(n20405), .Z(n20407) );
  XOR U21075 ( .A(n20408), .B(n20407), .Z(n20414) );
  XOR U21076 ( .A(n20413), .B(n20414), .Z(n20420) );
  XOR U21077 ( .A(n20419), .B(n20420), .Z(n20432) );
  XNOR U21078 ( .A(n20431), .B(n20432), .Z(n20363) );
  XNOR U21079 ( .A(n20364), .B(n20363), .Z(n20365) );
  XOR U21080 ( .A(n20366), .B(n20365), .Z(n20484) );
  XNOR U21081 ( .A(n20483), .B(n20484), .Z(n20485) );
  XNOR U21082 ( .A(n20486), .B(n20485), .Z(n20359) );
  XOR U21083 ( .A(n20360), .B(n20359), .Z(n20352) );
  NANDN U21084 ( .A(n20335), .B(n20334), .Z(n20339) );
  OR U21085 ( .A(n20337), .B(n20336), .Z(n20338) );
  AND U21086 ( .A(n20339), .B(n20338), .Z(n20351) );
  XNOR U21087 ( .A(n20352), .B(n20351), .Z(n20353) );
  XNOR U21088 ( .A(n20354), .B(n20353), .Z(n20345) );
  XNOR U21089 ( .A(n20346), .B(n20345), .Z(n20347) );
  XNOR U21090 ( .A(n20348), .B(n20347), .Z(n20489) );
  XNOR U21091 ( .A(sreg[375]), .B(n20489), .Z(n20491) );
  NANDN U21092 ( .A(sreg[374]), .B(n20340), .Z(n20344) );
  NAND U21093 ( .A(n20342), .B(n20341), .Z(n20343) );
  NAND U21094 ( .A(n20344), .B(n20343), .Z(n20490) );
  XNOR U21095 ( .A(n20491), .B(n20490), .Z(c[375]) );
  NANDN U21096 ( .A(n20346), .B(n20345), .Z(n20350) );
  NANDN U21097 ( .A(n20348), .B(n20347), .Z(n20349) );
  AND U21098 ( .A(n20350), .B(n20349), .Z(n20497) );
  NANDN U21099 ( .A(n20352), .B(n20351), .Z(n20356) );
  NANDN U21100 ( .A(n20354), .B(n20353), .Z(n20355) );
  AND U21101 ( .A(n20356), .B(n20355), .Z(n20495) );
  NANDN U21102 ( .A(n20358), .B(n20357), .Z(n20362) );
  NAND U21103 ( .A(n20360), .B(n20359), .Z(n20361) );
  AND U21104 ( .A(n20362), .B(n20361), .Z(n20502) );
  NANDN U21105 ( .A(n20364), .B(n20363), .Z(n20368) );
  NANDN U21106 ( .A(n20366), .B(n20365), .Z(n20367) );
  AND U21107 ( .A(n20368), .B(n20367), .Z(n20507) );
  NANDN U21108 ( .A(n20370), .B(n20369), .Z(n20374) );
  NAND U21109 ( .A(n20372), .B(n20371), .Z(n20373) );
  AND U21110 ( .A(n20374), .B(n20373), .Z(n20506) );
  XNOR U21111 ( .A(n20507), .B(n20506), .Z(n20509) );
  NANDN U21112 ( .A(n20376), .B(n20375), .Z(n20380) );
  NANDN U21113 ( .A(n20378), .B(n20377), .Z(n20379) );
  AND U21114 ( .A(n20380), .B(n20379), .Z(n20584) );
  NAND U21115 ( .A(n38385), .B(n20381), .Z(n20383) );
  XOR U21116 ( .A(b[27]), .B(a[126]), .Z(n20530) );
  NAND U21117 ( .A(n38343), .B(n20530), .Z(n20382) );
  AND U21118 ( .A(n20383), .B(n20382), .Z(n20591) );
  NAND U21119 ( .A(n183), .B(n20384), .Z(n20386) );
  XOR U21120 ( .A(b[5]), .B(a[148]), .Z(n20533) );
  NAND U21121 ( .A(n36296), .B(n20533), .Z(n20385) );
  AND U21122 ( .A(n20386), .B(n20385), .Z(n20589) );
  NAND U21123 ( .A(n190), .B(n20387), .Z(n20389) );
  XOR U21124 ( .A(b[19]), .B(a[134]), .Z(n20536) );
  NAND U21125 ( .A(n37821), .B(n20536), .Z(n20388) );
  NAND U21126 ( .A(n20389), .B(n20388), .Z(n20588) );
  XNOR U21127 ( .A(n20589), .B(n20588), .Z(n20590) );
  XNOR U21128 ( .A(n20591), .B(n20590), .Z(n20582) );
  NAND U21129 ( .A(n38470), .B(n20390), .Z(n20392) );
  XOR U21130 ( .A(b[31]), .B(a[122]), .Z(n20539) );
  NAND U21131 ( .A(n38453), .B(n20539), .Z(n20391) );
  AND U21132 ( .A(n20392), .B(n20391), .Z(n20551) );
  NAND U21133 ( .A(n181), .B(n20393), .Z(n20395) );
  XOR U21134 ( .A(b[3]), .B(a[150]), .Z(n20542) );
  NAND U21135 ( .A(n182), .B(n20542), .Z(n20394) );
  AND U21136 ( .A(n20395), .B(n20394), .Z(n20549) );
  NAND U21137 ( .A(n189), .B(n20396), .Z(n20398) );
  XOR U21138 ( .A(b[17]), .B(a[136]), .Z(n20545) );
  NAND U21139 ( .A(n37652), .B(n20545), .Z(n20397) );
  NAND U21140 ( .A(n20398), .B(n20397), .Z(n20548) );
  XNOR U21141 ( .A(n20549), .B(n20548), .Z(n20550) );
  XOR U21142 ( .A(n20551), .B(n20550), .Z(n20583) );
  XOR U21143 ( .A(n20582), .B(n20583), .Z(n20585) );
  XOR U21144 ( .A(n20584), .B(n20585), .Z(n20519) );
  NANDN U21145 ( .A(n20400), .B(n20399), .Z(n20404) );
  NANDN U21146 ( .A(n20402), .B(n20401), .Z(n20403) );
  AND U21147 ( .A(n20404), .B(n20403), .Z(n20572) );
  NANDN U21148 ( .A(n20406), .B(n20405), .Z(n20410) );
  NANDN U21149 ( .A(n20408), .B(n20407), .Z(n20409) );
  NAND U21150 ( .A(n20410), .B(n20409), .Z(n20573) );
  XNOR U21151 ( .A(n20572), .B(n20573), .Z(n20574) );
  NANDN U21152 ( .A(n20412), .B(n20411), .Z(n20416) );
  NANDN U21153 ( .A(n20414), .B(n20413), .Z(n20415) );
  NAND U21154 ( .A(n20416), .B(n20415), .Z(n20575) );
  XNOR U21155 ( .A(n20574), .B(n20575), .Z(n20518) );
  XNOR U21156 ( .A(n20519), .B(n20518), .Z(n20521) );
  NANDN U21157 ( .A(n20418), .B(n20417), .Z(n20422) );
  NANDN U21158 ( .A(n20420), .B(n20419), .Z(n20421) );
  AND U21159 ( .A(n20422), .B(n20421), .Z(n20520) );
  XOR U21160 ( .A(n20521), .B(n20520), .Z(n20633) );
  NANDN U21161 ( .A(n20424), .B(n20423), .Z(n20428) );
  NANDN U21162 ( .A(n20426), .B(n20425), .Z(n20427) );
  AND U21163 ( .A(n20428), .B(n20427), .Z(n20630) );
  NANDN U21164 ( .A(n20430), .B(n20429), .Z(n20434) );
  NANDN U21165 ( .A(n20432), .B(n20431), .Z(n20433) );
  AND U21166 ( .A(n20434), .B(n20433), .Z(n20515) );
  NANDN U21167 ( .A(n20436), .B(n20435), .Z(n20440) );
  OR U21168 ( .A(n20438), .B(n20437), .Z(n20439) );
  AND U21169 ( .A(n20440), .B(n20439), .Z(n20513) );
  NANDN U21170 ( .A(n20442), .B(n20441), .Z(n20446) );
  NANDN U21171 ( .A(n20444), .B(n20443), .Z(n20445) );
  AND U21172 ( .A(n20446), .B(n20445), .Z(n20579) );
  NANDN U21173 ( .A(n20448), .B(n20447), .Z(n20452) );
  NANDN U21174 ( .A(n20450), .B(n20449), .Z(n20451) );
  NAND U21175 ( .A(n20452), .B(n20451), .Z(n20578) );
  XNOR U21176 ( .A(n20579), .B(n20578), .Z(n20581) );
  NAND U21177 ( .A(b[0]), .B(a[152]), .Z(n20453) );
  XNOR U21178 ( .A(b[1]), .B(n20453), .Z(n20455) );
  NANDN U21179 ( .A(b[0]), .B(a[151]), .Z(n20454) );
  NAND U21180 ( .A(n20455), .B(n20454), .Z(n20527) );
  NAND U21181 ( .A(n194), .B(n20456), .Z(n20458) );
  XOR U21182 ( .A(b[29]), .B(a[124]), .Z(n20603) );
  NAND U21183 ( .A(n38456), .B(n20603), .Z(n20457) );
  AND U21184 ( .A(n20458), .B(n20457), .Z(n20525) );
  AND U21185 ( .A(b[31]), .B(a[120]), .Z(n20524) );
  XNOR U21186 ( .A(n20525), .B(n20524), .Z(n20526) );
  XNOR U21187 ( .A(n20527), .B(n20526), .Z(n20567) );
  NAND U21188 ( .A(n38185), .B(n20459), .Z(n20461) );
  XOR U21189 ( .A(b[23]), .B(a[130]), .Z(n20606) );
  NAND U21190 ( .A(n38132), .B(n20606), .Z(n20460) );
  AND U21191 ( .A(n20461), .B(n20460), .Z(n20596) );
  NAND U21192 ( .A(n184), .B(n20462), .Z(n20464) );
  XOR U21193 ( .A(b[7]), .B(a[146]), .Z(n20609) );
  NAND U21194 ( .A(n36592), .B(n20609), .Z(n20463) );
  AND U21195 ( .A(n20464), .B(n20463), .Z(n20595) );
  NAND U21196 ( .A(n38289), .B(n20465), .Z(n20467) );
  XOR U21197 ( .A(b[25]), .B(a[128]), .Z(n20612) );
  NAND U21198 ( .A(n38247), .B(n20612), .Z(n20466) );
  NAND U21199 ( .A(n20467), .B(n20466), .Z(n20594) );
  XOR U21200 ( .A(n20595), .B(n20594), .Z(n20597) );
  XOR U21201 ( .A(n20596), .B(n20597), .Z(n20566) );
  XOR U21202 ( .A(n20567), .B(n20566), .Z(n20569) );
  NAND U21203 ( .A(n187), .B(n20468), .Z(n20470) );
  XOR U21204 ( .A(b[13]), .B(a[140]), .Z(n20615) );
  NAND U21205 ( .A(n37295), .B(n20615), .Z(n20469) );
  AND U21206 ( .A(n20470), .B(n20469), .Z(n20561) );
  NAND U21207 ( .A(n186), .B(n20471), .Z(n20473) );
  XOR U21208 ( .A(b[11]), .B(a[142]), .Z(n20618) );
  NAND U21209 ( .A(n37097), .B(n20618), .Z(n20472) );
  NAND U21210 ( .A(n20473), .B(n20472), .Z(n20560) );
  XNOR U21211 ( .A(n20561), .B(n20560), .Z(n20563) );
  NAND U21212 ( .A(n188), .B(n20474), .Z(n20476) );
  XOR U21213 ( .A(b[15]), .B(a[138]), .Z(n20621) );
  NAND U21214 ( .A(n37382), .B(n20621), .Z(n20475) );
  AND U21215 ( .A(n20476), .B(n20475), .Z(n20557) );
  NAND U21216 ( .A(n38064), .B(n20477), .Z(n20479) );
  XOR U21217 ( .A(b[21]), .B(a[132]), .Z(n20624) );
  NAND U21218 ( .A(n37993), .B(n20624), .Z(n20478) );
  AND U21219 ( .A(n20479), .B(n20478), .Z(n20555) );
  NAND U21220 ( .A(n185), .B(n20480), .Z(n20482) );
  XOR U21221 ( .A(b[9]), .B(a[144]), .Z(n20627) );
  NAND U21222 ( .A(n36805), .B(n20627), .Z(n20481) );
  NAND U21223 ( .A(n20482), .B(n20481), .Z(n20554) );
  XNOR U21224 ( .A(n20555), .B(n20554), .Z(n20556) );
  XNOR U21225 ( .A(n20557), .B(n20556), .Z(n20562) );
  XOR U21226 ( .A(n20563), .B(n20562), .Z(n20568) );
  XNOR U21227 ( .A(n20569), .B(n20568), .Z(n20580) );
  XNOR U21228 ( .A(n20581), .B(n20580), .Z(n20512) );
  XNOR U21229 ( .A(n20513), .B(n20512), .Z(n20514) );
  XOR U21230 ( .A(n20515), .B(n20514), .Z(n20631) );
  XNOR U21231 ( .A(n20630), .B(n20631), .Z(n20632) );
  XNOR U21232 ( .A(n20633), .B(n20632), .Z(n20508) );
  XOR U21233 ( .A(n20509), .B(n20508), .Z(n20501) );
  NANDN U21234 ( .A(n20484), .B(n20483), .Z(n20488) );
  NANDN U21235 ( .A(n20486), .B(n20485), .Z(n20487) );
  AND U21236 ( .A(n20488), .B(n20487), .Z(n20500) );
  XOR U21237 ( .A(n20501), .B(n20500), .Z(n20503) );
  XNOR U21238 ( .A(n20502), .B(n20503), .Z(n20494) );
  XNOR U21239 ( .A(n20495), .B(n20494), .Z(n20496) );
  XNOR U21240 ( .A(n20497), .B(n20496), .Z(n20636) );
  XNOR U21241 ( .A(sreg[376]), .B(n20636), .Z(n20638) );
  NANDN U21242 ( .A(sreg[375]), .B(n20489), .Z(n20493) );
  NAND U21243 ( .A(n20491), .B(n20490), .Z(n20492) );
  NAND U21244 ( .A(n20493), .B(n20492), .Z(n20637) );
  XNOR U21245 ( .A(n20638), .B(n20637), .Z(c[376]) );
  NANDN U21246 ( .A(n20495), .B(n20494), .Z(n20499) );
  NANDN U21247 ( .A(n20497), .B(n20496), .Z(n20498) );
  AND U21248 ( .A(n20499), .B(n20498), .Z(n20644) );
  NANDN U21249 ( .A(n20501), .B(n20500), .Z(n20505) );
  NANDN U21250 ( .A(n20503), .B(n20502), .Z(n20504) );
  AND U21251 ( .A(n20505), .B(n20504), .Z(n20642) );
  NANDN U21252 ( .A(n20507), .B(n20506), .Z(n20511) );
  NAND U21253 ( .A(n20509), .B(n20508), .Z(n20510) );
  AND U21254 ( .A(n20511), .B(n20510), .Z(n20649) );
  NANDN U21255 ( .A(n20513), .B(n20512), .Z(n20517) );
  NANDN U21256 ( .A(n20515), .B(n20514), .Z(n20516) );
  AND U21257 ( .A(n20517), .B(n20516), .Z(n20778) );
  NANDN U21258 ( .A(n20519), .B(n20518), .Z(n20523) );
  NAND U21259 ( .A(n20521), .B(n20520), .Z(n20522) );
  AND U21260 ( .A(n20523), .B(n20522), .Z(n20777) );
  XNOR U21261 ( .A(n20778), .B(n20777), .Z(n20780) );
  NANDN U21262 ( .A(n20525), .B(n20524), .Z(n20529) );
  NANDN U21263 ( .A(n20527), .B(n20526), .Z(n20528) );
  AND U21264 ( .A(n20529), .B(n20528), .Z(n20713) );
  NAND U21265 ( .A(n38385), .B(n20530), .Z(n20532) );
  XOR U21266 ( .A(b[27]), .B(a[127]), .Z(n20659) );
  NAND U21267 ( .A(n38343), .B(n20659), .Z(n20531) );
  AND U21268 ( .A(n20532), .B(n20531), .Z(n20720) );
  NAND U21269 ( .A(n183), .B(n20533), .Z(n20535) );
  XOR U21270 ( .A(b[5]), .B(a[149]), .Z(n20662) );
  NAND U21271 ( .A(n36296), .B(n20662), .Z(n20534) );
  AND U21272 ( .A(n20535), .B(n20534), .Z(n20718) );
  NAND U21273 ( .A(n190), .B(n20536), .Z(n20538) );
  XOR U21274 ( .A(b[19]), .B(a[135]), .Z(n20665) );
  NAND U21275 ( .A(n37821), .B(n20665), .Z(n20537) );
  NAND U21276 ( .A(n20538), .B(n20537), .Z(n20717) );
  XNOR U21277 ( .A(n20718), .B(n20717), .Z(n20719) );
  XNOR U21278 ( .A(n20720), .B(n20719), .Z(n20711) );
  NAND U21279 ( .A(n38470), .B(n20539), .Z(n20541) );
  XOR U21280 ( .A(b[31]), .B(a[123]), .Z(n20668) );
  NAND U21281 ( .A(n38453), .B(n20668), .Z(n20540) );
  AND U21282 ( .A(n20541), .B(n20540), .Z(n20680) );
  NAND U21283 ( .A(n181), .B(n20542), .Z(n20544) );
  XOR U21284 ( .A(b[3]), .B(a[151]), .Z(n20671) );
  NAND U21285 ( .A(n182), .B(n20671), .Z(n20543) );
  AND U21286 ( .A(n20544), .B(n20543), .Z(n20678) );
  NAND U21287 ( .A(n189), .B(n20545), .Z(n20547) );
  XOR U21288 ( .A(b[17]), .B(a[137]), .Z(n20674) );
  NAND U21289 ( .A(n37652), .B(n20674), .Z(n20546) );
  NAND U21290 ( .A(n20547), .B(n20546), .Z(n20677) );
  XNOR U21291 ( .A(n20678), .B(n20677), .Z(n20679) );
  XOR U21292 ( .A(n20680), .B(n20679), .Z(n20712) );
  XOR U21293 ( .A(n20711), .B(n20712), .Z(n20714) );
  XOR U21294 ( .A(n20713), .B(n20714), .Z(n20760) );
  NANDN U21295 ( .A(n20549), .B(n20548), .Z(n20553) );
  NANDN U21296 ( .A(n20551), .B(n20550), .Z(n20552) );
  AND U21297 ( .A(n20553), .B(n20552), .Z(n20701) );
  NANDN U21298 ( .A(n20555), .B(n20554), .Z(n20559) );
  NANDN U21299 ( .A(n20557), .B(n20556), .Z(n20558) );
  NAND U21300 ( .A(n20559), .B(n20558), .Z(n20702) );
  XNOR U21301 ( .A(n20701), .B(n20702), .Z(n20703) );
  NANDN U21302 ( .A(n20561), .B(n20560), .Z(n20565) );
  NAND U21303 ( .A(n20563), .B(n20562), .Z(n20564) );
  NAND U21304 ( .A(n20565), .B(n20564), .Z(n20704) );
  XNOR U21305 ( .A(n20703), .B(n20704), .Z(n20759) );
  XNOR U21306 ( .A(n20760), .B(n20759), .Z(n20762) );
  NAND U21307 ( .A(n20567), .B(n20566), .Z(n20571) );
  NAND U21308 ( .A(n20569), .B(n20568), .Z(n20570) );
  AND U21309 ( .A(n20571), .B(n20570), .Z(n20761) );
  XOR U21310 ( .A(n20762), .B(n20761), .Z(n20774) );
  NANDN U21311 ( .A(n20573), .B(n20572), .Z(n20577) );
  NANDN U21312 ( .A(n20575), .B(n20574), .Z(n20576) );
  AND U21313 ( .A(n20577), .B(n20576), .Z(n20771) );
  NANDN U21314 ( .A(n20583), .B(n20582), .Z(n20587) );
  OR U21315 ( .A(n20585), .B(n20584), .Z(n20586) );
  AND U21316 ( .A(n20587), .B(n20586), .Z(n20766) );
  NANDN U21317 ( .A(n20589), .B(n20588), .Z(n20593) );
  NANDN U21318 ( .A(n20591), .B(n20590), .Z(n20592) );
  AND U21319 ( .A(n20593), .B(n20592), .Z(n20708) );
  NANDN U21320 ( .A(n20595), .B(n20594), .Z(n20599) );
  OR U21321 ( .A(n20597), .B(n20596), .Z(n20598) );
  NAND U21322 ( .A(n20599), .B(n20598), .Z(n20707) );
  XNOR U21323 ( .A(n20708), .B(n20707), .Z(n20710) );
  NAND U21324 ( .A(b[0]), .B(a[153]), .Z(n20600) );
  XNOR U21325 ( .A(b[1]), .B(n20600), .Z(n20602) );
  NANDN U21326 ( .A(b[0]), .B(a[152]), .Z(n20601) );
  NAND U21327 ( .A(n20602), .B(n20601), .Z(n20656) );
  NAND U21328 ( .A(n194), .B(n20603), .Z(n20605) );
  XOR U21329 ( .A(b[29]), .B(a[125]), .Z(n20732) );
  NAND U21330 ( .A(n38456), .B(n20732), .Z(n20604) );
  AND U21331 ( .A(n20605), .B(n20604), .Z(n20654) );
  AND U21332 ( .A(b[31]), .B(a[121]), .Z(n20653) );
  XNOR U21333 ( .A(n20654), .B(n20653), .Z(n20655) );
  XNOR U21334 ( .A(n20656), .B(n20655), .Z(n20696) );
  NAND U21335 ( .A(n38185), .B(n20606), .Z(n20608) );
  XOR U21336 ( .A(b[23]), .B(a[131]), .Z(n20735) );
  NAND U21337 ( .A(n38132), .B(n20735), .Z(n20607) );
  AND U21338 ( .A(n20608), .B(n20607), .Z(n20725) );
  NAND U21339 ( .A(n184), .B(n20609), .Z(n20611) );
  XOR U21340 ( .A(b[7]), .B(a[147]), .Z(n20738) );
  NAND U21341 ( .A(n36592), .B(n20738), .Z(n20610) );
  AND U21342 ( .A(n20611), .B(n20610), .Z(n20724) );
  NAND U21343 ( .A(n38289), .B(n20612), .Z(n20614) );
  XOR U21344 ( .A(b[25]), .B(a[129]), .Z(n20741) );
  NAND U21345 ( .A(n38247), .B(n20741), .Z(n20613) );
  NAND U21346 ( .A(n20614), .B(n20613), .Z(n20723) );
  XOR U21347 ( .A(n20724), .B(n20723), .Z(n20726) );
  XOR U21348 ( .A(n20725), .B(n20726), .Z(n20695) );
  XOR U21349 ( .A(n20696), .B(n20695), .Z(n20698) );
  NAND U21350 ( .A(n187), .B(n20615), .Z(n20617) );
  XOR U21351 ( .A(b[13]), .B(a[141]), .Z(n20744) );
  NAND U21352 ( .A(n37295), .B(n20744), .Z(n20616) );
  AND U21353 ( .A(n20617), .B(n20616), .Z(n20690) );
  NAND U21354 ( .A(n186), .B(n20618), .Z(n20620) );
  XOR U21355 ( .A(b[11]), .B(a[143]), .Z(n20747) );
  NAND U21356 ( .A(n37097), .B(n20747), .Z(n20619) );
  NAND U21357 ( .A(n20620), .B(n20619), .Z(n20689) );
  XNOR U21358 ( .A(n20690), .B(n20689), .Z(n20692) );
  NAND U21359 ( .A(n188), .B(n20621), .Z(n20623) );
  XOR U21360 ( .A(b[15]), .B(a[139]), .Z(n20750) );
  NAND U21361 ( .A(n37382), .B(n20750), .Z(n20622) );
  AND U21362 ( .A(n20623), .B(n20622), .Z(n20686) );
  NAND U21363 ( .A(n38064), .B(n20624), .Z(n20626) );
  XOR U21364 ( .A(b[21]), .B(a[133]), .Z(n20753) );
  NAND U21365 ( .A(n37993), .B(n20753), .Z(n20625) );
  AND U21366 ( .A(n20626), .B(n20625), .Z(n20684) );
  NAND U21367 ( .A(n185), .B(n20627), .Z(n20629) );
  XOR U21368 ( .A(b[9]), .B(a[145]), .Z(n20756) );
  NAND U21369 ( .A(n36805), .B(n20756), .Z(n20628) );
  NAND U21370 ( .A(n20629), .B(n20628), .Z(n20683) );
  XNOR U21371 ( .A(n20684), .B(n20683), .Z(n20685) );
  XNOR U21372 ( .A(n20686), .B(n20685), .Z(n20691) );
  XOR U21373 ( .A(n20692), .B(n20691), .Z(n20697) );
  XNOR U21374 ( .A(n20698), .B(n20697), .Z(n20709) );
  XNOR U21375 ( .A(n20710), .B(n20709), .Z(n20765) );
  XNOR U21376 ( .A(n20766), .B(n20765), .Z(n20767) );
  XOR U21377 ( .A(n20768), .B(n20767), .Z(n20772) );
  XNOR U21378 ( .A(n20771), .B(n20772), .Z(n20773) );
  XNOR U21379 ( .A(n20774), .B(n20773), .Z(n20779) );
  XOR U21380 ( .A(n20780), .B(n20779), .Z(n20648) );
  NANDN U21381 ( .A(n20631), .B(n20630), .Z(n20635) );
  NANDN U21382 ( .A(n20633), .B(n20632), .Z(n20634) );
  AND U21383 ( .A(n20635), .B(n20634), .Z(n20647) );
  XOR U21384 ( .A(n20648), .B(n20647), .Z(n20650) );
  XNOR U21385 ( .A(n20649), .B(n20650), .Z(n20641) );
  XNOR U21386 ( .A(n20642), .B(n20641), .Z(n20643) );
  XNOR U21387 ( .A(n20644), .B(n20643), .Z(n20783) );
  XNOR U21388 ( .A(sreg[377]), .B(n20783), .Z(n20785) );
  NANDN U21389 ( .A(sreg[376]), .B(n20636), .Z(n20640) );
  NAND U21390 ( .A(n20638), .B(n20637), .Z(n20639) );
  NAND U21391 ( .A(n20640), .B(n20639), .Z(n20784) );
  XNOR U21392 ( .A(n20785), .B(n20784), .Z(c[377]) );
  NANDN U21393 ( .A(n20642), .B(n20641), .Z(n20646) );
  NANDN U21394 ( .A(n20644), .B(n20643), .Z(n20645) );
  AND U21395 ( .A(n20646), .B(n20645), .Z(n20791) );
  NANDN U21396 ( .A(n20648), .B(n20647), .Z(n20652) );
  NANDN U21397 ( .A(n20650), .B(n20649), .Z(n20651) );
  AND U21398 ( .A(n20652), .B(n20651), .Z(n20789) );
  NANDN U21399 ( .A(n20654), .B(n20653), .Z(n20658) );
  NANDN U21400 ( .A(n20656), .B(n20655), .Z(n20657) );
  AND U21401 ( .A(n20658), .B(n20657), .Z(n20868) );
  NAND U21402 ( .A(n38385), .B(n20659), .Z(n20661) );
  XOR U21403 ( .A(b[27]), .B(a[128]), .Z(n20812) );
  NAND U21404 ( .A(n38343), .B(n20812), .Z(n20660) );
  AND U21405 ( .A(n20661), .B(n20660), .Z(n20875) );
  NAND U21406 ( .A(n183), .B(n20662), .Z(n20664) );
  XOR U21407 ( .A(b[5]), .B(a[150]), .Z(n20815) );
  NAND U21408 ( .A(n36296), .B(n20815), .Z(n20663) );
  AND U21409 ( .A(n20664), .B(n20663), .Z(n20873) );
  NAND U21410 ( .A(n190), .B(n20665), .Z(n20667) );
  XOR U21411 ( .A(b[19]), .B(a[136]), .Z(n20818) );
  NAND U21412 ( .A(n37821), .B(n20818), .Z(n20666) );
  NAND U21413 ( .A(n20667), .B(n20666), .Z(n20872) );
  XNOR U21414 ( .A(n20873), .B(n20872), .Z(n20874) );
  XNOR U21415 ( .A(n20875), .B(n20874), .Z(n20866) );
  NAND U21416 ( .A(n38470), .B(n20668), .Z(n20670) );
  XOR U21417 ( .A(b[31]), .B(a[124]), .Z(n20821) );
  NAND U21418 ( .A(n38453), .B(n20821), .Z(n20669) );
  AND U21419 ( .A(n20670), .B(n20669), .Z(n20833) );
  NAND U21420 ( .A(n181), .B(n20671), .Z(n20673) );
  XOR U21421 ( .A(b[3]), .B(a[152]), .Z(n20824) );
  NAND U21422 ( .A(n182), .B(n20824), .Z(n20672) );
  AND U21423 ( .A(n20673), .B(n20672), .Z(n20831) );
  NAND U21424 ( .A(n189), .B(n20674), .Z(n20676) );
  XOR U21425 ( .A(b[17]), .B(a[138]), .Z(n20827) );
  NAND U21426 ( .A(n37652), .B(n20827), .Z(n20675) );
  NAND U21427 ( .A(n20676), .B(n20675), .Z(n20830) );
  XNOR U21428 ( .A(n20831), .B(n20830), .Z(n20832) );
  XOR U21429 ( .A(n20833), .B(n20832), .Z(n20867) );
  XOR U21430 ( .A(n20866), .B(n20867), .Z(n20869) );
  XOR U21431 ( .A(n20868), .B(n20869), .Z(n20915) );
  NANDN U21432 ( .A(n20678), .B(n20677), .Z(n20682) );
  NANDN U21433 ( .A(n20680), .B(n20679), .Z(n20681) );
  AND U21434 ( .A(n20682), .B(n20681), .Z(n20854) );
  NANDN U21435 ( .A(n20684), .B(n20683), .Z(n20688) );
  NANDN U21436 ( .A(n20686), .B(n20685), .Z(n20687) );
  NAND U21437 ( .A(n20688), .B(n20687), .Z(n20855) );
  XNOR U21438 ( .A(n20854), .B(n20855), .Z(n20856) );
  NANDN U21439 ( .A(n20690), .B(n20689), .Z(n20694) );
  NAND U21440 ( .A(n20692), .B(n20691), .Z(n20693) );
  NAND U21441 ( .A(n20694), .B(n20693), .Z(n20857) );
  XNOR U21442 ( .A(n20856), .B(n20857), .Z(n20914) );
  XNOR U21443 ( .A(n20915), .B(n20914), .Z(n20917) );
  NAND U21444 ( .A(n20696), .B(n20695), .Z(n20700) );
  NAND U21445 ( .A(n20698), .B(n20697), .Z(n20699) );
  AND U21446 ( .A(n20700), .B(n20699), .Z(n20916) );
  XOR U21447 ( .A(n20917), .B(n20916), .Z(n20928) );
  NANDN U21448 ( .A(n20702), .B(n20701), .Z(n20706) );
  NANDN U21449 ( .A(n20704), .B(n20703), .Z(n20705) );
  AND U21450 ( .A(n20706), .B(n20705), .Z(n20926) );
  NANDN U21451 ( .A(n20712), .B(n20711), .Z(n20716) );
  OR U21452 ( .A(n20714), .B(n20713), .Z(n20715) );
  AND U21453 ( .A(n20716), .B(n20715), .Z(n20921) );
  NANDN U21454 ( .A(n20718), .B(n20717), .Z(n20722) );
  NANDN U21455 ( .A(n20720), .B(n20719), .Z(n20721) );
  AND U21456 ( .A(n20722), .B(n20721), .Z(n20861) );
  NANDN U21457 ( .A(n20724), .B(n20723), .Z(n20728) );
  OR U21458 ( .A(n20726), .B(n20725), .Z(n20727) );
  NAND U21459 ( .A(n20728), .B(n20727), .Z(n20860) );
  XNOR U21460 ( .A(n20861), .B(n20860), .Z(n20862) );
  NAND U21461 ( .A(b[0]), .B(a[154]), .Z(n20729) );
  XNOR U21462 ( .A(b[1]), .B(n20729), .Z(n20731) );
  NANDN U21463 ( .A(b[0]), .B(a[153]), .Z(n20730) );
  NAND U21464 ( .A(n20731), .B(n20730), .Z(n20809) );
  NAND U21465 ( .A(n194), .B(n20732), .Z(n20734) );
  XOR U21466 ( .A(b[29]), .B(a[126]), .Z(n20887) );
  NAND U21467 ( .A(n38456), .B(n20887), .Z(n20733) );
  AND U21468 ( .A(n20734), .B(n20733), .Z(n20807) );
  AND U21469 ( .A(b[31]), .B(a[122]), .Z(n20806) );
  XNOR U21470 ( .A(n20807), .B(n20806), .Z(n20808) );
  XNOR U21471 ( .A(n20809), .B(n20808), .Z(n20848) );
  NAND U21472 ( .A(n38185), .B(n20735), .Z(n20737) );
  XOR U21473 ( .A(b[23]), .B(a[132]), .Z(n20890) );
  NAND U21474 ( .A(n38132), .B(n20890), .Z(n20736) );
  AND U21475 ( .A(n20737), .B(n20736), .Z(n20881) );
  NAND U21476 ( .A(n184), .B(n20738), .Z(n20740) );
  XOR U21477 ( .A(b[7]), .B(a[148]), .Z(n20893) );
  NAND U21478 ( .A(n36592), .B(n20893), .Z(n20739) );
  AND U21479 ( .A(n20740), .B(n20739), .Z(n20879) );
  NAND U21480 ( .A(n38289), .B(n20741), .Z(n20743) );
  XOR U21481 ( .A(b[25]), .B(a[130]), .Z(n20896) );
  NAND U21482 ( .A(n38247), .B(n20896), .Z(n20742) );
  NAND U21483 ( .A(n20743), .B(n20742), .Z(n20878) );
  XNOR U21484 ( .A(n20879), .B(n20878), .Z(n20880) );
  XOR U21485 ( .A(n20881), .B(n20880), .Z(n20849) );
  XNOR U21486 ( .A(n20848), .B(n20849), .Z(n20850) );
  NAND U21487 ( .A(n187), .B(n20744), .Z(n20746) );
  XOR U21488 ( .A(b[13]), .B(a[142]), .Z(n20899) );
  NAND U21489 ( .A(n37295), .B(n20899), .Z(n20745) );
  AND U21490 ( .A(n20746), .B(n20745), .Z(n20843) );
  NAND U21491 ( .A(n186), .B(n20747), .Z(n20749) );
  XOR U21492 ( .A(b[11]), .B(a[144]), .Z(n20902) );
  NAND U21493 ( .A(n37097), .B(n20902), .Z(n20748) );
  NAND U21494 ( .A(n20749), .B(n20748), .Z(n20842) );
  XNOR U21495 ( .A(n20843), .B(n20842), .Z(n20844) );
  NAND U21496 ( .A(n188), .B(n20750), .Z(n20752) );
  XOR U21497 ( .A(b[15]), .B(a[140]), .Z(n20905) );
  NAND U21498 ( .A(n37382), .B(n20905), .Z(n20751) );
  AND U21499 ( .A(n20752), .B(n20751), .Z(n20839) );
  NAND U21500 ( .A(n38064), .B(n20753), .Z(n20755) );
  XOR U21501 ( .A(b[21]), .B(a[134]), .Z(n20908) );
  NAND U21502 ( .A(n37993), .B(n20908), .Z(n20754) );
  AND U21503 ( .A(n20755), .B(n20754), .Z(n20837) );
  NAND U21504 ( .A(n185), .B(n20756), .Z(n20758) );
  XOR U21505 ( .A(b[9]), .B(a[146]), .Z(n20911) );
  NAND U21506 ( .A(n36805), .B(n20911), .Z(n20757) );
  NAND U21507 ( .A(n20758), .B(n20757), .Z(n20836) );
  XNOR U21508 ( .A(n20837), .B(n20836), .Z(n20838) );
  XOR U21509 ( .A(n20839), .B(n20838), .Z(n20845) );
  XOR U21510 ( .A(n20844), .B(n20845), .Z(n20851) );
  XOR U21511 ( .A(n20850), .B(n20851), .Z(n20863) );
  XNOR U21512 ( .A(n20862), .B(n20863), .Z(n20920) );
  XNOR U21513 ( .A(n20921), .B(n20920), .Z(n20922) );
  XOR U21514 ( .A(n20923), .B(n20922), .Z(n20927) );
  XOR U21515 ( .A(n20926), .B(n20927), .Z(n20929) );
  XOR U21516 ( .A(n20928), .B(n20929), .Z(n20803) );
  NANDN U21517 ( .A(n20760), .B(n20759), .Z(n20764) );
  NAND U21518 ( .A(n20762), .B(n20761), .Z(n20763) );
  AND U21519 ( .A(n20764), .B(n20763), .Z(n20801) );
  NANDN U21520 ( .A(n20766), .B(n20765), .Z(n20770) );
  NANDN U21521 ( .A(n20768), .B(n20767), .Z(n20769) );
  AND U21522 ( .A(n20770), .B(n20769), .Z(n20800) );
  XNOR U21523 ( .A(n20801), .B(n20800), .Z(n20802) );
  XNOR U21524 ( .A(n20803), .B(n20802), .Z(n20794) );
  NANDN U21525 ( .A(n20772), .B(n20771), .Z(n20776) );
  NANDN U21526 ( .A(n20774), .B(n20773), .Z(n20775) );
  NAND U21527 ( .A(n20776), .B(n20775), .Z(n20795) );
  XNOR U21528 ( .A(n20794), .B(n20795), .Z(n20796) );
  NANDN U21529 ( .A(n20778), .B(n20777), .Z(n20782) );
  NAND U21530 ( .A(n20780), .B(n20779), .Z(n20781) );
  NAND U21531 ( .A(n20782), .B(n20781), .Z(n20797) );
  XNOR U21532 ( .A(n20796), .B(n20797), .Z(n20788) );
  XNOR U21533 ( .A(n20789), .B(n20788), .Z(n20790) );
  XNOR U21534 ( .A(n20791), .B(n20790), .Z(n20932) );
  XNOR U21535 ( .A(sreg[378]), .B(n20932), .Z(n20934) );
  NANDN U21536 ( .A(sreg[377]), .B(n20783), .Z(n20787) );
  NAND U21537 ( .A(n20785), .B(n20784), .Z(n20786) );
  NAND U21538 ( .A(n20787), .B(n20786), .Z(n20933) );
  XNOR U21539 ( .A(n20934), .B(n20933), .Z(c[378]) );
  NANDN U21540 ( .A(n20789), .B(n20788), .Z(n20793) );
  NANDN U21541 ( .A(n20791), .B(n20790), .Z(n20792) );
  AND U21542 ( .A(n20793), .B(n20792), .Z(n20940) );
  NANDN U21543 ( .A(n20795), .B(n20794), .Z(n20799) );
  NANDN U21544 ( .A(n20797), .B(n20796), .Z(n20798) );
  AND U21545 ( .A(n20799), .B(n20798), .Z(n20938) );
  NANDN U21546 ( .A(n20801), .B(n20800), .Z(n20805) );
  NANDN U21547 ( .A(n20803), .B(n20802), .Z(n20804) );
  AND U21548 ( .A(n20805), .B(n20804), .Z(n20946) );
  NANDN U21549 ( .A(n20807), .B(n20806), .Z(n20811) );
  NANDN U21550 ( .A(n20809), .B(n20808), .Z(n20810) );
  AND U21551 ( .A(n20811), .B(n20810), .Z(n21027) );
  NAND U21552 ( .A(n38385), .B(n20812), .Z(n20814) );
  XOR U21553 ( .A(b[27]), .B(a[129]), .Z(n20973) );
  NAND U21554 ( .A(n38343), .B(n20973), .Z(n20813) );
  AND U21555 ( .A(n20814), .B(n20813), .Z(n21034) );
  NAND U21556 ( .A(n183), .B(n20815), .Z(n20817) );
  XOR U21557 ( .A(b[5]), .B(a[151]), .Z(n20976) );
  NAND U21558 ( .A(n36296), .B(n20976), .Z(n20816) );
  AND U21559 ( .A(n20817), .B(n20816), .Z(n21032) );
  NAND U21560 ( .A(n190), .B(n20818), .Z(n20820) );
  XOR U21561 ( .A(b[19]), .B(a[137]), .Z(n20979) );
  NAND U21562 ( .A(n37821), .B(n20979), .Z(n20819) );
  NAND U21563 ( .A(n20820), .B(n20819), .Z(n21031) );
  XNOR U21564 ( .A(n21032), .B(n21031), .Z(n21033) );
  XNOR U21565 ( .A(n21034), .B(n21033), .Z(n21025) );
  NAND U21566 ( .A(n38470), .B(n20821), .Z(n20823) );
  XOR U21567 ( .A(b[31]), .B(a[125]), .Z(n20982) );
  NAND U21568 ( .A(n38453), .B(n20982), .Z(n20822) );
  AND U21569 ( .A(n20823), .B(n20822), .Z(n20994) );
  NAND U21570 ( .A(n181), .B(n20824), .Z(n20826) );
  XOR U21571 ( .A(b[3]), .B(a[153]), .Z(n20985) );
  NAND U21572 ( .A(n182), .B(n20985), .Z(n20825) );
  AND U21573 ( .A(n20826), .B(n20825), .Z(n20992) );
  NAND U21574 ( .A(n189), .B(n20827), .Z(n20829) );
  XOR U21575 ( .A(b[17]), .B(a[139]), .Z(n20988) );
  NAND U21576 ( .A(n37652), .B(n20988), .Z(n20828) );
  NAND U21577 ( .A(n20829), .B(n20828), .Z(n20991) );
  XNOR U21578 ( .A(n20992), .B(n20991), .Z(n20993) );
  XOR U21579 ( .A(n20994), .B(n20993), .Z(n21026) );
  XOR U21580 ( .A(n21025), .B(n21026), .Z(n21028) );
  XOR U21581 ( .A(n21027), .B(n21028), .Z(n20962) );
  NANDN U21582 ( .A(n20831), .B(n20830), .Z(n20835) );
  NANDN U21583 ( .A(n20833), .B(n20832), .Z(n20834) );
  AND U21584 ( .A(n20835), .B(n20834), .Z(n21015) );
  NANDN U21585 ( .A(n20837), .B(n20836), .Z(n20841) );
  NANDN U21586 ( .A(n20839), .B(n20838), .Z(n20840) );
  NAND U21587 ( .A(n20841), .B(n20840), .Z(n21016) );
  XNOR U21588 ( .A(n21015), .B(n21016), .Z(n21017) );
  NANDN U21589 ( .A(n20843), .B(n20842), .Z(n20847) );
  NANDN U21590 ( .A(n20845), .B(n20844), .Z(n20846) );
  NAND U21591 ( .A(n20847), .B(n20846), .Z(n21018) );
  XNOR U21592 ( .A(n21017), .B(n21018), .Z(n20961) );
  XNOR U21593 ( .A(n20962), .B(n20961), .Z(n20964) );
  NANDN U21594 ( .A(n20849), .B(n20848), .Z(n20853) );
  NANDN U21595 ( .A(n20851), .B(n20850), .Z(n20852) );
  AND U21596 ( .A(n20853), .B(n20852), .Z(n20963) );
  XOR U21597 ( .A(n20964), .B(n20963), .Z(n21075) );
  NANDN U21598 ( .A(n20855), .B(n20854), .Z(n20859) );
  NANDN U21599 ( .A(n20857), .B(n20856), .Z(n20858) );
  AND U21600 ( .A(n20859), .B(n20858), .Z(n21073) );
  NANDN U21601 ( .A(n20861), .B(n20860), .Z(n20865) );
  NANDN U21602 ( .A(n20863), .B(n20862), .Z(n20864) );
  AND U21603 ( .A(n20865), .B(n20864), .Z(n20958) );
  NANDN U21604 ( .A(n20867), .B(n20866), .Z(n20871) );
  OR U21605 ( .A(n20869), .B(n20868), .Z(n20870) );
  AND U21606 ( .A(n20871), .B(n20870), .Z(n20956) );
  NANDN U21607 ( .A(n20873), .B(n20872), .Z(n20877) );
  NANDN U21608 ( .A(n20875), .B(n20874), .Z(n20876) );
  AND U21609 ( .A(n20877), .B(n20876), .Z(n21022) );
  NANDN U21610 ( .A(n20879), .B(n20878), .Z(n20883) );
  NANDN U21611 ( .A(n20881), .B(n20880), .Z(n20882) );
  NAND U21612 ( .A(n20883), .B(n20882), .Z(n21021) );
  XNOR U21613 ( .A(n21022), .B(n21021), .Z(n21024) );
  NAND U21614 ( .A(b[0]), .B(a[155]), .Z(n20884) );
  XNOR U21615 ( .A(b[1]), .B(n20884), .Z(n20886) );
  NANDN U21616 ( .A(b[0]), .B(a[154]), .Z(n20885) );
  NAND U21617 ( .A(n20886), .B(n20885), .Z(n20970) );
  NAND U21618 ( .A(n194), .B(n20887), .Z(n20889) );
  XOR U21619 ( .A(b[29]), .B(a[127]), .Z(n21046) );
  NAND U21620 ( .A(n38456), .B(n21046), .Z(n20888) );
  AND U21621 ( .A(n20889), .B(n20888), .Z(n20968) );
  AND U21622 ( .A(b[31]), .B(a[123]), .Z(n20967) );
  XNOR U21623 ( .A(n20968), .B(n20967), .Z(n20969) );
  XNOR U21624 ( .A(n20970), .B(n20969), .Z(n21010) );
  NAND U21625 ( .A(n38185), .B(n20890), .Z(n20892) );
  XOR U21626 ( .A(b[23]), .B(a[133]), .Z(n21049) );
  NAND U21627 ( .A(n38132), .B(n21049), .Z(n20891) );
  AND U21628 ( .A(n20892), .B(n20891), .Z(n21039) );
  NAND U21629 ( .A(n184), .B(n20893), .Z(n20895) );
  XOR U21630 ( .A(b[7]), .B(a[149]), .Z(n21052) );
  NAND U21631 ( .A(n36592), .B(n21052), .Z(n20894) );
  AND U21632 ( .A(n20895), .B(n20894), .Z(n21038) );
  NAND U21633 ( .A(n38289), .B(n20896), .Z(n20898) );
  XOR U21634 ( .A(b[25]), .B(a[131]), .Z(n21055) );
  NAND U21635 ( .A(n38247), .B(n21055), .Z(n20897) );
  NAND U21636 ( .A(n20898), .B(n20897), .Z(n21037) );
  XOR U21637 ( .A(n21038), .B(n21037), .Z(n21040) );
  XOR U21638 ( .A(n21039), .B(n21040), .Z(n21009) );
  XOR U21639 ( .A(n21010), .B(n21009), .Z(n21012) );
  NAND U21640 ( .A(n187), .B(n20899), .Z(n20901) );
  XOR U21641 ( .A(b[13]), .B(a[143]), .Z(n21058) );
  NAND U21642 ( .A(n37295), .B(n21058), .Z(n20900) );
  AND U21643 ( .A(n20901), .B(n20900), .Z(n21004) );
  NAND U21644 ( .A(n186), .B(n20902), .Z(n20904) );
  XOR U21645 ( .A(b[11]), .B(a[145]), .Z(n21061) );
  NAND U21646 ( .A(n37097), .B(n21061), .Z(n20903) );
  NAND U21647 ( .A(n20904), .B(n20903), .Z(n21003) );
  XNOR U21648 ( .A(n21004), .B(n21003), .Z(n21006) );
  NAND U21649 ( .A(n188), .B(n20905), .Z(n20907) );
  XOR U21650 ( .A(b[15]), .B(a[141]), .Z(n21064) );
  NAND U21651 ( .A(n37382), .B(n21064), .Z(n20906) );
  AND U21652 ( .A(n20907), .B(n20906), .Z(n21000) );
  NAND U21653 ( .A(n38064), .B(n20908), .Z(n20910) );
  XOR U21654 ( .A(b[21]), .B(a[135]), .Z(n21067) );
  NAND U21655 ( .A(n37993), .B(n21067), .Z(n20909) );
  AND U21656 ( .A(n20910), .B(n20909), .Z(n20998) );
  NAND U21657 ( .A(n185), .B(n20911), .Z(n20913) );
  XOR U21658 ( .A(b[9]), .B(a[147]), .Z(n21070) );
  NAND U21659 ( .A(n36805), .B(n21070), .Z(n20912) );
  NAND U21660 ( .A(n20913), .B(n20912), .Z(n20997) );
  XNOR U21661 ( .A(n20998), .B(n20997), .Z(n20999) );
  XNOR U21662 ( .A(n21000), .B(n20999), .Z(n21005) );
  XOR U21663 ( .A(n21006), .B(n21005), .Z(n21011) );
  XNOR U21664 ( .A(n21012), .B(n21011), .Z(n21023) );
  XNOR U21665 ( .A(n21024), .B(n21023), .Z(n20955) );
  XNOR U21666 ( .A(n20956), .B(n20955), .Z(n20957) );
  XOR U21667 ( .A(n20958), .B(n20957), .Z(n21074) );
  XOR U21668 ( .A(n21073), .B(n21074), .Z(n21076) );
  XOR U21669 ( .A(n21075), .B(n21076), .Z(n20952) );
  NANDN U21670 ( .A(n20915), .B(n20914), .Z(n20919) );
  NAND U21671 ( .A(n20917), .B(n20916), .Z(n20918) );
  AND U21672 ( .A(n20919), .B(n20918), .Z(n20950) );
  NANDN U21673 ( .A(n20921), .B(n20920), .Z(n20925) );
  NANDN U21674 ( .A(n20923), .B(n20922), .Z(n20924) );
  AND U21675 ( .A(n20925), .B(n20924), .Z(n20949) );
  XNOR U21676 ( .A(n20950), .B(n20949), .Z(n20951) );
  XNOR U21677 ( .A(n20952), .B(n20951), .Z(n20943) );
  NANDN U21678 ( .A(n20927), .B(n20926), .Z(n20931) );
  OR U21679 ( .A(n20929), .B(n20928), .Z(n20930) );
  NAND U21680 ( .A(n20931), .B(n20930), .Z(n20944) );
  XNOR U21681 ( .A(n20943), .B(n20944), .Z(n20945) );
  XNOR U21682 ( .A(n20946), .B(n20945), .Z(n20937) );
  XNOR U21683 ( .A(n20938), .B(n20937), .Z(n20939) );
  XNOR U21684 ( .A(n20940), .B(n20939), .Z(n21079) );
  XNOR U21685 ( .A(sreg[379]), .B(n21079), .Z(n21081) );
  NANDN U21686 ( .A(sreg[378]), .B(n20932), .Z(n20936) );
  NAND U21687 ( .A(n20934), .B(n20933), .Z(n20935) );
  NAND U21688 ( .A(n20936), .B(n20935), .Z(n21080) );
  XNOR U21689 ( .A(n21081), .B(n21080), .Z(c[379]) );
  NANDN U21690 ( .A(n20938), .B(n20937), .Z(n20942) );
  NANDN U21691 ( .A(n20940), .B(n20939), .Z(n20941) );
  AND U21692 ( .A(n20942), .B(n20941), .Z(n21087) );
  NANDN U21693 ( .A(n20944), .B(n20943), .Z(n20948) );
  NANDN U21694 ( .A(n20946), .B(n20945), .Z(n20947) );
  AND U21695 ( .A(n20948), .B(n20947), .Z(n21085) );
  NANDN U21696 ( .A(n20950), .B(n20949), .Z(n20954) );
  NANDN U21697 ( .A(n20952), .B(n20951), .Z(n20953) );
  AND U21698 ( .A(n20954), .B(n20953), .Z(n21093) );
  NANDN U21699 ( .A(n20956), .B(n20955), .Z(n20960) );
  NANDN U21700 ( .A(n20958), .B(n20957), .Z(n20959) );
  AND U21701 ( .A(n20960), .B(n20959), .Z(n21223) );
  NANDN U21702 ( .A(n20962), .B(n20961), .Z(n20966) );
  NAND U21703 ( .A(n20964), .B(n20963), .Z(n20965) );
  AND U21704 ( .A(n20966), .B(n20965), .Z(n21222) );
  XNOR U21705 ( .A(n21223), .B(n21222), .Z(n21225) );
  NANDN U21706 ( .A(n20968), .B(n20967), .Z(n20972) );
  NANDN U21707 ( .A(n20970), .B(n20969), .Z(n20971) );
  AND U21708 ( .A(n20972), .B(n20971), .Z(n21158) );
  NAND U21709 ( .A(n38385), .B(n20973), .Z(n20975) );
  XOR U21710 ( .A(b[27]), .B(a[130]), .Z(n21102) );
  NAND U21711 ( .A(n38343), .B(n21102), .Z(n20974) );
  AND U21712 ( .A(n20975), .B(n20974), .Z(n21165) );
  NAND U21713 ( .A(n183), .B(n20976), .Z(n20978) );
  XOR U21714 ( .A(b[5]), .B(a[152]), .Z(n21105) );
  NAND U21715 ( .A(n36296), .B(n21105), .Z(n20977) );
  AND U21716 ( .A(n20978), .B(n20977), .Z(n21163) );
  NAND U21717 ( .A(n190), .B(n20979), .Z(n20981) );
  XOR U21718 ( .A(b[19]), .B(a[138]), .Z(n21108) );
  NAND U21719 ( .A(n37821), .B(n21108), .Z(n20980) );
  NAND U21720 ( .A(n20981), .B(n20980), .Z(n21162) );
  XNOR U21721 ( .A(n21163), .B(n21162), .Z(n21164) );
  XNOR U21722 ( .A(n21165), .B(n21164), .Z(n21156) );
  NAND U21723 ( .A(n38470), .B(n20982), .Z(n20984) );
  XOR U21724 ( .A(b[31]), .B(a[126]), .Z(n21111) );
  NAND U21725 ( .A(n38453), .B(n21111), .Z(n20983) );
  AND U21726 ( .A(n20984), .B(n20983), .Z(n21123) );
  NAND U21727 ( .A(n181), .B(n20985), .Z(n20987) );
  XOR U21728 ( .A(b[3]), .B(a[154]), .Z(n21114) );
  NAND U21729 ( .A(n182), .B(n21114), .Z(n20986) );
  AND U21730 ( .A(n20987), .B(n20986), .Z(n21121) );
  NAND U21731 ( .A(n189), .B(n20988), .Z(n20990) );
  XOR U21732 ( .A(b[17]), .B(a[140]), .Z(n21117) );
  NAND U21733 ( .A(n37652), .B(n21117), .Z(n20989) );
  NAND U21734 ( .A(n20990), .B(n20989), .Z(n21120) );
  XNOR U21735 ( .A(n21121), .B(n21120), .Z(n21122) );
  XOR U21736 ( .A(n21123), .B(n21122), .Z(n21157) );
  XOR U21737 ( .A(n21156), .B(n21157), .Z(n21159) );
  XOR U21738 ( .A(n21158), .B(n21159), .Z(n21205) );
  NANDN U21739 ( .A(n20992), .B(n20991), .Z(n20996) );
  NANDN U21740 ( .A(n20994), .B(n20993), .Z(n20995) );
  AND U21741 ( .A(n20996), .B(n20995), .Z(n21144) );
  NANDN U21742 ( .A(n20998), .B(n20997), .Z(n21002) );
  NANDN U21743 ( .A(n21000), .B(n20999), .Z(n21001) );
  NAND U21744 ( .A(n21002), .B(n21001), .Z(n21145) );
  XNOR U21745 ( .A(n21144), .B(n21145), .Z(n21146) );
  NANDN U21746 ( .A(n21004), .B(n21003), .Z(n21008) );
  NAND U21747 ( .A(n21006), .B(n21005), .Z(n21007) );
  NAND U21748 ( .A(n21008), .B(n21007), .Z(n21147) );
  XNOR U21749 ( .A(n21146), .B(n21147), .Z(n21204) );
  XNOR U21750 ( .A(n21205), .B(n21204), .Z(n21207) );
  NAND U21751 ( .A(n21010), .B(n21009), .Z(n21014) );
  NAND U21752 ( .A(n21012), .B(n21011), .Z(n21013) );
  AND U21753 ( .A(n21014), .B(n21013), .Z(n21206) );
  XOR U21754 ( .A(n21207), .B(n21206), .Z(n21219) );
  NANDN U21755 ( .A(n21016), .B(n21015), .Z(n21020) );
  NANDN U21756 ( .A(n21018), .B(n21017), .Z(n21019) );
  AND U21757 ( .A(n21020), .B(n21019), .Z(n21216) );
  NANDN U21758 ( .A(n21026), .B(n21025), .Z(n21030) );
  OR U21759 ( .A(n21028), .B(n21027), .Z(n21029) );
  AND U21760 ( .A(n21030), .B(n21029), .Z(n21211) );
  NANDN U21761 ( .A(n21032), .B(n21031), .Z(n21036) );
  NANDN U21762 ( .A(n21034), .B(n21033), .Z(n21035) );
  AND U21763 ( .A(n21036), .B(n21035), .Z(n21151) );
  NANDN U21764 ( .A(n21038), .B(n21037), .Z(n21042) );
  OR U21765 ( .A(n21040), .B(n21039), .Z(n21041) );
  NAND U21766 ( .A(n21042), .B(n21041), .Z(n21150) );
  XNOR U21767 ( .A(n21151), .B(n21150), .Z(n21152) );
  NAND U21768 ( .A(b[0]), .B(a[156]), .Z(n21043) );
  XNOR U21769 ( .A(b[1]), .B(n21043), .Z(n21045) );
  NANDN U21770 ( .A(b[0]), .B(a[155]), .Z(n21044) );
  NAND U21771 ( .A(n21045), .B(n21044), .Z(n21099) );
  NAND U21772 ( .A(n194), .B(n21046), .Z(n21048) );
  XOR U21773 ( .A(b[29]), .B(a[128]), .Z(n21177) );
  NAND U21774 ( .A(n38456), .B(n21177), .Z(n21047) );
  AND U21775 ( .A(n21048), .B(n21047), .Z(n21097) );
  AND U21776 ( .A(b[31]), .B(a[124]), .Z(n21096) );
  XNOR U21777 ( .A(n21097), .B(n21096), .Z(n21098) );
  XNOR U21778 ( .A(n21099), .B(n21098), .Z(n21138) );
  NAND U21779 ( .A(n38185), .B(n21049), .Z(n21051) );
  XOR U21780 ( .A(b[23]), .B(a[134]), .Z(n21180) );
  NAND U21781 ( .A(n38132), .B(n21180), .Z(n21050) );
  AND U21782 ( .A(n21051), .B(n21050), .Z(n21171) );
  NAND U21783 ( .A(n184), .B(n21052), .Z(n21054) );
  XOR U21784 ( .A(b[7]), .B(a[150]), .Z(n21183) );
  NAND U21785 ( .A(n36592), .B(n21183), .Z(n21053) );
  AND U21786 ( .A(n21054), .B(n21053), .Z(n21169) );
  NAND U21787 ( .A(n38289), .B(n21055), .Z(n21057) );
  XOR U21788 ( .A(b[25]), .B(a[132]), .Z(n21186) );
  NAND U21789 ( .A(n38247), .B(n21186), .Z(n21056) );
  NAND U21790 ( .A(n21057), .B(n21056), .Z(n21168) );
  XNOR U21791 ( .A(n21169), .B(n21168), .Z(n21170) );
  XOR U21792 ( .A(n21171), .B(n21170), .Z(n21139) );
  XNOR U21793 ( .A(n21138), .B(n21139), .Z(n21140) );
  NAND U21794 ( .A(n187), .B(n21058), .Z(n21060) );
  XOR U21795 ( .A(b[13]), .B(a[144]), .Z(n21189) );
  NAND U21796 ( .A(n37295), .B(n21189), .Z(n21059) );
  AND U21797 ( .A(n21060), .B(n21059), .Z(n21133) );
  NAND U21798 ( .A(n186), .B(n21061), .Z(n21063) );
  XOR U21799 ( .A(b[11]), .B(a[146]), .Z(n21192) );
  NAND U21800 ( .A(n37097), .B(n21192), .Z(n21062) );
  NAND U21801 ( .A(n21063), .B(n21062), .Z(n21132) );
  XNOR U21802 ( .A(n21133), .B(n21132), .Z(n21134) );
  NAND U21803 ( .A(n188), .B(n21064), .Z(n21066) );
  XOR U21804 ( .A(b[15]), .B(a[142]), .Z(n21195) );
  NAND U21805 ( .A(n37382), .B(n21195), .Z(n21065) );
  AND U21806 ( .A(n21066), .B(n21065), .Z(n21129) );
  NAND U21807 ( .A(n38064), .B(n21067), .Z(n21069) );
  XOR U21808 ( .A(b[21]), .B(a[136]), .Z(n21198) );
  NAND U21809 ( .A(n37993), .B(n21198), .Z(n21068) );
  AND U21810 ( .A(n21069), .B(n21068), .Z(n21127) );
  NAND U21811 ( .A(n185), .B(n21070), .Z(n21072) );
  XOR U21812 ( .A(b[9]), .B(a[148]), .Z(n21201) );
  NAND U21813 ( .A(n36805), .B(n21201), .Z(n21071) );
  NAND U21814 ( .A(n21072), .B(n21071), .Z(n21126) );
  XNOR U21815 ( .A(n21127), .B(n21126), .Z(n21128) );
  XOR U21816 ( .A(n21129), .B(n21128), .Z(n21135) );
  XOR U21817 ( .A(n21134), .B(n21135), .Z(n21141) );
  XOR U21818 ( .A(n21140), .B(n21141), .Z(n21153) );
  XNOR U21819 ( .A(n21152), .B(n21153), .Z(n21210) );
  XNOR U21820 ( .A(n21211), .B(n21210), .Z(n21212) );
  XOR U21821 ( .A(n21213), .B(n21212), .Z(n21217) );
  XNOR U21822 ( .A(n21216), .B(n21217), .Z(n21218) );
  XNOR U21823 ( .A(n21219), .B(n21218), .Z(n21224) );
  XOR U21824 ( .A(n21225), .B(n21224), .Z(n21091) );
  NANDN U21825 ( .A(n21074), .B(n21073), .Z(n21078) );
  OR U21826 ( .A(n21076), .B(n21075), .Z(n21077) );
  AND U21827 ( .A(n21078), .B(n21077), .Z(n21090) );
  XNOR U21828 ( .A(n21091), .B(n21090), .Z(n21092) );
  XNOR U21829 ( .A(n21093), .B(n21092), .Z(n21084) );
  XNOR U21830 ( .A(n21085), .B(n21084), .Z(n21086) );
  XNOR U21831 ( .A(n21087), .B(n21086), .Z(n21228) );
  XNOR U21832 ( .A(sreg[380]), .B(n21228), .Z(n21230) );
  NANDN U21833 ( .A(sreg[379]), .B(n21079), .Z(n21083) );
  NAND U21834 ( .A(n21081), .B(n21080), .Z(n21082) );
  NAND U21835 ( .A(n21083), .B(n21082), .Z(n21229) );
  XNOR U21836 ( .A(n21230), .B(n21229), .Z(c[380]) );
  NANDN U21837 ( .A(n21085), .B(n21084), .Z(n21089) );
  NANDN U21838 ( .A(n21087), .B(n21086), .Z(n21088) );
  AND U21839 ( .A(n21089), .B(n21088), .Z(n21236) );
  NANDN U21840 ( .A(n21091), .B(n21090), .Z(n21095) );
  NANDN U21841 ( .A(n21093), .B(n21092), .Z(n21094) );
  AND U21842 ( .A(n21095), .B(n21094), .Z(n21234) );
  NANDN U21843 ( .A(n21097), .B(n21096), .Z(n21101) );
  NANDN U21844 ( .A(n21099), .B(n21098), .Z(n21100) );
  AND U21845 ( .A(n21101), .B(n21100), .Z(n21325) );
  NAND U21846 ( .A(n38385), .B(n21102), .Z(n21104) );
  XOR U21847 ( .A(b[27]), .B(a[131]), .Z(n21269) );
  NAND U21848 ( .A(n38343), .B(n21269), .Z(n21103) );
  AND U21849 ( .A(n21104), .B(n21103), .Z(n21332) );
  NAND U21850 ( .A(n183), .B(n21105), .Z(n21107) );
  XOR U21851 ( .A(b[5]), .B(a[153]), .Z(n21272) );
  NAND U21852 ( .A(n36296), .B(n21272), .Z(n21106) );
  AND U21853 ( .A(n21107), .B(n21106), .Z(n21330) );
  NAND U21854 ( .A(n190), .B(n21108), .Z(n21110) );
  XOR U21855 ( .A(b[19]), .B(a[139]), .Z(n21275) );
  NAND U21856 ( .A(n37821), .B(n21275), .Z(n21109) );
  NAND U21857 ( .A(n21110), .B(n21109), .Z(n21329) );
  XNOR U21858 ( .A(n21330), .B(n21329), .Z(n21331) );
  XNOR U21859 ( .A(n21332), .B(n21331), .Z(n21323) );
  NAND U21860 ( .A(n38470), .B(n21111), .Z(n21113) );
  XOR U21861 ( .A(b[31]), .B(a[127]), .Z(n21278) );
  NAND U21862 ( .A(n38453), .B(n21278), .Z(n21112) );
  AND U21863 ( .A(n21113), .B(n21112), .Z(n21290) );
  NAND U21864 ( .A(n181), .B(n21114), .Z(n21116) );
  XOR U21865 ( .A(b[3]), .B(a[155]), .Z(n21281) );
  NAND U21866 ( .A(n182), .B(n21281), .Z(n21115) );
  AND U21867 ( .A(n21116), .B(n21115), .Z(n21288) );
  NAND U21868 ( .A(n189), .B(n21117), .Z(n21119) );
  XOR U21869 ( .A(b[17]), .B(a[141]), .Z(n21284) );
  NAND U21870 ( .A(n37652), .B(n21284), .Z(n21118) );
  NAND U21871 ( .A(n21119), .B(n21118), .Z(n21287) );
  XNOR U21872 ( .A(n21288), .B(n21287), .Z(n21289) );
  XOR U21873 ( .A(n21290), .B(n21289), .Z(n21324) );
  XOR U21874 ( .A(n21323), .B(n21324), .Z(n21326) );
  XOR U21875 ( .A(n21325), .B(n21326), .Z(n21258) );
  NANDN U21876 ( .A(n21121), .B(n21120), .Z(n21125) );
  NANDN U21877 ( .A(n21123), .B(n21122), .Z(n21124) );
  AND U21878 ( .A(n21125), .B(n21124), .Z(n21311) );
  NANDN U21879 ( .A(n21127), .B(n21126), .Z(n21131) );
  NANDN U21880 ( .A(n21129), .B(n21128), .Z(n21130) );
  NAND U21881 ( .A(n21131), .B(n21130), .Z(n21312) );
  XNOR U21882 ( .A(n21311), .B(n21312), .Z(n21313) );
  NANDN U21883 ( .A(n21133), .B(n21132), .Z(n21137) );
  NANDN U21884 ( .A(n21135), .B(n21134), .Z(n21136) );
  NAND U21885 ( .A(n21137), .B(n21136), .Z(n21314) );
  XNOR U21886 ( .A(n21313), .B(n21314), .Z(n21257) );
  XNOR U21887 ( .A(n21258), .B(n21257), .Z(n21260) );
  NANDN U21888 ( .A(n21139), .B(n21138), .Z(n21143) );
  NANDN U21889 ( .A(n21141), .B(n21140), .Z(n21142) );
  AND U21890 ( .A(n21143), .B(n21142), .Z(n21259) );
  XOR U21891 ( .A(n21260), .B(n21259), .Z(n21373) );
  NANDN U21892 ( .A(n21145), .B(n21144), .Z(n21149) );
  NANDN U21893 ( .A(n21147), .B(n21146), .Z(n21148) );
  AND U21894 ( .A(n21149), .B(n21148), .Z(n21371) );
  NANDN U21895 ( .A(n21151), .B(n21150), .Z(n21155) );
  NANDN U21896 ( .A(n21153), .B(n21152), .Z(n21154) );
  AND U21897 ( .A(n21155), .B(n21154), .Z(n21254) );
  NANDN U21898 ( .A(n21157), .B(n21156), .Z(n21161) );
  OR U21899 ( .A(n21159), .B(n21158), .Z(n21160) );
  AND U21900 ( .A(n21161), .B(n21160), .Z(n21252) );
  NANDN U21901 ( .A(n21163), .B(n21162), .Z(n21167) );
  NANDN U21902 ( .A(n21165), .B(n21164), .Z(n21166) );
  AND U21903 ( .A(n21167), .B(n21166), .Z(n21318) );
  NANDN U21904 ( .A(n21169), .B(n21168), .Z(n21173) );
  NANDN U21905 ( .A(n21171), .B(n21170), .Z(n21172) );
  NAND U21906 ( .A(n21173), .B(n21172), .Z(n21317) );
  XNOR U21907 ( .A(n21318), .B(n21317), .Z(n21319) );
  NAND U21908 ( .A(b[0]), .B(a[157]), .Z(n21174) );
  XNOR U21909 ( .A(b[1]), .B(n21174), .Z(n21176) );
  NANDN U21910 ( .A(b[0]), .B(a[156]), .Z(n21175) );
  NAND U21911 ( .A(n21176), .B(n21175), .Z(n21266) );
  NAND U21912 ( .A(n194), .B(n21177), .Z(n21179) );
  XOR U21913 ( .A(b[29]), .B(a[129]), .Z(n21344) );
  NAND U21914 ( .A(n38456), .B(n21344), .Z(n21178) );
  AND U21915 ( .A(n21179), .B(n21178), .Z(n21264) );
  AND U21916 ( .A(b[31]), .B(a[125]), .Z(n21263) );
  XNOR U21917 ( .A(n21264), .B(n21263), .Z(n21265) );
  XNOR U21918 ( .A(n21266), .B(n21265), .Z(n21305) );
  NAND U21919 ( .A(n38185), .B(n21180), .Z(n21182) );
  XOR U21920 ( .A(b[23]), .B(a[135]), .Z(n21347) );
  NAND U21921 ( .A(n38132), .B(n21347), .Z(n21181) );
  AND U21922 ( .A(n21182), .B(n21181), .Z(n21338) );
  NAND U21923 ( .A(n184), .B(n21183), .Z(n21185) );
  XOR U21924 ( .A(b[7]), .B(a[151]), .Z(n21350) );
  NAND U21925 ( .A(n36592), .B(n21350), .Z(n21184) );
  AND U21926 ( .A(n21185), .B(n21184), .Z(n21336) );
  NAND U21927 ( .A(n38289), .B(n21186), .Z(n21188) );
  XOR U21928 ( .A(b[25]), .B(a[133]), .Z(n21353) );
  NAND U21929 ( .A(n38247), .B(n21353), .Z(n21187) );
  NAND U21930 ( .A(n21188), .B(n21187), .Z(n21335) );
  XNOR U21931 ( .A(n21336), .B(n21335), .Z(n21337) );
  XOR U21932 ( .A(n21338), .B(n21337), .Z(n21306) );
  XNOR U21933 ( .A(n21305), .B(n21306), .Z(n21307) );
  NAND U21934 ( .A(n187), .B(n21189), .Z(n21191) );
  XOR U21935 ( .A(b[13]), .B(a[145]), .Z(n21356) );
  NAND U21936 ( .A(n37295), .B(n21356), .Z(n21190) );
  AND U21937 ( .A(n21191), .B(n21190), .Z(n21300) );
  NAND U21938 ( .A(n186), .B(n21192), .Z(n21194) );
  XOR U21939 ( .A(b[11]), .B(a[147]), .Z(n21359) );
  NAND U21940 ( .A(n37097), .B(n21359), .Z(n21193) );
  NAND U21941 ( .A(n21194), .B(n21193), .Z(n21299) );
  XNOR U21942 ( .A(n21300), .B(n21299), .Z(n21301) );
  NAND U21943 ( .A(n188), .B(n21195), .Z(n21197) );
  XOR U21944 ( .A(b[15]), .B(a[143]), .Z(n21362) );
  NAND U21945 ( .A(n37382), .B(n21362), .Z(n21196) );
  AND U21946 ( .A(n21197), .B(n21196), .Z(n21296) );
  NAND U21947 ( .A(n38064), .B(n21198), .Z(n21200) );
  XOR U21948 ( .A(b[21]), .B(a[137]), .Z(n21365) );
  NAND U21949 ( .A(n37993), .B(n21365), .Z(n21199) );
  AND U21950 ( .A(n21200), .B(n21199), .Z(n21294) );
  NAND U21951 ( .A(n185), .B(n21201), .Z(n21203) );
  XOR U21952 ( .A(b[9]), .B(a[149]), .Z(n21368) );
  NAND U21953 ( .A(n36805), .B(n21368), .Z(n21202) );
  NAND U21954 ( .A(n21203), .B(n21202), .Z(n21293) );
  XNOR U21955 ( .A(n21294), .B(n21293), .Z(n21295) );
  XOR U21956 ( .A(n21296), .B(n21295), .Z(n21302) );
  XOR U21957 ( .A(n21301), .B(n21302), .Z(n21308) );
  XOR U21958 ( .A(n21307), .B(n21308), .Z(n21320) );
  XNOR U21959 ( .A(n21319), .B(n21320), .Z(n21251) );
  XNOR U21960 ( .A(n21252), .B(n21251), .Z(n21253) );
  XOR U21961 ( .A(n21254), .B(n21253), .Z(n21372) );
  XOR U21962 ( .A(n21371), .B(n21372), .Z(n21374) );
  XOR U21963 ( .A(n21373), .B(n21374), .Z(n21248) );
  NANDN U21964 ( .A(n21205), .B(n21204), .Z(n21209) );
  NAND U21965 ( .A(n21207), .B(n21206), .Z(n21208) );
  AND U21966 ( .A(n21209), .B(n21208), .Z(n21246) );
  NANDN U21967 ( .A(n21211), .B(n21210), .Z(n21215) );
  NANDN U21968 ( .A(n21213), .B(n21212), .Z(n21214) );
  AND U21969 ( .A(n21215), .B(n21214), .Z(n21245) );
  XNOR U21970 ( .A(n21246), .B(n21245), .Z(n21247) );
  XNOR U21971 ( .A(n21248), .B(n21247), .Z(n21239) );
  NANDN U21972 ( .A(n21217), .B(n21216), .Z(n21221) );
  NANDN U21973 ( .A(n21219), .B(n21218), .Z(n21220) );
  NAND U21974 ( .A(n21221), .B(n21220), .Z(n21240) );
  XNOR U21975 ( .A(n21239), .B(n21240), .Z(n21241) );
  NANDN U21976 ( .A(n21223), .B(n21222), .Z(n21227) );
  NAND U21977 ( .A(n21225), .B(n21224), .Z(n21226) );
  NAND U21978 ( .A(n21227), .B(n21226), .Z(n21242) );
  XNOR U21979 ( .A(n21241), .B(n21242), .Z(n21233) );
  XNOR U21980 ( .A(n21234), .B(n21233), .Z(n21235) );
  XNOR U21981 ( .A(n21236), .B(n21235), .Z(n21377) );
  XNOR U21982 ( .A(sreg[381]), .B(n21377), .Z(n21379) );
  NANDN U21983 ( .A(sreg[380]), .B(n21228), .Z(n21232) );
  NAND U21984 ( .A(n21230), .B(n21229), .Z(n21231) );
  NAND U21985 ( .A(n21232), .B(n21231), .Z(n21378) );
  XNOR U21986 ( .A(n21379), .B(n21378), .Z(c[381]) );
  NANDN U21987 ( .A(n21234), .B(n21233), .Z(n21238) );
  NANDN U21988 ( .A(n21236), .B(n21235), .Z(n21237) );
  AND U21989 ( .A(n21238), .B(n21237), .Z(n21385) );
  NANDN U21990 ( .A(n21240), .B(n21239), .Z(n21244) );
  NANDN U21991 ( .A(n21242), .B(n21241), .Z(n21243) );
  AND U21992 ( .A(n21244), .B(n21243), .Z(n21383) );
  NANDN U21993 ( .A(n21246), .B(n21245), .Z(n21250) );
  NANDN U21994 ( .A(n21248), .B(n21247), .Z(n21249) );
  AND U21995 ( .A(n21250), .B(n21249), .Z(n21391) );
  NANDN U21996 ( .A(n21252), .B(n21251), .Z(n21256) );
  NANDN U21997 ( .A(n21254), .B(n21253), .Z(n21255) );
  AND U21998 ( .A(n21256), .B(n21255), .Z(n21395) );
  NANDN U21999 ( .A(n21258), .B(n21257), .Z(n21262) );
  NAND U22000 ( .A(n21260), .B(n21259), .Z(n21261) );
  AND U22001 ( .A(n21262), .B(n21261), .Z(n21394) );
  XNOR U22002 ( .A(n21395), .B(n21394), .Z(n21397) );
  NANDN U22003 ( .A(n21264), .B(n21263), .Z(n21268) );
  NANDN U22004 ( .A(n21266), .B(n21265), .Z(n21267) );
  AND U22005 ( .A(n21268), .B(n21267), .Z(n21474) );
  NAND U22006 ( .A(n38385), .B(n21269), .Z(n21271) );
  XOR U22007 ( .A(b[27]), .B(a[132]), .Z(n21418) );
  NAND U22008 ( .A(n38343), .B(n21418), .Z(n21270) );
  AND U22009 ( .A(n21271), .B(n21270), .Z(n21481) );
  NAND U22010 ( .A(n183), .B(n21272), .Z(n21274) );
  XOR U22011 ( .A(b[5]), .B(a[154]), .Z(n21421) );
  NAND U22012 ( .A(n36296), .B(n21421), .Z(n21273) );
  AND U22013 ( .A(n21274), .B(n21273), .Z(n21479) );
  NAND U22014 ( .A(n190), .B(n21275), .Z(n21277) );
  XOR U22015 ( .A(b[19]), .B(a[140]), .Z(n21424) );
  NAND U22016 ( .A(n37821), .B(n21424), .Z(n21276) );
  NAND U22017 ( .A(n21277), .B(n21276), .Z(n21478) );
  XNOR U22018 ( .A(n21479), .B(n21478), .Z(n21480) );
  XNOR U22019 ( .A(n21481), .B(n21480), .Z(n21472) );
  NAND U22020 ( .A(n38470), .B(n21278), .Z(n21280) );
  XOR U22021 ( .A(b[31]), .B(a[128]), .Z(n21427) );
  NAND U22022 ( .A(n38453), .B(n21427), .Z(n21279) );
  AND U22023 ( .A(n21280), .B(n21279), .Z(n21439) );
  NAND U22024 ( .A(n181), .B(n21281), .Z(n21283) );
  XOR U22025 ( .A(b[3]), .B(a[156]), .Z(n21430) );
  NAND U22026 ( .A(n182), .B(n21430), .Z(n21282) );
  AND U22027 ( .A(n21283), .B(n21282), .Z(n21437) );
  NAND U22028 ( .A(n189), .B(n21284), .Z(n21286) );
  XOR U22029 ( .A(b[17]), .B(a[142]), .Z(n21433) );
  NAND U22030 ( .A(n37652), .B(n21433), .Z(n21285) );
  NAND U22031 ( .A(n21286), .B(n21285), .Z(n21436) );
  XNOR U22032 ( .A(n21437), .B(n21436), .Z(n21438) );
  XOR U22033 ( .A(n21439), .B(n21438), .Z(n21473) );
  XOR U22034 ( .A(n21472), .B(n21473), .Z(n21475) );
  XOR U22035 ( .A(n21474), .B(n21475), .Z(n21407) );
  NANDN U22036 ( .A(n21288), .B(n21287), .Z(n21292) );
  NANDN U22037 ( .A(n21290), .B(n21289), .Z(n21291) );
  AND U22038 ( .A(n21292), .B(n21291), .Z(n21460) );
  NANDN U22039 ( .A(n21294), .B(n21293), .Z(n21298) );
  NANDN U22040 ( .A(n21296), .B(n21295), .Z(n21297) );
  NAND U22041 ( .A(n21298), .B(n21297), .Z(n21461) );
  XNOR U22042 ( .A(n21460), .B(n21461), .Z(n21462) );
  NANDN U22043 ( .A(n21300), .B(n21299), .Z(n21304) );
  NANDN U22044 ( .A(n21302), .B(n21301), .Z(n21303) );
  NAND U22045 ( .A(n21304), .B(n21303), .Z(n21463) );
  XNOR U22046 ( .A(n21462), .B(n21463), .Z(n21406) );
  XNOR U22047 ( .A(n21407), .B(n21406), .Z(n21409) );
  NANDN U22048 ( .A(n21306), .B(n21305), .Z(n21310) );
  NANDN U22049 ( .A(n21308), .B(n21307), .Z(n21309) );
  AND U22050 ( .A(n21310), .B(n21309), .Z(n21408) );
  XOR U22051 ( .A(n21409), .B(n21408), .Z(n21523) );
  NANDN U22052 ( .A(n21312), .B(n21311), .Z(n21316) );
  NANDN U22053 ( .A(n21314), .B(n21313), .Z(n21315) );
  AND U22054 ( .A(n21316), .B(n21315), .Z(n21520) );
  NANDN U22055 ( .A(n21318), .B(n21317), .Z(n21322) );
  NANDN U22056 ( .A(n21320), .B(n21319), .Z(n21321) );
  AND U22057 ( .A(n21322), .B(n21321), .Z(n21403) );
  NANDN U22058 ( .A(n21324), .B(n21323), .Z(n21328) );
  OR U22059 ( .A(n21326), .B(n21325), .Z(n21327) );
  AND U22060 ( .A(n21328), .B(n21327), .Z(n21401) );
  NANDN U22061 ( .A(n21330), .B(n21329), .Z(n21334) );
  NANDN U22062 ( .A(n21332), .B(n21331), .Z(n21333) );
  AND U22063 ( .A(n21334), .B(n21333), .Z(n21467) );
  NANDN U22064 ( .A(n21336), .B(n21335), .Z(n21340) );
  NANDN U22065 ( .A(n21338), .B(n21337), .Z(n21339) );
  NAND U22066 ( .A(n21340), .B(n21339), .Z(n21466) );
  XNOR U22067 ( .A(n21467), .B(n21466), .Z(n21468) );
  NAND U22068 ( .A(b[0]), .B(a[158]), .Z(n21341) );
  XNOR U22069 ( .A(b[1]), .B(n21341), .Z(n21343) );
  NANDN U22070 ( .A(b[0]), .B(a[157]), .Z(n21342) );
  NAND U22071 ( .A(n21343), .B(n21342), .Z(n21415) );
  NAND U22072 ( .A(n194), .B(n21344), .Z(n21346) );
  XOR U22073 ( .A(b[29]), .B(a[130]), .Z(n21493) );
  NAND U22074 ( .A(n38456), .B(n21493), .Z(n21345) );
  AND U22075 ( .A(n21346), .B(n21345), .Z(n21413) );
  AND U22076 ( .A(b[31]), .B(a[126]), .Z(n21412) );
  XNOR U22077 ( .A(n21413), .B(n21412), .Z(n21414) );
  XNOR U22078 ( .A(n21415), .B(n21414), .Z(n21454) );
  NAND U22079 ( .A(n38185), .B(n21347), .Z(n21349) );
  XOR U22080 ( .A(b[23]), .B(a[136]), .Z(n21496) );
  NAND U22081 ( .A(n38132), .B(n21496), .Z(n21348) );
  AND U22082 ( .A(n21349), .B(n21348), .Z(n21487) );
  NAND U22083 ( .A(n184), .B(n21350), .Z(n21352) );
  XOR U22084 ( .A(b[7]), .B(a[152]), .Z(n21499) );
  NAND U22085 ( .A(n36592), .B(n21499), .Z(n21351) );
  AND U22086 ( .A(n21352), .B(n21351), .Z(n21485) );
  NAND U22087 ( .A(n38289), .B(n21353), .Z(n21355) );
  XOR U22088 ( .A(b[25]), .B(a[134]), .Z(n21502) );
  NAND U22089 ( .A(n38247), .B(n21502), .Z(n21354) );
  NAND U22090 ( .A(n21355), .B(n21354), .Z(n21484) );
  XNOR U22091 ( .A(n21485), .B(n21484), .Z(n21486) );
  XOR U22092 ( .A(n21487), .B(n21486), .Z(n21455) );
  XNOR U22093 ( .A(n21454), .B(n21455), .Z(n21456) );
  NAND U22094 ( .A(n187), .B(n21356), .Z(n21358) );
  XOR U22095 ( .A(b[13]), .B(a[146]), .Z(n21505) );
  NAND U22096 ( .A(n37295), .B(n21505), .Z(n21357) );
  AND U22097 ( .A(n21358), .B(n21357), .Z(n21449) );
  NAND U22098 ( .A(n186), .B(n21359), .Z(n21361) );
  XOR U22099 ( .A(b[11]), .B(a[148]), .Z(n21508) );
  NAND U22100 ( .A(n37097), .B(n21508), .Z(n21360) );
  NAND U22101 ( .A(n21361), .B(n21360), .Z(n21448) );
  XNOR U22102 ( .A(n21449), .B(n21448), .Z(n21450) );
  NAND U22103 ( .A(n188), .B(n21362), .Z(n21364) );
  XOR U22104 ( .A(b[15]), .B(a[144]), .Z(n21511) );
  NAND U22105 ( .A(n37382), .B(n21511), .Z(n21363) );
  AND U22106 ( .A(n21364), .B(n21363), .Z(n21445) );
  NAND U22107 ( .A(n38064), .B(n21365), .Z(n21367) );
  XOR U22108 ( .A(b[21]), .B(a[138]), .Z(n21514) );
  NAND U22109 ( .A(n37993), .B(n21514), .Z(n21366) );
  AND U22110 ( .A(n21367), .B(n21366), .Z(n21443) );
  NAND U22111 ( .A(n185), .B(n21368), .Z(n21370) );
  XOR U22112 ( .A(b[9]), .B(a[150]), .Z(n21517) );
  NAND U22113 ( .A(n36805), .B(n21517), .Z(n21369) );
  NAND U22114 ( .A(n21370), .B(n21369), .Z(n21442) );
  XNOR U22115 ( .A(n21443), .B(n21442), .Z(n21444) );
  XOR U22116 ( .A(n21445), .B(n21444), .Z(n21451) );
  XOR U22117 ( .A(n21450), .B(n21451), .Z(n21457) );
  XOR U22118 ( .A(n21456), .B(n21457), .Z(n21469) );
  XNOR U22119 ( .A(n21468), .B(n21469), .Z(n21400) );
  XNOR U22120 ( .A(n21401), .B(n21400), .Z(n21402) );
  XOR U22121 ( .A(n21403), .B(n21402), .Z(n21521) );
  XNOR U22122 ( .A(n21520), .B(n21521), .Z(n21522) );
  XNOR U22123 ( .A(n21523), .B(n21522), .Z(n21396) );
  XOR U22124 ( .A(n21397), .B(n21396), .Z(n21389) );
  NANDN U22125 ( .A(n21372), .B(n21371), .Z(n21376) );
  OR U22126 ( .A(n21374), .B(n21373), .Z(n21375) );
  AND U22127 ( .A(n21376), .B(n21375), .Z(n21388) );
  XNOR U22128 ( .A(n21389), .B(n21388), .Z(n21390) );
  XNOR U22129 ( .A(n21391), .B(n21390), .Z(n21382) );
  XNOR U22130 ( .A(n21383), .B(n21382), .Z(n21384) );
  XNOR U22131 ( .A(n21385), .B(n21384), .Z(n21526) );
  XNOR U22132 ( .A(sreg[382]), .B(n21526), .Z(n21528) );
  NANDN U22133 ( .A(sreg[381]), .B(n21377), .Z(n21381) );
  NAND U22134 ( .A(n21379), .B(n21378), .Z(n21380) );
  NAND U22135 ( .A(n21381), .B(n21380), .Z(n21527) );
  XNOR U22136 ( .A(n21528), .B(n21527), .Z(c[382]) );
  NANDN U22137 ( .A(n21383), .B(n21382), .Z(n21387) );
  NANDN U22138 ( .A(n21385), .B(n21384), .Z(n21386) );
  AND U22139 ( .A(n21387), .B(n21386), .Z(n21534) );
  NANDN U22140 ( .A(n21389), .B(n21388), .Z(n21393) );
  NANDN U22141 ( .A(n21391), .B(n21390), .Z(n21392) );
  AND U22142 ( .A(n21393), .B(n21392), .Z(n21532) );
  NANDN U22143 ( .A(n21395), .B(n21394), .Z(n21399) );
  NAND U22144 ( .A(n21397), .B(n21396), .Z(n21398) );
  AND U22145 ( .A(n21399), .B(n21398), .Z(n21539) );
  NANDN U22146 ( .A(n21401), .B(n21400), .Z(n21405) );
  NANDN U22147 ( .A(n21403), .B(n21402), .Z(n21404) );
  AND U22148 ( .A(n21405), .B(n21404), .Z(n21670) );
  NANDN U22149 ( .A(n21407), .B(n21406), .Z(n21411) );
  NAND U22150 ( .A(n21409), .B(n21408), .Z(n21410) );
  AND U22151 ( .A(n21411), .B(n21410), .Z(n21669) );
  XNOR U22152 ( .A(n21670), .B(n21669), .Z(n21672) );
  NANDN U22153 ( .A(n21413), .B(n21412), .Z(n21417) );
  NANDN U22154 ( .A(n21415), .B(n21414), .Z(n21416) );
  AND U22155 ( .A(n21417), .B(n21416), .Z(n21617) );
  NAND U22156 ( .A(n38385), .B(n21418), .Z(n21420) );
  XOR U22157 ( .A(b[27]), .B(a[133]), .Z(n21561) );
  NAND U22158 ( .A(n38343), .B(n21561), .Z(n21419) );
  AND U22159 ( .A(n21420), .B(n21419), .Z(n21624) );
  NAND U22160 ( .A(n183), .B(n21421), .Z(n21423) );
  XOR U22161 ( .A(b[5]), .B(a[155]), .Z(n21564) );
  NAND U22162 ( .A(n36296), .B(n21564), .Z(n21422) );
  AND U22163 ( .A(n21423), .B(n21422), .Z(n21622) );
  NAND U22164 ( .A(n190), .B(n21424), .Z(n21426) );
  XOR U22165 ( .A(b[19]), .B(a[141]), .Z(n21567) );
  NAND U22166 ( .A(n37821), .B(n21567), .Z(n21425) );
  NAND U22167 ( .A(n21426), .B(n21425), .Z(n21621) );
  XNOR U22168 ( .A(n21622), .B(n21621), .Z(n21623) );
  XNOR U22169 ( .A(n21624), .B(n21623), .Z(n21615) );
  NAND U22170 ( .A(n38470), .B(n21427), .Z(n21429) );
  XOR U22171 ( .A(b[31]), .B(a[129]), .Z(n21570) );
  NAND U22172 ( .A(n38453), .B(n21570), .Z(n21428) );
  AND U22173 ( .A(n21429), .B(n21428), .Z(n21582) );
  NAND U22174 ( .A(n181), .B(n21430), .Z(n21432) );
  XOR U22175 ( .A(b[3]), .B(a[157]), .Z(n21573) );
  NAND U22176 ( .A(n182), .B(n21573), .Z(n21431) );
  AND U22177 ( .A(n21432), .B(n21431), .Z(n21580) );
  NAND U22178 ( .A(n189), .B(n21433), .Z(n21435) );
  XOR U22179 ( .A(b[17]), .B(a[143]), .Z(n21576) );
  NAND U22180 ( .A(n37652), .B(n21576), .Z(n21434) );
  NAND U22181 ( .A(n21435), .B(n21434), .Z(n21579) );
  XNOR U22182 ( .A(n21580), .B(n21579), .Z(n21581) );
  XOR U22183 ( .A(n21582), .B(n21581), .Z(n21616) );
  XOR U22184 ( .A(n21615), .B(n21616), .Z(n21618) );
  XOR U22185 ( .A(n21617), .B(n21618), .Z(n21550) );
  NANDN U22186 ( .A(n21437), .B(n21436), .Z(n21441) );
  NANDN U22187 ( .A(n21439), .B(n21438), .Z(n21440) );
  AND U22188 ( .A(n21441), .B(n21440), .Z(n21603) );
  NANDN U22189 ( .A(n21443), .B(n21442), .Z(n21447) );
  NANDN U22190 ( .A(n21445), .B(n21444), .Z(n21446) );
  NAND U22191 ( .A(n21447), .B(n21446), .Z(n21604) );
  XNOR U22192 ( .A(n21603), .B(n21604), .Z(n21605) );
  NANDN U22193 ( .A(n21449), .B(n21448), .Z(n21453) );
  NANDN U22194 ( .A(n21451), .B(n21450), .Z(n21452) );
  NAND U22195 ( .A(n21453), .B(n21452), .Z(n21606) );
  XNOR U22196 ( .A(n21605), .B(n21606), .Z(n21549) );
  XNOR U22197 ( .A(n21550), .B(n21549), .Z(n21552) );
  NANDN U22198 ( .A(n21455), .B(n21454), .Z(n21459) );
  NANDN U22199 ( .A(n21457), .B(n21456), .Z(n21458) );
  AND U22200 ( .A(n21459), .B(n21458), .Z(n21551) );
  XOR U22201 ( .A(n21552), .B(n21551), .Z(n21666) );
  NANDN U22202 ( .A(n21461), .B(n21460), .Z(n21465) );
  NANDN U22203 ( .A(n21463), .B(n21462), .Z(n21464) );
  AND U22204 ( .A(n21465), .B(n21464), .Z(n21663) );
  NANDN U22205 ( .A(n21467), .B(n21466), .Z(n21471) );
  NANDN U22206 ( .A(n21469), .B(n21468), .Z(n21470) );
  AND U22207 ( .A(n21471), .B(n21470), .Z(n21546) );
  NANDN U22208 ( .A(n21473), .B(n21472), .Z(n21477) );
  OR U22209 ( .A(n21475), .B(n21474), .Z(n21476) );
  AND U22210 ( .A(n21477), .B(n21476), .Z(n21544) );
  NANDN U22211 ( .A(n21479), .B(n21478), .Z(n21483) );
  NANDN U22212 ( .A(n21481), .B(n21480), .Z(n21482) );
  AND U22213 ( .A(n21483), .B(n21482), .Z(n21610) );
  NANDN U22214 ( .A(n21485), .B(n21484), .Z(n21489) );
  NANDN U22215 ( .A(n21487), .B(n21486), .Z(n21488) );
  NAND U22216 ( .A(n21489), .B(n21488), .Z(n21609) );
  XNOR U22217 ( .A(n21610), .B(n21609), .Z(n21611) );
  NAND U22218 ( .A(b[0]), .B(a[159]), .Z(n21490) );
  XNOR U22219 ( .A(b[1]), .B(n21490), .Z(n21492) );
  NANDN U22220 ( .A(b[0]), .B(a[158]), .Z(n21491) );
  NAND U22221 ( .A(n21492), .B(n21491), .Z(n21558) );
  NAND U22222 ( .A(n194), .B(n21493), .Z(n21495) );
  XOR U22223 ( .A(b[29]), .B(a[131]), .Z(n21633) );
  NAND U22224 ( .A(n38456), .B(n21633), .Z(n21494) );
  AND U22225 ( .A(n21495), .B(n21494), .Z(n21556) );
  AND U22226 ( .A(b[31]), .B(a[127]), .Z(n21555) );
  XNOR U22227 ( .A(n21556), .B(n21555), .Z(n21557) );
  XNOR U22228 ( .A(n21558), .B(n21557), .Z(n21597) );
  NAND U22229 ( .A(n38185), .B(n21496), .Z(n21498) );
  XOR U22230 ( .A(b[23]), .B(a[137]), .Z(n21639) );
  NAND U22231 ( .A(n38132), .B(n21639), .Z(n21497) );
  AND U22232 ( .A(n21498), .B(n21497), .Z(n21630) );
  NAND U22233 ( .A(n184), .B(n21499), .Z(n21501) );
  XOR U22234 ( .A(b[7]), .B(a[153]), .Z(n21642) );
  NAND U22235 ( .A(n36592), .B(n21642), .Z(n21500) );
  AND U22236 ( .A(n21501), .B(n21500), .Z(n21628) );
  NAND U22237 ( .A(n38289), .B(n21502), .Z(n21504) );
  XOR U22238 ( .A(b[25]), .B(a[135]), .Z(n21645) );
  NAND U22239 ( .A(n38247), .B(n21645), .Z(n21503) );
  NAND U22240 ( .A(n21504), .B(n21503), .Z(n21627) );
  XNOR U22241 ( .A(n21628), .B(n21627), .Z(n21629) );
  XOR U22242 ( .A(n21630), .B(n21629), .Z(n21598) );
  XNOR U22243 ( .A(n21597), .B(n21598), .Z(n21599) );
  NAND U22244 ( .A(n187), .B(n21505), .Z(n21507) );
  XOR U22245 ( .A(b[13]), .B(a[147]), .Z(n21648) );
  NAND U22246 ( .A(n37295), .B(n21648), .Z(n21506) );
  AND U22247 ( .A(n21507), .B(n21506), .Z(n21592) );
  NAND U22248 ( .A(n186), .B(n21508), .Z(n21510) );
  XOR U22249 ( .A(b[11]), .B(a[149]), .Z(n21651) );
  NAND U22250 ( .A(n37097), .B(n21651), .Z(n21509) );
  NAND U22251 ( .A(n21510), .B(n21509), .Z(n21591) );
  XNOR U22252 ( .A(n21592), .B(n21591), .Z(n21593) );
  NAND U22253 ( .A(n188), .B(n21511), .Z(n21513) );
  XOR U22254 ( .A(b[15]), .B(a[145]), .Z(n21654) );
  NAND U22255 ( .A(n37382), .B(n21654), .Z(n21512) );
  AND U22256 ( .A(n21513), .B(n21512), .Z(n21588) );
  NAND U22257 ( .A(n38064), .B(n21514), .Z(n21516) );
  XOR U22258 ( .A(b[21]), .B(a[139]), .Z(n21657) );
  NAND U22259 ( .A(n37993), .B(n21657), .Z(n21515) );
  AND U22260 ( .A(n21516), .B(n21515), .Z(n21586) );
  NAND U22261 ( .A(n185), .B(n21517), .Z(n21519) );
  XOR U22262 ( .A(b[9]), .B(a[151]), .Z(n21660) );
  NAND U22263 ( .A(n36805), .B(n21660), .Z(n21518) );
  NAND U22264 ( .A(n21519), .B(n21518), .Z(n21585) );
  XNOR U22265 ( .A(n21586), .B(n21585), .Z(n21587) );
  XOR U22266 ( .A(n21588), .B(n21587), .Z(n21594) );
  XOR U22267 ( .A(n21593), .B(n21594), .Z(n21600) );
  XOR U22268 ( .A(n21599), .B(n21600), .Z(n21612) );
  XNOR U22269 ( .A(n21611), .B(n21612), .Z(n21543) );
  XNOR U22270 ( .A(n21544), .B(n21543), .Z(n21545) );
  XOR U22271 ( .A(n21546), .B(n21545), .Z(n21664) );
  XNOR U22272 ( .A(n21663), .B(n21664), .Z(n21665) );
  XNOR U22273 ( .A(n21666), .B(n21665), .Z(n21671) );
  XOR U22274 ( .A(n21672), .B(n21671), .Z(n21538) );
  NANDN U22275 ( .A(n21521), .B(n21520), .Z(n21525) );
  NANDN U22276 ( .A(n21523), .B(n21522), .Z(n21524) );
  AND U22277 ( .A(n21525), .B(n21524), .Z(n21537) );
  XOR U22278 ( .A(n21538), .B(n21537), .Z(n21540) );
  XNOR U22279 ( .A(n21539), .B(n21540), .Z(n21531) );
  XNOR U22280 ( .A(n21532), .B(n21531), .Z(n21533) );
  XNOR U22281 ( .A(n21534), .B(n21533), .Z(n21675) );
  XNOR U22282 ( .A(sreg[383]), .B(n21675), .Z(n21677) );
  NANDN U22283 ( .A(sreg[382]), .B(n21526), .Z(n21530) );
  NAND U22284 ( .A(n21528), .B(n21527), .Z(n21529) );
  NAND U22285 ( .A(n21530), .B(n21529), .Z(n21676) );
  XNOR U22286 ( .A(n21677), .B(n21676), .Z(c[383]) );
  NANDN U22287 ( .A(n21532), .B(n21531), .Z(n21536) );
  NANDN U22288 ( .A(n21534), .B(n21533), .Z(n21535) );
  AND U22289 ( .A(n21536), .B(n21535), .Z(n21683) );
  NANDN U22290 ( .A(n21538), .B(n21537), .Z(n21542) );
  NANDN U22291 ( .A(n21540), .B(n21539), .Z(n21541) );
  AND U22292 ( .A(n21542), .B(n21541), .Z(n21681) );
  NANDN U22293 ( .A(n21544), .B(n21543), .Z(n21548) );
  NANDN U22294 ( .A(n21546), .B(n21545), .Z(n21547) );
  AND U22295 ( .A(n21548), .B(n21547), .Z(n21693) );
  NANDN U22296 ( .A(n21550), .B(n21549), .Z(n21554) );
  NAND U22297 ( .A(n21552), .B(n21551), .Z(n21553) );
  AND U22298 ( .A(n21554), .B(n21553), .Z(n21692) );
  XNOR U22299 ( .A(n21693), .B(n21692), .Z(n21695) );
  NANDN U22300 ( .A(n21556), .B(n21555), .Z(n21560) );
  NANDN U22301 ( .A(n21558), .B(n21557), .Z(n21559) );
  AND U22302 ( .A(n21560), .B(n21559), .Z(n21770) );
  NAND U22303 ( .A(n38385), .B(n21561), .Z(n21563) );
  XOR U22304 ( .A(b[27]), .B(a[134]), .Z(n21716) );
  NAND U22305 ( .A(n38343), .B(n21716), .Z(n21562) );
  AND U22306 ( .A(n21563), .B(n21562), .Z(n21777) );
  NAND U22307 ( .A(n183), .B(n21564), .Z(n21566) );
  XOR U22308 ( .A(b[5]), .B(a[156]), .Z(n21719) );
  NAND U22309 ( .A(n36296), .B(n21719), .Z(n21565) );
  AND U22310 ( .A(n21566), .B(n21565), .Z(n21775) );
  NAND U22311 ( .A(n190), .B(n21567), .Z(n21569) );
  XOR U22312 ( .A(b[19]), .B(a[142]), .Z(n21722) );
  NAND U22313 ( .A(n37821), .B(n21722), .Z(n21568) );
  NAND U22314 ( .A(n21569), .B(n21568), .Z(n21774) );
  XNOR U22315 ( .A(n21775), .B(n21774), .Z(n21776) );
  XNOR U22316 ( .A(n21777), .B(n21776), .Z(n21768) );
  NAND U22317 ( .A(n38470), .B(n21570), .Z(n21572) );
  XOR U22318 ( .A(b[31]), .B(a[130]), .Z(n21725) );
  NAND U22319 ( .A(n38453), .B(n21725), .Z(n21571) );
  AND U22320 ( .A(n21572), .B(n21571), .Z(n21737) );
  NAND U22321 ( .A(n181), .B(n21573), .Z(n21575) );
  XOR U22322 ( .A(b[3]), .B(a[158]), .Z(n21728) );
  NAND U22323 ( .A(n182), .B(n21728), .Z(n21574) );
  AND U22324 ( .A(n21575), .B(n21574), .Z(n21735) );
  NAND U22325 ( .A(n189), .B(n21576), .Z(n21578) );
  XOR U22326 ( .A(b[17]), .B(a[144]), .Z(n21731) );
  NAND U22327 ( .A(n37652), .B(n21731), .Z(n21577) );
  NAND U22328 ( .A(n21578), .B(n21577), .Z(n21734) );
  XNOR U22329 ( .A(n21735), .B(n21734), .Z(n21736) );
  XOR U22330 ( .A(n21737), .B(n21736), .Z(n21769) );
  XOR U22331 ( .A(n21768), .B(n21769), .Z(n21771) );
  XOR U22332 ( .A(n21770), .B(n21771), .Z(n21705) );
  NANDN U22333 ( .A(n21580), .B(n21579), .Z(n21584) );
  NANDN U22334 ( .A(n21582), .B(n21581), .Z(n21583) );
  AND U22335 ( .A(n21584), .B(n21583), .Z(n21758) );
  NANDN U22336 ( .A(n21586), .B(n21585), .Z(n21590) );
  NANDN U22337 ( .A(n21588), .B(n21587), .Z(n21589) );
  NAND U22338 ( .A(n21590), .B(n21589), .Z(n21759) );
  XNOR U22339 ( .A(n21758), .B(n21759), .Z(n21760) );
  NANDN U22340 ( .A(n21592), .B(n21591), .Z(n21596) );
  NANDN U22341 ( .A(n21594), .B(n21593), .Z(n21595) );
  NAND U22342 ( .A(n21596), .B(n21595), .Z(n21761) );
  XNOR U22343 ( .A(n21760), .B(n21761), .Z(n21704) );
  XNOR U22344 ( .A(n21705), .B(n21704), .Z(n21707) );
  NANDN U22345 ( .A(n21598), .B(n21597), .Z(n21602) );
  NANDN U22346 ( .A(n21600), .B(n21599), .Z(n21601) );
  AND U22347 ( .A(n21602), .B(n21601), .Z(n21706) );
  XOR U22348 ( .A(n21707), .B(n21706), .Z(n21819) );
  NANDN U22349 ( .A(n21604), .B(n21603), .Z(n21608) );
  NANDN U22350 ( .A(n21606), .B(n21605), .Z(n21607) );
  AND U22351 ( .A(n21608), .B(n21607), .Z(n21816) );
  NANDN U22352 ( .A(n21610), .B(n21609), .Z(n21614) );
  NANDN U22353 ( .A(n21612), .B(n21611), .Z(n21613) );
  AND U22354 ( .A(n21614), .B(n21613), .Z(n21701) );
  NANDN U22355 ( .A(n21616), .B(n21615), .Z(n21620) );
  OR U22356 ( .A(n21618), .B(n21617), .Z(n21619) );
  AND U22357 ( .A(n21620), .B(n21619), .Z(n21699) );
  NANDN U22358 ( .A(n21622), .B(n21621), .Z(n21626) );
  NANDN U22359 ( .A(n21624), .B(n21623), .Z(n21625) );
  AND U22360 ( .A(n21626), .B(n21625), .Z(n21765) );
  NANDN U22361 ( .A(n21628), .B(n21627), .Z(n21632) );
  NANDN U22362 ( .A(n21630), .B(n21629), .Z(n21631) );
  NAND U22363 ( .A(n21632), .B(n21631), .Z(n21764) );
  XNOR U22364 ( .A(n21765), .B(n21764), .Z(n21767) );
  NAND U22365 ( .A(n194), .B(n21633), .Z(n21635) );
  XOR U22366 ( .A(b[29]), .B(a[132]), .Z(n21789) );
  NAND U22367 ( .A(n38456), .B(n21789), .Z(n21634) );
  AND U22368 ( .A(n21635), .B(n21634), .Z(n21711) );
  AND U22369 ( .A(b[31]), .B(a[128]), .Z(n21710) );
  XNOR U22370 ( .A(n21711), .B(n21710), .Z(n21712) );
  NAND U22371 ( .A(b[0]), .B(a[160]), .Z(n21636) );
  XNOR U22372 ( .A(b[1]), .B(n21636), .Z(n21638) );
  NANDN U22373 ( .A(b[0]), .B(a[159]), .Z(n21637) );
  NAND U22374 ( .A(n21638), .B(n21637), .Z(n21713) );
  XNOR U22375 ( .A(n21712), .B(n21713), .Z(n21753) );
  NAND U22376 ( .A(n38185), .B(n21639), .Z(n21641) );
  XOR U22377 ( .A(b[23]), .B(a[138]), .Z(n21792) );
  NAND U22378 ( .A(n38132), .B(n21792), .Z(n21640) );
  AND U22379 ( .A(n21641), .B(n21640), .Z(n21782) );
  NAND U22380 ( .A(n184), .B(n21642), .Z(n21644) );
  XOR U22381 ( .A(b[7]), .B(a[154]), .Z(n21795) );
  NAND U22382 ( .A(n36592), .B(n21795), .Z(n21643) );
  AND U22383 ( .A(n21644), .B(n21643), .Z(n21781) );
  NAND U22384 ( .A(n38289), .B(n21645), .Z(n21647) );
  XOR U22385 ( .A(b[25]), .B(a[136]), .Z(n21798) );
  NAND U22386 ( .A(n38247), .B(n21798), .Z(n21646) );
  NAND U22387 ( .A(n21647), .B(n21646), .Z(n21780) );
  XOR U22388 ( .A(n21781), .B(n21780), .Z(n21783) );
  XOR U22389 ( .A(n21782), .B(n21783), .Z(n21752) );
  XOR U22390 ( .A(n21753), .B(n21752), .Z(n21755) );
  NAND U22391 ( .A(n187), .B(n21648), .Z(n21650) );
  XOR U22392 ( .A(b[13]), .B(a[148]), .Z(n21801) );
  NAND U22393 ( .A(n37295), .B(n21801), .Z(n21649) );
  AND U22394 ( .A(n21650), .B(n21649), .Z(n21747) );
  NAND U22395 ( .A(n186), .B(n21651), .Z(n21653) );
  XOR U22396 ( .A(b[11]), .B(a[150]), .Z(n21804) );
  NAND U22397 ( .A(n37097), .B(n21804), .Z(n21652) );
  NAND U22398 ( .A(n21653), .B(n21652), .Z(n21746) );
  XNOR U22399 ( .A(n21747), .B(n21746), .Z(n21749) );
  NAND U22400 ( .A(n188), .B(n21654), .Z(n21656) );
  XOR U22401 ( .A(b[15]), .B(a[146]), .Z(n21807) );
  NAND U22402 ( .A(n37382), .B(n21807), .Z(n21655) );
  AND U22403 ( .A(n21656), .B(n21655), .Z(n21743) );
  NAND U22404 ( .A(n38064), .B(n21657), .Z(n21659) );
  XOR U22405 ( .A(b[21]), .B(a[140]), .Z(n21810) );
  NAND U22406 ( .A(n37993), .B(n21810), .Z(n21658) );
  AND U22407 ( .A(n21659), .B(n21658), .Z(n21741) );
  NAND U22408 ( .A(n185), .B(n21660), .Z(n21662) );
  XOR U22409 ( .A(b[9]), .B(a[152]), .Z(n21813) );
  NAND U22410 ( .A(n36805), .B(n21813), .Z(n21661) );
  NAND U22411 ( .A(n21662), .B(n21661), .Z(n21740) );
  XNOR U22412 ( .A(n21741), .B(n21740), .Z(n21742) );
  XNOR U22413 ( .A(n21743), .B(n21742), .Z(n21748) );
  XOR U22414 ( .A(n21749), .B(n21748), .Z(n21754) );
  XNOR U22415 ( .A(n21755), .B(n21754), .Z(n21766) );
  XNOR U22416 ( .A(n21767), .B(n21766), .Z(n21698) );
  XNOR U22417 ( .A(n21699), .B(n21698), .Z(n21700) );
  XOR U22418 ( .A(n21701), .B(n21700), .Z(n21817) );
  XNOR U22419 ( .A(n21816), .B(n21817), .Z(n21818) );
  XNOR U22420 ( .A(n21819), .B(n21818), .Z(n21694) );
  XOR U22421 ( .A(n21695), .B(n21694), .Z(n21687) );
  NANDN U22422 ( .A(n21664), .B(n21663), .Z(n21668) );
  NANDN U22423 ( .A(n21666), .B(n21665), .Z(n21667) );
  AND U22424 ( .A(n21668), .B(n21667), .Z(n21686) );
  XNOR U22425 ( .A(n21687), .B(n21686), .Z(n21688) );
  NANDN U22426 ( .A(n21670), .B(n21669), .Z(n21674) );
  NAND U22427 ( .A(n21672), .B(n21671), .Z(n21673) );
  NAND U22428 ( .A(n21674), .B(n21673), .Z(n21689) );
  XNOR U22429 ( .A(n21688), .B(n21689), .Z(n21680) );
  XNOR U22430 ( .A(n21681), .B(n21680), .Z(n21682) );
  XNOR U22431 ( .A(n21683), .B(n21682), .Z(n21822) );
  XNOR U22432 ( .A(sreg[384]), .B(n21822), .Z(n21824) );
  NANDN U22433 ( .A(sreg[383]), .B(n21675), .Z(n21679) );
  NAND U22434 ( .A(n21677), .B(n21676), .Z(n21678) );
  NAND U22435 ( .A(n21679), .B(n21678), .Z(n21823) );
  XNOR U22436 ( .A(n21824), .B(n21823), .Z(c[384]) );
  NANDN U22437 ( .A(n21681), .B(n21680), .Z(n21685) );
  NANDN U22438 ( .A(n21683), .B(n21682), .Z(n21684) );
  AND U22439 ( .A(n21685), .B(n21684), .Z(n21830) );
  NANDN U22440 ( .A(n21687), .B(n21686), .Z(n21691) );
  NANDN U22441 ( .A(n21689), .B(n21688), .Z(n21690) );
  AND U22442 ( .A(n21691), .B(n21690), .Z(n21828) );
  NANDN U22443 ( .A(n21693), .B(n21692), .Z(n21697) );
  NAND U22444 ( .A(n21695), .B(n21694), .Z(n21696) );
  AND U22445 ( .A(n21697), .B(n21696), .Z(n21835) );
  NANDN U22446 ( .A(n21699), .B(n21698), .Z(n21703) );
  NANDN U22447 ( .A(n21701), .B(n21700), .Z(n21702) );
  AND U22448 ( .A(n21703), .B(n21702), .Z(n21840) );
  NANDN U22449 ( .A(n21705), .B(n21704), .Z(n21709) );
  NAND U22450 ( .A(n21707), .B(n21706), .Z(n21708) );
  AND U22451 ( .A(n21709), .B(n21708), .Z(n21839) );
  XNOR U22452 ( .A(n21840), .B(n21839), .Z(n21842) );
  NANDN U22453 ( .A(n21711), .B(n21710), .Z(n21715) );
  NANDN U22454 ( .A(n21713), .B(n21712), .Z(n21714) );
  AND U22455 ( .A(n21715), .B(n21714), .Z(n21907) );
  NAND U22456 ( .A(n38385), .B(n21716), .Z(n21718) );
  XOR U22457 ( .A(b[27]), .B(a[135]), .Z(n21851) );
  NAND U22458 ( .A(n38343), .B(n21851), .Z(n21717) );
  AND U22459 ( .A(n21718), .B(n21717), .Z(n21914) );
  NAND U22460 ( .A(n183), .B(n21719), .Z(n21721) );
  XOR U22461 ( .A(b[5]), .B(a[157]), .Z(n21854) );
  NAND U22462 ( .A(n36296), .B(n21854), .Z(n21720) );
  AND U22463 ( .A(n21721), .B(n21720), .Z(n21912) );
  NAND U22464 ( .A(n190), .B(n21722), .Z(n21724) );
  XOR U22465 ( .A(b[19]), .B(a[143]), .Z(n21857) );
  NAND U22466 ( .A(n37821), .B(n21857), .Z(n21723) );
  NAND U22467 ( .A(n21724), .B(n21723), .Z(n21911) );
  XNOR U22468 ( .A(n21912), .B(n21911), .Z(n21913) );
  XNOR U22469 ( .A(n21914), .B(n21913), .Z(n21905) );
  NAND U22470 ( .A(n38470), .B(n21725), .Z(n21727) );
  XOR U22471 ( .A(b[31]), .B(a[131]), .Z(n21860) );
  NAND U22472 ( .A(n38453), .B(n21860), .Z(n21726) );
  AND U22473 ( .A(n21727), .B(n21726), .Z(n21872) );
  NAND U22474 ( .A(n181), .B(n21728), .Z(n21730) );
  XOR U22475 ( .A(b[3]), .B(a[159]), .Z(n21863) );
  NAND U22476 ( .A(n182), .B(n21863), .Z(n21729) );
  AND U22477 ( .A(n21730), .B(n21729), .Z(n21870) );
  NAND U22478 ( .A(n189), .B(n21731), .Z(n21733) );
  XOR U22479 ( .A(b[17]), .B(a[145]), .Z(n21866) );
  NAND U22480 ( .A(n37652), .B(n21866), .Z(n21732) );
  NAND U22481 ( .A(n21733), .B(n21732), .Z(n21869) );
  XNOR U22482 ( .A(n21870), .B(n21869), .Z(n21871) );
  XOR U22483 ( .A(n21872), .B(n21871), .Z(n21906) );
  XOR U22484 ( .A(n21905), .B(n21906), .Z(n21908) );
  XOR U22485 ( .A(n21907), .B(n21908), .Z(n21954) );
  NANDN U22486 ( .A(n21735), .B(n21734), .Z(n21739) );
  NANDN U22487 ( .A(n21737), .B(n21736), .Z(n21738) );
  AND U22488 ( .A(n21739), .B(n21738), .Z(n21893) );
  NANDN U22489 ( .A(n21741), .B(n21740), .Z(n21745) );
  NANDN U22490 ( .A(n21743), .B(n21742), .Z(n21744) );
  NAND U22491 ( .A(n21745), .B(n21744), .Z(n21894) );
  XNOR U22492 ( .A(n21893), .B(n21894), .Z(n21895) );
  NANDN U22493 ( .A(n21747), .B(n21746), .Z(n21751) );
  NAND U22494 ( .A(n21749), .B(n21748), .Z(n21750) );
  NAND U22495 ( .A(n21751), .B(n21750), .Z(n21896) );
  XNOR U22496 ( .A(n21895), .B(n21896), .Z(n21953) );
  XNOR U22497 ( .A(n21954), .B(n21953), .Z(n21956) );
  NAND U22498 ( .A(n21753), .B(n21752), .Z(n21757) );
  NAND U22499 ( .A(n21755), .B(n21754), .Z(n21756) );
  AND U22500 ( .A(n21757), .B(n21756), .Z(n21955) );
  XOR U22501 ( .A(n21956), .B(n21955), .Z(n21968) );
  NANDN U22502 ( .A(n21759), .B(n21758), .Z(n21763) );
  NANDN U22503 ( .A(n21761), .B(n21760), .Z(n21762) );
  AND U22504 ( .A(n21763), .B(n21762), .Z(n21965) );
  NANDN U22505 ( .A(n21769), .B(n21768), .Z(n21773) );
  OR U22506 ( .A(n21771), .B(n21770), .Z(n21772) );
  AND U22507 ( .A(n21773), .B(n21772), .Z(n21960) );
  NANDN U22508 ( .A(n21775), .B(n21774), .Z(n21779) );
  NANDN U22509 ( .A(n21777), .B(n21776), .Z(n21778) );
  AND U22510 ( .A(n21779), .B(n21778), .Z(n21900) );
  NANDN U22511 ( .A(n21781), .B(n21780), .Z(n21785) );
  OR U22512 ( .A(n21783), .B(n21782), .Z(n21784) );
  NAND U22513 ( .A(n21785), .B(n21784), .Z(n21899) );
  XNOR U22514 ( .A(n21900), .B(n21899), .Z(n21901) );
  NAND U22515 ( .A(b[0]), .B(a[161]), .Z(n21786) );
  XNOR U22516 ( .A(b[1]), .B(n21786), .Z(n21788) );
  NANDN U22517 ( .A(b[0]), .B(a[160]), .Z(n21787) );
  NAND U22518 ( .A(n21788), .B(n21787), .Z(n21848) );
  NAND U22519 ( .A(n194), .B(n21789), .Z(n21791) );
  XOR U22520 ( .A(b[29]), .B(a[133]), .Z(n21926) );
  NAND U22521 ( .A(n38456), .B(n21926), .Z(n21790) );
  AND U22522 ( .A(n21791), .B(n21790), .Z(n21846) );
  AND U22523 ( .A(b[31]), .B(a[129]), .Z(n21845) );
  XNOR U22524 ( .A(n21846), .B(n21845), .Z(n21847) );
  XNOR U22525 ( .A(n21848), .B(n21847), .Z(n21887) );
  NAND U22526 ( .A(n38185), .B(n21792), .Z(n21794) );
  XOR U22527 ( .A(b[23]), .B(a[139]), .Z(n21929) );
  NAND U22528 ( .A(n38132), .B(n21929), .Z(n21793) );
  AND U22529 ( .A(n21794), .B(n21793), .Z(n21920) );
  NAND U22530 ( .A(n184), .B(n21795), .Z(n21797) );
  XOR U22531 ( .A(b[7]), .B(a[155]), .Z(n21932) );
  NAND U22532 ( .A(n36592), .B(n21932), .Z(n21796) );
  AND U22533 ( .A(n21797), .B(n21796), .Z(n21918) );
  NAND U22534 ( .A(n38289), .B(n21798), .Z(n21800) );
  XOR U22535 ( .A(b[25]), .B(a[137]), .Z(n21935) );
  NAND U22536 ( .A(n38247), .B(n21935), .Z(n21799) );
  NAND U22537 ( .A(n21800), .B(n21799), .Z(n21917) );
  XNOR U22538 ( .A(n21918), .B(n21917), .Z(n21919) );
  XOR U22539 ( .A(n21920), .B(n21919), .Z(n21888) );
  XNOR U22540 ( .A(n21887), .B(n21888), .Z(n21889) );
  NAND U22541 ( .A(n187), .B(n21801), .Z(n21803) );
  XOR U22542 ( .A(b[13]), .B(a[149]), .Z(n21938) );
  NAND U22543 ( .A(n37295), .B(n21938), .Z(n21802) );
  AND U22544 ( .A(n21803), .B(n21802), .Z(n21882) );
  NAND U22545 ( .A(n186), .B(n21804), .Z(n21806) );
  XOR U22546 ( .A(b[11]), .B(a[151]), .Z(n21941) );
  NAND U22547 ( .A(n37097), .B(n21941), .Z(n21805) );
  NAND U22548 ( .A(n21806), .B(n21805), .Z(n21881) );
  XNOR U22549 ( .A(n21882), .B(n21881), .Z(n21883) );
  NAND U22550 ( .A(n188), .B(n21807), .Z(n21809) );
  XOR U22551 ( .A(b[15]), .B(a[147]), .Z(n21944) );
  NAND U22552 ( .A(n37382), .B(n21944), .Z(n21808) );
  AND U22553 ( .A(n21809), .B(n21808), .Z(n21878) );
  NAND U22554 ( .A(n38064), .B(n21810), .Z(n21812) );
  XOR U22555 ( .A(b[21]), .B(a[141]), .Z(n21947) );
  NAND U22556 ( .A(n37993), .B(n21947), .Z(n21811) );
  AND U22557 ( .A(n21812), .B(n21811), .Z(n21876) );
  NAND U22558 ( .A(n185), .B(n21813), .Z(n21815) );
  XOR U22559 ( .A(b[9]), .B(a[153]), .Z(n21950) );
  NAND U22560 ( .A(n36805), .B(n21950), .Z(n21814) );
  NAND U22561 ( .A(n21815), .B(n21814), .Z(n21875) );
  XNOR U22562 ( .A(n21876), .B(n21875), .Z(n21877) );
  XOR U22563 ( .A(n21878), .B(n21877), .Z(n21884) );
  XOR U22564 ( .A(n21883), .B(n21884), .Z(n21890) );
  XOR U22565 ( .A(n21889), .B(n21890), .Z(n21902) );
  XNOR U22566 ( .A(n21901), .B(n21902), .Z(n21959) );
  XNOR U22567 ( .A(n21960), .B(n21959), .Z(n21961) );
  XOR U22568 ( .A(n21962), .B(n21961), .Z(n21966) );
  XNOR U22569 ( .A(n21965), .B(n21966), .Z(n21967) );
  XNOR U22570 ( .A(n21968), .B(n21967), .Z(n21841) );
  XOR U22571 ( .A(n21842), .B(n21841), .Z(n21834) );
  NANDN U22572 ( .A(n21817), .B(n21816), .Z(n21821) );
  NANDN U22573 ( .A(n21819), .B(n21818), .Z(n21820) );
  AND U22574 ( .A(n21821), .B(n21820), .Z(n21833) );
  XOR U22575 ( .A(n21834), .B(n21833), .Z(n21836) );
  XNOR U22576 ( .A(n21835), .B(n21836), .Z(n21827) );
  XNOR U22577 ( .A(n21828), .B(n21827), .Z(n21829) );
  XNOR U22578 ( .A(n21830), .B(n21829), .Z(n21971) );
  XNOR U22579 ( .A(sreg[385]), .B(n21971), .Z(n21973) );
  NANDN U22580 ( .A(sreg[384]), .B(n21822), .Z(n21826) );
  NAND U22581 ( .A(n21824), .B(n21823), .Z(n21825) );
  NAND U22582 ( .A(n21826), .B(n21825), .Z(n21972) );
  XNOR U22583 ( .A(n21973), .B(n21972), .Z(c[385]) );
  NANDN U22584 ( .A(n21828), .B(n21827), .Z(n21832) );
  NANDN U22585 ( .A(n21830), .B(n21829), .Z(n21831) );
  AND U22586 ( .A(n21832), .B(n21831), .Z(n21979) );
  NANDN U22587 ( .A(n21834), .B(n21833), .Z(n21838) );
  NANDN U22588 ( .A(n21836), .B(n21835), .Z(n21837) );
  AND U22589 ( .A(n21838), .B(n21837), .Z(n21977) );
  NANDN U22590 ( .A(n21840), .B(n21839), .Z(n21844) );
  NAND U22591 ( .A(n21842), .B(n21841), .Z(n21843) );
  AND U22592 ( .A(n21844), .B(n21843), .Z(n21984) );
  NANDN U22593 ( .A(n21846), .B(n21845), .Z(n21850) );
  NANDN U22594 ( .A(n21848), .B(n21847), .Z(n21849) );
  AND U22595 ( .A(n21850), .B(n21849), .Z(n22068) );
  NAND U22596 ( .A(n38385), .B(n21851), .Z(n21853) );
  XOR U22597 ( .A(b[27]), .B(a[136]), .Z(n22012) );
  NAND U22598 ( .A(n38343), .B(n22012), .Z(n21852) );
  AND U22599 ( .A(n21853), .B(n21852), .Z(n22075) );
  NAND U22600 ( .A(n183), .B(n21854), .Z(n21856) );
  XOR U22601 ( .A(b[5]), .B(a[158]), .Z(n22015) );
  NAND U22602 ( .A(n36296), .B(n22015), .Z(n21855) );
  AND U22603 ( .A(n21856), .B(n21855), .Z(n22073) );
  NAND U22604 ( .A(n190), .B(n21857), .Z(n21859) );
  XOR U22605 ( .A(b[19]), .B(a[144]), .Z(n22018) );
  NAND U22606 ( .A(n37821), .B(n22018), .Z(n21858) );
  NAND U22607 ( .A(n21859), .B(n21858), .Z(n22072) );
  XNOR U22608 ( .A(n22073), .B(n22072), .Z(n22074) );
  XNOR U22609 ( .A(n22075), .B(n22074), .Z(n22066) );
  NAND U22610 ( .A(n38470), .B(n21860), .Z(n21862) );
  XOR U22611 ( .A(b[31]), .B(a[132]), .Z(n22021) );
  NAND U22612 ( .A(n38453), .B(n22021), .Z(n21861) );
  AND U22613 ( .A(n21862), .B(n21861), .Z(n22033) );
  NAND U22614 ( .A(n181), .B(n21863), .Z(n21865) );
  XOR U22615 ( .A(b[3]), .B(a[160]), .Z(n22024) );
  NAND U22616 ( .A(n182), .B(n22024), .Z(n21864) );
  AND U22617 ( .A(n21865), .B(n21864), .Z(n22031) );
  NAND U22618 ( .A(n189), .B(n21866), .Z(n21868) );
  XOR U22619 ( .A(b[17]), .B(a[146]), .Z(n22027) );
  NAND U22620 ( .A(n37652), .B(n22027), .Z(n21867) );
  NAND U22621 ( .A(n21868), .B(n21867), .Z(n22030) );
  XNOR U22622 ( .A(n22031), .B(n22030), .Z(n22032) );
  XOR U22623 ( .A(n22033), .B(n22032), .Z(n22067) );
  XOR U22624 ( .A(n22066), .B(n22067), .Z(n22069) );
  XOR U22625 ( .A(n22068), .B(n22069), .Z(n22001) );
  NANDN U22626 ( .A(n21870), .B(n21869), .Z(n21874) );
  NANDN U22627 ( .A(n21872), .B(n21871), .Z(n21873) );
  AND U22628 ( .A(n21874), .B(n21873), .Z(n22054) );
  NANDN U22629 ( .A(n21876), .B(n21875), .Z(n21880) );
  NANDN U22630 ( .A(n21878), .B(n21877), .Z(n21879) );
  NAND U22631 ( .A(n21880), .B(n21879), .Z(n22055) );
  XNOR U22632 ( .A(n22054), .B(n22055), .Z(n22056) );
  NANDN U22633 ( .A(n21882), .B(n21881), .Z(n21886) );
  NANDN U22634 ( .A(n21884), .B(n21883), .Z(n21885) );
  NAND U22635 ( .A(n21886), .B(n21885), .Z(n22057) );
  XNOR U22636 ( .A(n22056), .B(n22057), .Z(n22000) );
  XNOR U22637 ( .A(n22001), .B(n22000), .Z(n22003) );
  NANDN U22638 ( .A(n21888), .B(n21887), .Z(n21892) );
  NANDN U22639 ( .A(n21890), .B(n21889), .Z(n21891) );
  AND U22640 ( .A(n21892), .B(n21891), .Z(n22002) );
  XOR U22641 ( .A(n22003), .B(n22002), .Z(n22116) );
  NANDN U22642 ( .A(n21894), .B(n21893), .Z(n21898) );
  NANDN U22643 ( .A(n21896), .B(n21895), .Z(n21897) );
  AND U22644 ( .A(n21898), .B(n21897), .Z(n22114) );
  NANDN U22645 ( .A(n21900), .B(n21899), .Z(n21904) );
  NANDN U22646 ( .A(n21902), .B(n21901), .Z(n21903) );
  AND U22647 ( .A(n21904), .B(n21903), .Z(n21997) );
  NANDN U22648 ( .A(n21906), .B(n21905), .Z(n21910) );
  OR U22649 ( .A(n21908), .B(n21907), .Z(n21909) );
  AND U22650 ( .A(n21910), .B(n21909), .Z(n21995) );
  NANDN U22651 ( .A(n21912), .B(n21911), .Z(n21916) );
  NANDN U22652 ( .A(n21914), .B(n21913), .Z(n21915) );
  AND U22653 ( .A(n21916), .B(n21915), .Z(n22061) );
  NANDN U22654 ( .A(n21918), .B(n21917), .Z(n21922) );
  NANDN U22655 ( .A(n21920), .B(n21919), .Z(n21921) );
  NAND U22656 ( .A(n21922), .B(n21921), .Z(n22060) );
  XNOR U22657 ( .A(n22061), .B(n22060), .Z(n22062) );
  NAND U22658 ( .A(b[0]), .B(a[162]), .Z(n21923) );
  XNOR U22659 ( .A(b[1]), .B(n21923), .Z(n21925) );
  NANDN U22660 ( .A(b[0]), .B(a[161]), .Z(n21924) );
  NAND U22661 ( .A(n21925), .B(n21924), .Z(n22009) );
  NAND U22662 ( .A(n194), .B(n21926), .Z(n21928) );
  XOR U22663 ( .A(b[29]), .B(a[134]), .Z(n22087) );
  NAND U22664 ( .A(n38456), .B(n22087), .Z(n21927) );
  AND U22665 ( .A(n21928), .B(n21927), .Z(n22007) );
  AND U22666 ( .A(b[31]), .B(a[130]), .Z(n22006) );
  XNOR U22667 ( .A(n22007), .B(n22006), .Z(n22008) );
  XNOR U22668 ( .A(n22009), .B(n22008), .Z(n22048) );
  NAND U22669 ( .A(n38185), .B(n21929), .Z(n21931) );
  XOR U22670 ( .A(b[23]), .B(a[140]), .Z(n22090) );
  NAND U22671 ( .A(n38132), .B(n22090), .Z(n21930) );
  AND U22672 ( .A(n21931), .B(n21930), .Z(n22081) );
  NAND U22673 ( .A(n184), .B(n21932), .Z(n21934) );
  XOR U22674 ( .A(b[7]), .B(a[156]), .Z(n22093) );
  NAND U22675 ( .A(n36592), .B(n22093), .Z(n21933) );
  AND U22676 ( .A(n21934), .B(n21933), .Z(n22079) );
  NAND U22677 ( .A(n38289), .B(n21935), .Z(n21937) );
  XOR U22678 ( .A(b[25]), .B(a[138]), .Z(n22096) );
  NAND U22679 ( .A(n38247), .B(n22096), .Z(n21936) );
  NAND U22680 ( .A(n21937), .B(n21936), .Z(n22078) );
  XNOR U22681 ( .A(n22079), .B(n22078), .Z(n22080) );
  XOR U22682 ( .A(n22081), .B(n22080), .Z(n22049) );
  XNOR U22683 ( .A(n22048), .B(n22049), .Z(n22050) );
  NAND U22684 ( .A(n187), .B(n21938), .Z(n21940) );
  XOR U22685 ( .A(b[13]), .B(a[150]), .Z(n22099) );
  NAND U22686 ( .A(n37295), .B(n22099), .Z(n21939) );
  AND U22687 ( .A(n21940), .B(n21939), .Z(n22043) );
  NAND U22688 ( .A(n186), .B(n21941), .Z(n21943) );
  XOR U22689 ( .A(b[11]), .B(a[152]), .Z(n22102) );
  NAND U22690 ( .A(n37097), .B(n22102), .Z(n21942) );
  NAND U22691 ( .A(n21943), .B(n21942), .Z(n22042) );
  XNOR U22692 ( .A(n22043), .B(n22042), .Z(n22044) );
  NAND U22693 ( .A(n188), .B(n21944), .Z(n21946) );
  XOR U22694 ( .A(b[15]), .B(a[148]), .Z(n22105) );
  NAND U22695 ( .A(n37382), .B(n22105), .Z(n21945) );
  AND U22696 ( .A(n21946), .B(n21945), .Z(n22039) );
  NAND U22697 ( .A(n38064), .B(n21947), .Z(n21949) );
  XOR U22698 ( .A(b[21]), .B(a[142]), .Z(n22108) );
  NAND U22699 ( .A(n37993), .B(n22108), .Z(n21948) );
  AND U22700 ( .A(n21949), .B(n21948), .Z(n22037) );
  NAND U22701 ( .A(n185), .B(n21950), .Z(n21952) );
  XOR U22702 ( .A(b[9]), .B(a[154]), .Z(n22111) );
  NAND U22703 ( .A(n36805), .B(n22111), .Z(n21951) );
  NAND U22704 ( .A(n21952), .B(n21951), .Z(n22036) );
  XNOR U22705 ( .A(n22037), .B(n22036), .Z(n22038) );
  XOR U22706 ( .A(n22039), .B(n22038), .Z(n22045) );
  XOR U22707 ( .A(n22044), .B(n22045), .Z(n22051) );
  XOR U22708 ( .A(n22050), .B(n22051), .Z(n22063) );
  XNOR U22709 ( .A(n22062), .B(n22063), .Z(n21994) );
  XNOR U22710 ( .A(n21995), .B(n21994), .Z(n21996) );
  XOR U22711 ( .A(n21997), .B(n21996), .Z(n22115) );
  XOR U22712 ( .A(n22114), .B(n22115), .Z(n22117) );
  XOR U22713 ( .A(n22116), .B(n22117), .Z(n21991) );
  NANDN U22714 ( .A(n21954), .B(n21953), .Z(n21958) );
  NAND U22715 ( .A(n21956), .B(n21955), .Z(n21957) );
  AND U22716 ( .A(n21958), .B(n21957), .Z(n21989) );
  NANDN U22717 ( .A(n21960), .B(n21959), .Z(n21964) );
  NANDN U22718 ( .A(n21962), .B(n21961), .Z(n21963) );
  AND U22719 ( .A(n21964), .B(n21963), .Z(n21988) );
  XNOR U22720 ( .A(n21989), .B(n21988), .Z(n21990) );
  XNOR U22721 ( .A(n21991), .B(n21990), .Z(n21982) );
  NANDN U22722 ( .A(n21966), .B(n21965), .Z(n21970) );
  NANDN U22723 ( .A(n21968), .B(n21967), .Z(n21969) );
  NAND U22724 ( .A(n21970), .B(n21969), .Z(n21983) );
  XOR U22725 ( .A(n21982), .B(n21983), .Z(n21985) );
  XNOR U22726 ( .A(n21984), .B(n21985), .Z(n21976) );
  XNOR U22727 ( .A(n21977), .B(n21976), .Z(n21978) );
  XNOR U22728 ( .A(n21979), .B(n21978), .Z(n22120) );
  XNOR U22729 ( .A(sreg[386]), .B(n22120), .Z(n22122) );
  NANDN U22730 ( .A(sreg[385]), .B(n21971), .Z(n21975) );
  NAND U22731 ( .A(n21973), .B(n21972), .Z(n21974) );
  NAND U22732 ( .A(n21975), .B(n21974), .Z(n22121) );
  XNOR U22733 ( .A(n22122), .B(n22121), .Z(c[386]) );
  NANDN U22734 ( .A(n21977), .B(n21976), .Z(n21981) );
  NANDN U22735 ( .A(n21979), .B(n21978), .Z(n21980) );
  AND U22736 ( .A(n21981), .B(n21980), .Z(n22128) );
  NANDN U22737 ( .A(n21983), .B(n21982), .Z(n21987) );
  NANDN U22738 ( .A(n21985), .B(n21984), .Z(n21986) );
  AND U22739 ( .A(n21987), .B(n21986), .Z(n22126) );
  NANDN U22740 ( .A(n21989), .B(n21988), .Z(n21993) );
  NANDN U22741 ( .A(n21991), .B(n21990), .Z(n21992) );
  AND U22742 ( .A(n21993), .B(n21992), .Z(n22134) );
  NANDN U22743 ( .A(n21995), .B(n21994), .Z(n21999) );
  NANDN U22744 ( .A(n21997), .B(n21996), .Z(n21998) );
  AND U22745 ( .A(n21999), .B(n21998), .Z(n22138) );
  NANDN U22746 ( .A(n22001), .B(n22000), .Z(n22005) );
  NAND U22747 ( .A(n22003), .B(n22002), .Z(n22004) );
  AND U22748 ( .A(n22005), .B(n22004), .Z(n22137) );
  XNOR U22749 ( .A(n22138), .B(n22137), .Z(n22140) );
  NANDN U22750 ( .A(n22007), .B(n22006), .Z(n22011) );
  NANDN U22751 ( .A(n22009), .B(n22008), .Z(n22010) );
  AND U22752 ( .A(n22011), .B(n22010), .Z(n22215) );
  NAND U22753 ( .A(n38385), .B(n22012), .Z(n22014) );
  XOR U22754 ( .A(b[27]), .B(a[137]), .Z(n22161) );
  NAND U22755 ( .A(n38343), .B(n22161), .Z(n22013) );
  AND U22756 ( .A(n22014), .B(n22013), .Z(n22222) );
  NAND U22757 ( .A(n183), .B(n22015), .Z(n22017) );
  XOR U22758 ( .A(b[5]), .B(a[159]), .Z(n22164) );
  NAND U22759 ( .A(n36296), .B(n22164), .Z(n22016) );
  AND U22760 ( .A(n22017), .B(n22016), .Z(n22220) );
  NAND U22761 ( .A(n190), .B(n22018), .Z(n22020) );
  XOR U22762 ( .A(b[19]), .B(a[145]), .Z(n22167) );
  NAND U22763 ( .A(n37821), .B(n22167), .Z(n22019) );
  NAND U22764 ( .A(n22020), .B(n22019), .Z(n22219) );
  XNOR U22765 ( .A(n22220), .B(n22219), .Z(n22221) );
  XNOR U22766 ( .A(n22222), .B(n22221), .Z(n22213) );
  NAND U22767 ( .A(n38470), .B(n22021), .Z(n22023) );
  XOR U22768 ( .A(b[31]), .B(a[133]), .Z(n22170) );
  NAND U22769 ( .A(n38453), .B(n22170), .Z(n22022) );
  AND U22770 ( .A(n22023), .B(n22022), .Z(n22182) );
  NAND U22771 ( .A(n181), .B(n22024), .Z(n22026) );
  XOR U22772 ( .A(b[3]), .B(a[161]), .Z(n22173) );
  NAND U22773 ( .A(n182), .B(n22173), .Z(n22025) );
  AND U22774 ( .A(n22026), .B(n22025), .Z(n22180) );
  NAND U22775 ( .A(n189), .B(n22027), .Z(n22029) );
  XOR U22776 ( .A(b[17]), .B(a[147]), .Z(n22176) );
  NAND U22777 ( .A(n37652), .B(n22176), .Z(n22028) );
  NAND U22778 ( .A(n22029), .B(n22028), .Z(n22179) );
  XNOR U22779 ( .A(n22180), .B(n22179), .Z(n22181) );
  XOR U22780 ( .A(n22182), .B(n22181), .Z(n22214) );
  XOR U22781 ( .A(n22213), .B(n22214), .Z(n22216) );
  XOR U22782 ( .A(n22215), .B(n22216), .Z(n22150) );
  NANDN U22783 ( .A(n22031), .B(n22030), .Z(n22035) );
  NANDN U22784 ( .A(n22033), .B(n22032), .Z(n22034) );
  AND U22785 ( .A(n22035), .B(n22034), .Z(n22203) );
  NANDN U22786 ( .A(n22037), .B(n22036), .Z(n22041) );
  NANDN U22787 ( .A(n22039), .B(n22038), .Z(n22040) );
  NAND U22788 ( .A(n22041), .B(n22040), .Z(n22204) );
  XNOR U22789 ( .A(n22203), .B(n22204), .Z(n22205) );
  NANDN U22790 ( .A(n22043), .B(n22042), .Z(n22047) );
  NANDN U22791 ( .A(n22045), .B(n22044), .Z(n22046) );
  NAND U22792 ( .A(n22047), .B(n22046), .Z(n22206) );
  XNOR U22793 ( .A(n22205), .B(n22206), .Z(n22149) );
  XNOR U22794 ( .A(n22150), .B(n22149), .Z(n22152) );
  NANDN U22795 ( .A(n22049), .B(n22048), .Z(n22053) );
  NANDN U22796 ( .A(n22051), .B(n22050), .Z(n22052) );
  AND U22797 ( .A(n22053), .B(n22052), .Z(n22151) );
  XOR U22798 ( .A(n22152), .B(n22151), .Z(n22264) );
  NANDN U22799 ( .A(n22055), .B(n22054), .Z(n22059) );
  NANDN U22800 ( .A(n22057), .B(n22056), .Z(n22058) );
  AND U22801 ( .A(n22059), .B(n22058), .Z(n22261) );
  NANDN U22802 ( .A(n22061), .B(n22060), .Z(n22065) );
  NANDN U22803 ( .A(n22063), .B(n22062), .Z(n22064) );
  AND U22804 ( .A(n22065), .B(n22064), .Z(n22146) );
  NANDN U22805 ( .A(n22067), .B(n22066), .Z(n22071) );
  OR U22806 ( .A(n22069), .B(n22068), .Z(n22070) );
  AND U22807 ( .A(n22071), .B(n22070), .Z(n22144) );
  NANDN U22808 ( .A(n22073), .B(n22072), .Z(n22077) );
  NANDN U22809 ( .A(n22075), .B(n22074), .Z(n22076) );
  AND U22810 ( .A(n22077), .B(n22076), .Z(n22210) );
  NANDN U22811 ( .A(n22079), .B(n22078), .Z(n22083) );
  NANDN U22812 ( .A(n22081), .B(n22080), .Z(n22082) );
  NAND U22813 ( .A(n22083), .B(n22082), .Z(n22209) );
  XNOR U22814 ( .A(n22210), .B(n22209), .Z(n22212) );
  NAND U22815 ( .A(b[0]), .B(a[163]), .Z(n22084) );
  XNOR U22816 ( .A(b[1]), .B(n22084), .Z(n22086) );
  NANDN U22817 ( .A(b[0]), .B(a[162]), .Z(n22085) );
  NAND U22818 ( .A(n22086), .B(n22085), .Z(n22158) );
  NAND U22819 ( .A(n194), .B(n22087), .Z(n22089) );
  XOR U22820 ( .A(b[29]), .B(a[135]), .Z(n22234) );
  NAND U22821 ( .A(n38456), .B(n22234), .Z(n22088) );
  AND U22822 ( .A(n22089), .B(n22088), .Z(n22156) );
  AND U22823 ( .A(b[31]), .B(a[131]), .Z(n22155) );
  XNOR U22824 ( .A(n22156), .B(n22155), .Z(n22157) );
  XNOR U22825 ( .A(n22158), .B(n22157), .Z(n22198) );
  NAND U22826 ( .A(n38185), .B(n22090), .Z(n22092) );
  XOR U22827 ( .A(b[23]), .B(a[141]), .Z(n22237) );
  NAND U22828 ( .A(n38132), .B(n22237), .Z(n22091) );
  AND U22829 ( .A(n22092), .B(n22091), .Z(n22227) );
  NAND U22830 ( .A(n184), .B(n22093), .Z(n22095) );
  XOR U22831 ( .A(b[7]), .B(a[157]), .Z(n22240) );
  NAND U22832 ( .A(n36592), .B(n22240), .Z(n22094) );
  AND U22833 ( .A(n22095), .B(n22094), .Z(n22226) );
  NAND U22834 ( .A(n38289), .B(n22096), .Z(n22098) );
  XOR U22835 ( .A(b[25]), .B(a[139]), .Z(n22243) );
  NAND U22836 ( .A(n38247), .B(n22243), .Z(n22097) );
  NAND U22837 ( .A(n22098), .B(n22097), .Z(n22225) );
  XOR U22838 ( .A(n22226), .B(n22225), .Z(n22228) );
  XOR U22839 ( .A(n22227), .B(n22228), .Z(n22197) );
  XOR U22840 ( .A(n22198), .B(n22197), .Z(n22200) );
  NAND U22841 ( .A(n187), .B(n22099), .Z(n22101) );
  XOR U22842 ( .A(b[13]), .B(a[151]), .Z(n22246) );
  NAND U22843 ( .A(n37295), .B(n22246), .Z(n22100) );
  AND U22844 ( .A(n22101), .B(n22100), .Z(n22192) );
  NAND U22845 ( .A(n186), .B(n22102), .Z(n22104) );
  XOR U22846 ( .A(b[11]), .B(a[153]), .Z(n22249) );
  NAND U22847 ( .A(n37097), .B(n22249), .Z(n22103) );
  NAND U22848 ( .A(n22104), .B(n22103), .Z(n22191) );
  XNOR U22849 ( .A(n22192), .B(n22191), .Z(n22194) );
  NAND U22850 ( .A(n188), .B(n22105), .Z(n22107) );
  XOR U22851 ( .A(b[15]), .B(a[149]), .Z(n22252) );
  NAND U22852 ( .A(n37382), .B(n22252), .Z(n22106) );
  AND U22853 ( .A(n22107), .B(n22106), .Z(n22188) );
  NAND U22854 ( .A(n38064), .B(n22108), .Z(n22110) );
  XOR U22855 ( .A(b[21]), .B(a[143]), .Z(n22255) );
  NAND U22856 ( .A(n37993), .B(n22255), .Z(n22109) );
  AND U22857 ( .A(n22110), .B(n22109), .Z(n22186) );
  NAND U22858 ( .A(n185), .B(n22111), .Z(n22113) );
  XOR U22859 ( .A(b[9]), .B(a[155]), .Z(n22258) );
  NAND U22860 ( .A(n36805), .B(n22258), .Z(n22112) );
  NAND U22861 ( .A(n22113), .B(n22112), .Z(n22185) );
  XNOR U22862 ( .A(n22186), .B(n22185), .Z(n22187) );
  XNOR U22863 ( .A(n22188), .B(n22187), .Z(n22193) );
  XOR U22864 ( .A(n22194), .B(n22193), .Z(n22199) );
  XNOR U22865 ( .A(n22200), .B(n22199), .Z(n22211) );
  XNOR U22866 ( .A(n22212), .B(n22211), .Z(n22143) );
  XNOR U22867 ( .A(n22144), .B(n22143), .Z(n22145) );
  XOR U22868 ( .A(n22146), .B(n22145), .Z(n22262) );
  XNOR U22869 ( .A(n22261), .B(n22262), .Z(n22263) );
  XNOR U22870 ( .A(n22264), .B(n22263), .Z(n22139) );
  XOR U22871 ( .A(n22140), .B(n22139), .Z(n22132) );
  NANDN U22872 ( .A(n22115), .B(n22114), .Z(n22119) );
  OR U22873 ( .A(n22117), .B(n22116), .Z(n22118) );
  AND U22874 ( .A(n22119), .B(n22118), .Z(n22131) );
  XNOR U22875 ( .A(n22132), .B(n22131), .Z(n22133) );
  XNOR U22876 ( .A(n22134), .B(n22133), .Z(n22125) );
  XNOR U22877 ( .A(n22126), .B(n22125), .Z(n22127) );
  XNOR U22878 ( .A(n22128), .B(n22127), .Z(n22267) );
  XNOR U22879 ( .A(sreg[387]), .B(n22267), .Z(n22269) );
  NANDN U22880 ( .A(sreg[386]), .B(n22120), .Z(n22124) );
  NAND U22881 ( .A(n22122), .B(n22121), .Z(n22123) );
  NAND U22882 ( .A(n22124), .B(n22123), .Z(n22268) );
  XNOR U22883 ( .A(n22269), .B(n22268), .Z(c[387]) );
  NANDN U22884 ( .A(n22126), .B(n22125), .Z(n22130) );
  NANDN U22885 ( .A(n22128), .B(n22127), .Z(n22129) );
  AND U22886 ( .A(n22130), .B(n22129), .Z(n22275) );
  NANDN U22887 ( .A(n22132), .B(n22131), .Z(n22136) );
  NANDN U22888 ( .A(n22134), .B(n22133), .Z(n22135) );
  AND U22889 ( .A(n22136), .B(n22135), .Z(n22273) );
  NANDN U22890 ( .A(n22138), .B(n22137), .Z(n22142) );
  NAND U22891 ( .A(n22140), .B(n22139), .Z(n22141) );
  AND U22892 ( .A(n22142), .B(n22141), .Z(n22280) );
  NANDN U22893 ( .A(n22144), .B(n22143), .Z(n22148) );
  NANDN U22894 ( .A(n22146), .B(n22145), .Z(n22147) );
  AND U22895 ( .A(n22148), .B(n22147), .Z(n22411) );
  NANDN U22896 ( .A(n22150), .B(n22149), .Z(n22154) );
  NAND U22897 ( .A(n22152), .B(n22151), .Z(n22153) );
  AND U22898 ( .A(n22154), .B(n22153), .Z(n22410) );
  XNOR U22899 ( .A(n22411), .B(n22410), .Z(n22413) );
  NANDN U22900 ( .A(n22156), .B(n22155), .Z(n22160) );
  NANDN U22901 ( .A(n22158), .B(n22157), .Z(n22159) );
  AND U22902 ( .A(n22160), .B(n22159), .Z(n22346) );
  NAND U22903 ( .A(n38385), .B(n22161), .Z(n22163) );
  XOR U22904 ( .A(b[27]), .B(a[138]), .Z(n22290) );
  NAND U22905 ( .A(n38343), .B(n22290), .Z(n22162) );
  AND U22906 ( .A(n22163), .B(n22162), .Z(n22353) );
  NAND U22907 ( .A(n183), .B(n22164), .Z(n22166) );
  XOR U22908 ( .A(b[5]), .B(a[160]), .Z(n22293) );
  NAND U22909 ( .A(n36296), .B(n22293), .Z(n22165) );
  AND U22910 ( .A(n22166), .B(n22165), .Z(n22351) );
  NAND U22911 ( .A(n190), .B(n22167), .Z(n22169) );
  XOR U22912 ( .A(b[19]), .B(a[146]), .Z(n22296) );
  NAND U22913 ( .A(n37821), .B(n22296), .Z(n22168) );
  NAND U22914 ( .A(n22169), .B(n22168), .Z(n22350) );
  XNOR U22915 ( .A(n22351), .B(n22350), .Z(n22352) );
  XNOR U22916 ( .A(n22353), .B(n22352), .Z(n22344) );
  NAND U22917 ( .A(n38470), .B(n22170), .Z(n22172) );
  XOR U22918 ( .A(b[31]), .B(a[134]), .Z(n22299) );
  NAND U22919 ( .A(n38453), .B(n22299), .Z(n22171) );
  AND U22920 ( .A(n22172), .B(n22171), .Z(n22311) );
  NAND U22921 ( .A(n181), .B(n22173), .Z(n22175) );
  XOR U22922 ( .A(b[3]), .B(a[162]), .Z(n22302) );
  NAND U22923 ( .A(n182), .B(n22302), .Z(n22174) );
  AND U22924 ( .A(n22175), .B(n22174), .Z(n22309) );
  NAND U22925 ( .A(n189), .B(n22176), .Z(n22178) );
  XOR U22926 ( .A(b[17]), .B(a[148]), .Z(n22305) );
  NAND U22927 ( .A(n37652), .B(n22305), .Z(n22177) );
  NAND U22928 ( .A(n22178), .B(n22177), .Z(n22308) );
  XNOR U22929 ( .A(n22309), .B(n22308), .Z(n22310) );
  XOR U22930 ( .A(n22311), .B(n22310), .Z(n22345) );
  XOR U22931 ( .A(n22344), .B(n22345), .Z(n22347) );
  XOR U22932 ( .A(n22346), .B(n22347), .Z(n22393) );
  NANDN U22933 ( .A(n22180), .B(n22179), .Z(n22184) );
  NANDN U22934 ( .A(n22182), .B(n22181), .Z(n22183) );
  AND U22935 ( .A(n22184), .B(n22183), .Z(n22332) );
  NANDN U22936 ( .A(n22186), .B(n22185), .Z(n22190) );
  NANDN U22937 ( .A(n22188), .B(n22187), .Z(n22189) );
  NAND U22938 ( .A(n22190), .B(n22189), .Z(n22333) );
  XNOR U22939 ( .A(n22332), .B(n22333), .Z(n22334) );
  NANDN U22940 ( .A(n22192), .B(n22191), .Z(n22196) );
  NAND U22941 ( .A(n22194), .B(n22193), .Z(n22195) );
  NAND U22942 ( .A(n22196), .B(n22195), .Z(n22335) );
  XNOR U22943 ( .A(n22334), .B(n22335), .Z(n22392) );
  XNOR U22944 ( .A(n22393), .B(n22392), .Z(n22395) );
  NAND U22945 ( .A(n22198), .B(n22197), .Z(n22202) );
  NAND U22946 ( .A(n22200), .B(n22199), .Z(n22201) );
  AND U22947 ( .A(n22202), .B(n22201), .Z(n22394) );
  XOR U22948 ( .A(n22395), .B(n22394), .Z(n22407) );
  NANDN U22949 ( .A(n22204), .B(n22203), .Z(n22208) );
  NANDN U22950 ( .A(n22206), .B(n22205), .Z(n22207) );
  AND U22951 ( .A(n22208), .B(n22207), .Z(n22404) );
  NANDN U22952 ( .A(n22214), .B(n22213), .Z(n22218) );
  OR U22953 ( .A(n22216), .B(n22215), .Z(n22217) );
  AND U22954 ( .A(n22218), .B(n22217), .Z(n22399) );
  NANDN U22955 ( .A(n22220), .B(n22219), .Z(n22224) );
  NANDN U22956 ( .A(n22222), .B(n22221), .Z(n22223) );
  AND U22957 ( .A(n22224), .B(n22223), .Z(n22339) );
  NANDN U22958 ( .A(n22226), .B(n22225), .Z(n22230) );
  OR U22959 ( .A(n22228), .B(n22227), .Z(n22229) );
  NAND U22960 ( .A(n22230), .B(n22229), .Z(n22338) );
  XNOR U22961 ( .A(n22339), .B(n22338), .Z(n22340) );
  NAND U22962 ( .A(b[0]), .B(a[164]), .Z(n22231) );
  XNOR U22963 ( .A(b[1]), .B(n22231), .Z(n22233) );
  NANDN U22964 ( .A(b[0]), .B(a[163]), .Z(n22232) );
  NAND U22965 ( .A(n22233), .B(n22232), .Z(n22287) );
  NAND U22966 ( .A(n194), .B(n22234), .Z(n22236) );
  XOR U22967 ( .A(b[29]), .B(a[136]), .Z(n22365) );
  NAND U22968 ( .A(n38456), .B(n22365), .Z(n22235) );
  AND U22969 ( .A(n22236), .B(n22235), .Z(n22285) );
  AND U22970 ( .A(b[31]), .B(a[132]), .Z(n22284) );
  XNOR U22971 ( .A(n22285), .B(n22284), .Z(n22286) );
  XNOR U22972 ( .A(n22287), .B(n22286), .Z(n22326) );
  NAND U22973 ( .A(n38185), .B(n22237), .Z(n22239) );
  XOR U22974 ( .A(b[23]), .B(a[142]), .Z(n22368) );
  NAND U22975 ( .A(n38132), .B(n22368), .Z(n22238) );
  AND U22976 ( .A(n22239), .B(n22238), .Z(n22359) );
  NAND U22977 ( .A(n184), .B(n22240), .Z(n22242) );
  XOR U22978 ( .A(b[7]), .B(a[158]), .Z(n22371) );
  NAND U22979 ( .A(n36592), .B(n22371), .Z(n22241) );
  AND U22980 ( .A(n22242), .B(n22241), .Z(n22357) );
  NAND U22981 ( .A(n38289), .B(n22243), .Z(n22245) );
  XOR U22982 ( .A(b[25]), .B(a[140]), .Z(n22374) );
  NAND U22983 ( .A(n38247), .B(n22374), .Z(n22244) );
  NAND U22984 ( .A(n22245), .B(n22244), .Z(n22356) );
  XNOR U22985 ( .A(n22357), .B(n22356), .Z(n22358) );
  XOR U22986 ( .A(n22359), .B(n22358), .Z(n22327) );
  XNOR U22987 ( .A(n22326), .B(n22327), .Z(n22328) );
  NAND U22988 ( .A(n187), .B(n22246), .Z(n22248) );
  XOR U22989 ( .A(b[13]), .B(a[152]), .Z(n22377) );
  NAND U22990 ( .A(n37295), .B(n22377), .Z(n22247) );
  AND U22991 ( .A(n22248), .B(n22247), .Z(n22321) );
  NAND U22992 ( .A(n186), .B(n22249), .Z(n22251) );
  XOR U22993 ( .A(b[11]), .B(a[154]), .Z(n22380) );
  NAND U22994 ( .A(n37097), .B(n22380), .Z(n22250) );
  NAND U22995 ( .A(n22251), .B(n22250), .Z(n22320) );
  XNOR U22996 ( .A(n22321), .B(n22320), .Z(n22322) );
  NAND U22997 ( .A(n188), .B(n22252), .Z(n22254) );
  XOR U22998 ( .A(b[15]), .B(a[150]), .Z(n22383) );
  NAND U22999 ( .A(n37382), .B(n22383), .Z(n22253) );
  AND U23000 ( .A(n22254), .B(n22253), .Z(n22317) );
  NAND U23001 ( .A(n38064), .B(n22255), .Z(n22257) );
  XOR U23002 ( .A(b[21]), .B(a[144]), .Z(n22386) );
  NAND U23003 ( .A(n37993), .B(n22386), .Z(n22256) );
  AND U23004 ( .A(n22257), .B(n22256), .Z(n22315) );
  NAND U23005 ( .A(n185), .B(n22258), .Z(n22260) );
  XOR U23006 ( .A(b[9]), .B(a[156]), .Z(n22389) );
  NAND U23007 ( .A(n36805), .B(n22389), .Z(n22259) );
  NAND U23008 ( .A(n22260), .B(n22259), .Z(n22314) );
  XNOR U23009 ( .A(n22315), .B(n22314), .Z(n22316) );
  XOR U23010 ( .A(n22317), .B(n22316), .Z(n22323) );
  XOR U23011 ( .A(n22322), .B(n22323), .Z(n22329) );
  XOR U23012 ( .A(n22328), .B(n22329), .Z(n22341) );
  XNOR U23013 ( .A(n22340), .B(n22341), .Z(n22398) );
  XNOR U23014 ( .A(n22399), .B(n22398), .Z(n22400) );
  XOR U23015 ( .A(n22401), .B(n22400), .Z(n22405) );
  XNOR U23016 ( .A(n22404), .B(n22405), .Z(n22406) );
  XNOR U23017 ( .A(n22407), .B(n22406), .Z(n22412) );
  XOR U23018 ( .A(n22413), .B(n22412), .Z(n22279) );
  NANDN U23019 ( .A(n22262), .B(n22261), .Z(n22266) );
  NANDN U23020 ( .A(n22264), .B(n22263), .Z(n22265) );
  AND U23021 ( .A(n22266), .B(n22265), .Z(n22278) );
  XOR U23022 ( .A(n22279), .B(n22278), .Z(n22281) );
  XNOR U23023 ( .A(n22280), .B(n22281), .Z(n22272) );
  XNOR U23024 ( .A(n22273), .B(n22272), .Z(n22274) );
  XNOR U23025 ( .A(n22275), .B(n22274), .Z(n22416) );
  XNOR U23026 ( .A(sreg[388]), .B(n22416), .Z(n22418) );
  NANDN U23027 ( .A(sreg[387]), .B(n22267), .Z(n22271) );
  NAND U23028 ( .A(n22269), .B(n22268), .Z(n22270) );
  NAND U23029 ( .A(n22271), .B(n22270), .Z(n22417) );
  XNOR U23030 ( .A(n22418), .B(n22417), .Z(c[388]) );
  NANDN U23031 ( .A(n22273), .B(n22272), .Z(n22277) );
  NANDN U23032 ( .A(n22275), .B(n22274), .Z(n22276) );
  AND U23033 ( .A(n22277), .B(n22276), .Z(n22424) );
  NANDN U23034 ( .A(n22279), .B(n22278), .Z(n22283) );
  NANDN U23035 ( .A(n22281), .B(n22280), .Z(n22282) );
  AND U23036 ( .A(n22283), .B(n22282), .Z(n22422) );
  NANDN U23037 ( .A(n22285), .B(n22284), .Z(n22289) );
  NANDN U23038 ( .A(n22287), .B(n22286), .Z(n22288) );
  AND U23039 ( .A(n22289), .B(n22288), .Z(n22513) );
  NAND U23040 ( .A(n38385), .B(n22290), .Z(n22292) );
  XOR U23041 ( .A(b[27]), .B(a[139]), .Z(n22457) );
  NAND U23042 ( .A(n38343), .B(n22457), .Z(n22291) );
  AND U23043 ( .A(n22292), .B(n22291), .Z(n22520) );
  NAND U23044 ( .A(n183), .B(n22293), .Z(n22295) );
  XOR U23045 ( .A(b[5]), .B(a[161]), .Z(n22460) );
  NAND U23046 ( .A(n36296), .B(n22460), .Z(n22294) );
  AND U23047 ( .A(n22295), .B(n22294), .Z(n22518) );
  NAND U23048 ( .A(n190), .B(n22296), .Z(n22298) );
  XOR U23049 ( .A(b[19]), .B(a[147]), .Z(n22463) );
  NAND U23050 ( .A(n37821), .B(n22463), .Z(n22297) );
  NAND U23051 ( .A(n22298), .B(n22297), .Z(n22517) );
  XNOR U23052 ( .A(n22518), .B(n22517), .Z(n22519) );
  XNOR U23053 ( .A(n22520), .B(n22519), .Z(n22511) );
  NAND U23054 ( .A(n38470), .B(n22299), .Z(n22301) );
  XOR U23055 ( .A(b[31]), .B(a[135]), .Z(n22466) );
  NAND U23056 ( .A(n38453), .B(n22466), .Z(n22300) );
  AND U23057 ( .A(n22301), .B(n22300), .Z(n22478) );
  NAND U23058 ( .A(n181), .B(n22302), .Z(n22304) );
  XOR U23059 ( .A(b[3]), .B(a[163]), .Z(n22469) );
  NAND U23060 ( .A(n182), .B(n22469), .Z(n22303) );
  AND U23061 ( .A(n22304), .B(n22303), .Z(n22476) );
  NAND U23062 ( .A(n189), .B(n22305), .Z(n22307) );
  XOR U23063 ( .A(b[17]), .B(a[149]), .Z(n22472) );
  NAND U23064 ( .A(n37652), .B(n22472), .Z(n22306) );
  NAND U23065 ( .A(n22307), .B(n22306), .Z(n22475) );
  XNOR U23066 ( .A(n22476), .B(n22475), .Z(n22477) );
  XOR U23067 ( .A(n22478), .B(n22477), .Z(n22512) );
  XOR U23068 ( .A(n22511), .B(n22512), .Z(n22514) );
  XOR U23069 ( .A(n22513), .B(n22514), .Z(n22446) );
  NANDN U23070 ( .A(n22309), .B(n22308), .Z(n22313) );
  NANDN U23071 ( .A(n22311), .B(n22310), .Z(n22312) );
  AND U23072 ( .A(n22313), .B(n22312), .Z(n22499) );
  NANDN U23073 ( .A(n22315), .B(n22314), .Z(n22319) );
  NANDN U23074 ( .A(n22317), .B(n22316), .Z(n22318) );
  NAND U23075 ( .A(n22319), .B(n22318), .Z(n22500) );
  XNOR U23076 ( .A(n22499), .B(n22500), .Z(n22501) );
  NANDN U23077 ( .A(n22321), .B(n22320), .Z(n22325) );
  NANDN U23078 ( .A(n22323), .B(n22322), .Z(n22324) );
  NAND U23079 ( .A(n22325), .B(n22324), .Z(n22502) );
  XNOR U23080 ( .A(n22501), .B(n22502), .Z(n22445) );
  XNOR U23081 ( .A(n22446), .B(n22445), .Z(n22448) );
  NANDN U23082 ( .A(n22327), .B(n22326), .Z(n22331) );
  NANDN U23083 ( .A(n22329), .B(n22328), .Z(n22330) );
  AND U23084 ( .A(n22331), .B(n22330), .Z(n22447) );
  XOR U23085 ( .A(n22448), .B(n22447), .Z(n22561) );
  NANDN U23086 ( .A(n22333), .B(n22332), .Z(n22337) );
  NANDN U23087 ( .A(n22335), .B(n22334), .Z(n22336) );
  AND U23088 ( .A(n22337), .B(n22336), .Z(n22559) );
  NANDN U23089 ( .A(n22339), .B(n22338), .Z(n22343) );
  NANDN U23090 ( .A(n22341), .B(n22340), .Z(n22342) );
  AND U23091 ( .A(n22343), .B(n22342), .Z(n22442) );
  NANDN U23092 ( .A(n22345), .B(n22344), .Z(n22349) );
  OR U23093 ( .A(n22347), .B(n22346), .Z(n22348) );
  AND U23094 ( .A(n22349), .B(n22348), .Z(n22440) );
  NANDN U23095 ( .A(n22351), .B(n22350), .Z(n22355) );
  NANDN U23096 ( .A(n22353), .B(n22352), .Z(n22354) );
  AND U23097 ( .A(n22355), .B(n22354), .Z(n22506) );
  NANDN U23098 ( .A(n22357), .B(n22356), .Z(n22361) );
  NANDN U23099 ( .A(n22359), .B(n22358), .Z(n22360) );
  NAND U23100 ( .A(n22361), .B(n22360), .Z(n22505) );
  XNOR U23101 ( .A(n22506), .B(n22505), .Z(n22507) );
  NAND U23102 ( .A(b[0]), .B(a[165]), .Z(n22362) );
  XNOR U23103 ( .A(b[1]), .B(n22362), .Z(n22364) );
  NANDN U23104 ( .A(b[0]), .B(a[164]), .Z(n22363) );
  NAND U23105 ( .A(n22364), .B(n22363), .Z(n22454) );
  NAND U23106 ( .A(n194), .B(n22365), .Z(n22367) );
  XOR U23107 ( .A(b[29]), .B(a[137]), .Z(n22532) );
  NAND U23108 ( .A(n38456), .B(n22532), .Z(n22366) );
  AND U23109 ( .A(n22367), .B(n22366), .Z(n22452) );
  AND U23110 ( .A(b[31]), .B(a[133]), .Z(n22451) );
  XNOR U23111 ( .A(n22452), .B(n22451), .Z(n22453) );
  XNOR U23112 ( .A(n22454), .B(n22453), .Z(n22493) );
  NAND U23113 ( .A(n38185), .B(n22368), .Z(n22370) );
  XOR U23114 ( .A(b[23]), .B(a[143]), .Z(n22535) );
  NAND U23115 ( .A(n38132), .B(n22535), .Z(n22369) );
  AND U23116 ( .A(n22370), .B(n22369), .Z(n22526) );
  NAND U23117 ( .A(n184), .B(n22371), .Z(n22373) );
  XOR U23118 ( .A(b[7]), .B(a[159]), .Z(n22538) );
  NAND U23119 ( .A(n36592), .B(n22538), .Z(n22372) );
  AND U23120 ( .A(n22373), .B(n22372), .Z(n22524) );
  NAND U23121 ( .A(n38289), .B(n22374), .Z(n22376) );
  XOR U23122 ( .A(b[25]), .B(a[141]), .Z(n22541) );
  NAND U23123 ( .A(n38247), .B(n22541), .Z(n22375) );
  NAND U23124 ( .A(n22376), .B(n22375), .Z(n22523) );
  XNOR U23125 ( .A(n22524), .B(n22523), .Z(n22525) );
  XOR U23126 ( .A(n22526), .B(n22525), .Z(n22494) );
  XNOR U23127 ( .A(n22493), .B(n22494), .Z(n22495) );
  NAND U23128 ( .A(n187), .B(n22377), .Z(n22379) );
  XOR U23129 ( .A(b[13]), .B(a[153]), .Z(n22544) );
  NAND U23130 ( .A(n37295), .B(n22544), .Z(n22378) );
  AND U23131 ( .A(n22379), .B(n22378), .Z(n22488) );
  NAND U23132 ( .A(n186), .B(n22380), .Z(n22382) );
  XOR U23133 ( .A(b[11]), .B(a[155]), .Z(n22547) );
  NAND U23134 ( .A(n37097), .B(n22547), .Z(n22381) );
  NAND U23135 ( .A(n22382), .B(n22381), .Z(n22487) );
  XNOR U23136 ( .A(n22488), .B(n22487), .Z(n22489) );
  NAND U23137 ( .A(n188), .B(n22383), .Z(n22385) );
  XOR U23138 ( .A(b[15]), .B(a[151]), .Z(n22550) );
  NAND U23139 ( .A(n37382), .B(n22550), .Z(n22384) );
  AND U23140 ( .A(n22385), .B(n22384), .Z(n22484) );
  NAND U23141 ( .A(n38064), .B(n22386), .Z(n22388) );
  XOR U23142 ( .A(b[21]), .B(a[145]), .Z(n22553) );
  NAND U23143 ( .A(n37993), .B(n22553), .Z(n22387) );
  AND U23144 ( .A(n22388), .B(n22387), .Z(n22482) );
  NAND U23145 ( .A(n185), .B(n22389), .Z(n22391) );
  XOR U23146 ( .A(b[9]), .B(a[157]), .Z(n22556) );
  NAND U23147 ( .A(n36805), .B(n22556), .Z(n22390) );
  NAND U23148 ( .A(n22391), .B(n22390), .Z(n22481) );
  XNOR U23149 ( .A(n22482), .B(n22481), .Z(n22483) );
  XOR U23150 ( .A(n22484), .B(n22483), .Z(n22490) );
  XOR U23151 ( .A(n22489), .B(n22490), .Z(n22496) );
  XOR U23152 ( .A(n22495), .B(n22496), .Z(n22508) );
  XNOR U23153 ( .A(n22507), .B(n22508), .Z(n22439) );
  XNOR U23154 ( .A(n22440), .B(n22439), .Z(n22441) );
  XOR U23155 ( .A(n22442), .B(n22441), .Z(n22560) );
  XOR U23156 ( .A(n22559), .B(n22560), .Z(n22562) );
  XOR U23157 ( .A(n22561), .B(n22562), .Z(n22436) );
  NANDN U23158 ( .A(n22393), .B(n22392), .Z(n22397) );
  NAND U23159 ( .A(n22395), .B(n22394), .Z(n22396) );
  AND U23160 ( .A(n22397), .B(n22396), .Z(n22434) );
  NANDN U23161 ( .A(n22399), .B(n22398), .Z(n22403) );
  NANDN U23162 ( .A(n22401), .B(n22400), .Z(n22402) );
  AND U23163 ( .A(n22403), .B(n22402), .Z(n22433) );
  XNOR U23164 ( .A(n22434), .B(n22433), .Z(n22435) );
  XNOR U23165 ( .A(n22436), .B(n22435), .Z(n22427) );
  NANDN U23166 ( .A(n22405), .B(n22404), .Z(n22409) );
  NANDN U23167 ( .A(n22407), .B(n22406), .Z(n22408) );
  NAND U23168 ( .A(n22409), .B(n22408), .Z(n22428) );
  XNOR U23169 ( .A(n22427), .B(n22428), .Z(n22429) );
  NANDN U23170 ( .A(n22411), .B(n22410), .Z(n22415) );
  NAND U23171 ( .A(n22413), .B(n22412), .Z(n22414) );
  NAND U23172 ( .A(n22415), .B(n22414), .Z(n22430) );
  XNOR U23173 ( .A(n22429), .B(n22430), .Z(n22421) );
  XNOR U23174 ( .A(n22422), .B(n22421), .Z(n22423) );
  XNOR U23175 ( .A(n22424), .B(n22423), .Z(n22565) );
  XNOR U23176 ( .A(sreg[389]), .B(n22565), .Z(n22567) );
  NANDN U23177 ( .A(sreg[388]), .B(n22416), .Z(n22420) );
  NAND U23178 ( .A(n22418), .B(n22417), .Z(n22419) );
  NAND U23179 ( .A(n22420), .B(n22419), .Z(n22566) );
  XNOR U23180 ( .A(n22567), .B(n22566), .Z(c[389]) );
  NANDN U23181 ( .A(n22422), .B(n22421), .Z(n22426) );
  NANDN U23182 ( .A(n22424), .B(n22423), .Z(n22425) );
  AND U23183 ( .A(n22426), .B(n22425), .Z(n22573) );
  NANDN U23184 ( .A(n22428), .B(n22427), .Z(n22432) );
  NANDN U23185 ( .A(n22430), .B(n22429), .Z(n22431) );
  AND U23186 ( .A(n22432), .B(n22431), .Z(n22571) );
  NANDN U23187 ( .A(n22434), .B(n22433), .Z(n22438) );
  NANDN U23188 ( .A(n22436), .B(n22435), .Z(n22437) );
  AND U23189 ( .A(n22438), .B(n22437), .Z(n22579) );
  NANDN U23190 ( .A(n22440), .B(n22439), .Z(n22444) );
  NANDN U23191 ( .A(n22442), .B(n22441), .Z(n22443) );
  AND U23192 ( .A(n22444), .B(n22443), .Z(n22583) );
  NANDN U23193 ( .A(n22446), .B(n22445), .Z(n22450) );
  NAND U23194 ( .A(n22448), .B(n22447), .Z(n22449) );
  AND U23195 ( .A(n22450), .B(n22449), .Z(n22582) );
  XNOR U23196 ( .A(n22583), .B(n22582), .Z(n22585) );
  NANDN U23197 ( .A(n22452), .B(n22451), .Z(n22456) );
  NANDN U23198 ( .A(n22454), .B(n22453), .Z(n22455) );
  AND U23199 ( .A(n22456), .B(n22455), .Z(n22662) );
  NAND U23200 ( .A(n38385), .B(n22457), .Z(n22459) );
  XOR U23201 ( .A(b[27]), .B(a[140]), .Z(n22606) );
  NAND U23202 ( .A(n38343), .B(n22606), .Z(n22458) );
  AND U23203 ( .A(n22459), .B(n22458), .Z(n22669) );
  NAND U23204 ( .A(n183), .B(n22460), .Z(n22462) );
  XOR U23205 ( .A(b[5]), .B(a[162]), .Z(n22609) );
  NAND U23206 ( .A(n36296), .B(n22609), .Z(n22461) );
  AND U23207 ( .A(n22462), .B(n22461), .Z(n22667) );
  NAND U23208 ( .A(n190), .B(n22463), .Z(n22465) );
  XOR U23209 ( .A(b[19]), .B(a[148]), .Z(n22612) );
  NAND U23210 ( .A(n37821), .B(n22612), .Z(n22464) );
  NAND U23211 ( .A(n22465), .B(n22464), .Z(n22666) );
  XNOR U23212 ( .A(n22667), .B(n22666), .Z(n22668) );
  XNOR U23213 ( .A(n22669), .B(n22668), .Z(n22660) );
  NAND U23214 ( .A(n38470), .B(n22466), .Z(n22468) );
  XOR U23215 ( .A(b[31]), .B(a[136]), .Z(n22615) );
  NAND U23216 ( .A(n38453), .B(n22615), .Z(n22467) );
  AND U23217 ( .A(n22468), .B(n22467), .Z(n22627) );
  NAND U23218 ( .A(n181), .B(n22469), .Z(n22471) );
  XOR U23219 ( .A(b[3]), .B(a[164]), .Z(n22618) );
  NAND U23220 ( .A(n182), .B(n22618), .Z(n22470) );
  AND U23221 ( .A(n22471), .B(n22470), .Z(n22625) );
  NAND U23222 ( .A(n189), .B(n22472), .Z(n22474) );
  XOR U23223 ( .A(b[17]), .B(a[150]), .Z(n22621) );
  NAND U23224 ( .A(n37652), .B(n22621), .Z(n22473) );
  NAND U23225 ( .A(n22474), .B(n22473), .Z(n22624) );
  XNOR U23226 ( .A(n22625), .B(n22624), .Z(n22626) );
  XOR U23227 ( .A(n22627), .B(n22626), .Z(n22661) );
  XOR U23228 ( .A(n22660), .B(n22661), .Z(n22663) );
  XOR U23229 ( .A(n22662), .B(n22663), .Z(n22595) );
  NANDN U23230 ( .A(n22476), .B(n22475), .Z(n22480) );
  NANDN U23231 ( .A(n22478), .B(n22477), .Z(n22479) );
  AND U23232 ( .A(n22480), .B(n22479), .Z(n22648) );
  NANDN U23233 ( .A(n22482), .B(n22481), .Z(n22486) );
  NANDN U23234 ( .A(n22484), .B(n22483), .Z(n22485) );
  NAND U23235 ( .A(n22486), .B(n22485), .Z(n22649) );
  XNOR U23236 ( .A(n22648), .B(n22649), .Z(n22650) );
  NANDN U23237 ( .A(n22488), .B(n22487), .Z(n22492) );
  NANDN U23238 ( .A(n22490), .B(n22489), .Z(n22491) );
  NAND U23239 ( .A(n22492), .B(n22491), .Z(n22651) );
  XNOR U23240 ( .A(n22650), .B(n22651), .Z(n22594) );
  XNOR U23241 ( .A(n22595), .B(n22594), .Z(n22597) );
  NANDN U23242 ( .A(n22494), .B(n22493), .Z(n22498) );
  NANDN U23243 ( .A(n22496), .B(n22495), .Z(n22497) );
  AND U23244 ( .A(n22498), .B(n22497), .Z(n22596) );
  XOR U23245 ( .A(n22597), .B(n22596), .Z(n22711) );
  NANDN U23246 ( .A(n22500), .B(n22499), .Z(n22504) );
  NANDN U23247 ( .A(n22502), .B(n22501), .Z(n22503) );
  AND U23248 ( .A(n22504), .B(n22503), .Z(n22708) );
  NANDN U23249 ( .A(n22506), .B(n22505), .Z(n22510) );
  NANDN U23250 ( .A(n22508), .B(n22507), .Z(n22509) );
  AND U23251 ( .A(n22510), .B(n22509), .Z(n22591) );
  NANDN U23252 ( .A(n22512), .B(n22511), .Z(n22516) );
  OR U23253 ( .A(n22514), .B(n22513), .Z(n22515) );
  AND U23254 ( .A(n22516), .B(n22515), .Z(n22589) );
  NANDN U23255 ( .A(n22518), .B(n22517), .Z(n22522) );
  NANDN U23256 ( .A(n22520), .B(n22519), .Z(n22521) );
  AND U23257 ( .A(n22522), .B(n22521), .Z(n22655) );
  NANDN U23258 ( .A(n22524), .B(n22523), .Z(n22528) );
  NANDN U23259 ( .A(n22526), .B(n22525), .Z(n22527) );
  NAND U23260 ( .A(n22528), .B(n22527), .Z(n22654) );
  XNOR U23261 ( .A(n22655), .B(n22654), .Z(n22656) );
  NAND U23262 ( .A(b[0]), .B(a[166]), .Z(n22529) );
  XNOR U23263 ( .A(b[1]), .B(n22529), .Z(n22531) );
  NANDN U23264 ( .A(b[0]), .B(a[165]), .Z(n22530) );
  NAND U23265 ( .A(n22531), .B(n22530), .Z(n22603) );
  NAND U23266 ( .A(n194), .B(n22532), .Z(n22534) );
  XOR U23267 ( .A(b[29]), .B(a[138]), .Z(n22681) );
  NAND U23268 ( .A(n38456), .B(n22681), .Z(n22533) );
  AND U23269 ( .A(n22534), .B(n22533), .Z(n22601) );
  AND U23270 ( .A(b[31]), .B(a[134]), .Z(n22600) );
  XNOR U23271 ( .A(n22601), .B(n22600), .Z(n22602) );
  XNOR U23272 ( .A(n22603), .B(n22602), .Z(n22642) );
  NAND U23273 ( .A(n38185), .B(n22535), .Z(n22537) );
  XOR U23274 ( .A(b[23]), .B(a[144]), .Z(n22684) );
  NAND U23275 ( .A(n38132), .B(n22684), .Z(n22536) );
  AND U23276 ( .A(n22537), .B(n22536), .Z(n22675) );
  NAND U23277 ( .A(n184), .B(n22538), .Z(n22540) );
  XOR U23278 ( .A(b[7]), .B(a[160]), .Z(n22687) );
  NAND U23279 ( .A(n36592), .B(n22687), .Z(n22539) );
  AND U23280 ( .A(n22540), .B(n22539), .Z(n22673) );
  NAND U23281 ( .A(n38289), .B(n22541), .Z(n22543) );
  XOR U23282 ( .A(b[25]), .B(a[142]), .Z(n22690) );
  NAND U23283 ( .A(n38247), .B(n22690), .Z(n22542) );
  NAND U23284 ( .A(n22543), .B(n22542), .Z(n22672) );
  XNOR U23285 ( .A(n22673), .B(n22672), .Z(n22674) );
  XOR U23286 ( .A(n22675), .B(n22674), .Z(n22643) );
  XNOR U23287 ( .A(n22642), .B(n22643), .Z(n22644) );
  NAND U23288 ( .A(n187), .B(n22544), .Z(n22546) );
  XOR U23289 ( .A(b[13]), .B(a[154]), .Z(n22693) );
  NAND U23290 ( .A(n37295), .B(n22693), .Z(n22545) );
  AND U23291 ( .A(n22546), .B(n22545), .Z(n22637) );
  NAND U23292 ( .A(n186), .B(n22547), .Z(n22549) );
  XOR U23293 ( .A(b[11]), .B(a[156]), .Z(n22696) );
  NAND U23294 ( .A(n37097), .B(n22696), .Z(n22548) );
  NAND U23295 ( .A(n22549), .B(n22548), .Z(n22636) );
  XNOR U23296 ( .A(n22637), .B(n22636), .Z(n22638) );
  NAND U23297 ( .A(n188), .B(n22550), .Z(n22552) );
  XOR U23298 ( .A(b[15]), .B(a[152]), .Z(n22699) );
  NAND U23299 ( .A(n37382), .B(n22699), .Z(n22551) );
  AND U23300 ( .A(n22552), .B(n22551), .Z(n22633) );
  NAND U23301 ( .A(n38064), .B(n22553), .Z(n22555) );
  XOR U23302 ( .A(b[21]), .B(a[146]), .Z(n22702) );
  NAND U23303 ( .A(n37993), .B(n22702), .Z(n22554) );
  AND U23304 ( .A(n22555), .B(n22554), .Z(n22631) );
  NAND U23305 ( .A(n185), .B(n22556), .Z(n22558) );
  XOR U23306 ( .A(b[9]), .B(a[158]), .Z(n22705) );
  NAND U23307 ( .A(n36805), .B(n22705), .Z(n22557) );
  NAND U23308 ( .A(n22558), .B(n22557), .Z(n22630) );
  XNOR U23309 ( .A(n22631), .B(n22630), .Z(n22632) );
  XOR U23310 ( .A(n22633), .B(n22632), .Z(n22639) );
  XOR U23311 ( .A(n22638), .B(n22639), .Z(n22645) );
  XOR U23312 ( .A(n22644), .B(n22645), .Z(n22657) );
  XNOR U23313 ( .A(n22656), .B(n22657), .Z(n22588) );
  XNOR U23314 ( .A(n22589), .B(n22588), .Z(n22590) );
  XOR U23315 ( .A(n22591), .B(n22590), .Z(n22709) );
  XNOR U23316 ( .A(n22708), .B(n22709), .Z(n22710) );
  XNOR U23317 ( .A(n22711), .B(n22710), .Z(n22584) );
  XOR U23318 ( .A(n22585), .B(n22584), .Z(n22577) );
  NANDN U23319 ( .A(n22560), .B(n22559), .Z(n22564) );
  OR U23320 ( .A(n22562), .B(n22561), .Z(n22563) );
  AND U23321 ( .A(n22564), .B(n22563), .Z(n22576) );
  XNOR U23322 ( .A(n22577), .B(n22576), .Z(n22578) );
  XNOR U23323 ( .A(n22579), .B(n22578), .Z(n22570) );
  XNOR U23324 ( .A(n22571), .B(n22570), .Z(n22572) );
  XNOR U23325 ( .A(n22573), .B(n22572), .Z(n22714) );
  XNOR U23326 ( .A(sreg[390]), .B(n22714), .Z(n22716) );
  NANDN U23327 ( .A(sreg[389]), .B(n22565), .Z(n22569) );
  NAND U23328 ( .A(n22567), .B(n22566), .Z(n22568) );
  NAND U23329 ( .A(n22569), .B(n22568), .Z(n22715) );
  XNOR U23330 ( .A(n22716), .B(n22715), .Z(c[390]) );
  NANDN U23331 ( .A(n22571), .B(n22570), .Z(n22575) );
  NANDN U23332 ( .A(n22573), .B(n22572), .Z(n22574) );
  AND U23333 ( .A(n22575), .B(n22574), .Z(n22722) );
  NANDN U23334 ( .A(n22577), .B(n22576), .Z(n22581) );
  NANDN U23335 ( .A(n22579), .B(n22578), .Z(n22580) );
  AND U23336 ( .A(n22581), .B(n22580), .Z(n22720) );
  NANDN U23337 ( .A(n22583), .B(n22582), .Z(n22587) );
  NAND U23338 ( .A(n22585), .B(n22584), .Z(n22586) );
  AND U23339 ( .A(n22587), .B(n22586), .Z(n22727) );
  NANDN U23340 ( .A(n22589), .B(n22588), .Z(n22593) );
  NANDN U23341 ( .A(n22591), .B(n22590), .Z(n22592) );
  AND U23342 ( .A(n22593), .B(n22592), .Z(n22732) );
  NANDN U23343 ( .A(n22595), .B(n22594), .Z(n22599) );
  NAND U23344 ( .A(n22597), .B(n22596), .Z(n22598) );
  AND U23345 ( .A(n22599), .B(n22598), .Z(n22731) );
  XNOR U23346 ( .A(n22732), .B(n22731), .Z(n22734) );
  NANDN U23347 ( .A(n22601), .B(n22600), .Z(n22605) );
  NANDN U23348 ( .A(n22603), .B(n22602), .Z(n22604) );
  AND U23349 ( .A(n22605), .B(n22604), .Z(n22811) );
  NAND U23350 ( .A(n38385), .B(n22606), .Z(n22608) );
  XOR U23351 ( .A(b[27]), .B(a[141]), .Z(n22755) );
  NAND U23352 ( .A(n38343), .B(n22755), .Z(n22607) );
  AND U23353 ( .A(n22608), .B(n22607), .Z(n22818) );
  NAND U23354 ( .A(n183), .B(n22609), .Z(n22611) );
  XOR U23355 ( .A(b[5]), .B(a[163]), .Z(n22758) );
  NAND U23356 ( .A(n36296), .B(n22758), .Z(n22610) );
  AND U23357 ( .A(n22611), .B(n22610), .Z(n22816) );
  NAND U23358 ( .A(n190), .B(n22612), .Z(n22614) );
  XOR U23359 ( .A(b[19]), .B(a[149]), .Z(n22761) );
  NAND U23360 ( .A(n37821), .B(n22761), .Z(n22613) );
  NAND U23361 ( .A(n22614), .B(n22613), .Z(n22815) );
  XNOR U23362 ( .A(n22816), .B(n22815), .Z(n22817) );
  XNOR U23363 ( .A(n22818), .B(n22817), .Z(n22809) );
  NAND U23364 ( .A(n38470), .B(n22615), .Z(n22617) );
  XOR U23365 ( .A(b[31]), .B(a[137]), .Z(n22764) );
  NAND U23366 ( .A(n38453), .B(n22764), .Z(n22616) );
  AND U23367 ( .A(n22617), .B(n22616), .Z(n22776) );
  NAND U23368 ( .A(n181), .B(n22618), .Z(n22620) );
  XOR U23369 ( .A(b[3]), .B(a[165]), .Z(n22767) );
  NAND U23370 ( .A(n182), .B(n22767), .Z(n22619) );
  AND U23371 ( .A(n22620), .B(n22619), .Z(n22774) );
  NAND U23372 ( .A(n189), .B(n22621), .Z(n22623) );
  XOR U23373 ( .A(b[17]), .B(a[151]), .Z(n22770) );
  NAND U23374 ( .A(n37652), .B(n22770), .Z(n22622) );
  NAND U23375 ( .A(n22623), .B(n22622), .Z(n22773) );
  XNOR U23376 ( .A(n22774), .B(n22773), .Z(n22775) );
  XOR U23377 ( .A(n22776), .B(n22775), .Z(n22810) );
  XOR U23378 ( .A(n22809), .B(n22810), .Z(n22812) );
  XOR U23379 ( .A(n22811), .B(n22812), .Z(n22744) );
  NANDN U23380 ( .A(n22625), .B(n22624), .Z(n22629) );
  NANDN U23381 ( .A(n22627), .B(n22626), .Z(n22628) );
  AND U23382 ( .A(n22629), .B(n22628), .Z(n22797) );
  NANDN U23383 ( .A(n22631), .B(n22630), .Z(n22635) );
  NANDN U23384 ( .A(n22633), .B(n22632), .Z(n22634) );
  NAND U23385 ( .A(n22635), .B(n22634), .Z(n22798) );
  XNOR U23386 ( .A(n22797), .B(n22798), .Z(n22799) );
  NANDN U23387 ( .A(n22637), .B(n22636), .Z(n22641) );
  NANDN U23388 ( .A(n22639), .B(n22638), .Z(n22640) );
  NAND U23389 ( .A(n22641), .B(n22640), .Z(n22800) );
  XNOR U23390 ( .A(n22799), .B(n22800), .Z(n22743) );
  XNOR U23391 ( .A(n22744), .B(n22743), .Z(n22746) );
  NANDN U23392 ( .A(n22643), .B(n22642), .Z(n22647) );
  NANDN U23393 ( .A(n22645), .B(n22644), .Z(n22646) );
  AND U23394 ( .A(n22647), .B(n22646), .Z(n22745) );
  XOR U23395 ( .A(n22746), .B(n22745), .Z(n22860) );
  NANDN U23396 ( .A(n22649), .B(n22648), .Z(n22653) );
  NANDN U23397 ( .A(n22651), .B(n22650), .Z(n22652) );
  AND U23398 ( .A(n22653), .B(n22652), .Z(n22857) );
  NANDN U23399 ( .A(n22655), .B(n22654), .Z(n22659) );
  NANDN U23400 ( .A(n22657), .B(n22656), .Z(n22658) );
  AND U23401 ( .A(n22659), .B(n22658), .Z(n22740) );
  NANDN U23402 ( .A(n22661), .B(n22660), .Z(n22665) );
  OR U23403 ( .A(n22663), .B(n22662), .Z(n22664) );
  AND U23404 ( .A(n22665), .B(n22664), .Z(n22738) );
  NANDN U23405 ( .A(n22667), .B(n22666), .Z(n22671) );
  NANDN U23406 ( .A(n22669), .B(n22668), .Z(n22670) );
  AND U23407 ( .A(n22671), .B(n22670), .Z(n22804) );
  NANDN U23408 ( .A(n22673), .B(n22672), .Z(n22677) );
  NANDN U23409 ( .A(n22675), .B(n22674), .Z(n22676) );
  NAND U23410 ( .A(n22677), .B(n22676), .Z(n22803) );
  XNOR U23411 ( .A(n22804), .B(n22803), .Z(n22805) );
  NAND U23412 ( .A(b[0]), .B(a[167]), .Z(n22678) );
  XNOR U23413 ( .A(b[1]), .B(n22678), .Z(n22680) );
  NANDN U23414 ( .A(b[0]), .B(a[166]), .Z(n22679) );
  NAND U23415 ( .A(n22680), .B(n22679), .Z(n22752) );
  NAND U23416 ( .A(n194), .B(n22681), .Z(n22683) );
  XOR U23417 ( .A(b[29]), .B(a[139]), .Z(n22830) );
  NAND U23418 ( .A(n38456), .B(n22830), .Z(n22682) );
  AND U23419 ( .A(n22683), .B(n22682), .Z(n22750) );
  AND U23420 ( .A(b[31]), .B(a[135]), .Z(n22749) );
  XNOR U23421 ( .A(n22750), .B(n22749), .Z(n22751) );
  XNOR U23422 ( .A(n22752), .B(n22751), .Z(n22791) );
  NAND U23423 ( .A(n38185), .B(n22684), .Z(n22686) );
  XOR U23424 ( .A(b[23]), .B(a[145]), .Z(n22833) );
  NAND U23425 ( .A(n38132), .B(n22833), .Z(n22685) );
  AND U23426 ( .A(n22686), .B(n22685), .Z(n22824) );
  NAND U23427 ( .A(n184), .B(n22687), .Z(n22689) );
  XOR U23428 ( .A(b[7]), .B(a[161]), .Z(n22836) );
  NAND U23429 ( .A(n36592), .B(n22836), .Z(n22688) );
  AND U23430 ( .A(n22689), .B(n22688), .Z(n22822) );
  NAND U23431 ( .A(n38289), .B(n22690), .Z(n22692) );
  XOR U23432 ( .A(b[25]), .B(a[143]), .Z(n22839) );
  NAND U23433 ( .A(n38247), .B(n22839), .Z(n22691) );
  NAND U23434 ( .A(n22692), .B(n22691), .Z(n22821) );
  XNOR U23435 ( .A(n22822), .B(n22821), .Z(n22823) );
  XOR U23436 ( .A(n22824), .B(n22823), .Z(n22792) );
  XNOR U23437 ( .A(n22791), .B(n22792), .Z(n22793) );
  NAND U23438 ( .A(n187), .B(n22693), .Z(n22695) );
  XOR U23439 ( .A(b[13]), .B(a[155]), .Z(n22842) );
  NAND U23440 ( .A(n37295), .B(n22842), .Z(n22694) );
  AND U23441 ( .A(n22695), .B(n22694), .Z(n22786) );
  NAND U23442 ( .A(n186), .B(n22696), .Z(n22698) );
  XOR U23443 ( .A(b[11]), .B(a[157]), .Z(n22845) );
  NAND U23444 ( .A(n37097), .B(n22845), .Z(n22697) );
  NAND U23445 ( .A(n22698), .B(n22697), .Z(n22785) );
  XNOR U23446 ( .A(n22786), .B(n22785), .Z(n22787) );
  NAND U23447 ( .A(n188), .B(n22699), .Z(n22701) );
  XOR U23448 ( .A(b[15]), .B(a[153]), .Z(n22848) );
  NAND U23449 ( .A(n37382), .B(n22848), .Z(n22700) );
  AND U23450 ( .A(n22701), .B(n22700), .Z(n22782) );
  NAND U23451 ( .A(n38064), .B(n22702), .Z(n22704) );
  XOR U23452 ( .A(b[21]), .B(a[147]), .Z(n22851) );
  NAND U23453 ( .A(n37993), .B(n22851), .Z(n22703) );
  AND U23454 ( .A(n22704), .B(n22703), .Z(n22780) );
  NAND U23455 ( .A(n185), .B(n22705), .Z(n22707) );
  XOR U23456 ( .A(b[9]), .B(a[159]), .Z(n22854) );
  NAND U23457 ( .A(n36805), .B(n22854), .Z(n22706) );
  NAND U23458 ( .A(n22707), .B(n22706), .Z(n22779) );
  XNOR U23459 ( .A(n22780), .B(n22779), .Z(n22781) );
  XOR U23460 ( .A(n22782), .B(n22781), .Z(n22788) );
  XOR U23461 ( .A(n22787), .B(n22788), .Z(n22794) );
  XOR U23462 ( .A(n22793), .B(n22794), .Z(n22806) );
  XNOR U23463 ( .A(n22805), .B(n22806), .Z(n22737) );
  XNOR U23464 ( .A(n22738), .B(n22737), .Z(n22739) );
  XOR U23465 ( .A(n22740), .B(n22739), .Z(n22858) );
  XNOR U23466 ( .A(n22857), .B(n22858), .Z(n22859) );
  XNOR U23467 ( .A(n22860), .B(n22859), .Z(n22733) );
  XOR U23468 ( .A(n22734), .B(n22733), .Z(n22726) );
  NANDN U23469 ( .A(n22709), .B(n22708), .Z(n22713) );
  NANDN U23470 ( .A(n22711), .B(n22710), .Z(n22712) );
  AND U23471 ( .A(n22713), .B(n22712), .Z(n22725) );
  XOR U23472 ( .A(n22726), .B(n22725), .Z(n22728) );
  XNOR U23473 ( .A(n22727), .B(n22728), .Z(n22719) );
  XNOR U23474 ( .A(n22720), .B(n22719), .Z(n22721) );
  XNOR U23475 ( .A(n22722), .B(n22721), .Z(n22863) );
  XNOR U23476 ( .A(sreg[391]), .B(n22863), .Z(n22865) );
  NANDN U23477 ( .A(sreg[390]), .B(n22714), .Z(n22718) );
  NAND U23478 ( .A(n22716), .B(n22715), .Z(n22717) );
  NAND U23479 ( .A(n22718), .B(n22717), .Z(n22864) );
  XNOR U23480 ( .A(n22865), .B(n22864), .Z(c[391]) );
  NANDN U23481 ( .A(n22720), .B(n22719), .Z(n22724) );
  NANDN U23482 ( .A(n22722), .B(n22721), .Z(n22723) );
  AND U23483 ( .A(n22724), .B(n22723), .Z(n22871) );
  NANDN U23484 ( .A(n22726), .B(n22725), .Z(n22730) );
  NANDN U23485 ( .A(n22728), .B(n22727), .Z(n22729) );
  AND U23486 ( .A(n22730), .B(n22729), .Z(n22869) );
  NANDN U23487 ( .A(n22732), .B(n22731), .Z(n22736) );
  NAND U23488 ( .A(n22734), .B(n22733), .Z(n22735) );
  AND U23489 ( .A(n22736), .B(n22735), .Z(n22876) );
  NANDN U23490 ( .A(n22738), .B(n22737), .Z(n22742) );
  NANDN U23491 ( .A(n22740), .B(n22739), .Z(n22741) );
  AND U23492 ( .A(n22742), .B(n22741), .Z(n22881) );
  NANDN U23493 ( .A(n22744), .B(n22743), .Z(n22748) );
  NAND U23494 ( .A(n22746), .B(n22745), .Z(n22747) );
  AND U23495 ( .A(n22748), .B(n22747), .Z(n22880) );
  XNOR U23496 ( .A(n22881), .B(n22880), .Z(n22883) );
  NANDN U23497 ( .A(n22750), .B(n22749), .Z(n22754) );
  NANDN U23498 ( .A(n22752), .B(n22751), .Z(n22753) );
  AND U23499 ( .A(n22754), .B(n22753), .Z(n22960) );
  NAND U23500 ( .A(n38385), .B(n22755), .Z(n22757) );
  XOR U23501 ( .A(b[27]), .B(a[142]), .Z(n22904) );
  NAND U23502 ( .A(n38343), .B(n22904), .Z(n22756) );
  AND U23503 ( .A(n22757), .B(n22756), .Z(n22967) );
  NAND U23504 ( .A(n183), .B(n22758), .Z(n22760) );
  XOR U23505 ( .A(b[5]), .B(a[164]), .Z(n22907) );
  NAND U23506 ( .A(n36296), .B(n22907), .Z(n22759) );
  AND U23507 ( .A(n22760), .B(n22759), .Z(n22965) );
  NAND U23508 ( .A(n190), .B(n22761), .Z(n22763) );
  XOR U23509 ( .A(b[19]), .B(a[150]), .Z(n22910) );
  NAND U23510 ( .A(n37821), .B(n22910), .Z(n22762) );
  NAND U23511 ( .A(n22763), .B(n22762), .Z(n22964) );
  XNOR U23512 ( .A(n22965), .B(n22964), .Z(n22966) );
  XNOR U23513 ( .A(n22967), .B(n22966), .Z(n22958) );
  NAND U23514 ( .A(n38470), .B(n22764), .Z(n22766) );
  XOR U23515 ( .A(b[31]), .B(a[138]), .Z(n22913) );
  NAND U23516 ( .A(n38453), .B(n22913), .Z(n22765) );
  AND U23517 ( .A(n22766), .B(n22765), .Z(n22925) );
  NAND U23518 ( .A(n181), .B(n22767), .Z(n22769) );
  XOR U23519 ( .A(b[3]), .B(a[166]), .Z(n22916) );
  NAND U23520 ( .A(n182), .B(n22916), .Z(n22768) );
  AND U23521 ( .A(n22769), .B(n22768), .Z(n22923) );
  NAND U23522 ( .A(n189), .B(n22770), .Z(n22772) );
  XOR U23523 ( .A(b[17]), .B(a[152]), .Z(n22919) );
  NAND U23524 ( .A(n37652), .B(n22919), .Z(n22771) );
  NAND U23525 ( .A(n22772), .B(n22771), .Z(n22922) );
  XNOR U23526 ( .A(n22923), .B(n22922), .Z(n22924) );
  XOR U23527 ( .A(n22925), .B(n22924), .Z(n22959) );
  XOR U23528 ( .A(n22958), .B(n22959), .Z(n22961) );
  XOR U23529 ( .A(n22960), .B(n22961), .Z(n22893) );
  NANDN U23530 ( .A(n22774), .B(n22773), .Z(n22778) );
  NANDN U23531 ( .A(n22776), .B(n22775), .Z(n22777) );
  AND U23532 ( .A(n22778), .B(n22777), .Z(n22946) );
  NANDN U23533 ( .A(n22780), .B(n22779), .Z(n22784) );
  NANDN U23534 ( .A(n22782), .B(n22781), .Z(n22783) );
  NAND U23535 ( .A(n22784), .B(n22783), .Z(n22947) );
  XNOR U23536 ( .A(n22946), .B(n22947), .Z(n22948) );
  NANDN U23537 ( .A(n22786), .B(n22785), .Z(n22790) );
  NANDN U23538 ( .A(n22788), .B(n22787), .Z(n22789) );
  NAND U23539 ( .A(n22790), .B(n22789), .Z(n22949) );
  XNOR U23540 ( .A(n22948), .B(n22949), .Z(n22892) );
  XNOR U23541 ( .A(n22893), .B(n22892), .Z(n22895) );
  NANDN U23542 ( .A(n22792), .B(n22791), .Z(n22796) );
  NANDN U23543 ( .A(n22794), .B(n22793), .Z(n22795) );
  AND U23544 ( .A(n22796), .B(n22795), .Z(n22894) );
  XOR U23545 ( .A(n22895), .B(n22894), .Z(n23009) );
  NANDN U23546 ( .A(n22798), .B(n22797), .Z(n22802) );
  NANDN U23547 ( .A(n22800), .B(n22799), .Z(n22801) );
  AND U23548 ( .A(n22802), .B(n22801), .Z(n23006) );
  NANDN U23549 ( .A(n22804), .B(n22803), .Z(n22808) );
  NANDN U23550 ( .A(n22806), .B(n22805), .Z(n22807) );
  AND U23551 ( .A(n22808), .B(n22807), .Z(n22889) );
  NANDN U23552 ( .A(n22810), .B(n22809), .Z(n22814) );
  OR U23553 ( .A(n22812), .B(n22811), .Z(n22813) );
  AND U23554 ( .A(n22814), .B(n22813), .Z(n22887) );
  NANDN U23555 ( .A(n22816), .B(n22815), .Z(n22820) );
  NANDN U23556 ( .A(n22818), .B(n22817), .Z(n22819) );
  AND U23557 ( .A(n22820), .B(n22819), .Z(n22953) );
  NANDN U23558 ( .A(n22822), .B(n22821), .Z(n22826) );
  NANDN U23559 ( .A(n22824), .B(n22823), .Z(n22825) );
  NAND U23560 ( .A(n22826), .B(n22825), .Z(n22952) );
  XNOR U23561 ( .A(n22953), .B(n22952), .Z(n22954) );
  NAND U23562 ( .A(b[0]), .B(a[168]), .Z(n22827) );
  XNOR U23563 ( .A(b[1]), .B(n22827), .Z(n22829) );
  NANDN U23564 ( .A(b[0]), .B(a[167]), .Z(n22828) );
  NAND U23565 ( .A(n22829), .B(n22828), .Z(n22901) );
  NAND U23566 ( .A(n194), .B(n22830), .Z(n22832) );
  XOR U23567 ( .A(b[29]), .B(a[140]), .Z(n22976) );
  NAND U23568 ( .A(n38456), .B(n22976), .Z(n22831) );
  AND U23569 ( .A(n22832), .B(n22831), .Z(n22899) );
  AND U23570 ( .A(b[31]), .B(a[136]), .Z(n22898) );
  XNOR U23571 ( .A(n22899), .B(n22898), .Z(n22900) );
  XNOR U23572 ( .A(n22901), .B(n22900), .Z(n22940) );
  NAND U23573 ( .A(n38185), .B(n22833), .Z(n22835) );
  XOR U23574 ( .A(b[23]), .B(a[146]), .Z(n22982) );
  NAND U23575 ( .A(n38132), .B(n22982), .Z(n22834) );
  AND U23576 ( .A(n22835), .B(n22834), .Z(n22973) );
  NAND U23577 ( .A(n184), .B(n22836), .Z(n22838) );
  XOR U23578 ( .A(b[7]), .B(a[162]), .Z(n22985) );
  NAND U23579 ( .A(n36592), .B(n22985), .Z(n22837) );
  AND U23580 ( .A(n22838), .B(n22837), .Z(n22971) );
  NAND U23581 ( .A(n38289), .B(n22839), .Z(n22841) );
  XOR U23582 ( .A(b[25]), .B(a[144]), .Z(n22988) );
  NAND U23583 ( .A(n38247), .B(n22988), .Z(n22840) );
  NAND U23584 ( .A(n22841), .B(n22840), .Z(n22970) );
  XNOR U23585 ( .A(n22971), .B(n22970), .Z(n22972) );
  XOR U23586 ( .A(n22973), .B(n22972), .Z(n22941) );
  XNOR U23587 ( .A(n22940), .B(n22941), .Z(n22942) );
  NAND U23588 ( .A(n187), .B(n22842), .Z(n22844) );
  XOR U23589 ( .A(b[13]), .B(a[156]), .Z(n22991) );
  NAND U23590 ( .A(n37295), .B(n22991), .Z(n22843) );
  AND U23591 ( .A(n22844), .B(n22843), .Z(n22935) );
  NAND U23592 ( .A(n186), .B(n22845), .Z(n22847) );
  XOR U23593 ( .A(b[11]), .B(a[158]), .Z(n22994) );
  NAND U23594 ( .A(n37097), .B(n22994), .Z(n22846) );
  NAND U23595 ( .A(n22847), .B(n22846), .Z(n22934) );
  XNOR U23596 ( .A(n22935), .B(n22934), .Z(n22936) );
  NAND U23597 ( .A(n188), .B(n22848), .Z(n22850) );
  XOR U23598 ( .A(b[15]), .B(a[154]), .Z(n22997) );
  NAND U23599 ( .A(n37382), .B(n22997), .Z(n22849) );
  AND U23600 ( .A(n22850), .B(n22849), .Z(n22931) );
  NAND U23601 ( .A(n38064), .B(n22851), .Z(n22853) );
  XOR U23602 ( .A(b[21]), .B(a[148]), .Z(n23000) );
  NAND U23603 ( .A(n37993), .B(n23000), .Z(n22852) );
  AND U23604 ( .A(n22853), .B(n22852), .Z(n22929) );
  NAND U23605 ( .A(n185), .B(n22854), .Z(n22856) );
  XOR U23606 ( .A(b[9]), .B(a[160]), .Z(n23003) );
  NAND U23607 ( .A(n36805), .B(n23003), .Z(n22855) );
  NAND U23608 ( .A(n22856), .B(n22855), .Z(n22928) );
  XNOR U23609 ( .A(n22929), .B(n22928), .Z(n22930) );
  XOR U23610 ( .A(n22931), .B(n22930), .Z(n22937) );
  XOR U23611 ( .A(n22936), .B(n22937), .Z(n22943) );
  XOR U23612 ( .A(n22942), .B(n22943), .Z(n22955) );
  XNOR U23613 ( .A(n22954), .B(n22955), .Z(n22886) );
  XNOR U23614 ( .A(n22887), .B(n22886), .Z(n22888) );
  XOR U23615 ( .A(n22889), .B(n22888), .Z(n23007) );
  XNOR U23616 ( .A(n23006), .B(n23007), .Z(n23008) );
  XNOR U23617 ( .A(n23009), .B(n23008), .Z(n22882) );
  XOR U23618 ( .A(n22883), .B(n22882), .Z(n22875) );
  NANDN U23619 ( .A(n22858), .B(n22857), .Z(n22862) );
  NANDN U23620 ( .A(n22860), .B(n22859), .Z(n22861) );
  AND U23621 ( .A(n22862), .B(n22861), .Z(n22874) );
  XOR U23622 ( .A(n22875), .B(n22874), .Z(n22877) );
  XNOR U23623 ( .A(n22876), .B(n22877), .Z(n22868) );
  XNOR U23624 ( .A(n22869), .B(n22868), .Z(n22870) );
  XNOR U23625 ( .A(n22871), .B(n22870), .Z(n23012) );
  XNOR U23626 ( .A(sreg[392]), .B(n23012), .Z(n23014) );
  NANDN U23627 ( .A(sreg[391]), .B(n22863), .Z(n22867) );
  NAND U23628 ( .A(n22865), .B(n22864), .Z(n22866) );
  NAND U23629 ( .A(n22867), .B(n22866), .Z(n23013) );
  XNOR U23630 ( .A(n23014), .B(n23013), .Z(c[392]) );
  NANDN U23631 ( .A(n22869), .B(n22868), .Z(n22873) );
  NANDN U23632 ( .A(n22871), .B(n22870), .Z(n22872) );
  AND U23633 ( .A(n22873), .B(n22872), .Z(n23020) );
  NANDN U23634 ( .A(n22875), .B(n22874), .Z(n22879) );
  NANDN U23635 ( .A(n22877), .B(n22876), .Z(n22878) );
  AND U23636 ( .A(n22879), .B(n22878), .Z(n23018) );
  NANDN U23637 ( .A(n22881), .B(n22880), .Z(n22885) );
  NAND U23638 ( .A(n22883), .B(n22882), .Z(n22884) );
  AND U23639 ( .A(n22885), .B(n22884), .Z(n23025) );
  NANDN U23640 ( .A(n22887), .B(n22886), .Z(n22891) );
  NANDN U23641 ( .A(n22889), .B(n22888), .Z(n22890) );
  AND U23642 ( .A(n22891), .B(n22890), .Z(n23030) );
  NANDN U23643 ( .A(n22893), .B(n22892), .Z(n22897) );
  NAND U23644 ( .A(n22895), .B(n22894), .Z(n22896) );
  AND U23645 ( .A(n22897), .B(n22896), .Z(n23029) );
  XNOR U23646 ( .A(n23030), .B(n23029), .Z(n23032) );
  NANDN U23647 ( .A(n22899), .B(n22898), .Z(n22903) );
  NANDN U23648 ( .A(n22901), .B(n22900), .Z(n22902) );
  AND U23649 ( .A(n22903), .B(n22902), .Z(n23109) );
  NAND U23650 ( .A(n38385), .B(n22904), .Z(n22906) );
  XOR U23651 ( .A(b[27]), .B(a[143]), .Z(n23053) );
  NAND U23652 ( .A(n38343), .B(n23053), .Z(n22905) );
  AND U23653 ( .A(n22906), .B(n22905), .Z(n23116) );
  NAND U23654 ( .A(n183), .B(n22907), .Z(n22909) );
  XOR U23655 ( .A(b[5]), .B(a[165]), .Z(n23056) );
  NAND U23656 ( .A(n36296), .B(n23056), .Z(n22908) );
  AND U23657 ( .A(n22909), .B(n22908), .Z(n23114) );
  NAND U23658 ( .A(n190), .B(n22910), .Z(n22912) );
  XOR U23659 ( .A(b[19]), .B(a[151]), .Z(n23059) );
  NAND U23660 ( .A(n37821), .B(n23059), .Z(n22911) );
  NAND U23661 ( .A(n22912), .B(n22911), .Z(n23113) );
  XNOR U23662 ( .A(n23114), .B(n23113), .Z(n23115) );
  XNOR U23663 ( .A(n23116), .B(n23115), .Z(n23107) );
  NAND U23664 ( .A(n38470), .B(n22913), .Z(n22915) );
  XOR U23665 ( .A(b[31]), .B(a[139]), .Z(n23062) );
  NAND U23666 ( .A(n38453), .B(n23062), .Z(n22914) );
  AND U23667 ( .A(n22915), .B(n22914), .Z(n23074) );
  NAND U23668 ( .A(n181), .B(n22916), .Z(n22918) );
  XOR U23669 ( .A(b[3]), .B(a[167]), .Z(n23065) );
  NAND U23670 ( .A(n182), .B(n23065), .Z(n22917) );
  AND U23671 ( .A(n22918), .B(n22917), .Z(n23072) );
  NAND U23672 ( .A(n189), .B(n22919), .Z(n22921) );
  XOR U23673 ( .A(b[17]), .B(a[153]), .Z(n23068) );
  NAND U23674 ( .A(n37652), .B(n23068), .Z(n22920) );
  NAND U23675 ( .A(n22921), .B(n22920), .Z(n23071) );
  XNOR U23676 ( .A(n23072), .B(n23071), .Z(n23073) );
  XOR U23677 ( .A(n23074), .B(n23073), .Z(n23108) );
  XOR U23678 ( .A(n23107), .B(n23108), .Z(n23110) );
  XOR U23679 ( .A(n23109), .B(n23110), .Z(n23042) );
  NANDN U23680 ( .A(n22923), .B(n22922), .Z(n22927) );
  NANDN U23681 ( .A(n22925), .B(n22924), .Z(n22926) );
  AND U23682 ( .A(n22927), .B(n22926), .Z(n23095) );
  NANDN U23683 ( .A(n22929), .B(n22928), .Z(n22933) );
  NANDN U23684 ( .A(n22931), .B(n22930), .Z(n22932) );
  NAND U23685 ( .A(n22933), .B(n22932), .Z(n23096) );
  XNOR U23686 ( .A(n23095), .B(n23096), .Z(n23097) );
  NANDN U23687 ( .A(n22935), .B(n22934), .Z(n22939) );
  NANDN U23688 ( .A(n22937), .B(n22936), .Z(n22938) );
  NAND U23689 ( .A(n22939), .B(n22938), .Z(n23098) );
  XNOR U23690 ( .A(n23097), .B(n23098), .Z(n23041) );
  XNOR U23691 ( .A(n23042), .B(n23041), .Z(n23044) );
  NANDN U23692 ( .A(n22941), .B(n22940), .Z(n22945) );
  NANDN U23693 ( .A(n22943), .B(n22942), .Z(n22944) );
  AND U23694 ( .A(n22945), .B(n22944), .Z(n23043) );
  XOR U23695 ( .A(n23044), .B(n23043), .Z(n23158) );
  NANDN U23696 ( .A(n22947), .B(n22946), .Z(n22951) );
  NANDN U23697 ( .A(n22949), .B(n22948), .Z(n22950) );
  AND U23698 ( .A(n22951), .B(n22950), .Z(n23155) );
  NANDN U23699 ( .A(n22953), .B(n22952), .Z(n22957) );
  NANDN U23700 ( .A(n22955), .B(n22954), .Z(n22956) );
  AND U23701 ( .A(n22957), .B(n22956), .Z(n23038) );
  NANDN U23702 ( .A(n22959), .B(n22958), .Z(n22963) );
  OR U23703 ( .A(n22961), .B(n22960), .Z(n22962) );
  AND U23704 ( .A(n22963), .B(n22962), .Z(n23036) );
  NANDN U23705 ( .A(n22965), .B(n22964), .Z(n22969) );
  NANDN U23706 ( .A(n22967), .B(n22966), .Z(n22968) );
  AND U23707 ( .A(n22969), .B(n22968), .Z(n23102) );
  NANDN U23708 ( .A(n22971), .B(n22970), .Z(n22975) );
  NANDN U23709 ( .A(n22973), .B(n22972), .Z(n22974) );
  NAND U23710 ( .A(n22975), .B(n22974), .Z(n23101) );
  XNOR U23711 ( .A(n23102), .B(n23101), .Z(n23103) );
  NAND U23712 ( .A(n194), .B(n22976), .Z(n22978) );
  XOR U23713 ( .A(b[29]), .B(a[141]), .Z(n23128) );
  NAND U23714 ( .A(n38456), .B(n23128), .Z(n22977) );
  AND U23715 ( .A(n22978), .B(n22977), .Z(n23048) );
  AND U23716 ( .A(b[31]), .B(a[137]), .Z(n23047) );
  XNOR U23717 ( .A(n23048), .B(n23047), .Z(n23049) );
  NAND U23718 ( .A(b[0]), .B(a[169]), .Z(n22979) );
  XNOR U23719 ( .A(b[1]), .B(n22979), .Z(n22981) );
  NANDN U23720 ( .A(b[0]), .B(a[168]), .Z(n22980) );
  NAND U23721 ( .A(n22981), .B(n22980), .Z(n23050) );
  XNOR U23722 ( .A(n23049), .B(n23050), .Z(n23089) );
  NAND U23723 ( .A(n38185), .B(n22982), .Z(n22984) );
  XOR U23724 ( .A(b[23]), .B(a[147]), .Z(n23131) );
  NAND U23725 ( .A(n38132), .B(n23131), .Z(n22983) );
  AND U23726 ( .A(n22984), .B(n22983), .Z(n23122) );
  NAND U23727 ( .A(n184), .B(n22985), .Z(n22987) );
  XOR U23728 ( .A(b[7]), .B(a[163]), .Z(n23134) );
  NAND U23729 ( .A(n36592), .B(n23134), .Z(n22986) );
  AND U23730 ( .A(n22987), .B(n22986), .Z(n23120) );
  NAND U23731 ( .A(n38289), .B(n22988), .Z(n22990) );
  XOR U23732 ( .A(b[25]), .B(a[145]), .Z(n23137) );
  NAND U23733 ( .A(n38247), .B(n23137), .Z(n22989) );
  NAND U23734 ( .A(n22990), .B(n22989), .Z(n23119) );
  XNOR U23735 ( .A(n23120), .B(n23119), .Z(n23121) );
  XOR U23736 ( .A(n23122), .B(n23121), .Z(n23090) );
  XNOR U23737 ( .A(n23089), .B(n23090), .Z(n23091) );
  NAND U23738 ( .A(n187), .B(n22991), .Z(n22993) );
  XOR U23739 ( .A(b[13]), .B(a[157]), .Z(n23140) );
  NAND U23740 ( .A(n37295), .B(n23140), .Z(n22992) );
  AND U23741 ( .A(n22993), .B(n22992), .Z(n23084) );
  NAND U23742 ( .A(n186), .B(n22994), .Z(n22996) );
  XOR U23743 ( .A(b[11]), .B(a[159]), .Z(n23143) );
  NAND U23744 ( .A(n37097), .B(n23143), .Z(n22995) );
  NAND U23745 ( .A(n22996), .B(n22995), .Z(n23083) );
  XNOR U23746 ( .A(n23084), .B(n23083), .Z(n23085) );
  NAND U23747 ( .A(n188), .B(n22997), .Z(n22999) );
  XOR U23748 ( .A(b[15]), .B(a[155]), .Z(n23146) );
  NAND U23749 ( .A(n37382), .B(n23146), .Z(n22998) );
  AND U23750 ( .A(n22999), .B(n22998), .Z(n23080) );
  NAND U23751 ( .A(n38064), .B(n23000), .Z(n23002) );
  XOR U23752 ( .A(b[21]), .B(a[149]), .Z(n23149) );
  NAND U23753 ( .A(n37993), .B(n23149), .Z(n23001) );
  AND U23754 ( .A(n23002), .B(n23001), .Z(n23078) );
  NAND U23755 ( .A(n185), .B(n23003), .Z(n23005) );
  XOR U23756 ( .A(b[9]), .B(a[161]), .Z(n23152) );
  NAND U23757 ( .A(n36805), .B(n23152), .Z(n23004) );
  NAND U23758 ( .A(n23005), .B(n23004), .Z(n23077) );
  XNOR U23759 ( .A(n23078), .B(n23077), .Z(n23079) );
  XOR U23760 ( .A(n23080), .B(n23079), .Z(n23086) );
  XOR U23761 ( .A(n23085), .B(n23086), .Z(n23092) );
  XOR U23762 ( .A(n23091), .B(n23092), .Z(n23104) );
  XNOR U23763 ( .A(n23103), .B(n23104), .Z(n23035) );
  XNOR U23764 ( .A(n23036), .B(n23035), .Z(n23037) );
  XOR U23765 ( .A(n23038), .B(n23037), .Z(n23156) );
  XNOR U23766 ( .A(n23155), .B(n23156), .Z(n23157) );
  XNOR U23767 ( .A(n23158), .B(n23157), .Z(n23031) );
  XOR U23768 ( .A(n23032), .B(n23031), .Z(n23024) );
  NANDN U23769 ( .A(n23007), .B(n23006), .Z(n23011) );
  NANDN U23770 ( .A(n23009), .B(n23008), .Z(n23010) );
  AND U23771 ( .A(n23011), .B(n23010), .Z(n23023) );
  XOR U23772 ( .A(n23024), .B(n23023), .Z(n23026) );
  XNOR U23773 ( .A(n23025), .B(n23026), .Z(n23017) );
  XNOR U23774 ( .A(n23018), .B(n23017), .Z(n23019) );
  XNOR U23775 ( .A(n23020), .B(n23019), .Z(n23161) );
  XNOR U23776 ( .A(sreg[393]), .B(n23161), .Z(n23163) );
  NANDN U23777 ( .A(sreg[392]), .B(n23012), .Z(n23016) );
  NAND U23778 ( .A(n23014), .B(n23013), .Z(n23015) );
  NAND U23779 ( .A(n23016), .B(n23015), .Z(n23162) );
  XNOR U23780 ( .A(n23163), .B(n23162), .Z(c[393]) );
  NANDN U23781 ( .A(n23018), .B(n23017), .Z(n23022) );
  NANDN U23782 ( .A(n23020), .B(n23019), .Z(n23021) );
  AND U23783 ( .A(n23022), .B(n23021), .Z(n23169) );
  NANDN U23784 ( .A(n23024), .B(n23023), .Z(n23028) );
  NANDN U23785 ( .A(n23026), .B(n23025), .Z(n23027) );
  AND U23786 ( .A(n23028), .B(n23027), .Z(n23167) );
  NANDN U23787 ( .A(n23030), .B(n23029), .Z(n23034) );
  NAND U23788 ( .A(n23032), .B(n23031), .Z(n23033) );
  AND U23789 ( .A(n23034), .B(n23033), .Z(n23174) );
  NANDN U23790 ( .A(n23036), .B(n23035), .Z(n23040) );
  NANDN U23791 ( .A(n23038), .B(n23037), .Z(n23039) );
  AND U23792 ( .A(n23040), .B(n23039), .Z(n23305) );
  NANDN U23793 ( .A(n23042), .B(n23041), .Z(n23046) );
  NAND U23794 ( .A(n23044), .B(n23043), .Z(n23045) );
  AND U23795 ( .A(n23046), .B(n23045), .Z(n23304) );
  XNOR U23796 ( .A(n23305), .B(n23304), .Z(n23307) );
  NANDN U23797 ( .A(n23048), .B(n23047), .Z(n23052) );
  NANDN U23798 ( .A(n23050), .B(n23049), .Z(n23051) );
  AND U23799 ( .A(n23052), .B(n23051), .Z(n23252) );
  NAND U23800 ( .A(n38385), .B(n23053), .Z(n23055) );
  XOR U23801 ( .A(b[27]), .B(a[144]), .Z(n23196) );
  NAND U23802 ( .A(n38343), .B(n23196), .Z(n23054) );
  AND U23803 ( .A(n23055), .B(n23054), .Z(n23259) );
  NAND U23804 ( .A(n183), .B(n23056), .Z(n23058) );
  XOR U23805 ( .A(b[5]), .B(a[166]), .Z(n23199) );
  NAND U23806 ( .A(n36296), .B(n23199), .Z(n23057) );
  AND U23807 ( .A(n23058), .B(n23057), .Z(n23257) );
  NAND U23808 ( .A(n190), .B(n23059), .Z(n23061) );
  XOR U23809 ( .A(b[19]), .B(a[152]), .Z(n23202) );
  NAND U23810 ( .A(n37821), .B(n23202), .Z(n23060) );
  NAND U23811 ( .A(n23061), .B(n23060), .Z(n23256) );
  XNOR U23812 ( .A(n23257), .B(n23256), .Z(n23258) );
  XNOR U23813 ( .A(n23259), .B(n23258), .Z(n23250) );
  NAND U23814 ( .A(n38470), .B(n23062), .Z(n23064) );
  XOR U23815 ( .A(b[31]), .B(a[140]), .Z(n23205) );
  NAND U23816 ( .A(n38453), .B(n23205), .Z(n23063) );
  AND U23817 ( .A(n23064), .B(n23063), .Z(n23217) );
  NAND U23818 ( .A(n181), .B(n23065), .Z(n23067) );
  XOR U23819 ( .A(b[3]), .B(a[168]), .Z(n23208) );
  NAND U23820 ( .A(n182), .B(n23208), .Z(n23066) );
  AND U23821 ( .A(n23067), .B(n23066), .Z(n23215) );
  NAND U23822 ( .A(n189), .B(n23068), .Z(n23070) );
  XOR U23823 ( .A(b[17]), .B(a[154]), .Z(n23211) );
  NAND U23824 ( .A(n37652), .B(n23211), .Z(n23069) );
  NAND U23825 ( .A(n23070), .B(n23069), .Z(n23214) );
  XNOR U23826 ( .A(n23215), .B(n23214), .Z(n23216) );
  XOR U23827 ( .A(n23217), .B(n23216), .Z(n23251) );
  XOR U23828 ( .A(n23250), .B(n23251), .Z(n23253) );
  XOR U23829 ( .A(n23252), .B(n23253), .Z(n23185) );
  NANDN U23830 ( .A(n23072), .B(n23071), .Z(n23076) );
  NANDN U23831 ( .A(n23074), .B(n23073), .Z(n23075) );
  AND U23832 ( .A(n23076), .B(n23075), .Z(n23238) );
  NANDN U23833 ( .A(n23078), .B(n23077), .Z(n23082) );
  NANDN U23834 ( .A(n23080), .B(n23079), .Z(n23081) );
  NAND U23835 ( .A(n23082), .B(n23081), .Z(n23239) );
  XNOR U23836 ( .A(n23238), .B(n23239), .Z(n23240) );
  NANDN U23837 ( .A(n23084), .B(n23083), .Z(n23088) );
  NANDN U23838 ( .A(n23086), .B(n23085), .Z(n23087) );
  NAND U23839 ( .A(n23088), .B(n23087), .Z(n23241) );
  XNOR U23840 ( .A(n23240), .B(n23241), .Z(n23184) );
  XNOR U23841 ( .A(n23185), .B(n23184), .Z(n23187) );
  NANDN U23842 ( .A(n23090), .B(n23089), .Z(n23094) );
  NANDN U23843 ( .A(n23092), .B(n23091), .Z(n23093) );
  AND U23844 ( .A(n23094), .B(n23093), .Z(n23186) );
  XOR U23845 ( .A(n23187), .B(n23186), .Z(n23301) );
  NANDN U23846 ( .A(n23096), .B(n23095), .Z(n23100) );
  NANDN U23847 ( .A(n23098), .B(n23097), .Z(n23099) );
  AND U23848 ( .A(n23100), .B(n23099), .Z(n23298) );
  NANDN U23849 ( .A(n23102), .B(n23101), .Z(n23106) );
  NANDN U23850 ( .A(n23104), .B(n23103), .Z(n23105) );
  AND U23851 ( .A(n23106), .B(n23105), .Z(n23181) );
  NANDN U23852 ( .A(n23108), .B(n23107), .Z(n23112) );
  OR U23853 ( .A(n23110), .B(n23109), .Z(n23111) );
  AND U23854 ( .A(n23112), .B(n23111), .Z(n23179) );
  NANDN U23855 ( .A(n23114), .B(n23113), .Z(n23118) );
  NANDN U23856 ( .A(n23116), .B(n23115), .Z(n23117) );
  AND U23857 ( .A(n23118), .B(n23117), .Z(n23245) );
  NANDN U23858 ( .A(n23120), .B(n23119), .Z(n23124) );
  NANDN U23859 ( .A(n23122), .B(n23121), .Z(n23123) );
  NAND U23860 ( .A(n23124), .B(n23123), .Z(n23244) );
  XNOR U23861 ( .A(n23245), .B(n23244), .Z(n23246) );
  NAND U23862 ( .A(b[0]), .B(a[170]), .Z(n23125) );
  XNOR U23863 ( .A(b[1]), .B(n23125), .Z(n23127) );
  NANDN U23864 ( .A(b[0]), .B(a[169]), .Z(n23126) );
  NAND U23865 ( .A(n23127), .B(n23126), .Z(n23193) );
  NAND U23866 ( .A(n194), .B(n23128), .Z(n23130) );
  XOR U23867 ( .A(b[29]), .B(a[142]), .Z(n23271) );
  NAND U23868 ( .A(n38456), .B(n23271), .Z(n23129) );
  AND U23869 ( .A(n23130), .B(n23129), .Z(n23191) );
  AND U23870 ( .A(b[31]), .B(a[138]), .Z(n23190) );
  XNOR U23871 ( .A(n23191), .B(n23190), .Z(n23192) );
  XNOR U23872 ( .A(n23193), .B(n23192), .Z(n23232) );
  NAND U23873 ( .A(n38185), .B(n23131), .Z(n23133) );
  XOR U23874 ( .A(b[23]), .B(a[148]), .Z(n23274) );
  NAND U23875 ( .A(n38132), .B(n23274), .Z(n23132) );
  AND U23876 ( .A(n23133), .B(n23132), .Z(n23265) );
  NAND U23877 ( .A(n184), .B(n23134), .Z(n23136) );
  XOR U23878 ( .A(b[7]), .B(a[164]), .Z(n23277) );
  NAND U23879 ( .A(n36592), .B(n23277), .Z(n23135) );
  AND U23880 ( .A(n23136), .B(n23135), .Z(n23263) );
  NAND U23881 ( .A(n38289), .B(n23137), .Z(n23139) );
  XOR U23882 ( .A(b[25]), .B(a[146]), .Z(n23280) );
  NAND U23883 ( .A(n38247), .B(n23280), .Z(n23138) );
  NAND U23884 ( .A(n23139), .B(n23138), .Z(n23262) );
  XNOR U23885 ( .A(n23263), .B(n23262), .Z(n23264) );
  XOR U23886 ( .A(n23265), .B(n23264), .Z(n23233) );
  XNOR U23887 ( .A(n23232), .B(n23233), .Z(n23234) );
  NAND U23888 ( .A(n187), .B(n23140), .Z(n23142) );
  XOR U23889 ( .A(b[13]), .B(a[158]), .Z(n23283) );
  NAND U23890 ( .A(n37295), .B(n23283), .Z(n23141) );
  AND U23891 ( .A(n23142), .B(n23141), .Z(n23227) );
  NAND U23892 ( .A(n186), .B(n23143), .Z(n23145) );
  XOR U23893 ( .A(b[11]), .B(a[160]), .Z(n23286) );
  NAND U23894 ( .A(n37097), .B(n23286), .Z(n23144) );
  NAND U23895 ( .A(n23145), .B(n23144), .Z(n23226) );
  XNOR U23896 ( .A(n23227), .B(n23226), .Z(n23228) );
  NAND U23897 ( .A(n188), .B(n23146), .Z(n23148) );
  XOR U23898 ( .A(b[15]), .B(a[156]), .Z(n23289) );
  NAND U23899 ( .A(n37382), .B(n23289), .Z(n23147) );
  AND U23900 ( .A(n23148), .B(n23147), .Z(n23223) );
  NAND U23901 ( .A(n38064), .B(n23149), .Z(n23151) );
  XOR U23902 ( .A(b[21]), .B(a[150]), .Z(n23292) );
  NAND U23903 ( .A(n37993), .B(n23292), .Z(n23150) );
  AND U23904 ( .A(n23151), .B(n23150), .Z(n23221) );
  NAND U23905 ( .A(n185), .B(n23152), .Z(n23154) );
  XOR U23906 ( .A(b[9]), .B(a[162]), .Z(n23295) );
  NAND U23907 ( .A(n36805), .B(n23295), .Z(n23153) );
  NAND U23908 ( .A(n23154), .B(n23153), .Z(n23220) );
  XNOR U23909 ( .A(n23221), .B(n23220), .Z(n23222) );
  XOR U23910 ( .A(n23223), .B(n23222), .Z(n23229) );
  XOR U23911 ( .A(n23228), .B(n23229), .Z(n23235) );
  XOR U23912 ( .A(n23234), .B(n23235), .Z(n23247) );
  XNOR U23913 ( .A(n23246), .B(n23247), .Z(n23178) );
  XNOR U23914 ( .A(n23179), .B(n23178), .Z(n23180) );
  XOR U23915 ( .A(n23181), .B(n23180), .Z(n23299) );
  XNOR U23916 ( .A(n23298), .B(n23299), .Z(n23300) );
  XNOR U23917 ( .A(n23301), .B(n23300), .Z(n23306) );
  XOR U23918 ( .A(n23307), .B(n23306), .Z(n23173) );
  NANDN U23919 ( .A(n23156), .B(n23155), .Z(n23160) );
  NANDN U23920 ( .A(n23158), .B(n23157), .Z(n23159) );
  AND U23921 ( .A(n23160), .B(n23159), .Z(n23172) );
  XOR U23922 ( .A(n23173), .B(n23172), .Z(n23175) );
  XNOR U23923 ( .A(n23174), .B(n23175), .Z(n23166) );
  XNOR U23924 ( .A(n23167), .B(n23166), .Z(n23168) );
  XNOR U23925 ( .A(n23169), .B(n23168), .Z(n23310) );
  XNOR U23926 ( .A(sreg[394]), .B(n23310), .Z(n23312) );
  NANDN U23927 ( .A(sreg[393]), .B(n23161), .Z(n23165) );
  NAND U23928 ( .A(n23163), .B(n23162), .Z(n23164) );
  NAND U23929 ( .A(n23165), .B(n23164), .Z(n23311) );
  XNOR U23930 ( .A(n23312), .B(n23311), .Z(c[394]) );
  NANDN U23931 ( .A(n23167), .B(n23166), .Z(n23171) );
  NANDN U23932 ( .A(n23169), .B(n23168), .Z(n23170) );
  AND U23933 ( .A(n23171), .B(n23170), .Z(n23318) );
  NANDN U23934 ( .A(n23173), .B(n23172), .Z(n23177) );
  NANDN U23935 ( .A(n23175), .B(n23174), .Z(n23176) );
  AND U23936 ( .A(n23177), .B(n23176), .Z(n23316) );
  NANDN U23937 ( .A(n23179), .B(n23178), .Z(n23183) );
  NANDN U23938 ( .A(n23181), .B(n23180), .Z(n23182) );
  AND U23939 ( .A(n23183), .B(n23182), .Z(n23452) );
  NANDN U23940 ( .A(n23185), .B(n23184), .Z(n23189) );
  NAND U23941 ( .A(n23187), .B(n23186), .Z(n23188) );
  AND U23942 ( .A(n23189), .B(n23188), .Z(n23451) );
  XNOR U23943 ( .A(n23452), .B(n23451), .Z(n23454) );
  NANDN U23944 ( .A(n23191), .B(n23190), .Z(n23195) );
  NANDN U23945 ( .A(n23193), .B(n23192), .Z(n23194) );
  AND U23946 ( .A(n23195), .B(n23194), .Z(n23399) );
  NAND U23947 ( .A(n38385), .B(n23196), .Z(n23198) );
  XOR U23948 ( .A(b[27]), .B(a[145]), .Z(n23345) );
  NAND U23949 ( .A(n38343), .B(n23345), .Z(n23197) );
  AND U23950 ( .A(n23198), .B(n23197), .Z(n23406) );
  NAND U23951 ( .A(n183), .B(n23199), .Z(n23201) );
  XOR U23952 ( .A(b[5]), .B(a[167]), .Z(n23348) );
  NAND U23953 ( .A(n36296), .B(n23348), .Z(n23200) );
  AND U23954 ( .A(n23201), .B(n23200), .Z(n23404) );
  NAND U23955 ( .A(n190), .B(n23202), .Z(n23204) );
  XOR U23956 ( .A(b[19]), .B(a[153]), .Z(n23351) );
  NAND U23957 ( .A(n37821), .B(n23351), .Z(n23203) );
  NAND U23958 ( .A(n23204), .B(n23203), .Z(n23403) );
  XNOR U23959 ( .A(n23404), .B(n23403), .Z(n23405) );
  XNOR U23960 ( .A(n23406), .B(n23405), .Z(n23397) );
  NAND U23961 ( .A(n38470), .B(n23205), .Z(n23207) );
  XOR U23962 ( .A(b[31]), .B(a[141]), .Z(n23354) );
  NAND U23963 ( .A(n38453), .B(n23354), .Z(n23206) );
  AND U23964 ( .A(n23207), .B(n23206), .Z(n23366) );
  NAND U23965 ( .A(n181), .B(n23208), .Z(n23210) );
  XOR U23966 ( .A(b[3]), .B(a[169]), .Z(n23357) );
  NAND U23967 ( .A(n182), .B(n23357), .Z(n23209) );
  AND U23968 ( .A(n23210), .B(n23209), .Z(n23364) );
  NAND U23969 ( .A(n189), .B(n23211), .Z(n23213) );
  XOR U23970 ( .A(b[17]), .B(a[155]), .Z(n23360) );
  NAND U23971 ( .A(n37652), .B(n23360), .Z(n23212) );
  NAND U23972 ( .A(n23213), .B(n23212), .Z(n23363) );
  XNOR U23973 ( .A(n23364), .B(n23363), .Z(n23365) );
  XOR U23974 ( .A(n23366), .B(n23365), .Z(n23398) );
  XOR U23975 ( .A(n23397), .B(n23398), .Z(n23400) );
  XOR U23976 ( .A(n23399), .B(n23400), .Z(n23334) );
  NANDN U23977 ( .A(n23215), .B(n23214), .Z(n23219) );
  NANDN U23978 ( .A(n23217), .B(n23216), .Z(n23218) );
  AND U23979 ( .A(n23219), .B(n23218), .Z(n23387) );
  NANDN U23980 ( .A(n23221), .B(n23220), .Z(n23225) );
  NANDN U23981 ( .A(n23223), .B(n23222), .Z(n23224) );
  NAND U23982 ( .A(n23225), .B(n23224), .Z(n23388) );
  XNOR U23983 ( .A(n23387), .B(n23388), .Z(n23389) );
  NANDN U23984 ( .A(n23227), .B(n23226), .Z(n23231) );
  NANDN U23985 ( .A(n23229), .B(n23228), .Z(n23230) );
  NAND U23986 ( .A(n23231), .B(n23230), .Z(n23390) );
  XNOR U23987 ( .A(n23389), .B(n23390), .Z(n23333) );
  XNOR U23988 ( .A(n23334), .B(n23333), .Z(n23336) );
  NANDN U23989 ( .A(n23233), .B(n23232), .Z(n23237) );
  NANDN U23990 ( .A(n23235), .B(n23234), .Z(n23236) );
  AND U23991 ( .A(n23237), .B(n23236), .Z(n23335) );
  XOR U23992 ( .A(n23336), .B(n23335), .Z(n23448) );
  NANDN U23993 ( .A(n23239), .B(n23238), .Z(n23243) );
  NANDN U23994 ( .A(n23241), .B(n23240), .Z(n23242) );
  AND U23995 ( .A(n23243), .B(n23242), .Z(n23445) );
  NANDN U23996 ( .A(n23245), .B(n23244), .Z(n23249) );
  NANDN U23997 ( .A(n23247), .B(n23246), .Z(n23248) );
  AND U23998 ( .A(n23249), .B(n23248), .Z(n23330) );
  NANDN U23999 ( .A(n23251), .B(n23250), .Z(n23255) );
  OR U24000 ( .A(n23253), .B(n23252), .Z(n23254) );
  AND U24001 ( .A(n23255), .B(n23254), .Z(n23328) );
  NANDN U24002 ( .A(n23257), .B(n23256), .Z(n23261) );
  NANDN U24003 ( .A(n23259), .B(n23258), .Z(n23260) );
  AND U24004 ( .A(n23261), .B(n23260), .Z(n23394) );
  NANDN U24005 ( .A(n23263), .B(n23262), .Z(n23267) );
  NANDN U24006 ( .A(n23265), .B(n23264), .Z(n23266) );
  NAND U24007 ( .A(n23267), .B(n23266), .Z(n23393) );
  XNOR U24008 ( .A(n23394), .B(n23393), .Z(n23396) );
  NAND U24009 ( .A(b[0]), .B(a[171]), .Z(n23268) );
  XNOR U24010 ( .A(b[1]), .B(n23268), .Z(n23270) );
  NANDN U24011 ( .A(b[0]), .B(a[170]), .Z(n23269) );
  NAND U24012 ( .A(n23270), .B(n23269), .Z(n23342) );
  NAND U24013 ( .A(n194), .B(n23271), .Z(n23273) );
  XOR U24014 ( .A(b[29]), .B(a[143]), .Z(n23415) );
  NAND U24015 ( .A(n38456), .B(n23415), .Z(n23272) );
  AND U24016 ( .A(n23273), .B(n23272), .Z(n23340) );
  AND U24017 ( .A(b[31]), .B(a[139]), .Z(n23339) );
  XNOR U24018 ( .A(n23340), .B(n23339), .Z(n23341) );
  XNOR U24019 ( .A(n23342), .B(n23341), .Z(n23382) );
  NAND U24020 ( .A(n38185), .B(n23274), .Z(n23276) );
  XOR U24021 ( .A(b[23]), .B(a[149]), .Z(n23421) );
  NAND U24022 ( .A(n38132), .B(n23421), .Z(n23275) );
  AND U24023 ( .A(n23276), .B(n23275), .Z(n23411) );
  NAND U24024 ( .A(n184), .B(n23277), .Z(n23279) );
  XOR U24025 ( .A(b[7]), .B(a[165]), .Z(n23424) );
  NAND U24026 ( .A(n36592), .B(n23424), .Z(n23278) );
  AND U24027 ( .A(n23279), .B(n23278), .Z(n23410) );
  NAND U24028 ( .A(n38289), .B(n23280), .Z(n23282) );
  XOR U24029 ( .A(b[25]), .B(a[147]), .Z(n23427) );
  NAND U24030 ( .A(n38247), .B(n23427), .Z(n23281) );
  NAND U24031 ( .A(n23282), .B(n23281), .Z(n23409) );
  XOR U24032 ( .A(n23410), .B(n23409), .Z(n23412) );
  XOR U24033 ( .A(n23411), .B(n23412), .Z(n23381) );
  XOR U24034 ( .A(n23382), .B(n23381), .Z(n23384) );
  NAND U24035 ( .A(n187), .B(n23283), .Z(n23285) );
  XOR U24036 ( .A(b[13]), .B(a[159]), .Z(n23430) );
  NAND U24037 ( .A(n37295), .B(n23430), .Z(n23284) );
  AND U24038 ( .A(n23285), .B(n23284), .Z(n23376) );
  NAND U24039 ( .A(n186), .B(n23286), .Z(n23288) );
  XOR U24040 ( .A(b[11]), .B(a[161]), .Z(n23433) );
  NAND U24041 ( .A(n37097), .B(n23433), .Z(n23287) );
  NAND U24042 ( .A(n23288), .B(n23287), .Z(n23375) );
  XNOR U24043 ( .A(n23376), .B(n23375), .Z(n23378) );
  NAND U24044 ( .A(n188), .B(n23289), .Z(n23291) );
  XOR U24045 ( .A(b[15]), .B(a[157]), .Z(n23436) );
  NAND U24046 ( .A(n37382), .B(n23436), .Z(n23290) );
  AND U24047 ( .A(n23291), .B(n23290), .Z(n23372) );
  NAND U24048 ( .A(n38064), .B(n23292), .Z(n23294) );
  XOR U24049 ( .A(b[21]), .B(a[151]), .Z(n23439) );
  NAND U24050 ( .A(n37993), .B(n23439), .Z(n23293) );
  AND U24051 ( .A(n23294), .B(n23293), .Z(n23370) );
  NAND U24052 ( .A(n185), .B(n23295), .Z(n23297) );
  XOR U24053 ( .A(b[9]), .B(a[163]), .Z(n23442) );
  NAND U24054 ( .A(n36805), .B(n23442), .Z(n23296) );
  NAND U24055 ( .A(n23297), .B(n23296), .Z(n23369) );
  XNOR U24056 ( .A(n23370), .B(n23369), .Z(n23371) );
  XNOR U24057 ( .A(n23372), .B(n23371), .Z(n23377) );
  XOR U24058 ( .A(n23378), .B(n23377), .Z(n23383) );
  XNOR U24059 ( .A(n23384), .B(n23383), .Z(n23395) );
  XNOR U24060 ( .A(n23396), .B(n23395), .Z(n23327) );
  XNOR U24061 ( .A(n23328), .B(n23327), .Z(n23329) );
  XOR U24062 ( .A(n23330), .B(n23329), .Z(n23446) );
  XNOR U24063 ( .A(n23445), .B(n23446), .Z(n23447) );
  XNOR U24064 ( .A(n23448), .B(n23447), .Z(n23453) );
  XOR U24065 ( .A(n23454), .B(n23453), .Z(n23322) );
  NANDN U24066 ( .A(n23299), .B(n23298), .Z(n23303) );
  NANDN U24067 ( .A(n23301), .B(n23300), .Z(n23302) );
  AND U24068 ( .A(n23303), .B(n23302), .Z(n23321) );
  XNOR U24069 ( .A(n23322), .B(n23321), .Z(n23323) );
  NANDN U24070 ( .A(n23305), .B(n23304), .Z(n23309) );
  NAND U24071 ( .A(n23307), .B(n23306), .Z(n23308) );
  NAND U24072 ( .A(n23309), .B(n23308), .Z(n23324) );
  XNOR U24073 ( .A(n23323), .B(n23324), .Z(n23315) );
  XNOR U24074 ( .A(n23316), .B(n23315), .Z(n23317) );
  XNOR U24075 ( .A(n23318), .B(n23317), .Z(n23457) );
  XNOR U24076 ( .A(sreg[395]), .B(n23457), .Z(n23459) );
  NANDN U24077 ( .A(sreg[394]), .B(n23310), .Z(n23314) );
  NAND U24078 ( .A(n23312), .B(n23311), .Z(n23313) );
  NAND U24079 ( .A(n23314), .B(n23313), .Z(n23458) );
  XNOR U24080 ( .A(n23459), .B(n23458), .Z(c[395]) );
  NANDN U24081 ( .A(n23316), .B(n23315), .Z(n23320) );
  NANDN U24082 ( .A(n23318), .B(n23317), .Z(n23319) );
  AND U24083 ( .A(n23320), .B(n23319), .Z(n23465) );
  NANDN U24084 ( .A(n23322), .B(n23321), .Z(n23326) );
  NANDN U24085 ( .A(n23324), .B(n23323), .Z(n23325) );
  AND U24086 ( .A(n23326), .B(n23325), .Z(n23463) );
  NANDN U24087 ( .A(n23328), .B(n23327), .Z(n23332) );
  NANDN U24088 ( .A(n23330), .B(n23329), .Z(n23331) );
  AND U24089 ( .A(n23332), .B(n23331), .Z(n23599) );
  NANDN U24090 ( .A(n23334), .B(n23333), .Z(n23338) );
  NAND U24091 ( .A(n23336), .B(n23335), .Z(n23337) );
  AND U24092 ( .A(n23338), .B(n23337), .Z(n23598) );
  XNOR U24093 ( .A(n23599), .B(n23598), .Z(n23601) );
  NANDN U24094 ( .A(n23340), .B(n23339), .Z(n23344) );
  NANDN U24095 ( .A(n23342), .B(n23341), .Z(n23343) );
  AND U24096 ( .A(n23344), .B(n23343), .Z(n23534) );
  NAND U24097 ( .A(n38385), .B(n23345), .Z(n23347) );
  XOR U24098 ( .A(b[27]), .B(a[146]), .Z(n23480) );
  NAND U24099 ( .A(n38343), .B(n23480), .Z(n23346) );
  AND U24100 ( .A(n23347), .B(n23346), .Z(n23541) );
  NAND U24101 ( .A(n183), .B(n23348), .Z(n23350) );
  XOR U24102 ( .A(b[5]), .B(a[168]), .Z(n23483) );
  NAND U24103 ( .A(n36296), .B(n23483), .Z(n23349) );
  AND U24104 ( .A(n23350), .B(n23349), .Z(n23539) );
  NAND U24105 ( .A(n190), .B(n23351), .Z(n23353) );
  XOR U24106 ( .A(b[19]), .B(a[154]), .Z(n23486) );
  NAND U24107 ( .A(n37821), .B(n23486), .Z(n23352) );
  NAND U24108 ( .A(n23353), .B(n23352), .Z(n23538) );
  XNOR U24109 ( .A(n23539), .B(n23538), .Z(n23540) );
  XNOR U24110 ( .A(n23541), .B(n23540), .Z(n23532) );
  NAND U24111 ( .A(n38470), .B(n23354), .Z(n23356) );
  XOR U24112 ( .A(b[31]), .B(a[142]), .Z(n23489) );
  NAND U24113 ( .A(n38453), .B(n23489), .Z(n23355) );
  AND U24114 ( .A(n23356), .B(n23355), .Z(n23501) );
  NAND U24115 ( .A(n181), .B(n23357), .Z(n23359) );
  XOR U24116 ( .A(b[3]), .B(a[170]), .Z(n23492) );
  NAND U24117 ( .A(n182), .B(n23492), .Z(n23358) );
  AND U24118 ( .A(n23359), .B(n23358), .Z(n23499) );
  NAND U24119 ( .A(n189), .B(n23360), .Z(n23362) );
  XOR U24120 ( .A(b[17]), .B(a[156]), .Z(n23495) );
  NAND U24121 ( .A(n37652), .B(n23495), .Z(n23361) );
  NAND U24122 ( .A(n23362), .B(n23361), .Z(n23498) );
  XNOR U24123 ( .A(n23499), .B(n23498), .Z(n23500) );
  XOR U24124 ( .A(n23501), .B(n23500), .Z(n23533) );
  XOR U24125 ( .A(n23532), .B(n23533), .Z(n23535) );
  XOR U24126 ( .A(n23534), .B(n23535), .Z(n23581) );
  NANDN U24127 ( .A(n23364), .B(n23363), .Z(n23368) );
  NANDN U24128 ( .A(n23366), .B(n23365), .Z(n23367) );
  AND U24129 ( .A(n23368), .B(n23367), .Z(n23522) );
  NANDN U24130 ( .A(n23370), .B(n23369), .Z(n23374) );
  NANDN U24131 ( .A(n23372), .B(n23371), .Z(n23373) );
  NAND U24132 ( .A(n23374), .B(n23373), .Z(n23523) );
  XNOR U24133 ( .A(n23522), .B(n23523), .Z(n23524) );
  NANDN U24134 ( .A(n23376), .B(n23375), .Z(n23380) );
  NAND U24135 ( .A(n23378), .B(n23377), .Z(n23379) );
  NAND U24136 ( .A(n23380), .B(n23379), .Z(n23525) );
  XNOR U24137 ( .A(n23524), .B(n23525), .Z(n23580) );
  XNOR U24138 ( .A(n23581), .B(n23580), .Z(n23583) );
  NAND U24139 ( .A(n23382), .B(n23381), .Z(n23386) );
  NAND U24140 ( .A(n23384), .B(n23383), .Z(n23385) );
  AND U24141 ( .A(n23386), .B(n23385), .Z(n23582) );
  XOR U24142 ( .A(n23583), .B(n23582), .Z(n23595) );
  NANDN U24143 ( .A(n23388), .B(n23387), .Z(n23392) );
  NANDN U24144 ( .A(n23390), .B(n23389), .Z(n23391) );
  AND U24145 ( .A(n23392), .B(n23391), .Z(n23592) );
  NANDN U24146 ( .A(n23398), .B(n23397), .Z(n23402) );
  OR U24147 ( .A(n23400), .B(n23399), .Z(n23401) );
  AND U24148 ( .A(n23402), .B(n23401), .Z(n23587) );
  NANDN U24149 ( .A(n23404), .B(n23403), .Z(n23408) );
  NANDN U24150 ( .A(n23406), .B(n23405), .Z(n23407) );
  AND U24151 ( .A(n23408), .B(n23407), .Z(n23529) );
  NANDN U24152 ( .A(n23410), .B(n23409), .Z(n23414) );
  OR U24153 ( .A(n23412), .B(n23411), .Z(n23413) );
  NAND U24154 ( .A(n23414), .B(n23413), .Z(n23528) );
  XNOR U24155 ( .A(n23529), .B(n23528), .Z(n23531) );
  NAND U24156 ( .A(n194), .B(n23415), .Z(n23417) );
  XOR U24157 ( .A(b[29]), .B(a[144]), .Z(n23553) );
  NAND U24158 ( .A(n38456), .B(n23553), .Z(n23416) );
  AND U24159 ( .A(n23417), .B(n23416), .Z(n23475) );
  AND U24160 ( .A(b[31]), .B(a[140]), .Z(n23474) );
  XNOR U24161 ( .A(n23475), .B(n23474), .Z(n23476) );
  NAND U24162 ( .A(b[0]), .B(a[172]), .Z(n23418) );
  XNOR U24163 ( .A(b[1]), .B(n23418), .Z(n23420) );
  NANDN U24164 ( .A(b[0]), .B(a[171]), .Z(n23419) );
  NAND U24165 ( .A(n23420), .B(n23419), .Z(n23477) );
  XNOR U24166 ( .A(n23476), .B(n23477), .Z(n23517) );
  NAND U24167 ( .A(n38185), .B(n23421), .Z(n23423) );
  XOR U24168 ( .A(b[23]), .B(a[150]), .Z(n23556) );
  NAND U24169 ( .A(n38132), .B(n23556), .Z(n23422) );
  AND U24170 ( .A(n23423), .B(n23422), .Z(n23546) );
  NAND U24171 ( .A(n184), .B(n23424), .Z(n23426) );
  XOR U24172 ( .A(b[7]), .B(a[166]), .Z(n23559) );
  NAND U24173 ( .A(n36592), .B(n23559), .Z(n23425) );
  AND U24174 ( .A(n23426), .B(n23425), .Z(n23545) );
  NAND U24175 ( .A(n38289), .B(n23427), .Z(n23429) );
  XOR U24176 ( .A(b[25]), .B(a[148]), .Z(n23562) );
  NAND U24177 ( .A(n38247), .B(n23562), .Z(n23428) );
  NAND U24178 ( .A(n23429), .B(n23428), .Z(n23544) );
  XOR U24179 ( .A(n23545), .B(n23544), .Z(n23547) );
  XOR U24180 ( .A(n23546), .B(n23547), .Z(n23516) );
  XOR U24181 ( .A(n23517), .B(n23516), .Z(n23519) );
  NAND U24182 ( .A(n187), .B(n23430), .Z(n23432) );
  XOR U24183 ( .A(b[13]), .B(a[160]), .Z(n23565) );
  NAND U24184 ( .A(n37295), .B(n23565), .Z(n23431) );
  AND U24185 ( .A(n23432), .B(n23431), .Z(n23511) );
  NAND U24186 ( .A(n186), .B(n23433), .Z(n23435) );
  XOR U24187 ( .A(b[11]), .B(a[162]), .Z(n23568) );
  NAND U24188 ( .A(n37097), .B(n23568), .Z(n23434) );
  NAND U24189 ( .A(n23435), .B(n23434), .Z(n23510) );
  XNOR U24190 ( .A(n23511), .B(n23510), .Z(n23513) );
  NAND U24191 ( .A(n188), .B(n23436), .Z(n23438) );
  XOR U24192 ( .A(b[15]), .B(a[158]), .Z(n23571) );
  NAND U24193 ( .A(n37382), .B(n23571), .Z(n23437) );
  AND U24194 ( .A(n23438), .B(n23437), .Z(n23507) );
  NAND U24195 ( .A(n38064), .B(n23439), .Z(n23441) );
  XOR U24196 ( .A(b[21]), .B(a[152]), .Z(n23574) );
  NAND U24197 ( .A(n37993), .B(n23574), .Z(n23440) );
  AND U24198 ( .A(n23441), .B(n23440), .Z(n23505) );
  NAND U24199 ( .A(n185), .B(n23442), .Z(n23444) );
  XOR U24200 ( .A(b[9]), .B(a[164]), .Z(n23577) );
  NAND U24201 ( .A(n36805), .B(n23577), .Z(n23443) );
  NAND U24202 ( .A(n23444), .B(n23443), .Z(n23504) );
  XNOR U24203 ( .A(n23505), .B(n23504), .Z(n23506) );
  XNOR U24204 ( .A(n23507), .B(n23506), .Z(n23512) );
  XOR U24205 ( .A(n23513), .B(n23512), .Z(n23518) );
  XNOR U24206 ( .A(n23519), .B(n23518), .Z(n23530) );
  XNOR U24207 ( .A(n23531), .B(n23530), .Z(n23586) );
  XNOR U24208 ( .A(n23587), .B(n23586), .Z(n23588) );
  XOR U24209 ( .A(n23589), .B(n23588), .Z(n23593) );
  XNOR U24210 ( .A(n23592), .B(n23593), .Z(n23594) );
  XNOR U24211 ( .A(n23595), .B(n23594), .Z(n23600) );
  XOR U24212 ( .A(n23601), .B(n23600), .Z(n23469) );
  NANDN U24213 ( .A(n23446), .B(n23445), .Z(n23450) );
  NANDN U24214 ( .A(n23448), .B(n23447), .Z(n23449) );
  AND U24215 ( .A(n23450), .B(n23449), .Z(n23468) );
  XNOR U24216 ( .A(n23469), .B(n23468), .Z(n23470) );
  NANDN U24217 ( .A(n23452), .B(n23451), .Z(n23456) );
  NAND U24218 ( .A(n23454), .B(n23453), .Z(n23455) );
  NAND U24219 ( .A(n23456), .B(n23455), .Z(n23471) );
  XNOR U24220 ( .A(n23470), .B(n23471), .Z(n23462) );
  XNOR U24221 ( .A(n23463), .B(n23462), .Z(n23464) );
  XNOR U24222 ( .A(n23465), .B(n23464), .Z(n23604) );
  XNOR U24223 ( .A(sreg[396]), .B(n23604), .Z(n23606) );
  NANDN U24224 ( .A(sreg[395]), .B(n23457), .Z(n23461) );
  NAND U24225 ( .A(n23459), .B(n23458), .Z(n23460) );
  NAND U24226 ( .A(n23461), .B(n23460), .Z(n23605) );
  XNOR U24227 ( .A(n23606), .B(n23605), .Z(c[396]) );
  NANDN U24228 ( .A(n23463), .B(n23462), .Z(n23467) );
  NANDN U24229 ( .A(n23465), .B(n23464), .Z(n23466) );
  AND U24230 ( .A(n23467), .B(n23466), .Z(n23612) );
  NANDN U24231 ( .A(n23469), .B(n23468), .Z(n23473) );
  NANDN U24232 ( .A(n23471), .B(n23470), .Z(n23472) );
  AND U24233 ( .A(n23473), .B(n23472), .Z(n23610) );
  NANDN U24234 ( .A(n23475), .B(n23474), .Z(n23479) );
  NANDN U24235 ( .A(n23477), .B(n23476), .Z(n23478) );
  AND U24236 ( .A(n23479), .B(n23478), .Z(n23689) );
  NAND U24237 ( .A(n38385), .B(n23480), .Z(n23482) );
  XOR U24238 ( .A(b[27]), .B(a[147]), .Z(n23633) );
  NAND U24239 ( .A(n38343), .B(n23633), .Z(n23481) );
  AND U24240 ( .A(n23482), .B(n23481), .Z(n23696) );
  NAND U24241 ( .A(n183), .B(n23483), .Z(n23485) );
  XOR U24242 ( .A(b[5]), .B(a[169]), .Z(n23636) );
  NAND U24243 ( .A(n36296), .B(n23636), .Z(n23484) );
  AND U24244 ( .A(n23485), .B(n23484), .Z(n23694) );
  NAND U24245 ( .A(n190), .B(n23486), .Z(n23488) );
  XOR U24246 ( .A(b[19]), .B(a[155]), .Z(n23639) );
  NAND U24247 ( .A(n37821), .B(n23639), .Z(n23487) );
  NAND U24248 ( .A(n23488), .B(n23487), .Z(n23693) );
  XNOR U24249 ( .A(n23694), .B(n23693), .Z(n23695) );
  XNOR U24250 ( .A(n23696), .B(n23695), .Z(n23687) );
  NAND U24251 ( .A(n38470), .B(n23489), .Z(n23491) );
  XOR U24252 ( .A(b[31]), .B(a[143]), .Z(n23642) );
  NAND U24253 ( .A(n38453), .B(n23642), .Z(n23490) );
  AND U24254 ( .A(n23491), .B(n23490), .Z(n23654) );
  NAND U24255 ( .A(n181), .B(n23492), .Z(n23494) );
  XOR U24256 ( .A(b[3]), .B(a[171]), .Z(n23645) );
  NAND U24257 ( .A(n182), .B(n23645), .Z(n23493) );
  AND U24258 ( .A(n23494), .B(n23493), .Z(n23652) );
  NAND U24259 ( .A(n189), .B(n23495), .Z(n23497) );
  XOR U24260 ( .A(b[17]), .B(a[157]), .Z(n23648) );
  NAND U24261 ( .A(n37652), .B(n23648), .Z(n23496) );
  NAND U24262 ( .A(n23497), .B(n23496), .Z(n23651) );
  XNOR U24263 ( .A(n23652), .B(n23651), .Z(n23653) );
  XOR U24264 ( .A(n23654), .B(n23653), .Z(n23688) );
  XOR U24265 ( .A(n23687), .B(n23688), .Z(n23690) );
  XOR U24266 ( .A(n23689), .B(n23690), .Z(n23736) );
  NANDN U24267 ( .A(n23499), .B(n23498), .Z(n23503) );
  NANDN U24268 ( .A(n23501), .B(n23500), .Z(n23502) );
  AND U24269 ( .A(n23503), .B(n23502), .Z(n23675) );
  NANDN U24270 ( .A(n23505), .B(n23504), .Z(n23509) );
  NANDN U24271 ( .A(n23507), .B(n23506), .Z(n23508) );
  NAND U24272 ( .A(n23509), .B(n23508), .Z(n23676) );
  XNOR U24273 ( .A(n23675), .B(n23676), .Z(n23677) );
  NANDN U24274 ( .A(n23511), .B(n23510), .Z(n23515) );
  NAND U24275 ( .A(n23513), .B(n23512), .Z(n23514) );
  NAND U24276 ( .A(n23515), .B(n23514), .Z(n23678) );
  XNOR U24277 ( .A(n23677), .B(n23678), .Z(n23735) );
  XNOR U24278 ( .A(n23736), .B(n23735), .Z(n23738) );
  NAND U24279 ( .A(n23517), .B(n23516), .Z(n23521) );
  NAND U24280 ( .A(n23519), .B(n23518), .Z(n23520) );
  AND U24281 ( .A(n23521), .B(n23520), .Z(n23737) );
  XOR U24282 ( .A(n23738), .B(n23737), .Z(n23749) );
  NANDN U24283 ( .A(n23523), .B(n23522), .Z(n23527) );
  NANDN U24284 ( .A(n23525), .B(n23524), .Z(n23526) );
  AND U24285 ( .A(n23527), .B(n23526), .Z(n23747) );
  NANDN U24286 ( .A(n23533), .B(n23532), .Z(n23537) );
  OR U24287 ( .A(n23535), .B(n23534), .Z(n23536) );
  AND U24288 ( .A(n23537), .B(n23536), .Z(n23742) );
  NANDN U24289 ( .A(n23539), .B(n23538), .Z(n23543) );
  NANDN U24290 ( .A(n23541), .B(n23540), .Z(n23542) );
  AND U24291 ( .A(n23543), .B(n23542), .Z(n23682) );
  NANDN U24292 ( .A(n23545), .B(n23544), .Z(n23549) );
  OR U24293 ( .A(n23547), .B(n23546), .Z(n23548) );
  NAND U24294 ( .A(n23549), .B(n23548), .Z(n23681) );
  XNOR U24295 ( .A(n23682), .B(n23681), .Z(n23683) );
  NAND U24296 ( .A(b[0]), .B(a[173]), .Z(n23550) );
  XNOR U24297 ( .A(b[1]), .B(n23550), .Z(n23552) );
  NANDN U24298 ( .A(b[0]), .B(a[172]), .Z(n23551) );
  NAND U24299 ( .A(n23552), .B(n23551), .Z(n23630) );
  NAND U24300 ( .A(n194), .B(n23553), .Z(n23555) );
  XOR U24301 ( .A(b[29]), .B(a[145]), .Z(n23708) );
  NAND U24302 ( .A(n38456), .B(n23708), .Z(n23554) );
  AND U24303 ( .A(n23555), .B(n23554), .Z(n23628) );
  AND U24304 ( .A(b[31]), .B(a[141]), .Z(n23627) );
  XNOR U24305 ( .A(n23628), .B(n23627), .Z(n23629) );
  XNOR U24306 ( .A(n23630), .B(n23629), .Z(n23669) );
  NAND U24307 ( .A(n38185), .B(n23556), .Z(n23558) );
  XOR U24308 ( .A(b[23]), .B(a[151]), .Z(n23711) );
  NAND U24309 ( .A(n38132), .B(n23711), .Z(n23557) );
  AND U24310 ( .A(n23558), .B(n23557), .Z(n23702) );
  NAND U24311 ( .A(n184), .B(n23559), .Z(n23561) );
  XOR U24312 ( .A(b[7]), .B(a[167]), .Z(n23714) );
  NAND U24313 ( .A(n36592), .B(n23714), .Z(n23560) );
  AND U24314 ( .A(n23561), .B(n23560), .Z(n23700) );
  NAND U24315 ( .A(n38289), .B(n23562), .Z(n23564) );
  XOR U24316 ( .A(b[25]), .B(a[149]), .Z(n23717) );
  NAND U24317 ( .A(n38247), .B(n23717), .Z(n23563) );
  NAND U24318 ( .A(n23564), .B(n23563), .Z(n23699) );
  XNOR U24319 ( .A(n23700), .B(n23699), .Z(n23701) );
  XOR U24320 ( .A(n23702), .B(n23701), .Z(n23670) );
  XNOR U24321 ( .A(n23669), .B(n23670), .Z(n23671) );
  NAND U24322 ( .A(n187), .B(n23565), .Z(n23567) );
  XOR U24323 ( .A(b[13]), .B(a[161]), .Z(n23720) );
  NAND U24324 ( .A(n37295), .B(n23720), .Z(n23566) );
  AND U24325 ( .A(n23567), .B(n23566), .Z(n23664) );
  NAND U24326 ( .A(n186), .B(n23568), .Z(n23570) );
  XOR U24327 ( .A(b[11]), .B(a[163]), .Z(n23723) );
  NAND U24328 ( .A(n37097), .B(n23723), .Z(n23569) );
  NAND U24329 ( .A(n23570), .B(n23569), .Z(n23663) );
  XNOR U24330 ( .A(n23664), .B(n23663), .Z(n23665) );
  NAND U24331 ( .A(n188), .B(n23571), .Z(n23573) );
  XOR U24332 ( .A(b[15]), .B(a[159]), .Z(n23726) );
  NAND U24333 ( .A(n37382), .B(n23726), .Z(n23572) );
  AND U24334 ( .A(n23573), .B(n23572), .Z(n23660) );
  NAND U24335 ( .A(n38064), .B(n23574), .Z(n23576) );
  XOR U24336 ( .A(b[21]), .B(a[153]), .Z(n23729) );
  NAND U24337 ( .A(n37993), .B(n23729), .Z(n23575) );
  AND U24338 ( .A(n23576), .B(n23575), .Z(n23658) );
  NAND U24339 ( .A(n185), .B(n23577), .Z(n23579) );
  XOR U24340 ( .A(b[9]), .B(a[165]), .Z(n23732) );
  NAND U24341 ( .A(n36805), .B(n23732), .Z(n23578) );
  NAND U24342 ( .A(n23579), .B(n23578), .Z(n23657) );
  XNOR U24343 ( .A(n23658), .B(n23657), .Z(n23659) );
  XOR U24344 ( .A(n23660), .B(n23659), .Z(n23666) );
  XOR U24345 ( .A(n23665), .B(n23666), .Z(n23672) );
  XOR U24346 ( .A(n23671), .B(n23672), .Z(n23684) );
  XNOR U24347 ( .A(n23683), .B(n23684), .Z(n23741) );
  XNOR U24348 ( .A(n23742), .B(n23741), .Z(n23743) );
  XOR U24349 ( .A(n23744), .B(n23743), .Z(n23748) );
  XOR U24350 ( .A(n23747), .B(n23748), .Z(n23750) );
  XOR U24351 ( .A(n23749), .B(n23750), .Z(n23624) );
  NANDN U24352 ( .A(n23581), .B(n23580), .Z(n23585) );
  NAND U24353 ( .A(n23583), .B(n23582), .Z(n23584) );
  AND U24354 ( .A(n23585), .B(n23584), .Z(n23622) );
  NANDN U24355 ( .A(n23587), .B(n23586), .Z(n23591) );
  NANDN U24356 ( .A(n23589), .B(n23588), .Z(n23590) );
  AND U24357 ( .A(n23591), .B(n23590), .Z(n23621) );
  XNOR U24358 ( .A(n23622), .B(n23621), .Z(n23623) );
  XNOR U24359 ( .A(n23624), .B(n23623), .Z(n23615) );
  NANDN U24360 ( .A(n23593), .B(n23592), .Z(n23597) );
  NANDN U24361 ( .A(n23595), .B(n23594), .Z(n23596) );
  NAND U24362 ( .A(n23597), .B(n23596), .Z(n23616) );
  XNOR U24363 ( .A(n23615), .B(n23616), .Z(n23617) );
  NANDN U24364 ( .A(n23599), .B(n23598), .Z(n23603) );
  NAND U24365 ( .A(n23601), .B(n23600), .Z(n23602) );
  NAND U24366 ( .A(n23603), .B(n23602), .Z(n23618) );
  XNOR U24367 ( .A(n23617), .B(n23618), .Z(n23609) );
  XNOR U24368 ( .A(n23610), .B(n23609), .Z(n23611) );
  XNOR U24369 ( .A(n23612), .B(n23611), .Z(n23753) );
  XNOR U24370 ( .A(sreg[397]), .B(n23753), .Z(n23755) );
  NANDN U24371 ( .A(sreg[396]), .B(n23604), .Z(n23608) );
  NAND U24372 ( .A(n23606), .B(n23605), .Z(n23607) );
  NAND U24373 ( .A(n23608), .B(n23607), .Z(n23754) );
  XNOR U24374 ( .A(n23755), .B(n23754), .Z(c[397]) );
  NANDN U24375 ( .A(n23610), .B(n23609), .Z(n23614) );
  NANDN U24376 ( .A(n23612), .B(n23611), .Z(n23613) );
  AND U24377 ( .A(n23614), .B(n23613), .Z(n23761) );
  NANDN U24378 ( .A(n23616), .B(n23615), .Z(n23620) );
  NANDN U24379 ( .A(n23618), .B(n23617), .Z(n23619) );
  AND U24380 ( .A(n23620), .B(n23619), .Z(n23759) );
  NANDN U24381 ( .A(n23622), .B(n23621), .Z(n23626) );
  NANDN U24382 ( .A(n23624), .B(n23623), .Z(n23625) );
  AND U24383 ( .A(n23626), .B(n23625), .Z(n23767) );
  NANDN U24384 ( .A(n23628), .B(n23627), .Z(n23632) );
  NANDN U24385 ( .A(n23630), .B(n23629), .Z(n23631) );
  AND U24386 ( .A(n23632), .B(n23631), .Z(n23848) );
  NAND U24387 ( .A(n38385), .B(n23633), .Z(n23635) );
  XOR U24388 ( .A(b[27]), .B(a[148]), .Z(n23794) );
  NAND U24389 ( .A(n38343), .B(n23794), .Z(n23634) );
  AND U24390 ( .A(n23635), .B(n23634), .Z(n23855) );
  NAND U24391 ( .A(n183), .B(n23636), .Z(n23638) );
  XOR U24392 ( .A(b[5]), .B(a[170]), .Z(n23797) );
  NAND U24393 ( .A(n36296), .B(n23797), .Z(n23637) );
  AND U24394 ( .A(n23638), .B(n23637), .Z(n23853) );
  NAND U24395 ( .A(n190), .B(n23639), .Z(n23641) );
  XOR U24396 ( .A(b[19]), .B(a[156]), .Z(n23800) );
  NAND U24397 ( .A(n37821), .B(n23800), .Z(n23640) );
  NAND U24398 ( .A(n23641), .B(n23640), .Z(n23852) );
  XNOR U24399 ( .A(n23853), .B(n23852), .Z(n23854) );
  XNOR U24400 ( .A(n23855), .B(n23854), .Z(n23846) );
  NAND U24401 ( .A(n38470), .B(n23642), .Z(n23644) );
  XOR U24402 ( .A(b[31]), .B(a[144]), .Z(n23803) );
  NAND U24403 ( .A(n38453), .B(n23803), .Z(n23643) );
  AND U24404 ( .A(n23644), .B(n23643), .Z(n23815) );
  NAND U24405 ( .A(n181), .B(n23645), .Z(n23647) );
  XOR U24406 ( .A(b[3]), .B(a[172]), .Z(n23806) );
  NAND U24407 ( .A(n182), .B(n23806), .Z(n23646) );
  AND U24408 ( .A(n23647), .B(n23646), .Z(n23813) );
  NAND U24409 ( .A(n189), .B(n23648), .Z(n23650) );
  XOR U24410 ( .A(b[17]), .B(a[158]), .Z(n23809) );
  NAND U24411 ( .A(n37652), .B(n23809), .Z(n23649) );
  NAND U24412 ( .A(n23650), .B(n23649), .Z(n23812) );
  XNOR U24413 ( .A(n23813), .B(n23812), .Z(n23814) );
  XOR U24414 ( .A(n23815), .B(n23814), .Z(n23847) );
  XOR U24415 ( .A(n23846), .B(n23847), .Z(n23849) );
  XOR U24416 ( .A(n23848), .B(n23849), .Z(n23783) );
  NANDN U24417 ( .A(n23652), .B(n23651), .Z(n23656) );
  NANDN U24418 ( .A(n23654), .B(n23653), .Z(n23655) );
  AND U24419 ( .A(n23656), .B(n23655), .Z(n23836) );
  NANDN U24420 ( .A(n23658), .B(n23657), .Z(n23662) );
  NANDN U24421 ( .A(n23660), .B(n23659), .Z(n23661) );
  NAND U24422 ( .A(n23662), .B(n23661), .Z(n23837) );
  XNOR U24423 ( .A(n23836), .B(n23837), .Z(n23838) );
  NANDN U24424 ( .A(n23664), .B(n23663), .Z(n23668) );
  NANDN U24425 ( .A(n23666), .B(n23665), .Z(n23667) );
  NAND U24426 ( .A(n23668), .B(n23667), .Z(n23839) );
  XNOR U24427 ( .A(n23838), .B(n23839), .Z(n23782) );
  XNOR U24428 ( .A(n23783), .B(n23782), .Z(n23785) );
  NANDN U24429 ( .A(n23670), .B(n23669), .Z(n23674) );
  NANDN U24430 ( .A(n23672), .B(n23671), .Z(n23673) );
  AND U24431 ( .A(n23674), .B(n23673), .Z(n23784) );
  XOR U24432 ( .A(n23785), .B(n23784), .Z(n23896) );
  NANDN U24433 ( .A(n23676), .B(n23675), .Z(n23680) );
  NANDN U24434 ( .A(n23678), .B(n23677), .Z(n23679) );
  AND U24435 ( .A(n23680), .B(n23679), .Z(n23894) );
  NANDN U24436 ( .A(n23682), .B(n23681), .Z(n23686) );
  NANDN U24437 ( .A(n23684), .B(n23683), .Z(n23685) );
  AND U24438 ( .A(n23686), .B(n23685), .Z(n23779) );
  NANDN U24439 ( .A(n23688), .B(n23687), .Z(n23692) );
  OR U24440 ( .A(n23690), .B(n23689), .Z(n23691) );
  AND U24441 ( .A(n23692), .B(n23691), .Z(n23777) );
  NANDN U24442 ( .A(n23694), .B(n23693), .Z(n23698) );
  NANDN U24443 ( .A(n23696), .B(n23695), .Z(n23697) );
  AND U24444 ( .A(n23698), .B(n23697), .Z(n23843) );
  NANDN U24445 ( .A(n23700), .B(n23699), .Z(n23704) );
  NANDN U24446 ( .A(n23702), .B(n23701), .Z(n23703) );
  NAND U24447 ( .A(n23704), .B(n23703), .Z(n23842) );
  XNOR U24448 ( .A(n23843), .B(n23842), .Z(n23845) );
  NAND U24449 ( .A(b[0]), .B(a[174]), .Z(n23705) );
  XNOR U24450 ( .A(b[1]), .B(n23705), .Z(n23707) );
  NANDN U24451 ( .A(b[0]), .B(a[173]), .Z(n23706) );
  NAND U24452 ( .A(n23707), .B(n23706), .Z(n23791) );
  NAND U24453 ( .A(n194), .B(n23708), .Z(n23710) );
  XOR U24454 ( .A(b[29]), .B(a[146]), .Z(n23867) );
  NAND U24455 ( .A(n38456), .B(n23867), .Z(n23709) );
  AND U24456 ( .A(n23710), .B(n23709), .Z(n23789) );
  AND U24457 ( .A(b[31]), .B(a[142]), .Z(n23788) );
  XNOR U24458 ( .A(n23789), .B(n23788), .Z(n23790) );
  XNOR U24459 ( .A(n23791), .B(n23790), .Z(n23831) );
  NAND U24460 ( .A(n38185), .B(n23711), .Z(n23713) );
  XOR U24461 ( .A(b[23]), .B(a[152]), .Z(n23870) );
  NAND U24462 ( .A(n38132), .B(n23870), .Z(n23712) );
  AND U24463 ( .A(n23713), .B(n23712), .Z(n23860) );
  NAND U24464 ( .A(n184), .B(n23714), .Z(n23716) );
  XOR U24465 ( .A(b[7]), .B(a[168]), .Z(n23873) );
  NAND U24466 ( .A(n36592), .B(n23873), .Z(n23715) );
  AND U24467 ( .A(n23716), .B(n23715), .Z(n23859) );
  NAND U24468 ( .A(n38289), .B(n23717), .Z(n23719) );
  XOR U24469 ( .A(b[25]), .B(a[150]), .Z(n23876) );
  NAND U24470 ( .A(n38247), .B(n23876), .Z(n23718) );
  NAND U24471 ( .A(n23719), .B(n23718), .Z(n23858) );
  XOR U24472 ( .A(n23859), .B(n23858), .Z(n23861) );
  XOR U24473 ( .A(n23860), .B(n23861), .Z(n23830) );
  XOR U24474 ( .A(n23831), .B(n23830), .Z(n23833) );
  NAND U24475 ( .A(n187), .B(n23720), .Z(n23722) );
  XOR U24476 ( .A(b[13]), .B(a[162]), .Z(n23879) );
  NAND U24477 ( .A(n37295), .B(n23879), .Z(n23721) );
  AND U24478 ( .A(n23722), .B(n23721), .Z(n23825) );
  NAND U24479 ( .A(n186), .B(n23723), .Z(n23725) );
  XOR U24480 ( .A(b[11]), .B(a[164]), .Z(n23882) );
  NAND U24481 ( .A(n37097), .B(n23882), .Z(n23724) );
  NAND U24482 ( .A(n23725), .B(n23724), .Z(n23824) );
  XNOR U24483 ( .A(n23825), .B(n23824), .Z(n23827) );
  NAND U24484 ( .A(n188), .B(n23726), .Z(n23728) );
  XOR U24485 ( .A(b[15]), .B(a[160]), .Z(n23885) );
  NAND U24486 ( .A(n37382), .B(n23885), .Z(n23727) );
  AND U24487 ( .A(n23728), .B(n23727), .Z(n23821) );
  NAND U24488 ( .A(n38064), .B(n23729), .Z(n23731) );
  XOR U24489 ( .A(b[21]), .B(a[154]), .Z(n23888) );
  NAND U24490 ( .A(n37993), .B(n23888), .Z(n23730) );
  AND U24491 ( .A(n23731), .B(n23730), .Z(n23819) );
  NAND U24492 ( .A(n185), .B(n23732), .Z(n23734) );
  XOR U24493 ( .A(b[9]), .B(a[166]), .Z(n23891) );
  NAND U24494 ( .A(n36805), .B(n23891), .Z(n23733) );
  NAND U24495 ( .A(n23734), .B(n23733), .Z(n23818) );
  XNOR U24496 ( .A(n23819), .B(n23818), .Z(n23820) );
  XNOR U24497 ( .A(n23821), .B(n23820), .Z(n23826) );
  XOR U24498 ( .A(n23827), .B(n23826), .Z(n23832) );
  XNOR U24499 ( .A(n23833), .B(n23832), .Z(n23844) );
  XNOR U24500 ( .A(n23845), .B(n23844), .Z(n23776) );
  XNOR U24501 ( .A(n23777), .B(n23776), .Z(n23778) );
  XOR U24502 ( .A(n23779), .B(n23778), .Z(n23895) );
  XOR U24503 ( .A(n23894), .B(n23895), .Z(n23897) );
  XOR U24504 ( .A(n23896), .B(n23897), .Z(n23773) );
  NANDN U24505 ( .A(n23736), .B(n23735), .Z(n23740) );
  NAND U24506 ( .A(n23738), .B(n23737), .Z(n23739) );
  AND U24507 ( .A(n23740), .B(n23739), .Z(n23771) );
  NANDN U24508 ( .A(n23742), .B(n23741), .Z(n23746) );
  NANDN U24509 ( .A(n23744), .B(n23743), .Z(n23745) );
  AND U24510 ( .A(n23746), .B(n23745), .Z(n23770) );
  XNOR U24511 ( .A(n23771), .B(n23770), .Z(n23772) );
  XNOR U24512 ( .A(n23773), .B(n23772), .Z(n23764) );
  NANDN U24513 ( .A(n23748), .B(n23747), .Z(n23752) );
  OR U24514 ( .A(n23750), .B(n23749), .Z(n23751) );
  NAND U24515 ( .A(n23752), .B(n23751), .Z(n23765) );
  XNOR U24516 ( .A(n23764), .B(n23765), .Z(n23766) );
  XNOR U24517 ( .A(n23767), .B(n23766), .Z(n23758) );
  XNOR U24518 ( .A(n23759), .B(n23758), .Z(n23760) );
  XNOR U24519 ( .A(n23761), .B(n23760), .Z(n23900) );
  XNOR U24520 ( .A(sreg[398]), .B(n23900), .Z(n23902) );
  NANDN U24521 ( .A(sreg[397]), .B(n23753), .Z(n23757) );
  NAND U24522 ( .A(n23755), .B(n23754), .Z(n23756) );
  NAND U24523 ( .A(n23757), .B(n23756), .Z(n23901) );
  XNOR U24524 ( .A(n23902), .B(n23901), .Z(c[398]) );
  NANDN U24525 ( .A(n23759), .B(n23758), .Z(n23763) );
  NANDN U24526 ( .A(n23761), .B(n23760), .Z(n23762) );
  AND U24527 ( .A(n23763), .B(n23762), .Z(n23908) );
  NANDN U24528 ( .A(n23765), .B(n23764), .Z(n23769) );
  NANDN U24529 ( .A(n23767), .B(n23766), .Z(n23768) );
  AND U24530 ( .A(n23769), .B(n23768), .Z(n23906) );
  NANDN U24531 ( .A(n23771), .B(n23770), .Z(n23775) );
  NANDN U24532 ( .A(n23773), .B(n23772), .Z(n23774) );
  AND U24533 ( .A(n23775), .B(n23774), .Z(n23914) );
  NANDN U24534 ( .A(n23777), .B(n23776), .Z(n23781) );
  NANDN U24535 ( .A(n23779), .B(n23778), .Z(n23780) );
  AND U24536 ( .A(n23781), .B(n23780), .Z(n23918) );
  NANDN U24537 ( .A(n23783), .B(n23782), .Z(n23787) );
  NAND U24538 ( .A(n23785), .B(n23784), .Z(n23786) );
  AND U24539 ( .A(n23787), .B(n23786), .Z(n23917) );
  XNOR U24540 ( .A(n23918), .B(n23917), .Z(n23920) );
  NANDN U24541 ( .A(n23789), .B(n23788), .Z(n23793) );
  NANDN U24542 ( .A(n23791), .B(n23790), .Z(n23792) );
  AND U24543 ( .A(n23793), .B(n23792), .Z(n23985) );
  NAND U24544 ( .A(n38385), .B(n23794), .Z(n23796) );
  XOR U24545 ( .A(b[27]), .B(a[149]), .Z(n23929) );
  NAND U24546 ( .A(n38343), .B(n23929), .Z(n23795) );
  AND U24547 ( .A(n23796), .B(n23795), .Z(n23992) );
  NAND U24548 ( .A(n183), .B(n23797), .Z(n23799) );
  XOR U24549 ( .A(b[5]), .B(a[171]), .Z(n23932) );
  NAND U24550 ( .A(n36296), .B(n23932), .Z(n23798) );
  AND U24551 ( .A(n23799), .B(n23798), .Z(n23990) );
  NAND U24552 ( .A(n190), .B(n23800), .Z(n23802) );
  XOR U24553 ( .A(b[19]), .B(a[157]), .Z(n23935) );
  NAND U24554 ( .A(n37821), .B(n23935), .Z(n23801) );
  NAND U24555 ( .A(n23802), .B(n23801), .Z(n23989) );
  XNOR U24556 ( .A(n23990), .B(n23989), .Z(n23991) );
  XNOR U24557 ( .A(n23992), .B(n23991), .Z(n23983) );
  NAND U24558 ( .A(n38470), .B(n23803), .Z(n23805) );
  XOR U24559 ( .A(b[31]), .B(a[145]), .Z(n23938) );
  NAND U24560 ( .A(n38453), .B(n23938), .Z(n23804) );
  AND U24561 ( .A(n23805), .B(n23804), .Z(n23950) );
  NAND U24562 ( .A(n181), .B(n23806), .Z(n23808) );
  XOR U24563 ( .A(b[3]), .B(a[173]), .Z(n23941) );
  NAND U24564 ( .A(n182), .B(n23941), .Z(n23807) );
  AND U24565 ( .A(n23808), .B(n23807), .Z(n23948) );
  NAND U24566 ( .A(n189), .B(n23809), .Z(n23811) );
  XOR U24567 ( .A(b[17]), .B(a[159]), .Z(n23944) );
  NAND U24568 ( .A(n37652), .B(n23944), .Z(n23810) );
  NAND U24569 ( .A(n23811), .B(n23810), .Z(n23947) );
  XNOR U24570 ( .A(n23948), .B(n23947), .Z(n23949) );
  XOR U24571 ( .A(n23950), .B(n23949), .Z(n23984) );
  XOR U24572 ( .A(n23983), .B(n23984), .Z(n23986) );
  XOR U24573 ( .A(n23985), .B(n23986), .Z(n24032) );
  NANDN U24574 ( .A(n23813), .B(n23812), .Z(n23817) );
  NANDN U24575 ( .A(n23815), .B(n23814), .Z(n23816) );
  AND U24576 ( .A(n23817), .B(n23816), .Z(n23971) );
  NANDN U24577 ( .A(n23819), .B(n23818), .Z(n23823) );
  NANDN U24578 ( .A(n23821), .B(n23820), .Z(n23822) );
  NAND U24579 ( .A(n23823), .B(n23822), .Z(n23972) );
  XNOR U24580 ( .A(n23971), .B(n23972), .Z(n23973) );
  NANDN U24581 ( .A(n23825), .B(n23824), .Z(n23829) );
  NAND U24582 ( .A(n23827), .B(n23826), .Z(n23828) );
  NAND U24583 ( .A(n23829), .B(n23828), .Z(n23974) );
  XNOR U24584 ( .A(n23973), .B(n23974), .Z(n24031) );
  XNOR U24585 ( .A(n24032), .B(n24031), .Z(n24034) );
  NAND U24586 ( .A(n23831), .B(n23830), .Z(n23835) );
  NAND U24587 ( .A(n23833), .B(n23832), .Z(n23834) );
  AND U24588 ( .A(n23835), .B(n23834), .Z(n24033) );
  XOR U24589 ( .A(n24034), .B(n24033), .Z(n24046) );
  NANDN U24590 ( .A(n23837), .B(n23836), .Z(n23841) );
  NANDN U24591 ( .A(n23839), .B(n23838), .Z(n23840) );
  AND U24592 ( .A(n23841), .B(n23840), .Z(n24043) );
  NANDN U24593 ( .A(n23847), .B(n23846), .Z(n23851) );
  OR U24594 ( .A(n23849), .B(n23848), .Z(n23850) );
  AND U24595 ( .A(n23851), .B(n23850), .Z(n24038) );
  NANDN U24596 ( .A(n23853), .B(n23852), .Z(n23857) );
  NANDN U24597 ( .A(n23855), .B(n23854), .Z(n23856) );
  AND U24598 ( .A(n23857), .B(n23856), .Z(n23978) );
  NANDN U24599 ( .A(n23859), .B(n23858), .Z(n23863) );
  OR U24600 ( .A(n23861), .B(n23860), .Z(n23862) );
  NAND U24601 ( .A(n23863), .B(n23862), .Z(n23977) );
  XNOR U24602 ( .A(n23978), .B(n23977), .Z(n23979) );
  NAND U24603 ( .A(b[0]), .B(a[175]), .Z(n23864) );
  XNOR U24604 ( .A(b[1]), .B(n23864), .Z(n23866) );
  NANDN U24605 ( .A(b[0]), .B(a[174]), .Z(n23865) );
  NAND U24606 ( .A(n23866), .B(n23865), .Z(n23926) );
  NAND U24607 ( .A(n194), .B(n23867), .Z(n23869) );
  XOR U24608 ( .A(b[29]), .B(a[147]), .Z(n24001) );
  NAND U24609 ( .A(n38456), .B(n24001), .Z(n23868) );
  AND U24610 ( .A(n23869), .B(n23868), .Z(n23924) );
  AND U24611 ( .A(b[31]), .B(a[143]), .Z(n23923) );
  XNOR U24612 ( .A(n23924), .B(n23923), .Z(n23925) );
  XNOR U24613 ( .A(n23926), .B(n23925), .Z(n23965) );
  NAND U24614 ( .A(n38185), .B(n23870), .Z(n23872) );
  XOR U24615 ( .A(b[23]), .B(a[153]), .Z(n24007) );
  NAND U24616 ( .A(n38132), .B(n24007), .Z(n23871) );
  AND U24617 ( .A(n23872), .B(n23871), .Z(n23998) );
  NAND U24618 ( .A(n184), .B(n23873), .Z(n23875) );
  XOR U24619 ( .A(b[7]), .B(a[169]), .Z(n24010) );
  NAND U24620 ( .A(n36592), .B(n24010), .Z(n23874) );
  AND U24621 ( .A(n23875), .B(n23874), .Z(n23996) );
  NAND U24622 ( .A(n38289), .B(n23876), .Z(n23878) );
  XOR U24623 ( .A(b[25]), .B(a[151]), .Z(n24013) );
  NAND U24624 ( .A(n38247), .B(n24013), .Z(n23877) );
  NAND U24625 ( .A(n23878), .B(n23877), .Z(n23995) );
  XNOR U24626 ( .A(n23996), .B(n23995), .Z(n23997) );
  XOR U24627 ( .A(n23998), .B(n23997), .Z(n23966) );
  XNOR U24628 ( .A(n23965), .B(n23966), .Z(n23967) );
  NAND U24629 ( .A(n187), .B(n23879), .Z(n23881) );
  XOR U24630 ( .A(b[13]), .B(a[163]), .Z(n24016) );
  NAND U24631 ( .A(n37295), .B(n24016), .Z(n23880) );
  AND U24632 ( .A(n23881), .B(n23880), .Z(n23960) );
  NAND U24633 ( .A(n186), .B(n23882), .Z(n23884) );
  XOR U24634 ( .A(b[11]), .B(a[165]), .Z(n24019) );
  NAND U24635 ( .A(n37097), .B(n24019), .Z(n23883) );
  NAND U24636 ( .A(n23884), .B(n23883), .Z(n23959) );
  XNOR U24637 ( .A(n23960), .B(n23959), .Z(n23961) );
  NAND U24638 ( .A(n188), .B(n23885), .Z(n23887) );
  XOR U24639 ( .A(b[15]), .B(a[161]), .Z(n24022) );
  NAND U24640 ( .A(n37382), .B(n24022), .Z(n23886) );
  AND U24641 ( .A(n23887), .B(n23886), .Z(n23956) );
  NAND U24642 ( .A(n38064), .B(n23888), .Z(n23890) );
  XOR U24643 ( .A(b[21]), .B(a[155]), .Z(n24025) );
  NAND U24644 ( .A(n37993), .B(n24025), .Z(n23889) );
  AND U24645 ( .A(n23890), .B(n23889), .Z(n23954) );
  NAND U24646 ( .A(n185), .B(n23891), .Z(n23893) );
  XOR U24647 ( .A(b[9]), .B(a[167]), .Z(n24028) );
  NAND U24648 ( .A(n36805), .B(n24028), .Z(n23892) );
  NAND U24649 ( .A(n23893), .B(n23892), .Z(n23953) );
  XNOR U24650 ( .A(n23954), .B(n23953), .Z(n23955) );
  XOR U24651 ( .A(n23956), .B(n23955), .Z(n23962) );
  XOR U24652 ( .A(n23961), .B(n23962), .Z(n23968) );
  XOR U24653 ( .A(n23967), .B(n23968), .Z(n23980) );
  XNOR U24654 ( .A(n23979), .B(n23980), .Z(n24037) );
  XNOR U24655 ( .A(n24038), .B(n24037), .Z(n24039) );
  XOR U24656 ( .A(n24040), .B(n24039), .Z(n24044) );
  XNOR U24657 ( .A(n24043), .B(n24044), .Z(n24045) );
  XNOR U24658 ( .A(n24046), .B(n24045), .Z(n23919) );
  XOR U24659 ( .A(n23920), .B(n23919), .Z(n23912) );
  NANDN U24660 ( .A(n23895), .B(n23894), .Z(n23899) );
  OR U24661 ( .A(n23897), .B(n23896), .Z(n23898) );
  AND U24662 ( .A(n23899), .B(n23898), .Z(n23911) );
  XNOR U24663 ( .A(n23912), .B(n23911), .Z(n23913) );
  XNOR U24664 ( .A(n23914), .B(n23913), .Z(n23905) );
  XNOR U24665 ( .A(n23906), .B(n23905), .Z(n23907) );
  XNOR U24666 ( .A(n23908), .B(n23907), .Z(n24049) );
  XNOR U24667 ( .A(sreg[399]), .B(n24049), .Z(n24051) );
  NANDN U24668 ( .A(sreg[398]), .B(n23900), .Z(n23904) );
  NAND U24669 ( .A(n23902), .B(n23901), .Z(n23903) );
  NAND U24670 ( .A(n23904), .B(n23903), .Z(n24050) );
  XNOR U24671 ( .A(n24051), .B(n24050), .Z(c[399]) );
  NANDN U24672 ( .A(n23906), .B(n23905), .Z(n23910) );
  NANDN U24673 ( .A(n23908), .B(n23907), .Z(n23909) );
  AND U24674 ( .A(n23910), .B(n23909), .Z(n24057) );
  NANDN U24675 ( .A(n23912), .B(n23911), .Z(n23916) );
  NANDN U24676 ( .A(n23914), .B(n23913), .Z(n23915) );
  AND U24677 ( .A(n23916), .B(n23915), .Z(n24055) );
  NANDN U24678 ( .A(n23918), .B(n23917), .Z(n23922) );
  NAND U24679 ( .A(n23920), .B(n23919), .Z(n23921) );
  AND U24680 ( .A(n23922), .B(n23921), .Z(n24062) );
  NANDN U24681 ( .A(n23924), .B(n23923), .Z(n23928) );
  NANDN U24682 ( .A(n23926), .B(n23925), .Z(n23927) );
  AND U24683 ( .A(n23928), .B(n23927), .Z(n24144) );
  NAND U24684 ( .A(n38385), .B(n23929), .Z(n23931) );
  XOR U24685 ( .A(b[27]), .B(a[150]), .Z(n24090) );
  NAND U24686 ( .A(n38343), .B(n24090), .Z(n23930) );
  AND U24687 ( .A(n23931), .B(n23930), .Z(n24151) );
  NAND U24688 ( .A(n183), .B(n23932), .Z(n23934) );
  XOR U24689 ( .A(b[5]), .B(a[172]), .Z(n24093) );
  NAND U24690 ( .A(n36296), .B(n24093), .Z(n23933) );
  AND U24691 ( .A(n23934), .B(n23933), .Z(n24149) );
  NAND U24692 ( .A(n190), .B(n23935), .Z(n23937) );
  XOR U24693 ( .A(b[19]), .B(a[158]), .Z(n24096) );
  NAND U24694 ( .A(n37821), .B(n24096), .Z(n23936) );
  NAND U24695 ( .A(n23937), .B(n23936), .Z(n24148) );
  XNOR U24696 ( .A(n24149), .B(n24148), .Z(n24150) );
  XNOR U24697 ( .A(n24151), .B(n24150), .Z(n24142) );
  NAND U24698 ( .A(n38470), .B(n23938), .Z(n23940) );
  XOR U24699 ( .A(b[31]), .B(a[146]), .Z(n24099) );
  NAND U24700 ( .A(n38453), .B(n24099), .Z(n23939) );
  AND U24701 ( .A(n23940), .B(n23939), .Z(n24111) );
  NAND U24702 ( .A(n181), .B(n23941), .Z(n23943) );
  XOR U24703 ( .A(b[3]), .B(a[174]), .Z(n24102) );
  NAND U24704 ( .A(n182), .B(n24102), .Z(n23942) );
  AND U24705 ( .A(n23943), .B(n23942), .Z(n24109) );
  NAND U24706 ( .A(n189), .B(n23944), .Z(n23946) );
  XOR U24707 ( .A(b[17]), .B(a[160]), .Z(n24105) );
  NAND U24708 ( .A(n37652), .B(n24105), .Z(n23945) );
  NAND U24709 ( .A(n23946), .B(n23945), .Z(n24108) );
  XNOR U24710 ( .A(n24109), .B(n24108), .Z(n24110) );
  XOR U24711 ( .A(n24111), .B(n24110), .Z(n24143) );
  XOR U24712 ( .A(n24142), .B(n24143), .Z(n24145) );
  XOR U24713 ( .A(n24144), .B(n24145), .Z(n24079) );
  NANDN U24714 ( .A(n23948), .B(n23947), .Z(n23952) );
  NANDN U24715 ( .A(n23950), .B(n23949), .Z(n23951) );
  AND U24716 ( .A(n23952), .B(n23951), .Z(n24132) );
  NANDN U24717 ( .A(n23954), .B(n23953), .Z(n23958) );
  NANDN U24718 ( .A(n23956), .B(n23955), .Z(n23957) );
  NAND U24719 ( .A(n23958), .B(n23957), .Z(n24133) );
  XNOR U24720 ( .A(n24132), .B(n24133), .Z(n24134) );
  NANDN U24721 ( .A(n23960), .B(n23959), .Z(n23964) );
  NANDN U24722 ( .A(n23962), .B(n23961), .Z(n23963) );
  NAND U24723 ( .A(n23964), .B(n23963), .Z(n24135) );
  XNOR U24724 ( .A(n24134), .B(n24135), .Z(n24078) );
  XNOR U24725 ( .A(n24079), .B(n24078), .Z(n24081) );
  NANDN U24726 ( .A(n23966), .B(n23965), .Z(n23970) );
  NANDN U24727 ( .A(n23968), .B(n23967), .Z(n23969) );
  AND U24728 ( .A(n23970), .B(n23969), .Z(n24080) );
  XOR U24729 ( .A(n24081), .B(n24080), .Z(n24192) );
  NANDN U24730 ( .A(n23972), .B(n23971), .Z(n23976) );
  NANDN U24731 ( .A(n23974), .B(n23973), .Z(n23975) );
  AND U24732 ( .A(n23976), .B(n23975), .Z(n24190) );
  NANDN U24733 ( .A(n23978), .B(n23977), .Z(n23982) );
  NANDN U24734 ( .A(n23980), .B(n23979), .Z(n23981) );
  AND U24735 ( .A(n23982), .B(n23981), .Z(n24075) );
  NANDN U24736 ( .A(n23984), .B(n23983), .Z(n23988) );
  OR U24737 ( .A(n23986), .B(n23985), .Z(n23987) );
  AND U24738 ( .A(n23988), .B(n23987), .Z(n24073) );
  NANDN U24739 ( .A(n23990), .B(n23989), .Z(n23994) );
  NANDN U24740 ( .A(n23992), .B(n23991), .Z(n23993) );
  AND U24741 ( .A(n23994), .B(n23993), .Z(n24139) );
  NANDN U24742 ( .A(n23996), .B(n23995), .Z(n24000) );
  NANDN U24743 ( .A(n23998), .B(n23997), .Z(n23999) );
  NAND U24744 ( .A(n24000), .B(n23999), .Z(n24138) );
  XNOR U24745 ( .A(n24139), .B(n24138), .Z(n24141) );
  NAND U24746 ( .A(n194), .B(n24001), .Z(n24003) );
  XOR U24747 ( .A(b[29]), .B(a[148]), .Z(n24163) );
  NAND U24748 ( .A(n38456), .B(n24163), .Z(n24002) );
  AND U24749 ( .A(n24003), .B(n24002), .Z(n24085) );
  AND U24750 ( .A(b[31]), .B(a[144]), .Z(n24084) );
  XNOR U24751 ( .A(n24085), .B(n24084), .Z(n24086) );
  NAND U24752 ( .A(b[0]), .B(a[176]), .Z(n24004) );
  XNOR U24753 ( .A(b[1]), .B(n24004), .Z(n24006) );
  NANDN U24754 ( .A(b[0]), .B(a[175]), .Z(n24005) );
  NAND U24755 ( .A(n24006), .B(n24005), .Z(n24087) );
  XNOR U24756 ( .A(n24086), .B(n24087), .Z(n24127) );
  NAND U24757 ( .A(n38185), .B(n24007), .Z(n24009) );
  XOR U24758 ( .A(b[23]), .B(a[154]), .Z(n24166) );
  NAND U24759 ( .A(n38132), .B(n24166), .Z(n24008) );
  AND U24760 ( .A(n24009), .B(n24008), .Z(n24156) );
  NAND U24761 ( .A(n184), .B(n24010), .Z(n24012) );
  XOR U24762 ( .A(b[7]), .B(a[170]), .Z(n24169) );
  NAND U24763 ( .A(n36592), .B(n24169), .Z(n24011) );
  AND U24764 ( .A(n24012), .B(n24011), .Z(n24155) );
  NAND U24765 ( .A(n38289), .B(n24013), .Z(n24015) );
  XOR U24766 ( .A(b[25]), .B(a[152]), .Z(n24172) );
  NAND U24767 ( .A(n38247), .B(n24172), .Z(n24014) );
  NAND U24768 ( .A(n24015), .B(n24014), .Z(n24154) );
  XOR U24769 ( .A(n24155), .B(n24154), .Z(n24157) );
  XOR U24770 ( .A(n24156), .B(n24157), .Z(n24126) );
  XOR U24771 ( .A(n24127), .B(n24126), .Z(n24129) );
  NAND U24772 ( .A(n187), .B(n24016), .Z(n24018) );
  XOR U24773 ( .A(b[13]), .B(a[164]), .Z(n24175) );
  NAND U24774 ( .A(n37295), .B(n24175), .Z(n24017) );
  AND U24775 ( .A(n24018), .B(n24017), .Z(n24121) );
  NAND U24776 ( .A(n186), .B(n24019), .Z(n24021) );
  XOR U24777 ( .A(b[11]), .B(a[166]), .Z(n24178) );
  NAND U24778 ( .A(n37097), .B(n24178), .Z(n24020) );
  NAND U24779 ( .A(n24021), .B(n24020), .Z(n24120) );
  XNOR U24780 ( .A(n24121), .B(n24120), .Z(n24123) );
  NAND U24781 ( .A(n188), .B(n24022), .Z(n24024) );
  XOR U24782 ( .A(b[15]), .B(a[162]), .Z(n24181) );
  NAND U24783 ( .A(n37382), .B(n24181), .Z(n24023) );
  AND U24784 ( .A(n24024), .B(n24023), .Z(n24117) );
  NAND U24785 ( .A(n38064), .B(n24025), .Z(n24027) );
  XOR U24786 ( .A(b[21]), .B(a[156]), .Z(n24184) );
  NAND U24787 ( .A(n37993), .B(n24184), .Z(n24026) );
  AND U24788 ( .A(n24027), .B(n24026), .Z(n24115) );
  NAND U24789 ( .A(n185), .B(n24028), .Z(n24030) );
  XOR U24790 ( .A(b[9]), .B(a[168]), .Z(n24187) );
  NAND U24791 ( .A(n36805), .B(n24187), .Z(n24029) );
  NAND U24792 ( .A(n24030), .B(n24029), .Z(n24114) );
  XNOR U24793 ( .A(n24115), .B(n24114), .Z(n24116) );
  XNOR U24794 ( .A(n24117), .B(n24116), .Z(n24122) );
  XOR U24795 ( .A(n24123), .B(n24122), .Z(n24128) );
  XNOR U24796 ( .A(n24129), .B(n24128), .Z(n24140) );
  XNOR U24797 ( .A(n24141), .B(n24140), .Z(n24072) );
  XNOR U24798 ( .A(n24073), .B(n24072), .Z(n24074) );
  XOR U24799 ( .A(n24075), .B(n24074), .Z(n24191) );
  XOR U24800 ( .A(n24190), .B(n24191), .Z(n24193) );
  XOR U24801 ( .A(n24192), .B(n24193), .Z(n24069) );
  NANDN U24802 ( .A(n24032), .B(n24031), .Z(n24036) );
  NAND U24803 ( .A(n24034), .B(n24033), .Z(n24035) );
  AND U24804 ( .A(n24036), .B(n24035), .Z(n24067) );
  NANDN U24805 ( .A(n24038), .B(n24037), .Z(n24042) );
  NANDN U24806 ( .A(n24040), .B(n24039), .Z(n24041) );
  AND U24807 ( .A(n24042), .B(n24041), .Z(n24066) );
  XNOR U24808 ( .A(n24067), .B(n24066), .Z(n24068) );
  XNOR U24809 ( .A(n24069), .B(n24068), .Z(n24060) );
  NANDN U24810 ( .A(n24044), .B(n24043), .Z(n24048) );
  NANDN U24811 ( .A(n24046), .B(n24045), .Z(n24047) );
  NAND U24812 ( .A(n24048), .B(n24047), .Z(n24061) );
  XOR U24813 ( .A(n24060), .B(n24061), .Z(n24063) );
  XNOR U24814 ( .A(n24062), .B(n24063), .Z(n24054) );
  XNOR U24815 ( .A(n24055), .B(n24054), .Z(n24056) );
  XNOR U24816 ( .A(n24057), .B(n24056), .Z(n24196) );
  XNOR U24817 ( .A(sreg[400]), .B(n24196), .Z(n24198) );
  NANDN U24818 ( .A(sreg[399]), .B(n24049), .Z(n24053) );
  NAND U24819 ( .A(n24051), .B(n24050), .Z(n24052) );
  NAND U24820 ( .A(n24053), .B(n24052), .Z(n24197) );
  XNOR U24821 ( .A(n24198), .B(n24197), .Z(c[400]) );
  NANDN U24822 ( .A(n24055), .B(n24054), .Z(n24059) );
  NANDN U24823 ( .A(n24057), .B(n24056), .Z(n24058) );
  AND U24824 ( .A(n24059), .B(n24058), .Z(n24204) );
  NANDN U24825 ( .A(n24061), .B(n24060), .Z(n24065) );
  NANDN U24826 ( .A(n24063), .B(n24062), .Z(n24064) );
  AND U24827 ( .A(n24065), .B(n24064), .Z(n24202) );
  NANDN U24828 ( .A(n24067), .B(n24066), .Z(n24071) );
  NANDN U24829 ( .A(n24069), .B(n24068), .Z(n24070) );
  AND U24830 ( .A(n24071), .B(n24070), .Z(n24210) );
  NANDN U24831 ( .A(n24073), .B(n24072), .Z(n24077) );
  NANDN U24832 ( .A(n24075), .B(n24074), .Z(n24076) );
  AND U24833 ( .A(n24077), .B(n24076), .Z(n24338) );
  NANDN U24834 ( .A(n24079), .B(n24078), .Z(n24083) );
  NAND U24835 ( .A(n24081), .B(n24080), .Z(n24082) );
  AND U24836 ( .A(n24083), .B(n24082), .Z(n24337) );
  XNOR U24837 ( .A(n24338), .B(n24337), .Z(n24340) );
  NANDN U24838 ( .A(n24085), .B(n24084), .Z(n24089) );
  NANDN U24839 ( .A(n24087), .B(n24086), .Z(n24088) );
  AND U24840 ( .A(n24089), .B(n24088), .Z(n24273) );
  NAND U24841 ( .A(n38385), .B(n24090), .Z(n24092) );
  XOR U24842 ( .A(b[27]), .B(a[151]), .Z(n24219) );
  NAND U24843 ( .A(n38343), .B(n24219), .Z(n24091) );
  AND U24844 ( .A(n24092), .B(n24091), .Z(n24280) );
  NAND U24845 ( .A(n183), .B(n24093), .Z(n24095) );
  XOR U24846 ( .A(b[5]), .B(a[173]), .Z(n24222) );
  NAND U24847 ( .A(n36296), .B(n24222), .Z(n24094) );
  AND U24848 ( .A(n24095), .B(n24094), .Z(n24278) );
  NAND U24849 ( .A(n190), .B(n24096), .Z(n24098) );
  XOR U24850 ( .A(b[19]), .B(a[159]), .Z(n24225) );
  NAND U24851 ( .A(n37821), .B(n24225), .Z(n24097) );
  NAND U24852 ( .A(n24098), .B(n24097), .Z(n24277) );
  XNOR U24853 ( .A(n24278), .B(n24277), .Z(n24279) );
  XNOR U24854 ( .A(n24280), .B(n24279), .Z(n24271) );
  NAND U24855 ( .A(n38470), .B(n24099), .Z(n24101) );
  XOR U24856 ( .A(b[31]), .B(a[147]), .Z(n24228) );
  NAND U24857 ( .A(n38453), .B(n24228), .Z(n24100) );
  AND U24858 ( .A(n24101), .B(n24100), .Z(n24240) );
  NAND U24859 ( .A(n181), .B(n24102), .Z(n24104) );
  XOR U24860 ( .A(b[3]), .B(a[175]), .Z(n24231) );
  NAND U24861 ( .A(n182), .B(n24231), .Z(n24103) );
  AND U24862 ( .A(n24104), .B(n24103), .Z(n24238) );
  NAND U24863 ( .A(n189), .B(n24105), .Z(n24107) );
  XOR U24864 ( .A(b[17]), .B(a[161]), .Z(n24234) );
  NAND U24865 ( .A(n37652), .B(n24234), .Z(n24106) );
  NAND U24866 ( .A(n24107), .B(n24106), .Z(n24237) );
  XNOR U24867 ( .A(n24238), .B(n24237), .Z(n24239) );
  XOR U24868 ( .A(n24240), .B(n24239), .Z(n24272) );
  XOR U24869 ( .A(n24271), .B(n24272), .Z(n24274) );
  XOR U24870 ( .A(n24273), .B(n24274), .Z(n24320) );
  NANDN U24871 ( .A(n24109), .B(n24108), .Z(n24113) );
  NANDN U24872 ( .A(n24111), .B(n24110), .Z(n24112) );
  AND U24873 ( .A(n24113), .B(n24112), .Z(n24261) );
  NANDN U24874 ( .A(n24115), .B(n24114), .Z(n24119) );
  NANDN U24875 ( .A(n24117), .B(n24116), .Z(n24118) );
  NAND U24876 ( .A(n24119), .B(n24118), .Z(n24262) );
  XNOR U24877 ( .A(n24261), .B(n24262), .Z(n24263) );
  NANDN U24878 ( .A(n24121), .B(n24120), .Z(n24125) );
  NAND U24879 ( .A(n24123), .B(n24122), .Z(n24124) );
  NAND U24880 ( .A(n24125), .B(n24124), .Z(n24264) );
  XNOR U24881 ( .A(n24263), .B(n24264), .Z(n24319) );
  XNOR U24882 ( .A(n24320), .B(n24319), .Z(n24322) );
  NAND U24883 ( .A(n24127), .B(n24126), .Z(n24131) );
  NAND U24884 ( .A(n24129), .B(n24128), .Z(n24130) );
  AND U24885 ( .A(n24131), .B(n24130), .Z(n24321) );
  XOR U24886 ( .A(n24322), .B(n24321), .Z(n24334) );
  NANDN U24887 ( .A(n24133), .B(n24132), .Z(n24137) );
  NANDN U24888 ( .A(n24135), .B(n24134), .Z(n24136) );
  AND U24889 ( .A(n24137), .B(n24136), .Z(n24331) );
  NANDN U24890 ( .A(n24143), .B(n24142), .Z(n24147) );
  OR U24891 ( .A(n24145), .B(n24144), .Z(n24146) );
  AND U24892 ( .A(n24147), .B(n24146), .Z(n24326) );
  NANDN U24893 ( .A(n24149), .B(n24148), .Z(n24153) );
  NANDN U24894 ( .A(n24151), .B(n24150), .Z(n24152) );
  AND U24895 ( .A(n24153), .B(n24152), .Z(n24268) );
  NANDN U24896 ( .A(n24155), .B(n24154), .Z(n24159) );
  OR U24897 ( .A(n24157), .B(n24156), .Z(n24158) );
  NAND U24898 ( .A(n24159), .B(n24158), .Z(n24267) );
  XNOR U24899 ( .A(n24268), .B(n24267), .Z(n24270) );
  NAND U24900 ( .A(b[0]), .B(a[177]), .Z(n24160) );
  XNOR U24901 ( .A(b[1]), .B(n24160), .Z(n24162) );
  NANDN U24902 ( .A(b[0]), .B(a[176]), .Z(n24161) );
  NAND U24903 ( .A(n24162), .B(n24161), .Z(n24216) );
  NAND U24904 ( .A(n194), .B(n24163), .Z(n24165) );
  XOR U24905 ( .A(b[29]), .B(a[149]), .Z(n24289) );
  NAND U24906 ( .A(n38456), .B(n24289), .Z(n24164) );
  AND U24907 ( .A(n24165), .B(n24164), .Z(n24214) );
  AND U24908 ( .A(b[31]), .B(a[145]), .Z(n24213) );
  XNOR U24909 ( .A(n24214), .B(n24213), .Z(n24215) );
  XNOR U24910 ( .A(n24216), .B(n24215), .Z(n24256) );
  NAND U24911 ( .A(n38185), .B(n24166), .Z(n24168) );
  XOR U24912 ( .A(b[23]), .B(a[155]), .Z(n24295) );
  NAND U24913 ( .A(n38132), .B(n24295), .Z(n24167) );
  AND U24914 ( .A(n24168), .B(n24167), .Z(n24285) );
  NAND U24915 ( .A(n184), .B(n24169), .Z(n24171) );
  XOR U24916 ( .A(b[7]), .B(a[171]), .Z(n24298) );
  NAND U24917 ( .A(n36592), .B(n24298), .Z(n24170) );
  AND U24918 ( .A(n24171), .B(n24170), .Z(n24284) );
  NAND U24919 ( .A(n38289), .B(n24172), .Z(n24174) );
  XOR U24920 ( .A(b[25]), .B(a[153]), .Z(n24301) );
  NAND U24921 ( .A(n38247), .B(n24301), .Z(n24173) );
  NAND U24922 ( .A(n24174), .B(n24173), .Z(n24283) );
  XOR U24923 ( .A(n24284), .B(n24283), .Z(n24286) );
  XOR U24924 ( .A(n24285), .B(n24286), .Z(n24255) );
  XOR U24925 ( .A(n24256), .B(n24255), .Z(n24258) );
  NAND U24926 ( .A(n187), .B(n24175), .Z(n24177) );
  XOR U24927 ( .A(b[13]), .B(a[165]), .Z(n24304) );
  NAND U24928 ( .A(n37295), .B(n24304), .Z(n24176) );
  AND U24929 ( .A(n24177), .B(n24176), .Z(n24250) );
  NAND U24930 ( .A(n186), .B(n24178), .Z(n24180) );
  XOR U24931 ( .A(b[11]), .B(a[167]), .Z(n24307) );
  NAND U24932 ( .A(n37097), .B(n24307), .Z(n24179) );
  NAND U24933 ( .A(n24180), .B(n24179), .Z(n24249) );
  XNOR U24934 ( .A(n24250), .B(n24249), .Z(n24252) );
  NAND U24935 ( .A(n188), .B(n24181), .Z(n24183) );
  XOR U24936 ( .A(b[15]), .B(a[163]), .Z(n24310) );
  NAND U24937 ( .A(n37382), .B(n24310), .Z(n24182) );
  AND U24938 ( .A(n24183), .B(n24182), .Z(n24246) );
  NAND U24939 ( .A(n38064), .B(n24184), .Z(n24186) );
  XOR U24940 ( .A(b[21]), .B(a[157]), .Z(n24313) );
  NAND U24941 ( .A(n37993), .B(n24313), .Z(n24185) );
  AND U24942 ( .A(n24186), .B(n24185), .Z(n24244) );
  NAND U24943 ( .A(n185), .B(n24187), .Z(n24189) );
  XOR U24944 ( .A(b[9]), .B(a[169]), .Z(n24316) );
  NAND U24945 ( .A(n36805), .B(n24316), .Z(n24188) );
  NAND U24946 ( .A(n24189), .B(n24188), .Z(n24243) );
  XNOR U24947 ( .A(n24244), .B(n24243), .Z(n24245) );
  XNOR U24948 ( .A(n24246), .B(n24245), .Z(n24251) );
  XOR U24949 ( .A(n24252), .B(n24251), .Z(n24257) );
  XNOR U24950 ( .A(n24258), .B(n24257), .Z(n24269) );
  XNOR U24951 ( .A(n24270), .B(n24269), .Z(n24325) );
  XNOR U24952 ( .A(n24326), .B(n24325), .Z(n24327) );
  XOR U24953 ( .A(n24328), .B(n24327), .Z(n24332) );
  XNOR U24954 ( .A(n24331), .B(n24332), .Z(n24333) );
  XNOR U24955 ( .A(n24334), .B(n24333), .Z(n24339) );
  XOR U24956 ( .A(n24340), .B(n24339), .Z(n24208) );
  NANDN U24957 ( .A(n24191), .B(n24190), .Z(n24195) );
  OR U24958 ( .A(n24193), .B(n24192), .Z(n24194) );
  AND U24959 ( .A(n24195), .B(n24194), .Z(n24207) );
  XNOR U24960 ( .A(n24208), .B(n24207), .Z(n24209) );
  XNOR U24961 ( .A(n24210), .B(n24209), .Z(n24201) );
  XNOR U24962 ( .A(n24202), .B(n24201), .Z(n24203) );
  XNOR U24963 ( .A(n24204), .B(n24203), .Z(n24343) );
  XNOR U24964 ( .A(sreg[401]), .B(n24343), .Z(n24345) );
  NANDN U24965 ( .A(sreg[400]), .B(n24196), .Z(n24200) );
  NAND U24966 ( .A(n24198), .B(n24197), .Z(n24199) );
  NAND U24967 ( .A(n24200), .B(n24199), .Z(n24344) );
  XNOR U24968 ( .A(n24345), .B(n24344), .Z(c[401]) );
  NANDN U24969 ( .A(n24202), .B(n24201), .Z(n24206) );
  NANDN U24970 ( .A(n24204), .B(n24203), .Z(n24205) );
  AND U24971 ( .A(n24206), .B(n24205), .Z(n24351) );
  NANDN U24972 ( .A(n24208), .B(n24207), .Z(n24212) );
  NANDN U24973 ( .A(n24210), .B(n24209), .Z(n24211) );
  AND U24974 ( .A(n24212), .B(n24211), .Z(n24349) );
  NANDN U24975 ( .A(n24214), .B(n24213), .Z(n24218) );
  NANDN U24976 ( .A(n24216), .B(n24215), .Z(n24217) );
  AND U24977 ( .A(n24218), .B(n24217), .Z(n24426) );
  NAND U24978 ( .A(n38385), .B(n24219), .Z(n24221) );
  XOR U24979 ( .A(b[27]), .B(a[152]), .Z(n24372) );
  NAND U24980 ( .A(n38343), .B(n24372), .Z(n24220) );
  AND U24981 ( .A(n24221), .B(n24220), .Z(n24433) );
  NAND U24982 ( .A(n183), .B(n24222), .Z(n24224) );
  XOR U24983 ( .A(b[5]), .B(a[174]), .Z(n24375) );
  NAND U24984 ( .A(n36296), .B(n24375), .Z(n24223) );
  AND U24985 ( .A(n24224), .B(n24223), .Z(n24431) );
  NAND U24986 ( .A(n190), .B(n24225), .Z(n24227) );
  XOR U24987 ( .A(b[19]), .B(a[160]), .Z(n24378) );
  NAND U24988 ( .A(n37821), .B(n24378), .Z(n24226) );
  NAND U24989 ( .A(n24227), .B(n24226), .Z(n24430) );
  XNOR U24990 ( .A(n24431), .B(n24430), .Z(n24432) );
  XNOR U24991 ( .A(n24433), .B(n24432), .Z(n24424) );
  NAND U24992 ( .A(n38470), .B(n24228), .Z(n24230) );
  XOR U24993 ( .A(b[31]), .B(a[148]), .Z(n24381) );
  NAND U24994 ( .A(n38453), .B(n24381), .Z(n24229) );
  AND U24995 ( .A(n24230), .B(n24229), .Z(n24393) );
  NAND U24996 ( .A(n181), .B(n24231), .Z(n24233) );
  XOR U24997 ( .A(b[3]), .B(a[176]), .Z(n24384) );
  NAND U24998 ( .A(n182), .B(n24384), .Z(n24232) );
  AND U24999 ( .A(n24233), .B(n24232), .Z(n24391) );
  NAND U25000 ( .A(n189), .B(n24234), .Z(n24236) );
  XOR U25001 ( .A(b[17]), .B(a[162]), .Z(n24387) );
  NAND U25002 ( .A(n37652), .B(n24387), .Z(n24235) );
  NAND U25003 ( .A(n24236), .B(n24235), .Z(n24390) );
  XNOR U25004 ( .A(n24391), .B(n24390), .Z(n24392) );
  XOR U25005 ( .A(n24393), .B(n24392), .Z(n24425) );
  XOR U25006 ( .A(n24424), .B(n24425), .Z(n24427) );
  XOR U25007 ( .A(n24426), .B(n24427), .Z(n24473) );
  NANDN U25008 ( .A(n24238), .B(n24237), .Z(n24242) );
  NANDN U25009 ( .A(n24240), .B(n24239), .Z(n24241) );
  AND U25010 ( .A(n24242), .B(n24241), .Z(n24414) );
  NANDN U25011 ( .A(n24244), .B(n24243), .Z(n24248) );
  NANDN U25012 ( .A(n24246), .B(n24245), .Z(n24247) );
  NAND U25013 ( .A(n24248), .B(n24247), .Z(n24415) );
  XNOR U25014 ( .A(n24414), .B(n24415), .Z(n24416) );
  NANDN U25015 ( .A(n24250), .B(n24249), .Z(n24254) );
  NAND U25016 ( .A(n24252), .B(n24251), .Z(n24253) );
  NAND U25017 ( .A(n24254), .B(n24253), .Z(n24417) );
  XNOR U25018 ( .A(n24416), .B(n24417), .Z(n24472) );
  XNOR U25019 ( .A(n24473), .B(n24472), .Z(n24475) );
  NAND U25020 ( .A(n24256), .B(n24255), .Z(n24260) );
  NAND U25021 ( .A(n24258), .B(n24257), .Z(n24259) );
  AND U25022 ( .A(n24260), .B(n24259), .Z(n24474) );
  XOR U25023 ( .A(n24475), .B(n24474), .Z(n24486) );
  NANDN U25024 ( .A(n24262), .B(n24261), .Z(n24266) );
  NANDN U25025 ( .A(n24264), .B(n24263), .Z(n24265) );
  AND U25026 ( .A(n24266), .B(n24265), .Z(n24484) );
  NANDN U25027 ( .A(n24272), .B(n24271), .Z(n24276) );
  OR U25028 ( .A(n24274), .B(n24273), .Z(n24275) );
  AND U25029 ( .A(n24276), .B(n24275), .Z(n24479) );
  NANDN U25030 ( .A(n24278), .B(n24277), .Z(n24282) );
  NANDN U25031 ( .A(n24280), .B(n24279), .Z(n24281) );
  AND U25032 ( .A(n24282), .B(n24281), .Z(n24421) );
  NANDN U25033 ( .A(n24284), .B(n24283), .Z(n24288) );
  OR U25034 ( .A(n24286), .B(n24285), .Z(n24287) );
  NAND U25035 ( .A(n24288), .B(n24287), .Z(n24420) );
  XNOR U25036 ( .A(n24421), .B(n24420), .Z(n24423) );
  NAND U25037 ( .A(n194), .B(n24289), .Z(n24291) );
  XOR U25038 ( .A(b[29]), .B(a[150]), .Z(n24445) );
  NAND U25039 ( .A(n38456), .B(n24445), .Z(n24290) );
  AND U25040 ( .A(n24291), .B(n24290), .Z(n24367) );
  AND U25041 ( .A(b[31]), .B(a[146]), .Z(n24366) );
  XNOR U25042 ( .A(n24367), .B(n24366), .Z(n24368) );
  NAND U25043 ( .A(b[0]), .B(a[178]), .Z(n24292) );
  XNOR U25044 ( .A(b[1]), .B(n24292), .Z(n24294) );
  NANDN U25045 ( .A(b[0]), .B(a[177]), .Z(n24293) );
  NAND U25046 ( .A(n24294), .B(n24293), .Z(n24369) );
  XNOR U25047 ( .A(n24368), .B(n24369), .Z(n24409) );
  NAND U25048 ( .A(n38185), .B(n24295), .Z(n24297) );
  XOR U25049 ( .A(b[23]), .B(a[156]), .Z(n24448) );
  NAND U25050 ( .A(n38132), .B(n24448), .Z(n24296) );
  AND U25051 ( .A(n24297), .B(n24296), .Z(n24438) );
  NAND U25052 ( .A(n184), .B(n24298), .Z(n24300) );
  XOR U25053 ( .A(b[7]), .B(a[172]), .Z(n24451) );
  NAND U25054 ( .A(n36592), .B(n24451), .Z(n24299) );
  AND U25055 ( .A(n24300), .B(n24299), .Z(n24437) );
  NAND U25056 ( .A(n38289), .B(n24301), .Z(n24303) );
  XOR U25057 ( .A(b[25]), .B(a[154]), .Z(n24454) );
  NAND U25058 ( .A(n38247), .B(n24454), .Z(n24302) );
  NAND U25059 ( .A(n24303), .B(n24302), .Z(n24436) );
  XOR U25060 ( .A(n24437), .B(n24436), .Z(n24439) );
  XOR U25061 ( .A(n24438), .B(n24439), .Z(n24408) );
  XOR U25062 ( .A(n24409), .B(n24408), .Z(n24411) );
  NAND U25063 ( .A(n187), .B(n24304), .Z(n24306) );
  XOR U25064 ( .A(b[13]), .B(a[166]), .Z(n24457) );
  NAND U25065 ( .A(n37295), .B(n24457), .Z(n24305) );
  AND U25066 ( .A(n24306), .B(n24305), .Z(n24403) );
  NAND U25067 ( .A(n186), .B(n24307), .Z(n24309) );
  XOR U25068 ( .A(b[11]), .B(a[168]), .Z(n24460) );
  NAND U25069 ( .A(n37097), .B(n24460), .Z(n24308) );
  NAND U25070 ( .A(n24309), .B(n24308), .Z(n24402) );
  XNOR U25071 ( .A(n24403), .B(n24402), .Z(n24405) );
  NAND U25072 ( .A(n188), .B(n24310), .Z(n24312) );
  XOR U25073 ( .A(b[15]), .B(a[164]), .Z(n24463) );
  NAND U25074 ( .A(n37382), .B(n24463), .Z(n24311) );
  AND U25075 ( .A(n24312), .B(n24311), .Z(n24399) );
  NAND U25076 ( .A(n38064), .B(n24313), .Z(n24315) );
  XOR U25077 ( .A(b[21]), .B(a[158]), .Z(n24466) );
  NAND U25078 ( .A(n37993), .B(n24466), .Z(n24314) );
  AND U25079 ( .A(n24315), .B(n24314), .Z(n24397) );
  NAND U25080 ( .A(n185), .B(n24316), .Z(n24318) );
  XOR U25081 ( .A(b[9]), .B(a[170]), .Z(n24469) );
  NAND U25082 ( .A(n36805), .B(n24469), .Z(n24317) );
  NAND U25083 ( .A(n24318), .B(n24317), .Z(n24396) );
  XNOR U25084 ( .A(n24397), .B(n24396), .Z(n24398) );
  XNOR U25085 ( .A(n24399), .B(n24398), .Z(n24404) );
  XOR U25086 ( .A(n24405), .B(n24404), .Z(n24410) );
  XNOR U25087 ( .A(n24411), .B(n24410), .Z(n24422) );
  XNOR U25088 ( .A(n24423), .B(n24422), .Z(n24478) );
  XNOR U25089 ( .A(n24479), .B(n24478), .Z(n24480) );
  XOR U25090 ( .A(n24481), .B(n24480), .Z(n24485) );
  XOR U25091 ( .A(n24484), .B(n24485), .Z(n24487) );
  XOR U25092 ( .A(n24486), .B(n24487), .Z(n24363) );
  NANDN U25093 ( .A(n24320), .B(n24319), .Z(n24324) );
  NAND U25094 ( .A(n24322), .B(n24321), .Z(n24323) );
  AND U25095 ( .A(n24324), .B(n24323), .Z(n24361) );
  NANDN U25096 ( .A(n24326), .B(n24325), .Z(n24330) );
  NANDN U25097 ( .A(n24328), .B(n24327), .Z(n24329) );
  AND U25098 ( .A(n24330), .B(n24329), .Z(n24360) );
  XNOR U25099 ( .A(n24361), .B(n24360), .Z(n24362) );
  XNOR U25100 ( .A(n24363), .B(n24362), .Z(n24354) );
  NANDN U25101 ( .A(n24332), .B(n24331), .Z(n24336) );
  NANDN U25102 ( .A(n24334), .B(n24333), .Z(n24335) );
  NAND U25103 ( .A(n24336), .B(n24335), .Z(n24355) );
  XNOR U25104 ( .A(n24354), .B(n24355), .Z(n24356) );
  NANDN U25105 ( .A(n24338), .B(n24337), .Z(n24342) );
  NAND U25106 ( .A(n24340), .B(n24339), .Z(n24341) );
  NAND U25107 ( .A(n24342), .B(n24341), .Z(n24357) );
  XNOR U25108 ( .A(n24356), .B(n24357), .Z(n24348) );
  XNOR U25109 ( .A(n24349), .B(n24348), .Z(n24350) );
  XNOR U25110 ( .A(n24351), .B(n24350), .Z(n24490) );
  XNOR U25111 ( .A(sreg[402]), .B(n24490), .Z(n24492) );
  NANDN U25112 ( .A(sreg[401]), .B(n24343), .Z(n24347) );
  NAND U25113 ( .A(n24345), .B(n24344), .Z(n24346) );
  NAND U25114 ( .A(n24347), .B(n24346), .Z(n24491) );
  XNOR U25115 ( .A(n24492), .B(n24491), .Z(c[402]) );
  NANDN U25116 ( .A(n24349), .B(n24348), .Z(n24353) );
  NANDN U25117 ( .A(n24351), .B(n24350), .Z(n24352) );
  AND U25118 ( .A(n24353), .B(n24352), .Z(n24498) );
  NANDN U25119 ( .A(n24355), .B(n24354), .Z(n24359) );
  NANDN U25120 ( .A(n24357), .B(n24356), .Z(n24358) );
  AND U25121 ( .A(n24359), .B(n24358), .Z(n24496) );
  NANDN U25122 ( .A(n24361), .B(n24360), .Z(n24365) );
  NANDN U25123 ( .A(n24363), .B(n24362), .Z(n24364) );
  AND U25124 ( .A(n24365), .B(n24364), .Z(n24504) );
  NANDN U25125 ( .A(n24367), .B(n24366), .Z(n24371) );
  NANDN U25126 ( .A(n24369), .B(n24368), .Z(n24370) );
  AND U25127 ( .A(n24371), .B(n24370), .Z(n24575) );
  NAND U25128 ( .A(n38385), .B(n24372), .Z(n24374) );
  XOR U25129 ( .A(b[27]), .B(a[153]), .Z(n24519) );
  NAND U25130 ( .A(n38343), .B(n24519), .Z(n24373) );
  AND U25131 ( .A(n24374), .B(n24373), .Z(n24582) );
  NAND U25132 ( .A(n183), .B(n24375), .Z(n24377) );
  XOR U25133 ( .A(b[5]), .B(a[175]), .Z(n24522) );
  NAND U25134 ( .A(n36296), .B(n24522), .Z(n24376) );
  AND U25135 ( .A(n24377), .B(n24376), .Z(n24580) );
  NAND U25136 ( .A(n190), .B(n24378), .Z(n24380) );
  XOR U25137 ( .A(b[19]), .B(a[161]), .Z(n24525) );
  NAND U25138 ( .A(n37821), .B(n24525), .Z(n24379) );
  NAND U25139 ( .A(n24380), .B(n24379), .Z(n24579) );
  XNOR U25140 ( .A(n24580), .B(n24579), .Z(n24581) );
  XNOR U25141 ( .A(n24582), .B(n24581), .Z(n24573) );
  NAND U25142 ( .A(n38470), .B(n24381), .Z(n24383) );
  XOR U25143 ( .A(b[31]), .B(a[149]), .Z(n24528) );
  NAND U25144 ( .A(n38453), .B(n24528), .Z(n24382) );
  AND U25145 ( .A(n24383), .B(n24382), .Z(n24540) );
  NAND U25146 ( .A(n181), .B(n24384), .Z(n24386) );
  XOR U25147 ( .A(b[3]), .B(a[177]), .Z(n24531) );
  NAND U25148 ( .A(n182), .B(n24531), .Z(n24385) );
  AND U25149 ( .A(n24386), .B(n24385), .Z(n24538) );
  NAND U25150 ( .A(n189), .B(n24387), .Z(n24389) );
  XOR U25151 ( .A(b[17]), .B(a[163]), .Z(n24534) );
  NAND U25152 ( .A(n37652), .B(n24534), .Z(n24388) );
  NAND U25153 ( .A(n24389), .B(n24388), .Z(n24537) );
  XNOR U25154 ( .A(n24538), .B(n24537), .Z(n24539) );
  XOR U25155 ( .A(n24540), .B(n24539), .Z(n24574) );
  XOR U25156 ( .A(n24573), .B(n24574), .Z(n24576) );
  XOR U25157 ( .A(n24575), .B(n24576), .Z(n24622) );
  NANDN U25158 ( .A(n24391), .B(n24390), .Z(n24395) );
  NANDN U25159 ( .A(n24393), .B(n24392), .Z(n24394) );
  AND U25160 ( .A(n24395), .B(n24394), .Z(n24561) );
  NANDN U25161 ( .A(n24397), .B(n24396), .Z(n24401) );
  NANDN U25162 ( .A(n24399), .B(n24398), .Z(n24400) );
  NAND U25163 ( .A(n24401), .B(n24400), .Z(n24562) );
  XNOR U25164 ( .A(n24561), .B(n24562), .Z(n24563) );
  NANDN U25165 ( .A(n24403), .B(n24402), .Z(n24407) );
  NAND U25166 ( .A(n24405), .B(n24404), .Z(n24406) );
  NAND U25167 ( .A(n24407), .B(n24406), .Z(n24564) );
  XNOR U25168 ( .A(n24563), .B(n24564), .Z(n24621) );
  XNOR U25169 ( .A(n24622), .B(n24621), .Z(n24624) );
  NAND U25170 ( .A(n24409), .B(n24408), .Z(n24413) );
  NAND U25171 ( .A(n24411), .B(n24410), .Z(n24412) );
  AND U25172 ( .A(n24413), .B(n24412), .Z(n24623) );
  XOR U25173 ( .A(n24624), .B(n24623), .Z(n24635) );
  NANDN U25174 ( .A(n24415), .B(n24414), .Z(n24419) );
  NANDN U25175 ( .A(n24417), .B(n24416), .Z(n24418) );
  AND U25176 ( .A(n24419), .B(n24418), .Z(n24633) );
  NANDN U25177 ( .A(n24425), .B(n24424), .Z(n24429) );
  OR U25178 ( .A(n24427), .B(n24426), .Z(n24428) );
  AND U25179 ( .A(n24429), .B(n24428), .Z(n24628) );
  NANDN U25180 ( .A(n24431), .B(n24430), .Z(n24435) );
  NANDN U25181 ( .A(n24433), .B(n24432), .Z(n24434) );
  AND U25182 ( .A(n24435), .B(n24434), .Z(n24568) );
  NANDN U25183 ( .A(n24437), .B(n24436), .Z(n24441) );
  OR U25184 ( .A(n24439), .B(n24438), .Z(n24440) );
  NAND U25185 ( .A(n24441), .B(n24440), .Z(n24567) );
  XNOR U25186 ( .A(n24568), .B(n24567), .Z(n24569) );
  NAND U25187 ( .A(b[0]), .B(a[179]), .Z(n24442) );
  XNOR U25188 ( .A(b[1]), .B(n24442), .Z(n24444) );
  NANDN U25189 ( .A(b[0]), .B(a[178]), .Z(n24443) );
  NAND U25190 ( .A(n24444), .B(n24443), .Z(n24516) );
  NAND U25191 ( .A(n194), .B(n24445), .Z(n24447) );
  XOR U25192 ( .A(b[29]), .B(a[151]), .Z(n24594) );
  NAND U25193 ( .A(n38456), .B(n24594), .Z(n24446) );
  AND U25194 ( .A(n24447), .B(n24446), .Z(n24514) );
  AND U25195 ( .A(b[31]), .B(a[147]), .Z(n24513) );
  XNOR U25196 ( .A(n24514), .B(n24513), .Z(n24515) );
  XNOR U25197 ( .A(n24516), .B(n24515), .Z(n24555) );
  NAND U25198 ( .A(n38185), .B(n24448), .Z(n24450) );
  XOR U25199 ( .A(b[23]), .B(a[157]), .Z(n24597) );
  NAND U25200 ( .A(n38132), .B(n24597), .Z(n24449) );
  AND U25201 ( .A(n24450), .B(n24449), .Z(n24588) );
  NAND U25202 ( .A(n184), .B(n24451), .Z(n24453) );
  XOR U25203 ( .A(b[7]), .B(a[173]), .Z(n24600) );
  NAND U25204 ( .A(n36592), .B(n24600), .Z(n24452) );
  AND U25205 ( .A(n24453), .B(n24452), .Z(n24586) );
  NAND U25206 ( .A(n38289), .B(n24454), .Z(n24456) );
  XOR U25207 ( .A(b[25]), .B(a[155]), .Z(n24603) );
  NAND U25208 ( .A(n38247), .B(n24603), .Z(n24455) );
  NAND U25209 ( .A(n24456), .B(n24455), .Z(n24585) );
  XNOR U25210 ( .A(n24586), .B(n24585), .Z(n24587) );
  XOR U25211 ( .A(n24588), .B(n24587), .Z(n24556) );
  XNOR U25212 ( .A(n24555), .B(n24556), .Z(n24557) );
  NAND U25213 ( .A(n187), .B(n24457), .Z(n24459) );
  XOR U25214 ( .A(b[13]), .B(a[167]), .Z(n24606) );
  NAND U25215 ( .A(n37295), .B(n24606), .Z(n24458) );
  AND U25216 ( .A(n24459), .B(n24458), .Z(n24550) );
  NAND U25217 ( .A(n186), .B(n24460), .Z(n24462) );
  XOR U25218 ( .A(b[11]), .B(a[169]), .Z(n24609) );
  NAND U25219 ( .A(n37097), .B(n24609), .Z(n24461) );
  NAND U25220 ( .A(n24462), .B(n24461), .Z(n24549) );
  XNOR U25221 ( .A(n24550), .B(n24549), .Z(n24551) );
  NAND U25222 ( .A(n188), .B(n24463), .Z(n24465) );
  XOR U25223 ( .A(b[15]), .B(a[165]), .Z(n24612) );
  NAND U25224 ( .A(n37382), .B(n24612), .Z(n24464) );
  AND U25225 ( .A(n24465), .B(n24464), .Z(n24546) );
  NAND U25226 ( .A(n38064), .B(n24466), .Z(n24468) );
  XOR U25227 ( .A(b[21]), .B(a[159]), .Z(n24615) );
  NAND U25228 ( .A(n37993), .B(n24615), .Z(n24467) );
  AND U25229 ( .A(n24468), .B(n24467), .Z(n24544) );
  NAND U25230 ( .A(n185), .B(n24469), .Z(n24471) );
  XOR U25231 ( .A(b[9]), .B(a[171]), .Z(n24618) );
  NAND U25232 ( .A(n36805), .B(n24618), .Z(n24470) );
  NAND U25233 ( .A(n24471), .B(n24470), .Z(n24543) );
  XNOR U25234 ( .A(n24544), .B(n24543), .Z(n24545) );
  XOR U25235 ( .A(n24546), .B(n24545), .Z(n24552) );
  XOR U25236 ( .A(n24551), .B(n24552), .Z(n24558) );
  XOR U25237 ( .A(n24557), .B(n24558), .Z(n24570) );
  XNOR U25238 ( .A(n24569), .B(n24570), .Z(n24627) );
  XNOR U25239 ( .A(n24628), .B(n24627), .Z(n24629) );
  XOR U25240 ( .A(n24630), .B(n24629), .Z(n24634) );
  XOR U25241 ( .A(n24633), .B(n24634), .Z(n24636) );
  XOR U25242 ( .A(n24635), .B(n24636), .Z(n24510) );
  NANDN U25243 ( .A(n24473), .B(n24472), .Z(n24477) );
  NAND U25244 ( .A(n24475), .B(n24474), .Z(n24476) );
  AND U25245 ( .A(n24477), .B(n24476), .Z(n24508) );
  NANDN U25246 ( .A(n24479), .B(n24478), .Z(n24483) );
  NANDN U25247 ( .A(n24481), .B(n24480), .Z(n24482) );
  AND U25248 ( .A(n24483), .B(n24482), .Z(n24507) );
  XNOR U25249 ( .A(n24508), .B(n24507), .Z(n24509) );
  XNOR U25250 ( .A(n24510), .B(n24509), .Z(n24501) );
  NANDN U25251 ( .A(n24485), .B(n24484), .Z(n24489) );
  OR U25252 ( .A(n24487), .B(n24486), .Z(n24488) );
  NAND U25253 ( .A(n24489), .B(n24488), .Z(n24502) );
  XNOR U25254 ( .A(n24501), .B(n24502), .Z(n24503) );
  XNOR U25255 ( .A(n24504), .B(n24503), .Z(n24495) );
  XNOR U25256 ( .A(n24496), .B(n24495), .Z(n24497) );
  XNOR U25257 ( .A(n24498), .B(n24497), .Z(n24639) );
  XNOR U25258 ( .A(sreg[403]), .B(n24639), .Z(n24641) );
  NANDN U25259 ( .A(sreg[402]), .B(n24490), .Z(n24494) );
  NAND U25260 ( .A(n24492), .B(n24491), .Z(n24493) );
  NAND U25261 ( .A(n24494), .B(n24493), .Z(n24640) );
  XNOR U25262 ( .A(n24641), .B(n24640), .Z(c[403]) );
  NANDN U25263 ( .A(n24496), .B(n24495), .Z(n24500) );
  NANDN U25264 ( .A(n24498), .B(n24497), .Z(n24499) );
  AND U25265 ( .A(n24500), .B(n24499), .Z(n24647) );
  NANDN U25266 ( .A(n24502), .B(n24501), .Z(n24506) );
  NANDN U25267 ( .A(n24504), .B(n24503), .Z(n24505) );
  AND U25268 ( .A(n24506), .B(n24505), .Z(n24645) );
  NANDN U25269 ( .A(n24508), .B(n24507), .Z(n24512) );
  NANDN U25270 ( .A(n24510), .B(n24509), .Z(n24511) );
  AND U25271 ( .A(n24512), .B(n24511), .Z(n24653) );
  NANDN U25272 ( .A(n24514), .B(n24513), .Z(n24518) );
  NANDN U25273 ( .A(n24516), .B(n24515), .Z(n24517) );
  AND U25274 ( .A(n24518), .B(n24517), .Z(n24736) );
  NAND U25275 ( .A(n38385), .B(n24519), .Z(n24521) );
  XOR U25276 ( .A(b[27]), .B(a[154]), .Z(n24680) );
  NAND U25277 ( .A(n38343), .B(n24680), .Z(n24520) );
  AND U25278 ( .A(n24521), .B(n24520), .Z(n24743) );
  NAND U25279 ( .A(n183), .B(n24522), .Z(n24524) );
  XOR U25280 ( .A(b[5]), .B(a[176]), .Z(n24683) );
  NAND U25281 ( .A(n36296), .B(n24683), .Z(n24523) );
  AND U25282 ( .A(n24524), .B(n24523), .Z(n24741) );
  NAND U25283 ( .A(n190), .B(n24525), .Z(n24527) );
  XOR U25284 ( .A(b[19]), .B(a[162]), .Z(n24686) );
  NAND U25285 ( .A(n37821), .B(n24686), .Z(n24526) );
  NAND U25286 ( .A(n24527), .B(n24526), .Z(n24740) );
  XNOR U25287 ( .A(n24741), .B(n24740), .Z(n24742) );
  XNOR U25288 ( .A(n24743), .B(n24742), .Z(n24734) );
  NAND U25289 ( .A(n38470), .B(n24528), .Z(n24530) );
  XOR U25290 ( .A(b[31]), .B(a[150]), .Z(n24689) );
  NAND U25291 ( .A(n38453), .B(n24689), .Z(n24529) );
  AND U25292 ( .A(n24530), .B(n24529), .Z(n24701) );
  NAND U25293 ( .A(n181), .B(n24531), .Z(n24533) );
  XOR U25294 ( .A(b[3]), .B(a[178]), .Z(n24692) );
  NAND U25295 ( .A(n182), .B(n24692), .Z(n24532) );
  AND U25296 ( .A(n24533), .B(n24532), .Z(n24699) );
  NAND U25297 ( .A(n189), .B(n24534), .Z(n24536) );
  XOR U25298 ( .A(b[17]), .B(a[164]), .Z(n24695) );
  NAND U25299 ( .A(n37652), .B(n24695), .Z(n24535) );
  NAND U25300 ( .A(n24536), .B(n24535), .Z(n24698) );
  XNOR U25301 ( .A(n24699), .B(n24698), .Z(n24700) );
  XOR U25302 ( .A(n24701), .B(n24700), .Z(n24735) );
  XOR U25303 ( .A(n24734), .B(n24735), .Z(n24737) );
  XOR U25304 ( .A(n24736), .B(n24737), .Z(n24669) );
  NANDN U25305 ( .A(n24538), .B(n24537), .Z(n24542) );
  NANDN U25306 ( .A(n24540), .B(n24539), .Z(n24541) );
  AND U25307 ( .A(n24542), .B(n24541), .Z(n24722) );
  NANDN U25308 ( .A(n24544), .B(n24543), .Z(n24548) );
  NANDN U25309 ( .A(n24546), .B(n24545), .Z(n24547) );
  NAND U25310 ( .A(n24548), .B(n24547), .Z(n24723) );
  XNOR U25311 ( .A(n24722), .B(n24723), .Z(n24724) );
  NANDN U25312 ( .A(n24550), .B(n24549), .Z(n24554) );
  NANDN U25313 ( .A(n24552), .B(n24551), .Z(n24553) );
  NAND U25314 ( .A(n24554), .B(n24553), .Z(n24725) );
  XNOR U25315 ( .A(n24724), .B(n24725), .Z(n24668) );
  XNOR U25316 ( .A(n24669), .B(n24668), .Z(n24671) );
  NANDN U25317 ( .A(n24556), .B(n24555), .Z(n24560) );
  NANDN U25318 ( .A(n24558), .B(n24557), .Z(n24559) );
  AND U25319 ( .A(n24560), .B(n24559), .Z(n24670) );
  XOR U25320 ( .A(n24671), .B(n24670), .Z(n24784) );
  NANDN U25321 ( .A(n24562), .B(n24561), .Z(n24566) );
  NANDN U25322 ( .A(n24564), .B(n24563), .Z(n24565) );
  AND U25323 ( .A(n24566), .B(n24565), .Z(n24782) );
  NANDN U25324 ( .A(n24568), .B(n24567), .Z(n24572) );
  NANDN U25325 ( .A(n24570), .B(n24569), .Z(n24571) );
  AND U25326 ( .A(n24572), .B(n24571), .Z(n24665) );
  NANDN U25327 ( .A(n24574), .B(n24573), .Z(n24578) );
  OR U25328 ( .A(n24576), .B(n24575), .Z(n24577) );
  AND U25329 ( .A(n24578), .B(n24577), .Z(n24663) );
  NANDN U25330 ( .A(n24580), .B(n24579), .Z(n24584) );
  NANDN U25331 ( .A(n24582), .B(n24581), .Z(n24583) );
  AND U25332 ( .A(n24584), .B(n24583), .Z(n24729) );
  NANDN U25333 ( .A(n24586), .B(n24585), .Z(n24590) );
  NANDN U25334 ( .A(n24588), .B(n24587), .Z(n24589) );
  NAND U25335 ( .A(n24590), .B(n24589), .Z(n24728) );
  XNOR U25336 ( .A(n24729), .B(n24728), .Z(n24730) );
  NAND U25337 ( .A(b[0]), .B(a[180]), .Z(n24591) );
  XNOR U25338 ( .A(b[1]), .B(n24591), .Z(n24593) );
  NANDN U25339 ( .A(b[0]), .B(a[179]), .Z(n24592) );
  NAND U25340 ( .A(n24593), .B(n24592), .Z(n24677) );
  NAND U25341 ( .A(n194), .B(n24594), .Z(n24596) );
  XOR U25342 ( .A(b[29]), .B(a[152]), .Z(n24755) );
  NAND U25343 ( .A(n38456), .B(n24755), .Z(n24595) );
  AND U25344 ( .A(n24596), .B(n24595), .Z(n24675) );
  AND U25345 ( .A(b[31]), .B(a[148]), .Z(n24674) );
  XNOR U25346 ( .A(n24675), .B(n24674), .Z(n24676) );
  XNOR U25347 ( .A(n24677), .B(n24676), .Z(n24716) );
  NAND U25348 ( .A(n38185), .B(n24597), .Z(n24599) );
  XOR U25349 ( .A(b[23]), .B(a[158]), .Z(n24758) );
  NAND U25350 ( .A(n38132), .B(n24758), .Z(n24598) );
  AND U25351 ( .A(n24599), .B(n24598), .Z(n24749) );
  NAND U25352 ( .A(n184), .B(n24600), .Z(n24602) );
  XOR U25353 ( .A(b[7]), .B(a[174]), .Z(n24761) );
  NAND U25354 ( .A(n36592), .B(n24761), .Z(n24601) );
  AND U25355 ( .A(n24602), .B(n24601), .Z(n24747) );
  NAND U25356 ( .A(n38289), .B(n24603), .Z(n24605) );
  XOR U25357 ( .A(b[25]), .B(a[156]), .Z(n24764) );
  NAND U25358 ( .A(n38247), .B(n24764), .Z(n24604) );
  NAND U25359 ( .A(n24605), .B(n24604), .Z(n24746) );
  XNOR U25360 ( .A(n24747), .B(n24746), .Z(n24748) );
  XOR U25361 ( .A(n24749), .B(n24748), .Z(n24717) );
  XNOR U25362 ( .A(n24716), .B(n24717), .Z(n24718) );
  NAND U25363 ( .A(n187), .B(n24606), .Z(n24608) );
  XOR U25364 ( .A(b[13]), .B(a[168]), .Z(n24767) );
  NAND U25365 ( .A(n37295), .B(n24767), .Z(n24607) );
  AND U25366 ( .A(n24608), .B(n24607), .Z(n24711) );
  NAND U25367 ( .A(n186), .B(n24609), .Z(n24611) );
  XOR U25368 ( .A(b[11]), .B(a[170]), .Z(n24770) );
  NAND U25369 ( .A(n37097), .B(n24770), .Z(n24610) );
  NAND U25370 ( .A(n24611), .B(n24610), .Z(n24710) );
  XNOR U25371 ( .A(n24711), .B(n24710), .Z(n24712) );
  NAND U25372 ( .A(n188), .B(n24612), .Z(n24614) );
  XOR U25373 ( .A(b[15]), .B(a[166]), .Z(n24773) );
  NAND U25374 ( .A(n37382), .B(n24773), .Z(n24613) );
  AND U25375 ( .A(n24614), .B(n24613), .Z(n24707) );
  NAND U25376 ( .A(n38064), .B(n24615), .Z(n24617) );
  XOR U25377 ( .A(b[21]), .B(a[160]), .Z(n24776) );
  NAND U25378 ( .A(n37993), .B(n24776), .Z(n24616) );
  AND U25379 ( .A(n24617), .B(n24616), .Z(n24705) );
  NAND U25380 ( .A(n185), .B(n24618), .Z(n24620) );
  XOR U25381 ( .A(b[9]), .B(a[172]), .Z(n24779) );
  NAND U25382 ( .A(n36805), .B(n24779), .Z(n24619) );
  NAND U25383 ( .A(n24620), .B(n24619), .Z(n24704) );
  XNOR U25384 ( .A(n24705), .B(n24704), .Z(n24706) );
  XOR U25385 ( .A(n24707), .B(n24706), .Z(n24713) );
  XOR U25386 ( .A(n24712), .B(n24713), .Z(n24719) );
  XOR U25387 ( .A(n24718), .B(n24719), .Z(n24731) );
  XNOR U25388 ( .A(n24730), .B(n24731), .Z(n24662) );
  XNOR U25389 ( .A(n24663), .B(n24662), .Z(n24664) );
  XOR U25390 ( .A(n24665), .B(n24664), .Z(n24783) );
  XOR U25391 ( .A(n24782), .B(n24783), .Z(n24785) );
  XOR U25392 ( .A(n24784), .B(n24785), .Z(n24659) );
  NANDN U25393 ( .A(n24622), .B(n24621), .Z(n24626) );
  NAND U25394 ( .A(n24624), .B(n24623), .Z(n24625) );
  AND U25395 ( .A(n24626), .B(n24625), .Z(n24657) );
  NANDN U25396 ( .A(n24628), .B(n24627), .Z(n24632) );
  NANDN U25397 ( .A(n24630), .B(n24629), .Z(n24631) );
  AND U25398 ( .A(n24632), .B(n24631), .Z(n24656) );
  XNOR U25399 ( .A(n24657), .B(n24656), .Z(n24658) );
  XNOR U25400 ( .A(n24659), .B(n24658), .Z(n24650) );
  NANDN U25401 ( .A(n24634), .B(n24633), .Z(n24638) );
  OR U25402 ( .A(n24636), .B(n24635), .Z(n24637) );
  NAND U25403 ( .A(n24638), .B(n24637), .Z(n24651) );
  XNOR U25404 ( .A(n24650), .B(n24651), .Z(n24652) );
  XNOR U25405 ( .A(n24653), .B(n24652), .Z(n24644) );
  XNOR U25406 ( .A(n24645), .B(n24644), .Z(n24646) );
  XNOR U25407 ( .A(n24647), .B(n24646), .Z(n24788) );
  XNOR U25408 ( .A(sreg[404]), .B(n24788), .Z(n24790) );
  NANDN U25409 ( .A(sreg[403]), .B(n24639), .Z(n24643) );
  NAND U25410 ( .A(n24641), .B(n24640), .Z(n24642) );
  NAND U25411 ( .A(n24643), .B(n24642), .Z(n24789) );
  XNOR U25412 ( .A(n24790), .B(n24789), .Z(c[404]) );
  NANDN U25413 ( .A(n24645), .B(n24644), .Z(n24649) );
  NANDN U25414 ( .A(n24647), .B(n24646), .Z(n24648) );
  AND U25415 ( .A(n24649), .B(n24648), .Z(n24796) );
  NANDN U25416 ( .A(n24651), .B(n24650), .Z(n24655) );
  NANDN U25417 ( .A(n24653), .B(n24652), .Z(n24654) );
  AND U25418 ( .A(n24655), .B(n24654), .Z(n24794) );
  NANDN U25419 ( .A(n24657), .B(n24656), .Z(n24661) );
  NANDN U25420 ( .A(n24659), .B(n24658), .Z(n24660) );
  AND U25421 ( .A(n24661), .B(n24660), .Z(n24802) );
  NANDN U25422 ( .A(n24663), .B(n24662), .Z(n24667) );
  NANDN U25423 ( .A(n24665), .B(n24664), .Z(n24666) );
  AND U25424 ( .A(n24667), .B(n24666), .Z(n24806) );
  NANDN U25425 ( .A(n24669), .B(n24668), .Z(n24673) );
  NAND U25426 ( .A(n24671), .B(n24670), .Z(n24672) );
  AND U25427 ( .A(n24673), .B(n24672), .Z(n24805) );
  XNOR U25428 ( .A(n24806), .B(n24805), .Z(n24808) );
  NANDN U25429 ( .A(n24675), .B(n24674), .Z(n24679) );
  NANDN U25430 ( .A(n24677), .B(n24676), .Z(n24678) );
  AND U25431 ( .A(n24679), .B(n24678), .Z(n24883) );
  NAND U25432 ( .A(n38385), .B(n24680), .Z(n24682) );
  XOR U25433 ( .A(b[27]), .B(a[155]), .Z(n24829) );
  NAND U25434 ( .A(n38343), .B(n24829), .Z(n24681) );
  AND U25435 ( .A(n24682), .B(n24681), .Z(n24890) );
  NAND U25436 ( .A(n183), .B(n24683), .Z(n24685) );
  XOR U25437 ( .A(b[5]), .B(a[177]), .Z(n24832) );
  NAND U25438 ( .A(n36296), .B(n24832), .Z(n24684) );
  AND U25439 ( .A(n24685), .B(n24684), .Z(n24888) );
  NAND U25440 ( .A(n190), .B(n24686), .Z(n24688) );
  XOR U25441 ( .A(b[19]), .B(a[163]), .Z(n24835) );
  NAND U25442 ( .A(n37821), .B(n24835), .Z(n24687) );
  NAND U25443 ( .A(n24688), .B(n24687), .Z(n24887) );
  XNOR U25444 ( .A(n24888), .B(n24887), .Z(n24889) );
  XNOR U25445 ( .A(n24890), .B(n24889), .Z(n24881) );
  NAND U25446 ( .A(n38470), .B(n24689), .Z(n24691) );
  XOR U25447 ( .A(b[31]), .B(a[151]), .Z(n24838) );
  NAND U25448 ( .A(n38453), .B(n24838), .Z(n24690) );
  AND U25449 ( .A(n24691), .B(n24690), .Z(n24850) );
  NAND U25450 ( .A(n181), .B(n24692), .Z(n24694) );
  XOR U25451 ( .A(b[3]), .B(a[179]), .Z(n24841) );
  NAND U25452 ( .A(n182), .B(n24841), .Z(n24693) );
  AND U25453 ( .A(n24694), .B(n24693), .Z(n24848) );
  NAND U25454 ( .A(n189), .B(n24695), .Z(n24697) );
  XOR U25455 ( .A(b[17]), .B(a[165]), .Z(n24844) );
  NAND U25456 ( .A(n37652), .B(n24844), .Z(n24696) );
  NAND U25457 ( .A(n24697), .B(n24696), .Z(n24847) );
  XNOR U25458 ( .A(n24848), .B(n24847), .Z(n24849) );
  XOR U25459 ( .A(n24850), .B(n24849), .Z(n24882) );
  XOR U25460 ( .A(n24881), .B(n24882), .Z(n24884) );
  XOR U25461 ( .A(n24883), .B(n24884), .Z(n24818) );
  NANDN U25462 ( .A(n24699), .B(n24698), .Z(n24703) );
  NANDN U25463 ( .A(n24701), .B(n24700), .Z(n24702) );
  AND U25464 ( .A(n24703), .B(n24702), .Z(n24871) );
  NANDN U25465 ( .A(n24705), .B(n24704), .Z(n24709) );
  NANDN U25466 ( .A(n24707), .B(n24706), .Z(n24708) );
  NAND U25467 ( .A(n24709), .B(n24708), .Z(n24872) );
  XNOR U25468 ( .A(n24871), .B(n24872), .Z(n24873) );
  NANDN U25469 ( .A(n24711), .B(n24710), .Z(n24715) );
  NANDN U25470 ( .A(n24713), .B(n24712), .Z(n24714) );
  NAND U25471 ( .A(n24715), .B(n24714), .Z(n24874) );
  XNOR U25472 ( .A(n24873), .B(n24874), .Z(n24817) );
  XNOR U25473 ( .A(n24818), .B(n24817), .Z(n24820) );
  NANDN U25474 ( .A(n24717), .B(n24716), .Z(n24721) );
  NANDN U25475 ( .A(n24719), .B(n24718), .Z(n24720) );
  AND U25476 ( .A(n24721), .B(n24720), .Z(n24819) );
  XOR U25477 ( .A(n24820), .B(n24819), .Z(n24932) );
  NANDN U25478 ( .A(n24723), .B(n24722), .Z(n24727) );
  NANDN U25479 ( .A(n24725), .B(n24724), .Z(n24726) );
  AND U25480 ( .A(n24727), .B(n24726), .Z(n24929) );
  NANDN U25481 ( .A(n24729), .B(n24728), .Z(n24733) );
  NANDN U25482 ( .A(n24731), .B(n24730), .Z(n24732) );
  AND U25483 ( .A(n24733), .B(n24732), .Z(n24814) );
  NANDN U25484 ( .A(n24735), .B(n24734), .Z(n24739) );
  OR U25485 ( .A(n24737), .B(n24736), .Z(n24738) );
  AND U25486 ( .A(n24739), .B(n24738), .Z(n24812) );
  NANDN U25487 ( .A(n24741), .B(n24740), .Z(n24745) );
  NANDN U25488 ( .A(n24743), .B(n24742), .Z(n24744) );
  AND U25489 ( .A(n24745), .B(n24744), .Z(n24878) );
  NANDN U25490 ( .A(n24747), .B(n24746), .Z(n24751) );
  NANDN U25491 ( .A(n24749), .B(n24748), .Z(n24750) );
  NAND U25492 ( .A(n24751), .B(n24750), .Z(n24877) );
  XNOR U25493 ( .A(n24878), .B(n24877), .Z(n24880) );
  NAND U25494 ( .A(b[0]), .B(a[181]), .Z(n24752) );
  XNOR U25495 ( .A(b[1]), .B(n24752), .Z(n24754) );
  NANDN U25496 ( .A(b[0]), .B(a[180]), .Z(n24753) );
  NAND U25497 ( .A(n24754), .B(n24753), .Z(n24826) );
  NAND U25498 ( .A(n194), .B(n24755), .Z(n24757) );
  XOR U25499 ( .A(b[29]), .B(a[153]), .Z(n24902) );
  NAND U25500 ( .A(n38456), .B(n24902), .Z(n24756) );
  AND U25501 ( .A(n24757), .B(n24756), .Z(n24824) );
  AND U25502 ( .A(b[31]), .B(a[149]), .Z(n24823) );
  XNOR U25503 ( .A(n24824), .B(n24823), .Z(n24825) );
  XNOR U25504 ( .A(n24826), .B(n24825), .Z(n24866) );
  NAND U25505 ( .A(n38185), .B(n24758), .Z(n24760) );
  XOR U25506 ( .A(b[23]), .B(a[159]), .Z(n24905) );
  NAND U25507 ( .A(n38132), .B(n24905), .Z(n24759) );
  AND U25508 ( .A(n24760), .B(n24759), .Z(n24895) );
  NAND U25509 ( .A(n184), .B(n24761), .Z(n24763) );
  XOR U25510 ( .A(b[7]), .B(a[175]), .Z(n24908) );
  NAND U25511 ( .A(n36592), .B(n24908), .Z(n24762) );
  AND U25512 ( .A(n24763), .B(n24762), .Z(n24894) );
  NAND U25513 ( .A(n38289), .B(n24764), .Z(n24766) );
  XOR U25514 ( .A(b[25]), .B(a[157]), .Z(n24911) );
  NAND U25515 ( .A(n38247), .B(n24911), .Z(n24765) );
  NAND U25516 ( .A(n24766), .B(n24765), .Z(n24893) );
  XOR U25517 ( .A(n24894), .B(n24893), .Z(n24896) );
  XOR U25518 ( .A(n24895), .B(n24896), .Z(n24865) );
  XOR U25519 ( .A(n24866), .B(n24865), .Z(n24868) );
  NAND U25520 ( .A(n187), .B(n24767), .Z(n24769) );
  XOR U25521 ( .A(b[13]), .B(a[169]), .Z(n24914) );
  NAND U25522 ( .A(n37295), .B(n24914), .Z(n24768) );
  AND U25523 ( .A(n24769), .B(n24768), .Z(n24860) );
  NAND U25524 ( .A(n186), .B(n24770), .Z(n24772) );
  XOR U25525 ( .A(b[11]), .B(a[171]), .Z(n24917) );
  NAND U25526 ( .A(n37097), .B(n24917), .Z(n24771) );
  NAND U25527 ( .A(n24772), .B(n24771), .Z(n24859) );
  XNOR U25528 ( .A(n24860), .B(n24859), .Z(n24862) );
  NAND U25529 ( .A(n188), .B(n24773), .Z(n24775) );
  XOR U25530 ( .A(b[15]), .B(a[167]), .Z(n24920) );
  NAND U25531 ( .A(n37382), .B(n24920), .Z(n24774) );
  AND U25532 ( .A(n24775), .B(n24774), .Z(n24856) );
  NAND U25533 ( .A(n38064), .B(n24776), .Z(n24778) );
  XOR U25534 ( .A(b[21]), .B(a[161]), .Z(n24923) );
  NAND U25535 ( .A(n37993), .B(n24923), .Z(n24777) );
  AND U25536 ( .A(n24778), .B(n24777), .Z(n24854) );
  NAND U25537 ( .A(n185), .B(n24779), .Z(n24781) );
  XOR U25538 ( .A(b[9]), .B(a[173]), .Z(n24926) );
  NAND U25539 ( .A(n36805), .B(n24926), .Z(n24780) );
  NAND U25540 ( .A(n24781), .B(n24780), .Z(n24853) );
  XNOR U25541 ( .A(n24854), .B(n24853), .Z(n24855) );
  XNOR U25542 ( .A(n24856), .B(n24855), .Z(n24861) );
  XOR U25543 ( .A(n24862), .B(n24861), .Z(n24867) );
  XNOR U25544 ( .A(n24868), .B(n24867), .Z(n24879) );
  XNOR U25545 ( .A(n24880), .B(n24879), .Z(n24811) );
  XNOR U25546 ( .A(n24812), .B(n24811), .Z(n24813) );
  XOR U25547 ( .A(n24814), .B(n24813), .Z(n24930) );
  XNOR U25548 ( .A(n24929), .B(n24930), .Z(n24931) );
  XNOR U25549 ( .A(n24932), .B(n24931), .Z(n24807) );
  XOR U25550 ( .A(n24808), .B(n24807), .Z(n24800) );
  NANDN U25551 ( .A(n24783), .B(n24782), .Z(n24787) );
  OR U25552 ( .A(n24785), .B(n24784), .Z(n24786) );
  AND U25553 ( .A(n24787), .B(n24786), .Z(n24799) );
  XNOR U25554 ( .A(n24800), .B(n24799), .Z(n24801) );
  XNOR U25555 ( .A(n24802), .B(n24801), .Z(n24793) );
  XNOR U25556 ( .A(n24794), .B(n24793), .Z(n24795) );
  XNOR U25557 ( .A(n24796), .B(n24795), .Z(n24935) );
  XNOR U25558 ( .A(sreg[405]), .B(n24935), .Z(n24937) );
  NANDN U25559 ( .A(sreg[404]), .B(n24788), .Z(n24792) );
  NAND U25560 ( .A(n24790), .B(n24789), .Z(n24791) );
  NAND U25561 ( .A(n24792), .B(n24791), .Z(n24936) );
  XNOR U25562 ( .A(n24937), .B(n24936), .Z(c[405]) );
  NANDN U25563 ( .A(n24794), .B(n24793), .Z(n24798) );
  NANDN U25564 ( .A(n24796), .B(n24795), .Z(n24797) );
  AND U25565 ( .A(n24798), .B(n24797), .Z(n24943) );
  NANDN U25566 ( .A(n24800), .B(n24799), .Z(n24804) );
  NANDN U25567 ( .A(n24802), .B(n24801), .Z(n24803) );
  AND U25568 ( .A(n24804), .B(n24803), .Z(n24941) );
  NANDN U25569 ( .A(n24806), .B(n24805), .Z(n24810) );
  NAND U25570 ( .A(n24808), .B(n24807), .Z(n24809) );
  AND U25571 ( .A(n24810), .B(n24809), .Z(n24948) );
  NANDN U25572 ( .A(n24812), .B(n24811), .Z(n24816) );
  NANDN U25573 ( .A(n24814), .B(n24813), .Z(n24815) );
  AND U25574 ( .A(n24816), .B(n24815), .Z(n25079) );
  NANDN U25575 ( .A(n24818), .B(n24817), .Z(n24822) );
  NAND U25576 ( .A(n24820), .B(n24819), .Z(n24821) );
  AND U25577 ( .A(n24822), .B(n24821), .Z(n25078) );
  XNOR U25578 ( .A(n25079), .B(n25078), .Z(n25081) );
  NANDN U25579 ( .A(n24824), .B(n24823), .Z(n24828) );
  NANDN U25580 ( .A(n24826), .B(n24825), .Z(n24827) );
  AND U25581 ( .A(n24828), .B(n24827), .Z(n25014) );
  NAND U25582 ( .A(n38385), .B(n24829), .Z(n24831) );
  XOR U25583 ( .A(b[27]), .B(a[156]), .Z(n24958) );
  NAND U25584 ( .A(n38343), .B(n24958), .Z(n24830) );
  AND U25585 ( .A(n24831), .B(n24830), .Z(n25021) );
  NAND U25586 ( .A(n183), .B(n24832), .Z(n24834) );
  XOR U25587 ( .A(b[5]), .B(a[178]), .Z(n24961) );
  NAND U25588 ( .A(n36296), .B(n24961), .Z(n24833) );
  AND U25589 ( .A(n24834), .B(n24833), .Z(n25019) );
  NAND U25590 ( .A(n190), .B(n24835), .Z(n24837) );
  XOR U25591 ( .A(b[19]), .B(a[164]), .Z(n24964) );
  NAND U25592 ( .A(n37821), .B(n24964), .Z(n24836) );
  NAND U25593 ( .A(n24837), .B(n24836), .Z(n25018) );
  XNOR U25594 ( .A(n25019), .B(n25018), .Z(n25020) );
  XNOR U25595 ( .A(n25021), .B(n25020), .Z(n25012) );
  NAND U25596 ( .A(n38470), .B(n24838), .Z(n24840) );
  XOR U25597 ( .A(b[31]), .B(a[152]), .Z(n24967) );
  NAND U25598 ( .A(n38453), .B(n24967), .Z(n24839) );
  AND U25599 ( .A(n24840), .B(n24839), .Z(n24979) );
  NAND U25600 ( .A(n181), .B(n24841), .Z(n24843) );
  XOR U25601 ( .A(b[3]), .B(a[180]), .Z(n24970) );
  NAND U25602 ( .A(n182), .B(n24970), .Z(n24842) );
  AND U25603 ( .A(n24843), .B(n24842), .Z(n24977) );
  NAND U25604 ( .A(n189), .B(n24844), .Z(n24846) );
  XOR U25605 ( .A(b[17]), .B(a[166]), .Z(n24973) );
  NAND U25606 ( .A(n37652), .B(n24973), .Z(n24845) );
  NAND U25607 ( .A(n24846), .B(n24845), .Z(n24976) );
  XNOR U25608 ( .A(n24977), .B(n24976), .Z(n24978) );
  XOR U25609 ( .A(n24979), .B(n24978), .Z(n25013) );
  XOR U25610 ( .A(n25012), .B(n25013), .Z(n25015) );
  XOR U25611 ( .A(n25014), .B(n25015), .Z(n25061) );
  NANDN U25612 ( .A(n24848), .B(n24847), .Z(n24852) );
  NANDN U25613 ( .A(n24850), .B(n24849), .Z(n24851) );
  AND U25614 ( .A(n24852), .B(n24851), .Z(n25000) );
  NANDN U25615 ( .A(n24854), .B(n24853), .Z(n24858) );
  NANDN U25616 ( .A(n24856), .B(n24855), .Z(n24857) );
  NAND U25617 ( .A(n24858), .B(n24857), .Z(n25001) );
  XNOR U25618 ( .A(n25000), .B(n25001), .Z(n25002) );
  NANDN U25619 ( .A(n24860), .B(n24859), .Z(n24864) );
  NAND U25620 ( .A(n24862), .B(n24861), .Z(n24863) );
  NAND U25621 ( .A(n24864), .B(n24863), .Z(n25003) );
  XNOR U25622 ( .A(n25002), .B(n25003), .Z(n25060) );
  XNOR U25623 ( .A(n25061), .B(n25060), .Z(n25063) );
  NAND U25624 ( .A(n24866), .B(n24865), .Z(n24870) );
  NAND U25625 ( .A(n24868), .B(n24867), .Z(n24869) );
  AND U25626 ( .A(n24870), .B(n24869), .Z(n25062) );
  XOR U25627 ( .A(n25063), .B(n25062), .Z(n25075) );
  NANDN U25628 ( .A(n24872), .B(n24871), .Z(n24876) );
  NANDN U25629 ( .A(n24874), .B(n24873), .Z(n24875) );
  AND U25630 ( .A(n24876), .B(n24875), .Z(n25072) );
  NANDN U25631 ( .A(n24882), .B(n24881), .Z(n24886) );
  OR U25632 ( .A(n24884), .B(n24883), .Z(n24885) );
  AND U25633 ( .A(n24886), .B(n24885), .Z(n25067) );
  NANDN U25634 ( .A(n24888), .B(n24887), .Z(n24892) );
  NANDN U25635 ( .A(n24890), .B(n24889), .Z(n24891) );
  AND U25636 ( .A(n24892), .B(n24891), .Z(n25007) );
  NANDN U25637 ( .A(n24894), .B(n24893), .Z(n24898) );
  OR U25638 ( .A(n24896), .B(n24895), .Z(n24897) );
  NAND U25639 ( .A(n24898), .B(n24897), .Z(n25006) );
  XNOR U25640 ( .A(n25007), .B(n25006), .Z(n25008) );
  NAND U25641 ( .A(b[0]), .B(a[182]), .Z(n24899) );
  XNOR U25642 ( .A(b[1]), .B(n24899), .Z(n24901) );
  NANDN U25643 ( .A(b[0]), .B(a[181]), .Z(n24900) );
  NAND U25644 ( .A(n24901), .B(n24900), .Z(n24955) );
  NAND U25645 ( .A(n194), .B(n24902), .Z(n24904) );
  XOR U25646 ( .A(b[29]), .B(a[154]), .Z(n25033) );
  NAND U25647 ( .A(n38456), .B(n25033), .Z(n24903) );
  AND U25648 ( .A(n24904), .B(n24903), .Z(n24953) );
  AND U25649 ( .A(b[31]), .B(a[150]), .Z(n24952) );
  XNOR U25650 ( .A(n24953), .B(n24952), .Z(n24954) );
  XNOR U25651 ( .A(n24955), .B(n24954), .Z(n24994) );
  NAND U25652 ( .A(n38185), .B(n24905), .Z(n24907) );
  XOR U25653 ( .A(b[23]), .B(a[160]), .Z(n25036) );
  NAND U25654 ( .A(n38132), .B(n25036), .Z(n24906) );
  AND U25655 ( .A(n24907), .B(n24906), .Z(n25027) );
  NAND U25656 ( .A(n184), .B(n24908), .Z(n24910) );
  XOR U25657 ( .A(b[7]), .B(a[176]), .Z(n25039) );
  NAND U25658 ( .A(n36592), .B(n25039), .Z(n24909) );
  AND U25659 ( .A(n24910), .B(n24909), .Z(n25025) );
  NAND U25660 ( .A(n38289), .B(n24911), .Z(n24913) );
  XOR U25661 ( .A(b[25]), .B(a[158]), .Z(n25042) );
  NAND U25662 ( .A(n38247), .B(n25042), .Z(n24912) );
  NAND U25663 ( .A(n24913), .B(n24912), .Z(n25024) );
  XNOR U25664 ( .A(n25025), .B(n25024), .Z(n25026) );
  XOR U25665 ( .A(n25027), .B(n25026), .Z(n24995) );
  XNOR U25666 ( .A(n24994), .B(n24995), .Z(n24996) );
  NAND U25667 ( .A(n187), .B(n24914), .Z(n24916) );
  XOR U25668 ( .A(b[13]), .B(a[170]), .Z(n25045) );
  NAND U25669 ( .A(n37295), .B(n25045), .Z(n24915) );
  AND U25670 ( .A(n24916), .B(n24915), .Z(n24989) );
  NAND U25671 ( .A(n186), .B(n24917), .Z(n24919) );
  XOR U25672 ( .A(b[11]), .B(a[172]), .Z(n25048) );
  NAND U25673 ( .A(n37097), .B(n25048), .Z(n24918) );
  NAND U25674 ( .A(n24919), .B(n24918), .Z(n24988) );
  XNOR U25675 ( .A(n24989), .B(n24988), .Z(n24990) );
  NAND U25676 ( .A(n188), .B(n24920), .Z(n24922) );
  XOR U25677 ( .A(b[15]), .B(a[168]), .Z(n25051) );
  NAND U25678 ( .A(n37382), .B(n25051), .Z(n24921) );
  AND U25679 ( .A(n24922), .B(n24921), .Z(n24985) );
  NAND U25680 ( .A(n38064), .B(n24923), .Z(n24925) );
  XOR U25681 ( .A(b[21]), .B(a[162]), .Z(n25054) );
  NAND U25682 ( .A(n37993), .B(n25054), .Z(n24924) );
  AND U25683 ( .A(n24925), .B(n24924), .Z(n24983) );
  NAND U25684 ( .A(n185), .B(n24926), .Z(n24928) );
  XOR U25685 ( .A(b[9]), .B(a[174]), .Z(n25057) );
  NAND U25686 ( .A(n36805), .B(n25057), .Z(n24927) );
  NAND U25687 ( .A(n24928), .B(n24927), .Z(n24982) );
  XNOR U25688 ( .A(n24983), .B(n24982), .Z(n24984) );
  XOR U25689 ( .A(n24985), .B(n24984), .Z(n24991) );
  XOR U25690 ( .A(n24990), .B(n24991), .Z(n24997) );
  XOR U25691 ( .A(n24996), .B(n24997), .Z(n25009) );
  XNOR U25692 ( .A(n25008), .B(n25009), .Z(n25066) );
  XNOR U25693 ( .A(n25067), .B(n25066), .Z(n25068) );
  XOR U25694 ( .A(n25069), .B(n25068), .Z(n25073) );
  XNOR U25695 ( .A(n25072), .B(n25073), .Z(n25074) );
  XNOR U25696 ( .A(n25075), .B(n25074), .Z(n25080) );
  XOR U25697 ( .A(n25081), .B(n25080), .Z(n24947) );
  NANDN U25698 ( .A(n24930), .B(n24929), .Z(n24934) );
  NANDN U25699 ( .A(n24932), .B(n24931), .Z(n24933) );
  AND U25700 ( .A(n24934), .B(n24933), .Z(n24946) );
  XOR U25701 ( .A(n24947), .B(n24946), .Z(n24949) );
  XNOR U25702 ( .A(n24948), .B(n24949), .Z(n24940) );
  XNOR U25703 ( .A(n24941), .B(n24940), .Z(n24942) );
  XNOR U25704 ( .A(n24943), .B(n24942), .Z(n25084) );
  XNOR U25705 ( .A(sreg[406]), .B(n25084), .Z(n25086) );
  NANDN U25706 ( .A(sreg[405]), .B(n24935), .Z(n24939) );
  NAND U25707 ( .A(n24937), .B(n24936), .Z(n24938) );
  NAND U25708 ( .A(n24939), .B(n24938), .Z(n25085) );
  XNOR U25709 ( .A(n25086), .B(n25085), .Z(c[406]) );
  NANDN U25710 ( .A(n24941), .B(n24940), .Z(n24945) );
  NANDN U25711 ( .A(n24943), .B(n24942), .Z(n24944) );
  AND U25712 ( .A(n24945), .B(n24944), .Z(n25092) );
  NANDN U25713 ( .A(n24947), .B(n24946), .Z(n24951) );
  NANDN U25714 ( .A(n24949), .B(n24948), .Z(n24950) );
  AND U25715 ( .A(n24951), .B(n24950), .Z(n25090) );
  NANDN U25716 ( .A(n24953), .B(n24952), .Z(n24957) );
  NANDN U25717 ( .A(n24955), .B(n24954), .Z(n24956) );
  AND U25718 ( .A(n24957), .B(n24956), .Z(n25181) );
  NAND U25719 ( .A(n38385), .B(n24958), .Z(n24960) );
  XOR U25720 ( .A(b[27]), .B(a[157]), .Z(n25125) );
  NAND U25721 ( .A(n38343), .B(n25125), .Z(n24959) );
  AND U25722 ( .A(n24960), .B(n24959), .Z(n25188) );
  NAND U25723 ( .A(n183), .B(n24961), .Z(n24963) );
  XOR U25724 ( .A(b[5]), .B(a[179]), .Z(n25128) );
  NAND U25725 ( .A(n36296), .B(n25128), .Z(n24962) );
  AND U25726 ( .A(n24963), .B(n24962), .Z(n25186) );
  NAND U25727 ( .A(n190), .B(n24964), .Z(n24966) );
  XOR U25728 ( .A(b[19]), .B(a[165]), .Z(n25131) );
  NAND U25729 ( .A(n37821), .B(n25131), .Z(n24965) );
  NAND U25730 ( .A(n24966), .B(n24965), .Z(n25185) );
  XNOR U25731 ( .A(n25186), .B(n25185), .Z(n25187) );
  XNOR U25732 ( .A(n25188), .B(n25187), .Z(n25179) );
  NAND U25733 ( .A(n38470), .B(n24967), .Z(n24969) );
  XOR U25734 ( .A(b[31]), .B(a[153]), .Z(n25134) );
  NAND U25735 ( .A(n38453), .B(n25134), .Z(n24968) );
  AND U25736 ( .A(n24969), .B(n24968), .Z(n25146) );
  NAND U25737 ( .A(n181), .B(n24970), .Z(n24972) );
  XOR U25738 ( .A(b[3]), .B(a[181]), .Z(n25137) );
  NAND U25739 ( .A(n182), .B(n25137), .Z(n24971) );
  AND U25740 ( .A(n24972), .B(n24971), .Z(n25144) );
  NAND U25741 ( .A(n189), .B(n24973), .Z(n24975) );
  XOR U25742 ( .A(b[17]), .B(a[167]), .Z(n25140) );
  NAND U25743 ( .A(n37652), .B(n25140), .Z(n24974) );
  NAND U25744 ( .A(n24975), .B(n24974), .Z(n25143) );
  XNOR U25745 ( .A(n25144), .B(n25143), .Z(n25145) );
  XOR U25746 ( .A(n25146), .B(n25145), .Z(n25180) );
  XOR U25747 ( .A(n25179), .B(n25180), .Z(n25182) );
  XOR U25748 ( .A(n25181), .B(n25182), .Z(n25114) );
  NANDN U25749 ( .A(n24977), .B(n24976), .Z(n24981) );
  NANDN U25750 ( .A(n24979), .B(n24978), .Z(n24980) );
  AND U25751 ( .A(n24981), .B(n24980), .Z(n25167) );
  NANDN U25752 ( .A(n24983), .B(n24982), .Z(n24987) );
  NANDN U25753 ( .A(n24985), .B(n24984), .Z(n24986) );
  NAND U25754 ( .A(n24987), .B(n24986), .Z(n25168) );
  XNOR U25755 ( .A(n25167), .B(n25168), .Z(n25169) );
  NANDN U25756 ( .A(n24989), .B(n24988), .Z(n24993) );
  NANDN U25757 ( .A(n24991), .B(n24990), .Z(n24992) );
  NAND U25758 ( .A(n24993), .B(n24992), .Z(n25170) );
  XNOR U25759 ( .A(n25169), .B(n25170), .Z(n25113) );
  XNOR U25760 ( .A(n25114), .B(n25113), .Z(n25116) );
  NANDN U25761 ( .A(n24995), .B(n24994), .Z(n24999) );
  NANDN U25762 ( .A(n24997), .B(n24996), .Z(n24998) );
  AND U25763 ( .A(n24999), .B(n24998), .Z(n25115) );
  XOR U25764 ( .A(n25116), .B(n25115), .Z(n25229) );
  NANDN U25765 ( .A(n25001), .B(n25000), .Z(n25005) );
  NANDN U25766 ( .A(n25003), .B(n25002), .Z(n25004) );
  AND U25767 ( .A(n25005), .B(n25004), .Z(n25227) );
  NANDN U25768 ( .A(n25007), .B(n25006), .Z(n25011) );
  NANDN U25769 ( .A(n25009), .B(n25008), .Z(n25010) );
  AND U25770 ( .A(n25011), .B(n25010), .Z(n25110) );
  NANDN U25771 ( .A(n25013), .B(n25012), .Z(n25017) );
  OR U25772 ( .A(n25015), .B(n25014), .Z(n25016) );
  AND U25773 ( .A(n25017), .B(n25016), .Z(n25108) );
  NANDN U25774 ( .A(n25019), .B(n25018), .Z(n25023) );
  NANDN U25775 ( .A(n25021), .B(n25020), .Z(n25022) );
  AND U25776 ( .A(n25023), .B(n25022), .Z(n25174) );
  NANDN U25777 ( .A(n25025), .B(n25024), .Z(n25029) );
  NANDN U25778 ( .A(n25027), .B(n25026), .Z(n25028) );
  NAND U25779 ( .A(n25029), .B(n25028), .Z(n25173) );
  XNOR U25780 ( .A(n25174), .B(n25173), .Z(n25175) );
  NAND U25781 ( .A(b[0]), .B(a[183]), .Z(n25030) );
  XNOR U25782 ( .A(b[1]), .B(n25030), .Z(n25032) );
  NANDN U25783 ( .A(b[0]), .B(a[182]), .Z(n25031) );
  NAND U25784 ( .A(n25032), .B(n25031), .Z(n25122) );
  NAND U25785 ( .A(n194), .B(n25033), .Z(n25035) );
  XOR U25786 ( .A(b[29]), .B(a[155]), .Z(n25200) );
  NAND U25787 ( .A(n38456), .B(n25200), .Z(n25034) );
  AND U25788 ( .A(n25035), .B(n25034), .Z(n25120) );
  AND U25789 ( .A(b[31]), .B(a[151]), .Z(n25119) );
  XNOR U25790 ( .A(n25120), .B(n25119), .Z(n25121) );
  XNOR U25791 ( .A(n25122), .B(n25121), .Z(n25161) );
  NAND U25792 ( .A(n38185), .B(n25036), .Z(n25038) );
  XOR U25793 ( .A(b[23]), .B(a[161]), .Z(n25203) );
  NAND U25794 ( .A(n38132), .B(n25203), .Z(n25037) );
  AND U25795 ( .A(n25038), .B(n25037), .Z(n25194) );
  NAND U25796 ( .A(n184), .B(n25039), .Z(n25041) );
  XOR U25797 ( .A(b[7]), .B(a[177]), .Z(n25206) );
  NAND U25798 ( .A(n36592), .B(n25206), .Z(n25040) );
  AND U25799 ( .A(n25041), .B(n25040), .Z(n25192) );
  NAND U25800 ( .A(n38289), .B(n25042), .Z(n25044) );
  XOR U25801 ( .A(b[25]), .B(a[159]), .Z(n25209) );
  NAND U25802 ( .A(n38247), .B(n25209), .Z(n25043) );
  NAND U25803 ( .A(n25044), .B(n25043), .Z(n25191) );
  XNOR U25804 ( .A(n25192), .B(n25191), .Z(n25193) );
  XOR U25805 ( .A(n25194), .B(n25193), .Z(n25162) );
  XNOR U25806 ( .A(n25161), .B(n25162), .Z(n25163) );
  NAND U25807 ( .A(n187), .B(n25045), .Z(n25047) );
  XOR U25808 ( .A(b[13]), .B(a[171]), .Z(n25212) );
  NAND U25809 ( .A(n37295), .B(n25212), .Z(n25046) );
  AND U25810 ( .A(n25047), .B(n25046), .Z(n25156) );
  NAND U25811 ( .A(n186), .B(n25048), .Z(n25050) );
  XOR U25812 ( .A(b[11]), .B(a[173]), .Z(n25215) );
  NAND U25813 ( .A(n37097), .B(n25215), .Z(n25049) );
  NAND U25814 ( .A(n25050), .B(n25049), .Z(n25155) );
  XNOR U25815 ( .A(n25156), .B(n25155), .Z(n25157) );
  NAND U25816 ( .A(n188), .B(n25051), .Z(n25053) );
  XOR U25817 ( .A(b[15]), .B(a[169]), .Z(n25218) );
  NAND U25818 ( .A(n37382), .B(n25218), .Z(n25052) );
  AND U25819 ( .A(n25053), .B(n25052), .Z(n25152) );
  NAND U25820 ( .A(n38064), .B(n25054), .Z(n25056) );
  XOR U25821 ( .A(b[21]), .B(a[163]), .Z(n25221) );
  NAND U25822 ( .A(n37993), .B(n25221), .Z(n25055) );
  AND U25823 ( .A(n25056), .B(n25055), .Z(n25150) );
  NAND U25824 ( .A(n185), .B(n25057), .Z(n25059) );
  XOR U25825 ( .A(b[9]), .B(a[175]), .Z(n25224) );
  NAND U25826 ( .A(n36805), .B(n25224), .Z(n25058) );
  NAND U25827 ( .A(n25059), .B(n25058), .Z(n25149) );
  XNOR U25828 ( .A(n25150), .B(n25149), .Z(n25151) );
  XOR U25829 ( .A(n25152), .B(n25151), .Z(n25158) );
  XOR U25830 ( .A(n25157), .B(n25158), .Z(n25164) );
  XOR U25831 ( .A(n25163), .B(n25164), .Z(n25176) );
  XNOR U25832 ( .A(n25175), .B(n25176), .Z(n25107) );
  XNOR U25833 ( .A(n25108), .B(n25107), .Z(n25109) );
  XOR U25834 ( .A(n25110), .B(n25109), .Z(n25228) );
  XOR U25835 ( .A(n25227), .B(n25228), .Z(n25230) );
  XOR U25836 ( .A(n25229), .B(n25230), .Z(n25104) );
  NANDN U25837 ( .A(n25061), .B(n25060), .Z(n25065) );
  NAND U25838 ( .A(n25063), .B(n25062), .Z(n25064) );
  AND U25839 ( .A(n25065), .B(n25064), .Z(n25102) );
  NANDN U25840 ( .A(n25067), .B(n25066), .Z(n25071) );
  NANDN U25841 ( .A(n25069), .B(n25068), .Z(n25070) );
  AND U25842 ( .A(n25071), .B(n25070), .Z(n25101) );
  XNOR U25843 ( .A(n25102), .B(n25101), .Z(n25103) );
  XNOR U25844 ( .A(n25104), .B(n25103), .Z(n25095) );
  NANDN U25845 ( .A(n25073), .B(n25072), .Z(n25077) );
  NANDN U25846 ( .A(n25075), .B(n25074), .Z(n25076) );
  NAND U25847 ( .A(n25077), .B(n25076), .Z(n25096) );
  XNOR U25848 ( .A(n25095), .B(n25096), .Z(n25097) );
  NANDN U25849 ( .A(n25079), .B(n25078), .Z(n25083) );
  NAND U25850 ( .A(n25081), .B(n25080), .Z(n25082) );
  NAND U25851 ( .A(n25083), .B(n25082), .Z(n25098) );
  XNOR U25852 ( .A(n25097), .B(n25098), .Z(n25089) );
  XNOR U25853 ( .A(n25090), .B(n25089), .Z(n25091) );
  XNOR U25854 ( .A(n25092), .B(n25091), .Z(n25233) );
  XNOR U25855 ( .A(sreg[407]), .B(n25233), .Z(n25235) );
  NANDN U25856 ( .A(sreg[406]), .B(n25084), .Z(n25088) );
  NAND U25857 ( .A(n25086), .B(n25085), .Z(n25087) );
  NAND U25858 ( .A(n25088), .B(n25087), .Z(n25234) );
  XNOR U25859 ( .A(n25235), .B(n25234), .Z(c[407]) );
  NANDN U25860 ( .A(n25090), .B(n25089), .Z(n25094) );
  NANDN U25861 ( .A(n25092), .B(n25091), .Z(n25093) );
  AND U25862 ( .A(n25094), .B(n25093), .Z(n25241) );
  NANDN U25863 ( .A(n25096), .B(n25095), .Z(n25100) );
  NANDN U25864 ( .A(n25098), .B(n25097), .Z(n25099) );
  AND U25865 ( .A(n25100), .B(n25099), .Z(n25239) );
  NANDN U25866 ( .A(n25102), .B(n25101), .Z(n25106) );
  NANDN U25867 ( .A(n25104), .B(n25103), .Z(n25105) );
  AND U25868 ( .A(n25106), .B(n25105), .Z(n25247) );
  NANDN U25869 ( .A(n25108), .B(n25107), .Z(n25112) );
  NANDN U25870 ( .A(n25110), .B(n25109), .Z(n25111) );
  AND U25871 ( .A(n25112), .B(n25111), .Z(n25251) );
  NANDN U25872 ( .A(n25114), .B(n25113), .Z(n25118) );
  NAND U25873 ( .A(n25116), .B(n25115), .Z(n25117) );
  AND U25874 ( .A(n25118), .B(n25117), .Z(n25250) );
  XNOR U25875 ( .A(n25251), .B(n25250), .Z(n25253) );
  NANDN U25876 ( .A(n25120), .B(n25119), .Z(n25124) );
  NANDN U25877 ( .A(n25122), .B(n25121), .Z(n25123) );
  AND U25878 ( .A(n25124), .B(n25123), .Z(n25330) );
  NAND U25879 ( .A(n38385), .B(n25125), .Z(n25127) );
  XOR U25880 ( .A(b[27]), .B(a[158]), .Z(n25274) );
  NAND U25881 ( .A(n38343), .B(n25274), .Z(n25126) );
  AND U25882 ( .A(n25127), .B(n25126), .Z(n25337) );
  NAND U25883 ( .A(n183), .B(n25128), .Z(n25130) );
  XOR U25884 ( .A(b[5]), .B(a[180]), .Z(n25277) );
  NAND U25885 ( .A(n36296), .B(n25277), .Z(n25129) );
  AND U25886 ( .A(n25130), .B(n25129), .Z(n25335) );
  NAND U25887 ( .A(n190), .B(n25131), .Z(n25133) );
  XOR U25888 ( .A(b[19]), .B(a[166]), .Z(n25280) );
  NAND U25889 ( .A(n37821), .B(n25280), .Z(n25132) );
  NAND U25890 ( .A(n25133), .B(n25132), .Z(n25334) );
  XNOR U25891 ( .A(n25335), .B(n25334), .Z(n25336) );
  XNOR U25892 ( .A(n25337), .B(n25336), .Z(n25328) );
  NAND U25893 ( .A(n38470), .B(n25134), .Z(n25136) );
  XOR U25894 ( .A(b[31]), .B(a[154]), .Z(n25283) );
  NAND U25895 ( .A(n38453), .B(n25283), .Z(n25135) );
  AND U25896 ( .A(n25136), .B(n25135), .Z(n25295) );
  NAND U25897 ( .A(n181), .B(n25137), .Z(n25139) );
  XOR U25898 ( .A(b[3]), .B(a[182]), .Z(n25286) );
  NAND U25899 ( .A(n182), .B(n25286), .Z(n25138) );
  AND U25900 ( .A(n25139), .B(n25138), .Z(n25293) );
  NAND U25901 ( .A(n189), .B(n25140), .Z(n25142) );
  XOR U25902 ( .A(b[17]), .B(a[168]), .Z(n25289) );
  NAND U25903 ( .A(n37652), .B(n25289), .Z(n25141) );
  NAND U25904 ( .A(n25142), .B(n25141), .Z(n25292) );
  XNOR U25905 ( .A(n25293), .B(n25292), .Z(n25294) );
  XOR U25906 ( .A(n25295), .B(n25294), .Z(n25329) );
  XOR U25907 ( .A(n25328), .B(n25329), .Z(n25331) );
  XOR U25908 ( .A(n25330), .B(n25331), .Z(n25263) );
  NANDN U25909 ( .A(n25144), .B(n25143), .Z(n25148) );
  NANDN U25910 ( .A(n25146), .B(n25145), .Z(n25147) );
  AND U25911 ( .A(n25148), .B(n25147), .Z(n25316) );
  NANDN U25912 ( .A(n25150), .B(n25149), .Z(n25154) );
  NANDN U25913 ( .A(n25152), .B(n25151), .Z(n25153) );
  NAND U25914 ( .A(n25154), .B(n25153), .Z(n25317) );
  XNOR U25915 ( .A(n25316), .B(n25317), .Z(n25318) );
  NANDN U25916 ( .A(n25156), .B(n25155), .Z(n25160) );
  NANDN U25917 ( .A(n25158), .B(n25157), .Z(n25159) );
  NAND U25918 ( .A(n25160), .B(n25159), .Z(n25319) );
  XNOR U25919 ( .A(n25318), .B(n25319), .Z(n25262) );
  XNOR U25920 ( .A(n25263), .B(n25262), .Z(n25265) );
  NANDN U25921 ( .A(n25162), .B(n25161), .Z(n25166) );
  NANDN U25922 ( .A(n25164), .B(n25163), .Z(n25165) );
  AND U25923 ( .A(n25166), .B(n25165), .Z(n25264) );
  XOR U25924 ( .A(n25265), .B(n25264), .Z(n25379) );
  NANDN U25925 ( .A(n25168), .B(n25167), .Z(n25172) );
  NANDN U25926 ( .A(n25170), .B(n25169), .Z(n25171) );
  AND U25927 ( .A(n25172), .B(n25171), .Z(n25376) );
  NANDN U25928 ( .A(n25174), .B(n25173), .Z(n25178) );
  NANDN U25929 ( .A(n25176), .B(n25175), .Z(n25177) );
  AND U25930 ( .A(n25178), .B(n25177), .Z(n25259) );
  NANDN U25931 ( .A(n25180), .B(n25179), .Z(n25184) );
  OR U25932 ( .A(n25182), .B(n25181), .Z(n25183) );
  AND U25933 ( .A(n25184), .B(n25183), .Z(n25257) );
  NANDN U25934 ( .A(n25186), .B(n25185), .Z(n25190) );
  NANDN U25935 ( .A(n25188), .B(n25187), .Z(n25189) );
  AND U25936 ( .A(n25190), .B(n25189), .Z(n25323) );
  NANDN U25937 ( .A(n25192), .B(n25191), .Z(n25196) );
  NANDN U25938 ( .A(n25194), .B(n25193), .Z(n25195) );
  NAND U25939 ( .A(n25196), .B(n25195), .Z(n25322) );
  XNOR U25940 ( .A(n25323), .B(n25322), .Z(n25324) );
  NAND U25941 ( .A(b[0]), .B(a[184]), .Z(n25197) );
  XNOR U25942 ( .A(b[1]), .B(n25197), .Z(n25199) );
  NANDN U25943 ( .A(b[0]), .B(a[183]), .Z(n25198) );
  NAND U25944 ( .A(n25199), .B(n25198), .Z(n25271) );
  NAND U25945 ( .A(n194), .B(n25200), .Z(n25202) );
  XOR U25946 ( .A(b[29]), .B(a[156]), .Z(n25349) );
  NAND U25947 ( .A(n38456), .B(n25349), .Z(n25201) );
  AND U25948 ( .A(n25202), .B(n25201), .Z(n25269) );
  AND U25949 ( .A(b[31]), .B(a[152]), .Z(n25268) );
  XNOR U25950 ( .A(n25269), .B(n25268), .Z(n25270) );
  XNOR U25951 ( .A(n25271), .B(n25270), .Z(n25310) );
  NAND U25952 ( .A(n38185), .B(n25203), .Z(n25205) );
  XOR U25953 ( .A(b[23]), .B(a[162]), .Z(n25352) );
  NAND U25954 ( .A(n38132), .B(n25352), .Z(n25204) );
  AND U25955 ( .A(n25205), .B(n25204), .Z(n25343) );
  NAND U25956 ( .A(n184), .B(n25206), .Z(n25208) );
  XOR U25957 ( .A(b[7]), .B(a[178]), .Z(n25355) );
  NAND U25958 ( .A(n36592), .B(n25355), .Z(n25207) );
  AND U25959 ( .A(n25208), .B(n25207), .Z(n25341) );
  NAND U25960 ( .A(n38289), .B(n25209), .Z(n25211) );
  XOR U25961 ( .A(b[25]), .B(a[160]), .Z(n25358) );
  NAND U25962 ( .A(n38247), .B(n25358), .Z(n25210) );
  NAND U25963 ( .A(n25211), .B(n25210), .Z(n25340) );
  XNOR U25964 ( .A(n25341), .B(n25340), .Z(n25342) );
  XOR U25965 ( .A(n25343), .B(n25342), .Z(n25311) );
  XNOR U25966 ( .A(n25310), .B(n25311), .Z(n25312) );
  NAND U25967 ( .A(n187), .B(n25212), .Z(n25214) );
  XOR U25968 ( .A(b[13]), .B(a[172]), .Z(n25361) );
  NAND U25969 ( .A(n37295), .B(n25361), .Z(n25213) );
  AND U25970 ( .A(n25214), .B(n25213), .Z(n25305) );
  NAND U25971 ( .A(n186), .B(n25215), .Z(n25217) );
  XOR U25972 ( .A(b[11]), .B(a[174]), .Z(n25364) );
  NAND U25973 ( .A(n37097), .B(n25364), .Z(n25216) );
  NAND U25974 ( .A(n25217), .B(n25216), .Z(n25304) );
  XNOR U25975 ( .A(n25305), .B(n25304), .Z(n25306) );
  NAND U25976 ( .A(n188), .B(n25218), .Z(n25220) );
  XOR U25977 ( .A(b[15]), .B(a[170]), .Z(n25367) );
  NAND U25978 ( .A(n37382), .B(n25367), .Z(n25219) );
  AND U25979 ( .A(n25220), .B(n25219), .Z(n25301) );
  NAND U25980 ( .A(n38064), .B(n25221), .Z(n25223) );
  XOR U25981 ( .A(b[21]), .B(a[164]), .Z(n25370) );
  NAND U25982 ( .A(n37993), .B(n25370), .Z(n25222) );
  AND U25983 ( .A(n25223), .B(n25222), .Z(n25299) );
  NAND U25984 ( .A(n185), .B(n25224), .Z(n25226) );
  XOR U25985 ( .A(b[9]), .B(a[176]), .Z(n25373) );
  NAND U25986 ( .A(n36805), .B(n25373), .Z(n25225) );
  NAND U25987 ( .A(n25226), .B(n25225), .Z(n25298) );
  XNOR U25988 ( .A(n25299), .B(n25298), .Z(n25300) );
  XOR U25989 ( .A(n25301), .B(n25300), .Z(n25307) );
  XOR U25990 ( .A(n25306), .B(n25307), .Z(n25313) );
  XOR U25991 ( .A(n25312), .B(n25313), .Z(n25325) );
  XNOR U25992 ( .A(n25324), .B(n25325), .Z(n25256) );
  XNOR U25993 ( .A(n25257), .B(n25256), .Z(n25258) );
  XOR U25994 ( .A(n25259), .B(n25258), .Z(n25377) );
  XNOR U25995 ( .A(n25376), .B(n25377), .Z(n25378) );
  XNOR U25996 ( .A(n25379), .B(n25378), .Z(n25252) );
  XOR U25997 ( .A(n25253), .B(n25252), .Z(n25245) );
  NANDN U25998 ( .A(n25228), .B(n25227), .Z(n25232) );
  OR U25999 ( .A(n25230), .B(n25229), .Z(n25231) );
  AND U26000 ( .A(n25232), .B(n25231), .Z(n25244) );
  XNOR U26001 ( .A(n25245), .B(n25244), .Z(n25246) );
  XNOR U26002 ( .A(n25247), .B(n25246), .Z(n25238) );
  XNOR U26003 ( .A(n25239), .B(n25238), .Z(n25240) );
  XNOR U26004 ( .A(n25241), .B(n25240), .Z(n25382) );
  XNOR U26005 ( .A(sreg[408]), .B(n25382), .Z(n25384) );
  NANDN U26006 ( .A(sreg[407]), .B(n25233), .Z(n25237) );
  NAND U26007 ( .A(n25235), .B(n25234), .Z(n25236) );
  NAND U26008 ( .A(n25237), .B(n25236), .Z(n25383) );
  XNOR U26009 ( .A(n25384), .B(n25383), .Z(c[408]) );
  NANDN U26010 ( .A(n25239), .B(n25238), .Z(n25243) );
  NANDN U26011 ( .A(n25241), .B(n25240), .Z(n25242) );
  AND U26012 ( .A(n25243), .B(n25242), .Z(n25390) );
  NANDN U26013 ( .A(n25245), .B(n25244), .Z(n25249) );
  NANDN U26014 ( .A(n25247), .B(n25246), .Z(n25248) );
  AND U26015 ( .A(n25249), .B(n25248), .Z(n25388) );
  NANDN U26016 ( .A(n25251), .B(n25250), .Z(n25255) );
  NAND U26017 ( .A(n25253), .B(n25252), .Z(n25254) );
  AND U26018 ( .A(n25255), .B(n25254), .Z(n25395) );
  NANDN U26019 ( .A(n25257), .B(n25256), .Z(n25261) );
  NANDN U26020 ( .A(n25259), .B(n25258), .Z(n25260) );
  AND U26021 ( .A(n25261), .B(n25260), .Z(n25526) );
  NANDN U26022 ( .A(n25263), .B(n25262), .Z(n25267) );
  NAND U26023 ( .A(n25265), .B(n25264), .Z(n25266) );
  AND U26024 ( .A(n25267), .B(n25266), .Z(n25525) );
  XNOR U26025 ( .A(n25526), .B(n25525), .Z(n25528) );
  NANDN U26026 ( .A(n25269), .B(n25268), .Z(n25273) );
  NANDN U26027 ( .A(n25271), .B(n25270), .Z(n25272) );
  AND U26028 ( .A(n25273), .B(n25272), .Z(n25473) );
  NAND U26029 ( .A(n38385), .B(n25274), .Z(n25276) );
  XOR U26030 ( .A(b[27]), .B(a[159]), .Z(n25417) );
  NAND U26031 ( .A(n38343), .B(n25417), .Z(n25275) );
  AND U26032 ( .A(n25276), .B(n25275), .Z(n25480) );
  NAND U26033 ( .A(n183), .B(n25277), .Z(n25279) );
  XOR U26034 ( .A(b[5]), .B(a[181]), .Z(n25420) );
  NAND U26035 ( .A(n36296), .B(n25420), .Z(n25278) );
  AND U26036 ( .A(n25279), .B(n25278), .Z(n25478) );
  NAND U26037 ( .A(n190), .B(n25280), .Z(n25282) );
  XOR U26038 ( .A(b[19]), .B(a[167]), .Z(n25423) );
  NAND U26039 ( .A(n37821), .B(n25423), .Z(n25281) );
  NAND U26040 ( .A(n25282), .B(n25281), .Z(n25477) );
  XNOR U26041 ( .A(n25478), .B(n25477), .Z(n25479) );
  XNOR U26042 ( .A(n25480), .B(n25479), .Z(n25471) );
  NAND U26043 ( .A(n38470), .B(n25283), .Z(n25285) );
  XOR U26044 ( .A(b[31]), .B(a[155]), .Z(n25426) );
  NAND U26045 ( .A(n38453), .B(n25426), .Z(n25284) );
  AND U26046 ( .A(n25285), .B(n25284), .Z(n25438) );
  NAND U26047 ( .A(n181), .B(n25286), .Z(n25288) );
  XOR U26048 ( .A(b[3]), .B(a[183]), .Z(n25429) );
  NAND U26049 ( .A(n182), .B(n25429), .Z(n25287) );
  AND U26050 ( .A(n25288), .B(n25287), .Z(n25436) );
  NAND U26051 ( .A(n189), .B(n25289), .Z(n25291) );
  XOR U26052 ( .A(b[17]), .B(a[169]), .Z(n25432) );
  NAND U26053 ( .A(n37652), .B(n25432), .Z(n25290) );
  NAND U26054 ( .A(n25291), .B(n25290), .Z(n25435) );
  XNOR U26055 ( .A(n25436), .B(n25435), .Z(n25437) );
  XOR U26056 ( .A(n25438), .B(n25437), .Z(n25472) );
  XOR U26057 ( .A(n25471), .B(n25472), .Z(n25474) );
  XOR U26058 ( .A(n25473), .B(n25474), .Z(n25406) );
  NANDN U26059 ( .A(n25293), .B(n25292), .Z(n25297) );
  NANDN U26060 ( .A(n25295), .B(n25294), .Z(n25296) );
  AND U26061 ( .A(n25297), .B(n25296), .Z(n25459) );
  NANDN U26062 ( .A(n25299), .B(n25298), .Z(n25303) );
  NANDN U26063 ( .A(n25301), .B(n25300), .Z(n25302) );
  NAND U26064 ( .A(n25303), .B(n25302), .Z(n25460) );
  XNOR U26065 ( .A(n25459), .B(n25460), .Z(n25461) );
  NANDN U26066 ( .A(n25305), .B(n25304), .Z(n25309) );
  NANDN U26067 ( .A(n25307), .B(n25306), .Z(n25308) );
  NAND U26068 ( .A(n25309), .B(n25308), .Z(n25462) );
  XNOR U26069 ( .A(n25461), .B(n25462), .Z(n25405) );
  XNOR U26070 ( .A(n25406), .B(n25405), .Z(n25408) );
  NANDN U26071 ( .A(n25311), .B(n25310), .Z(n25315) );
  NANDN U26072 ( .A(n25313), .B(n25312), .Z(n25314) );
  AND U26073 ( .A(n25315), .B(n25314), .Z(n25407) );
  XOR U26074 ( .A(n25408), .B(n25407), .Z(n25522) );
  NANDN U26075 ( .A(n25317), .B(n25316), .Z(n25321) );
  NANDN U26076 ( .A(n25319), .B(n25318), .Z(n25320) );
  AND U26077 ( .A(n25321), .B(n25320), .Z(n25519) );
  NANDN U26078 ( .A(n25323), .B(n25322), .Z(n25327) );
  NANDN U26079 ( .A(n25325), .B(n25324), .Z(n25326) );
  AND U26080 ( .A(n25327), .B(n25326), .Z(n25402) );
  NANDN U26081 ( .A(n25329), .B(n25328), .Z(n25333) );
  OR U26082 ( .A(n25331), .B(n25330), .Z(n25332) );
  AND U26083 ( .A(n25333), .B(n25332), .Z(n25400) );
  NANDN U26084 ( .A(n25335), .B(n25334), .Z(n25339) );
  NANDN U26085 ( .A(n25337), .B(n25336), .Z(n25338) );
  AND U26086 ( .A(n25339), .B(n25338), .Z(n25466) );
  NANDN U26087 ( .A(n25341), .B(n25340), .Z(n25345) );
  NANDN U26088 ( .A(n25343), .B(n25342), .Z(n25344) );
  NAND U26089 ( .A(n25345), .B(n25344), .Z(n25465) );
  XNOR U26090 ( .A(n25466), .B(n25465), .Z(n25467) );
  NAND U26091 ( .A(b[0]), .B(a[185]), .Z(n25346) );
  XNOR U26092 ( .A(b[1]), .B(n25346), .Z(n25348) );
  NANDN U26093 ( .A(b[0]), .B(a[184]), .Z(n25347) );
  NAND U26094 ( .A(n25348), .B(n25347), .Z(n25414) );
  NAND U26095 ( .A(n194), .B(n25349), .Z(n25351) );
  XOR U26096 ( .A(b[29]), .B(a[157]), .Z(n25492) );
  NAND U26097 ( .A(n38456), .B(n25492), .Z(n25350) );
  AND U26098 ( .A(n25351), .B(n25350), .Z(n25412) );
  AND U26099 ( .A(b[31]), .B(a[153]), .Z(n25411) );
  XNOR U26100 ( .A(n25412), .B(n25411), .Z(n25413) );
  XNOR U26101 ( .A(n25414), .B(n25413), .Z(n25453) );
  NAND U26102 ( .A(n38185), .B(n25352), .Z(n25354) );
  XOR U26103 ( .A(b[23]), .B(a[163]), .Z(n25495) );
  NAND U26104 ( .A(n38132), .B(n25495), .Z(n25353) );
  AND U26105 ( .A(n25354), .B(n25353), .Z(n25486) );
  NAND U26106 ( .A(n184), .B(n25355), .Z(n25357) );
  XOR U26107 ( .A(b[7]), .B(a[179]), .Z(n25498) );
  NAND U26108 ( .A(n36592), .B(n25498), .Z(n25356) );
  AND U26109 ( .A(n25357), .B(n25356), .Z(n25484) );
  NAND U26110 ( .A(n38289), .B(n25358), .Z(n25360) );
  XOR U26111 ( .A(b[25]), .B(a[161]), .Z(n25501) );
  NAND U26112 ( .A(n38247), .B(n25501), .Z(n25359) );
  NAND U26113 ( .A(n25360), .B(n25359), .Z(n25483) );
  XNOR U26114 ( .A(n25484), .B(n25483), .Z(n25485) );
  XOR U26115 ( .A(n25486), .B(n25485), .Z(n25454) );
  XNOR U26116 ( .A(n25453), .B(n25454), .Z(n25455) );
  NAND U26117 ( .A(n187), .B(n25361), .Z(n25363) );
  XOR U26118 ( .A(b[13]), .B(a[173]), .Z(n25504) );
  NAND U26119 ( .A(n37295), .B(n25504), .Z(n25362) );
  AND U26120 ( .A(n25363), .B(n25362), .Z(n25448) );
  NAND U26121 ( .A(n186), .B(n25364), .Z(n25366) );
  XOR U26122 ( .A(b[11]), .B(a[175]), .Z(n25507) );
  NAND U26123 ( .A(n37097), .B(n25507), .Z(n25365) );
  NAND U26124 ( .A(n25366), .B(n25365), .Z(n25447) );
  XNOR U26125 ( .A(n25448), .B(n25447), .Z(n25449) );
  NAND U26126 ( .A(n188), .B(n25367), .Z(n25369) );
  XOR U26127 ( .A(b[15]), .B(a[171]), .Z(n25510) );
  NAND U26128 ( .A(n37382), .B(n25510), .Z(n25368) );
  AND U26129 ( .A(n25369), .B(n25368), .Z(n25444) );
  NAND U26130 ( .A(n38064), .B(n25370), .Z(n25372) );
  XOR U26131 ( .A(b[21]), .B(a[165]), .Z(n25513) );
  NAND U26132 ( .A(n37993), .B(n25513), .Z(n25371) );
  AND U26133 ( .A(n25372), .B(n25371), .Z(n25442) );
  NAND U26134 ( .A(n185), .B(n25373), .Z(n25375) );
  XOR U26135 ( .A(b[9]), .B(a[177]), .Z(n25516) );
  NAND U26136 ( .A(n36805), .B(n25516), .Z(n25374) );
  NAND U26137 ( .A(n25375), .B(n25374), .Z(n25441) );
  XNOR U26138 ( .A(n25442), .B(n25441), .Z(n25443) );
  XOR U26139 ( .A(n25444), .B(n25443), .Z(n25450) );
  XOR U26140 ( .A(n25449), .B(n25450), .Z(n25456) );
  XOR U26141 ( .A(n25455), .B(n25456), .Z(n25468) );
  XNOR U26142 ( .A(n25467), .B(n25468), .Z(n25399) );
  XNOR U26143 ( .A(n25400), .B(n25399), .Z(n25401) );
  XOR U26144 ( .A(n25402), .B(n25401), .Z(n25520) );
  XNOR U26145 ( .A(n25519), .B(n25520), .Z(n25521) );
  XNOR U26146 ( .A(n25522), .B(n25521), .Z(n25527) );
  XOR U26147 ( .A(n25528), .B(n25527), .Z(n25394) );
  NANDN U26148 ( .A(n25377), .B(n25376), .Z(n25381) );
  NANDN U26149 ( .A(n25379), .B(n25378), .Z(n25380) );
  AND U26150 ( .A(n25381), .B(n25380), .Z(n25393) );
  XOR U26151 ( .A(n25394), .B(n25393), .Z(n25396) );
  XNOR U26152 ( .A(n25395), .B(n25396), .Z(n25387) );
  XNOR U26153 ( .A(n25388), .B(n25387), .Z(n25389) );
  XNOR U26154 ( .A(n25390), .B(n25389), .Z(n25531) );
  XNOR U26155 ( .A(sreg[409]), .B(n25531), .Z(n25533) );
  NANDN U26156 ( .A(sreg[408]), .B(n25382), .Z(n25386) );
  NAND U26157 ( .A(n25384), .B(n25383), .Z(n25385) );
  NAND U26158 ( .A(n25386), .B(n25385), .Z(n25532) );
  XNOR U26159 ( .A(n25533), .B(n25532), .Z(c[409]) );
  NANDN U26160 ( .A(n25388), .B(n25387), .Z(n25392) );
  NANDN U26161 ( .A(n25390), .B(n25389), .Z(n25391) );
  AND U26162 ( .A(n25392), .B(n25391), .Z(n25539) );
  NANDN U26163 ( .A(n25394), .B(n25393), .Z(n25398) );
  NANDN U26164 ( .A(n25396), .B(n25395), .Z(n25397) );
  AND U26165 ( .A(n25398), .B(n25397), .Z(n25537) );
  NANDN U26166 ( .A(n25400), .B(n25399), .Z(n25404) );
  NANDN U26167 ( .A(n25402), .B(n25401), .Z(n25403) );
  AND U26168 ( .A(n25404), .B(n25403), .Z(n25549) );
  NANDN U26169 ( .A(n25406), .B(n25405), .Z(n25410) );
  NAND U26170 ( .A(n25408), .B(n25407), .Z(n25409) );
  AND U26171 ( .A(n25410), .B(n25409), .Z(n25548) );
  XNOR U26172 ( .A(n25549), .B(n25548), .Z(n25551) );
  NANDN U26173 ( .A(n25412), .B(n25411), .Z(n25416) );
  NANDN U26174 ( .A(n25414), .B(n25413), .Z(n25415) );
  AND U26175 ( .A(n25416), .B(n25415), .Z(n25628) );
  NAND U26176 ( .A(n38385), .B(n25417), .Z(n25419) );
  XOR U26177 ( .A(b[27]), .B(a[160]), .Z(n25572) );
  NAND U26178 ( .A(n38343), .B(n25572), .Z(n25418) );
  AND U26179 ( .A(n25419), .B(n25418), .Z(n25635) );
  NAND U26180 ( .A(n183), .B(n25420), .Z(n25422) );
  XOR U26181 ( .A(b[5]), .B(a[182]), .Z(n25575) );
  NAND U26182 ( .A(n36296), .B(n25575), .Z(n25421) );
  AND U26183 ( .A(n25422), .B(n25421), .Z(n25633) );
  NAND U26184 ( .A(n190), .B(n25423), .Z(n25425) );
  XOR U26185 ( .A(b[19]), .B(a[168]), .Z(n25578) );
  NAND U26186 ( .A(n37821), .B(n25578), .Z(n25424) );
  NAND U26187 ( .A(n25425), .B(n25424), .Z(n25632) );
  XNOR U26188 ( .A(n25633), .B(n25632), .Z(n25634) );
  XNOR U26189 ( .A(n25635), .B(n25634), .Z(n25626) );
  NAND U26190 ( .A(n38470), .B(n25426), .Z(n25428) );
  XOR U26191 ( .A(b[31]), .B(a[156]), .Z(n25581) );
  NAND U26192 ( .A(n38453), .B(n25581), .Z(n25427) );
  AND U26193 ( .A(n25428), .B(n25427), .Z(n25593) );
  NAND U26194 ( .A(n181), .B(n25429), .Z(n25431) );
  XOR U26195 ( .A(b[3]), .B(a[184]), .Z(n25584) );
  NAND U26196 ( .A(n182), .B(n25584), .Z(n25430) );
  AND U26197 ( .A(n25431), .B(n25430), .Z(n25591) );
  NAND U26198 ( .A(n189), .B(n25432), .Z(n25434) );
  XOR U26199 ( .A(b[17]), .B(a[170]), .Z(n25587) );
  NAND U26200 ( .A(n37652), .B(n25587), .Z(n25433) );
  NAND U26201 ( .A(n25434), .B(n25433), .Z(n25590) );
  XNOR U26202 ( .A(n25591), .B(n25590), .Z(n25592) );
  XOR U26203 ( .A(n25593), .B(n25592), .Z(n25627) );
  XOR U26204 ( .A(n25626), .B(n25627), .Z(n25629) );
  XOR U26205 ( .A(n25628), .B(n25629), .Z(n25561) );
  NANDN U26206 ( .A(n25436), .B(n25435), .Z(n25440) );
  NANDN U26207 ( .A(n25438), .B(n25437), .Z(n25439) );
  AND U26208 ( .A(n25440), .B(n25439), .Z(n25614) );
  NANDN U26209 ( .A(n25442), .B(n25441), .Z(n25446) );
  NANDN U26210 ( .A(n25444), .B(n25443), .Z(n25445) );
  NAND U26211 ( .A(n25446), .B(n25445), .Z(n25615) );
  XNOR U26212 ( .A(n25614), .B(n25615), .Z(n25616) );
  NANDN U26213 ( .A(n25448), .B(n25447), .Z(n25452) );
  NANDN U26214 ( .A(n25450), .B(n25449), .Z(n25451) );
  NAND U26215 ( .A(n25452), .B(n25451), .Z(n25617) );
  XNOR U26216 ( .A(n25616), .B(n25617), .Z(n25560) );
  XNOR U26217 ( .A(n25561), .B(n25560), .Z(n25563) );
  NANDN U26218 ( .A(n25454), .B(n25453), .Z(n25458) );
  NANDN U26219 ( .A(n25456), .B(n25455), .Z(n25457) );
  AND U26220 ( .A(n25458), .B(n25457), .Z(n25562) );
  XOR U26221 ( .A(n25563), .B(n25562), .Z(n25677) );
  NANDN U26222 ( .A(n25460), .B(n25459), .Z(n25464) );
  NANDN U26223 ( .A(n25462), .B(n25461), .Z(n25463) );
  AND U26224 ( .A(n25464), .B(n25463), .Z(n25674) );
  NANDN U26225 ( .A(n25466), .B(n25465), .Z(n25470) );
  NANDN U26226 ( .A(n25468), .B(n25467), .Z(n25469) );
  AND U26227 ( .A(n25470), .B(n25469), .Z(n25557) );
  NANDN U26228 ( .A(n25472), .B(n25471), .Z(n25476) );
  OR U26229 ( .A(n25474), .B(n25473), .Z(n25475) );
  AND U26230 ( .A(n25476), .B(n25475), .Z(n25555) );
  NANDN U26231 ( .A(n25478), .B(n25477), .Z(n25482) );
  NANDN U26232 ( .A(n25480), .B(n25479), .Z(n25481) );
  AND U26233 ( .A(n25482), .B(n25481), .Z(n25621) );
  NANDN U26234 ( .A(n25484), .B(n25483), .Z(n25488) );
  NANDN U26235 ( .A(n25486), .B(n25485), .Z(n25487) );
  NAND U26236 ( .A(n25488), .B(n25487), .Z(n25620) );
  XNOR U26237 ( .A(n25621), .B(n25620), .Z(n25622) );
  NAND U26238 ( .A(b[0]), .B(a[186]), .Z(n25489) );
  XNOR U26239 ( .A(b[1]), .B(n25489), .Z(n25491) );
  NANDN U26240 ( .A(b[0]), .B(a[185]), .Z(n25490) );
  NAND U26241 ( .A(n25491), .B(n25490), .Z(n25569) );
  NAND U26242 ( .A(n194), .B(n25492), .Z(n25494) );
  XOR U26243 ( .A(b[29]), .B(a[158]), .Z(n25647) );
  NAND U26244 ( .A(n38456), .B(n25647), .Z(n25493) );
  AND U26245 ( .A(n25494), .B(n25493), .Z(n25567) );
  AND U26246 ( .A(b[31]), .B(a[154]), .Z(n25566) );
  XNOR U26247 ( .A(n25567), .B(n25566), .Z(n25568) );
  XNOR U26248 ( .A(n25569), .B(n25568), .Z(n25608) );
  NAND U26249 ( .A(n38185), .B(n25495), .Z(n25497) );
  XOR U26250 ( .A(b[23]), .B(a[164]), .Z(n25650) );
  NAND U26251 ( .A(n38132), .B(n25650), .Z(n25496) );
  AND U26252 ( .A(n25497), .B(n25496), .Z(n25641) );
  NAND U26253 ( .A(n184), .B(n25498), .Z(n25500) );
  XOR U26254 ( .A(b[7]), .B(a[180]), .Z(n25653) );
  NAND U26255 ( .A(n36592), .B(n25653), .Z(n25499) );
  AND U26256 ( .A(n25500), .B(n25499), .Z(n25639) );
  NAND U26257 ( .A(n38289), .B(n25501), .Z(n25503) );
  XOR U26258 ( .A(b[25]), .B(a[162]), .Z(n25656) );
  NAND U26259 ( .A(n38247), .B(n25656), .Z(n25502) );
  NAND U26260 ( .A(n25503), .B(n25502), .Z(n25638) );
  XNOR U26261 ( .A(n25639), .B(n25638), .Z(n25640) );
  XOR U26262 ( .A(n25641), .B(n25640), .Z(n25609) );
  XNOR U26263 ( .A(n25608), .B(n25609), .Z(n25610) );
  NAND U26264 ( .A(n187), .B(n25504), .Z(n25506) );
  XOR U26265 ( .A(b[13]), .B(a[174]), .Z(n25659) );
  NAND U26266 ( .A(n37295), .B(n25659), .Z(n25505) );
  AND U26267 ( .A(n25506), .B(n25505), .Z(n25603) );
  NAND U26268 ( .A(n186), .B(n25507), .Z(n25509) );
  XOR U26269 ( .A(b[11]), .B(a[176]), .Z(n25662) );
  NAND U26270 ( .A(n37097), .B(n25662), .Z(n25508) );
  NAND U26271 ( .A(n25509), .B(n25508), .Z(n25602) );
  XNOR U26272 ( .A(n25603), .B(n25602), .Z(n25604) );
  NAND U26273 ( .A(n188), .B(n25510), .Z(n25512) );
  XOR U26274 ( .A(b[15]), .B(a[172]), .Z(n25665) );
  NAND U26275 ( .A(n37382), .B(n25665), .Z(n25511) );
  AND U26276 ( .A(n25512), .B(n25511), .Z(n25599) );
  NAND U26277 ( .A(n38064), .B(n25513), .Z(n25515) );
  XOR U26278 ( .A(b[21]), .B(a[166]), .Z(n25668) );
  NAND U26279 ( .A(n37993), .B(n25668), .Z(n25514) );
  AND U26280 ( .A(n25515), .B(n25514), .Z(n25597) );
  NAND U26281 ( .A(n185), .B(n25516), .Z(n25518) );
  XOR U26282 ( .A(b[9]), .B(a[178]), .Z(n25671) );
  NAND U26283 ( .A(n36805), .B(n25671), .Z(n25517) );
  NAND U26284 ( .A(n25518), .B(n25517), .Z(n25596) );
  XNOR U26285 ( .A(n25597), .B(n25596), .Z(n25598) );
  XOR U26286 ( .A(n25599), .B(n25598), .Z(n25605) );
  XOR U26287 ( .A(n25604), .B(n25605), .Z(n25611) );
  XOR U26288 ( .A(n25610), .B(n25611), .Z(n25623) );
  XNOR U26289 ( .A(n25622), .B(n25623), .Z(n25554) );
  XNOR U26290 ( .A(n25555), .B(n25554), .Z(n25556) );
  XOR U26291 ( .A(n25557), .B(n25556), .Z(n25675) );
  XNOR U26292 ( .A(n25674), .B(n25675), .Z(n25676) );
  XNOR U26293 ( .A(n25677), .B(n25676), .Z(n25550) );
  XOR U26294 ( .A(n25551), .B(n25550), .Z(n25543) );
  NANDN U26295 ( .A(n25520), .B(n25519), .Z(n25524) );
  NANDN U26296 ( .A(n25522), .B(n25521), .Z(n25523) );
  AND U26297 ( .A(n25524), .B(n25523), .Z(n25542) );
  XNOR U26298 ( .A(n25543), .B(n25542), .Z(n25544) );
  NANDN U26299 ( .A(n25526), .B(n25525), .Z(n25530) );
  NAND U26300 ( .A(n25528), .B(n25527), .Z(n25529) );
  NAND U26301 ( .A(n25530), .B(n25529), .Z(n25545) );
  XNOR U26302 ( .A(n25544), .B(n25545), .Z(n25536) );
  XNOR U26303 ( .A(n25537), .B(n25536), .Z(n25538) );
  XNOR U26304 ( .A(n25539), .B(n25538), .Z(n25680) );
  XNOR U26305 ( .A(sreg[410]), .B(n25680), .Z(n25682) );
  NANDN U26306 ( .A(sreg[409]), .B(n25531), .Z(n25535) );
  NAND U26307 ( .A(n25533), .B(n25532), .Z(n25534) );
  NAND U26308 ( .A(n25535), .B(n25534), .Z(n25681) );
  XNOR U26309 ( .A(n25682), .B(n25681), .Z(c[410]) );
  NANDN U26310 ( .A(n25537), .B(n25536), .Z(n25541) );
  NANDN U26311 ( .A(n25539), .B(n25538), .Z(n25540) );
  AND U26312 ( .A(n25541), .B(n25540), .Z(n25688) );
  NANDN U26313 ( .A(n25543), .B(n25542), .Z(n25547) );
  NANDN U26314 ( .A(n25545), .B(n25544), .Z(n25546) );
  AND U26315 ( .A(n25547), .B(n25546), .Z(n25686) );
  NANDN U26316 ( .A(n25549), .B(n25548), .Z(n25553) );
  NAND U26317 ( .A(n25551), .B(n25550), .Z(n25552) );
  AND U26318 ( .A(n25553), .B(n25552), .Z(n25693) );
  NANDN U26319 ( .A(n25555), .B(n25554), .Z(n25559) );
  NANDN U26320 ( .A(n25557), .B(n25556), .Z(n25558) );
  AND U26321 ( .A(n25559), .B(n25558), .Z(n25698) );
  NANDN U26322 ( .A(n25561), .B(n25560), .Z(n25565) );
  NAND U26323 ( .A(n25563), .B(n25562), .Z(n25564) );
  AND U26324 ( .A(n25565), .B(n25564), .Z(n25697) );
  XNOR U26325 ( .A(n25698), .B(n25697), .Z(n25700) );
  NANDN U26326 ( .A(n25567), .B(n25566), .Z(n25571) );
  NANDN U26327 ( .A(n25569), .B(n25568), .Z(n25570) );
  AND U26328 ( .A(n25571), .B(n25570), .Z(n25777) );
  NAND U26329 ( .A(n38385), .B(n25572), .Z(n25574) );
  XOR U26330 ( .A(b[27]), .B(a[161]), .Z(n25721) );
  NAND U26331 ( .A(n38343), .B(n25721), .Z(n25573) );
  AND U26332 ( .A(n25574), .B(n25573), .Z(n25784) );
  NAND U26333 ( .A(n183), .B(n25575), .Z(n25577) );
  XOR U26334 ( .A(b[5]), .B(a[183]), .Z(n25724) );
  NAND U26335 ( .A(n36296), .B(n25724), .Z(n25576) );
  AND U26336 ( .A(n25577), .B(n25576), .Z(n25782) );
  NAND U26337 ( .A(n190), .B(n25578), .Z(n25580) );
  XOR U26338 ( .A(b[19]), .B(a[169]), .Z(n25727) );
  NAND U26339 ( .A(n37821), .B(n25727), .Z(n25579) );
  NAND U26340 ( .A(n25580), .B(n25579), .Z(n25781) );
  XNOR U26341 ( .A(n25782), .B(n25781), .Z(n25783) );
  XNOR U26342 ( .A(n25784), .B(n25783), .Z(n25775) );
  NAND U26343 ( .A(n38470), .B(n25581), .Z(n25583) );
  XOR U26344 ( .A(b[31]), .B(a[157]), .Z(n25730) );
  NAND U26345 ( .A(n38453), .B(n25730), .Z(n25582) );
  AND U26346 ( .A(n25583), .B(n25582), .Z(n25742) );
  NAND U26347 ( .A(n181), .B(n25584), .Z(n25586) );
  XOR U26348 ( .A(b[3]), .B(a[185]), .Z(n25733) );
  NAND U26349 ( .A(n182), .B(n25733), .Z(n25585) );
  AND U26350 ( .A(n25586), .B(n25585), .Z(n25740) );
  NAND U26351 ( .A(n189), .B(n25587), .Z(n25589) );
  XOR U26352 ( .A(b[17]), .B(a[171]), .Z(n25736) );
  NAND U26353 ( .A(n37652), .B(n25736), .Z(n25588) );
  NAND U26354 ( .A(n25589), .B(n25588), .Z(n25739) );
  XNOR U26355 ( .A(n25740), .B(n25739), .Z(n25741) );
  XOR U26356 ( .A(n25742), .B(n25741), .Z(n25776) );
  XOR U26357 ( .A(n25775), .B(n25776), .Z(n25778) );
  XOR U26358 ( .A(n25777), .B(n25778), .Z(n25710) );
  NANDN U26359 ( .A(n25591), .B(n25590), .Z(n25595) );
  NANDN U26360 ( .A(n25593), .B(n25592), .Z(n25594) );
  AND U26361 ( .A(n25595), .B(n25594), .Z(n25763) );
  NANDN U26362 ( .A(n25597), .B(n25596), .Z(n25601) );
  NANDN U26363 ( .A(n25599), .B(n25598), .Z(n25600) );
  NAND U26364 ( .A(n25601), .B(n25600), .Z(n25764) );
  XNOR U26365 ( .A(n25763), .B(n25764), .Z(n25765) );
  NANDN U26366 ( .A(n25603), .B(n25602), .Z(n25607) );
  NANDN U26367 ( .A(n25605), .B(n25604), .Z(n25606) );
  NAND U26368 ( .A(n25607), .B(n25606), .Z(n25766) );
  XNOR U26369 ( .A(n25765), .B(n25766), .Z(n25709) );
  XNOR U26370 ( .A(n25710), .B(n25709), .Z(n25712) );
  NANDN U26371 ( .A(n25609), .B(n25608), .Z(n25613) );
  NANDN U26372 ( .A(n25611), .B(n25610), .Z(n25612) );
  AND U26373 ( .A(n25613), .B(n25612), .Z(n25711) );
  XOR U26374 ( .A(n25712), .B(n25711), .Z(n25826) );
  NANDN U26375 ( .A(n25615), .B(n25614), .Z(n25619) );
  NANDN U26376 ( .A(n25617), .B(n25616), .Z(n25618) );
  AND U26377 ( .A(n25619), .B(n25618), .Z(n25823) );
  NANDN U26378 ( .A(n25621), .B(n25620), .Z(n25625) );
  NANDN U26379 ( .A(n25623), .B(n25622), .Z(n25624) );
  AND U26380 ( .A(n25625), .B(n25624), .Z(n25706) );
  NANDN U26381 ( .A(n25627), .B(n25626), .Z(n25631) );
  OR U26382 ( .A(n25629), .B(n25628), .Z(n25630) );
  AND U26383 ( .A(n25631), .B(n25630), .Z(n25704) );
  NANDN U26384 ( .A(n25633), .B(n25632), .Z(n25637) );
  NANDN U26385 ( .A(n25635), .B(n25634), .Z(n25636) );
  AND U26386 ( .A(n25637), .B(n25636), .Z(n25770) );
  NANDN U26387 ( .A(n25639), .B(n25638), .Z(n25643) );
  NANDN U26388 ( .A(n25641), .B(n25640), .Z(n25642) );
  NAND U26389 ( .A(n25643), .B(n25642), .Z(n25769) );
  XNOR U26390 ( .A(n25770), .B(n25769), .Z(n25771) );
  NAND U26391 ( .A(b[0]), .B(a[187]), .Z(n25644) );
  XNOR U26392 ( .A(b[1]), .B(n25644), .Z(n25646) );
  NANDN U26393 ( .A(b[0]), .B(a[186]), .Z(n25645) );
  NAND U26394 ( .A(n25646), .B(n25645), .Z(n25718) );
  NAND U26395 ( .A(n194), .B(n25647), .Z(n25649) );
  XOR U26396 ( .A(b[29]), .B(a[159]), .Z(n25796) );
  NAND U26397 ( .A(n38456), .B(n25796), .Z(n25648) );
  AND U26398 ( .A(n25649), .B(n25648), .Z(n25716) );
  AND U26399 ( .A(b[31]), .B(a[155]), .Z(n25715) );
  XNOR U26400 ( .A(n25716), .B(n25715), .Z(n25717) );
  XNOR U26401 ( .A(n25718), .B(n25717), .Z(n25757) );
  NAND U26402 ( .A(n38185), .B(n25650), .Z(n25652) );
  XOR U26403 ( .A(b[23]), .B(a[165]), .Z(n25799) );
  NAND U26404 ( .A(n38132), .B(n25799), .Z(n25651) );
  AND U26405 ( .A(n25652), .B(n25651), .Z(n25790) );
  NAND U26406 ( .A(n184), .B(n25653), .Z(n25655) );
  XOR U26407 ( .A(b[7]), .B(a[181]), .Z(n25802) );
  NAND U26408 ( .A(n36592), .B(n25802), .Z(n25654) );
  AND U26409 ( .A(n25655), .B(n25654), .Z(n25788) );
  NAND U26410 ( .A(n38289), .B(n25656), .Z(n25658) );
  XOR U26411 ( .A(b[25]), .B(a[163]), .Z(n25805) );
  NAND U26412 ( .A(n38247), .B(n25805), .Z(n25657) );
  NAND U26413 ( .A(n25658), .B(n25657), .Z(n25787) );
  XNOR U26414 ( .A(n25788), .B(n25787), .Z(n25789) );
  XOR U26415 ( .A(n25790), .B(n25789), .Z(n25758) );
  XNOR U26416 ( .A(n25757), .B(n25758), .Z(n25759) );
  NAND U26417 ( .A(n187), .B(n25659), .Z(n25661) );
  XOR U26418 ( .A(b[13]), .B(a[175]), .Z(n25808) );
  NAND U26419 ( .A(n37295), .B(n25808), .Z(n25660) );
  AND U26420 ( .A(n25661), .B(n25660), .Z(n25752) );
  NAND U26421 ( .A(n186), .B(n25662), .Z(n25664) );
  XOR U26422 ( .A(b[11]), .B(a[177]), .Z(n25811) );
  NAND U26423 ( .A(n37097), .B(n25811), .Z(n25663) );
  NAND U26424 ( .A(n25664), .B(n25663), .Z(n25751) );
  XNOR U26425 ( .A(n25752), .B(n25751), .Z(n25753) );
  NAND U26426 ( .A(n188), .B(n25665), .Z(n25667) );
  XOR U26427 ( .A(b[15]), .B(a[173]), .Z(n25814) );
  NAND U26428 ( .A(n37382), .B(n25814), .Z(n25666) );
  AND U26429 ( .A(n25667), .B(n25666), .Z(n25748) );
  NAND U26430 ( .A(n38064), .B(n25668), .Z(n25670) );
  XOR U26431 ( .A(b[21]), .B(a[167]), .Z(n25817) );
  NAND U26432 ( .A(n37993), .B(n25817), .Z(n25669) );
  AND U26433 ( .A(n25670), .B(n25669), .Z(n25746) );
  NAND U26434 ( .A(n185), .B(n25671), .Z(n25673) );
  XOR U26435 ( .A(b[9]), .B(a[179]), .Z(n25820) );
  NAND U26436 ( .A(n36805), .B(n25820), .Z(n25672) );
  NAND U26437 ( .A(n25673), .B(n25672), .Z(n25745) );
  XNOR U26438 ( .A(n25746), .B(n25745), .Z(n25747) );
  XOR U26439 ( .A(n25748), .B(n25747), .Z(n25754) );
  XOR U26440 ( .A(n25753), .B(n25754), .Z(n25760) );
  XOR U26441 ( .A(n25759), .B(n25760), .Z(n25772) );
  XNOR U26442 ( .A(n25771), .B(n25772), .Z(n25703) );
  XNOR U26443 ( .A(n25704), .B(n25703), .Z(n25705) );
  XOR U26444 ( .A(n25706), .B(n25705), .Z(n25824) );
  XNOR U26445 ( .A(n25823), .B(n25824), .Z(n25825) );
  XNOR U26446 ( .A(n25826), .B(n25825), .Z(n25699) );
  XOR U26447 ( .A(n25700), .B(n25699), .Z(n25692) );
  NANDN U26448 ( .A(n25675), .B(n25674), .Z(n25679) );
  NANDN U26449 ( .A(n25677), .B(n25676), .Z(n25678) );
  AND U26450 ( .A(n25679), .B(n25678), .Z(n25691) );
  XOR U26451 ( .A(n25692), .B(n25691), .Z(n25694) );
  XNOR U26452 ( .A(n25693), .B(n25694), .Z(n25685) );
  XNOR U26453 ( .A(n25686), .B(n25685), .Z(n25687) );
  XNOR U26454 ( .A(n25688), .B(n25687), .Z(n25829) );
  XNOR U26455 ( .A(sreg[411]), .B(n25829), .Z(n25831) );
  NANDN U26456 ( .A(sreg[410]), .B(n25680), .Z(n25684) );
  NAND U26457 ( .A(n25682), .B(n25681), .Z(n25683) );
  NAND U26458 ( .A(n25684), .B(n25683), .Z(n25830) );
  XNOR U26459 ( .A(n25831), .B(n25830), .Z(c[411]) );
  NANDN U26460 ( .A(n25686), .B(n25685), .Z(n25690) );
  NANDN U26461 ( .A(n25688), .B(n25687), .Z(n25689) );
  AND U26462 ( .A(n25690), .B(n25689), .Z(n25837) );
  NANDN U26463 ( .A(n25692), .B(n25691), .Z(n25696) );
  NANDN U26464 ( .A(n25694), .B(n25693), .Z(n25695) );
  AND U26465 ( .A(n25696), .B(n25695), .Z(n25835) );
  NANDN U26466 ( .A(n25698), .B(n25697), .Z(n25702) );
  NAND U26467 ( .A(n25700), .B(n25699), .Z(n25701) );
  AND U26468 ( .A(n25702), .B(n25701), .Z(n25842) );
  NANDN U26469 ( .A(n25704), .B(n25703), .Z(n25708) );
  NANDN U26470 ( .A(n25706), .B(n25705), .Z(n25707) );
  AND U26471 ( .A(n25708), .B(n25707), .Z(n25847) );
  NANDN U26472 ( .A(n25710), .B(n25709), .Z(n25714) );
  NAND U26473 ( .A(n25712), .B(n25711), .Z(n25713) );
  AND U26474 ( .A(n25714), .B(n25713), .Z(n25846) );
  XNOR U26475 ( .A(n25847), .B(n25846), .Z(n25849) );
  NANDN U26476 ( .A(n25716), .B(n25715), .Z(n25720) );
  NANDN U26477 ( .A(n25718), .B(n25717), .Z(n25719) );
  AND U26478 ( .A(n25720), .B(n25719), .Z(n25924) );
  NAND U26479 ( .A(n38385), .B(n25721), .Z(n25723) );
  XOR U26480 ( .A(b[27]), .B(a[162]), .Z(n25870) );
  NAND U26481 ( .A(n38343), .B(n25870), .Z(n25722) );
  AND U26482 ( .A(n25723), .B(n25722), .Z(n25931) );
  NAND U26483 ( .A(n183), .B(n25724), .Z(n25726) );
  XOR U26484 ( .A(b[5]), .B(a[184]), .Z(n25873) );
  NAND U26485 ( .A(n36296), .B(n25873), .Z(n25725) );
  AND U26486 ( .A(n25726), .B(n25725), .Z(n25929) );
  NAND U26487 ( .A(n190), .B(n25727), .Z(n25729) );
  XOR U26488 ( .A(b[19]), .B(a[170]), .Z(n25876) );
  NAND U26489 ( .A(n37821), .B(n25876), .Z(n25728) );
  NAND U26490 ( .A(n25729), .B(n25728), .Z(n25928) );
  XNOR U26491 ( .A(n25929), .B(n25928), .Z(n25930) );
  XNOR U26492 ( .A(n25931), .B(n25930), .Z(n25922) );
  NAND U26493 ( .A(n38470), .B(n25730), .Z(n25732) );
  XOR U26494 ( .A(b[31]), .B(a[158]), .Z(n25879) );
  NAND U26495 ( .A(n38453), .B(n25879), .Z(n25731) );
  AND U26496 ( .A(n25732), .B(n25731), .Z(n25891) );
  NAND U26497 ( .A(n181), .B(n25733), .Z(n25735) );
  XOR U26498 ( .A(b[3]), .B(a[186]), .Z(n25882) );
  NAND U26499 ( .A(n182), .B(n25882), .Z(n25734) );
  AND U26500 ( .A(n25735), .B(n25734), .Z(n25889) );
  NAND U26501 ( .A(n189), .B(n25736), .Z(n25738) );
  XOR U26502 ( .A(b[17]), .B(a[172]), .Z(n25885) );
  NAND U26503 ( .A(n37652), .B(n25885), .Z(n25737) );
  NAND U26504 ( .A(n25738), .B(n25737), .Z(n25888) );
  XNOR U26505 ( .A(n25889), .B(n25888), .Z(n25890) );
  XOR U26506 ( .A(n25891), .B(n25890), .Z(n25923) );
  XOR U26507 ( .A(n25922), .B(n25923), .Z(n25925) );
  XOR U26508 ( .A(n25924), .B(n25925), .Z(n25859) );
  NANDN U26509 ( .A(n25740), .B(n25739), .Z(n25744) );
  NANDN U26510 ( .A(n25742), .B(n25741), .Z(n25743) );
  AND U26511 ( .A(n25744), .B(n25743), .Z(n25912) );
  NANDN U26512 ( .A(n25746), .B(n25745), .Z(n25750) );
  NANDN U26513 ( .A(n25748), .B(n25747), .Z(n25749) );
  NAND U26514 ( .A(n25750), .B(n25749), .Z(n25913) );
  XNOR U26515 ( .A(n25912), .B(n25913), .Z(n25914) );
  NANDN U26516 ( .A(n25752), .B(n25751), .Z(n25756) );
  NANDN U26517 ( .A(n25754), .B(n25753), .Z(n25755) );
  NAND U26518 ( .A(n25756), .B(n25755), .Z(n25915) );
  XNOR U26519 ( .A(n25914), .B(n25915), .Z(n25858) );
  XNOR U26520 ( .A(n25859), .B(n25858), .Z(n25861) );
  NANDN U26521 ( .A(n25758), .B(n25757), .Z(n25762) );
  NANDN U26522 ( .A(n25760), .B(n25759), .Z(n25761) );
  AND U26523 ( .A(n25762), .B(n25761), .Z(n25860) );
  XOR U26524 ( .A(n25861), .B(n25860), .Z(n25973) );
  NANDN U26525 ( .A(n25764), .B(n25763), .Z(n25768) );
  NANDN U26526 ( .A(n25766), .B(n25765), .Z(n25767) );
  AND U26527 ( .A(n25768), .B(n25767), .Z(n25970) );
  NANDN U26528 ( .A(n25770), .B(n25769), .Z(n25774) );
  NANDN U26529 ( .A(n25772), .B(n25771), .Z(n25773) );
  AND U26530 ( .A(n25774), .B(n25773), .Z(n25855) );
  NANDN U26531 ( .A(n25776), .B(n25775), .Z(n25780) );
  OR U26532 ( .A(n25778), .B(n25777), .Z(n25779) );
  AND U26533 ( .A(n25780), .B(n25779), .Z(n25853) );
  NANDN U26534 ( .A(n25782), .B(n25781), .Z(n25786) );
  NANDN U26535 ( .A(n25784), .B(n25783), .Z(n25785) );
  AND U26536 ( .A(n25786), .B(n25785), .Z(n25919) );
  NANDN U26537 ( .A(n25788), .B(n25787), .Z(n25792) );
  NANDN U26538 ( .A(n25790), .B(n25789), .Z(n25791) );
  NAND U26539 ( .A(n25792), .B(n25791), .Z(n25918) );
  XNOR U26540 ( .A(n25919), .B(n25918), .Z(n25921) );
  NAND U26541 ( .A(b[0]), .B(a[188]), .Z(n25793) );
  XNOR U26542 ( .A(b[1]), .B(n25793), .Z(n25795) );
  NANDN U26543 ( .A(b[0]), .B(a[187]), .Z(n25794) );
  NAND U26544 ( .A(n25795), .B(n25794), .Z(n25867) );
  NAND U26545 ( .A(n194), .B(n25796), .Z(n25798) );
  XOR U26546 ( .A(b[29]), .B(a[160]), .Z(n25943) );
  NAND U26547 ( .A(n38456), .B(n25943), .Z(n25797) );
  AND U26548 ( .A(n25798), .B(n25797), .Z(n25865) );
  AND U26549 ( .A(b[31]), .B(a[156]), .Z(n25864) );
  XNOR U26550 ( .A(n25865), .B(n25864), .Z(n25866) );
  XNOR U26551 ( .A(n25867), .B(n25866), .Z(n25907) );
  NAND U26552 ( .A(n38185), .B(n25799), .Z(n25801) );
  XOR U26553 ( .A(b[23]), .B(a[166]), .Z(n25946) );
  NAND U26554 ( .A(n38132), .B(n25946), .Z(n25800) );
  AND U26555 ( .A(n25801), .B(n25800), .Z(n25936) );
  NAND U26556 ( .A(n184), .B(n25802), .Z(n25804) );
  XOR U26557 ( .A(b[7]), .B(a[182]), .Z(n25949) );
  NAND U26558 ( .A(n36592), .B(n25949), .Z(n25803) );
  AND U26559 ( .A(n25804), .B(n25803), .Z(n25935) );
  NAND U26560 ( .A(n38289), .B(n25805), .Z(n25807) );
  XOR U26561 ( .A(b[25]), .B(a[164]), .Z(n25952) );
  NAND U26562 ( .A(n38247), .B(n25952), .Z(n25806) );
  NAND U26563 ( .A(n25807), .B(n25806), .Z(n25934) );
  XOR U26564 ( .A(n25935), .B(n25934), .Z(n25937) );
  XOR U26565 ( .A(n25936), .B(n25937), .Z(n25906) );
  XOR U26566 ( .A(n25907), .B(n25906), .Z(n25909) );
  NAND U26567 ( .A(n187), .B(n25808), .Z(n25810) );
  XOR U26568 ( .A(b[13]), .B(a[176]), .Z(n25955) );
  NAND U26569 ( .A(n37295), .B(n25955), .Z(n25809) );
  AND U26570 ( .A(n25810), .B(n25809), .Z(n25901) );
  NAND U26571 ( .A(n186), .B(n25811), .Z(n25813) );
  XOR U26572 ( .A(b[11]), .B(a[178]), .Z(n25958) );
  NAND U26573 ( .A(n37097), .B(n25958), .Z(n25812) );
  NAND U26574 ( .A(n25813), .B(n25812), .Z(n25900) );
  XNOR U26575 ( .A(n25901), .B(n25900), .Z(n25903) );
  NAND U26576 ( .A(n188), .B(n25814), .Z(n25816) );
  XOR U26577 ( .A(b[15]), .B(a[174]), .Z(n25961) );
  NAND U26578 ( .A(n37382), .B(n25961), .Z(n25815) );
  AND U26579 ( .A(n25816), .B(n25815), .Z(n25897) );
  NAND U26580 ( .A(n38064), .B(n25817), .Z(n25819) );
  XOR U26581 ( .A(b[21]), .B(a[168]), .Z(n25964) );
  NAND U26582 ( .A(n37993), .B(n25964), .Z(n25818) );
  AND U26583 ( .A(n25819), .B(n25818), .Z(n25895) );
  NAND U26584 ( .A(n185), .B(n25820), .Z(n25822) );
  XOR U26585 ( .A(b[9]), .B(a[180]), .Z(n25967) );
  NAND U26586 ( .A(n36805), .B(n25967), .Z(n25821) );
  NAND U26587 ( .A(n25822), .B(n25821), .Z(n25894) );
  XNOR U26588 ( .A(n25895), .B(n25894), .Z(n25896) );
  XNOR U26589 ( .A(n25897), .B(n25896), .Z(n25902) );
  XOR U26590 ( .A(n25903), .B(n25902), .Z(n25908) );
  XNOR U26591 ( .A(n25909), .B(n25908), .Z(n25920) );
  XNOR U26592 ( .A(n25921), .B(n25920), .Z(n25852) );
  XNOR U26593 ( .A(n25853), .B(n25852), .Z(n25854) );
  XOR U26594 ( .A(n25855), .B(n25854), .Z(n25971) );
  XNOR U26595 ( .A(n25970), .B(n25971), .Z(n25972) );
  XNOR U26596 ( .A(n25973), .B(n25972), .Z(n25848) );
  XOR U26597 ( .A(n25849), .B(n25848), .Z(n25841) );
  NANDN U26598 ( .A(n25824), .B(n25823), .Z(n25828) );
  NANDN U26599 ( .A(n25826), .B(n25825), .Z(n25827) );
  AND U26600 ( .A(n25828), .B(n25827), .Z(n25840) );
  XOR U26601 ( .A(n25841), .B(n25840), .Z(n25843) );
  XNOR U26602 ( .A(n25842), .B(n25843), .Z(n25834) );
  XNOR U26603 ( .A(n25835), .B(n25834), .Z(n25836) );
  XNOR U26604 ( .A(n25837), .B(n25836), .Z(n25976) );
  XNOR U26605 ( .A(sreg[412]), .B(n25976), .Z(n25978) );
  NANDN U26606 ( .A(sreg[411]), .B(n25829), .Z(n25833) );
  NAND U26607 ( .A(n25831), .B(n25830), .Z(n25832) );
  NAND U26608 ( .A(n25833), .B(n25832), .Z(n25977) );
  XNOR U26609 ( .A(n25978), .B(n25977), .Z(c[412]) );
  NANDN U26610 ( .A(n25835), .B(n25834), .Z(n25839) );
  NANDN U26611 ( .A(n25837), .B(n25836), .Z(n25838) );
  AND U26612 ( .A(n25839), .B(n25838), .Z(n25984) );
  NANDN U26613 ( .A(n25841), .B(n25840), .Z(n25845) );
  NANDN U26614 ( .A(n25843), .B(n25842), .Z(n25844) );
  AND U26615 ( .A(n25845), .B(n25844), .Z(n25982) );
  NANDN U26616 ( .A(n25847), .B(n25846), .Z(n25851) );
  NAND U26617 ( .A(n25849), .B(n25848), .Z(n25850) );
  AND U26618 ( .A(n25851), .B(n25850), .Z(n25989) );
  NANDN U26619 ( .A(n25853), .B(n25852), .Z(n25857) );
  NANDN U26620 ( .A(n25855), .B(n25854), .Z(n25856) );
  AND U26621 ( .A(n25857), .B(n25856), .Z(n26118) );
  NANDN U26622 ( .A(n25859), .B(n25858), .Z(n25863) );
  NAND U26623 ( .A(n25861), .B(n25860), .Z(n25862) );
  AND U26624 ( .A(n25863), .B(n25862), .Z(n26117) );
  XNOR U26625 ( .A(n26118), .B(n26117), .Z(n26120) );
  NANDN U26626 ( .A(n25865), .B(n25864), .Z(n25869) );
  NANDN U26627 ( .A(n25867), .B(n25866), .Z(n25868) );
  AND U26628 ( .A(n25869), .B(n25868), .Z(n26053) );
  NAND U26629 ( .A(n38385), .B(n25870), .Z(n25872) );
  XOR U26630 ( .A(b[27]), .B(a[163]), .Z(n25999) );
  NAND U26631 ( .A(n38343), .B(n25999), .Z(n25871) );
  AND U26632 ( .A(n25872), .B(n25871), .Z(n26060) );
  NAND U26633 ( .A(n183), .B(n25873), .Z(n25875) );
  XOR U26634 ( .A(b[5]), .B(a[185]), .Z(n26002) );
  NAND U26635 ( .A(n36296), .B(n26002), .Z(n25874) );
  AND U26636 ( .A(n25875), .B(n25874), .Z(n26058) );
  NAND U26637 ( .A(n190), .B(n25876), .Z(n25878) );
  XOR U26638 ( .A(b[19]), .B(a[171]), .Z(n26005) );
  NAND U26639 ( .A(n37821), .B(n26005), .Z(n25877) );
  NAND U26640 ( .A(n25878), .B(n25877), .Z(n26057) );
  XNOR U26641 ( .A(n26058), .B(n26057), .Z(n26059) );
  XNOR U26642 ( .A(n26060), .B(n26059), .Z(n26051) );
  NAND U26643 ( .A(n38470), .B(n25879), .Z(n25881) );
  XOR U26644 ( .A(b[31]), .B(a[159]), .Z(n26008) );
  NAND U26645 ( .A(n38453), .B(n26008), .Z(n25880) );
  AND U26646 ( .A(n25881), .B(n25880), .Z(n26020) );
  NAND U26647 ( .A(n181), .B(n25882), .Z(n25884) );
  XOR U26648 ( .A(b[3]), .B(a[187]), .Z(n26011) );
  NAND U26649 ( .A(n182), .B(n26011), .Z(n25883) );
  AND U26650 ( .A(n25884), .B(n25883), .Z(n26018) );
  NAND U26651 ( .A(n189), .B(n25885), .Z(n25887) );
  XOR U26652 ( .A(b[17]), .B(a[173]), .Z(n26014) );
  NAND U26653 ( .A(n37652), .B(n26014), .Z(n25886) );
  NAND U26654 ( .A(n25887), .B(n25886), .Z(n26017) );
  XNOR U26655 ( .A(n26018), .B(n26017), .Z(n26019) );
  XOR U26656 ( .A(n26020), .B(n26019), .Z(n26052) );
  XOR U26657 ( .A(n26051), .B(n26052), .Z(n26054) );
  XOR U26658 ( .A(n26053), .B(n26054), .Z(n26100) );
  NANDN U26659 ( .A(n25889), .B(n25888), .Z(n25893) );
  NANDN U26660 ( .A(n25891), .B(n25890), .Z(n25892) );
  AND U26661 ( .A(n25893), .B(n25892), .Z(n26041) );
  NANDN U26662 ( .A(n25895), .B(n25894), .Z(n25899) );
  NANDN U26663 ( .A(n25897), .B(n25896), .Z(n25898) );
  NAND U26664 ( .A(n25899), .B(n25898), .Z(n26042) );
  XNOR U26665 ( .A(n26041), .B(n26042), .Z(n26043) );
  NANDN U26666 ( .A(n25901), .B(n25900), .Z(n25905) );
  NAND U26667 ( .A(n25903), .B(n25902), .Z(n25904) );
  NAND U26668 ( .A(n25905), .B(n25904), .Z(n26044) );
  XNOR U26669 ( .A(n26043), .B(n26044), .Z(n26099) );
  XNOR U26670 ( .A(n26100), .B(n26099), .Z(n26102) );
  NAND U26671 ( .A(n25907), .B(n25906), .Z(n25911) );
  NAND U26672 ( .A(n25909), .B(n25908), .Z(n25910) );
  AND U26673 ( .A(n25911), .B(n25910), .Z(n26101) );
  XOR U26674 ( .A(n26102), .B(n26101), .Z(n26114) );
  NANDN U26675 ( .A(n25913), .B(n25912), .Z(n25917) );
  NANDN U26676 ( .A(n25915), .B(n25914), .Z(n25916) );
  AND U26677 ( .A(n25917), .B(n25916), .Z(n26111) );
  NANDN U26678 ( .A(n25923), .B(n25922), .Z(n25927) );
  OR U26679 ( .A(n25925), .B(n25924), .Z(n25926) );
  AND U26680 ( .A(n25927), .B(n25926), .Z(n26106) );
  NANDN U26681 ( .A(n25929), .B(n25928), .Z(n25933) );
  NANDN U26682 ( .A(n25931), .B(n25930), .Z(n25932) );
  AND U26683 ( .A(n25933), .B(n25932), .Z(n26048) );
  NANDN U26684 ( .A(n25935), .B(n25934), .Z(n25939) );
  OR U26685 ( .A(n25937), .B(n25936), .Z(n25938) );
  NAND U26686 ( .A(n25939), .B(n25938), .Z(n26047) );
  XNOR U26687 ( .A(n26048), .B(n26047), .Z(n26050) );
  NAND U26688 ( .A(b[0]), .B(a[189]), .Z(n25940) );
  XNOR U26689 ( .A(b[1]), .B(n25940), .Z(n25942) );
  NANDN U26690 ( .A(b[0]), .B(a[188]), .Z(n25941) );
  NAND U26691 ( .A(n25942), .B(n25941), .Z(n25996) );
  NAND U26692 ( .A(n194), .B(n25943), .Z(n25945) );
  XOR U26693 ( .A(b[29]), .B(a[161]), .Z(n26072) );
  NAND U26694 ( .A(n38456), .B(n26072), .Z(n25944) );
  AND U26695 ( .A(n25945), .B(n25944), .Z(n25994) );
  AND U26696 ( .A(b[31]), .B(a[157]), .Z(n25993) );
  XNOR U26697 ( .A(n25994), .B(n25993), .Z(n25995) );
  XNOR U26698 ( .A(n25996), .B(n25995), .Z(n26036) );
  NAND U26699 ( .A(n38185), .B(n25946), .Z(n25948) );
  XOR U26700 ( .A(b[23]), .B(a[167]), .Z(n26075) );
  NAND U26701 ( .A(n38132), .B(n26075), .Z(n25947) );
  AND U26702 ( .A(n25948), .B(n25947), .Z(n26065) );
  NAND U26703 ( .A(n184), .B(n25949), .Z(n25951) );
  XOR U26704 ( .A(b[7]), .B(a[183]), .Z(n26078) );
  NAND U26705 ( .A(n36592), .B(n26078), .Z(n25950) );
  AND U26706 ( .A(n25951), .B(n25950), .Z(n26064) );
  NAND U26707 ( .A(n38289), .B(n25952), .Z(n25954) );
  XOR U26708 ( .A(b[25]), .B(a[165]), .Z(n26081) );
  NAND U26709 ( .A(n38247), .B(n26081), .Z(n25953) );
  NAND U26710 ( .A(n25954), .B(n25953), .Z(n26063) );
  XOR U26711 ( .A(n26064), .B(n26063), .Z(n26066) );
  XOR U26712 ( .A(n26065), .B(n26066), .Z(n26035) );
  XOR U26713 ( .A(n26036), .B(n26035), .Z(n26038) );
  NAND U26714 ( .A(n187), .B(n25955), .Z(n25957) );
  XOR U26715 ( .A(b[13]), .B(a[177]), .Z(n26084) );
  NAND U26716 ( .A(n37295), .B(n26084), .Z(n25956) );
  AND U26717 ( .A(n25957), .B(n25956), .Z(n26030) );
  NAND U26718 ( .A(n186), .B(n25958), .Z(n25960) );
  XOR U26719 ( .A(b[11]), .B(a[179]), .Z(n26087) );
  NAND U26720 ( .A(n37097), .B(n26087), .Z(n25959) );
  NAND U26721 ( .A(n25960), .B(n25959), .Z(n26029) );
  XNOR U26722 ( .A(n26030), .B(n26029), .Z(n26032) );
  NAND U26723 ( .A(n188), .B(n25961), .Z(n25963) );
  XOR U26724 ( .A(b[15]), .B(a[175]), .Z(n26090) );
  NAND U26725 ( .A(n37382), .B(n26090), .Z(n25962) );
  AND U26726 ( .A(n25963), .B(n25962), .Z(n26026) );
  NAND U26727 ( .A(n38064), .B(n25964), .Z(n25966) );
  XOR U26728 ( .A(b[21]), .B(a[169]), .Z(n26093) );
  NAND U26729 ( .A(n37993), .B(n26093), .Z(n25965) );
  AND U26730 ( .A(n25966), .B(n25965), .Z(n26024) );
  NAND U26731 ( .A(n185), .B(n25967), .Z(n25969) );
  XOR U26732 ( .A(b[9]), .B(a[181]), .Z(n26096) );
  NAND U26733 ( .A(n36805), .B(n26096), .Z(n25968) );
  NAND U26734 ( .A(n25969), .B(n25968), .Z(n26023) );
  XNOR U26735 ( .A(n26024), .B(n26023), .Z(n26025) );
  XNOR U26736 ( .A(n26026), .B(n26025), .Z(n26031) );
  XOR U26737 ( .A(n26032), .B(n26031), .Z(n26037) );
  XNOR U26738 ( .A(n26038), .B(n26037), .Z(n26049) );
  XNOR U26739 ( .A(n26050), .B(n26049), .Z(n26105) );
  XNOR U26740 ( .A(n26106), .B(n26105), .Z(n26107) );
  XOR U26741 ( .A(n26108), .B(n26107), .Z(n26112) );
  XNOR U26742 ( .A(n26111), .B(n26112), .Z(n26113) );
  XNOR U26743 ( .A(n26114), .B(n26113), .Z(n26119) );
  XOR U26744 ( .A(n26120), .B(n26119), .Z(n25988) );
  NANDN U26745 ( .A(n25971), .B(n25970), .Z(n25975) );
  NANDN U26746 ( .A(n25973), .B(n25972), .Z(n25974) );
  AND U26747 ( .A(n25975), .B(n25974), .Z(n25987) );
  XOR U26748 ( .A(n25988), .B(n25987), .Z(n25990) );
  XNOR U26749 ( .A(n25989), .B(n25990), .Z(n25981) );
  XNOR U26750 ( .A(n25982), .B(n25981), .Z(n25983) );
  XNOR U26751 ( .A(n25984), .B(n25983), .Z(n26123) );
  XNOR U26752 ( .A(sreg[413]), .B(n26123), .Z(n26125) );
  NANDN U26753 ( .A(sreg[412]), .B(n25976), .Z(n25980) );
  NAND U26754 ( .A(n25978), .B(n25977), .Z(n25979) );
  NAND U26755 ( .A(n25980), .B(n25979), .Z(n26124) );
  XNOR U26756 ( .A(n26125), .B(n26124), .Z(c[413]) );
  NANDN U26757 ( .A(n25982), .B(n25981), .Z(n25986) );
  NANDN U26758 ( .A(n25984), .B(n25983), .Z(n25985) );
  AND U26759 ( .A(n25986), .B(n25985), .Z(n26131) );
  NANDN U26760 ( .A(n25988), .B(n25987), .Z(n25992) );
  NANDN U26761 ( .A(n25990), .B(n25989), .Z(n25991) );
  AND U26762 ( .A(n25992), .B(n25991), .Z(n26129) );
  NANDN U26763 ( .A(n25994), .B(n25993), .Z(n25998) );
  NANDN U26764 ( .A(n25996), .B(n25995), .Z(n25997) );
  AND U26765 ( .A(n25998), .B(n25997), .Z(n26208) );
  NAND U26766 ( .A(n38385), .B(n25999), .Z(n26001) );
  XOR U26767 ( .A(b[27]), .B(a[164]), .Z(n26152) );
  NAND U26768 ( .A(n38343), .B(n26152), .Z(n26000) );
  AND U26769 ( .A(n26001), .B(n26000), .Z(n26215) );
  NAND U26770 ( .A(n183), .B(n26002), .Z(n26004) );
  XOR U26771 ( .A(b[5]), .B(a[186]), .Z(n26155) );
  NAND U26772 ( .A(n36296), .B(n26155), .Z(n26003) );
  AND U26773 ( .A(n26004), .B(n26003), .Z(n26213) );
  NAND U26774 ( .A(n190), .B(n26005), .Z(n26007) );
  XOR U26775 ( .A(b[19]), .B(a[172]), .Z(n26158) );
  NAND U26776 ( .A(n37821), .B(n26158), .Z(n26006) );
  NAND U26777 ( .A(n26007), .B(n26006), .Z(n26212) );
  XNOR U26778 ( .A(n26213), .B(n26212), .Z(n26214) );
  XNOR U26779 ( .A(n26215), .B(n26214), .Z(n26206) );
  NAND U26780 ( .A(n38470), .B(n26008), .Z(n26010) );
  XOR U26781 ( .A(b[31]), .B(a[160]), .Z(n26161) );
  NAND U26782 ( .A(n38453), .B(n26161), .Z(n26009) );
  AND U26783 ( .A(n26010), .B(n26009), .Z(n26173) );
  NAND U26784 ( .A(n181), .B(n26011), .Z(n26013) );
  XOR U26785 ( .A(b[3]), .B(a[188]), .Z(n26164) );
  NAND U26786 ( .A(n182), .B(n26164), .Z(n26012) );
  AND U26787 ( .A(n26013), .B(n26012), .Z(n26171) );
  NAND U26788 ( .A(n189), .B(n26014), .Z(n26016) );
  XOR U26789 ( .A(b[17]), .B(a[174]), .Z(n26167) );
  NAND U26790 ( .A(n37652), .B(n26167), .Z(n26015) );
  NAND U26791 ( .A(n26016), .B(n26015), .Z(n26170) );
  XNOR U26792 ( .A(n26171), .B(n26170), .Z(n26172) );
  XOR U26793 ( .A(n26173), .B(n26172), .Z(n26207) );
  XOR U26794 ( .A(n26206), .B(n26207), .Z(n26209) );
  XOR U26795 ( .A(n26208), .B(n26209), .Z(n26255) );
  NANDN U26796 ( .A(n26018), .B(n26017), .Z(n26022) );
  NANDN U26797 ( .A(n26020), .B(n26019), .Z(n26021) );
  AND U26798 ( .A(n26022), .B(n26021), .Z(n26194) );
  NANDN U26799 ( .A(n26024), .B(n26023), .Z(n26028) );
  NANDN U26800 ( .A(n26026), .B(n26025), .Z(n26027) );
  NAND U26801 ( .A(n26028), .B(n26027), .Z(n26195) );
  XNOR U26802 ( .A(n26194), .B(n26195), .Z(n26196) );
  NANDN U26803 ( .A(n26030), .B(n26029), .Z(n26034) );
  NAND U26804 ( .A(n26032), .B(n26031), .Z(n26033) );
  NAND U26805 ( .A(n26034), .B(n26033), .Z(n26197) );
  XNOR U26806 ( .A(n26196), .B(n26197), .Z(n26254) );
  XNOR U26807 ( .A(n26255), .B(n26254), .Z(n26257) );
  NAND U26808 ( .A(n26036), .B(n26035), .Z(n26040) );
  NAND U26809 ( .A(n26038), .B(n26037), .Z(n26039) );
  AND U26810 ( .A(n26040), .B(n26039), .Z(n26256) );
  XOR U26811 ( .A(n26257), .B(n26256), .Z(n26268) );
  NANDN U26812 ( .A(n26042), .B(n26041), .Z(n26046) );
  NANDN U26813 ( .A(n26044), .B(n26043), .Z(n26045) );
  AND U26814 ( .A(n26046), .B(n26045), .Z(n26266) );
  NANDN U26815 ( .A(n26052), .B(n26051), .Z(n26056) );
  OR U26816 ( .A(n26054), .B(n26053), .Z(n26055) );
  AND U26817 ( .A(n26056), .B(n26055), .Z(n26261) );
  NANDN U26818 ( .A(n26058), .B(n26057), .Z(n26062) );
  NANDN U26819 ( .A(n26060), .B(n26059), .Z(n26061) );
  AND U26820 ( .A(n26062), .B(n26061), .Z(n26201) );
  NANDN U26821 ( .A(n26064), .B(n26063), .Z(n26068) );
  OR U26822 ( .A(n26066), .B(n26065), .Z(n26067) );
  NAND U26823 ( .A(n26068), .B(n26067), .Z(n26200) );
  XNOR U26824 ( .A(n26201), .B(n26200), .Z(n26202) );
  NAND U26825 ( .A(b[0]), .B(a[190]), .Z(n26069) );
  XNOR U26826 ( .A(b[1]), .B(n26069), .Z(n26071) );
  NANDN U26827 ( .A(b[0]), .B(a[189]), .Z(n26070) );
  NAND U26828 ( .A(n26071), .B(n26070), .Z(n26149) );
  NAND U26829 ( .A(n194), .B(n26072), .Z(n26074) );
  XOR U26830 ( .A(b[29]), .B(a[162]), .Z(n26227) );
  NAND U26831 ( .A(n38456), .B(n26227), .Z(n26073) );
  AND U26832 ( .A(n26074), .B(n26073), .Z(n26147) );
  AND U26833 ( .A(b[31]), .B(a[158]), .Z(n26146) );
  XNOR U26834 ( .A(n26147), .B(n26146), .Z(n26148) );
  XNOR U26835 ( .A(n26149), .B(n26148), .Z(n26188) );
  NAND U26836 ( .A(n38185), .B(n26075), .Z(n26077) );
  XOR U26837 ( .A(b[23]), .B(a[168]), .Z(n26230) );
  NAND U26838 ( .A(n38132), .B(n26230), .Z(n26076) );
  AND U26839 ( .A(n26077), .B(n26076), .Z(n26221) );
  NAND U26840 ( .A(n184), .B(n26078), .Z(n26080) );
  XOR U26841 ( .A(b[7]), .B(a[184]), .Z(n26233) );
  NAND U26842 ( .A(n36592), .B(n26233), .Z(n26079) );
  AND U26843 ( .A(n26080), .B(n26079), .Z(n26219) );
  NAND U26844 ( .A(n38289), .B(n26081), .Z(n26083) );
  XOR U26845 ( .A(b[25]), .B(a[166]), .Z(n26236) );
  NAND U26846 ( .A(n38247), .B(n26236), .Z(n26082) );
  NAND U26847 ( .A(n26083), .B(n26082), .Z(n26218) );
  XNOR U26848 ( .A(n26219), .B(n26218), .Z(n26220) );
  XOR U26849 ( .A(n26221), .B(n26220), .Z(n26189) );
  XNOR U26850 ( .A(n26188), .B(n26189), .Z(n26190) );
  NAND U26851 ( .A(n187), .B(n26084), .Z(n26086) );
  XOR U26852 ( .A(b[13]), .B(a[178]), .Z(n26239) );
  NAND U26853 ( .A(n37295), .B(n26239), .Z(n26085) );
  AND U26854 ( .A(n26086), .B(n26085), .Z(n26183) );
  NAND U26855 ( .A(n186), .B(n26087), .Z(n26089) );
  XOR U26856 ( .A(b[11]), .B(a[180]), .Z(n26242) );
  NAND U26857 ( .A(n37097), .B(n26242), .Z(n26088) );
  NAND U26858 ( .A(n26089), .B(n26088), .Z(n26182) );
  XNOR U26859 ( .A(n26183), .B(n26182), .Z(n26184) );
  NAND U26860 ( .A(n188), .B(n26090), .Z(n26092) );
  XOR U26861 ( .A(b[15]), .B(a[176]), .Z(n26245) );
  NAND U26862 ( .A(n37382), .B(n26245), .Z(n26091) );
  AND U26863 ( .A(n26092), .B(n26091), .Z(n26179) );
  NAND U26864 ( .A(n38064), .B(n26093), .Z(n26095) );
  XOR U26865 ( .A(b[21]), .B(a[170]), .Z(n26248) );
  NAND U26866 ( .A(n37993), .B(n26248), .Z(n26094) );
  AND U26867 ( .A(n26095), .B(n26094), .Z(n26177) );
  NAND U26868 ( .A(n185), .B(n26096), .Z(n26098) );
  XOR U26869 ( .A(b[9]), .B(a[182]), .Z(n26251) );
  NAND U26870 ( .A(n36805), .B(n26251), .Z(n26097) );
  NAND U26871 ( .A(n26098), .B(n26097), .Z(n26176) );
  XNOR U26872 ( .A(n26177), .B(n26176), .Z(n26178) );
  XOR U26873 ( .A(n26179), .B(n26178), .Z(n26185) );
  XOR U26874 ( .A(n26184), .B(n26185), .Z(n26191) );
  XOR U26875 ( .A(n26190), .B(n26191), .Z(n26203) );
  XNOR U26876 ( .A(n26202), .B(n26203), .Z(n26260) );
  XNOR U26877 ( .A(n26261), .B(n26260), .Z(n26262) );
  XOR U26878 ( .A(n26263), .B(n26262), .Z(n26267) );
  XOR U26879 ( .A(n26266), .B(n26267), .Z(n26269) );
  XOR U26880 ( .A(n26268), .B(n26269), .Z(n26143) );
  NANDN U26881 ( .A(n26100), .B(n26099), .Z(n26104) );
  NAND U26882 ( .A(n26102), .B(n26101), .Z(n26103) );
  AND U26883 ( .A(n26104), .B(n26103), .Z(n26141) );
  NANDN U26884 ( .A(n26106), .B(n26105), .Z(n26110) );
  NANDN U26885 ( .A(n26108), .B(n26107), .Z(n26109) );
  AND U26886 ( .A(n26110), .B(n26109), .Z(n26140) );
  XNOR U26887 ( .A(n26141), .B(n26140), .Z(n26142) );
  XNOR U26888 ( .A(n26143), .B(n26142), .Z(n26134) );
  NANDN U26889 ( .A(n26112), .B(n26111), .Z(n26116) );
  NANDN U26890 ( .A(n26114), .B(n26113), .Z(n26115) );
  NAND U26891 ( .A(n26116), .B(n26115), .Z(n26135) );
  XNOR U26892 ( .A(n26134), .B(n26135), .Z(n26136) );
  NANDN U26893 ( .A(n26118), .B(n26117), .Z(n26122) );
  NAND U26894 ( .A(n26120), .B(n26119), .Z(n26121) );
  NAND U26895 ( .A(n26122), .B(n26121), .Z(n26137) );
  XNOR U26896 ( .A(n26136), .B(n26137), .Z(n26128) );
  XNOR U26897 ( .A(n26129), .B(n26128), .Z(n26130) );
  XNOR U26898 ( .A(n26131), .B(n26130), .Z(n26272) );
  XNOR U26899 ( .A(sreg[414]), .B(n26272), .Z(n26274) );
  NANDN U26900 ( .A(sreg[413]), .B(n26123), .Z(n26127) );
  NAND U26901 ( .A(n26125), .B(n26124), .Z(n26126) );
  NAND U26902 ( .A(n26127), .B(n26126), .Z(n26273) );
  XNOR U26903 ( .A(n26274), .B(n26273), .Z(c[414]) );
  NANDN U26904 ( .A(n26129), .B(n26128), .Z(n26133) );
  NANDN U26905 ( .A(n26131), .B(n26130), .Z(n26132) );
  AND U26906 ( .A(n26133), .B(n26132), .Z(n26280) );
  NANDN U26907 ( .A(n26135), .B(n26134), .Z(n26139) );
  NANDN U26908 ( .A(n26137), .B(n26136), .Z(n26138) );
  AND U26909 ( .A(n26139), .B(n26138), .Z(n26278) );
  NANDN U26910 ( .A(n26141), .B(n26140), .Z(n26145) );
  NANDN U26911 ( .A(n26143), .B(n26142), .Z(n26144) );
  AND U26912 ( .A(n26145), .B(n26144), .Z(n26286) );
  NANDN U26913 ( .A(n26147), .B(n26146), .Z(n26151) );
  NANDN U26914 ( .A(n26149), .B(n26148), .Z(n26150) );
  AND U26915 ( .A(n26151), .B(n26150), .Z(n26369) );
  NAND U26916 ( .A(n38385), .B(n26152), .Z(n26154) );
  XOR U26917 ( .A(b[27]), .B(a[165]), .Z(n26313) );
  NAND U26918 ( .A(n38343), .B(n26313), .Z(n26153) );
  AND U26919 ( .A(n26154), .B(n26153), .Z(n26376) );
  NAND U26920 ( .A(n183), .B(n26155), .Z(n26157) );
  XOR U26921 ( .A(b[5]), .B(a[187]), .Z(n26316) );
  NAND U26922 ( .A(n36296), .B(n26316), .Z(n26156) );
  AND U26923 ( .A(n26157), .B(n26156), .Z(n26374) );
  NAND U26924 ( .A(n190), .B(n26158), .Z(n26160) );
  XOR U26925 ( .A(b[19]), .B(a[173]), .Z(n26319) );
  NAND U26926 ( .A(n37821), .B(n26319), .Z(n26159) );
  NAND U26927 ( .A(n26160), .B(n26159), .Z(n26373) );
  XNOR U26928 ( .A(n26374), .B(n26373), .Z(n26375) );
  XNOR U26929 ( .A(n26376), .B(n26375), .Z(n26367) );
  NAND U26930 ( .A(n38470), .B(n26161), .Z(n26163) );
  XOR U26931 ( .A(b[31]), .B(a[161]), .Z(n26322) );
  NAND U26932 ( .A(n38453), .B(n26322), .Z(n26162) );
  AND U26933 ( .A(n26163), .B(n26162), .Z(n26334) );
  NAND U26934 ( .A(n181), .B(n26164), .Z(n26166) );
  XOR U26935 ( .A(b[3]), .B(a[189]), .Z(n26325) );
  NAND U26936 ( .A(n182), .B(n26325), .Z(n26165) );
  AND U26937 ( .A(n26166), .B(n26165), .Z(n26332) );
  NAND U26938 ( .A(n189), .B(n26167), .Z(n26169) );
  XOR U26939 ( .A(b[17]), .B(a[175]), .Z(n26328) );
  NAND U26940 ( .A(n37652), .B(n26328), .Z(n26168) );
  NAND U26941 ( .A(n26169), .B(n26168), .Z(n26331) );
  XNOR U26942 ( .A(n26332), .B(n26331), .Z(n26333) );
  XOR U26943 ( .A(n26334), .B(n26333), .Z(n26368) );
  XOR U26944 ( .A(n26367), .B(n26368), .Z(n26370) );
  XOR U26945 ( .A(n26369), .B(n26370), .Z(n26302) );
  NANDN U26946 ( .A(n26171), .B(n26170), .Z(n26175) );
  NANDN U26947 ( .A(n26173), .B(n26172), .Z(n26174) );
  AND U26948 ( .A(n26175), .B(n26174), .Z(n26355) );
  NANDN U26949 ( .A(n26177), .B(n26176), .Z(n26181) );
  NANDN U26950 ( .A(n26179), .B(n26178), .Z(n26180) );
  NAND U26951 ( .A(n26181), .B(n26180), .Z(n26356) );
  XNOR U26952 ( .A(n26355), .B(n26356), .Z(n26357) );
  NANDN U26953 ( .A(n26183), .B(n26182), .Z(n26187) );
  NANDN U26954 ( .A(n26185), .B(n26184), .Z(n26186) );
  NAND U26955 ( .A(n26187), .B(n26186), .Z(n26358) );
  XNOR U26956 ( .A(n26357), .B(n26358), .Z(n26301) );
  XNOR U26957 ( .A(n26302), .B(n26301), .Z(n26304) );
  NANDN U26958 ( .A(n26189), .B(n26188), .Z(n26193) );
  NANDN U26959 ( .A(n26191), .B(n26190), .Z(n26192) );
  AND U26960 ( .A(n26193), .B(n26192), .Z(n26303) );
  XOR U26961 ( .A(n26304), .B(n26303), .Z(n26417) );
  NANDN U26962 ( .A(n26195), .B(n26194), .Z(n26199) );
  NANDN U26963 ( .A(n26197), .B(n26196), .Z(n26198) );
  AND U26964 ( .A(n26199), .B(n26198), .Z(n26415) );
  NANDN U26965 ( .A(n26201), .B(n26200), .Z(n26205) );
  NANDN U26966 ( .A(n26203), .B(n26202), .Z(n26204) );
  AND U26967 ( .A(n26205), .B(n26204), .Z(n26298) );
  NANDN U26968 ( .A(n26207), .B(n26206), .Z(n26211) );
  OR U26969 ( .A(n26209), .B(n26208), .Z(n26210) );
  AND U26970 ( .A(n26211), .B(n26210), .Z(n26296) );
  NANDN U26971 ( .A(n26213), .B(n26212), .Z(n26217) );
  NANDN U26972 ( .A(n26215), .B(n26214), .Z(n26216) );
  AND U26973 ( .A(n26217), .B(n26216), .Z(n26362) );
  NANDN U26974 ( .A(n26219), .B(n26218), .Z(n26223) );
  NANDN U26975 ( .A(n26221), .B(n26220), .Z(n26222) );
  NAND U26976 ( .A(n26223), .B(n26222), .Z(n26361) );
  XNOR U26977 ( .A(n26362), .B(n26361), .Z(n26363) );
  NAND U26978 ( .A(b[0]), .B(a[191]), .Z(n26224) );
  XNOR U26979 ( .A(b[1]), .B(n26224), .Z(n26226) );
  NANDN U26980 ( .A(b[0]), .B(a[190]), .Z(n26225) );
  NAND U26981 ( .A(n26226), .B(n26225), .Z(n26310) );
  NAND U26982 ( .A(n194), .B(n26227), .Z(n26229) );
  XOR U26983 ( .A(b[29]), .B(a[163]), .Z(n26388) );
  NAND U26984 ( .A(n38456), .B(n26388), .Z(n26228) );
  AND U26985 ( .A(n26229), .B(n26228), .Z(n26308) );
  AND U26986 ( .A(b[31]), .B(a[159]), .Z(n26307) );
  XNOR U26987 ( .A(n26308), .B(n26307), .Z(n26309) );
  XNOR U26988 ( .A(n26310), .B(n26309), .Z(n26349) );
  NAND U26989 ( .A(n38185), .B(n26230), .Z(n26232) );
  XOR U26990 ( .A(b[23]), .B(a[169]), .Z(n26391) );
  NAND U26991 ( .A(n38132), .B(n26391), .Z(n26231) );
  AND U26992 ( .A(n26232), .B(n26231), .Z(n26382) );
  NAND U26993 ( .A(n184), .B(n26233), .Z(n26235) );
  XOR U26994 ( .A(b[7]), .B(a[185]), .Z(n26394) );
  NAND U26995 ( .A(n36592), .B(n26394), .Z(n26234) );
  AND U26996 ( .A(n26235), .B(n26234), .Z(n26380) );
  NAND U26997 ( .A(n38289), .B(n26236), .Z(n26238) );
  XOR U26998 ( .A(b[25]), .B(a[167]), .Z(n26397) );
  NAND U26999 ( .A(n38247), .B(n26397), .Z(n26237) );
  NAND U27000 ( .A(n26238), .B(n26237), .Z(n26379) );
  XNOR U27001 ( .A(n26380), .B(n26379), .Z(n26381) );
  XOR U27002 ( .A(n26382), .B(n26381), .Z(n26350) );
  XNOR U27003 ( .A(n26349), .B(n26350), .Z(n26351) );
  NAND U27004 ( .A(n187), .B(n26239), .Z(n26241) );
  XOR U27005 ( .A(b[13]), .B(a[179]), .Z(n26400) );
  NAND U27006 ( .A(n37295), .B(n26400), .Z(n26240) );
  AND U27007 ( .A(n26241), .B(n26240), .Z(n26344) );
  NAND U27008 ( .A(n186), .B(n26242), .Z(n26244) );
  XOR U27009 ( .A(b[11]), .B(a[181]), .Z(n26403) );
  NAND U27010 ( .A(n37097), .B(n26403), .Z(n26243) );
  NAND U27011 ( .A(n26244), .B(n26243), .Z(n26343) );
  XNOR U27012 ( .A(n26344), .B(n26343), .Z(n26345) );
  NAND U27013 ( .A(n188), .B(n26245), .Z(n26247) );
  XOR U27014 ( .A(b[15]), .B(a[177]), .Z(n26406) );
  NAND U27015 ( .A(n37382), .B(n26406), .Z(n26246) );
  AND U27016 ( .A(n26247), .B(n26246), .Z(n26340) );
  NAND U27017 ( .A(n38064), .B(n26248), .Z(n26250) );
  XOR U27018 ( .A(b[21]), .B(a[171]), .Z(n26409) );
  NAND U27019 ( .A(n37993), .B(n26409), .Z(n26249) );
  AND U27020 ( .A(n26250), .B(n26249), .Z(n26338) );
  NAND U27021 ( .A(n185), .B(n26251), .Z(n26253) );
  XOR U27022 ( .A(b[9]), .B(a[183]), .Z(n26412) );
  NAND U27023 ( .A(n36805), .B(n26412), .Z(n26252) );
  NAND U27024 ( .A(n26253), .B(n26252), .Z(n26337) );
  XNOR U27025 ( .A(n26338), .B(n26337), .Z(n26339) );
  XOR U27026 ( .A(n26340), .B(n26339), .Z(n26346) );
  XOR U27027 ( .A(n26345), .B(n26346), .Z(n26352) );
  XOR U27028 ( .A(n26351), .B(n26352), .Z(n26364) );
  XNOR U27029 ( .A(n26363), .B(n26364), .Z(n26295) );
  XNOR U27030 ( .A(n26296), .B(n26295), .Z(n26297) );
  XOR U27031 ( .A(n26298), .B(n26297), .Z(n26416) );
  XOR U27032 ( .A(n26415), .B(n26416), .Z(n26418) );
  XOR U27033 ( .A(n26417), .B(n26418), .Z(n26292) );
  NANDN U27034 ( .A(n26255), .B(n26254), .Z(n26259) );
  NAND U27035 ( .A(n26257), .B(n26256), .Z(n26258) );
  AND U27036 ( .A(n26259), .B(n26258), .Z(n26290) );
  NANDN U27037 ( .A(n26261), .B(n26260), .Z(n26265) );
  NANDN U27038 ( .A(n26263), .B(n26262), .Z(n26264) );
  AND U27039 ( .A(n26265), .B(n26264), .Z(n26289) );
  XNOR U27040 ( .A(n26290), .B(n26289), .Z(n26291) );
  XNOR U27041 ( .A(n26292), .B(n26291), .Z(n26283) );
  NANDN U27042 ( .A(n26267), .B(n26266), .Z(n26271) );
  OR U27043 ( .A(n26269), .B(n26268), .Z(n26270) );
  NAND U27044 ( .A(n26271), .B(n26270), .Z(n26284) );
  XNOR U27045 ( .A(n26283), .B(n26284), .Z(n26285) );
  XNOR U27046 ( .A(n26286), .B(n26285), .Z(n26277) );
  XNOR U27047 ( .A(n26278), .B(n26277), .Z(n26279) );
  XNOR U27048 ( .A(n26280), .B(n26279), .Z(n26421) );
  XNOR U27049 ( .A(sreg[415]), .B(n26421), .Z(n26423) );
  NANDN U27050 ( .A(sreg[414]), .B(n26272), .Z(n26276) );
  NAND U27051 ( .A(n26274), .B(n26273), .Z(n26275) );
  NAND U27052 ( .A(n26276), .B(n26275), .Z(n26422) );
  XNOR U27053 ( .A(n26423), .B(n26422), .Z(c[415]) );
  NANDN U27054 ( .A(n26278), .B(n26277), .Z(n26282) );
  NANDN U27055 ( .A(n26280), .B(n26279), .Z(n26281) );
  AND U27056 ( .A(n26282), .B(n26281), .Z(n26429) );
  NANDN U27057 ( .A(n26284), .B(n26283), .Z(n26288) );
  NANDN U27058 ( .A(n26286), .B(n26285), .Z(n26287) );
  AND U27059 ( .A(n26288), .B(n26287), .Z(n26427) );
  NANDN U27060 ( .A(n26290), .B(n26289), .Z(n26294) );
  NANDN U27061 ( .A(n26292), .B(n26291), .Z(n26293) );
  AND U27062 ( .A(n26294), .B(n26293), .Z(n26435) );
  NANDN U27063 ( .A(n26296), .B(n26295), .Z(n26300) );
  NANDN U27064 ( .A(n26298), .B(n26297), .Z(n26299) );
  AND U27065 ( .A(n26300), .B(n26299), .Z(n26439) );
  NANDN U27066 ( .A(n26302), .B(n26301), .Z(n26306) );
  NAND U27067 ( .A(n26304), .B(n26303), .Z(n26305) );
  AND U27068 ( .A(n26306), .B(n26305), .Z(n26438) );
  XNOR U27069 ( .A(n26439), .B(n26438), .Z(n26441) );
  NANDN U27070 ( .A(n26308), .B(n26307), .Z(n26312) );
  NANDN U27071 ( .A(n26310), .B(n26309), .Z(n26311) );
  AND U27072 ( .A(n26312), .B(n26311), .Z(n26518) );
  NAND U27073 ( .A(n38385), .B(n26313), .Z(n26315) );
  XOR U27074 ( .A(b[27]), .B(a[166]), .Z(n26462) );
  NAND U27075 ( .A(n38343), .B(n26462), .Z(n26314) );
  AND U27076 ( .A(n26315), .B(n26314), .Z(n26525) );
  NAND U27077 ( .A(n183), .B(n26316), .Z(n26318) );
  XOR U27078 ( .A(b[5]), .B(a[188]), .Z(n26465) );
  NAND U27079 ( .A(n36296), .B(n26465), .Z(n26317) );
  AND U27080 ( .A(n26318), .B(n26317), .Z(n26523) );
  NAND U27081 ( .A(n190), .B(n26319), .Z(n26321) );
  XOR U27082 ( .A(b[19]), .B(a[174]), .Z(n26468) );
  NAND U27083 ( .A(n37821), .B(n26468), .Z(n26320) );
  NAND U27084 ( .A(n26321), .B(n26320), .Z(n26522) );
  XNOR U27085 ( .A(n26523), .B(n26522), .Z(n26524) );
  XNOR U27086 ( .A(n26525), .B(n26524), .Z(n26516) );
  NAND U27087 ( .A(n38470), .B(n26322), .Z(n26324) );
  XOR U27088 ( .A(b[31]), .B(a[162]), .Z(n26471) );
  NAND U27089 ( .A(n38453), .B(n26471), .Z(n26323) );
  AND U27090 ( .A(n26324), .B(n26323), .Z(n26483) );
  NAND U27091 ( .A(n181), .B(n26325), .Z(n26327) );
  XOR U27092 ( .A(b[3]), .B(a[190]), .Z(n26474) );
  NAND U27093 ( .A(n182), .B(n26474), .Z(n26326) );
  AND U27094 ( .A(n26327), .B(n26326), .Z(n26481) );
  NAND U27095 ( .A(n189), .B(n26328), .Z(n26330) );
  XOR U27096 ( .A(b[17]), .B(a[176]), .Z(n26477) );
  NAND U27097 ( .A(n37652), .B(n26477), .Z(n26329) );
  NAND U27098 ( .A(n26330), .B(n26329), .Z(n26480) );
  XNOR U27099 ( .A(n26481), .B(n26480), .Z(n26482) );
  XOR U27100 ( .A(n26483), .B(n26482), .Z(n26517) );
  XOR U27101 ( .A(n26516), .B(n26517), .Z(n26519) );
  XOR U27102 ( .A(n26518), .B(n26519), .Z(n26451) );
  NANDN U27103 ( .A(n26332), .B(n26331), .Z(n26336) );
  NANDN U27104 ( .A(n26334), .B(n26333), .Z(n26335) );
  AND U27105 ( .A(n26336), .B(n26335), .Z(n26504) );
  NANDN U27106 ( .A(n26338), .B(n26337), .Z(n26342) );
  NANDN U27107 ( .A(n26340), .B(n26339), .Z(n26341) );
  NAND U27108 ( .A(n26342), .B(n26341), .Z(n26505) );
  XNOR U27109 ( .A(n26504), .B(n26505), .Z(n26506) );
  NANDN U27110 ( .A(n26344), .B(n26343), .Z(n26348) );
  NANDN U27111 ( .A(n26346), .B(n26345), .Z(n26347) );
  NAND U27112 ( .A(n26348), .B(n26347), .Z(n26507) );
  XNOR U27113 ( .A(n26506), .B(n26507), .Z(n26450) );
  XNOR U27114 ( .A(n26451), .B(n26450), .Z(n26453) );
  NANDN U27115 ( .A(n26350), .B(n26349), .Z(n26354) );
  NANDN U27116 ( .A(n26352), .B(n26351), .Z(n26353) );
  AND U27117 ( .A(n26354), .B(n26353), .Z(n26452) );
  XOR U27118 ( .A(n26453), .B(n26452), .Z(n26567) );
  NANDN U27119 ( .A(n26356), .B(n26355), .Z(n26360) );
  NANDN U27120 ( .A(n26358), .B(n26357), .Z(n26359) );
  AND U27121 ( .A(n26360), .B(n26359), .Z(n26564) );
  NANDN U27122 ( .A(n26362), .B(n26361), .Z(n26366) );
  NANDN U27123 ( .A(n26364), .B(n26363), .Z(n26365) );
  AND U27124 ( .A(n26366), .B(n26365), .Z(n26447) );
  NANDN U27125 ( .A(n26368), .B(n26367), .Z(n26372) );
  OR U27126 ( .A(n26370), .B(n26369), .Z(n26371) );
  AND U27127 ( .A(n26372), .B(n26371), .Z(n26445) );
  NANDN U27128 ( .A(n26374), .B(n26373), .Z(n26378) );
  NANDN U27129 ( .A(n26376), .B(n26375), .Z(n26377) );
  AND U27130 ( .A(n26378), .B(n26377), .Z(n26511) );
  NANDN U27131 ( .A(n26380), .B(n26379), .Z(n26384) );
  NANDN U27132 ( .A(n26382), .B(n26381), .Z(n26383) );
  NAND U27133 ( .A(n26384), .B(n26383), .Z(n26510) );
  XNOR U27134 ( .A(n26511), .B(n26510), .Z(n26512) );
  NAND U27135 ( .A(b[0]), .B(a[192]), .Z(n26385) );
  XNOR U27136 ( .A(b[1]), .B(n26385), .Z(n26387) );
  NANDN U27137 ( .A(b[0]), .B(a[191]), .Z(n26386) );
  NAND U27138 ( .A(n26387), .B(n26386), .Z(n26459) );
  NAND U27139 ( .A(n194), .B(n26388), .Z(n26390) );
  XOR U27140 ( .A(b[29]), .B(a[164]), .Z(n26537) );
  NAND U27141 ( .A(n38456), .B(n26537), .Z(n26389) );
  AND U27142 ( .A(n26390), .B(n26389), .Z(n26457) );
  AND U27143 ( .A(b[31]), .B(a[160]), .Z(n26456) );
  XNOR U27144 ( .A(n26457), .B(n26456), .Z(n26458) );
  XNOR U27145 ( .A(n26459), .B(n26458), .Z(n26498) );
  NAND U27146 ( .A(n38185), .B(n26391), .Z(n26393) );
  XOR U27147 ( .A(b[23]), .B(a[170]), .Z(n26540) );
  NAND U27148 ( .A(n38132), .B(n26540), .Z(n26392) );
  AND U27149 ( .A(n26393), .B(n26392), .Z(n26531) );
  NAND U27150 ( .A(n184), .B(n26394), .Z(n26396) );
  XOR U27151 ( .A(b[7]), .B(a[186]), .Z(n26543) );
  NAND U27152 ( .A(n36592), .B(n26543), .Z(n26395) );
  AND U27153 ( .A(n26396), .B(n26395), .Z(n26529) );
  NAND U27154 ( .A(n38289), .B(n26397), .Z(n26399) );
  XOR U27155 ( .A(b[25]), .B(a[168]), .Z(n26546) );
  NAND U27156 ( .A(n38247), .B(n26546), .Z(n26398) );
  NAND U27157 ( .A(n26399), .B(n26398), .Z(n26528) );
  XNOR U27158 ( .A(n26529), .B(n26528), .Z(n26530) );
  XOR U27159 ( .A(n26531), .B(n26530), .Z(n26499) );
  XNOR U27160 ( .A(n26498), .B(n26499), .Z(n26500) );
  NAND U27161 ( .A(n187), .B(n26400), .Z(n26402) );
  XOR U27162 ( .A(b[13]), .B(a[180]), .Z(n26549) );
  NAND U27163 ( .A(n37295), .B(n26549), .Z(n26401) );
  AND U27164 ( .A(n26402), .B(n26401), .Z(n26493) );
  NAND U27165 ( .A(n186), .B(n26403), .Z(n26405) );
  XOR U27166 ( .A(b[11]), .B(a[182]), .Z(n26552) );
  NAND U27167 ( .A(n37097), .B(n26552), .Z(n26404) );
  NAND U27168 ( .A(n26405), .B(n26404), .Z(n26492) );
  XNOR U27169 ( .A(n26493), .B(n26492), .Z(n26494) );
  NAND U27170 ( .A(n188), .B(n26406), .Z(n26408) );
  XOR U27171 ( .A(b[15]), .B(a[178]), .Z(n26555) );
  NAND U27172 ( .A(n37382), .B(n26555), .Z(n26407) );
  AND U27173 ( .A(n26408), .B(n26407), .Z(n26489) );
  NAND U27174 ( .A(n38064), .B(n26409), .Z(n26411) );
  XOR U27175 ( .A(b[21]), .B(a[172]), .Z(n26558) );
  NAND U27176 ( .A(n37993), .B(n26558), .Z(n26410) );
  AND U27177 ( .A(n26411), .B(n26410), .Z(n26487) );
  NAND U27178 ( .A(n185), .B(n26412), .Z(n26414) );
  XOR U27179 ( .A(b[9]), .B(a[184]), .Z(n26561) );
  NAND U27180 ( .A(n36805), .B(n26561), .Z(n26413) );
  NAND U27181 ( .A(n26414), .B(n26413), .Z(n26486) );
  XNOR U27182 ( .A(n26487), .B(n26486), .Z(n26488) );
  XOR U27183 ( .A(n26489), .B(n26488), .Z(n26495) );
  XOR U27184 ( .A(n26494), .B(n26495), .Z(n26501) );
  XOR U27185 ( .A(n26500), .B(n26501), .Z(n26513) );
  XNOR U27186 ( .A(n26512), .B(n26513), .Z(n26444) );
  XNOR U27187 ( .A(n26445), .B(n26444), .Z(n26446) );
  XOR U27188 ( .A(n26447), .B(n26446), .Z(n26565) );
  XNOR U27189 ( .A(n26564), .B(n26565), .Z(n26566) );
  XNOR U27190 ( .A(n26567), .B(n26566), .Z(n26440) );
  XOR U27191 ( .A(n26441), .B(n26440), .Z(n26433) );
  NANDN U27192 ( .A(n26416), .B(n26415), .Z(n26420) );
  OR U27193 ( .A(n26418), .B(n26417), .Z(n26419) );
  AND U27194 ( .A(n26420), .B(n26419), .Z(n26432) );
  XNOR U27195 ( .A(n26433), .B(n26432), .Z(n26434) );
  XNOR U27196 ( .A(n26435), .B(n26434), .Z(n26426) );
  XNOR U27197 ( .A(n26427), .B(n26426), .Z(n26428) );
  XNOR U27198 ( .A(n26429), .B(n26428), .Z(n26570) );
  XNOR U27199 ( .A(sreg[416]), .B(n26570), .Z(n26572) );
  NANDN U27200 ( .A(sreg[415]), .B(n26421), .Z(n26425) );
  NAND U27201 ( .A(n26423), .B(n26422), .Z(n26424) );
  NAND U27202 ( .A(n26425), .B(n26424), .Z(n26571) );
  XNOR U27203 ( .A(n26572), .B(n26571), .Z(c[416]) );
  NANDN U27204 ( .A(n26427), .B(n26426), .Z(n26431) );
  NANDN U27205 ( .A(n26429), .B(n26428), .Z(n26430) );
  AND U27206 ( .A(n26431), .B(n26430), .Z(n26578) );
  NANDN U27207 ( .A(n26433), .B(n26432), .Z(n26437) );
  NANDN U27208 ( .A(n26435), .B(n26434), .Z(n26436) );
  AND U27209 ( .A(n26437), .B(n26436), .Z(n26576) );
  NANDN U27210 ( .A(n26439), .B(n26438), .Z(n26443) );
  NAND U27211 ( .A(n26441), .B(n26440), .Z(n26442) );
  AND U27212 ( .A(n26443), .B(n26442), .Z(n26583) );
  NANDN U27213 ( .A(n26445), .B(n26444), .Z(n26449) );
  NANDN U27214 ( .A(n26447), .B(n26446), .Z(n26448) );
  AND U27215 ( .A(n26449), .B(n26448), .Z(n26588) );
  NANDN U27216 ( .A(n26451), .B(n26450), .Z(n26455) );
  NAND U27217 ( .A(n26453), .B(n26452), .Z(n26454) );
  AND U27218 ( .A(n26455), .B(n26454), .Z(n26587) );
  XNOR U27219 ( .A(n26588), .B(n26587), .Z(n26590) );
  NANDN U27220 ( .A(n26457), .B(n26456), .Z(n26461) );
  NANDN U27221 ( .A(n26459), .B(n26458), .Z(n26460) );
  AND U27222 ( .A(n26461), .B(n26460), .Z(n26667) );
  NAND U27223 ( .A(n38385), .B(n26462), .Z(n26464) );
  XOR U27224 ( .A(b[27]), .B(a[167]), .Z(n26611) );
  NAND U27225 ( .A(n38343), .B(n26611), .Z(n26463) );
  AND U27226 ( .A(n26464), .B(n26463), .Z(n26674) );
  NAND U27227 ( .A(n183), .B(n26465), .Z(n26467) );
  XOR U27228 ( .A(b[5]), .B(a[189]), .Z(n26614) );
  NAND U27229 ( .A(n36296), .B(n26614), .Z(n26466) );
  AND U27230 ( .A(n26467), .B(n26466), .Z(n26672) );
  NAND U27231 ( .A(n190), .B(n26468), .Z(n26470) );
  XOR U27232 ( .A(b[19]), .B(a[175]), .Z(n26617) );
  NAND U27233 ( .A(n37821), .B(n26617), .Z(n26469) );
  NAND U27234 ( .A(n26470), .B(n26469), .Z(n26671) );
  XNOR U27235 ( .A(n26672), .B(n26671), .Z(n26673) );
  XNOR U27236 ( .A(n26674), .B(n26673), .Z(n26665) );
  NAND U27237 ( .A(n38470), .B(n26471), .Z(n26473) );
  XOR U27238 ( .A(b[31]), .B(a[163]), .Z(n26620) );
  NAND U27239 ( .A(n38453), .B(n26620), .Z(n26472) );
  AND U27240 ( .A(n26473), .B(n26472), .Z(n26632) );
  NAND U27241 ( .A(n181), .B(n26474), .Z(n26476) );
  XOR U27242 ( .A(b[3]), .B(a[191]), .Z(n26623) );
  NAND U27243 ( .A(n182), .B(n26623), .Z(n26475) );
  AND U27244 ( .A(n26476), .B(n26475), .Z(n26630) );
  NAND U27245 ( .A(n189), .B(n26477), .Z(n26479) );
  XOR U27246 ( .A(b[17]), .B(a[177]), .Z(n26626) );
  NAND U27247 ( .A(n37652), .B(n26626), .Z(n26478) );
  NAND U27248 ( .A(n26479), .B(n26478), .Z(n26629) );
  XNOR U27249 ( .A(n26630), .B(n26629), .Z(n26631) );
  XOR U27250 ( .A(n26632), .B(n26631), .Z(n26666) );
  XOR U27251 ( .A(n26665), .B(n26666), .Z(n26668) );
  XOR U27252 ( .A(n26667), .B(n26668), .Z(n26600) );
  NANDN U27253 ( .A(n26481), .B(n26480), .Z(n26485) );
  NANDN U27254 ( .A(n26483), .B(n26482), .Z(n26484) );
  AND U27255 ( .A(n26485), .B(n26484), .Z(n26653) );
  NANDN U27256 ( .A(n26487), .B(n26486), .Z(n26491) );
  NANDN U27257 ( .A(n26489), .B(n26488), .Z(n26490) );
  NAND U27258 ( .A(n26491), .B(n26490), .Z(n26654) );
  XNOR U27259 ( .A(n26653), .B(n26654), .Z(n26655) );
  NANDN U27260 ( .A(n26493), .B(n26492), .Z(n26497) );
  NANDN U27261 ( .A(n26495), .B(n26494), .Z(n26496) );
  NAND U27262 ( .A(n26497), .B(n26496), .Z(n26656) );
  XNOR U27263 ( .A(n26655), .B(n26656), .Z(n26599) );
  XNOR U27264 ( .A(n26600), .B(n26599), .Z(n26602) );
  NANDN U27265 ( .A(n26499), .B(n26498), .Z(n26503) );
  NANDN U27266 ( .A(n26501), .B(n26500), .Z(n26502) );
  AND U27267 ( .A(n26503), .B(n26502), .Z(n26601) );
  XOR U27268 ( .A(n26602), .B(n26601), .Z(n26716) );
  NANDN U27269 ( .A(n26505), .B(n26504), .Z(n26509) );
  NANDN U27270 ( .A(n26507), .B(n26506), .Z(n26508) );
  AND U27271 ( .A(n26509), .B(n26508), .Z(n26713) );
  NANDN U27272 ( .A(n26511), .B(n26510), .Z(n26515) );
  NANDN U27273 ( .A(n26513), .B(n26512), .Z(n26514) );
  AND U27274 ( .A(n26515), .B(n26514), .Z(n26596) );
  NANDN U27275 ( .A(n26517), .B(n26516), .Z(n26521) );
  OR U27276 ( .A(n26519), .B(n26518), .Z(n26520) );
  AND U27277 ( .A(n26521), .B(n26520), .Z(n26594) );
  NANDN U27278 ( .A(n26523), .B(n26522), .Z(n26527) );
  NANDN U27279 ( .A(n26525), .B(n26524), .Z(n26526) );
  AND U27280 ( .A(n26527), .B(n26526), .Z(n26660) );
  NANDN U27281 ( .A(n26529), .B(n26528), .Z(n26533) );
  NANDN U27282 ( .A(n26531), .B(n26530), .Z(n26532) );
  NAND U27283 ( .A(n26533), .B(n26532), .Z(n26659) );
  XNOR U27284 ( .A(n26660), .B(n26659), .Z(n26661) );
  NAND U27285 ( .A(b[0]), .B(a[193]), .Z(n26534) );
  XNOR U27286 ( .A(b[1]), .B(n26534), .Z(n26536) );
  NANDN U27287 ( .A(b[0]), .B(a[192]), .Z(n26535) );
  NAND U27288 ( .A(n26536), .B(n26535), .Z(n26608) );
  NAND U27289 ( .A(n194), .B(n26537), .Z(n26539) );
  XOR U27290 ( .A(b[29]), .B(a[165]), .Z(n26686) );
  NAND U27291 ( .A(n38456), .B(n26686), .Z(n26538) );
  AND U27292 ( .A(n26539), .B(n26538), .Z(n26606) );
  AND U27293 ( .A(b[31]), .B(a[161]), .Z(n26605) );
  XNOR U27294 ( .A(n26606), .B(n26605), .Z(n26607) );
  XNOR U27295 ( .A(n26608), .B(n26607), .Z(n26647) );
  NAND U27296 ( .A(n38185), .B(n26540), .Z(n26542) );
  XOR U27297 ( .A(b[23]), .B(a[171]), .Z(n26689) );
  NAND U27298 ( .A(n38132), .B(n26689), .Z(n26541) );
  AND U27299 ( .A(n26542), .B(n26541), .Z(n26680) );
  NAND U27300 ( .A(n184), .B(n26543), .Z(n26545) );
  XOR U27301 ( .A(b[7]), .B(a[187]), .Z(n26692) );
  NAND U27302 ( .A(n36592), .B(n26692), .Z(n26544) );
  AND U27303 ( .A(n26545), .B(n26544), .Z(n26678) );
  NAND U27304 ( .A(n38289), .B(n26546), .Z(n26548) );
  XOR U27305 ( .A(b[25]), .B(a[169]), .Z(n26695) );
  NAND U27306 ( .A(n38247), .B(n26695), .Z(n26547) );
  NAND U27307 ( .A(n26548), .B(n26547), .Z(n26677) );
  XNOR U27308 ( .A(n26678), .B(n26677), .Z(n26679) );
  XOR U27309 ( .A(n26680), .B(n26679), .Z(n26648) );
  XNOR U27310 ( .A(n26647), .B(n26648), .Z(n26649) );
  NAND U27311 ( .A(n187), .B(n26549), .Z(n26551) );
  XOR U27312 ( .A(b[13]), .B(a[181]), .Z(n26698) );
  NAND U27313 ( .A(n37295), .B(n26698), .Z(n26550) );
  AND U27314 ( .A(n26551), .B(n26550), .Z(n26642) );
  NAND U27315 ( .A(n186), .B(n26552), .Z(n26554) );
  XOR U27316 ( .A(b[11]), .B(a[183]), .Z(n26701) );
  NAND U27317 ( .A(n37097), .B(n26701), .Z(n26553) );
  NAND U27318 ( .A(n26554), .B(n26553), .Z(n26641) );
  XNOR U27319 ( .A(n26642), .B(n26641), .Z(n26643) );
  NAND U27320 ( .A(n188), .B(n26555), .Z(n26557) );
  XOR U27321 ( .A(b[15]), .B(a[179]), .Z(n26704) );
  NAND U27322 ( .A(n37382), .B(n26704), .Z(n26556) );
  AND U27323 ( .A(n26557), .B(n26556), .Z(n26638) );
  NAND U27324 ( .A(n38064), .B(n26558), .Z(n26560) );
  XOR U27325 ( .A(b[21]), .B(a[173]), .Z(n26707) );
  NAND U27326 ( .A(n37993), .B(n26707), .Z(n26559) );
  AND U27327 ( .A(n26560), .B(n26559), .Z(n26636) );
  NAND U27328 ( .A(n185), .B(n26561), .Z(n26563) );
  XOR U27329 ( .A(b[9]), .B(a[185]), .Z(n26710) );
  NAND U27330 ( .A(n36805), .B(n26710), .Z(n26562) );
  NAND U27331 ( .A(n26563), .B(n26562), .Z(n26635) );
  XNOR U27332 ( .A(n26636), .B(n26635), .Z(n26637) );
  XOR U27333 ( .A(n26638), .B(n26637), .Z(n26644) );
  XOR U27334 ( .A(n26643), .B(n26644), .Z(n26650) );
  XOR U27335 ( .A(n26649), .B(n26650), .Z(n26662) );
  XNOR U27336 ( .A(n26661), .B(n26662), .Z(n26593) );
  XNOR U27337 ( .A(n26594), .B(n26593), .Z(n26595) );
  XOR U27338 ( .A(n26596), .B(n26595), .Z(n26714) );
  XNOR U27339 ( .A(n26713), .B(n26714), .Z(n26715) );
  XNOR U27340 ( .A(n26716), .B(n26715), .Z(n26589) );
  XOR U27341 ( .A(n26590), .B(n26589), .Z(n26582) );
  NANDN U27342 ( .A(n26565), .B(n26564), .Z(n26569) );
  NANDN U27343 ( .A(n26567), .B(n26566), .Z(n26568) );
  AND U27344 ( .A(n26569), .B(n26568), .Z(n26581) );
  XOR U27345 ( .A(n26582), .B(n26581), .Z(n26584) );
  XNOR U27346 ( .A(n26583), .B(n26584), .Z(n26575) );
  XNOR U27347 ( .A(n26576), .B(n26575), .Z(n26577) );
  XNOR U27348 ( .A(n26578), .B(n26577), .Z(n26719) );
  XNOR U27349 ( .A(sreg[417]), .B(n26719), .Z(n26721) );
  NANDN U27350 ( .A(sreg[416]), .B(n26570), .Z(n26574) );
  NAND U27351 ( .A(n26572), .B(n26571), .Z(n26573) );
  NAND U27352 ( .A(n26574), .B(n26573), .Z(n26720) );
  XNOR U27353 ( .A(n26721), .B(n26720), .Z(c[417]) );
  NANDN U27354 ( .A(n26576), .B(n26575), .Z(n26580) );
  NANDN U27355 ( .A(n26578), .B(n26577), .Z(n26579) );
  AND U27356 ( .A(n26580), .B(n26579), .Z(n26727) );
  NANDN U27357 ( .A(n26582), .B(n26581), .Z(n26586) );
  NANDN U27358 ( .A(n26584), .B(n26583), .Z(n26585) );
  AND U27359 ( .A(n26586), .B(n26585), .Z(n26725) );
  NANDN U27360 ( .A(n26588), .B(n26587), .Z(n26592) );
  NAND U27361 ( .A(n26590), .B(n26589), .Z(n26591) );
  AND U27362 ( .A(n26592), .B(n26591), .Z(n26732) );
  NANDN U27363 ( .A(n26594), .B(n26593), .Z(n26598) );
  NANDN U27364 ( .A(n26596), .B(n26595), .Z(n26597) );
  AND U27365 ( .A(n26598), .B(n26597), .Z(n26737) );
  NANDN U27366 ( .A(n26600), .B(n26599), .Z(n26604) );
  NAND U27367 ( .A(n26602), .B(n26601), .Z(n26603) );
  AND U27368 ( .A(n26604), .B(n26603), .Z(n26736) );
  XNOR U27369 ( .A(n26737), .B(n26736), .Z(n26739) );
  NANDN U27370 ( .A(n26606), .B(n26605), .Z(n26610) );
  NANDN U27371 ( .A(n26608), .B(n26607), .Z(n26609) );
  AND U27372 ( .A(n26610), .B(n26609), .Z(n26816) );
  NAND U27373 ( .A(n38385), .B(n26611), .Z(n26613) );
  XOR U27374 ( .A(b[27]), .B(a[168]), .Z(n26760) );
  NAND U27375 ( .A(n38343), .B(n26760), .Z(n26612) );
  AND U27376 ( .A(n26613), .B(n26612), .Z(n26823) );
  NAND U27377 ( .A(n183), .B(n26614), .Z(n26616) );
  XOR U27378 ( .A(b[5]), .B(a[190]), .Z(n26763) );
  NAND U27379 ( .A(n36296), .B(n26763), .Z(n26615) );
  AND U27380 ( .A(n26616), .B(n26615), .Z(n26821) );
  NAND U27381 ( .A(n190), .B(n26617), .Z(n26619) );
  XOR U27382 ( .A(b[19]), .B(a[176]), .Z(n26766) );
  NAND U27383 ( .A(n37821), .B(n26766), .Z(n26618) );
  NAND U27384 ( .A(n26619), .B(n26618), .Z(n26820) );
  XNOR U27385 ( .A(n26821), .B(n26820), .Z(n26822) );
  XNOR U27386 ( .A(n26823), .B(n26822), .Z(n26814) );
  NAND U27387 ( .A(n38470), .B(n26620), .Z(n26622) );
  XOR U27388 ( .A(b[31]), .B(a[164]), .Z(n26769) );
  NAND U27389 ( .A(n38453), .B(n26769), .Z(n26621) );
  AND U27390 ( .A(n26622), .B(n26621), .Z(n26781) );
  NAND U27391 ( .A(n181), .B(n26623), .Z(n26625) );
  XOR U27392 ( .A(b[3]), .B(a[192]), .Z(n26772) );
  NAND U27393 ( .A(n182), .B(n26772), .Z(n26624) );
  AND U27394 ( .A(n26625), .B(n26624), .Z(n26779) );
  NAND U27395 ( .A(n189), .B(n26626), .Z(n26628) );
  XOR U27396 ( .A(b[17]), .B(a[178]), .Z(n26775) );
  NAND U27397 ( .A(n37652), .B(n26775), .Z(n26627) );
  NAND U27398 ( .A(n26628), .B(n26627), .Z(n26778) );
  XNOR U27399 ( .A(n26779), .B(n26778), .Z(n26780) );
  XOR U27400 ( .A(n26781), .B(n26780), .Z(n26815) );
  XOR U27401 ( .A(n26814), .B(n26815), .Z(n26817) );
  XOR U27402 ( .A(n26816), .B(n26817), .Z(n26749) );
  NANDN U27403 ( .A(n26630), .B(n26629), .Z(n26634) );
  NANDN U27404 ( .A(n26632), .B(n26631), .Z(n26633) );
  AND U27405 ( .A(n26634), .B(n26633), .Z(n26802) );
  NANDN U27406 ( .A(n26636), .B(n26635), .Z(n26640) );
  NANDN U27407 ( .A(n26638), .B(n26637), .Z(n26639) );
  NAND U27408 ( .A(n26640), .B(n26639), .Z(n26803) );
  XNOR U27409 ( .A(n26802), .B(n26803), .Z(n26804) );
  NANDN U27410 ( .A(n26642), .B(n26641), .Z(n26646) );
  NANDN U27411 ( .A(n26644), .B(n26643), .Z(n26645) );
  NAND U27412 ( .A(n26646), .B(n26645), .Z(n26805) );
  XNOR U27413 ( .A(n26804), .B(n26805), .Z(n26748) );
  XNOR U27414 ( .A(n26749), .B(n26748), .Z(n26751) );
  NANDN U27415 ( .A(n26648), .B(n26647), .Z(n26652) );
  NANDN U27416 ( .A(n26650), .B(n26649), .Z(n26651) );
  AND U27417 ( .A(n26652), .B(n26651), .Z(n26750) );
  XOR U27418 ( .A(n26751), .B(n26750), .Z(n26865) );
  NANDN U27419 ( .A(n26654), .B(n26653), .Z(n26658) );
  NANDN U27420 ( .A(n26656), .B(n26655), .Z(n26657) );
  AND U27421 ( .A(n26658), .B(n26657), .Z(n26862) );
  NANDN U27422 ( .A(n26660), .B(n26659), .Z(n26664) );
  NANDN U27423 ( .A(n26662), .B(n26661), .Z(n26663) );
  AND U27424 ( .A(n26664), .B(n26663), .Z(n26745) );
  NANDN U27425 ( .A(n26666), .B(n26665), .Z(n26670) );
  OR U27426 ( .A(n26668), .B(n26667), .Z(n26669) );
  AND U27427 ( .A(n26670), .B(n26669), .Z(n26743) );
  NANDN U27428 ( .A(n26672), .B(n26671), .Z(n26676) );
  NANDN U27429 ( .A(n26674), .B(n26673), .Z(n26675) );
  AND U27430 ( .A(n26676), .B(n26675), .Z(n26809) );
  NANDN U27431 ( .A(n26678), .B(n26677), .Z(n26682) );
  NANDN U27432 ( .A(n26680), .B(n26679), .Z(n26681) );
  NAND U27433 ( .A(n26682), .B(n26681), .Z(n26808) );
  XNOR U27434 ( .A(n26809), .B(n26808), .Z(n26810) );
  NAND U27435 ( .A(b[0]), .B(a[194]), .Z(n26683) );
  XNOR U27436 ( .A(b[1]), .B(n26683), .Z(n26685) );
  NANDN U27437 ( .A(b[0]), .B(a[193]), .Z(n26684) );
  NAND U27438 ( .A(n26685), .B(n26684), .Z(n26757) );
  NAND U27439 ( .A(n194), .B(n26686), .Z(n26688) );
  XOR U27440 ( .A(b[29]), .B(a[166]), .Z(n26835) );
  NAND U27441 ( .A(n38456), .B(n26835), .Z(n26687) );
  AND U27442 ( .A(n26688), .B(n26687), .Z(n26755) );
  AND U27443 ( .A(b[31]), .B(a[162]), .Z(n26754) );
  XNOR U27444 ( .A(n26755), .B(n26754), .Z(n26756) );
  XNOR U27445 ( .A(n26757), .B(n26756), .Z(n26796) );
  NAND U27446 ( .A(n38185), .B(n26689), .Z(n26691) );
  XOR U27447 ( .A(b[23]), .B(a[172]), .Z(n26838) );
  NAND U27448 ( .A(n38132), .B(n26838), .Z(n26690) );
  AND U27449 ( .A(n26691), .B(n26690), .Z(n26829) );
  NAND U27450 ( .A(n184), .B(n26692), .Z(n26694) );
  XOR U27451 ( .A(b[7]), .B(a[188]), .Z(n26841) );
  NAND U27452 ( .A(n36592), .B(n26841), .Z(n26693) );
  AND U27453 ( .A(n26694), .B(n26693), .Z(n26827) );
  NAND U27454 ( .A(n38289), .B(n26695), .Z(n26697) );
  XOR U27455 ( .A(b[25]), .B(a[170]), .Z(n26844) );
  NAND U27456 ( .A(n38247), .B(n26844), .Z(n26696) );
  NAND U27457 ( .A(n26697), .B(n26696), .Z(n26826) );
  XNOR U27458 ( .A(n26827), .B(n26826), .Z(n26828) );
  XOR U27459 ( .A(n26829), .B(n26828), .Z(n26797) );
  XNOR U27460 ( .A(n26796), .B(n26797), .Z(n26798) );
  NAND U27461 ( .A(n187), .B(n26698), .Z(n26700) );
  XOR U27462 ( .A(b[13]), .B(a[182]), .Z(n26847) );
  NAND U27463 ( .A(n37295), .B(n26847), .Z(n26699) );
  AND U27464 ( .A(n26700), .B(n26699), .Z(n26791) );
  NAND U27465 ( .A(n186), .B(n26701), .Z(n26703) );
  XOR U27466 ( .A(b[11]), .B(a[184]), .Z(n26850) );
  NAND U27467 ( .A(n37097), .B(n26850), .Z(n26702) );
  NAND U27468 ( .A(n26703), .B(n26702), .Z(n26790) );
  XNOR U27469 ( .A(n26791), .B(n26790), .Z(n26792) );
  NAND U27470 ( .A(n188), .B(n26704), .Z(n26706) );
  XOR U27471 ( .A(b[15]), .B(a[180]), .Z(n26853) );
  NAND U27472 ( .A(n37382), .B(n26853), .Z(n26705) );
  AND U27473 ( .A(n26706), .B(n26705), .Z(n26787) );
  NAND U27474 ( .A(n38064), .B(n26707), .Z(n26709) );
  XOR U27475 ( .A(b[21]), .B(a[174]), .Z(n26856) );
  NAND U27476 ( .A(n37993), .B(n26856), .Z(n26708) );
  AND U27477 ( .A(n26709), .B(n26708), .Z(n26785) );
  NAND U27478 ( .A(n185), .B(n26710), .Z(n26712) );
  XOR U27479 ( .A(b[9]), .B(a[186]), .Z(n26859) );
  NAND U27480 ( .A(n36805), .B(n26859), .Z(n26711) );
  NAND U27481 ( .A(n26712), .B(n26711), .Z(n26784) );
  XNOR U27482 ( .A(n26785), .B(n26784), .Z(n26786) );
  XOR U27483 ( .A(n26787), .B(n26786), .Z(n26793) );
  XOR U27484 ( .A(n26792), .B(n26793), .Z(n26799) );
  XOR U27485 ( .A(n26798), .B(n26799), .Z(n26811) );
  XNOR U27486 ( .A(n26810), .B(n26811), .Z(n26742) );
  XNOR U27487 ( .A(n26743), .B(n26742), .Z(n26744) );
  XOR U27488 ( .A(n26745), .B(n26744), .Z(n26863) );
  XNOR U27489 ( .A(n26862), .B(n26863), .Z(n26864) );
  XNOR U27490 ( .A(n26865), .B(n26864), .Z(n26738) );
  XOR U27491 ( .A(n26739), .B(n26738), .Z(n26731) );
  NANDN U27492 ( .A(n26714), .B(n26713), .Z(n26718) );
  NANDN U27493 ( .A(n26716), .B(n26715), .Z(n26717) );
  AND U27494 ( .A(n26718), .B(n26717), .Z(n26730) );
  XOR U27495 ( .A(n26731), .B(n26730), .Z(n26733) );
  XNOR U27496 ( .A(n26732), .B(n26733), .Z(n26724) );
  XNOR U27497 ( .A(n26725), .B(n26724), .Z(n26726) );
  XNOR U27498 ( .A(n26727), .B(n26726), .Z(n26868) );
  XNOR U27499 ( .A(sreg[418]), .B(n26868), .Z(n26870) );
  NANDN U27500 ( .A(sreg[417]), .B(n26719), .Z(n26723) );
  NAND U27501 ( .A(n26721), .B(n26720), .Z(n26722) );
  NAND U27502 ( .A(n26723), .B(n26722), .Z(n26869) );
  XNOR U27503 ( .A(n26870), .B(n26869), .Z(c[418]) );
  NANDN U27504 ( .A(n26725), .B(n26724), .Z(n26729) );
  NANDN U27505 ( .A(n26727), .B(n26726), .Z(n26728) );
  AND U27506 ( .A(n26729), .B(n26728), .Z(n26876) );
  NANDN U27507 ( .A(n26731), .B(n26730), .Z(n26735) );
  NANDN U27508 ( .A(n26733), .B(n26732), .Z(n26734) );
  AND U27509 ( .A(n26735), .B(n26734), .Z(n26874) );
  NANDN U27510 ( .A(n26737), .B(n26736), .Z(n26741) );
  NAND U27511 ( .A(n26739), .B(n26738), .Z(n26740) );
  AND U27512 ( .A(n26741), .B(n26740), .Z(n26881) );
  NANDN U27513 ( .A(n26743), .B(n26742), .Z(n26747) );
  NANDN U27514 ( .A(n26745), .B(n26744), .Z(n26746) );
  AND U27515 ( .A(n26747), .B(n26746), .Z(n26886) );
  NANDN U27516 ( .A(n26749), .B(n26748), .Z(n26753) );
  NAND U27517 ( .A(n26751), .B(n26750), .Z(n26752) );
  AND U27518 ( .A(n26753), .B(n26752), .Z(n26885) );
  XNOR U27519 ( .A(n26886), .B(n26885), .Z(n26888) );
  NANDN U27520 ( .A(n26755), .B(n26754), .Z(n26759) );
  NANDN U27521 ( .A(n26757), .B(n26756), .Z(n26758) );
  AND U27522 ( .A(n26759), .B(n26758), .Z(n26963) );
  NAND U27523 ( .A(n38385), .B(n26760), .Z(n26762) );
  XOR U27524 ( .A(b[27]), .B(a[169]), .Z(n26909) );
  NAND U27525 ( .A(n38343), .B(n26909), .Z(n26761) );
  AND U27526 ( .A(n26762), .B(n26761), .Z(n26970) );
  NAND U27527 ( .A(n183), .B(n26763), .Z(n26765) );
  XOR U27528 ( .A(b[5]), .B(a[191]), .Z(n26912) );
  NAND U27529 ( .A(n36296), .B(n26912), .Z(n26764) );
  AND U27530 ( .A(n26765), .B(n26764), .Z(n26968) );
  NAND U27531 ( .A(n190), .B(n26766), .Z(n26768) );
  XOR U27532 ( .A(b[19]), .B(a[177]), .Z(n26915) );
  NAND U27533 ( .A(n37821), .B(n26915), .Z(n26767) );
  NAND U27534 ( .A(n26768), .B(n26767), .Z(n26967) );
  XNOR U27535 ( .A(n26968), .B(n26967), .Z(n26969) );
  XNOR U27536 ( .A(n26970), .B(n26969), .Z(n26961) );
  NAND U27537 ( .A(n38470), .B(n26769), .Z(n26771) );
  XOR U27538 ( .A(b[31]), .B(a[165]), .Z(n26918) );
  NAND U27539 ( .A(n38453), .B(n26918), .Z(n26770) );
  AND U27540 ( .A(n26771), .B(n26770), .Z(n26930) );
  NAND U27541 ( .A(n181), .B(n26772), .Z(n26774) );
  XOR U27542 ( .A(b[3]), .B(a[193]), .Z(n26921) );
  NAND U27543 ( .A(n182), .B(n26921), .Z(n26773) );
  AND U27544 ( .A(n26774), .B(n26773), .Z(n26928) );
  NAND U27545 ( .A(n189), .B(n26775), .Z(n26777) );
  XOR U27546 ( .A(b[17]), .B(a[179]), .Z(n26924) );
  NAND U27547 ( .A(n37652), .B(n26924), .Z(n26776) );
  NAND U27548 ( .A(n26777), .B(n26776), .Z(n26927) );
  XNOR U27549 ( .A(n26928), .B(n26927), .Z(n26929) );
  XOR U27550 ( .A(n26930), .B(n26929), .Z(n26962) );
  XOR U27551 ( .A(n26961), .B(n26962), .Z(n26964) );
  XOR U27552 ( .A(n26963), .B(n26964), .Z(n26898) );
  NANDN U27553 ( .A(n26779), .B(n26778), .Z(n26783) );
  NANDN U27554 ( .A(n26781), .B(n26780), .Z(n26782) );
  AND U27555 ( .A(n26783), .B(n26782), .Z(n26951) );
  NANDN U27556 ( .A(n26785), .B(n26784), .Z(n26789) );
  NANDN U27557 ( .A(n26787), .B(n26786), .Z(n26788) );
  NAND U27558 ( .A(n26789), .B(n26788), .Z(n26952) );
  XNOR U27559 ( .A(n26951), .B(n26952), .Z(n26953) );
  NANDN U27560 ( .A(n26791), .B(n26790), .Z(n26795) );
  NANDN U27561 ( .A(n26793), .B(n26792), .Z(n26794) );
  NAND U27562 ( .A(n26795), .B(n26794), .Z(n26954) );
  XNOR U27563 ( .A(n26953), .B(n26954), .Z(n26897) );
  XNOR U27564 ( .A(n26898), .B(n26897), .Z(n26900) );
  NANDN U27565 ( .A(n26797), .B(n26796), .Z(n26801) );
  NANDN U27566 ( .A(n26799), .B(n26798), .Z(n26800) );
  AND U27567 ( .A(n26801), .B(n26800), .Z(n26899) );
  XOR U27568 ( .A(n26900), .B(n26899), .Z(n27012) );
  NANDN U27569 ( .A(n26803), .B(n26802), .Z(n26807) );
  NANDN U27570 ( .A(n26805), .B(n26804), .Z(n26806) );
  AND U27571 ( .A(n26807), .B(n26806), .Z(n27009) );
  NANDN U27572 ( .A(n26809), .B(n26808), .Z(n26813) );
  NANDN U27573 ( .A(n26811), .B(n26810), .Z(n26812) );
  AND U27574 ( .A(n26813), .B(n26812), .Z(n26894) );
  NANDN U27575 ( .A(n26815), .B(n26814), .Z(n26819) );
  OR U27576 ( .A(n26817), .B(n26816), .Z(n26818) );
  AND U27577 ( .A(n26819), .B(n26818), .Z(n26892) );
  NANDN U27578 ( .A(n26821), .B(n26820), .Z(n26825) );
  NANDN U27579 ( .A(n26823), .B(n26822), .Z(n26824) );
  AND U27580 ( .A(n26825), .B(n26824), .Z(n26958) );
  NANDN U27581 ( .A(n26827), .B(n26826), .Z(n26831) );
  NANDN U27582 ( .A(n26829), .B(n26828), .Z(n26830) );
  NAND U27583 ( .A(n26831), .B(n26830), .Z(n26957) );
  XNOR U27584 ( .A(n26958), .B(n26957), .Z(n26960) );
  NAND U27585 ( .A(b[0]), .B(a[195]), .Z(n26832) );
  XNOR U27586 ( .A(b[1]), .B(n26832), .Z(n26834) );
  NANDN U27587 ( .A(b[0]), .B(a[194]), .Z(n26833) );
  NAND U27588 ( .A(n26834), .B(n26833), .Z(n26906) );
  NAND U27589 ( .A(n194), .B(n26835), .Z(n26837) );
  XOR U27590 ( .A(b[29]), .B(a[167]), .Z(n26979) );
  NAND U27591 ( .A(n38456), .B(n26979), .Z(n26836) );
  AND U27592 ( .A(n26837), .B(n26836), .Z(n26904) );
  AND U27593 ( .A(b[31]), .B(a[163]), .Z(n26903) );
  XNOR U27594 ( .A(n26904), .B(n26903), .Z(n26905) );
  XNOR U27595 ( .A(n26906), .B(n26905), .Z(n26946) );
  NAND U27596 ( .A(n38185), .B(n26838), .Z(n26840) );
  XOR U27597 ( .A(b[23]), .B(a[173]), .Z(n26985) );
  NAND U27598 ( .A(n38132), .B(n26985), .Z(n26839) );
  AND U27599 ( .A(n26840), .B(n26839), .Z(n26975) );
  NAND U27600 ( .A(n184), .B(n26841), .Z(n26843) );
  XOR U27601 ( .A(b[7]), .B(a[189]), .Z(n26988) );
  NAND U27602 ( .A(n36592), .B(n26988), .Z(n26842) );
  AND U27603 ( .A(n26843), .B(n26842), .Z(n26974) );
  NAND U27604 ( .A(n38289), .B(n26844), .Z(n26846) );
  XOR U27605 ( .A(b[25]), .B(a[171]), .Z(n26991) );
  NAND U27606 ( .A(n38247), .B(n26991), .Z(n26845) );
  NAND U27607 ( .A(n26846), .B(n26845), .Z(n26973) );
  XOR U27608 ( .A(n26974), .B(n26973), .Z(n26976) );
  XOR U27609 ( .A(n26975), .B(n26976), .Z(n26945) );
  XOR U27610 ( .A(n26946), .B(n26945), .Z(n26948) );
  NAND U27611 ( .A(n187), .B(n26847), .Z(n26849) );
  XOR U27612 ( .A(b[13]), .B(a[183]), .Z(n26994) );
  NAND U27613 ( .A(n37295), .B(n26994), .Z(n26848) );
  AND U27614 ( .A(n26849), .B(n26848), .Z(n26940) );
  NAND U27615 ( .A(n186), .B(n26850), .Z(n26852) );
  XOR U27616 ( .A(b[11]), .B(a[185]), .Z(n26997) );
  NAND U27617 ( .A(n37097), .B(n26997), .Z(n26851) );
  NAND U27618 ( .A(n26852), .B(n26851), .Z(n26939) );
  XNOR U27619 ( .A(n26940), .B(n26939), .Z(n26942) );
  NAND U27620 ( .A(n188), .B(n26853), .Z(n26855) );
  XOR U27621 ( .A(b[15]), .B(a[181]), .Z(n27000) );
  NAND U27622 ( .A(n37382), .B(n27000), .Z(n26854) );
  AND U27623 ( .A(n26855), .B(n26854), .Z(n26936) );
  NAND U27624 ( .A(n38064), .B(n26856), .Z(n26858) );
  XOR U27625 ( .A(b[21]), .B(a[175]), .Z(n27003) );
  NAND U27626 ( .A(n37993), .B(n27003), .Z(n26857) );
  AND U27627 ( .A(n26858), .B(n26857), .Z(n26934) );
  NAND U27628 ( .A(n185), .B(n26859), .Z(n26861) );
  XOR U27629 ( .A(b[9]), .B(a[187]), .Z(n27006) );
  NAND U27630 ( .A(n36805), .B(n27006), .Z(n26860) );
  NAND U27631 ( .A(n26861), .B(n26860), .Z(n26933) );
  XNOR U27632 ( .A(n26934), .B(n26933), .Z(n26935) );
  XNOR U27633 ( .A(n26936), .B(n26935), .Z(n26941) );
  XOR U27634 ( .A(n26942), .B(n26941), .Z(n26947) );
  XNOR U27635 ( .A(n26948), .B(n26947), .Z(n26959) );
  XNOR U27636 ( .A(n26960), .B(n26959), .Z(n26891) );
  XNOR U27637 ( .A(n26892), .B(n26891), .Z(n26893) );
  XOR U27638 ( .A(n26894), .B(n26893), .Z(n27010) );
  XNOR U27639 ( .A(n27009), .B(n27010), .Z(n27011) );
  XNOR U27640 ( .A(n27012), .B(n27011), .Z(n26887) );
  XOR U27641 ( .A(n26888), .B(n26887), .Z(n26880) );
  NANDN U27642 ( .A(n26863), .B(n26862), .Z(n26867) );
  NANDN U27643 ( .A(n26865), .B(n26864), .Z(n26866) );
  AND U27644 ( .A(n26867), .B(n26866), .Z(n26879) );
  XOR U27645 ( .A(n26880), .B(n26879), .Z(n26882) );
  XNOR U27646 ( .A(n26881), .B(n26882), .Z(n26873) );
  XNOR U27647 ( .A(n26874), .B(n26873), .Z(n26875) );
  XNOR U27648 ( .A(n26876), .B(n26875), .Z(n27015) );
  XNOR U27649 ( .A(sreg[419]), .B(n27015), .Z(n27017) );
  NANDN U27650 ( .A(sreg[418]), .B(n26868), .Z(n26872) );
  NAND U27651 ( .A(n26870), .B(n26869), .Z(n26871) );
  NAND U27652 ( .A(n26872), .B(n26871), .Z(n27016) );
  XNOR U27653 ( .A(n27017), .B(n27016), .Z(c[419]) );
  NANDN U27654 ( .A(n26874), .B(n26873), .Z(n26878) );
  NANDN U27655 ( .A(n26876), .B(n26875), .Z(n26877) );
  AND U27656 ( .A(n26878), .B(n26877), .Z(n27023) );
  NANDN U27657 ( .A(n26880), .B(n26879), .Z(n26884) );
  NANDN U27658 ( .A(n26882), .B(n26881), .Z(n26883) );
  AND U27659 ( .A(n26884), .B(n26883), .Z(n27021) );
  NANDN U27660 ( .A(n26886), .B(n26885), .Z(n26890) );
  NAND U27661 ( .A(n26888), .B(n26887), .Z(n26889) );
  AND U27662 ( .A(n26890), .B(n26889), .Z(n27028) );
  NANDN U27663 ( .A(n26892), .B(n26891), .Z(n26896) );
  NANDN U27664 ( .A(n26894), .B(n26893), .Z(n26895) );
  AND U27665 ( .A(n26896), .B(n26895), .Z(n27033) );
  NANDN U27666 ( .A(n26898), .B(n26897), .Z(n26902) );
  NAND U27667 ( .A(n26900), .B(n26899), .Z(n26901) );
  AND U27668 ( .A(n26902), .B(n26901), .Z(n27032) );
  XNOR U27669 ( .A(n27033), .B(n27032), .Z(n27035) );
  NANDN U27670 ( .A(n26904), .B(n26903), .Z(n26908) );
  NANDN U27671 ( .A(n26906), .B(n26905), .Z(n26907) );
  AND U27672 ( .A(n26908), .B(n26907), .Z(n27100) );
  NAND U27673 ( .A(n38385), .B(n26909), .Z(n26911) );
  XOR U27674 ( .A(b[27]), .B(a[170]), .Z(n27044) );
  NAND U27675 ( .A(n38343), .B(n27044), .Z(n26910) );
  AND U27676 ( .A(n26911), .B(n26910), .Z(n27107) );
  NAND U27677 ( .A(n183), .B(n26912), .Z(n26914) );
  XOR U27678 ( .A(b[5]), .B(a[192]), .Z(n27047) );
  NAND U27679 ( .A(n36296), .B(n27047), .Z(n26913) );
  AND U27680 ( .A(n26914), .B(n26913), .Z(n27105) );
  NAND U27681 ( .A(n190), .B(n26915), .Z(n26917) );
  XOR U27682 ( .A(b[19]), .B(a[178]), .Z(n27050) );
  NAND U27683 ( .A(n37821), .B(n27050), .Z(n26916) );
  NAND U27684 ( .A(n26917), .B(n26916), .Z(n27104) );
  XNOR U27685 ( .A(n27105), .B(n27104), .Z(n27106) );
  XNOR U27686 ( .A(n27107), .B(n27106), .Z(n27098) );
  NAND U27687 ( .A(n38470), .B(n26918), .Z(n26920) );
  XOR U27688 ( .A(b[31]), .B(a[166]), .Z(n27053) );
  NAND U27689 ( .A(n38453), .B(n27053), .Z(n26919) );
  AND U27690 ( .A(n26920), .B(n26919), .Z(n27065) );
  NAND U27691 ( .A(n181), .B(n26921), .Z(n26923) );
  XOR U27692 ( .A(b[3]), .B(a[194]), .Z(n27056) );
  NAND U27693 ( .A(n182), .B(n27056), .Z(n26922) );
  AND U27694 ( .A(n26923), .B(n26922), .Z(n27063) );
  NAND U27695 ( .A(n189), .B(n26924), .Z(n26926) );
  XOR U27696 ( .A(b[17]), .B(a[180]), .Z(n27059) );
  NAND U27697 ( .A(n37652), .B(n27059), .Z(n26925) );
  NAND U27698 ( .A(n26926), .B(n26925), .Z(n27062) );
  XNOR U27699 ( .A(n27063), .B(n27062), .Z(n27064) );
  XOR U27700 ( .A(n27065), .B(n27064), .Z(n27099) );
  XOR U27701 ( .A(n27098), .B(n27099), .Z(n27101) );
  XOR U27702 ( .A(n27100), .B(n27101), .Z(n27147) );
  NANDN U27703 ( .A(n26928), .B(n26927), .Z(n26932) );
  NANDN U27704 ( .A(n26930), .B(n26929), .Z(n26931) );
  AND U27705 ( .A(n26932), .B(n26931), .Z(n27086) );
  NANDN U27706 ( .A(n26934), .B(n26933), .Z(n26938) );
  NANDN U27707 ( .A(n26936), .B(n26935), .Z(n26937) );
  NAND U27708 ( .A(n26938), .B(n26937), .Z(n27087) );
  XNOR U27709 ( .A(n27086), .B(n27087), .Z(n27088) );
  NANDN U27710 ( .A(n26940), .B(n26939), .Z(n26944) );
  NAND U27711 ( .A(n26942), .B(n26941), .Z(n26943) );
  NAND U27712 ( .A(n26944), .B(n26943), .Z(n27089) );
  XNOR U27713 ( .A(n27088), .B(n27089), .Z(n27146) );
  XNOR U27714 ( .A(n27147), .B(n27146), .Z(n27149) );
  NAND U27715 ( .A(n26946), .B(n26945), .Z(n26950) );
  NAND U27716 ( .A(n26948), .B(n26947), .Z(n26949) );
  AND U27717 ( .A(n26950), .B(n26949), .Z(n27148) );
  XOR U27718 ( .A(n27149), .B(n27148), .Z(n27161) );
  NANDN U27719 ( .A(n26952), .B(n26951), .Z(n26956) );
  NANDN U27720 ( .A(n26954), .B(n26953), .Z(n26955) );
  AND U27721 ( .A(n26956), .B(n26955), .Z(n27158) );
  NANDN U27722 ( .A(n26962), .B(n26961), .Z(n26966) );
  OR U27723 ( .A(n26964), .B(n26963), .Z(n26965) );
  AND U27724 ( .A(n26966), .B(n26965), .Z(n27153) );
  NANDN U27725 ( .A(n26968), .B(n26967), .Z(n26972) );
  NANDN U27726 ( .A(n26970), .B(n26969), .Z(n26971) );
  AND U27727 ( .A(n26972), .B(n26971), .Z(n27093) );
  NANDN U27728 ( .A(n26974), .B(n26973), .Z(n26978) );
  OR U27729 ( .A(n26976), .B(n26975), .Z(n26977) );
  NAND U27730 ( .A(n26978), .B(n26977), .Z(n27092) );
  XNOR U27731 ( .A(n27093), .B(n27092), .Z(n27094) );
  NAND U27732 ( .A(n194), .B(n26979), .Z(n26981) );
  XOR U27733 ( .A(b[29]), .B(a[168]), .Z(n27116) );
  NAND U27734 ( .A(n38456), .B(n27116), .Z(n26980) );
  AND U27735 ( .A(n26981), .B(n26980), .Z(n27039) );
  AND U27736 ( .A(b[31]), .B(a[164]), .Z(n27038) );
  XNOR U27737 ( .A(n27039), .B(n27038), .Z(n27040) );
  NAND U27738 ( .A(b[0]), .B(a[196]), .Z(n26982) );
  XNOR U27739 ( .A(b[1]), .B(n26982), .Z(n26984) );
  NANDN U27740 ( .A(b[0]), .B(a[195]), .Z(n26983) );
  NAND U27741 ( .A(n26984), .B(n26983), .Z(n27041) );
  XNOR U27742 ( .A(n27040), .B(n27041), .Z(n27080) );
  NAND U27743 ( .A(n38185), .B(n26985), .Z(n26987) );
  XOR U27744 ( .A(b[23]), .B(a[174]), .Z(n27122) );
  NAND U27745 ( .A(n38132), .B(n27122), .Z(n26986) );
  AND U27746 ( .A(n26987), .B(n26986), .Z(n27113) );
  NAND U27747 ( .A(n184), .B(n26988), .Z(n26990) );
  XOR U27748 ( .A(b[7]), .B(a[190]), .Z(n27125) );
  NAND U27749 ( .A(n36592), .B(n27125), .Z(n26989) );
  AND U27750 ( .A(n26990), .B(n26989), .Z(n27111) );
  NAND U27751 ( .A(n38289), .B(n26991), .Z(n26993) );
  XOR U27752 ( .A(b[25]), .B(a[172]), .Z(n27128) );
  NAND U27753 ( .A(n38247), .B(n27128), .Z(n26992) );
  NAND U27754 ( .A(n26993), .B(n26992), .Z(n27110) );
  XNOR U27755 ( .A(n27111), .B(n27110), .Z(n27112) );
  XOR U27756 ( .A(n27113), .B(n27112), .Z(n27081) );
  XNOR U27757 ( .A(n27080), .B(n27081), .Z(n27082) );
  NAND U27758 ( .A(n187), .B(n26994), .Z(n26996) );
  XOR U27759 ( .A(b[13]), .B(a[184]), .Z(n27131) );
  NAND U27760 ( .A(n37295), .B(n27131), .Z(n26995) );
  AND U27761 ( .A(n26996), .B(n26995), .Z(n27075) );
  NAND U27762 ( .A(n186), .B(n26997), .Z(n26999) );
  XOR U27763 ( .A(b[11]), .B(a[186]), .Z(n27134) );
  NAND U27764 ( .A(n37097), .B(n27134), .Z(n26998) );
  NAND U27765 ( .A(n26999), .B(n26998), .Z(n27074) );
  XNOR U27766 ( .A(n27075), .B(n27074), .Z(n27076) );
  NAND U27767 ( .A(n188), .B(n27000), .Z(n27002) );
  XOR U27768 ( .A(b[15]), .B(a[182]), .Z(n27137) );
  NAND U27769 ( .A(n37382), .B(n27137), .Z(n27001) );
  AND U27770 ( .A(n27002), .B(n27001), .Z(n27071) );
  NAND U27771 ( .A(n38064), .B(n27003), .Z(n27005) );
  XOR U27772 ( .A(b[21]), .B(a[176]), .Z(n27140) );
  NAND U27773 ( .A(n37993), .B(n27140), .Z(n27004) );
  AND U27774 ( .A(n27005), .B(n27004), .Z(n27069) );
  NAND U27775 ( .A(n185), .B(n27006), .Z(n27008) );
  XOR U27776 ( .A(b[9]), .B(a[188]), .Z(n27143) );
  NAND U27777 ( .A(n36805), .B(n27143), .Z(n27007) );
  NAND U27778 ( .A(n27008), .B(n27007), .Z(n27068) );
  XNOR U27779 ( .A(n27069), .B(n27068), .Z(n27070) );
  XOR U27780 ( .A(n27071), .B(n27070), .Z(n27077) );
  XOR U27781 ( .A(n27076), .B(n27077), .Z(n27083) );
  XOR U27782 ( .A(n27082), .B(n27083), .Z(n27095) );
  XNOR U27783 ( .A(n27094), .B(n27095), .Z(n27152) );
  XNOR U27784 ( .A(n27153), .B(n27152), .Z(n27154) );
  XOR U27785 ( .A(n27155), .B(n27154), .Z(n27159) );
  XNOR U27786 ( .A(n27158), .B(n27159), .Z(n27160) );
  XNOR U27787 ( .A(n27161), .B(n27160), .Z(n27034) );
  XOR U27788 ( .A(n27035), .B(n27034), .Z(n27027) );
  NANDN U27789 ( .A(n27010), .B(n27009), .Z(n27014) );
  NANDN U27790 ( .A(n27012), .B(n27011), .Z(n27013) );
  AND U27791 ( .A(n27014), .B(n27013), .Z(n27026) );
  XOR U27792 ( .A(n27027), .B(n27026), .Z(n27029) );
  XNOR U27793 ( .A(n27028), .B(n27029), .Z(n27020) );
  XNOR U27794 ( .A(n27021), .B(n27020), .Z(n27022) );
  XNOR U27795 ( .A(n27023), .B(n27022), .Z(n27164) );
  XNOR U27796 ( .A(sreg[420]), .B(n27164), .Z(n27166) );
  NANDN U27797 ( .A(sreg[419]), .B(n27015), .Z(n27019) );
  NAND U27798 ( .A(n27017), .B(n27016), .Z(n27018) );
  NAND U27799 ( .A(n27019), .B(n27018), .Z(n27165) );
  XNOR U27800 ( .A(n27166), .B(n27165), .Z(c[420]) );
  NANDN U27801 ( .A(n27021), .B(n27020), .Z(n27025) );
  NANDN U27802 ( .A(n27023), .B(n27022), .Z(n27024) );
  AND U27803 ( .A(n27025), .B(n27024), .Z(n27172) );
  NANDN U27804 ( .A(n27027), .B(n27026), .Z(n27031) );
  NANDN U27805 ( .A(n27029), .B(n27028), .Z(n27030) );
  AND U27806 ( .A(n27031), .B(n27030), .Z(n27170) );
  NANDN U27807 ( .A(n27033), .B(n27032), .Z(n27037) );
  NAND U27808 ( .A(n27035), .B(n27034), .Z(n27036) );
  AND U27809 ( .A(n27037), .B(n27036), .Z(n27177) );
  NANDN U27810 ( .A(n27039), .B(n27038), .Z(n27043) );
  NANDN U27811 ( .A(n27041), .B(n27040), .Z(n27042) );
  AND U27812 ( .A(n27043), .B(n27042), .Z(n27261) );
  NAND U27813 ( .A(n38385), .B(n27044), .Z(n27046) );
  XOR U27814 ( .A(b[27]), .B(a[171]), .Z(n27205) );
  NAND U27815 ( .A(n38343), .B(n27205), .Z(n27045) );
  AND U27816 ( .A(n27046), .B(n27045), .Z(n27268) );
  NAND U27817 ( .A(n183), .B(n27047), .Z(n27049) );
  XOR U27818 ( .A(b[5]), .B(a[193]), .Z(n27208) );
  NAND U27819 ( .A(n36296), .B(n27208), .Z(n27048) );
  AND U27820 ( .A(n27049), .B(n27048), .Z(n27266) );
  NAND U27821 ( .A(n190), .B(n27050), .Z(n27052) );
  XOR U27822 ( .A(b[19]), .B(a[179]), .Z(n27211) );
  NAND U27823 ( .A(n37821), .B(n27211), .Z(n27051) );
  NAND U27824 ( .A(n27052), .B(n27051), .Z(n27265) );
  XNOR U27825 ( .A(n27266), .B(n27265), .Z(n27267) );
  XNOR U27826 ( .A(n27268), .B(n27267), .Z(n27259) );
  NAND U27827 ( .A(n38470), .B(n27053), .Z(n27055) );
  XOR U27828 ( .A(b[31]), .B(a[167]), .Z(n27214) );
  NAND U27829 ( .A(n38453), .B(n27214), .Z(n27054) );
  AND U27830 ( .A(n27055), .B(n27054), .Z(n27226) );
  NAND U27831 ( .A(n181), .B(n27056), .Z(n27058) );
  XOR U27832 ( .A(b[3]), .B(a[195]), .Z(n27217) );
  NAND U27833 ( .A(n182), .B(n27217), .Z(n27057) );
  AND U27834 ( .A(n27058), .B(n27057), .Z(n27224) );
  NAND U27835 ( .A(n189), .B(n27059), .Z(n27061) );
  XOR U27836 ( .A(b[17]), .B(a[181]), .Z(n27220) );
  NAND U27837 ( .A(n37652), .B(n27220), .Z(n27060) );
  NAND U27838 ( .A(n27061), .B(n27060), .Z(n27223) );
  XNOR U27839 ( .A(n27224), .B(n27223), .Z(n27225) );
  XOR U27840 ( .A(n27226), .B(n27225), .Z(n27260) );
  XOR U27841 ( .A(n27259), .B(n27260), .Z(n27262) );
  XOR U27842 ( .A(n27261), .B(n27262), .Z(n27194) );
  NANDN U27843 ( .A(n27063), .B(n27062), .Z(n27067) );
  NANDN U27844 ( .A(n27065), .B(n27064), .Z(n27066) );
  AND U27845 ( .A(n27067), .B(n27066), .Z(n27247) );
  NANDN U27846 ( .A(n27069), .B(n27068), .Z(n27073) );
  NANDN U27847 ( .A(n27071), .B(n27070), .Z(n27072) );
  NAND U27848 ( .A(n27073), .B(n27072), .Z(n27248) );
  XNOR U27849 ( .A(n27247), .B(n27248), .Z(n27249) );
  NANDN U27850 ( .A(n27075), .B(n27074), .Z(n27079) );
  NANDN U27851 ( .A(n27077), .B(n27076), .Z(n27078) );
  NAND U27852 ( .A(n27079), .B(n27078), .Z(n27250) );
  XNOR U27853 ( .A(n27249), .B(n27250), .Z(n27193) );
  XNOR U27854 ( .A(n27194), .B(n27193), .Z(n27196) );
  NANDN U27855 ( .A(n27081), .B(n27080), .Z(n27085) );
  NANDN U27856 ( .A(n27083), .B(n27082), .Z(n27084) );
  AND U27857 ( .A(n27085), .B(n27084), .Z(n27195) );
  XOR U27858 ( .A(n27196), .B(n27195), .Z(n27309) );
  NANDN U27859 ( .A(n27087), .B(n27086), .Z(n27091) );
  NANDN U27860 ( .A(n27089), .B(n27088), .Z(n27090) );
  AND U27861 ( .A(n27091), .B(n27090), .Z(n27307) );
  NANDN U27862 ( .A(n27093), .B(n27092), .Z(n27097) );
  NANDN U27863 ( .A(n27095), .B(n27094), .Z(n27096) );
  AND U27864 ( .A(n27097), .B(n27096), .Z(n27190) );
  NANDN U27865 ( .A(n27099), .B(n27098), .Z(n27103) );
  OR U27866 ( .A(n27101), .B(n27100), .Z(n27102) );
  AND U27867 ( .A(n27103), .B(n27102), .Z(n27188) );
  NANDN U27868 ( .A(n27105), .B(n27104), .Z(n27109) );
  NANDN U27869 ( .A(n27107), .B(n27106), .Z(n27108) );
  AND U27870 ( .A(n27109), .B(n27108), .Z(n27254) );
  NANDN U27871 ( .A(n27111), .B(n27110), .Z(n27115) );
  NANDN U27872 ( .A(n27113), .B(n27112), .Z(n27114) );
  NAND U27873 ( .A(n27115), .B(n27114), .Z(n27253) );
  XNOR U27874 ( .A(n27254), .B(n27253), .Z(n27255) );
  NAND U27875 ( .A(n194), .B(n27116), .Z(n27118) );
  XOR U27876 ( .A(b[29]), .B(a[169]), .Z(n27277) );
  NAND U27877 ( .A(n38456), .B(n27277), .Z(n27117) );
  AND U27878 ( .A(n27118), .B(n27117), .Z(n27200) );
  AND U27879 ( .A(b[31]), .B(a[165]), .Z(n27199) );
  XNOR U27880 ( .A(n27200), .B(n27199), .Z(n27201) );
  NAND U27881 ( .A(b[0]), .B(a[197]), .Z(n27119) );
  XNOR U27882 ( .A(b[1]), .B(n27119), .Z(n27121) );
  NANDN U27883 ( .A(b[0]), .B(a[196]), .Z(n27120) );
  NAND U27884 ( .A(n27121), .B(n27120), .Z(n27202) );
  XNOR U27885 ( .A(n27201), .B(n27202), .Z(n27241) );
  NAND U27886 ( .A(n38185), .B(n27122), .Z(n27124) );
  XOR U27887 ( .A(b[23]), .B(a[175]), .Z(n27283) );
  NAND U27888 ( .A(n38132), .B(n27283), .Z(n27123) );
  AND U27889 ( .A(n27124), .B(n27123), .Z(n27274) );
  NAND U27890 ( .A(n184), .B(n27125), .Z(n27127) );
  XOR U27891 ( .A(b[7]), .B(a[191]), .Z(n27286) );
  NAND U27892 ( .A(n36592), .B(n27286), .Z(n27126) );
  AND U27893 ( .A(n27127), .B(n27126), .Z(n27272) );
  NAND U27894 ( .A(n38289), .B(n27128), .Z(n27130) );
  XOR U27895 ( .A(b[25]), .B(a[173]), .Z(n27289) );
  NAND U27896 ( .A(n38247), .B(n27289), .Z(n27129) );
  NAND U27897 ( .A(n27130), .B(n27129), .Z(n27271) );
  XNOR U27898 ( .A(n27272), .B(n27271), .Z(n27273) );
  XOR U27899 ( .A(n27274), .B(n27273), .Z(n27242) );
  XNOR U27900 ( .A(n27241), .B(n27242), .Z(n27243) );
  NAND U27901 ( .A(n187), .B(n27131), .Z(n27133) );
  XOR U27902 ( .A(b[13]), .B(a[185]), .Z(n27292) );
  NAND U27903 ( .A(n37295), .B(n27292), .Z(n27132) );
  AND U27904 ( .A(n27133), .B(n27132), .Z(n27236) );
  NAND U27905 ( .A(n186), .B(n27134), .Z(n27136) );
  XOR U27906 ( .A(b[11]), .B(a[187]), .Z(n27295) );
  NAND U27907 ( .A(n37097), .B(n27295), .Z(n27135) );
  NAND U27908 ( .A(n27136), .B(n27135), .Z(n27235) );
  XNOR U27909 ( .A(n27236), .B(n27235), .Z(n27237) );
  NAND U27910 ( .A(n188), .B(n27137), .Z(n27139) );
  XOR U27911 ( .A(b[15]), .B(a[183]), .Z(n27298) );
  NAND U27912 ( .A(n37382), .B(n27298), .Z(n27138) );
  AND U27913 ( .A(n27139), .B(n27138), .Z(n27232) );
  NAND U27914 ( .A(n38064), .B(n27140), .Z(n27142) );
  XOR U27915 ( .A(b[21]), .B(a[177]), .Z(n27301) );
  NAND U27916 ( .A(n37993), .B(n27301), .Z(n27141) );
  AND U27917 ( .A(n27142), .B(n27141), .Z(n27230) );
  NAND U27918 ( .A(n185), .B(n27143), .Z(n27145) );
  XOR U27919 ( .A(b[9]), .B(a[189]), .Z(n27304) );
  NAND U27920 ( .A(n36805), .B(n27304), .Z(n27144) );
  NAND U27921 ( .A(n27145), .B(n27144), .Z(n27229) );
  XNOR U27922 ( .A(n27230), .B(n27229), .Z(n27231) );
  XOR U27923 ( .A(n27232), .B(n27231), .Z(n27238) );
  XOR U27924 ( .A(n27237), .B(n27238), .Z(n27244) );
  XOR U27925 ( .A(n27243), .B(n27244), .Z(n27256) );
  XNOR U27926 ( .A(n27255), .B(n27256), .Z(n27187) );
  XNOR U27927 ( .A(n27188), .B(n27187), .Z(n27189) );
  XOR U27928 ( .A(n27190), .B(n27189), .Z(n27308) );
  XOR U27929 ( .A(n27307), .B(n27308), .Z(n27310) );
  XOR U27930 ( .A(n27309), .B(n27310), .Z(n27184) );
  NANDN U27931 ( .A(n27147), .B(n27146), .Z(n27151) );
  NAND U27932 ( .A(n27149), .B(n27148), .Z(n27150) );
  AND U27933 ( .A(n27151), .B(n27150), .Z(n27182) );
  NANDN U27934 ( .A(n27153), .B(n27152), .Z(n27157) );
  NANDN U27935 ( .A(n27155), .B(n27154), .Z(n27156) );
  AND U27936 ( .A(n27157), .B(n27156), .Z(n27181) );
  XNOR U27937 ( .A(n27182), .B(n27181), .Z(n27183) );
  XNOR U27938 ( .A(n27184), .B(n27183), .Z(n27175) );
  NANDN U27939 ( .A(n27159), .B(n27158), .Z(n27163) );
  NANDN U27940 ( .A(n27161), .B(n27160), .Z(n27162) );
  NAND U27941 ( .A(n27163), .B(n27162), .Z(n27176) );
  XOR U27942 ( .A(n27175), .B(n27176), .Z(n27178) );
  XNOR U27943 ( .A(n27177), .B(n27178), .Z(n27169) );
  XNOR U27944 ( .A(n27170), .B(n27169), .Z(n27171) );
  XNOR U27945 ( .A(n27172), .B(n27171), .Z(n27313) );
  XNOR U27946 ( .A(sreg[421]), .B(n27313), .Z(n27315) );
  NANDN U27947 ( .A(sreg[420]), .B(n27164), .Z(n27168) );
  NAND U27948 ( .A(n27166), .B(n27165), .Z(n27167) );
  NAND U27949 ( .A(n27168), .B(n27167), .Z(n27314) );
  XNOR U27950 ( .A(n27315), .B(n27314), .Z(c[421]) );
  NANDN U27951 ( .A(n27170), .B(n27169), .Z(n27174) );
  NANDN U27952 ( .A(n27172), .B(n27171), .Z(n27173) );
  AND U27953 ( .A(n27174), .B(n27173), .Z(n27321) );
  NANDN U27954 ( .A(n27176), .B(n27175), .Z(n27180) );
  NANDN U27955 ( .A(n27178), .B(n27177), .Z(n27179) );
  AND U27956 ( .A(n27180), .B(n27179), .Z(n27319) );
  NANDN U27957 ( .A(n27182), .B(n27181), .Z(n27186) );
  NANDN U27958 ( .A(n27184), .B(n27183), .Z(n27185) );
  AND U27959 ( .A(n27186), .B(n27185), .Z(n27327) );
  NANDN U27960 ( .A(n27188), .B(n27187), .Z(n27192) );
  NANDN U27961 ( .A(n27190), .B(n27189), .Z(n27191) );
  AND U27962 ( .A(n27192), .B(n27191), .Z(n27331) );
  NANDN U27963 ( .A(n27194), .B(n27193), .Z(n27198) );
  NAND U27964 ( .A(n27196), .B(n27195), .Z(n27197) );
  AND U27965 ( .A(n27198), .B(n27197), .Z(n27330) );
  XNOR U27966 ( .A(n27331), .B(n27330), .Z(n27333) );
  NANDN U27967 ( .A(n27200), .B(n27199), .Z(n27204) );
  NANDN U27968 ( .A(n27202), .B(n27201), .Z(n27203) );
  AND U27969 ( .A(n27204), .B(n27203), .Z(n27410) );
  NAND U27970 ( .A(n38385), .B(n27205), .Z(n27207) );
  XOR U27971 ( .A(b[27]), .B(a[172]), .Z(n27354) );
  NAND U27972 ( .A(n38343), .B(n27354), .Z(n27206) );
  AND U27973 ( .A(n27207), .B(n27206), .Z(n27417) );
  NAND U27974 ( .A(n183), .B(n27208), .Z(n27210) );
  XOR U27975 ( .A(b[5]), .B(a[194]), .Z(n27357) );
  NAND U27976 ( .A(n36296), .B(n27357), .Z(n27209) );
  AND U27977 ( .A(n27210), .B(n27209), .Z(n27415) );
  NAND U27978 ( .A(n190), .B(n27211), .Z(n27213) );
  XOR U27979 ( .A(b[19]), .B(a[180]), .Z(n27360) );
  NAND U27980 ( .A(n37821), .B(n27360), .Z(n27212) );
  NAND U27981 ( .A(n27213), .B(n27212), .Z(n27414) );
  XNOR U27982 ( .A(n27415), .B(n27414), .Z(n27416) );
  XNOR U27983 ( .A(n27417), .B(n27416), .Z(n27408) );
  NAND U27984 ( .A(n38470), .B(n27214), .Z(n27216) );
  XOR U27985 ( .A(b[31]), .B(a[168]), .Z(n27363) );
  NAND U27986 ( .A(n38453), .B(n27363), .Z(n27215) );
  AND U27987 ( .A(n27216), .B(n27215), .Z(n27375) );
  NAND U27988 ( .A(n181), .B(n27217), .Z(n27219) );
  XOR U27989 ( .A(b[3]), .B(a[196]), .Z(n27366) );
  NAND U27990 ( .A(n182), .B(n27366), .Z(n27218) );
  AND U27991 ( .A(n27219), .B(n27218), .Z(n27373) );
  NAND U27992 ( .A(n189), .B(n27220), .Z(n27222) );
  XOR U27993 ( .A(b[17]), .B(a[182]), .Z(n27369) );
  NAND U27994 ( .A(n37652), .B(n27369), .Z(n27221) );
  NAND U27995 ( .A(n27222), .B(n27221), .Z(n27372) );
  XNOR U27996 ( .A(n27373), .B(n27372), .Z(n27374) );
  XOR U27997 ( .A(n27375), .B(n27374), .Z(n27409) );
  XOR U27998 ( .A(n27408), .B(n27409), .Z(n27411) );
  XOR U27999 ( .A(n27410), .B(n27411), .Z(n27343) );
  NANDN U28000 ( .A(n27224), .B(n27223), .Z(n27228) );
  NANDN U28001 ( .A(n27226), .B(n27225), .Z(n27227) );
  AND U28002 ( .A(n27228), .B(n27227), .Z(n27396) );
  NANDN U28003 ( .A(n27230), .B(n27229), .Z(n27234) );
  NANDN U28004 ( .A(n27232), .B(n27231), .Z(n27233) );
  NAND U28005 ( .A(n27234), .B(n27233), .Z(n27397) );
  XNOR U28006 ( .A(n27396), .B(n27397), .Z(n27398) );
  NANDN U28007 ( .A(n27236), .B(n27235), .Z(n27240) );
  NANDN U28008 ( .A(n27238), .B(n27237), .Z(n27239) );
  NAND U28009 ( .A(n27240), .B(n27239), .Z(n27399) );
  XNOR U28010 ( .A(n27398), .B(n27399), .Z(n27342) );
  XNOR U28011 ( .A(n27343), .B(n27342), .Z(n27345) );
  NANDN U28012 ( .A(n27242), .B(n27241), .Z(n27246) );
  NANDN U28013 ( .A(n27244), .B(n27243), .Z(n27245) );
  AND U28014 ( .A(n27246), .B(n27245), .Z(n27344) );
  XOR U28015 ( .A(n27345), .B(n27344), .Z(n27459) );
  NANDN U28016 ( .A(n27248), .B(n27247), .Z(n27252) );
  NANDN U28017 ( .A(n27250), .B(n27249), .Z(n27251) );
  AND U28018 ( .A(n27252), .B(n27251), .Z(n27456) );
  NANDN U28019 ( .A(n27254), .B(n27253), .Z(n27258) );
  NANDN U28020 ( .A(n27256), .B(n27255), .Z(n27257) );
  AND U28021 ( .A(n27258), .B(n27257), .Z(n27339) );
  NANDN U28022 ( .A(n27260), .B(n27259), .Z(n27264) );
  OR U28023 ( .A(n27262), .B(n27261), .Z(n27263) );
  AND U28024 ( .A(n27264), .B(n27263), .Z(n27337) );
  NANDN U28025 ( .A(n27266), .B(n27265), .Z(n27270) );
  NANDN U28026 ( .A(n27268), .B(n27267), .Z(n27269) );
  AND U28027 ( .A(n27270), .B(n27269), .Z(n27403) );
  NANDN U28028 ( .A(n27272), .B(n27271), .Z(n27276) );
  NANDN U28029 ( .A(n27274), .B(n27273), .Z(n27275) );
  NAND U28030 ( .A(n27276), .B(n27275), .Z(n27402) );
  XNOR U28031 ( .A(n27403), .B(n27402), .Z(n27404) );
  NAND U28032 ( .A(n194), .B(n27277), .Z(n27279) );
  XOR U28033 ( .A(b[29]), .B(a[170]), .Z(n27429) );
  NAND U28034 ( .A(n38456), .B(n27429), .Z(n27278) );
  AND U28035 ( .A(n27279), .B(n27278), .Z(n27349) );
  AND U28036 ( .A(b[31]), .B(a[166]), .Z(n27348) );
  XNOR U28037 ( .A(n27349), .B(n27348), .Z(n27350) );
  NAND U28038 ( .A(b[0]), .B(a[198]), .Z(n27280) );
  XNOR U28039 ( .A(b[1]), .B(n27280), .Z(n27282) );
  NANDN U28040 ( .A(b[0]), .B(a[197]), .Z(n27281) );
  NAND U28041 ( .A(n27282), .B(n27281), .Z(n27351) );
  XNOR U28042 ( .A(n27350), .B(n27351), .Z(n27390) );
  NAND U28043 ( .A(n38185), .B(n27283), .Z(n27285) );
  XOR U28044 ( .A(b[23]), .B(a[176]), .Z(n27432) );
  NAND U28045 ( .A(n38132), .B(n27432), .Z(n27284) );
  AND U28046 ( .A(n27285), .B(n27284), .Z(n27423) );
  NAND U28047 ( .A(n184), .B(n27286), .Z(n27288) );
  XOR U28048 ( .A(b[7]), .B(a[192]), .Z(n27435) );
  NAND U28049 ( .A(n36592), .B(n27435), .Z(n27287) );
  AND U28050 ( .A(n27288), .B(n27287), .Z(n27421) );
  NAND U28051 ( .A(n38289), .B(n27289), .Z(n27291) );
  XOR U28052 ( .A(b[25]), .B(a[174]), .Z(n27438) );
  NAND U28053 ( .A(n38247), .B(n27438), .Z(n27290) );
  NAND U28054 ( .A(n27291), .B(n27290), .Z(n27420) );
  XNOR U28055 ( .A(n27421), .B(n27420), .Z(n27422) );
  XOR U28056 ( .A(n27423), .B(n27422), .Z(n27391) );
  XNOR U28057 ( .A(n27390), .B(n27391), .Z(n27392) );
  NAND U28058 ( .A(n187), .B(n27292), .Z(n27294) );
  XOR U28059 ( .A(b[13]), .B(a[186]), .Z(n27441) );
  NAND U28060 ( .A(n37295), .B(n27441), .Z(n27293) );
  AND U28061 ( .A(n27294), .B(n27293), .Z(n27385) );
  NAND U28062 ( .A(n186), .B(n27295), .Z(n27297) );
  XOR U28063 ( .A(b[11]), .B(a[188]), .Z(n27444) );
  NAND U28064 ( .A(n37097), .B(n27444), .Z(n27296) );
  NAND U28065 ( .A(n27297), .B(n27296), .Z(n27384) );
  XNOR U28066 ( .A(n27385), .B(n27384), .Z(n27386) );
  NAND U28067 ( .A(n188), .B(n27298), .Z(n27300) );
  XOR U28068 ( .A(b[15]), .B(a[184]), .Z(n27447) );
  NAND U28069 ( .A(n37382), .B(n27447), .Z(n27299) );
  AND U28070 ( .A(n27300), .B(n27299), .Z(n27381) );
  NAND U28071 ( .A(n38064), .B(n27301), .Z(n27303) );
  XOR U28072 ( .A(b[21]), .B(a[178]), .Z(n27450) );
  NAND U28073 ( .A(n37993), .B(n27450), .Z(n27302) );
  AND U28074 ( .A(n27303), .B(n27302), .Z(n27379) );
  NAND U28075 ( .A(n185), .B(n27304), .Z(n27306) );
  XOR U28076 ( .A(b[9]), .B(a[190]), .Z(n27453) );
  NAND U28077 ( .A(n36805), .B(n27453), .Z(n27305) );
  NAND U28078 ( .A(n27306), .B(n27305), .Z(n27378) );
  XNOR U28079 ( .A(n27379), .B(n27378), .Z(n27380) );
  XOR U28080 ( .A(n27381), .B(n27380), .Z(n27387) );
  XOR U28081 ( .A(n27386), .B(n27387), .Z(n27393) );
  XOR U28082 ( .A(n27392), .B(n27393), .Z(n27405) );
  XNOR U28083 ( .A(n27404), .B(n27405), .Z(n27336) );
  XNOR U28084 ( .A(n27337), .B(n27336), .Z(n27338) );
  XOR U28085 ( .A(n27339), .B(n27338), .Z(n27457) );
  XNOR U28086 ( .A(n27456), .B(n27457), .Z(n27458) );
  XNOR U28087 ( .A(n27459), .B(n27458), .Z(n27332) );
  XOR U28088 ( .A(n27333), .B(n27332), .Z(n27325) );
  NANDN U28089 ( .A(n27308), .B(n27307), .Z(n27312) );
  OR U28090 ( .A(n27310), .B(n27309), .Z(n27311) );
  AND U28091 ( .A(n27312), .B(n27311), .Z(n27324) );
  XNOR U28092 ( .A(n27325), .B(n27324), .Z(n27326) );
  XNOR U28093 ( .A(n27327), .B(n27326), .Z(n27318) );
  XNOR U28094 ( .A(n27319), .B(n27318), .Z(n27320) );
  XNOR U28095 ( .A(n27321), .B(n27320), .Z(n27462) );
  XNOR U28096 ( .A(sreg[422]), .B(n27462), .Z(n27464) );
  NANDN U28097 ( .A(sreg[421]), .B(n27313), .Z(n27317) );
  NAND U28098 ( .A(n27315), .B(n27314), .Z(n27316) );
  NAND U28099 ( .A(n27317), .B(n27316), .Z(n27463) );
  XNOR U28100 ( .A(n27464), .B(n27463), .Z(c[422]) );
  NANDN U28101 ( .A(n27319), .B(n27318), .Z(n27323) );
  NANDN U28102 ( .A(n27321), .B(n27320), .Z(n27322) );
  AND U28103 ( .A(n27323), .B(n27322), .Z(n27470) );
  NANDN U28104 ( .A(n27325), .B(n27324), .Z(n27329) );
  NANDN U28105 ( .A(n27327), .B(n27326), .Z(n27328) );
  AND U28106 ( .A(n27329), .B(n27328), .Z(n27468) );
  NANDN U28107 ( .A(n27331), .B(n27330), .Z(n27335) );
  NAND U28108 ( .A(n27333), .B(n27332), .Z(n27334) );
  AND U28109 ( .A(n27335), .B(n27334), .Z(n27475) );
  NANDN U28110 ( .A(n27337), .B(n27336), .Z(n27341) );
  NANDN U28111 ( .A(n27339), .B(n27338), .Z(n27340) );
  AND U28112 ( .A(n27341), .B(n27340), .Z(n27606) );
  NANDN U28113 ( .A(n27343), .B(n27342), .Z(n27347) );
  NAND U28114 ( .A(n27345), .B(n27344), .Z(n27346) );
  AND U28115 ( .A(n27347), .B(n27346), .Z(n27605) );
  XNOR U28116 ( .A(n27606), .B(n27605), .Z(n27608) );
  NANDN U28117 ( .A(n27349), .B(n27348), .Z(n27353) );
  NANDN U28118 ( .A(n27351), .B(n27350), .Z(n27352) );
  AND U28119 ( .A(n27353), .B(n27352), .Z(n27553) );
  NAND U28120 ( .A(n38385), .B(n27354), .Z(n27356) );
  XOR U28121 ( .A(b[27]), .B(a[173]), .Z(n27497) );
  NAND U28122 ( .A(n38343), .B(n27497), .Z(n27355) );
  AND U28123 ( .A(n27356), .B(n27355), .Z(n27560) );
  NAND U28124 ( .A(n183), .B(n27357), .Z(n27359) );
  XOR U28125 ( .A(b[5]), .B(a[195]), .Z(n27500) );
  NAND U28126 ( .A(n36296), .B(n27500), .Z(n27358) );
  AND U28127 ( .A(n27359), .B(n27358), .Z(n27558) );
  NAND U28128 ( .A(n190), .B(n27360), .Z(n27362) );
  XOR U28129 ( .A(b[19]), .B(a[181]), .Z(n27503) );
  NAND U28130 ( .A(n37821), .B(n27503), .Z(n27361) );
  NAND U28131 ( .A(n27362), .B(n27361), .Z(n27557) );
  XNOR U28132 ( .A(n27558), .B(n27557), .Z(n27559) );
  XNOR U28133 ( .A(n27560), .B(n27559), .Z(n27551) );
  NAND U28134 ( .A(n38470), .B(n27363), .Z(n27365) );
  XOR U28135 ( .A(b[31]), .B(a[169]), .Z(n27506) );
  NAND U28136 ( .A(n38453), .B(n27506), .Z(n27364) );
  AND U28137 ( .A(n27365), .B(n27364), .Z(n27518) );
  NAND U28138 ( .A(n181), .B(n27366), .Z(n27368) );
  XOR U28139 ( .A(b[3]), .B(a[197]), .Z(n27509) );
  NAND U28140 ( .A(n182), .B(n27509), .Z(n27367) );
  AND U28141 ( .A(n27368), .B(n27367), .Z(n27516) );
  NAND U28142 ( .A(n189), .B(n27369), .Z(n27371) );
  XOR U28143 ( .A(b[17]), .B(a[183]), .Z(n27512) );
  NAND U28144 ( .A(n37652), .B(n27512), .Z(n27370) );
  NAND U28145 ( .A(n27371), .B(n27370), .Z(n27515) );
  XNOR U28146 ( .A(n27516), .B(n27515), .Z(n27517) );
  XOR U28147 ( .A(n27518), .B(n27517), .Z(n27552) );
  XOR U28148 ( .A(n27551), .B(n27552), .Z(n27554) );
  XOR U28149 ( .A(n27553), .B(n27554), .Z(n27486) );
  NANDN U28150 ( .A(n27373), .B(n27372), .Z(n27377) );
  NANDN U28151 ( .A(n27375), .B(n27374), .Z(n27376) );
  AND U28152 ( .A(n27377), .B(n27376), .Z(n27539) );
  NANDN U28153 ( .A(n27379), .B(n27378), .Z(n27383) );
  NANDN U28154 ( .A(n27381), .B(n27380), .Z(n27382) );
  NAND U28155 ( .A(n27383), .B(n27382), .Z(n27540) );
  XNOR U28156 ( .A(n27539), .B(n27540), .Z(n27541) );
  NANDN U28157 ( .A(n27385), .B(n27384), .Z(n27389) );
  NANDN U28158 ( .A(n27387), .B(n27386), .Z(n27388) );
  NAND U28159 ( .A(n27389), .B(n27388), .Z(n27542) );
  XNOR U28160 ( .A(n27541), .B(n27542), .Z(n27485) );
  XNOR U28161 ( .A(n27486), .B(n27485), .Z(n27488) );
  NANDN U28162 ( .A(n27391), .B(n27390), .Z(n27395) );
  NANDN U28163 ( .A(n27393), .B(n27392), .Z(n27394) );
  AND U28164 ( .A(n27395), .B(n27394), .Z(n27487) );
  XOR U28165 ( .A(n27488), .B(n27487), .Z(n27602) );
  NANDN U28166 ( .A(n27397), .B(n27396), .Z(n27401) );
  NANDN U28167 ( .A(n27399), .B(n27398), .Z(n27400) );
  AND U28168 ( .A(n27401), .B(n27400), .Z(n27599) );
  NANDN U28169 ( .A(n27403), .B(n27402), .Z(n27407) );
  NANDN U28170 ( .A(n27405), .B(n27404), .Z(n27406) );
  AND U28171 ( .A(n27407), .B(n27406), .Z(n27482) );
  NANDN U28172 ( .A(n27409), .B(n27408), .Z(n27413) );
  OR U28173 ( .A(n27411), .B(n27410), .Z(n27412) );
  AND U28174 ( .A(n27413), .B(n27412), .Z(n27480) );
  NANDN U28175 ( .A(n27415), .B(n27414), .Z(n27419) );
  NANDN U28176 ( .A(n27417), .B(n27416), .Z(n27418) );
  AND U28177 ( .A(n27419), .B(n27418), .Z(n27546) );
  NANDN U28178 ( .A(n27421), .B(n27420), .Z(n27425) );
  NANDN U28179 ( .A(n27423), .B(n27422), .Z(n27424) );
  NAND U28180 ( .A(n27425), .B(n27424), .Z(n27545) );
  XNOR U28181 ( .A(n27546), .B(n27545), .Z(n27547) );
  NAND U28182 ( .A(b[0]), .B(a[199]), .Z(n27426) );
  XNOR U28183 ( .A(b[1]), .B(n27426), .Z(n27428) );
  NANDN U28184 ( .A(b[0]), .B(a[198]), .Z(n27427) );
  NAND U28185 ( .A(n27428), .B(n27427), .Z(n27494) );
  NAND U28186 ( .A(n194), .B(n27429), .Z(n27431) );
  XOR U28187 ( .A(b[29]), .B(a[171]), .Z(n27572) );
  NAND U28188 ( .A(n38456), .B(n27572), .Z(n27430) );
  AND U28189 ( .A(n27431), .B(n27430), .Z(n27492) );
  AND U28190 ( .A(b[31]), .B(a[167]), .Z(n27491) );
  XNOR U28191 ( .A(n27492), .B(n27491), .Z(n27493) );
  XNOR U28192 ( .A(n27494), .B(n27493), .Z(n27533) );
  NAND U28193 ( .A(n38185), .B(n27432), .Z(n27434) );
  XOR U28194 ( .A(b[23]), .B(a[177]), .Z(n27575) );
  NAND U28195 ( .A(n38132), .B(n27575), .Z(n27433) );
  AND U28196 ( .A(n27434), .B(n27433), .Z(n27566) );
  NAND U28197 ( .A(n184), .B(n27435), .Z(n27437) );
  XOR U28198 ( .A(b[7]), .B(a[193]), .Z(n27578) );
  NAND U28199 ( .A(n36592), .B(n27578), .Z(n27436) );
  AND U28200 ( .A(n27437), .B(n27436), .Z(n27564) );
  NAND U28201 ( .A(n38289), .B(n27438), .Z(n27440) );
  XOR U28202 ( .A(b[25]), .B(a[175]), .Z(n27581) );
  NAND U28203 ( .A(n38247), .B(n27581), .Z(n27439) );
  NAND U28204 ( .A(n27440), .B(n27439), .Z(n27563) );
  XNOR U28205 ( .A(n27564), .B(n27563), .Z(n27565) );
  XOR U28206 ( .A(n27566), .B(n27565), .Z(n27534) );
  XNOR U28207 ( .A(n27533), .B(n27534), .Z(n27535) );
  NAND U28208 ( .A(n187), .B(n27441), .Z(n27443) );
  XOR U28209 ( .A(b[13]), .B(a[187]), .Z(n27584) );
  NAND U28210 ( .A(n37295), .B(n27584), .Z(n27442) );
  AND U28211 ( .A(n27443), .B(n27442), .Z(n27528) );
  NAND U28212 ( .A(n186), .B(n27444), .Z(n27446) );
  XOR U28213 ( .A(b[11]), .B(a[189]), .Z(n27587) );
  NAND U28214 ( .A(n37097), .B(n27587), .Z(n27445) );
  NAND U28215 ( .A(n27446), .B(n27445), .Z(n27527) );
  XNOR U28216 ( .A(n27528), .B(n27527), .Z(n27529) );
  NAND U28217 ( .A(n188), .B(n27447), .Z(n27449) );
  XOR U28218 ( .A(b[15]), .B(a[185]), .Z(n27590) );
  NAND U28219 ( .A(n37382), .B(n27590), .Z(n27448) );
  AND U28220 ( .A(n27449), .B(n27448), .Z(n27524) );
  NAND U28221 ( .A(n38064), .B(n27450), .Z(n27452) );
  XOR U28222 ( .A(b[21]), .B(a[179]), .Z(n27593) );
  NAND U28223 ( .A(n37993), .B(n27593), .Z(n27451) );
  AND U28224 ( .A(n27452), .B(n27451), .Z(n27522) );
  NAND U28225 ( .A(n185), .B(n27453), .Z(n27455) );
  XOR U28226 ( .A(b[9]), .B(a[191]), .Z(n27596) );
  NAND U28227 ( .A(n36805), .B(n27596), .Z(n27454) );
  NAND U28228 ( .A(n27455), .B(n27454), .Z(n27521) );
  XNOR U28229 ( .A(n27522), .B(n27521), .Z(n27523) );
  XOR U28230 ( .A(n27524), .B(n27523), .Z(n27530) );
  XOR U28231 ( .A(n27529), .B(n27530), .Z(n27536) );
  XOR U28232 ( .A(n27535), .B(n27536), .Z(n27548) );
  XNOR U28233 ( .A(n27547), .B(n27548), .Z(n27479) );
  XNOR U28234 ( .A(n27480), .B(n27479), .Z(n27481) );
  XOR U28235 ( .A(n27482), .B(n27481), .Z(n27600) );
  XNOR U28236 ( .A(n27599), .B(n27600), .Z(n27601) );
  XNOR U28237 ( .A(n27602), .B(n27601), .Z(n27607) );
  XOR U28238 ( .A(n27608), .B(n27607), .Z(n27474) );
  NANDN U28239 ( .A(n27457), .B(n27456), .Z(n27461) );
  NANDN U28240 ( .A(n27459), .B(n27458), .Z(n27460) );
  AND U28241 ( .A(n27461), .B(n27460), .Z(n27473) );
  XOR U28242 ( .A(n27474), .B(n27473), .Z(n27476) );
  XNOR U28243 ( .A(n27475), .B(n27476), .Z(n27467) );
  XNOR U28244 ( .A(n27468), .B(n27467), .Z(n27469) );
  XNOR U28245 ( .A(n27470), .B(n27469), .Z(n27611) );
  XNOR U28246 ( .A(sreg[423]), .B(n27611), .Z(n27613) );
  NANDN U28247 ( .A(sreg[422]), .B(n27462), .Z(n27466) );
  NAND U28248 ( .A(n27464), .B(n27463), .Z(n27465) );
  NAND U28249 ( .A(n27466), .B(n27465), .Z(n27612) );
  XNOR U28250 ( .A(n27613), .B(n27612), .Z(c[423]) );
  NANDN U28251 ( .A(n27468), .B(n27467), .Z(n27472) );
  NANDN U28252 ( .A(n27470), .B(n27469), .Z(n27471) );
  AND U28253 ( .A(n27472), .B(n27471), .Z(n27619) );
  NANDN U28254 ( .A(n27474), .B(n27473), .Z(n27478) );
  NANDN U28255 ( .A(n27476), .B(n27475), .Z(n27477) );
  AND U28256 ( .A(n27478), .B(n27477), .Z(n27617) );
  NANDN U28257 ( .A(n27480), .B(n27479), .Z(n27484) );
  NANDN U28258 ( .A(n27482), .B(n27481), .Z(n27483) );
  AND U28259 ( .A(n27484), .B(n27483), .Z(n27629) );
  NANDN U28260 ( .A(n27486), .B(n27485), .Z(n27490) );
  NAND U28261 ( .A(n27488), .B(n27487), .Z(n27489) );
  AND U28262 ( .A(n27490), .B(n27489), .Z(n27628) );
  XNOR U28263 ( .A(n27629), .B(n27628), .Z(n27631) );
  NANDN U28264 ( .A(n27492), .B(n27491), .Z(n27496) );
  NANDN U28265 ( .A(n27494), .B(n27493), .Z(n27495) );
  AND U28266 ( .A(n27496), .B(n27495), .Z(n27708) );
  NAND U28267 ( .A(n38385), .B(n27497), .Z(n27499) );
  XOR U28268 ( .A(b[27]), .B(a[174]), .Z(n27652) );
  NAND U28269 ( .A(n38343), .B(n27652), .Z(n27498) );
  AND U28270 ( .A(n27499), .B(n27498), .Z(n27715) );
  NAND U28271 ( .A(n183), .B(n27500), .Z(n27502) );
  XOR U28272 ( .A(b[5]), .B(a[196]), .Z(n27655) );
  NAND U28273 ( .A(n36296), .B(n27655), .Z(n27501) );
  AND U28274 ( .A(n27502), .B(n27501), .Z(n27713) );
  NAND U28275 ( .A(n190), .B(n27503), .Z(n27505) );
  XOR U28276 ( .A(b[19]), .B(a[182]), .Z(n27658) );
  NAND U28277 ( .A(n37821), .B(n27658), .Z(n27504) );
  NAND U28278 ( .A(n27505), .B(n27504), .Z(n27712) );
  XNOR U28279 ( .A(n27713), .B(n27712), .Z(n27714) );
  XNOR U28280 ( .A(n27715), .B(n27714), .Z(n27706) );
  NAND U28281 ( .A(n38470), .B(n27506), .Z(n27508) );
  XOR U28282 ( .A(b[31]), .B(a[170]), .Z(n27661) );
  NAND U28283 ( .A(n38453), .B(n27661), .Z(n27507) );
  AND U28284 ( .A(n27508), .B(n27507), .Z(n27673) );
  NAND U28285 ( .A(n181), .B(n27509), .Z(n27511) );
  XOR U28286 ( .A(b[3]), .B(a[198]), .Z(n27664) );
  NAND U28287 ( .A(n182), .B(n27664), .Z(n27510) );
  AND U28288 ( .A(n27511), .B(n27510), .Z(n27671) );
  NAND U28289 ( .A(n189), .B(n27512), .Z(n27514) );
  XOR U28290 ( .A(b[17]), .B(a[184]), .Z(n27667) );
  NAND U28291 ( .A(n37652), .B(n27667), .Z(n27513) );
  NAND U28292 ( .A(n27514), .B(n27513), .Z(n27670) );
  XNOR U28293 ( .A(n27671), .B(n27670), .Z(n27672) );
  XOR U28294 ( .A(n27673), .B(n27672), .Z(n27707) );
  XOR U28295 ( .A(n27706), .B(n27707), .Z(n27709) );
  XOR U28296 ( .A(n27708), .B(n27709), .Z(n27641) );
  NANDN U28297 ( .A(n27516), .B(n27515), .Z(n27520) );
  NANDN U28298 ( .A(n27518), .B(n27517), .Z(n27519) );
  AND U28299 ( .A(n27520), .B(n27519), .Z(n27694) );
  NANDN U28300 ( .A(n27522), .B(n27521), .Z(n27526) );
  NANDN U28301 ( .A(n27524), .B(n27523), .Z(n27525) );
  NAND U28302 ( .A(n27526), .B(n27525), .Z(n27695) );
  XNOR U28303 ( .A(n27694), .B(n27695), .Z(n27696) );
  NANDN U28304 ( .A(n27528), .B(n27527), .Z(n27532) );
  NANDN U28305 ( .A(n27530), .B(n27529), .Z(n27531) );
  NAND U28306 ( .A(n27532), .B(n27531), .Z(n27697) );
  XNOR U28307 ( .A(n27696), .B(n27697), .Z(n27640) );
  XNOR U28308 ( .A(n27641), .B(n27640), .Z(n27643) );
  NANDN U28309 ( .A(n27534), .B(n27533), .Z(n27538) );
  NANDN U28310 ( .A(n27536), .B(n27535), .Z(n27537) );
  AND U28311 ( .A(n27538), .B(n27537), .Z(n27642) );
  XOR U28312 ( .A(n27643), .B(n27642), .Z(n27757) );
  NANDN U28313 ( .A(n27540), .B(n27539), .Z(n27544) );
  NANDN U28314 ( .A(n27542), .B(n27541), .Z(n27543) );
  AND U28315 ( .A(n27544), .B(n27543), .Z(n27754) );
  NANDN U28316 ( .A(n27546), .B(n27545), .Z(n27550) );
  NANDN U28317 ( .A(n27548), .B(n27547), .Z(n27549) );
  AND U28318 ( .A(n27550), .B(n27549), .Z(n27637) );
  NANDN U28319 ( .A(n27552), .B(n27551), .Z(n27556) );
  OR U28320 ( .A(n27554), .B(n27553), .Z(n27555) );
  AND U28321 ( .A(n27556), .B(n27555), .Z(n27635) );
  NANDN U28322 ( .A(n27558), .B(n27557), .Z(n27562) );
  NANDN U28323 ( .A(n27560), .B(n27559), .Z(n27561) );
  AND U28324 ( .A(n27562), .B(n27561), .Z(n27701) );
  NANDN U28325 ( .A(n27564), .B(n27563), .Z(n27568) );
  NANDN U28326 ( .A(n27566), .B(n27565), .Z(n27567) );
  NAND U28327 ( .A(n27568), .B(n27567), .Z(n27700) );
  XNOR U28328 ( .A(n27701), .B(n27700), .Z(n27702) );
  NAND U28329 ( .A(b[0]), .B(a[200]), .Z(n27569) );
  XNOR U28330 ( .A(b[1]), .B(n27569), .Z(n27571) );
  NANDN U28331 ( .A(b[0]), .B(a[199]), .Z(n27570) );
  NAND U28332 ( .A(n27571), .B(n27570), .Z(n27649) );
  NAND U28333 ( .A(n194), .B(n27572), .Z(n27574) );
  XOR U28334 ( .A(b[29]), .B(a[172]), .Z(n27724) );
  NAND U28335 ( .A(n38456), .B(n27724), .Z(n27573) );
  AND U28336 ( .A(n27574), .B(n27573), .Z(n27647) );
  AND U28337 ( .A(b[31]), .B(a[168]), .Z(n27646) );
  XNOR U28338 ( .A(n27647), .B(n27646), .Z(n27648) );
  XNOR U28339 ( .A(n27649), .B(n27648), .Z(n27688) );
  NAND U28340 ( .A(n38185), .B(n27575), .Z(n27577) );
  XOR U28341 ( .A(b[23]), .B(a[178]), .Z(n27730) );
  NAND U28342 ( .A(n38132), .B(n27730), .Z(n27576) );
  AND U28343 ( .A(n27577), .B(n27576), .Z(n27721) );
  NAND U28344 ( .A(n184), .B(n27578), .Z(n27580) );
  XOR U28345 ( .A(b[7]), .B(a[194]), .Z(n27733) );
  NAND U28346 ( .A(n36592), .B(n27733), .Z(n27579) );
  AND U28347 ( .A(n27580), .B(n27579), .Z(n27719) );
  NAND U28348 ( .A(n38289), .B(n27581), .Z(n27583) );
  XOR U28349 ( .A(b[25]), .B(a[176]), .Z(n27736) );
  NAND U28350 ( .A(n38247), .B(n27736), .Z(n27582) );
  NAND U28351 ( .A(n27583), .B(n27582), .Z(n27718) );
  XNOR U28352 ( .A(n27719), .B(n27718), .Z(n27720) );
  XOR U28353 ( .A(n27721), .B(n27720), .Z(n27689) );
  XNOR U28354 ( .A(n27688), .B(n27689), .Z(n27690) );
  NAND U28355 ( .A(n187), .B(n27584), .Z(n27586) );
  XOR U28356 ( .A(b[13]), .B(a[188]), .Z(n27739) );
  NAND U28357 ( .A(n37295), .B(n27739), .Z(n27585) );
  AND U28358 ( .A(n27586), .B(n27585), .Z(n27683) );
  NAND U28359 ( .A(n186), .B(n27587), .Z(n27589) );
  XOR U28360 ( .A(b[11]), .B(a[190]), .Z(n27742) );
  NAND U28361 ( .A(n37097), .B(n27742), .Z(n27588) );
  NAND U28362 ( .A(n27589), .B(n27588), .Z(n27682) );
  XNOR U28363 ( .A(n27683), .B(n27682), .Z(n27684) );
  NAND U28364 ( .A(n188), .B(n27590), .Z(n27592) );
  XOR U28365 ( .A(b[15]), .B(a[186]), .Z(n27745) );
  NAND U28366 ( .A(n37382), .B(n27745), .Z(n27591) );
  AND U28367 ( .A(n27592), .B(n27591), .Z(n27679) );
  NAND U28368 ( .A(n38064), .B(n27593), .Z(n27595) );
  XOR U28369 ( .A(b[21]), .B(a[180]), .Z(n27748) );
  NAND U28370 ( .A(n37993), .B(n27748), .Z(n27594) );
  AND U28371 ( .A(n27595), .B(n27594), .Z(n27677) );
  NAND U28372 ( .A(n185), .B(n27596), .Z(n27598) );
  XOR U28373 ( .A(b[9]), .B(a[192]), .Z(n27751) );
  NAND U28374 ( .A(n36805), .B(n27751), .Z(n27597) );
  NAND U28375 ( .A(n27598), .B(n27597), .Z(n27676) );
  XNOR U28376 ( .A(n27677), .B(n27676), .Z(n27678) );
  XOR U28377 ( .A(n27679), .B(n27678), .Z(n27685) );
  XOR U28378 ( .A(n27684), .B(n27685), .Z(n27691) );
  XOR U28379 ( .A(n27690), .B(n27691), .Z(n27703) );
  XNOR U28380 ( .A(n27702), .B(n27703), .Z(n27634) );
  XNOR U28381 ( .A(n27635), .B(n27634), .Z(n27636) );
  XOR U28382 ( .A(n27637), .B(n27636), .Z(n27755) );
  XNOR U28383 ( .A(n27754), .B(n27755), .Z(n27756) );
  XNOR U28384 ( .A(n27757), .B(n27756), .Z(n27630) );
  XOR U28385 ( .A(n27631), .B(n27630), .Z(n27623) );
  NANDN U28386 ( .A(n27600), .B(n27599), .Z(n27604) );
  NANDN U28387 ( .A(n27602), .B(n27601), .Z(n27603) );
  AND U28388 ( .A(n27604), .B(n27603), .Z(n27622) );
  XNOR U28389 ( .A(n27623), .B(n27622), .Z(n27624) );
  NANDN U28390 ( .A(n27606), .B(n27605), .Z(n27610) );
  NAND U28391 ( .A(n27608), .B(n27607), .Z(n27609) );
  NAND U28392 ( .A(n27610), .B(n27609), .Z(n27625) );
  XNOR U28393 ( .A(n27624), .B(n27625), .Z(n27616) );
  XNOR U28394 ( .A(n27617), .B(n27616), .Z(n27618) );
  XNOR U28395 ( .A(n27619), .B(n27618), .Z(n27760) );
  XNOR U28396 ( .A(sreg[424]), .B(n27760), .Z(n27762) );
  NANDN U28397 ( .A(sreg[423]), .B(n27611), .Z(n27615) );
  NAND U28398 ( .A(n27613), .B(n27612), .Z(n27614) );
  NAND U28399 ( .A(n27615), .B(n27614), .Z(n27761) );
  XNOR U28400 ( .A(n27762), .B(n27761), .Z(c[424]) );
  NANDN U28401 ( .A(n27617), .B(n27616), .Z(n27621) );
  NANDN U28402 ( .A(n27619), .B(n27618), .Z(n27620) );
  AND U28403 ( .A(n27621), .B(n27620), .Z(n27768) );
  NANDN U28404 ( .A(n27623), .B(n27622), .Z(n27627) );
  NANDN U28405 ( .A(n27625), .B(n27624), .Z(n27626) );
  AND U28406 ( .A(n27627), .B(n27626), .Z(n27766) );
  NANDN U28407 ( .A(n27629), .B(n27628), .Z(n27633) );
  NAND U28408 ( .A(n27631), .B(n27630), .Z(n27632) );
  AND U28409 ( .A(n27633), .B(n27632), .Z(n27773) );
  NANDN U28410 ( .A(n27635), .B(n27634), .Z(n27639) );
  NANDN U28411 ( .A(n27637), .B(n27636), .Z(n27638) );
  AND U28412 ( .A(n27639), .B(n27638), .Z(n27778) );
  NANDN U28413 ( .A(n27641), .B(n27640), .Z(n27645) );
  NAND U28414 ( .A(n27643), .B(n27642), .Z(n27644) );
  AND U28415 ( .A(n27645), .B(n27644), .Z(n27777) );
  XNOR U28416 ( .A(n27778), .B(n27777), .Z(n27780) );
  NANDN U28417 ( .A(n27647), .B(n27646), .Z(n27651) );
  NANDN U28418 ( .A(n27649), .B(n27648), .Z(n27650) );
  AND U28419 ( .A(n27651), .B(n27650), .Z(n27857) );
  NAND U28420 ( .A(n38385), .B(n27652), .Z(n27654) );
  XOR U28421 ( .A(b[27]), .B(a[175]), .Z(n27801) );
  NAND U28422 ( .A(n38343), .B(n27801), .Z(n27653) );
  AND U28423 ( .A(n27654), .B(n27653), .Z(n27864) );
  NAND U28424 ( .A(n183), .B(n27655), .Z(n27657) );
  XOR U28425 ( .A(b[5]), .B(a[197]), .Z(n27804) );
  NAND U28426 ( .A(n36296), .B(n27804), .Z(n27656) );
  AND U28427 ( .A(n27657), .B(n27656), .Z(n27862) );
  NAND U28428 ( .A(n190), .B(n27658), .Z(n27660) );
  XOR U28429 ( .A(b[19]), .B(a[183]), .Z(n27807) );
  NAND U28430 ( .A(n37821), .B(n27807), .Z(n27659) );
  NAND U28431 ( .A(n27660), .B(n27659), .Z(n27861) );
  XNOR U28432 ( .A(n27862), .B(n27861), .Z(n27863) );
  XNOR U28433 ( .A(n27864), .B(n27863), .Z(n27855) );
  NAND U28434 ( .A(n38470), .B(n27661), .Z(n27663) );
  XOR U28435 ( .A(b[31]), .B(a[171]), .Z(n27810) );
  NAND U28436 ( .A(n38453), .B(n27810), .Z(n27662) );
  AND U28437 ( .A(n27663), .B(n27662), .Z(n27822) );
  NAND U28438 ( .A(n181), .B(n27664), .Z(n27666) );
  XOR U28439 ( .A(b[3]), .B(a[199]), .Z(n27813) );
  NAND U28440 ( .A(n182), .B(n27813), .Z(n27665) );
  AND U28441 ( .A(n27666), .B(n27665), .Z(n27820) );
  NAND U28442 ( .A(n189), .B(n27667), .Z(n27669) );
  XOR U28443 ( .A(b[17]), .B(a[185]), .Z(n27816) );
  NAND U28444 ( .A(n37652), .B(n27816), .Z(n27668) );
  NAND U28445 ( .A(n27669), .B(n27668), .Z(n27819) );
  XNOR U28446 ( .A(n27820), .B(n27819), .Z(n27821) );
  XOR U28447 ( .A(n27822), .B(n27821), .Z(n27856) );
  XOR U28448 ( .A(n27855), .B(n27856), .Z(n27858) );
  XOR U28449 ( .A(n27857), .B(n27858), .Z(n27790) );
  NANDN U28450 ( .A(n27671), .B(n27670), .Z(n27675) );
  NANDN U28451 ( .A(n27673), .B(n27672), .Z(n27674) );
  AND U28452 ( .A(n27675), .B(n27674), .Z(n27843) );
  NANDN U28453 ( .A(n27677), .B(n27676), .Z(n27681) );
  NANDN U28454 ( .A(n27679), .B(n27678), .Z(n27680) );
  NAND U28455 ( .A(n27681), .B(n27680), .Z(n27844) );
  XNOR U28456 ( .A(n27843), .B(n27844), .Z(n27845) );
  NANDN U28457 ( .A(n27683), .B(n27682), .Z(n27687) );
  NANDN U28458 ( .A(n27685), .B(n27684), .Z(n27686) );
  NAND U28459 ( .A(n27687), .B(n27686), .Z(n27846) );
  XNOR U28460 ( .A(n27845), .B(n27846), .Z(n27789) );
  XNOR U28461 ( .A(n27790), .B(n27789), .Z(n27792) );
  NANDN U28462 ( .A(n27689), .B(n27688), .Z(n27693) );
  NANDN U28463 ( .A(n27691), .B(n27690), .Z(n27692) );
  AND U28464 ( .A(n27693), .B(n27692), .Z(n27791) );
  XOR U28465 ( .A(n27792), .B(n27791), .Z(n27906) );
  NANDN U28466 ( .A(n27695), .B(n27694), .Z(n27699) );
  NANDN U28467 ( .A(n27697), .B(n27696), .Z(n27698) );
  AND U28468 ( .A(n27699), .B(n27698), .Z(n27903) );
  NANDN U28469 ( .A(n27701), .B(n27700), .Z(n27705) );
  NANDN U28470 ( .A(n27703), .B(n27702), .Z(n27704) );
  AND U28471 ( .A(n27705), .B(n27704), .Z(n27786) );
  NANDN U28472 ( .A(n27707), .B(n27706), .Z(n27711) );
  OR U28473 ( .A(n27709), .B(n27708), .Z(n27710) );
  AND U28474 ( .A(n27711), .B(n27710), .Z(n27784) );
  NANDN U28475 ( .A(n27713), .B(n27712), .Z(n27717) );
  NANDN U28476 ( .A(n27715), .B(n27714), .Z(n27716) );
  AND U28477 ( .A(n27717), .B(n27716), .Z(n27850) );
  NANDN U28478 ( .A(n27719), .B(n27718), .Z(n27723) );
  NANDN U28479 ( .A(n27721), .B(n27720), .Z(n27722) );
  NAND U28480 ( .A(n27723), .B(n27722), .Z(n27849) );
  XNOR U28481 ( .A(n27850), .B(n27849), .Z(n27851) );
  NAND U28482 ( .A(n194), .B(n27724), .Z(n27726) );
  XOR U28483 ( .A(b[29]), .B(a[173]), .Z(n27873) );
  NAND U28484 ( .A(n38456), .B(n27873), .Z(n27725) );
  AND U28485 ( .A(n27726), .B(n27725), .Z(n27796) );
  AND U28486 ( .A(b[31]), .B(a[169]), .Z(n27795) );
  XNOR U28487 ( .A(n27796), .B(n27795), .Z(n27797) );
  NAND U28488 ( .A(b[0]), .B(a[201]), .Z(n27727) );
  XNOR U28489 ( .A(b[1]), .B(n27727), .Z(n27729) );
  NANDN U28490 ( .A(b[0]), .B(a[200]), .Z(n27728) );
  NAND U28491 ( .A(n27729), .B(n27728), .Z(n27798) );
  XNOR U28492 ( .A(n27797), .B(n27798), .Z(n27837) );
  NAND U28493 ( .A(n38185), .B(n27730), .Z(n27732) );
  XOR U28494 ( .A(b[23]), .B(a[179]), .Z(n27879) );
  NAND U28495 ( .A(n38132), .B(n27879), .Z(n27731) );
  AND U28496 ( .A(n27732), .B(n27731), .Z(n27870) );
  NAND U28497 ( .A(n184), .B(n27733), .Z(n27735) );
  XOR U28498 ( .A(b[7]), .B(a[195]), .Z(n27882) );
  NAND U28499 ( .A(n36592), .B(n27882), .Z(n27734) );
  AND U28500 ( .A(n27735), .B(n27734), .Z(n27868) );
  NAND U28501 ( .A(n38289), .B(n27736), .Z(n27738) );
  XOR U28502 ( .A(b[25]), .B(a[177]), .Z(n27885) );
  NAND U28503 ( .A(n38247), .B(n27885), .Z(n27737) );
  NAND U28504 ( .A(n27738), .B(n27737), .Z(n27867) );
  XNOR U28505 ( .A(n27868), .B(n27867), .Z(n27869) );
  XOR U28506 ( .A(n27870), .B(n27869), .Z(n27838) );
  XNOR U28507 ( .A(n27837), .B(n27838), .Z(n27839) );
  NAND U28508 ( .A(n187), .B(n27739), .Z(n27741) );
  XOR U28509 ( .A(b[13]), .B(a[189]), .Z(n27888) );
  NAND U28510 ( .A(n37295), .B(n27888), .Z(n27740) );
  AND U28511 ( .A(n27741), .B(n27740), .Z(n27832) );
  NAND U28512 ( .A(n186), .B(n27742), .Z(n27744) );
  XOR U28513 ( .A(b[11]), .B(a[191]), .Z(n27891) );
  NAND U28514 ( .A(n37097), .B(n27891), .Z(n27743) );
  NAND U28515 ( .A(n27744), .B(n27743), .Z(n27831) );
  XNOR U28516 ( .A(n27832), .B(n27831), .Z(n27833) );
  NAND U28517 ( .A(n188), .B(n27745), .Z(n27747) );
  XOR U28518 ( .A(b[15]), .B(a[187]), .Z(n27894) );
  NAND U28519 ( .A(n37382), .B(n27894), .Z(n27746) );
  AND U28520 ( .A(n27747), .B(n27746), .Z(n27828) );
  NAND U28521 ( .A(n38064), .B(n27748), .Z(n27750) );
  XOR U28522 ( .A(b[21]), .B(a[181]), .Z(n27897) );
  NAND U28523 ( .A(n37993), .B(n27897), .Z(n27749) );
  AND U28524 ( .A(n27750), .B(n27749), .Z(n27826) );
  NAND U28525 ( .A(n185), .B(n27751), .Z(n27753) );
  XOR U28526 ( .A(b[9]), .B(a[193]), .Z(n27900) );
  NAND U28527 ( .A(n36805), .B(n27900), .Z(n27752) );
  NAND U28528 ( .A(n27753), .B(n27752), .Z(n27825) );
  XNOR U28529 ( .A(n27826), .B(n27825), .Z(n27827) );
  XOR U28530 ( .A(n27828), .B(n27827), .Z(n27834) );
  XOR U28531 ( .A(n27833), .B(n27834), .Z(n27840) );
  XOR U28532 ( .A(n27839), .B(n27840), .Z(n27852) );
  XNOR U28533 ( .A(n27851), .B(n27852), .Z(n27783) );
  XNOR U28534 ( .A(n27784), .B(n27783), .Z(n27785) );
  XOR U28535 ( .A(n27786), .B(n27785), .Z(n27904) );
  XNOR U28536 ( .A(n27903), .B(n27904), .Z(n27905) );
  XNOR U28537 ( .A(n27906), .B(n27905), .Z(n27779) );
  XOR U28538 ( .A(n27780), .B(n27779), .Z(n27772) );
  NANDN U28539 ( .A(n27755), .B(n27754), .Z(n27759) );
  NANDN U28540 ( .A(n27757), .B(n27756), .Z(n27758) );
  AND U28541 ( .A(n27759), .B(n27758), .Z(n27771) );
  XOR U28542 ( .A(n27772), .B(n27771), .Z(n27774) );
  XNOR U28543 ( .A(n27773), .B(n27774), .Z(n27765) );
  XNOR U28544 ( .A(n27766), .B(n27765), .Z(n27767) );
  XNOR U28545 ( .A(n27768), .B(n27767), .Z(n27909) );
  XNOR U28546 ( .A(sreg[425]), .B(n27909), .Z(n27911) );
  NANDN U28547 ( .A(sreg[424]), .B(n27760), .Z(n27764) );
  NAND U28548 ( .A(n27762), .B(n27761), .Z(n27763) );
  NAND U28549 ( .A(n27764), .B(n27763), .Z(n27910) );
  XNOR U28550 ( .A(n27911), .B(n27910), .Z(c[425]) );
  NANDN U28551 ( .A(n27766), .B(n27765), .Z(n27770) );
  NANDN U28552 ( .A(n27768), .B(n27767), .Z(n27769) );
  AND U28553 ( .A(n27770), .B(n27769), .Z(n27917) );
  NANDN U28554 ( .A(n27772), .B(n27771), .Z(n27776) );
  NANDN U28555 ( .A(n27774), .B(n27773), .Z(n27775) );
  AND U28556 ( .A(n27776), .B(n27775), .Z(n27915) );
  NANDN U28557 ( .A(n27778), .B(n27777), .Z(n27782) );
  NAND U28558 ( .A(n27780), .B(n27779), .Z(n27781) );
  AND U28559 ( .A(n27782), .B(n27781), .Z(n27922) );
  NANDN U28560 ( .A(n27784), .B(n27783), .Z(n27788) );
  NANDN U28561 ( .A(n27786), .B(n27785), .Z(n27787) );
  AND U28562 ( .A(n27788), .B(n27787), .Z(n27927) );
  NANDN U28563 ( .A(n27790), .B(n27789), .Z(n27794) );
  NAND U28564 ( .A(n27792), .B(n27791), .Z(n27793) );
  AND U28565 ( .A(n27794), .B(n27793), .Z(n27926) );
  XNOR U28566 ( .A(n27927), .B(n27926), .Z(n27929) );
  NANDN U28567 ( .A(n27796), .B(n27795), .Z(n27800) );
  NANDN U28568 ( .A(n27798), .B(n27797), .Z(n27799) );
  AND U28569 ( .A(n27800), .B(n27799), .Z(n28006) );
  NAND U28570 ( .A(n38385), .B(n27801), .Z(n27803) );
  XOR U28571 ( .A(b[27]), .B(a[176]), .Z(n27950) );
  NAND U28572 ( .A(n38343), .B(n27950), .Z(n27802) );
  AND U28573 ( .A(n27803), .B(n27802), .Z(n28013) );
  NAND U28574 ( .A(n183), .B(n27804), .Z(n27806) );
  XOR U28575 ( .A(b[5]), .B(a[198]), .Z(n27953) );
  NAND U28576 ( .A(n36296), .B(n27953), .Z(n27805) );
  AND U28577 ( .A(n27806), .B(n27805), .Z(n28011) );
  NAND U28578 ( .A(n190), .B(n27807), .Z(n27809) );
  XOR U28579 ( .A(b[19]), .B(a[184]), .Z(n27956) );
  NAND U28580 ( .A(n37821), .B(n27956), .Z(n27808) );
  NAND U28581 ( .A(n27809), .B(n27808), .Z(n28010) );
  XNOR U28582 ( .A(n28011), .B(n28010), .Z(n28012) );
  XNOR U28583 ( .A(n28013), .B(n28012), .Z(n28004) );
  NAND U28584 ( .A(n38470), .B(n27810), .Z(n27812) );
  XOR U28585 ( .A(b[31]), .B(a[172]), .Z(n27959) );
  NAND U28586 ( .A(n38453), .B(n27959), .Z(n27811) );
  AND U28587 ( .A(n27812), .B(n27811), .Z(n27971) );
  NAND U28588 ( .A(n181), .B(n27813), .Z(n27815) );
  XOR U28589 ( .A(b[3]), .B(a[200]), .Z(n27962) );
  NAND U28590 ( .A(n182), .B(n27962), .Z(n27814) );
  AND U28591 ( .A(n27815), .B(n27814), .Z(n27969) );
  NAND U28592 ( .A(n189), .B(n27816), .Z(n27818) );
  XOR U28593 ( .A(b[17]), .B(a[186]), .Z(n27965) );
  NAND U28594 ( .A(n37652), .B(n27965), .Z(n27817) );
  NAND U28595 ( .A(n27818), .B(n27817), .Z(n27968) );
  XNOR U28596 ( .A(n27969), .B(n27968), .Z(n27970) );
  XOR U28597 ( .A(n27971), .B(n27970), .Z(n28005) );
  XOR U28598 ( .A(n28004), .B(n28005), .Z(n28007) );
  XOR U28599 ( .A(n28006), .B(n28007), .Z(n27939) );
  NANDN U28600 ( .A(n27820), .B(n27819), .Z(n27824) );
  NANDN U28601 ( .A(n27822), .B(n27821), .Z(n27823) );
  AND U28602 ( .A(n27824), .B(n27823), .Z(n27992) );
  NANDN U28603 ( .A(n27826), .B(n27825), .Z(n27830) );
  NANDN U28604 ( .A(n27828), .B(n27827), .Z(n27829) );
  NAND U28605 ( .A(n27830), .B(n27829), .Z(n27993) );
  XNOR U28606 ( .A(n27992), .B(n27993), .Z(n27994) );
  NANDN U28607 ( .A(n27832), .B(n27831), .Z(n27836) );
  NANDN U28608 ( .A(n27834), .B(n27833), .Z(n27835) );
  NAND U28609 ( .A(n27836), .B(n27835), .Z(n27995) );
  XNOR U28610 ( .A(n27994), .B(n27995), .Z(n27938) );
  XNOR U28611 ( .A(n27939), .B(n27938), .Z(n27941) );
  NANDN U28612 ( .A(n27838), .B(n27837), .Z(n27842) );
  NANDN U28613 ( .A(n27840), .B(n27839), .Z(n27841) );
  AND U28614 ( .A(n27842), .B(n27841), .Z(n27940) );
  XOR U28615 ( .A(n27941), .B(n27940), .Z(n28055) );
  NANDN U28616 ( .A(n27844), .B(n27843), .Z(n27848) );
  NANDN U28617 ( .A(n27846), .B(n27845), .Z(n27847) );
  AND U28618 ( .A(n27848), .B(n27847), .Z(n28052) );
  NANDN U28619 ( .A(n27850), .B(n27849), .Z(n27854) );
  NANDN U28620 ( .A(n27852), .B(n27851), .Z(n27853) );
  AND U28621 ( .A(n27854), .B(n27853), .Z(n27935) );
  NANDN U28622 ( .A(n27856), .B(n27855), .Z(n27860) );
  OR U28623 ( .A(n27858), .B(n27857), .Z(n27859) );
  AND U28624 ( .A(n27860), .B(n27859), .Z(n27933) );
  NANDN U28625 ( .A(n27862), .B(n27861), .Z(n27866) );
  NANDN U28626 ( .A(n27864), .B(n27863), .Z(n27865) );
  AND U28627 ( .A(n27866), .B(n27865), .Z(n27999) );
  NANDN U28628 ( .A(n27868), .B(n27867), .Z(n27872) );
  NANDN U28629 ( .A(n27870), .B(n27869), .Z(n27871) );
  NAND U28630 ( .A(n27872), .B(n27871), .Z(n27998) );
  XNOR U28631 ( .A(n27999), .B(n27998), .Z(n28000) );
  NAND U28632 ( .A(n194), .B(n27873), .Z(n27875) );
  XOR U28633 ( .A(b[29]), .B(a[174]), .Z(n28025) );
  NAND U28634 ( .A(n38456), .B(n28025), .Z(n27874) );
  AND U28635 ( .A(n27875), .B(n27874), .Z(n27945) );
  AND U28636 ( .A(b[31]), .B(a[170]), .Z(n27944) );
  XNOR U28637 ( .A(n27945), .B(n27944), .Z(n27946) );
  NAND U28638 ( .A(b[0]), .B(a[202]), .Z(n27876) );
  XNOR U28639 ( .A(b[1]), .B(n27876), .Z(n27878) );
  NANDN U28640 ( .A(b[0]), .B(a[201]), .Z(n27877) );
  NAND U28641 ( .A(n27878), .B(n27877), .Z(n27947) );
  XNOR U28642 ( .A(n27946), .B(n27947), .Z(n27986) );
  NAND U28643 ( .A(n38185), .B(n27879), .Z(n27881) );
  XOR U28644 ( .A(b[23]), .B(a[180]), .Z(n28028) );
  NAND U28645 ( .A(n38132), .B(n28028), .Z(n27880) );
  AND U28646 ( .A(n27881), .B(n27880), .Z(n28019) );
  NAND U28647 ( .A(n184), .B(n27882), .Z(n27884) );
  XOR U28648 ( .A(b[7]), .B(a[196]), .Z(n28031) );
  NAND U28649 ( .A(n36592), .B(n28031), .Z(n27883) );
  AND U28650 ( .A(n27884), .B(n27883), .Z(n28017) );
  NAND U28651 ( .A(n38289), .B(n27885), .Z(n27887) );
  XOR U28652 ( .A(b[25]), .B(a[178]), .Z(n28034) );
  NAND U28653 ( .A(n38247), .B(n28034), .Z(n27886) );
  NAND U28654 ( .A(n27887), .B(n27886), .Z(n28016) );
  XNOR U28655 ( .A(n28017), .B(n28016), .Z(n28018) );
  XOR U28656 ( .A(n28019), .B(n28018), .Z(n27987) );
  XNOR U28657 ( .A(n27986), .B(n27987), .Z(n27988) );
  NAND U28658 ( .A(n187), .B(n27888), .Z(n27890) );
  XOR U28659 ( .A(b[13]), .B(a[190]), .Z(n28037) );
  NAND U28660 ( .A(n37295), .B(n28037), .Z(n27889) );
  AND U28661 ( .A(n27890), .B(n27889), .Z(n27981) );
  NAND U28662 ( .A(n186), .B(n27891), .Z(n27893) );
  XOR U28663 ( .A(b[11]), .B(a[192]), .Z(n28040) );
  NAND U28664 ( .A(n37097), .B(n28040), .Z(n27892) );
  NAND U28665 ( .A(n27893), .B(n27892), .Z(n27980) );
  XNOR U28666 ( .A(n27981), .B(n27980), .Z(n27982) );
  NAND U28667 ( .A(n188), .B(n27894), .Z(n27896) );
  XOR U28668 ( .A(b[15]), .B(a[188]), .Z(n28043) );
  NAND U28669 ( .A(n37382), .B(n28043), .Z(n27895) );
  AND U28670 ( .A(n27896), .B(n27895), .Z(n27977) );
  NAND U28671 ( .A(n38064), .B(n27897), .Z(n27899) );
  XOR U28672 ( .A(b[21]), .B(a[182]), .Z(n28046) );
  NAND U28673 ( .A(n37993), .B(n28046), .Z(n27898) );
  AND U28674 ( .A(n27899), .B(n27898), .Z(n27975) );
  NAND U28675 ( .A(n185), .B(n27900), .Z(n27902) );
  XOR U28676 ( .A(b[9]), .B(a[194]), .Z(n28049) );
  NAND U28677 ( .A(n36805), .B(n28049), .Z(n27901) );
  NAND U28678 ( .A(n27902), .B(n27901), .Z(n27974) );
  XNOR U28679 ( .A(n27975), .B(n27974), .Z(n27976) );
  XOR U28680 ( .A(n27977), .B(n27976), .Z(n27983) );
  XOR U28681 ( .A(n27982), .B(n27983), .Z(n27989) );
  XOR U28682 ( .A(n27988), .B(n27989), .Z(n28001) );
  XNOR U28683 ( .A(n28000), .B(n28001), .Z(n27932) );
  XNOR U28684 ( .A(n27933), .B(n27932), .Z(n27934) );
  XOR U28685 ( .A(n27935), .B(n27934), .Z(n28053) );
  XNOR U28686 ( .A(n28052), .B(n28053), .Z(n28054) );
  XNOR U28687 ( .A(n28055), .B(n28054), .Z(n27928) );
  XOR U28688 ( .A(n27929), .B(n27928), .Z(n27921) );
  NANDN U28689 ( .A(n27904), .B(n27903), .Z(n27908) );
  NANDN U28690 ( .A(n27906), .B(n27905), .Z(n27907) );
  AND U28691 ( .A(n27908), .B(n27907), .Z(n27920) );
  XOR U28692 ( .A(n27921), .B(n27920), .Z(n27923) );
  XNOR U28693 ( .A(n27922), .B(n27923), .Z(n27914) );
  XNOR U28694 ( .A(n27915), .B(n27914), .Z(n27916) );
  XNOR U28695 ( .A(n27917), .B(n27916), .Z(n28058) );
  XNOR U28696 ( .A(sreg[426]), .B(n28058), .Z(n28060) );
  NANDN U28697 ( .A(sreg[425]), .B(n27909), .Z(n27913) );
  NAND U28698 ( .A(n27911), .B(n27910), .Z(n27912) );
  NAND U28699 ( .A(n27913), .B(n27912), .Z(n28059) );
  XNOR U28700 ( .A(n28060), .B(n28059), .Z(c[426]) );
  NANDN U28701 ( .A(n27915), .B(n27914), .Z(n27919) );
  NANDN U28702 ( .A(n27917), .B(n27916), .Z(n27918) );
  AND U28703 ( .A(n27919), .B(n27918), .Z(n28066) );
  NANDN U28704 ( .A(n27921), .B(n27920), .Z(n27925) );
  NANDN U28705 ( .A(n27923), .B(n27922), .Z(n27924) );
  AND U28706 ( .A(n27925), .B(n27924), .Z(n28064) );
  NANDN U28707 ( .A(n27927), .B(n27926), .Z(n27931) );
  NAND U28708 ( .A(n27929), .B(n27928), .Z(n27930) );
  AND U28709 ( .A(n27931), .B(n27930), .Z(n28071) );
  NANDN U28710 ( .A(n27933), .B(n27932), .Z(n27937) );
  NANDN U28711 ( .A(n27935), .B(n27934), .Z(n27936) );
  AND U28712 ( .A(n27937), .B(n27936), .Z(n28076) );
  NANDN U28713 ( .A(n27939), .B(n27938), .Z(n27943) );
  NAND U28714 ( .A(n27941), .B(n27940), .Z(n27942) );
  AND U28715 ( .A(n27943), .B(n27942), .Z(n28075) );
  XNOR U28716 ( .A(n28076), .B(n28075), .Z(n28078) );
  NANDN U28717 ( .A(n27945), .B(n27944), .Z(n27949) );
  NANDN U28718 ( .A(n27947), .B(n27946), .Z(n27948) );
  AND U28719 ( .A(n27949), .B(n27948), .Z(n28155) );
  NAND U28720 ( .A(n38385), .B(n27950), .Z(n27952) );
  XOR U28721 ( .A(b[27]), .B(a[177]), .Z(n28099) );
  NAND U28722 ( .A(n38343), .B(n28099), .Z(n27951) );
  AND U28723 ( .A(n27952), .B(n27951), .Z(n28162) );
  NAND U28724 ( .A(n183), .B(n27953), .Z(n27955) );
  XOR U28725 ( .A(b[5]), .B(a[199]), .Z(n28102) );
  NAND U28726 ( .A(n36296), .B(n28102), .Z(n27954) );
  AND U28727 ( .A(n27955), .B(n27954), .Z(n28160) );
  NAND U28728 ( .A(n190), .B(n27956), .Z(n27958) );
  XOR U28729 ( .A(b[19]), .B(a[185]), .Z(n28105) );
  NAND U28730 ( .A(n37821), .B(n28105), .Z(n27957) );
  NAND U28731 ( .A(n27958), .B(n27957), .Z(n28159) );
  XNOR U28732 ( .A(n28160), .B(n28159), .Z(n28161) );
  XNOR U28733 ( .A(n28162), .B(n28161), .Z(n28153) );
  NAND U28734 ( .A(n38470), .B(n27959), .Z(n27961) );
  XOR U28735 ( .A(b[31]), .B(a[173]), .Z(n28108) );
  NAND U28736 ( .A(n38453), .B(n28108), .Z(n27960) );
  AND U28737 ( .A(n27961), .B(n27960), .Z(n28120) );
  NAND U28738 ( .A(n181), .B(n27962), .Z(n27964) );
  XOR U28739 ( .A(b[3]), .B(a[201]), .Z(n28111) );
  NAND U28740 ( .A(n182), .B(n28111), .Z(n27963) );
  AND U28741 ( .A(n27964), .B(n27963), .Z(n28118) );
  NAND U28742 ( .A(n189), .B(n27965), .Z(n27967) );
  XOR U28743 ( .A(b[17]), .B(a[187]), .Z(n28114) );
  NAND U28744 ( .A(n37652), .B(n28114), .Z(n27966) );
  NAND U28745 ( .A(n27967), .B(n27966), .Z(n28117) );
  XNOR U28746 ( .A(n28118), .B(n28117), .Z(n28119) );
  XOR U28747 ( .A(n28120), .B(n28119), .Z(n28154) );
  XOR U28748 ( .A(n28153), .B(n28154), .Z(n28156) );
  XOR U28749 ( .A(n28155), .B(n28156), .Z(n28088) );
  NANDN U28750 ( .A(n27969), .B(n27968), .Z(n27973) );
  NANDN U28751 ( .A(n27971), .B(n27970), .Z(n27972) );
  AND U28752 ( .A(n27973), .B(n27972), .Z(n28141) );
  NANDN U28753 ( .A(n27975), .B(n27974), .Z(n27979) );
  NANDN U28754 ( .A(n27977), .B(n27976), .Z(n27978) );
  NAND U28755 ( .A(n27979), .B(n27978), .Z(n28142) );
  XNOR U28756 ( .A(n28141), .B(n28142), .Z(n28143) );
  NANDN U28757 ( .A(n27981), .B(n27980), .Z(n27985) );
  NANDN U28758 ( .A(n27983), .B(n27982), .Z(n27984) );
  NAND U28759 ( .A(n27985), .B(n27984), .Z(n28144) );
  XNOR U28760 ( .A(n28143), .B(n28144), .Z(n28087) );
  XNOR U28761 ( .A(n28088), .B(n28087), .Z(n28090) );
  NANDN U28762 ( .A(n27987), .B(n27986), .Z(n27991) );
  NANDN U28763 ( .A(n27989), .B(n27988), .Z(n27990) );
  AND U28764 ( .A(n27991), .B(n27990), .Z(n28089) );
  XOR U28765 ( .A(n28090), .B(n28089), .Z(n28204) );
  NANDN U28766 ( .A(n27993), .B(n27992), .Z(n27997) );
  NANDN U28767 ( .A(n27995), .B(n27994), .Z(n27996) );
  AND U28768 ( .A(n27997), .B(n27996), .Z(n28201) );
  NANDN U28769 ( .A(n27999), .B(n27998), .Z(n28003) );
  NANDN U28770 ( .A(n28001), .B(n28000), .Z(n28002) );
  AND U28771 ( .A(n28003), .B(n28002), .Z(n28084) );
  NANDN U28772 ( .A(n28005), .B(n28004), .Z(n28009) );
  OR U28773 ( .A(n28007), .B(n28006), .Z(n28008) );
  AND U28774 ( .A(n28009), .B(n28008), .Z(n28082) );
  NANDN U28775 ( .A(n28011), .B(n28010), .Z(n28015) );
  NANDN U28776 ( .A(n28013), .B(n28012), .Z(n28014) );
  AND U28777 ( .A(n28015), .B(n28014), .Z(n28148) );
  NANDN U28778 ( .A(n28017), .B(n28016), .Z(n28021) );
  NANDN U28779 ( .A(n28019), .B(n28018), .Z(n28020) );
  NAND U28780 ( .A(n28021), .B(n28020), .Z(n28147) );
  XNOR U28781 ( .A(n28148), .B(n28147), .Z(n28149) );
  NAND U28782 ( .A(b[0]), .B(a[203]), .Z(n28022) );
  XNOR U28783 ( .A(b[1]), .B(n28022), .Z(n28024) );
  NANDN U28784 ( .A(b[0]), .B(a[202]), .Z(n28023) );
  NAND U28785 ( .A(n28024), .B(n28023), .Z(n28096) );
  NAND U28786 ( .A(n194), .B(n28025), .Z(n28027) );
  XOR U28787 ( .A(b[29]), .B(a[175]), .Z(n28174) );
  NAND U28788 ( .A(n38456), .B(n28174), .Z(n28026) );
  AND U28789 ( .A(n28027), .B(n28026), .Z(n28094) );
  AND U28790 ( .A(b[31]), .B(a[171]), .Z(n28093) );
  XNOR U28791 ( .A(n28094), .B(n28093), .Z(n28095) );
  XNOR U28792 ( .A(n28096), .B(n28095), .Z(n28135) );
  NAND U28793 ( .A(n38185), .B(n28028), .Z(n28030) );
  XOR U28794 ( .A(b[23]), .B(a[181]), .Z(n28177) );
  NAND U28795 ( .A(n38132), .B(n28177), .Z(n28029) );
  AND U28796 ( .A(n28030), .B(n28029), .Z(n28168) );
  NAND U28797 ( .A(n184), .B(n28031), .Z(n28033) );
  XOR U28798 ( .A(b[7]), .B(a[197]), .Z(n28180) );
  NAND U28799 ( .A(n36592), .B(n28180), .Z(n28032) );
  AND U28800 ( .A(n28033), .B(n28032), .Z(n28166) );
  NAND U28801 ( .A(n38289), .B(n28034), .Z(n28036) );
  XOR U28802 ( .A(b[25]), .B(a[179]), .Z(n28183) );
  NAND U28803 ( .A(n38247), .B(n28183), .Z(n28035) );
  NAND U28804 ( .A(n28036), .B(n28035), .Z(n28165) );
  XNOR U28805 ( .A(n28166), .B(n28165), .Z(n28167) );
  XOR U28806 ( .A(n28168), .B(n28167), .Z(n28136) );
  XNOR U28807 ( .A(n28135), .B(n28136), .Z(n28137) );
  NAND U28808 ( .A(n187), .B(n28037), .Z(n28039) );
  XOR U28809 ( .A(b[13]), .B(a[191]), .Z(n28186) );
  NAND U28810 ( .A(n37295), .B(n28186), .Z(n28038) );
  AND U28811 ( .A(n28039), .B(n28038), .Z(n28130) );
  NAND U28812 ( .A(n186), .B(n28040), .Z(n28042) );
  XOR U28813 ( .A(b[11]), .B(a[193]), .Z(n28189) );
  NAND U28814 ( .A(n37097), .B(n28189), .Z(n28041) );
  NAND U28815 ( .A(n28042), .B(n28041), .Z(n28129) );
  XNOR U28816 ( .A(n28130), .B(n28129), .Z(n28131) );
  NAND U28817 ( .A(n188), .B(n28043), .Z(n28045) );
  XOR U28818 ( .A(b[15]), .B(a[189]), .Z(n28192) );
  NAND U28819 ( .A(n37382), .B(n28192), .Z(n28044) );
  AND U28820 ( .A(n28045), .B(n28044), .Z(n28126) );
  NAND U28821 ( .A(n38064), .B(n28046), .Z(n28048) );
  XOR U28822 ( .A(b[21]), .B(a[183]), .Z(n28195) );
  NAND U28823 ( .A(n37993), .B(n28195), .Z(n28047) );
  AND U28824 ( .A(n28048), .B(n28047), .Z(n28124) );
  NAND U28825 ( .A(n185), .B(n28049), .Z(n28051) );
  XOR U28826 ( .A(b[9]), .B(a[195]), .Z(n28198) );
  NAND U28827 ( .A(n36805), .B(n28198), .Z(n28050) );
  NAND U28828 ( .A(n28051), .B(n28050), .Z(n28123) );
  XNOR U28829 ( .A(n28124), .B(n28123), .Z(n28125) );
  XOR U28830 ( .A(n28126), .B(n28125), .Z(n28132) );
  XOR U28831 ( .A(n28131), .B(n28132), .Z(n28138) );
  XOR U28832 ( .A(n28137), .B(n28138), .Z(n28150) );
  XNOR U28833 ( .A(n28149), .B(n28150), .Z(n28081) );
  XNOR U28834 ( .A(n28082), .B(n28081), .Z(n28083) );
  XOR U28835 ( .A(n28084), .B(n28083), .Z(n28202) );
  XNOR U28836 ( .A(n28201), .B(n28202), .Z(n28203) );
  XNOR U28837 ( .A(n28204), .B(n28203), .Z(n28077) );
  XOR U28838 ( .A(n28078), .B(n28077), .Z(n28070) );
  NANDN U28839 ( .A(n28053), .B(n28052), .Z(n28057) );
  NANDN U28840 ( .A(n28055), .B(n28054), .Z(n28056) );
  AND U28841 ( .A(n28057), .B(n28056), .Z(n28069) );
  XOR U28842 ( .A(n28070), .B(n28069), .Z(n28072) );
  XNOR U28843 ( .A(n28071), .B(n28072), .Z(n28063) );
  XNOR U28844 ( .A(n28064), .B(n28063), .Z(n28065) );
  XNOR U28845 ( .A(n28066), .B(n28065), .Z(n28207) );
  XNOR U28846 ( .A(sreg[427]), .B(n28207), .Z(n28209) );
  NANDN U28847 ( .A(sreg[426]), .B(n28058), .Z(n28062) );
  NAND U28848 ( .A(n28060), .B(n28059), .Z(n28061) );
  NAND U28849 ( .A(n28062), .B(n28061), .Z(n28208) );
  XNOR U28850 ( .A(n28209), .B(n28208), .Z(c[427]) );
  NANDN U28851 ( .A(n28064), .B(n28063), .Z(n28068) );
  NANDN U28852 ( .A(n28066), .B(n28065), .Z(n28067) );
  AND U28853 ( .A(n28068), .B(n28067), .Z(n28215) );
  NANDN U28854 ( .A(n28070), .B(n28069), .Z(n28074) );
  NANDN U28855 ( .A(n28072), .B(n28071), .Z(n28073) );
  AND U28856 ( .A(n28074), .B(n28073), .Z(n28213) );
  NANDN U28857 ( .A(n28076), .B(n28075), .Z(n28080) );
  NAND U28858 ( .A(n28078), .B(n28077), .Z(n28079) );
  AND U28859 ( .A(n28080), .B(n28079), .Z(n28220) );
  NANDN U28860 ( .A(n28082), .B(n28081), .Z(n28086) );
  NANDN U28861 ( .A(n28084), .B(n28083), .Z(n28085) );
  AND U28862 ( .A(n28086), .B(n28085), .Z(n28351) );
  NANDN U28863 ( .A(n28088), .B(n28087), .Z(n28092) );
  NAND U28864 ( .A(n28090), .B(n28089), .Z(n28091) );
  AND U28865 ( .A(n28092), .B(n28091), .Z(n28350) );
  XNOR U28866 ( .A(n28351), .B(n28350), .Z(n28353) );
  NANDN U28867 ( .A(n28094), .B(n28093), .Z(n28098) );
  NANDN U28868 ( .A(n28096), .B(n28095), .Z(n28097) );
  AND U28869 ( .A(n28098), .B(n28097), .Z(n28298) );
  NAND U28870 ( .A(n38385), .B(n28099), .Z(n28101) );
  XOR U28871 ( .A(b[27]), .B(a[178]), .Z(n28242) );
  NAND U28872 ( .A(n38343), .B(n28242), .Z(n28100) );
  AND U28873 ( .A(n28101), .B(n28100), .Z(n28305) );
  NAND U28874 ( .A(n183), .B(n28102), .Z(n28104) );
  XOR U28875 ( .A(b[5]), .B(a[200]), .Z(n28245) );
  NAND U28876 ( .A(n36296), .B(n28245), .Z(n28103) );
  AND U28877 ( .A(n28104), .B(n28103), .Z(n28303) );
  NAND U28878 ( .A(n190), .B(n28105), .Z(n28107) );
  XOR U28879 ( .A(b[19]), .B(a[186]), .Z(n28248) );
  NAND U28880 ( .A(n37821), .B(n28248), .Z(n28106) );
  NAND U28881 ( .A(n28107), .B(n28106), .Z(n28302) );
  XNOR U28882 ( .A(n28303), .B(n28302), .Z(n28304) );
  XNOR U28883 ( .A(n28305), .B(n28304), .Z(n28296) );
  NAND U28884 ( .A(n38470), .B(n28108), .Z(n28110) );
  XOR U28885 ( .A(b[31]), .B(a[174]), .Z(n28251) );
  NAND U28886 ( .A(n38453), .B(n28251), .Z(n28109) );
  AND U28887 ( .A(n28110), .B(n28109), .Z(n28263) );
  NAND U28888 ( .A(n181), .B(n28111), .Z(n28113) );
  XOR U28889 ( .A(b[3]), .B(a[202]), .Z(n28254) );
  NAND U28890 ( .A(n182), .B(n28254), .Z(n28112) );
  AND U28891 ( .A(n28113), .B(n28112), .Z(n28261) );
  NAND U28892 ( .A(n189), .B(n28114), .Z(n28116) );
  XOR U28893 ( .A(b[17]), .B(a[188]), .Z(n28257) );
  NAND U28894 ( .A(n37652), .B(n28257), .Z(n28115) );
  NAND U28895 ( .A(n28116), .B(n28115), .Z(n28260) );
  XNOR U28896 ( .A(n28261), .B(n28260), .Z(n28262) );
  XOR U28897 ( .A(n28263), .B(n28262), .Z(n28297) );
  XOR U28898 ( .A(n28296), .B(n28297), .Z(n28299) );
  XOR U28899 ( .A(n28298), .B(n28299), .Z(n28231) );
  NANDN U28900 ( .A(n28118), .B(n28117), .Z(n28122) );
  NANDN U28901 ( .A(n28120), .B(n28119), .Z(n28121) );
  AND U28902 ( .A(n28122), .B(n28121), .Z(n28284) );
  NANDN U28903 ( .A(n28124), .B(n28123), .Z(n28128) );
  NANDN U28904 ( .A(n28126), .B(n28125), .Z(n28127) );
  NAND U28905 ( .A(n28128), .B(n28127), .Z(n28285) );
  XNOR U28906 ( .A(n28284), .B(n28285), .Z(n28286) );
  NANDN U28907 ( .A(n28130), .B(n28129), .Z(n28134) );
  NANDN U28908 ( .A(n28132), .B(n28131), .Z(n28133) );
  NAND U28909 ( .A(n28134), .B(n28133), .Z(n28287) );
  XNOR U28910 ( .A(n28286), .B(n28287), .Z(n28230) );
  XNOR U28911 ( .A(n28231), .B(n28230), .Z(n28233) );
  NANDN U28912 ( .A(n28136), .B(n28135), .Z(n28140) );
  NANDN U28913 ( .A(n28138), .B(n28137), .Z(n28139) );
  AND U28914 ( .A(n28140), .B(n28139), .Z(n28232) );
  XOR U28915 ( .A(n28233), .B(n28232), .Z(n28347) );
  NANDN U28916 ( .A(n28142), .B(n28141), .Z(n28146) );
  NANDN U28917 ( .A(n28144), .B(n28143), .Z(n28145) );
  AND U28918 ( .A(n28146), .B(n28145), .Z(n28344) );
  NANDN U28919 ( .A(n28148), .B(n28147), .Z(n28152) );
  NANDN U28920 ( .A(n28150), .B(n28149), .Z(n28151) );
  AND U28921 ( .A(n28152), .B(n28151), .Z(n28227) );
  NANDN U28922 ( .A(n28154), .B(n28153), .Z(n28158) );
  OR U28923 ( .A(n28156), .B(n28155), .Z(n28157) );
  AND U28924 ( .A(n28158), .B(n28157), .Z(n28225) );
  NANDN U28925 ( .A(n28160), .B(n28159), .Z(n28164) );
  NANDN U28926 ( .A(n28162), .B(n28161), .Z(n28163) );
  AND U28927 ( .A(n28164), .B(n28163), .Z(n28291) );
  NANDN U28928 ( .A(n28166), .B(n28165), .Z(n28170) );
  NANDN U28929 ( .A(n28168), .B(n28167), .Z(n28169) );
  NAND U28930 ( .A(n28170), .B(n28169), .Z(n28290) );
  XNOR U28931 ( .A(n28291), .B(n28290), .Z(n28292) );
  NAND U28932 ( .A(b[0]), .B(a[204]), .Z(n28171) );
  XNOR U28933 ( .A(b[1]), .B(n28171), .Z(n28173) );
  NANDN U28934 ( .A(b[0]), .B(a[203]), .Z(n28172) );
  NAND U28935 ( .A(n28173), .B(n28172), .Z(n28239) );
  NAND U28936 ( .A(n194), .B(n28174), .Z(n28176) );
  XOR U28937 ( .A(b[29]), .B(a[176]), .Z(n28317) );
  NAND U28938 ( .A(n38456), .B(n28317), .Z(n28175) );
  AND U28939 ( .A(n28176), .B(n28175), .Z(n28237) );
  AND U28940 ( .A(b[31]), .B(a[172]), .Z(n28236) );
  XNOR U28941 ( .A(n28237), .B(n28236), .Z(n28238) );
  XNOR U28942 ( .A(n28239), .B(n28238), .Z(n28278) );
  NAND U28943 ( .A(n38185), .B(n28177), .Z(n28179) );
  XOR U28944 ( .A(b[23]), .B(a[182]), .Z(n28320) );
  NAND U28945 ( .A(n38132), .B(n28320), .Z(n28178) );
  AND U28946 ( .A(n28179), .B(n28178), .Z(n28311) );
  NAND U28947 ( .A(n184), .B(n28180), .Z(n28182) );
  XOR U28948 ( .A(b[7]), .B(a[198]), .Z(n28323) );
  NAND U28949 ( .A(n36592), .B(n28323), .Z(n28181) );
  AND U28950 ( .A(n28182), .B(n28181), .Z(n28309) );
  NAND U28951 ( .A(n38289), .B(n28183), .Z(n28185) );
  XOR U28952 ( .A(b[25]), .B(a[180]), .Z(n28326) );
  NAND U28953 ( .A(n38247), .B(n28326), .Z(n28184) );
  NAND U28954 ( .A(n28185), .B(n28184), .Z(n28308) );
  XNOR U28955 ( .A(n28309), .B(n28308), .Z(n28310) );
  XOR U28956 ( .A(n28311), .B(n28310), .Z(n28279) );
  XNOR U28957 ( .A(n28278), .B(n28279), .Z(n28280) );
  NAND U28958 ( .A(n187), .B(n28186), .Z(n28188) );
  XOR U28959 ( .A(b[13]), .B(a[192]), .Z(n28329) );
  NAND U28960 ( .A(n37295), .B(n28329), .Z(n28187) );
  AND U28961 ( .A(n28188), .B(n28187), .Z(n28273) );
  NAND U28962 ( .A(n186), .B(n28189), .Z(n28191) );
  XOR U28963 ( .A(b[11]), .B(a[194]), .Z(n28332) );
  NAND U28964 ( .A(n37097), .B(n28332), .Z(n28190) );
  NAND U28965 ( .A(n28191), .B(n28190), .Z(n28272) );
  XNOR U28966 ( .A(n28273), .B(n28272), .Z(n28274) );
  NAND U28967 ( .A(n188), .B(n28192), .Z(n28194) );
  XOR U28968 ( .A(b[15]), .B(a[190]), .Z(n28335) );
  NAND U28969 ( .A(n37382), .B(n28335), .Z(n28193) );
  AND U28970 ( .A(n28194), .B(n28193), .Z(n28269) );
  NAND U28971 ( .A(n38064), .B(n28195), .Z(n28197) );
  XOR U28972 ( .A(b[21]), .B(a[184]), .Z(n28338) );
  NAND U28973 ( .A(n37993), .B(n28338), .Z(n28196) );
  AND U28974 ( .A(n28197), .B(n28196), .Z(n28267) );
  NAND U28975 ( .A(n185), .B(n28198), .Z(n28200) );
  XOR U28976 ( .A(b[9]), .B(a[196]), .Z(n28341) );
  NAND U28977 ( .A(n36805), .B(n28341), .Z(n28199) );
  NAND U28978 ( .A(n28200), .B(n28199), .Z(n28266) );
  XNOR U28979 ( .A(n28267), .B(n28266), .Z(n28268) );
  XOR U28980 ( .A(n28269), .B(n28268), .Z(n28275) );
  XOR U28981 ( .A(n28274), .B(n28275), .Z(n28281) );
  XOR U28982 ( .A(n28280), .B(n28281), .Z(n28293) );
  XNOR U28983 ( .A(n28292), .B(n28293), .Z(n28224) );
  XNOR U28984 ( .A(n28225), .B(n28224), .Z(n28226) );
  XOR U28985 ( .A(n28227), .B(n28226), .Z(n28345) );
  XNOR U28986 ( .A(n28344), .B(n28345), .Z(n28346) );
  XNOR U28987 ( .A(n28347), .B(n28346), .Z(n28352) );
  XOR U28988 ( .A(n28353), .B(n28352), .Z(n28219) );
  NANDN U28989 ( .A(n28202), .B(n28201), .Z(n28206) );
  NANDN U28990 ( .A(n28204), .B(n28203), .Z(n28205) );
  AND U28991 ( .A(n28206), .B(n28205), .Z(n28218) );
  XOR U28992 ( .A(n28219), .B(n28218), .Z(n28221) );
  XNOR U28993 ( .A(n28220), .B(n28221), .Z(n28212) );
  XNOR U28994 ( .A(n28213), .B(n28212), .Z(n28214) );
  XNOR U28995 ( .A(n28215), .B(n28214), .Z(n28356) );
  XNOR U28996 ( .A(sreg[428]), .B(n28356), .Z(n28358) );
  NANDN U28997 ( .A(sreg[427]), .B(n28207), .Z(n28211) );
  NAND U28998 ( .A(n28209), .B(n28208), .Z(n28210) );
  NAND U28999 ( .A(n28211), .B(n28210), .Z(n28357) );
  XNOR U29000 ( .A(n28358), .B(n28357), .Z(c[428]) );
  NANDN U29001 ( .A(n28213), .B(n28212), .Z(n28217) );
  NANDN U29002 ( .A(n28215), .B(n28214), .Z(n28216) );
  AND U29003 ( .A(n28217), .B(n28216), .Z(n28364) );
  NANDN U29004 ( .A(n28219), .B(n28218), .Z(n28223) );
  NANDN U29005 ( .A(n28221), .B(n28220), .Z(n28222) );
  AND U29006 ( .A(n28223), .B(n28222), .Z(n28362) );
  NANDN U29007 ( .A(n28225), .B(n28224), .Z(n28229) );
  NANDN U29008 ( .A(n28227), .B(n28226), .Z(n28228) );
  AND U29009 ( .A(n28229), .B(n28228), .Z(n28500) );
  NANDN U29010 ( .A(n28231), .B(n28230), .Z(n28235) );
  NAND U29011 ( .A(n28233), .B(n28232), .Z(n28234) );
  AND U29012 ( .A(n28235), .B(n28234), .Z(n28499) );
  XNOR U29013 ( .A(n28500), .B(n28499), .Z(n28502) );
  NANDN U29014 ( .A(n28237), .B(n28236), .Z(n28241) );
  NANDN U29015 ( .A(n28239), .B(n28238), .Z(n28240) );
  AND U29016 ( .A(n28241), .B(n28240), .Z(n28447) );
  NAND U29017 ( .A(n38385), .B(n28242), .Z(n28244) );
  XOR U29018 ( .A(b[27]), .B(a[179]), .Z(n28391) );
  NAND U29019 ( .A(n38343), .B(n28391), .Z(n28243) );
  AND U29020 ( .A(n28244), .B(n28243), .Z(n28454) );
  NAND U29021 ( .A(n183), .B(n28245), .Z(n28247) );
  XOR U29022 ( .A(b[5]), .B(a[201]), .Z(n28394) );
  NAND U29023 ( .A(n36296), .B(n28394), .Z(n28246) );
  AND U29024 ( .A(n28247), .B(n28246), .Z(n28452) );
  NAND U29025 ( .A(n190), .B(n28248), .Z(n28250) );
  XOR U29026 ( .A(b[19]), .B(a[187]), .Z(n28397) );
  NAND U29027 ( .A(n37821), .B(n28397), .Z(n28249) );
  NAND U29028 ( .A(n28250), .B(n28249), .Z(n28451) );
  XNOR U29029 ( .A(n28452), .B(n28451), .Z(n28453) );
  XNOR U29030 ( .A(n28454), .B(n28453), .Z(n28445) );
  NAND U29031 ( .A(n38470), .B(n28251), .Z(n28253) );
  XOR U29032 ( .A(b[31]), .B(a[175]), .Z(n28400) );
  NAND U29033 ( .A(n38453), .B(n28400), .Z(n28252) );
  AND U29034 ( .A(n28253), .B(n28252), .Z(n28412) );
  NAND U29035 ( .A(n181), .B(n28254), .Z(n28256) );
  XOR U29036 ( .A(b[3]), .B(a[203]), .Z(n28403) );
  NAND U29037 ( .A(n182), .B(n28403), .Z(n28255) );
  AND U29038 ( .A(n28256), .B(n28255), .Z(n28410) );
  NAND U29039 ( .A(n189), .B(n28257), .Z(n28259) );
  XOR U29040 ( .A(b[17]), .B(a[189]), .Z(n28406) );
  NAND U29041 ( .A(n37652), .B(n28406), .Z(n28258) );
  NAND U29042 ( .A(n28259), .B(n28258), .Z(n28409) );
  XNOR U29043 ( .A(n28410), .B(n28409), .Z(n28411) );
  XOR U29044 ( .A(n28412), .B(n28411), .Z(n28446) );
  XOR U29045 ( .A(n28445), .B(n28446), .Z(n28448) );
  XOR U29046 ( .A(n28447), .B(n28448), .Z(n28380) );
  NANDN U29047 ( .A(n28261), .B(n28260), .Z(n28265) );
  NANDN U29048 ( .A(n28263), .B(n28262), .Z(n28264) );
  AND U29049 ( .A(n28265), .B(n28264), .Z(n28433) );
  NANDN U29050 ( .A(n28267), .B(n28266), .Z(n28271) );
  NANDN U29051 ( .A(n28269), .B(n28268), .Z(n28270) );
  NAND U29052 ( .A(n28271), .B(n28270), .Z(n28434) );
  XNOR U29053 ( .A(n28433), .B(n28434), .Z(n28435) );
  NANDN U29054 ( .A(n28273), .B(n28272), .Z(n28277) );
  NANDN U29055 ( .A(n28275), .B(n28274), .Z(n28276) );
  NAND U29056 ( .A(n28277), .B(n28276), .Z(n28436) );
  XNOR U29057 ( .A(n28435), .B(n28436), .Z(n28379) );
  XNOR U29058 ( .A(n28380), .B(n28379), .Z(n28382) );
  NANDN U29059 ( .A(n28279), .B(n28278), .Z(n28283) );
  NANDN U29060 ( .A(n28281), .B(n28280), .Z(n28282) );
  AND U29061 ( .A(n28283), .B(n28282), .Z(n28381) );
  XOR U29062 ( .A(n28382), .B(n28381), .Z(n28496) );
  NANDN U29063 ( .A(n28285), .B(n28284), .Z(n28289) );
  NANDN U29064 ( .A(n28287), .B(n28286), .Z(n28288) );
  AND U29065 ( .A(n28289), .B(n28288), .Z(n28493) );
  NANDN U29066 ( .A(n28291), .B(n28290), .Z(n28295) );
  NANDN U29067 ( .A(n28293), .B(n28292), .Z(n28294) );
  AND U29068 ( .A(n28295), .B(n28294), .Z(n28376) );
  NANDN U29069 ( .A(n28297), .B(n28296), .Z(n28301) );
  OR U29070 ( .A(n28299), .B(n28298), .Z(n28300) );
  AND U29071 ( .A(n28301), .B(n28300), .Z(n28374) );
  NANDN U29072 ( .A(n28303), .B(n28302), .Z(n28307) );
  NANDN U29073 ( .A(n28305), .B(n28304), .Z(n28306) );
  AND U29074 ( .A(n28307), .B(n28306), .Z(n28440) );
  NANDN U29075 ( .A(n28309), .B(n28308), .Z(n28313) );
  NANDN U29076 ( .A(n28311), .B(n28310), .Z(n28312) );
  NAND U29077 ( .A(n28313), .B(n28312), .Z(n28439) );
  XNOR U29078 ( .A(n28440), .B(n28439), .Z(n28441) );
  NAND U29079 ( .A(b[0]), .B(a[205]), .Z(n28314) );
  XNOR U29080 ( .A(b[1]), .B(n28314), .Z(n28316) );
  NANDN U29081 ( .A(b[0]), .B(a[204]), .Z(n28315) );
  NAND U29082 ( .A(n28316), .B(n28315), .Z(n28388) );
  NAND U29083 ( .A(n194), .B(n28317), .Z(n28319) );
  XOR U29084 ( .A(b[29]), .B(a[177]), .Z(n28466) );
  NAND U29085 ( .A(n38456), .B(n28466), .Z(n28318) );
  AND U29086 ( .A(n28319), .B(n28318), .Z(n28386) );
  AND U29087 ( .A(b[31]), .B(a[173]), .Z(n28385) );
  XNOR U29088 ( .A(n28386), .B(n28385), .Z(n28387) );
  XNOR U29089 ( .A(n28388), .B(n28387), .Z(n28427) );
  NAND U29090 ( .A(n38185), .B(n28320), .Z(n28322) );
  XOR U29091 ( .A(b[23]), .B(a[183]), .Z(n28469) );
  NAND U29092 ( .A(n38132), .B(n28469), .Z(n28321) );
  AND U29093 ( .A(n28322), .B(n28321), .Z(n28460) );
  NAND U29094 ( .A(n184), .B(n28323), .Z(n28325) );
  XOR U29095 ( .A(b[7]), .B(a[199]), .Z(n28472) );
  NAND U29096 ( .A(n36592), .B(n28472), .Z(n28324) );
  AND U29097 ( .A(n28325), .B(n28324), .Z(n28458) );
  NAND U29098 ( .A(n38289), .B(n28326), .Z(n28328) );
  XOR U29099 ( .A(b[25]), .B(a[181]), .Z(n28475) );
  NAND U29100 ( .A(n38247), .B(n28475), .Z(n28327) );
  NAND U29101 ( .A(n28328), .B(n28327), .Z(n28457) );
  XNOR U29102 ( .A(n28458), .B(n28457), .Z(n28459) );
  XOR U29103 ( .A(n28460), .B(n28459), .Z(n28428) );
  XNOR U29104 ( .A(n28427), .B(n28428), .Z(n28429) );
  NAND U29105 ( .A(n187), .B(n28329), .Z(n28331) );
  XOR U29106 ( .A(b[13]), .B(a[193]), .Z(n28478) );
  NAND U29107 ( .A(n37295), .B(n28478), .Z(n28330) );
  AND U29108 ( .A(n28331), .B(n28330), .Z(n28422) );
  NAND U29109 ( .A(n186), .B(n28332), .Z(n28334) );
  XOR U29110 ( .A(b[11]), .B(a[195]), .Z(n28481) );
  NAND U29111 ( .A(n37097), .B(n28481), .Z(n28333) );
  NAND U29112 ( .A(n28334), .B(n28333), .Z(n28421) );
  XNOR U29113 ( .A(n28422), .B(n28421), .Z(n28423) );
  NAND U29114 ( .A(n188), .B(n28335), .Z(n28337) );
  XOR U29115 ( .A(b[15]), .B(a[191]), .Z(n28484) );
  NAND U29116 ( .A(n37382), .B(n28484), .Z(n28336) );
  AND U29117 ( .A(n28337), .B(n28336), .Z(n28418) );
  NAND U29118 ( .A(n38064), .B(n28338), .Z(n28340) );
  XOR U29119 ( .A(b[21]), .B(a[185]), .Z(n28487) );
  NAND U29120 ( .A(n37993), .B(n28487), .Z(n28339) );
  AND U29121 ( .A(n28340), .B(n28339), .Z(n28416) );
  NAND U29122 ( .A(n185), .B(n28341), .Z(n28343) );
  XOR U29123 ( .A(b[9]), .B(a[197]), .Z(n28490) );
  NAND U29124 ( .A(n36805), .B(n28490), .Z(n28342) );
  NAND U29125 ( .A(n28343), .B(n28342), .Z(n28415) );
  XNOR U29126 ( .A(n28416), .B(n28415), .Z(n28417) );
  XOR U29127 ( .A(n28418), .B(n28417), .Z(n28424) );
  XOR U29128 ( .A(n28423), .B(n28424), .Z(n28430) );
  XOR U29129 ( .A(n28429), .B(n28430), .Z(n28442) );
  XNOR U29130 ( .A(n28441), .B(n28442), .Z(n28373) );
  XNOR U29131 ( .A(n28374), .B(n28373), .Z(n28375) );
  XOR U29132 ( .A(n28376), .B(n28375), .Z(n28494) );
  XNOR U29133 ( .A(n28493), .B(n28494), .Z(n28495) );
  XNOR U29134 ( .A(n28496), .B(n28495), .Z(n28501) );
  XOR U29135 ( .A(n28502), .B(n28501), .Z(n28368) );
  NANDN U29136 ( .A(n28345), .B(n28344), .Z(n28349) );
  NANDN U29137 ( .A(n28347), .B(n28346), .Z(n28348) );
  AND U29138 ( .A(n28349), .B(n28348), .Z(n28367) );
  XNOR U29139 ( .A(n28368), .B(n28367), .Z(n28369) );
  NANDN U29140 ( .A(n28351), .B(n28350), .Z(n28355) );
  NAND U29141 ( .A(n28353), .B(n28352), .Z(n28354) );
  NAND U29142 ( .A(n28355), .B(n28354), .Z(n28370) );
  XNOR U29143 ( .A(n28369), .B(n28370), .Z(n28361) );
  XNOR U29144 ( .A(n28362), .B(n28361), .Z(n28363) );
  XNOR U29145 ( .A(n28364), .B(n28363), .Z(n28505) );
  XNOR U29146 ( .A(sreg[429]), .B(n28505), .Z(n28507) );
  NANDN U29147 ( .A(sreg[428]), .B(n28356), .Z(n28360) );
  NAND U29148 ( .A(n28358), .B(n28357), .Z(n28359) );
  NAND U29149 ( .A(n28360), .B(n28359), .Z(n28506) );
  XNOR U29150 ( .A(n28507), .B(n28506), .Z(c[429]) );
  NANDN U29151 ( .A(n28362), .B(n28361), .Z(n28366) );
  NANDN U29152 ( .A(n28364), .B(n28363), .Z(n28365) );
  AND U29153 ( .A(n28366), .B(n28365), .Z(n28513) );
  NANDN U29154 ( .A(n28368), .B(n28367), .Z(n28372) );
  NANDN U29155 ( .A(n28370), .B(n28369), .Z(n28371) );
  AND U29156 ( .A(n28372), .B(n28371), .Z(n28511) );
  NANDN U29157 ( .A(n28374), .B(n28373), .Z(n28378) );
  NANDN U29158 ( .A(n28376), .B(n28375), .Z(n28377) );
  AND U29159 ( .A(n28378), .B(n28377), .Z(n28523) );
  NANDN U29160 ( .A(n28380), .B(n28379), .Z(n28384) );
  NAND U29161 ( .A(n28382), .B(n28381), .Z(n28383) );
  AND U29162 ( .A(n28384), .B(n28383), .Z(n28522) );
  XNOR U29163 ( .A(n28523), .B(n28522), .Z(n28525) );
  NANDN U29164 ( .A(n28386), .B(n28385), .Z(n28390) );
  NANDN U29165 ( .A(n28388), .B(n28387), .Z(n28389) );
  AND U29166 ( .A(n28390), .B(n28389), .Z(n28600) );
  NAND U29167 ( .A(n38385), .B(n28391), .Z(n28393) );
  XOR U29168 ( .A(b[27]), .B(a[180]), .Z(n28546) );
  NAND U29169 ( .A(n38343), .B(n28546), .Z(n28392) );
  AND U29170 ( .A(n28393), .B(n28392), .Z(n28607) );
  NAND U29171 ( .A(n183), .B(n28394), .Z(n28396) );
  XOR U29172 ( .A(b[5]), .B(a[202]), .Z(n28549) );
  NAND U29173 ( .A(n36296), .B(n28549), .Z(n28395) );
  AND U29174 ( .A(n28396), .B(n28395), .Z(n28605) );
  NAND U29175 ( .A(n190), .B(n28397), .Z(n28399) );
  XOR U29176 ( .A(b[19]), .B(a[188]), .Z(n28552) );
  NAND U29177 ( .A(n37821), .B(n28552), .Z(n28398) );
  NAND U29178 ( .A(n28399), .B(n28398), .Z(n28604) );
  XNOR U29179 ( .A(n28605), .B(n28604), .Z(n28606) );
  XNOR U29180 ( .A(n28607), .B(n28606), .Z(n28598) );
  NAND U29181 ( .A(n38470), .B(n28400), .Z(n28402) );
  XOR U29182 ( .A(b[31]), .B(a[176]), .Z(n28555) );
  NAND U29183 ( .A(n38453), .B(n28555), .Z(n28401) );
  AND U29184 ( .A(n28402), .B(n28401), .Z(n28567) );
  NAND U29185 ( .A(n181), .B(n28403), .Z(n28405) );
  XOR U29186 ( .A(b[3]), .B(a[204]), .Z(n28558) );
  NAND U29187 ( .A(n182), .B(n28558), .Z(n28404) );
  AND U29188 ( .A(n28405), .B(n28404), .Z(n28565) );
  NAND U29189 ( .A(n189), .B(n28406), .Z(n28408) );
  XOR U29190 ( .A(b[17]), .B(a[190]), .Z(n28561) );
  NAND U29191 ( .A(n37652), .B(n28561), .Z(n28407) );
  NAND U29192 ( .A(n28408), .B(n28407), .Z(n28564) );
  XNOR U29193 ( .A(n28565), .B(n28564), .Z(n28566) );
  XOR U29194 ( .A(n28567), .B(n28566), .Z(n28599) );
  XOR U29195 ( .A(n28598), .B(n28599), .Z(n28601) );
  XOR U29196 ( .A(n28600), .B(n28601), .Z(n28535) );
  NANDN U29197 ( .A(n28410), .B(n28409), .Z(n28414) );
  NANDN U29198 ( .A(n28412), .B(n28411), .Z(n28413) );
  AND U29199 ( .A(n28414), .B(n28413), .Z(n28588) );
  NANDN U29200 ( .A(n28416), .B(n28415), .Z(n28420) );
  NANDN U29201 ( .A(n28418), .B(n28417), .Z(n28419) );
  NAND U29202 ( .A(n28420), .B(n28419), .Z(n28589) );
  XNOR U29203 ( .A(n28588), .B(n28589), .Z(n28590) );
  NANDN U29204 ( .A(n28422), .B(n28421), .Z(n28426) );
  NANDN U29205 ( .A(n28424), .B(n28423), .Z(n28425) );
  NAND U29206 ( .A(n28426), .B(n28425), .Z(n28591) );
  XNOR U29207 ( .A(n28590), .B(n28591), .Z(n28534) );
  XNOR U29208 ( .A(n28535), .B(n28534), .Z(n28537) );
  NANDN U29209 ( .A(n28428), .B(n28427), .Z(n28432) );
  NANDN U29210 ( .A(n28430), .B(n28429), .Z(n28431) );
  AND U29211 ( .A(n28432), .B(n28431), .Z(n28536) );
  XOR U29212 ( .A(n28537), .B(n28536), .Z(n28649) );
  NANDN U29213 ( .A(n28434), .B(n28433), .Z(n28438) );
  NANDN U29214 ( .A(n28436), .B(n28435), .Z(n28437) );
  AND U29215 ( .A(n28438), .B(n28437), .Z(n28646) );
  NANDN U29216 ( .A(n28440), .B(n28439), .Z(n28444) );
  NANDN U29217 ( .A(n28442), .B(n28441), .Z(n28443) );
  AND U29218 ( .A(n28444), .B(n28443), .Z(n28531) );
  NANDN U29219 ( .A(n28446), .B(n28445), .Z(n28450) );
  OR U29220 ( .A(n28448), .B(n28447), .Z(n28449) );
  AND U29221 ( .A(n28450), .B(n28449), .Z(n28529) );
  NANDN U29222 ( .A(n28452), .B(n28451), .Z(n28456) );
  NANDN U29223 ( .A(n28454), .B(n28453), .Z(n28455) );
  AND U29224 ( .A(n28456), .B(n28455), .Z(n28595) );
  NANDN U29225 ( .A(n28458), .B(n28457), .Z(n28462) );
  NANDN U29226 ( .A(n28460), .B(n28459), .Z(n28461) );
  NAND U29227 ( .A(n28462), .B(n28461), .Z(n28594) );
  XNOR U29228 ( .A(n28595), .B(n28594), .Z(n28597) );
  AND U29229 ( .A(b[0]), .B(a[206]), .Z(n28463) );
  XOR U29230 ( .A(b[1]), .B(n28463), .Z(n28465) );
  NANDN U29231 ( .A(b[0]), .B(a[205]), .Z(n28464) );
  AND U29232 ( .A(n28465), .B(n28464), .Z(n28542) );
  NAND U29233 ( .A(n194), .B(n28466), .Z(n28468) );
  XOR U29234 ( .A(b[29]), .B(a[178]), .Z(n28619) );
  NAND U29235 ( .A(n38456), .B(n28619), .Z(n28467) );
  AND U29236 ( .A(n28468), .B(n28467), .Z(n28541) );
  AND U29237 ( .A(b[31]), .B(a[174]), .Z(n28540) );
  XOR U29238 ( .A(n28541), .B(n28540), .Z(n28543) );
  XNOR U29239 ( .A(n28542), .B(n28543), .Z(n28583) );
  NAND U29240 ( .A(n38185), .B(n28469), .Z(n28471) );
  XOR U29241 ( .A(b[23]), .B(a[184]), .Z(n28622) );
  NAND U29242 ( .A(n38132), .B(n28622), .Z(n28470) );
  AND U29243 ( .A(n28471), .B(n28470), .Z(n28612) );
  NAND U29244 ( .A(n184), .B(n28472), .Z(n28474) );
  XOR U29245 ( .A(b[7]), .B(a[200]), .Z(n28625) );
  NAND U29246 ( .A(n36592), .B(n28625), .Z(n28473) );
  AND U29247 ( .A(n28474), .B(n28473), .Z(n28611) );
  NAND U29248 ( .A(n38289), .B(n28475), .Z(n28477) );
  XOR U29249 ( .A(b[25]), .B(a[182]), .Z(n28628) );
  NAND U29250 ( .A(n38247), .B(n28628), .Z(n28476) );
  NAND U29251 ( .A(n28477), .B(n28476), .Z(n28610) );
  XOR U29252 ( .A(n28611), .B(n28610), .Z(n28613) );
  XOR U29253 ( .A(n28612), .B(n28613), .Z(n28582) );
  XOR U29254 ( .A(n28583), .B(n28582), .Z(n28585) );
  NAND U29255 ( .A(n187), .B(n28478), .Z(n28480) );
  XOR U29256 ( .A(b[13]), .B(a[194]), .Z(n28631) );
  NAND U29257 ( .A(n37295), .B(n28631), .Z(n28479) );
  AND U29258 ( .A(n28480), .B(n28479), .Z(n28577) );
  NAND U29259 ( .A(n186), .B(n28481), .Z(n28483) );
  XOR U29260 ( .A(b[11]), .B(a[196]), .Z(n28634) );
  NAND U29261 ( .A(n37097), .B(n28634), .Z(n28482) );
  NAND U29262 ( .A(n28483), .B(n28482), .Z(n28576) );
  XNOR U29263 ( .A(n28577), .B(n28576), .Z(n28579) );
  NAND U29264 ( .A(n188), .B(n28484), .Z(n28486) );
  XOR U29265 ( .A(b[15]), .B(a[192]), .Z(n28637) );
  NAND U29266 ( .A(n37382), .B(n28637), .Z(n28485) );
  AND U29267 ( .A(n28486), .B(n28485), .Z(n28573) );
  NAND U29268 ( .A(n38064), .B(n28487), .Z(n28489) );
  XOR U29269 ( .A(b[21]), .B(a[186]), .Z(n28640) );
  NAND U29270 ( .A(n37993), .B(n28640), .Z(n28488) );
  AND U29271 ( .A(n28489), .B(n28488), .Z(n28571) );
  NAND U29272 ( .A(n185), .B(n28490), .Z(n28492) );
  XOR U29273 ( .A(b[9]), .B(a[198]), .Z(n28643) );
  NAND U29274 ( .A(n36805), .B(n28643), .Z(n28491) );
  NAND U29275 ( .A(n28492), .B(n28491), .Z(n28570) );
  XNOR U29276 ( .A(n28571), .B(n28570), .Z(n28572) );
  XNOR U29277 ( .A(n28573), .B(n28572), .Z(n28578) );
  XOR U29278 ( .A(n28579), .B(n28578), .Z(n28584) );
  XNOR U29279 ( .A(n28585), .B(n28584), .Z(n28596) );
  XNOR U29280 ( .A(n28597), .B(n28596), .Z(n28528) );
  XNOR U29281 ( .A(n28529), .B(n28528), .Z(n28530) );
  XOR U29282 ( .A(n28531), .B(n28530), .Z(n28647) );
  XNOR U29283 ( .A(n28646), .B(n28647), .Z(n28648) );
  XNOR U29284 ( .A(n28649), .B(n28648), .Z(n28524) );
  XOR U29285 ( .A(n28525), .B(n28524), .Z(n28517) );
  NANDN U29286 ( .A(n28494), .B(n28493), .Z(n28498) );
  NANDN U29287 ( .A(n28496), .B(n28495), .Z(n28497) );
  AND U29288 ( .A(n28498), .B(n28497), .Z(n28516) );
  XNOR U29289 ( .A(n28517), .B(n28516), .Z(n28518) );
  NANDN U29290 ( .A(n28500), .B(n28499), .Z(n28504) );
  NAND U29291 ( .A(n28502), .B(n28501), .Z(n28503) );
  NAND U29292 ( .A(n28504), .B(n28503), .Z(n28519) );
  XNOR U29293 ( .A(n28518), .B(n28519), .Z(n28510) );
  XNOR U29294 ( .A(n28511), .B(n28510), .Z(n28512) );
  XNOR U29295 ( .A(n28513), .B(n28512), .Z(n28652) );
  XNOR U29296 ( .A(sreg[430]), .B(n28652), .Z(n28654) );
  NANDN U29297 ( .A(sreg[429]), .B(n28505), .Z(n28509) );
  NAND U29298 ( .A(n28507), .B(n28506), .Z(n28508) );
  NAND U29299 ( .A(n28509), .B(n28508), .Z(n28653) );
  XNOR U29300 ( .A(n28654), .B(n28653), .Z(c[430]) );
  NANDN U29301 ( .A(n28511), .B(n28510), .Z(n28515) );
  NANDN U29302 ( .A(n28513), .B(n28512), .Z(n28514) );
  AND U29303 ( .A(n28515), .B(n28514), .Z(n28660) );
  NANDN U29304 ( .A(n28517), .B(n28516), .Z(n28521) );
  NANDN U29305 ( .A(n28519), .B(n28518), .Z(n28520) );
  AND U29306 ( .A(n28521), .B(n28520), .Z(n28658) );
  NANDN U29307 ( .A(n28523), .B(n28522), .Z(n28527) );
  NAND U29308 ( .A(n28525), .B(n28524), .Z(n28526) );
  AND U29309 ( .A(n28527), .B(n28526), .Z(n28665) );
  NANDN U29310 ( .A(n28529), .B(n28528), .Z(n28533) );
  NANDN U29311 ( .A(n28531), .B(n28530), .Z(n28532) );
  AND U29312 ( .A(n28533), .B(n28532), .Z(n28670) );
  NANDN U29313 ( .A(n28535), .B(n28534), .Z(n28539) );
  NAND U29314 ( .A(n28537), .B(n28536), .Z(n28538) );
  AND U29315 ( .A(n28539), .B(n28538), .Z(n28669) );
  XNOR U29316 ( .A(n28670), .B(n28669), .Z(n28672) );
  NANDN U29317 ( .A(n28541), .B(n28540), .Z(n28545) );
  NANDN U29318 ( .A(n28543), .B(n28542), .Z(n28544) );
  AND U29319 ( .A(n28545), .B(n28544), .Z(n28735) );
  NAND U29320 ( .A(n38385), .B(n28546), .Z(n28548) );
  XOR U29321 ( .A(b[27]), .B(a[181]), .Z(n28681) );
  NAND U29322 ( .A(n38343), .B(n28681), .Z(n28547) );
  AND U29323 ( .A(n28548), .B(n28547), .Z(n28742) );
  NAND U29324 ( .A(n183), .B(n28549), .Z(n28551) );
  XOR U29325 ( .A(b[5]), .B(a[203]), .Z(n28684) );
  NAND U29326 ( .A(n36296), .B(n28684), .Z(n28550) );
  AND U29327 ( .A(n28551), .B(n28550), .Z(n28740) );
  NAND U29328 ( .A(n190), .B(n28552), .Z(n28554) );
  XOR U29329 ( .A(b[19]), .B(a[189]), .Z(n28687) );
  NAND U29330 ( .A(n37821), .B(n28687), .Z(n28553) );
  NAND U29331 ( .A(n28554), .B(n28553), .Z(n28739) );
  XNOR U29332 ( .A(n28740), .B(n28739), .Z(n28741) );
  XNOR U29333 ( .A(n28742), .B(n28741), .Z(n28733) );
  NAND U29334 ( .A(n38470), .B(n28555), .Z(n28557) );
  XOR U29335 ( .A(b[31]), .B(a[177]), .Z(n28690) );
  NAND U29336 ( .A(n38453), .B(n28690), .Z(n28556) );
  AND U29337 ( .A(n28557), .B(n28556), .Z(n28702) );
  NAND U29338 ( .A(n181), .B(n28558), .Z(n28560) );
  XOR U29339 ( .A(b[3]), .B(a[205]), .Z(n28693) );
  NAND U29340 ( .A(n182), .B(n28693), .Z(n28559) );
  AND U29341 ( .A(n28560), .B(n28559), .Z(n28700) );
  NAND U29342 ( .A(n189), .B(n28561), .Z(n28563) );
  XOR U29343 ( .A(b[17]), .B(a[191]), .Z(n28696) );
  NAND U29344 ( .A(n37652), .B(n28696), .Z(n28562) );
  NAND U29345 ( .A(n28563), .B(n28562), .Z(n28699) );
  XNOR U29346 ( .A(n28700), .B(n28699), .Z(n28701) );
  XOR U29347 ( .A(n28702), .B(n28701), .Z(n28734) );
  XOR U29348 ( .A(n28733), .B(n28734), .Z(n28736) );
  XOR U29349 ( .A(n28735), .B(n28736), .Z(n28782) );
  NANDN U29350 ( .A(n28565), .B(n28564), .Z(n28569) );
  NANDN U29351 ( .A(n28567), .B(n28566), .Z(n28568) );
  AND U29352 ( .A(n28569), .B(n28568), .Z(n28723) );
  NANDN U29353 ( .A(n28571), .B(n28570), .Z(n28575) );
  NANDN U29354 ( .A(n28573), .B(n28572), .Z(n28574) );
  NAND U29355 ( .A(n28575), .B(n28574), .Z(n28724) );
  XNOR U29356 ( .A(n28723), .B(n28724), .Z(n28725) );
  NANDN U29357 ( .A(n28577), .B(n28576), .Z(n28581) );
  NAND U29358 ( .A(n28579), .B(n28578), .Z(n28580) );
  NAND U29359 ( .A(n28581), .B(n28580), .Z(n28726) );
  XNOR U29360 ( .A(n28725), .B(n28726), .Z(n28781) );
  XNOR U29361 ( .A(n28782), .B(n28781), .Z(n28784) );
  NAND U29362 ( .A(n28583), .B(n28582), .Z(n28587) );
  NAND U29363 ( .A(n28585), .B(n28584), .Z(n28586) );
  AND U29364 ( .A(n28587), .B(n28586), .Z(n28783) );
  XOR U29365 ( .A(n28784), .B(n28783), .Z(n28796) );
  NANDN U29366 ( .A(n28589), .B(n28588), .Z(n28593) );
  NANDN U29367 ( .A(n28591), .B(n28590), .Z(n28592) );
  AND U29368 ( .A(n28593), .B(n28592), .Z(n28793) );
  NANDN U29369 ( .A(n28599), .B(n28598), .Z(n28603) );
  OR U29370 ( .A(n28601), .B(n28600), .Z(n28602) );
  AND U29371 ( .A(n28603), .B(n28602), .Z(n28788) );
  NANDN U29372 ( .A(n28605), .B(n28604), .Z(n28609) );
  NANDN U29373 ( .A(n28607), .B(n28606), .Z(n28608) );
  AND U29374 ( .A(n28609), .B(n28608), .Z(n28730) );
  NANDN U29375 ( .A(n28611), .B(n28610), .Z(n28615) );
  OR U29376 ( .A(n28613), .B(n28612), .Z(n28614) );
  NAND U29377 ( .A(n28615), .B(n28614), .Z(n28729) );
  XNOR U29378 ( .A(n28730), .B(n28729), .Z(n28732) );
  NAND U29379 ( .A(b[0]), .B(a[207]), .Z(n28616) );
  XNOR U29380 ( .A(b[1]), .B(n28616), .Z(n28618) );
  NANDN U29381 ( .A(b[0]), .B(a[206]), .Z(n28617) );
  NAND U29382 ( .A(n28618), .B(n28617), .Z(n28678) );
  NAND U29383 ( .A(n194), .B(n28619), .Z(n28621) );
  XOR U29384 ( .A(b[29]), .B(a[179]), .Z(n28754) );
  NAND U29385 ( .A(n38456), .B(n28754), .Z(n28620) );
  AND U29386 ( .A(n28621), .B(n28620), .Z(n28676) );
  AND U29387 ( .A(b[31]), .B(a[175]), .Z(n28675) );
  XNOR U29388 ( .A(n28676), .B(n28675), .Z(n28677) );
  XNOR U29389 ( .A(n28678), .B(n28677), .Z(n28718) );
  NAND U29390 ( .A(n38185), .B(n28622), .Z(n28624) );
  XOR U29391 ( .A(b[23]), .B(a[185]), .Z(n28757) );
  NAND U29392 ( .A(n38132), .B(n28757), .Z(n28623) );
  AND U29393 ( .A(n28624), .B(n28623), .Z(n28747) );
  NAND U29394 ( .A(n184), .B(n28625), .Z(n28627) );
  XOR U29395 ( .A(b[7]), .B(a[201]), .Z(n28760) );
  NAND U29396 ( .A(n36592), .B(n28760), .Z(n28626) );
  AND U29397 ( .A(n28627), .B(n28626), .Z(n28746) );
  NAND U29398 ( .A(n38289), .B(n28628), .Z(n28630) );
  XOR U29399 ( .A(b[25]), .B(a[183]), .Z(n28763) );
  NAND U29400 ( .A(n38247), .B(n28763), .Z(n28629) );
  NAND U29401 ( .A(n28630), .B(n28629), .Z(n28745) );
  XOR U29402 ( .A(n28746), .B(n28745), .Z(n28748) );
  XOR U29403 ( .A(n28747), .B(n28748), .Z(n28717) );
  XOR U29404 ( .A(n28718), .B(n28717), .Z(n28720) );
  NAND U29405 ( .A(n187), .B(n28631), .Z(n28633) );
  XOR U29406 ( .A(b[13]), .B(a[195]), .Z(n28766) );
  NAND U29407 ( .A(n37295), .B(n28766), .Z(n28632) );
  AND U29408 ( .A(n28633), .B(n28632), .Z(n28712) );
  NAND U29409 ( .A(n186), .B(n28634), .Z(n28636) );
  XOR U29410 ( .A(b[11]), .B(a[197]), .Z(n28769) );
  NAND U29411 ( .A(n37097), .B(n28769), .Z(n28635) );
  NAND U29412 ( .A(n28636), .B(n28635), .Z(n28711) );
  XNOR U29413 ( .A(n28712), .B(n28711), .Z(n28714) );
  NAND U29414 ( .A(n188), .B(n28637), .Z(n28639) );
  XOR U29415 ( .A(b[15]), .B(a[193]), .Z(n28772) );
  NAND U29416 ( .A(n37382), .B(n28772), .Z(n28638) );
  AND U29417 ( .A(n28639), .B(n28638), .Z(n28708) );
  NAND U29418 ( .A(n38064), .B(n28640), .Z(n28642) );
  XOR U29419 ( .A(b[21]), .B(a[187]), .Z(n28775) );
  NAND U29420 ( .A(n37993), .B(n28775), .Z(n28641) );
  AND U29421 ( .A(n28642), .B(n28641), .Z(n28706) );
  NAND U29422 ( .A(n185), .B(n28643), .Z(n28645) );
  XOR U29423 ( .A(b[9]), .B(a[199]), .Z(n28778) );
  NAND U29424 ( .A(n36805), .B(n28778), .Z(n28644) );
  NAND U29425 ( .A(n28645), .B(n28644), .Z(n28705) );
  XNOR U29426 ( .A(n28706), .B(n28705), .Z(n28707) );
  XNOR U29427 ( .A(n28708), .B(n28707), .Z(n28713) );
  XOR U29428 ( .A(n28714), .B(n28713), .Z(n28719) );
  XNOR U29429 ( .A(n28720), .B(n28719), .Z(n28731) );
  XNOR U29430 ( .A(n28732), .B(n28731), .Z(n28787) );
  XNOR U29431 ( .A(n28788), .B(n28787), .Z(n28789) );
  XOR U29432 ( .A(n28790), .B(n28789), .Z(n28794) );
  XNOR U29433 ( .A(n28793), .B(n28794), .Z(n28795) );
  XNOR U29434 ( .A(n28796), .B(n28795), .Z(n28671) );
  XOR U29435 ( .A(n28672), .B(n28671), .Z(n28664) );
  NANDN U29436 ( .A(n28647), .B(n28646), .Z(n28651) );
  NANDN U29437 ( .A(n28649), .B(n28648), .Z(n28650) );
  AND U29438 ( .A(n28651), .B(n28650), .Z(n28663) );
  XOR U29439 ( .A(n28664), .B(n28663), .Z(n28666) );
  XNOR U29440 ( .A(n28665), .B(n28666), .Z(n28657) );
  XNOR U29441 ( .A(n28658), .B(n28657), .Z(n28659) );
  XNOR U29442 ( .A(n28660), .B(n28659), .Z(n28799) );
  XNOR U29443 ( .A(sreg[431]), .B(n28799), .Z(n28801) );
  NANDN U29444 ( .A(sreg[430]), .B(n28652), .Z(n28656) );
  NAND U29445 ( .A(n28654), .B(n28653), .Z(n28655) );
  NAND U29446 ( .A(n28656), .B(n28655), .Z(n28800) );
  XNOR U29447 ( .A(n28801), .B(n28800), .Z(c[431]) );
  NANDN U29448 ( .A(n28658), .B(n28657), .Z(n28662) );
  NANDN U29449 ( .A(n28660), .B(n28659), .Z(n28661) );
  AND U29450 ( .A(n28662), .B(n28661), .Z(n28807) );
  NANDN U29451 ( .A(n28664), .B(n28663), .Z(n28668) );
  NANDN U29452 ( .A(n28666), .B(n28665), .Z(n28667) );
  AND U29453 ( .A(n28668), .B(n28667), .Z(n28805) );
  NANDN U29454 ( .A(n28670), .B(n28669), .Z(n28674) );
  NAND U29455 ( .A(n28672), .B(n28671), .Z(n28673) );
  AND U29456 ( .A(n28674), .B(n28673), .Z(n28812) );
  NANDN U29457 ( .A(n28676), .B(n28675), .Z(n28680) );
  NANDN U29458 ( .A(n28678), .B(n28677), .Z(n28679) );
  AND U29459 ( .A(n28680), .B(n28679), .Z(n28884) );
  NAND U29460 ( .A(n38385), .B(n28681), .Z(n28683) );
  XOR U29461 ( .A(b[27]), .B(a[182]), .Z(n28828) );
  NAND U29462 ( .A(n38343), .B(n28828), .Z(n28682) );
  AND U29463 ( .A(n28683), .B(n28682), .Z(n28891) );
  NAND U29464 ( .A(n183), .B(n28684), .Z(n28686) );
  XOR U29465 ( .A(b[5]), .B(a[204]), .Z(n28831) );
  NAND U29466 ( .A(n36296), .B(n28831), .Z(n28685) );
  AND U29467 ( .A(n28686), .B(n28685), .Z(n28889) );
  NAND U29468 ( .A(n190), .B(n28687), .Z(n28689) );
  XOR U29469 ( .A(b[19]), .B(a[190]), .Z(n28834) );
  NAND U29470 ( .A(n37821), .B(n28834), .Z(n28688) );
  NAND U29471 ( .A(n28689), .B(n28688), .Z(n28888) );
  XNOR U29472 ( .A(n28889), .B(n28888), .Z(n28890) );
  XNOR U29473 ( .A(n28891), .B(n28890), .Z(n28882) );
  NAND U29474 ( .A(n38470), .B(n28690), .Z(n28692) );
  XOR U29475 ( .A(b[31]), .B(a[178]), .Z(n28837) );
  NAND U29476 ( .A(n38453), .B(n28837), .Z(n28691) );
  AND U29477 ( .A(n28692), .B(n28691), .Z(n28849) );
  NAND U29478 ( .A(n181), .B(n28693), .Z(n28695) );
  XOR U29479 ( .A(b[3]), .B(a[206]), .Z(n28840) );
  NAND U29480 ( .A(n182), .B(n28840), .Z(n28694) );
  AND U29481 ( .A(n28695), .B(n28694), .Z(n28847) );
  NAND U29482 ( .A(n189), .B(n28696), .Z(n28698) );
  XOR U29483 ( .A(b[17]), .B(a[192]), .Z(n28843) );
  NAND U29484 ( .A(n37652), .B(n28843), .Z(n28697) );
  NAND U29485 ( .A(n28698), .B(n28697), .Z(n28846) );
  XNOR U29486 ( .A(n28847), .B(n28846), .Z(n28848) );
  XOR U29487 ( .A(n28849), .B(n28848), .Z(n28883) );
  XOR U29488 ( .A(n28882), .B(n28883), .Z(n28885) );
  XOR U29489 ( .A(n28884), .B(n28885), .Z(n28931) );
  NANDN U29490 ( .A(n28700), .B(n28699), .Z(n28704) );
  NANDN U29491 ( .A(n28702), .B(n28701), .Z(n28703) );
  AND U29492 ( .A(n28704), .B(n28703), .Z(n28870) );
  NANDN U29493 ( .A(n28706), .B(n28705), .Z(n28710) );
  NANDN U29494 ( .A(n28708), .B(n28707), .Z(n28709) );
  NAND U29495 ( .A(n28710), .B(n28709), .Z(n28871) );
  XNOR U29496 ( .A(n28870), .B(n28871), .Z(n28872) );
  NANDN U29497 ( .A(n28712), .B(n28711), .Z(n28716) );
  NAND U29498 ( .A(n28714), .B(n28713), .Z(n28715) );
  NAND U29499 ( .A(n28716), .B(n28715), .Z(n28873) );
  XNOR U29500 ( .A(n28872), .B(n28873), .Z(n28930) );
  XNOR U29501 ( .A(n28931), .B(n28930), .Z(n28933) );
  NAND U29502 ( .A(n28718), .B(n28717), .Z(n28722) );
  NAND U29503 ( .A(n28720), .B(n28719), .Z(n28721) );
  AND U29504 ( .A(n28722), .B(n28721), .Z(n28932) );
  XOR U29505 ( .A(n28933), .B(n28932), .Z(n28944) );
  NANDN U29506 ( .A(n28724), .B(n28723), .Z(n28728) );
  NANDN U29507 ( .A(n28726), .B(n28725), .Z(n28727) );
  AND U29508 ( .A(n28728), .B(n28727), .Z(n28942) );
  NANDN U29509 ( .A(n28734), .B(n28733), .Z(n28738) );
  OR U29510 ( .A(n28736), .B(n28735), .Z(n28737) );
  AND U29511 ( .A(n28738), .B(n28737), .Z(n28937) );
  NANDN U29512 ( .A(n28740), .B(n28739), .Z(n28744) );
  NANDN U29513 ( .A(n28742), .B(n28741), .Z(n28743) );
  AND U29514 ( .A(n28744), .B(n28743), .Z(n28877) );
  NANDN U29515 ( .A(n28746), .B(n28745), .Z(n28750) );
  OR U29516 ( .A(n28748), .B(n28747), .Z(n28749) );
  NAND U29517 ( .A(n28750), .B(n28749), .Z(n28876) );
  XNOR U29518 ( .A(n28877), .B(n28876), .Z(n28878) );
  AND U29519 ( .A(b[0]), .B(a[208]), .Z(n28751) );
  XOR U29520 ( .A(b[1]), .B(n28751), .Z(n28753) );
  NANDN U29521 ( .A(b[0]), .B(a[207]), .Z(n28752) );
  AND U29522 ( .A(n28753), .B(n28752), .Z(n28824) );
  NAND U29523 ( .A(n194), .B(n28754), .Z(n28756) );
  XOR U29524 ( .A(b[29]), .B(a[180]), .Z(n28903) );
  NAND U29525 ( .A(n38456), .B(n28903), .Z(n28755) );
  AND U29526 ( .A(n28756), .B(n28755), .Z(n28823) );
  AND U29527 ( .A(b[31]), .B(a[176]), .Z(n28822) );
  XOR U29528 ( .A(n28823), .B(n28822), .Z(n28825) );
  XNOR U29529 ( .A(n28824), .B(n28825), .Z(n28864) );
  NAND U29530 ( .A(n38185), .B(n28757), .Z(n28759) );
  XOR U29531 ( .A(b[23]), .B(a[186]), .Z(n28906) );
  NAND U29532 ( .A(n38132), .B(n28906), .Z(n28758) );
  AND U29533 ( .A(n28759), .B(n28758), .Z(n28897) );
  NAND U29534 ( .A(n184), .B(n28760), .Z(n28762) );
  XOR U29535 ( .A(b[7]), .B(a[202]), .Z(n28909) );
  NAND U29536 ( .A(n36592), .B(n28909), .Z(n28761) );
  AND U29537 ( .A(n28762), .B(n28761), .Z(n28895) );
  NAND U29538 ( .A(n38289), .B(n28763), .Z(n28765) );
  XOR U29539 ( .A(b[25]), .B(a[184]), .Z(n28912) );
  NAND U29540 ( .A(n38247), .B(n28912), .Z(n28764) );
  NAND U29541 ( .A(n28765), .B(n28764), .Z(n28894) );
  XNOR U29542 ( .A(n28895), .B(n28894), .Z(n28896) );
  XOR U29543 ( .A(n28897), .B(n28896), .Z(n28865) );
  XNOR U29544 ( .A(n28864), .B(n28865), .Z(n28866) );
  NAND U29545 ( .A(n187), .B(n28766), .Z(n28768) );
  XOR U29546 ( .A(b[13]), .B(a[196]), .Z(n28915) );
  NAND U29547 ( .A(n37295), .B(n28915), .Z(n28767) );
  AND U29548 ( .A(n28768), .B(n28767), .Z(n28859) );
  NAND U29549 ( .A(n186), .B(n28769), .Z(n28771) );
  XOR U29550 ( .A(b[11]), .B(a[198]), .Z(n28918) );
  NAND U29551 ( .A(n37097), .B(n28918), .Z(n28770) );
  NAND U29552 ( .A(n28771), .B(n28770), .Z(n28858) );
  XNOR U29553 ( .A(n28859), .B(n28858), .Z(n28860) );
  NAND U29554 ( .A(n188), .B(n28772), .Z(n28774) );
  XOR U29555 ( .A(b[15]), .B(a[194]), .Z(n28921) );
  NAND U29556 ( .A(n37382), .B(n28921), .Z(n28773) );
  AND U29557 ( .A(n28774), .B(n28773), .Z(n28855) );
  NAND U29558 ( .A(n38064), .B(n28775), .Z(n28777) );
  XOR U29559 ( .A(b[21]), .B(a[188]), .Z(n28924) );
  NAND U29560 ( .A(n37993), .B(n28924), .Z(n28776) );
  AND U29561 ( .A(n28777), .B(n28776), .Z(n28853) );
  NAND U29562 ( .A(n185), .B(n28778), .Z(n28780) );
  XOR U29563 ( .A(b[9]), .B(a[200]), .Z(n28927) );
  NAND U29564 ( .A(n36805), .B(n28927), .Z(n28779) );
  NAND U29565 ( .A(n28780), .B(n28779), .Z(n28852) );
  XNOR U29566 ( .A(n28853), .B(n28852), .Z(n28854) );
  XOR U29567 ( .A(n28855), .B(n28854), .Z(n28861) );
  XOR U29568 ( .A(n28860), .B(n28861), .Z(n28867) );
  XOR U29569 ( .A(n28866), .B(n28867), .Z(n28879) );
  XNOR U29570 ( .A(n28878), .B(n28879), .Z(n28936) );
  XNOR U29571 ( .A(n28937), .B(n28936), .Z(n28938) );
  XOR U29572 ( .A(n28939), .B(n28938), .Z(n28943) );
  XOR U29573 ( .A(n28942), .B(n28943), .Z(n28945) );
  XOR U29574 ( .A(n28944), .B(n28945), .Z(n28819) );
  NANDN U29575 ( .A(n28782), .B(n28781), .Z(n28786) );
  NAND U29576 ( .A(n28784), .B(n28783), .Z(n28785) );
  AND U29577 ( .A(n28786), .B(n28785), .Z(n28817) );
  NANDN U29578 ( .A(n28788), .B(n28787), .Z(n28792) );
  NANDN U29579 ( .A(n28790), .B(n28789), .Z(n28791) );
  AND U29580 ( .A(n28792), .B(n28791), .Z(n28816) );
  XNOR U29581 ( .A(n28817), .B(n28816), .Z(n28818) );
  XNOR U29582 ( .A(n28819), .B(n28818), .Z(n28810) );
  NANDN U29583 ( .A(n28794), .B(n28793), .Z(n28798) );
  NANDN U29584 ( .A(n28796), .B(n28795), .Z(n28797) );
  NAND U29585 ( .A(n28798), .B(n28797), .Z(n28811) );
  XOR U29586 ( .A(n28810), .B(n28811), .Z(n28813) );
  XNOR U29587 ( .A(n28812), .B(n28813), .Z(n28804) );
  XNOR U29588 ( .A(n28805), .B(n28804), .Z(n28806) );
  XNOR U29589 ( .A(n28807), .B(n28806), .Z(n28948) );
  XNOR U29590 ( .A(sreg[432]), .B(n28948), .Z(n28950) );
  NANDN U29591 ( .A(sreg[431]), .B(n28799), .Z(n28803) );
  NAND U29592 ( .A(n28801), .B(n28800), .Z(n28802) );
  NAND U29593 ( .A(n28803), .B(n28802), .Z(n28949) );
  XNOR U29594 ( .A(n28950), .B(n28949), .Z(c[432]) );
  NANDN U29595 ( .A(n28805), .B(n28804), .Z(n28809) );
  NANDN U29596 ( .A(n28807), .B(n28806), .Z(n28808) );
  AND U29597 ( .A(n28809), .B(n28808), .Z(n28956) );
  NANDN U29598 ( .A(n28811), .B(n28810), .Z(n28815) );
  NANDN U29599 ( .A(n28813), .B(n28812), .Z(n28814) );
  AND U29600 ( .A(n28815), .B(n28814), .Z(n28954) );
  NANDN U29601 ( .A(n28817), .B(n28816), .Z(n28821) );
  NANDN U29602 ( .A(n28819), .B(n28818), .Z(n28820) );
  AND U29603 ( .A(n28821), .B(n28820), .Z(n28962) );
  NANDN U29604 ( .A(n28823), .B(n28822), .Z(n28827) );
  NANDN U29605 ( .A(n28825), .B(n28824), .Z(n28826) );
  AND U29606 ( .A(n28827), .B(n28826), .Z(n29045) );
  NAND U29607 ( .A(n38385), .B(n28828), .Z(n28830) );
  XOR U29608 ( .A(b[27]), .B(a[183]), .Z(n28989) );
  NAND U29609 ( .A(n38343), .B(n28989), .Z(n28829) );
  AND U29610 ( .A(n28830), .B(n28829), .Z(n29052) );
  NAND U29611 ( .A(n183), .B(n28831), .Z(n28833) );
  XOR U29612 ( .A(b[5]), .B(a[205]), .Z(n28992) );
  NAND U29613 ( .A(n36296), .B(n28992), .Z(n28832) );
  AND U29614 ( .A(n28833), .B(n28832), .Z(n29050) );
  NAND U29615 ( .A(n190), .B(n28834), .Z(n28836) );
  XOR U29616 ( .A(b[19]), .B(a[191]), .Z(n28995) );
  NAND U29617 ( .A(n37821), .B(n28995), .Z(n28835) );
  NAND U29618 ( .A(n28836), .B(n28835), .Z(n29049) );
  XNOR U29619 ( .A(n29050), .B(n29049), .Z(n29051) );
  XNOR U29620 ( .A(n29052), .B(n29051), .Z(n29043) );
  NAND U29621 ( .A(n38470), .B(n28837), .Z(n28839) );
  XOR U29622 ( .A(b[31]), .B(a[179]), .Z(n28998) );
  NAND U29623 ( .A(n38453), .B(n28998), .Z(n28838) );
  AND U29624 ( .A(n28839), .B(n28838), .Z(n29010) );
  NAND U29625 ( .A(n181), .B(n28840), .Z(n28842) );
  XOR U29626 ( .A(b[3]), .B(a[207]), .Z(n29001) );
  NAND U29627 ( .A(n182), .B(n29001), .Z(n28841) );
  AND U29628 ( .A(n28842), .B(n28841), .Z(n29008) );
  NAND U29629 ( .A(n189), .B(n28843), .Z(n28845) );
  XOR U29630 ( .A(b[17]), .B(a[193]), .Z(n29004) );
  NAND U29631 ( .A(n37652), .B(n29004), .Z(n28844) );
  NAND U29632 ( .A(n28845), .B(n28844), .Z(n29007) );
  XNOR U29633 ( .A(n29008), .B(n29007), .Z(n29009) );
  XOR U29634 ( .A(n29010), .B(n29009), .Z(n29044) );
  XOR U29635 ( .A(n29043), .B(n29044), .Z(n29046) );
  XOR U29636 ( .A(n29045), .B(n29046), .Z(n28978) );
  NANDN U29637 ( .A(n28847), .B(n28846), .Z(n28851) );
  NANDN U29638 ( .A(n28849), .B(n28848), .Z(n28850) );
  AND U29639 ( .A(n28851), .B(n28850), .Z(n29031) );
  NANDN U29640 ( .A(n28853), .B(n28852), .Z(n28857) );
  NANDN U29641 ( .A(n28855), .B(n28854), .Z(n28856) );
  NAND U29642 ( .A(n28857), .B(n28856), .Z(n29032) );
  XNOR U29643 ( .A(n29031), .B(n29032), .Z(n29033) );
  NANDN U29644 ( .A(n28859), .B(n28858), .Z(n28863) );
  NANDN U29645 ( .A(n28861), .B(n28860), .Z(n28862) );
  NAND U29646 ( .A(n28863), .B(n28862), .Z(n29034) );
  XNOR U29647 ( .A(n29033), .B(n29034), .Z(n28977) );
  XNOR U29648 ( .A(n28978), .B(n28977), .Z(n28980) );
  NANDN U29649 ( .A(n28865), .B(n28864), .Z(n28869) );
  NANDN U29650 ( .A(n28867), .B(n28866), .Z(n28868) );
  AND U29651 ( .A(n28869), .B(n28868), .Z(n28979) );
  XOR U29652 ( .A(n28980), .B(n28979), .Z(n29093) );
  NANDN U29653 ( .A(n28871), .B(n28870), .Z(n28875) );
  NANDN U29654 ( .A(n28873), .B(n28872), .Z(n28874) );
  AND U29655 ( .A(n28875), .B(n28874), .Z(n29091) );
  NANDN U29656 ( .A(n28877), .B(n28876), .Z(n28881) );
  NANDN U29657 ( .A(n28879), .B(n28878), .Z(n28880) );
  AND U29658 ( .A(n28881), .B(n28880), .Z(n28974) );
  NANDN U29659 ( .A(n28883), .B(n28882), .Z(n28887) );
  OR U29660 ( .A(n28885), .B(n28884), .Z(n28886) );
  AND U29661 ( .A(n28887), .B(n28886), .Z(n28972) );
  NANDN U29662 ( .A(n28889), .B(n28888), .Z(n28893) );
  NANDN U29663 ( .A(n28891), .B(n28890), .Z(n28892) );
  AND U29664 ( .A(n28893), .B(n28892), .Z(n29038) );
  NANDN U29665 ( .A(n28895), .B(n28894), .Z(n28899) );
  NANDN U29666 ( .A(n28897), .B(n28896), .Z(n28898) );
  NAND U29667 ( .A(n28899), .B(n28898), .Z(n29037) );
  XNOR U29668 ( .A(n29038), .B(n29037), .Z(n29039) );
  NAND U29669 ( .A(b[0]), .B(a[209]), .Z(n28900) );
  XNOR U29670 ( .A(b[1]), .B(n28900), .Z(n28902) );
  NANDN U29671 ( .A(b[0]), .B(a[208]), .Z(n28901) );
  NAND U29672 ( .A(n28902), .B(n28901), .Z(n28986) );
  NAND U29673 ( .A(n194), .B(n28903), .Z(n28905) );
  XOR U29674 ( .A(b[29]), .B(a[181]), .Z(n29061) );
  NAND U29675 ( .A(n38456), .B(n29061), .Z(n28904) );
  AND U29676 ( .A(n28905), .B(n28904), .Z(n28984) );
  AND U29677 ( .A(b[31]), .B(a[177]), .Z(n28983) );
  XNOR U29678 ( .A(n28984), .B(n28983), .Z(n28985) );
  XNOR U29679 ( .A(n28986), .B(n28985), .Z(n29025) );
  NAND U29680 ( .A(n38185), .B(n28906), .Z(n28908) );
  XOR U29681 ( .A(b[23]), .B(a[187]), .Z(n29067) );
  NAND U29682 ( .A(n38132), .B(n29067), .Z(n28907) );
  AND U29683 ( .A(n28908), .B(n28907), .Z(n29058) );
  NAND U29684 ( .A(n184), .B(n28909), .Z(n28911) );
  XOR U29685 ( .A(b[7]), .B(a[203]), .Z(n29070) );
  NAND U29686 ( .A(n36592), .B(n29070), .Z(n28910) );
  AND U29687 ( .A(n28911), .B(n28910), .Z(n29056) );
  NAND U29688 ( .A(n38289), .B(n28912), .Z(n28914) );
  XOR U29689 ( .A(b[25]), .B(a[185]), .Z(n29073) );
  NAND U29690 ( .A(n38247), .B(n29073), .Z(n28913) );
  NAND U29691 ( .A(n28914), .B(n28913), .Z(n29055) );
  XNOR U29692 ( .A(n29056), .B(n29055), .Z(n29057) );
  XOR U29693 ( .A(n29058), .B(n29057), .Z(n29026) );
  XNOR U29694 ( .A(n29025), .B(n29026), .Z(n29027) );
  NAND U29695 ( .A(n187), .B(n28915), .Z(n28917) );
  XOR U29696 ( .A(b[13]), .B(a[197]), .Z(n29076) );
  NAND U29697 ( .A(n37295), .B(n29076), .Z(n28916) );
  AND U29698 ( .A(n28917), .B(n28916), .Z(n29020) );
  NAND U29699 ( .A(n186), .B(n28918), .Z(n28920) );
  XOR U29700 ( .A(b[11]), .B(a[199]), .Z(n29079) );
  NAND U29701 ( .A(n37097), .B(n29079), .Z(n28919) );
  NAND U29702 ( .A(n28920), .B(n28919), .Z(n29019) );
  XNOR U29703 ( .A(n29020), .B(n29019), .Z(n29021) );
  NAND U29704 ( .A(n188), .B(n28921), .Z(n28923) );
  XOR U29705 ( .A(b[15]), .B(a[195]), .Z(n29082) );
  NAND U29706 ( .A(n37382), .B(n29082), .Z(n28922) );
  AND U29707 ( .A(n28923), .B(n28922), .Z(n29016) );
  NAND U29708 ( .A(n38064), .B(n28924), .Z(n28926) );
  XOR U29709 ( .A(b[21]), .B(a[189]), .Z(n29085) );
  NAND U29710 ( .A(n37993), .B(n29085), .Z(n28925) );
  AND U29711 ( .A(n28926), .B(n28925), .Z(n29014) );
  NAND U29712 ( .A(n185), .B(n28927), .Z(n28929) );
  XOR U29713 ( .A(b[9]), .B(a[201]), .Z(n29088) );
  NAND U29714 ( .A(n36805), .B(n29088), .Z(n28928) );
  NAND U29715 ( .A(n28929), .B(n28928), .Z(n29013) );
  XNOR U29716 ( .A(n29014), .B(n29013), .Z(n29015) );
  XOR U29717 ( .A(n29016), .B(n29015), .Z(n29022) );
  XOR U29718 ( .A(n29021), .B(n29022), .Z(n29028) );
  XOR U29719 ( .A(n29027), .B(n29028), .Z(n29040) );
  XNOR U29720 ( .A(n29039), .B(n29040), .Z(n28971) );
  XNOR U29721 ( .A(n28972), .B(n28971), .Z(n28973) );
  XOR U29722 ( .A(n28974), .B(n28973), .Z(n29092) );
  XOR U29723 ( .A(n29091), .B(n29092), .Z(n29094) );
  XOR U29724 ( .A(n29093), .B(n29094), .Z(n28968) );
  NANDN U29725 ( .A(n28931), .B(n28930), .Z(n28935) );
  NAND U29726 ( .A(n28933), .B(n28932), .Z(n28934) );
  AND U29727 ( .A(n28935), .B(n28934), .Z(n28966) );
  NANDN U29728 ( .A(n28937), .B(n28936), .Z(n28941) );
  NANDN U29729 ( .A(n28939), .B(n28938), .Z(n28940) );
  AND U29730 ( .A(n28941), .B(n28940), .Z(n28965) );
  XNOR U29731 ( .A(n28966), .B(n28965), .Z(n28967) );
  XNOR U29732 ( .A(n28968), .B(n28967), .Z(n28959) );
  NANDN U29733 ( .A(n28943), .B(n28942), .Z(n28947) );
  OR U29734 ( .A(n28945), .B(n28944), .Z(n28946) );
  NAND U29735 ( .A(n28947), .B(n28946), .Z(n28960) );
  XNOR U29736 ( .A(n28959), .B(n28960), .Z(n28961) );
  XNOR U29737 ( .A(n28962), .B(n28961), .Z(n28953) );
  XNOR U29738 ( .A(n28954), .B(n28953), .Z(n28955) );
  XNOR U29739 ( .A(n28956), .B(n28955), .Z(n29097) );
  XNOR U29740 ( .A(sreg[433]), .B(n29097), .Z(n29099) );
  NANDN U29741 ( .A(sreg[432]), .B(n28948), .Z(n28952) );
  NAND U29742 ( .A(n28950), .B(n28949), .Z(n28951) );
  NAND U29743 ( .A(n28952), .B(n28951), .Z(n29098) );
  XNOR U29744 ( .A(n29099), .B(n29098), .Z(c[433]) );
  NANDN U29745 ( .A(n28954), .B(n28953), .Z(n28958) );
  NANDN U29746 ( .A(n28956), .B(n28955), .Z(n28957) );
  AND U29747 ( .A(n28958), .B(n28957), .Z(n29105) );
  NANDN U29748 ( .A(n28960), .B(n28959), .Z(n28964) );
  NANDN U29749 ( .A(n28962), .B(n28961), .Z(n28963) );
  AND U29750 ( .A(n28964), .B(n28963), .Z(n29103) );
  NANDN U29751 ( .A(n28966), .B(n28965), .Z(n28970) );
  NANDN U29752 ( .A(n28968), .B(n28967), .Z(n28969) );
  AND U29753 ( .A(n28970), .B(n28969), .Z(n29111) );
  NANDN U29754 ( .A(n28972), .B(n28971), .Z(n28976) );
  NANDN U29755 ( .A(n28974), .B(n28973), .Z(n28975) );
  AND U29756 ( .A(n28976), .B(n28975), .Z(n29115) );
  NANDN U29757 ( .A(n28978), .B(n28977), .Z(n28982) );
  NAND U29758 ( .A(n28980), .B(n28979), .Z(n28981) );
  AND U29759 ( .A(n28982), .B(n28981), .Z(n29114) );
  XNOR U29760 ( .A(n29115), .B(n29114), .Z(n29117) );
  NANDN U29761 ( .A(n28984), .B(n28983), .Z(n28988) );
  NANDN U29762 ( .A(n28986), .B(n28985), .Z(n28987) );
  AND U29763 ( .A(n28988), .B(n28987), .Z(n29192) );
  NAND U29764 ( .A(n38385), .B(n28989), .Z(n28991) );
  XOR U29765 ( .A(b[27]), .B(a[184]), .Z(n29138) );
  NAND U29766 ( .A(n38343), .B(n29138), .Z(n28990) );
  AND U29767 ( .A(n28991), .B(n28990), .Z(n29199) );
  NAND U29768 ( .A(n183), .B(n28992), .Z(n28994) );
  XOR U29769 ( .A(b[5]), .B(a[206]), .Z(n29141) );
  NAND U29770 ( .A(n36296), .B(n29141), .Z(n28993) );
  AND U29771 ( .A(n28994), .B(n28993), .Z(n29197) );
  NAND U29772 ( .A(n190), .B(n28995), .Z(n28997) );
  XOR U29773 ( .A(b[19]), .B(a[192]), .Z(n29144) );
  NAND U29774 ( .A(n37821), .B(n29144), .Z(n28996) );
  NAND U29775 ( .A(n28997), .B(n28996), .Z(n29196) );
  XNOR U29776 ( .A(n29197), .B(n29196), .Z(n29198) );
  XNOR U29777 ( .A(n29199), .B(n29198), .Z(n29190) );
  NAND U29778 ( .A(n38470), .B(n28998), .Z(n29000) );
  XOR U29779 ( .A(b[31]), .B(a[180]), .Z(n29147) );
  NAND U29780 ( .A(n38453), .B(n29147), .Z(n28999) );
  AND U29781 ( .A(n29000), .B(n28999), .Z(n29159) );
  NAND U29782 ( .A(n181), .B(n29001), .Z(n29003) );
  XOR U29783 ( .A(b[3]), .B(a[208]), .Z(n29150) );
  NAND U29784 ( .A(n182), .B(n29150), .Z(n29002) );
  AND U29785 ( .A(n29003), .B(n29002), .Z(n29157) );
  NAND U29786 ( .A(n189), .B(n29004), .Z(n29006) );
  XOR U29787 ( .A(b[17]), .B(a[194]), .Z(n29153) );
  NAND U29788 ( .A(n37652), .B(n29153), .Z(n29005) );
  NAND U29789 ( .A(n29006), .B(n29005), .Z(n29156) );
  XNOR U29790 ( .A(n29157), .B(n29156), .Z(n29158) );
  XOR U29791 ( .A(n29159), .B(n29158), .Z(n29191) );
  XOR U29792 ( .A(n29190), .B(n29191), .Z(n29193) );
  XOR U29793 ( .A(n29192), .B(n29193), .Z(n29127) );
  NANDN U29794 ( .A(n29008), .B(n29007), .Z(n29012) );
  NANDN U29795 ( .A(n29010), .B(n29009), .Z(n29011) );
  AND U29796 ( .A(n29012), .B(n29011), .Z(n29180) );
  NANDN U29797 ( .A(n29014), .B(n29013), .Z(n29018) );
  NANDN U29798 ( .A(n29016), .B(n29015), .Z(n29017) );
  NAND U29799 ( .A(n29018), .B(n29017), .Z(n29181) );
  XNOR U29800 ( .A(n29180), .B(n29181), .Z(n29182) );
  NANDN U29801 ( .A(n29020), .B(n29019), .Z(n29024) );
  NANDN U29802 ( .A(n29022), .B(n29021), .Z(n29023) );
  NAND U29803 ( .A(n29024), .B(n29023), .Z(n29183) );
  XNOR U29804 ( .A(n29182), .B(n29183), .Z(n29126) );
  XNOR U29805 ( .A(n29127), .B(n29126), .Z(n29129) );
  NANDN U29806 ( .A(n29026), .B(n29025), .Z(n29030) );
  NANDN U29807 ( .A(n29028), .B(n29027), .Z(n29029) );
  AND U29808 ( .A(n29030), .B(n29029), .Z(n29128) );
  XOR U29809 ( .A(n29129), .B(n29128), .Z(n29241) );
  NANDN U29810 ( .A(n29032), .B(n29031), .Z(n29036) );
  NANDN U29811 ( .A(n29034), .B(n29033), .Z(n29035) );
  AND U29812 ( .A(n29036), .B(n29035), .Z(n29238) );
  NANDN U29813 ( .A(n29038), .B(n29037), .Z(n29042) );
  NANDN U29814 ( .A(n29040), .B(n29039), .Z(n29041) );
  AND U29815 ( .A(n29042), .B(n29041), .Z(n29123) );
  NANDN U29816 ( .A(n29044), .B(n29043), .Z(n29048) );
  OR U29817 ( .A(n29046), .B(n29045), .Z(n29047) );
  AND U29818 ( .A(n29048), .B(n29047), .Z(n29121) );
  NANDN U29819 ( .A(n29050), .B(n29049), .Z(n29054) );
  NANDN U29820 ( .A(n29052), .B(n29051), .Z(n29053) );
  AND U29821 ( .A(n29054), .B(n29053), .Z(n29187) );
  NANDN U29822 ( .A(n29056), .B(n29055), .Z(n29060) );
  NANDN U29823 ( .A(n29058), .B(n29057), .Z(n29059) );
  NAND U29824 ( .A(n29060), .B(n29059), .Z(n29186) );
  XNOR U29825 ( .A(n29187), .B(n29186), .Z(n29189) );
  NAND U29826 ( .A(n194), .B(n29061), .Z(n29063) );
  XOR U29827 ( .A(b[29]), .B(a[182]), .Z(n29211) );
  NAND U29828 ( .A(n38456), .B(n29211), .Z(n29062) );
  AND U29829 ( .A(n29063), .B(n29062), .Z(n29133) );
  AND U29830 ( .A(b[31]), .B(a[178]), .Z(n29132) );
  XNOR U29831 ( .A(n29133), .B(n29132), .Z(n29134) );
  NAND U29832 ( .A(b[0]), .B(a[210]), .Z(n29064) );
  XNOR U29833 ( .A(b[1]), .B(n29064), .Z(n29066) );
  NANDN U29834 ( .A(b[0]), .B(a[209]), .Z(n29065) );
  NAND U29835 ( .A(n29066), .B(n29065), .Z(n29135) );
  XNOR U29836 ( .A(n29134), .B(n29135), .Z(n29175) );
  NAND U29837 ( .A(n38185), .B(n29067), .Z(n29069) );
  XOR U29838 ( .A(b[23]), .B(a[188]), .Z(n29214) );
  NAND U29839 ( .A(n38132), .B(n29214), .Z(n29068) );
  AND U29840 ( .A(n29069), .B(n29068), .Z(n29204) );
  NAND U29841 ( .A(n184), .B(n29070), .Z(n29072) );
  XOR U29842 ( .A(b[7]), .B(a[204]), .Z(n29217) );
  NAND U29843 ( .A(n36592), .B(n29217), .Z(n29071) );
  AND U29844 ( .A(n29072), .B(n29071), .Z(n29203) );
  NAND U29845 ( .A(n38289), .B(n29073), .Z(n29075) );
  XOR U29846 ( .A(b[25]), .B(a[186]), .Z(n29220) );
  NAND U29847 ( .A(n38247), .B(n29220), .Z(n29074) );
  NAND U29848 ( .A(n29075), .B(n29074), .Z(n29202) );
  XOR U29849 ( .A(n29203), .B(n29202), .Z(n29205) );
  XOR U29850 ( .A(n29204), .B(n29205), .Z(n29174) );
  XOR U29851 ( .A(n29175), .B(n29174), .Z(n29177) );
  NAND U29852 ( .A(n187), .B(n29076), .Z(n29078) );
  XOR U29853 ( .A(b[13]), .B(a[198]), .Z(n29223) );
  NAND U29854 ( .A(n37295), .B(n29223), .Z(n29077) );
  AND U29855 ( .A(n29078), .B(n29077), .Z(n29169) );
  NAND U29856 ( .A(n186), .B(n29079), .Z(n29081) );
  XOR U29857 ( .A(b[11]), .B(a[200]), .Z(n29226) );
  NAND U29858 ( .A(n37097), .B(n29226), .Z(n29080) );
  NAND U29859 ( .A(n29081), .B(n29080), .Z(n29168) );
  XNOR U29860 ( .A(n29169), .B(n29168), .Z(n29171) );
  NAND U29861 ( .A(n188), .B(n29082), .Z(n29084) );
  XOR U29862 ( .A(b[15]), .B(a[196]), .Z(n29229) );
  NAND U29863 ( .A(n37382), .B(n29229), .Z(n29083) );
  AND U29864 ( .A(n29084), .B(n29083), .Z(n29165) );
  NAND U29865 ( .A(n38064), .B(n29085), .Z(n29087) );
  XOR U29866 ( .A(b[21]), .B(a[190]), .Z(n29232) );
  NAND U29867 ( .A(n37993), .B(n29232), .Z(n29086) );
  AND U29868 ( .A(n29087), .B(n29086), .Z(n29163) );
  NAND U29869 ( .A(n185), .B(n29088), .Z(n29090) );
  XOR U29870 ( .A(b[9]), .B(a[202]), .Z(n29235) );
  NAND U29871 ( .A(n36805), .B(n29235), .Z(n29089) );
  NAND U29872 ( .A(n29090), .B(n29089), .Z(n29162) );
  XNOR U29873 ( .A(n29163), .B(n29162), .Z(n29164) );
  XNOR U29874 ( .A(n29165), .B(n29164), .Z(n29170) );
  XOR U29875 ( .A(n29171), .B(n29170), .Z(n29176) );
  XNOR U29876 ( .A(n29177), .B(n29176), .Z(n29188) );
  XNOR U29877 ( .A(n29189), .B(n29188), .Z(n29120) );
  XNOR U29878 ( .A(n29121), .B(n29120), .Z(n29122) );
  XOR U29879 ( .A(n29123), .B(n29122), .Z(n29239) );
  XNOR U29880 ( .A(n29238), .B(n29239), .Z(n29240) );
  XNOR U29881 ( .A(n29241), .B(n29240), .Z(n29116) );
  XOR U29882 ( .A(n29117), .B(n29116), .Z(n29109) );
  NANDN U29883 ( .A(n29092), .B(n29091), .Z(n29096) );
  OR U29884 ( .A(n29094), .B(n29093), .Z(n29095) );
  AND U29885 ( .A(n29096), .B(n29095), .Z(n29108) );
  XNOR U29886 ( .A(n29109), .B(n29108), .Z(n29110) );
  XNOR U29887 ( .A(n29111), .B(n29110), .Z(n29102) );
  XNOR U29888 ( .A(n29103), .B(n29102), .Z(n29104) );
  XNOR U29889 ( .A(n29105), .B(n29104), .Z(n29244) );
  XNOR U29890 ( .A(sreg[434]), .B(n29244), .Z(n29246) );
  NANDN U29891 ( .A(sreg[433]), .B(n29097), .Z(n29101) );
  NAND U29892 ( .A(n29099), .B(n29098), .Z(n29100) );
  NAND U29893 ( .A(n29101), .B(n29100), .Z(n29245) );
  XNOR U29894 ( .A(n29246), .B(n29245), .Z(c[434]) );
  NANDN U29895 ( .A(n29103), .B(n29102), .Z(n29107) );
  NANDN U29896 ( .A(n29105), .B(n29104), .Z(n29106) );
  AND U29897 ( .A(n29107), .B(n29106), .Z(n29252) );
  NANDN U29898 ( .A(n29109), .B(n29108), .Z(n29113) );
  NANDN U29899 ( .A(n29111), .B(n29110), .Z(n29112) );
  AND U29900 ( .A(n29113), .B(n29112), .Z(n29250) );
  NANDN U29901 ( .A(n29115), .B(n29114), .Z(n29119) );
  NAND U29902 ( .A(n29117), .B(n29116), .Z(n29118) );
  AND U29903 ( .A(n29119), .B(n29118), .Z(n29257) );
  NANDN U29904 ( .A(n29121), .B(n29120), .Z(n29125) );
  NANDN U29905 ( .A(n29123), .B(n29122), .Z(n29124) );
  AND U29906 ( .A(n29125), .B(n29124), .Z(n29262) );
  NANDN U29907 ( .A(n29127), .B(n29126), .Z(n29131) );
  NAND U29908 ( .A(n29129), .B(n29128), .Z(n29130) );
  AND U29909 ( .A(n29131), .B(n29130), .Z(n29261) );
  XNOR U29910 ( .A(n29262), .B(n29261), .Z(n29264) );
  NANDN U29911 ( .A(n29133), .B(n29132), .Z(n29137) );
  NANDN U29912 ( .A(n29135), .B(n29134), .Z(n29136) );
  AND U29913 ( .A(n29137), .B(n29136), .Z(n29327) );
  NAND U29914 ( .A(n38385), .B(n29138), .Z(n29140) );
  XOR U29915 ( .A(b[27]), .B(a[185]), .Z(n29273) );
  NAND U29916 ( .A(n38343), .B(n29273), .Z(n29139) );
  AND U29917 ( .A(n29140), .B(n29139), .Z(n29334) );
  NAND U29918 ( .A(n183), .B(n29141), .Z(n29143) );
  XOR U29919 ( .A(b[5]), .B(a[207]), .Z(n29276) );
  NAND U29920 ( .A(n36296), .B(n29276), .Z(n29142) );
  AND U29921 ( .A(n29143), .B(n29142), .Z(n29332) );
  NAND U29922 ( .A(n190), .B(n29144), .Z(n29146) );
  XOR U29923 ( .A(b[19]), .B(a[193]), .Z(n29279) );
  NAND U29924 ( .A(n37821), .B(n29279), .Z(n29145) );
  NAND U29925 ( .A(n29146), .B(n29145), .Z(n29331) );
  XNOR U29926 ( .A(n29332), .B(n29331), .Z(n29333) );
  XNOR U29927 ( .A(n29334), .B(n29333), .Z(n29325) );
  NAND U29928 ( .A(n38470), .B(n29147), .Z(n29149) );
  XOR U29929 ( .A(b[31]), .B(a[181]), .Z(n29282) );
  NAND U29930 ( .A(n38453), .B(n29282), .Z(n29148) );
  AND U29931 ( .A(n29149), .B(n29148), .Z(n29294) );
  NAND U29932 ( .A(n181), .B(n29150), .Z(n29152) );
  XOR U29933 ( .A(b[3]), .B(a[209]), .Z(n29285) );
  NAND U29934 ( .A(n182), .B(n29285), .Z(n29151) );
  AND U29935 ( .A(n29152), .B(n29151), .Z(n29292) );
  NAND U29936 ( .A(n189), .B(n29153), .Z(n29155) );
  XOR U29937 ( .A(b[17]), .B(a[195]), .Z(n29288) );
  NAND U29938 ( .A(n37652), .B(n29288), .Z(n29154) );
  NAND U29939 ( .A(n29155), .B(n29154), .Z(n29291) );
  XNOR U29940 ( .A(n29292), .B(n29291), .Z(n29293) );
  XOR U29941 ( .A(n29294), .B(n29293), .Z(n29326) );
  XOR U29942 ( .A(n29325), .B(n29326), .Z(n29328) );
  XOR U29943 ( .A(n29327), .B(n29328), .Z(n29374) );
  NANDN U29944 ( .A(n29157), .B(n29156), .Z(n29161) );
  NANDN U29945 ( .A(n29159), .B(n29158), .Z(n29160) );
  AND U29946 ( .A(n29161), .B(n29160), .Z(n29315) );
  NANDN U29947 ( .A(n29163), .B(n29162), .Z(n29167) );
  NANDN U29948 ( .A(n29165), .B(n29164), .Z(n29166) );
  NAND U29949 ( .A(n29167), .B(n29166), .Z(n29316) );
  XNOR U29950 ( .A(n29315), .B(n29316), .Z(n29317) );
  NANDN U29951 ( .A(n29169), .B(n29168), .Z(n29173) );
  NAND U29952 ( .A(n29171), .B(n29170), .Z(n29172) );
  NAND U29953 ( .A(n29173), .B(n29172), .Z(n29318) );
  XNOR U29954 ( .A(n29317), .B(n29318), .Z(n29373) );
  XNOR U29955 ( .A(n29374), .B(n29373), .Z(n29376) );
  NAND U29956 ( .A(n29175), .B(n29174), .Z(n29179) );
  NAND U29957 ( .A(n29177), .B(n29176), .Z(n29178) );
  AND U29958 ( .A(n29179), .B(n29178), .Z(n29375) );
  XOR U29959 ( .A(n29376), .B(n29375), .Z(n29388) );
  NANDN U29960 ( .A(n29181), .B(n29180), .Z(n29185) );
  NANDN U29961 ( .A(n29183), .B(n29182), .Z(n29184) );
  AND U29962 ( .A(n29185), .B(n29184), .Z(n29385) );
  NANDN U29963 ( .A(n29191), .B(n29190), .Z(n29195) );
  OR U29964 ( .A(n29193), .B(n29192), .Z(n29194) );
  AND U29965 ( .A(n29195), .B(n29194), .Z(n29380) );
  NANDN U29966 ( .A(n29197), .B(n29196), .Z(n29201) );
  NANDN U29967 ( .A(n29199), .B(n29198), .Z(n29200) );
  AND U29968 ( .A(n29201), .B(n29200), .Z(n29322) );
  NANDN U29969 ( .A(n29203), .B(n29202), .Z(n29207) );
  OR U29970 ( .A(n29205), .B(n29204), .Z(n29206) );
  NAND U29971 ( .A(n29207), .B(n29206), .Z(n29321) );
  XNOR U29972 ( .A(n29322), .B(n29321), .Z(n29324) );
  NAND U29973 ( .A(b[0]), .B(a[211]), .Z(n29208) );
  XNOR U29974 ( .A(b[1]), .B(n29208), .Z(n29210) );
  NANDN U29975 ( .A(b[0]), .B(a[210]), .Z(n29209) );
  NAND U29976 ( .A(n29210), .B(n29209), .Z(n29270) );
  NAND U29977 ( .A(n194), .B(n29211), .Z(n29213) );
  XOR U29978 ( .A(b[29]), .B(a[183]), .Z(n29346) );
  NAND U29979 ( .A(n38456), .B(n29346), .Z(n29212) );
  AND U29980 ( .A(n29213), .B(n29212), .Z(n29268) );
  AND U29981 ( .A(b[31]), .B(a[179]), .Z(n29267) );
  XNOR U29982 ( .A(n29268), .B(n29267), .Z(n29269) );
  XNOR U29983 ( .A(n29270), .B(n29269), .Z(n29310) );
  NAND U29984 ( .A(n38185), .B(n29214), .Z(n29216) );
  XOR U29985 ( .A(b[23]), .B(a[189]), .Z(n29349) );
  NAND U29986 ( .A(n38132), .B(n29349), .Z(n29215) );
  AND U29987 ( .A(n29216), .B(n29215), .Z(n29339) );
  NAND U29988 ( .A(n184), .B(n29217), .Z(n29219) );
  XOR U29989 ( .A(b[7]), .B(a[205]), .Z(n29352) );
  NAND U29990 ( .A(n36592), .B(n29352), .Z(n29218) );
  AND U29991 ( .A(n29219), .B(n29218), .Z(n29338) );
  NAND U29992 ( .A(n38289), .B(n29220), .Z(n29222) );
  XOR U29993 ( .A(b[25]), .B(a[187]), .Z(n29355) );
  NAND U29994 ( .A(n38247), .B(n29355), .Z(n29221) );
  NAND U29995 ( .A(n29222), .B(n29221), .Z(n29337) );
  XOR U29996 ( .A(n29338), .B(n29337), .Z(n29340) );
  XOR U29997 ( .A(n29339), .B(n29340), .Z(n29309) );
  XOR U29998 ( .A(n29310), .B(n29309), .Z(n29312) );
  NAND U29999 ( .A(n187), .B(n29223), .Z(n29225) );
  XOR U30000 ( .A(b[13]), .B(a[199]), .Z(n29358) );
  NAND U30001 ( .A(n37295), .B(n29358), .Z(n29224) );
  AND U30002 ( .A(n29225), .B(n29224), .Z(n29304) );
  NAND U30003 ( .A(n186), .B(n29226), .Z(n29228) );
  XOR U30004 ( .A(b[11]), .B(a[201]), .Z(n29361) );
  NAND U30005 ( .A(n37097), .B(n29361), .Z(n29227) );
  NAND U30006 ( .A(n29228), .B(n29227), .Z(n29303) );
  XNOR U30007 ( .A(n29304), .B(n29303), .Z(n29306) );
  NAND U30008 ( .A(n188), .B(n29229), .Z(n29231) );
  XOR U30009 ( .A(b[15]), .B(a[197]), .Z(n29364) );
  NAND U30010 ( .A(n37382), .B(n29364), .Z(n29230) );
  AND U30011 ( .A(n29231), .B(n29230), .Z(n29300) );
  NAND U30012 ( .A(n38064), .B(n29232), .Z(n29234) );
  XOR U30013 ( .A(b[21]), .B(a[191]), .Z(n29367) );
  NAND U30014 ( .A(n37993), .B(n29367), .Z(n29233) );
  AND U30015 ( .A(n29234), .B(n29233), .Z(n29298) );
  NAND U30016 ( .A(n185), .B(n29235), .Z(n29237) );
  XOR U30017 ( .A(b[9]), .B(a[203]), .Z(n29370) );
  NAND U30018 ( .A(n36805), .B(n29370), .Z(n29236) );
  NAND U30019 ( .A(n29237), .B(n29236), .Z(n29297) );
  XNOR U30020 ( .A(n29298), .B(n29297), .Z(n29299) );
  XNOR U30021 ( .A(n29300), .B(n29299), .Z(n29305) );
  XOR U30022 ( .A(n29306), .B(n29305), .Z(n29311) );
  XNOR U30023 ( .A(n29312), .B(n29311), .Z(n29323) );
  XNOR U30024 ( .A(n29324), .B(n29323), .Z(n29379) );
  XNOR U30025 ( .A(n29380), .B(n29379), .Z(n29381) );
  XOR U30026 ( .A(n29382), .B(n29381), .Z(n29386) );
  XNOR U30027 ( .A(n29385), .B(n29386), .Z(n29387) );
  XNOR U30028 ( .A(n29388), .B(n29387), .Z(n29263) );
  XOR U30029 ( .A(n29264), .B(n29263), .Z(n29256) );
  NANDN U30030 ( .A(n29239), .B(n29238), .Z(n29243) );
  NANDN U30031 ( .A(n29241), .B(n29240), .Z(n29242) );
  AND U30032 ( .A(n29243), .B(n29242), .Z(n29255) );
  XOR U30033 ( .A(n29256), .B(n29255), .Z(n29258) );
  XNOR U30034 ( .A(n29257), .B(n29258), .Z(n29249) );
  XNOR U30035 ( .A(n29250), .B(n29249), .Z(n29251) );
  XNOR U30036 ( .A(n29252), .B(n29251), .Z(n29391) );
  XNOR U30037 ( .A(sreg[435]), .B(n29391), .Z(n29393) );
  NANDN U30038 ( .A(sreg[434]), .B(n29244), .Z(n29248) );
  NAND U30039 ( .A(n29246), .B(n29245), .Z(n29247) );
  NAND U30040 ( .A(n29248), .B(n29247), .Z(n29392) );
  XNOR U30041 ( .A(n29393), .B(n29392), .Z(c[435]) );
  NANDN U30042 ( .A(n29250), .B(n29249), .Z(n29254) );
  NANDN U30043 ( .A(n29252), .B(n29251), .Z(n29253) );
  AND U30044 ( .A(n29254), .B(n29253), .Z(n29399) );
  NANDN U30045 ( .A(n29256), .B(n29255), .Z(n29260) );
  NANDN U30046 ( .A(n29258), .B(n29257), .Z(n29259) );
  AND U30047 ( .A(n29260), .B(n29259), .Z(n29397) );
  NANDN U30048 ( .A(n29262), .B(n29261), .Z(n29266) );
  NAND U30049 ( .A(n29264), .B(n29263), .Z(n29265) );
  AND U30050 ( .A(n29266), .B(n29265), .Z(n29404) );
  NANDN U30051 ( .A(n29268), .B(n29267), .Z(n29272) );
  NANDN U30052 ( .A(n29270), .B(n29269), .Z(n29271) );
  AND U30053 ( .A(n29272), .B(n29271), .Z(n29474) );
  NAND U30054 ( .A(n38385), .B(n29273), .Z(n29275) );
  XOR U30055 ( .A(b[27]), .B(a[186]), .Z(n29420) );
  NAND U30056 ( .A(n38343), .B(n29420), .Z(n29274) );
  AND U30057 ( .A(n29275), .B(n29274), .Z(n29481) );
  NAND U30058 ( .A(n183), .B(n29276), .Z(n29278) );
  XOR U30059 ( .A(b[5]), .B(a[208]), .Z(n29423) );
  NAND U30060 ( .A(n36296), .B(n29423), .Z(n29277) );
  AND U30061 ( .A(n29278), .B(n29277), .Z(n29479) );
  NAND U30062 ( .A(n190), .B(n29279), .Z(n29281) );
  XOR U30063 ( .A(b[19]), .B(a[194]), .Z(n29426) );
  NAND U30064 ( .A(n37821), .B(n29426), .Z(n29280) );
  NAND U30065 ( .A(n29281), .B(n29280), .Z(n29478) );
  XNOR U30066 ( .A(n29479), .B(n29478), .Z(n29480) );
  XNOR U30067 ( .A(n29481), .B(n29480), .Z(n29472) );
  NAND U30068 ( .A(n38470), .B(n29282), .Z(n29284) );
  XOR U30069 ( .A(b[31]), .B(a[182]), .Z(n29429) );
  NAND U30070 ( .A(n38453), .B(n29429), .Z(n29283) );
  AND U30071 ( .A(n29284), .B(n29283), .Z(n29441) );
  NAND U30072 ( .A(n181), .B(n29285), .Z(n29287) );
  XOR U30073 ( .A(b[3]), .B(a[210]), .Z(n29432) );
  NAND U30074 ( .A(n182), .B(n29432), .Z(n29286) );
  AND U30075 ( .A(n29287), .B(n29286), .Z(n29439) );
  NAND U30076 ( .A(n189), .B(n29288), .Z(n29290) );
  XOR U30077 ( .A(b[17]), .B(a[196]), .Z(n29435) );
  NAND U30078 ( .A(n37652), .B(n29435), .Z(n29289) );
  NAND U30079 ( .A(n29290), .B(n29289), .Z(n29438) );
  XNOR U30080 ( .A(n29439), .B(n29438), .Z(n29440) );
  XOR U30081 ( .A(n29441), .B(n29440), .Z(n29473) );
  XOR U30082 ( .A(n29472), .B(n29473), .Z(n29475) );
  XOR U30083 ( .A(n29474), .B(n29475), .Z(n29521) );
  NANDN U30084 ( .A(n29292), .B(n29291), .Z(n29296) );
  NANDN U30085 ( .A(n29294), .B(n29293), .Z(n29295) );
  AND U30086 ( .A(n29296), .B(n29295), .Z(n29462) );
  NANDN U30087 ( .A(n29298), .B(n29297), .Z(n29302) );
  NANDN U30088 ( .A(n29300), .B(n29299), .Z(n29301) );
  NAND U30089 ( .A(n29302), .B(n29301), .Z(n29463) );
  XNOR U30090 ( .A(n29462), .B(n29463), .Z(n29464) );
  NANDN U30091 ( .A(n29304), .B(n29303), .Z(n29308) );
  NAND U30092 ( .A(n29306), .B(n29305), .Z(n29307) );
  NAND U30093 ( .A(n29308), .B(n29307), .Z(n29465) );
  XNOR U30094 ( .A(n29464), .B(n29465), .Z(n29520) );
  XNOR U30095 ( .A(n29521), .B(n29520), .Z(n29523) );
  NAND U30096 ( .A(n29310), .B(n29309), .Z(n29314) );
  NAND U30097 ( .A(n29312), .B(n29311), .Z(n29313) );
  AND U30098 ( .A(n29314), .B(n29313), .Z(n29522) );
  XOR U30099 ( .A(n29523), .B(n29522), .Z(n29534) );
  NANDN U30100 ( .A(n29316), .B(n29315), .Z(n29320) );
  NANDN U30101 ( .A(n29318), .B(n29317), .Z(n29319) );
  AND U30102 ( .A(n29320), .B(n29319), .Z(n29532) );
  NANDN U30103 ( .A(n29326), .B(n29325), .Z(n29330) );
  OR U30104 ( .A(n29328), .B(n29327), .Z(n29329) );
  AND U30105 ( .A(n29330), .B(n29329), .Z(n29527) );
  NANDN U30106 ( .A(n29332), .B(n29331), .Z(n29336) );
  NANDN U30107 ( .A(n29334), .B(n29333), .Z(n29335) );
  AND U30108 ( .A(n29336), .B(n29335), .Z(n29469) );
  NANDN U30109 ( .A(n29338), .B(n29337), .Z(n29342) );
  OR U30110 ( .A(n29340), .B(n29339), .Z(n29341) );
  NAND U30111 ( .A(n29342), .B(n29341), .Z(n29468) );
  XNOR U30112 ( .A(n29469), .B(n29468), .Z(n29471) );
  NAND U30113 ( .A(b[0]), .B(a[212]), .Z(n29343) );
  XNOR U30114 ( .A(b[1]), .B(n29343), .Z(n29345) );
  NANDN U30115 ( .A(b[0]), .B(a[211]), .Z(n29344) );
  NAND U30116 ( .A(n29345), .B(n29344), .Z(n29417) );
  NAND U30117 ( .A(n194), .B(n29346), .Z(n29348) );
  XOR U30118 ( .A(b[29]), .B(a[184]), .Z(n29493) );
  NAND U30119 ( .A(n38456), .B(n29493), .Z(n29347) );
  AND U30120 ( .A(n29348), .B(n29347), .Z(n29415) );
  AND U30121 ( .A(b[31]), .B(a[180]), .Z(n29414) );
  XNOR U30122 ( .A(n29415), .B(n29414), .Z(n29416) );
  XNOR U30123 ( .A(n29417), .B(n29416), .Z(n29457) );
  NAND U30124 ( .A(n38185), .B(n29349), .Z(n29351) );
  XOR U30125 ( .A(b[23]), .B(a[190]), .Z(n29496) );
  NAND U30126 ( .A(n38132), .B(n29496), .Z(n29350) );
  AND U30127 ( .A(n29351), .B(n29350), .Z(n29486) );
  NAND U30128 ( .A(n184), .B(n29352), .Z(n29354) );
  XOR U30129 ( .A(b[7]), .B(a[206]), .Z(n29499) );
  NAND U30130 ( .A(n36592), .B(n29499), .Z(n29353) );
  AND U30131 ( .A(n29354), .B(n29353), .Z(n29485) );
  NAND U30132 ( .A(n38289), .B(n29355), .Z(n29357) );
  XOR U30133 ( .A(b[25]), .B(a[188]), .Z(n29502) );
  NAND U30134 ( .A(n38247), .B(n29502), .Z(n29356) );
  NAND U30135 ( .A(n29357), .B(n29356), .Z(n29484) );
  XOR U30136 ( .A(n29485), .B(n29484), .Z(n29487) );
  XOR U30137 ( .A(n29486), .B(n29487), .Z(n29456) );
  XOR U30138 ( .A(n29457), .B(n29456), .Z(n29459) );
  NAND U30139 ( .A(n187), .B(n29358), .Z(n29360) );
  XOR U30140 ( .A(b[13]), .B(a[200]), .Z(n29505) );
  NAND U30141 ( .A(n37295), .B(n29505), .Z(n29359) );
  AND U30142 ( .A(n29360), .B(n29359), .Z(n29451) );
  NAND U30143 ( .A(n186), .B(n29361), .Z(n29363) );
  XOR U30144 ( .A(b[11]), .B(a[202]), .Z(n29508) );
  NAND U30145 ( .A(n37097), .B(n29508), .Z(n29362) );
  NAND U30146 ( .A(n29363), .B(n29362), .Z(n29450) );
  XNOR U30147 ( .A(n29451), .B(n29450), .Z(n29453) );
  NAND U30148 ( .A(n188), .B(n29364), .Z(n29366) );
  XOR U30149 ( .A(b[15]), .B(a[198]), .Z(n29511) );
  NAND U30150 ( .A(n37382), .B(n29511), .Z(n29365) );
  AND U30151 ( .A(n29366), .B(n29365), .Z(n29447) );
  NAND U30152 ( .A(n38064), .B(n29367), .Z(n29369) );
  XOR U30153 ( .A(b[21]), .B(a[192]), .Z(n29514) );
  NAND U30154 ( .A(n37993), .B(n29514), .Z(n29368) );
  AND U30155 ( .A(n29369), .B(n29368), .Z(n29445) );
  NAND U30156 ( .A(n185), .B(n29370), .Z(n29372) );
  XOR U30157 ( .A(b[9]), .B(a[204]), .Z(n29517) );
  NAND U30158 ( .A(n36805), .B(n29517), .Z(n29371) );
  NAND U30159 ( .A(n29372), .B(n29371), .Z(n29444) );
  XNOR U30160 ( .A(n29445), .B(n29444), .Z(n29446) );
  XNOR U30161 ( .A(n29447), .B(n29446), .Z(n29452) );
  XOR U30162 ( .A(n29453), .B(n29452), .Z(n29458) );
  XNOR U30163 ( .A(n29459), .B(n29458), .Z(n29470) );
  XNOR U30164 ( .A(n29471), .B(n29470), .Z(n29526) );
  XNOR U30165 ( .A(n29527), .B(n29526), .Z(n29528) );
  XOR U30166 ( .A(n29529), .B(n29528), .Z(n29533) );
  XOR U30167 ( .A(n29532), .B(n29533), .Z(n29535) );
  XOR U30168 ( .A(n29534), .B(n29535), .Z(n29411) );
  NANDN U30169 ( .A(n29374), .B(n29373), .Z(n29378) );
  NAND U30170 ( .A(n29376), .B(n29375), .Z(n29377) );
  AND U30171 ( .A(n29378), .B(n29377), .Z(n29409) );
  NANDN U30172 ( .A(n29380), .B(n29379), .Z(n29384) );
  NANDN U30173 ( .A(n29382), .B(n29381), .Z(n29383) );
  AND U30174 ( .A(n29384), .B(n29383), .Z(n29408) );
  XNOR U30175 ( .A(n29409), .B(n29408), .Z(n29410) );
  XNOR U30176 ( .A(n29411), .B(n29410), .Z(n29402) );
  NANDN U30177 ( .A(n29386), .B(n29385), .Z(n29390) );
  NANDN U30178 ( .A(n29388), .B(n29387), .Z(n29389) );
  NAND U30179 ( .A(n29390), .B(n29389), .Z(n29403) );
  XOR U30180 ( .A(n29402), .B(n29403), .Z(n29405) );
  XNOR U30181 ( .A(n29404), .B(n29405), .Z(n29396) );
  XNOR U30182 ( .A(n29397), .B(n29396), .Z(n29398) );
  XNOR U30183 ( .A(n29399), .B(n29398), .Z(n29538) );
  XNOR U30184 ( .A(sreg[436]), .B(n29538), .Z(n29540) );
  NANDN U30185 ( .A(sreg[435]), .B(n29391), .Z(n29395) );
  NAND U30186 ( .A(n29393), .B(n29392), .Z(n29394) );
  NAND U30187 ( .A(n29395), .B(n29394), .Z(n29539) );
  XNOR U30188 ( .A(n29540), .B(n29539), .Z(c[436]) );
  NANDN U30189 ( .A(n29397), .B(n29396), .Z(n29401) );
  NANDN U30190 ( .A(n29399), .B(n29398), .Z(n29400) );
  AND U30191 ( .A(n29401), .B(n29400), .Z(n29546) );
  NANDN U30192 ( .A(n29403), .B(n29402), .Z(n29407) );
  NANDN U30193 ( .A(n29405), .B(n29404), .Z(n29406) );
  AND U30194 ( .A(n29407), .B(n29406), .Z(n29544) );
  NANDN U30195 ( .A(n29409), .B(n29408), .Z(n29413) );
  NANDN U30196 ( .A(n29411), .B(n29410), .Z(n29412) );
  AND U30197 ( .A(n29413), .B(n29412), .Z(n29552) );
  NANDN U30198 ( .A(n29415), .B(n29414), .Z(n29419) );
  NANDN U30199 ( .A(n29417), .B(n29416), .Z(n29418) );
  AND U30200 ( .A(n29419), .B(n29418), .Z(n29623) );
  NAND U30201 ( .A(n38385), .B(n29420), .Z(n29422) );
  XOR U30202 ( .A(b[27]), .B(a[187]), .Z(n29567) );
  NAND U30203 ( .A(n38343), .B(n29567), .Z(n29421) );
  AND U30204 ( .A(n29422), .B(n29421), .Z(n29630) );
  NAND U30205 ( .A(n183), .B(n29423), .Z(n29425) );
  XOR U30206 ( .A(b[5]), .B(a[209]), .Z(n29570) );
  NAND U30207 ( .A(n36296), .B(n29570), .Z(n29424) );
  AND U30208 ( .A(n29425), .B(n29424), .Z(n29628) );
  NAND U30209 ( .A(n190), .B(n29426), .Z(n29428) );
  XOR U30210 ( .A(b[19]), .B(a[195]), .Z(n29573) );
  NAND U30211 ( .A(n37821), .B(n29573), .Z(n29427) );
  NAND U30212 ( .A(n29428), .B(n29427), .Z(n29627) );
  XNOR U30213 ( .A(n29628), .B(n29627), .Z(n29629) );
  XNOR U30214 ( .A(n29630), .B(n29629), .Z(n29621) );
  NAND U30215 ( .A(n38470), .B(n29429), .Z(n29431) );
  XOR U30216 ( .A(b[31]), .B(a[183]), .Z(n29576) );
  NAND U30217 ( .A(n38453), .B(n29576), .Z(n29430) );
  AND U30218 ( .A(n29431), .B(n29430), .Z(n29588) );
  NAND U30219 ( .A(n181), .B(n29432), .Z(n29434) );
  XOR U30220 ( .A(b[3]), .B(a[211]), .Z(n29579) );
  NAND U30221 ( .A(n182), .B(n29579), .Z(n29433) );
  AND U30222 ( .A(n29434), .B(n29433), .Z(n29586) );
  NAND U30223 ( .A(n189), .B(n29435), .Z(n29437) );
  XOR U30224 ( .A(b[17]), .B(a[197]), .Z(n29582) );
  NAND U30225 ( .A(n37652), .B(n29582), .Z(n29436) );
  NAND U30226 ( .A(n29437), .B(n29436), .Z(n29585) );
  XNOR U30227 ( .A(n29586), .B(n29585), .Z(n29587) );
  XOR U30228 ( .A(n29588), .B(n29587), .Z(n29622) );
  XOR U30229 ( .A(n29621), .B(n29622), .Z(n29624) );
  XOR U30230 ( .A(n29623), .B(n29624), .Z(n29670) );
  NANDN U30231 ( .A(n29439), .B(n29438), .Z(n29443) );
  NANDN U30232 ( .A(n29441), .B(n29440), .Z(n29442) );
  AND U30233 ( .A(n29443), .B(n29442), .Z(n29609) );
  NANDN U30234 ( .A(n29445), .B(n29444), .Z(n29449) );
  NANDN U30235 ( .A(n29447), .B(n29446), .Z(n29448) );
  NAND U30236 ( .A(n29449), .B(n29448), .Z(n29610) );
  XNOR U30237 ( .A(n29609), .B(n29610), .Z(n29611) );
  NANDN U30238 ( .A(n29451), .B(n29450), .Z(n29455) );
  NAND U30239 ( .A(n29453), .B(n29452), .Z(n29454) );
  NAND U30240 ( .A(n29455), .B(n29454), .Z(n29612) );
  XNOR U30241 ( .A(n29611), .B(n29612), .Z(n29669) );
  XNOR U30242 ( .A(n29670), .B(n29669), .Z(n29672) );
  NAND U30243 ( .A(n29457), .B(n29456), .Z(n29461) );
  NAND U30244 ( .A(n29459), .B(n29458), .Z(n29460) );
  AND U30245 ( .A(n29461), .B(n29460), .Z(n29671) );
  XOR U30246 ( .A(n29672), .B(n29671), .Z(n29683) );
  NANDN U30247 ( .A(n29463), .B(n29462), .Z(n29467) );
  NANDN U30248 ( .A(n29465), .B(n29464), .Z(n29466) );
  AND U30249 ( .A(n29467), .B(n29466), .Z(n29681) );
  NANDN U30250 ( .A(n29473), .B(n29472), .Z(n29477) );
  OR U30251 ( .A(n29475), .B(n29474), .Z(n29476) );
  AND U30252 ( .A(n29477), .B(n29476), .Z(n29676) );
  NANDN U30253 ( .A(n29479), .B(n29478), .Z(n29483) );
  NANDN U30254 ( .A(n29481), .B(n29480), .Z(n29482) );
  AND U30255 ( .A(n29483), .B(n29482), .Z(n29616) );
  NANDN U30256 ( .A(n29485), .B(n29484), .Z(n29489) );
  OR U30257 ( .A(n29487), .B(n29486), .Z(n29488) );
  NAND U30258 ( .A(n29489), .B(n29488), .Z(n29615) );
  XNOR U30259 ( .A(n29616), .B(n29615), .Z(n29617) );
  NAND U30260 ( .A(b[0]), .B(a[213]), .Z(n29490) );
  XNOR U30261 ( .A(b[1]), .B(n29490), .Z(n29492) );
  NANDN U30262 ( .A(b[0]), .B(a[212]), .Z(n29491) );
  NAND U30263 ( .A(n29492), .B(n29491), .Z(n29564) );
  NAND U30264 ( .A(n194), .B(n29493), .Z(n29495) );
  XOR U30265 ( .A(b[29]), .B(a[185]), .Z(n29642) );
  NAND U30266 ( .A(n38456), .B(n29642), .Z(n29494) );
  AND U30267 ( .A(n29495), .B(n29494), .Z(n29562) );
  AND U30268 ( .A(b[31]), .B(a[181]), .Z(n29561) );
  XNOR U30269 ( .A(n29562), .B(n29561), .Z(n29563) );
  XNOR U30270 ( .A(n29564), .B(n29563), .Z(n29603) );
  NAND U30271 ( .A(n38185), .B(n29496), .Z(n29498) );
  XOR U30272 ( .A(b[23]), .B(a[191]), .Z(n29645) );
  NAND U30273 ( .A(n38132), .B(n29645), .Z(n29497) );
  AND U30274 ( .A(n29498), .B(n29497), .Z(n29636) );
  NAND U30275 ( .A(n184), .B(n29499), .Z(n29501) );
  XOR U30276 ( .A(b[7]), .B(a[207]), .Z(n29648) );
  NAND U30277 ( .A(n36592), .B(n29648), .Z(n29500) );
  AND U30278 ( .A(n29501), .B(n29500), .Z(n29634) );
  NAND U30279 ( .A(n38289), .B(n29502), .Z(n29504) );
  XOR U30280 ( .A(b[25]), .B(a[189]), .Z(n29651) );
  NAND U30281 ( .A(n38247), .B(n29651), .Z(n29503) );
  NAND U30282 ( .A(n29504), .B(n29503), .Z(n29633) );
  XNOR U30283 ( .A(n29634), .B(n29633), .Z(n29635) );
  XOR U30284 ( .A(n29636), .B(n29635), .Z(n29604) );
  XNOR U30285 ( .A(n29603), .B(n29604), .Z(n29605) );
  NAND U30286 ( .A(n187), .B(n29505), .Z(n29507) );
  XOR U30287 ( .A(b[13]), .B(a[201]), .Z(n29654) );
  NAND U30288 ( .A(n37295), .B(n29654), .Z(n29506) );
  AND U30289 ( .A(n29507), .B(n29506), .Z(n29598) );
  NAND U30290 ( .A(n186), .B(n29508), .Z(n29510) );
  XOR U30291 ( .A(b[11]), .B(a[203]), .Z(n29657) );
  NAND U30292 ( .A(n37097), .B(n29657), .Z(n29509) );
  NAND U30293 ( .A(n29510), .B(n29509), .Z(n29597) );
  XNOR U30294 ( .A(n29598), .B(n29597), .Z(n29599) );
  NAND U30295 ( .A(n188), .B(n29511), .Z(n29513) );
  XOR U30296 ( .A(b[15]), .B(a[199]), .Z(n29660) );
  NAND U30297 ( .A(n37382), .B(n29660), .Z(n29512) );
  AND U30298 ( .A(n29513), .B(n29512), .Z(n29594) );
  NAND U30299 ( .A(n38064), .B(n29514), .Z(n29516) );
  XOR U30300 ( .A(b[21]), .B(a[193]), .Z(n29663) );
  NAND U30301 ( .A(n37993), .B(n29663), .Z(n29515) );
  AND U30302 ( .A(n29516), .B(n29515), .Z(n29592) );
  NAND U30303 ( .A(n185), .B(n29517), .Z(n29519) );
  XOR U30304 ( .A(b[9]), .B(a[205]), .Z(n29666) );
  NAND U30305 ( .A(n36805), .B(n29666), .Z(n29518) );
  NAND U30306 ( .A(n29519), .B(n29518), .Z(n29591) );
  XNOR U30307 ( .A(n29592), .B(n29591), .Z(n29593) );
  XOR U30308 ( .A(n29594), .B(n29593), .Z(n29600) );
  XOR U30309 ( .A(n29599), .B(n29600), .Z(n29606) );
  XOR U30310 ( .A(n29605), .B(n29606), .Z(n29618) );
  XNOR U30311 ( .A(n29617), .B(n29618), .Z(n29675) );
  XNOR U30312 ( .A(n29676), .B(n29675), .Z(n29677) );
  XOR U30313 ( .A(n29678), .B(n29677), .Z(n29682) );
  XOR U30314 ( .A(n29681), .B(n29682), .Z(n29684) );
  XOR U30315 ( .A(n29683), .B(n29684), .Z(n29558) );
  NANDN U30316 ( .A(n29521), .B(n29520), .Z(n29525) );
  NAND U30317 ( .A(n29523), .B(n29522), .Z(n29524) );
  AND U30318 ( .A(n29525), .B(n29524), .Z(n29556) );
  NANDN U30319 ( .A(n29527), .B(n29526), .Z(n29531) );
  NANDN U30320 ( .A(n29529), .B(n29528), .Z(n29530) );
  AND U30321 ( .A(n29531), .B(n29530), .Z(n29555) );
  XNOR U30322 ( .A(n29556), .B(n29555), .Z(n29557) );
  XNOR U30323 ( .A(n29558), .B(n29557), .Z(n29549) );
  NANDN U30324 ( .A(n29533), .B(n29532), .Z(n29537) );
  OR U30325 ( .A(n29535), .B(n29534), .Z(n29536) );
  NAND U30326 ( .A(n29537), .B(n29536), .Z(n29550) );
  XNOR U30327 ( .A(n29549), .B(n29550), .Z(n29551) );
  XNOR U30328 ( .A(n29552), .B(n29551), .Z(n29543) );
  XNOR U30329 ( .A(n29544), .B(n29543), .Z(n29545) );
  XNOR U30330 ( .A(n29546), .B(n29545), .Z(n29687) );
  XNOR U30331 ( .A(sreg[437]), .B(n29687), .Z(n29689) );
  NANDN U30332 ( .A(sreg[436]), .B(n29538), .Z(n29542) );
  NAND U30333 ( .A(n29540), .B(n29539), .Z(n29541) );
  NAND U30334 ( .A(n29542), .B(n29541), .Z(n29688) );
  XNOR U30335 ( .A(n29689), .B(n29688), .Z(c[437]) );
  NANDN U30336 ( .A(n29544), .B(n29543), .Z(n29548) );
  NANDN U30337 ( .A(n29546), .B(n29545), .Z(n29547) );
  AND U30338 ( .A(n29548), .B(n29547), .Z(n29695) );
  NANDN U30339 ( .A(n29550), .B(n29549), .Z(n29554) );
  NANDN U30340 ( .A(n29552), .B(n29551), .Z(n29553) );
  AND U30341 ( .A(n29554), .B(n29553), .Z(n29693) );
  NANDN U30342 ( .A(n29556), .B(n29555), .Z(n29560) );
  NANDN U30343 ( .A(n29558), .B(n29557), .Z(n29559) );
  AND U30344 ( .A(n29560), .B(n29559), .Z(n29701) );
  NANDN U30345 ( .A(n29562), .B(n29561), .Z(n29566) );
  NANDN U30346 ( .A(n29564), .B(n29563), .Z(n29565) );
  AND U30347 ( .A(n29566), .B(n29565), .Z(n29782) );
  NAND U30348 ( .A(n38385), .B(n29567), .Z(n29569) );
  XOR U30349 ( .A(b[27]), .B(a[188]), .Z(n29728) );
  NAND U30350 ( .A(n38343), .B(n29728), .Z(n29568) );
  AND U30351 ( .A(n29569), .B(n29568), .Z(n29789) );
  NAND U30352 ( .A(n183), .B(n29570), .Z(n29572) );
  XOR U30353 ( .A(b[5]), .B(a[210]), .Z(n29731) );
  NAND U30354 ( .A(n36296), .B(n29731), .Z(n29571) );
  AND U30355 ( .A(n29572), .B(n29571), .Z(n29787) );
  NAND U30356 ( .A(n190), .B(n29573), .Z(n29575) );
  XOR U30357 ( .A(b[19]), .B(a[196]), .Z(n29734) );
  NAND U30358 ( .A(n37821), .B(n29734), .Z(n29574) );
  NAND U30359 ( .A(n29575), .B(n29574), .Z(n29786) );
  XNOR U30360 ( .A(n29787), .B(n29786), .Z(n29788) );
  XNOR U30361 ( .A(n29789), .B(n29788), .Z(n29780) );
  NAND U30362 ( .A(n38470), .B(n29576), .Z(n29578) );
  XOR U30363 ( .A(b[31]), .B(a[184]), .Z(n29737) );
  NAND U30364 ( .A(n38453), .B(n29737), .Z(n29577) );
  AND U30365 ( .A(n29578), .B(n29577), .Z(n29749) );
  NAND U30366 ( .A(n181), .B(n29579), .Z(n29581) );
  XOR U30367 ( .A(b[3]), .B(a[212]), .Z(n29740) );
  NAND U30368 ( .A(n182), .B(n29740), .Z(n29580) );
  AND U30369 ( .A(n29581), .B(n29580), .Z(n29747) );
  NAND U30370 ( .A(n189), .B(n29582), .Z(n29584) );
  XOR U30371 ( .A(b[17]), .B(a[198]), .Z(n29743) );
  NAND U30372 ( .A(n37652), .B(n29743), .Z(n29583) );
  NAND U30373 ( .A(n29584), .B(n29583), .Z(n29746) );
  XNOR U30374 ( .A(n29747), .B(n29746), .Z(n29748) );
  XOR U30375 ( .A(n29749), .B(n29748), .Z(n29781) );
  XOR U30376 ( .A(n29780), .B(n29781), .Z(n29783) );
  XOR U30377 ( .A(n29782), .B(n29783), .Z(n29717) );
  NANDN U30378 ( .A(n29586), .B(n29585), .Z(n29590) );
  NANDN U30379 ( .A(n29588), .B(n29587), .Z(n29589) );
  AND U30380 ( .A(n29590), .B(n29589), .Z(n29770) );
  NANDN U30381 ( .A(n29592), .B(n29591), .Z(n29596) );
  NANDN U30382 ( .A(n29594), .B(n29593), .Z(n29595) );
  NAND U30383 ( .A(n29596), .B(n29595), .Z(n29771) );
  XNOR U30384 ( .A(n29770), .B(n29771), .Z(n29772) );
  NANDN U30385 ( .A(n29598), .B(n29597), .Z(n29602) );
  NANDN U30386 ( .A(n29600), .B(n29599), .Z(n29601) );
  NAND U30387 ( .A(n29602), .B(n29601), .Z(n29773) );
  XNOR U30388 ( .A(n29772), .B(n29773), .Z(n29716) );
  XNOR U30389 ( .A(n29717), .B(n29716), .Z(n29719) );
  NANDN U30390 ( .A(n29604), .B(n29603), .Z(n29608) );
  NANDN U30391 ( .A(n29606), .B(n29605), .Z(n29607) );
  AND U30392 ( .A(n29608), .B(n29607), .Z(n29718) );
  XOR U30393 ( .A(n29719), .B(n29718), .Z(n29830) );
  NANDN U30394 ( .A(n29610), .B(n29609), .Z(n29614) );
  NANDN U30395 ( .A(n29612), .B(n29611), .Z(n29613) );
  AND U30396 ( .A(n29614), .B(n29613), .Z(n29828) );
  NANDN U30397 ( .A(n29616), .B(n29615), .Z(n29620) );
  NANDN U30398 ( .A(n29618), .B(n29617), .Z(n29619) );
  AND U30399 ( .A(n29620), .B(n29619), .Z(n29713) );
  NANDN U30400 ( .A(n29622), .B(n29621), .Z(n29626) );
  OR U30401 ( .A(n29624), .B(n29623), .Z(n29625) );
  AND U30402 ( .A(n29626), .B(n29625), .Z(n29711) );
  NANDN U30403 ( .A(n29628), .B(n29627), .Z(n29632) );
  NANDN U30404 ( .A(n29630), .B(n29629), .Z(n29631) );
  AND U30405 ( .A(n29632), .B(n29631), .Z(n29777) );
  NANDN U30406 ( .A(n29634), .B(n29633), .Z(n29638) );
  NANDN U30407 ( .A(n29636), .B(n29635), .Z(n29637) );
  NAND U30408 ( .A(n29638), .B(n29637), .Z(n29776) );
  XNOR U30409 ( .A(n29777), .B(n29776), .Z(n29779) );
  NAND U30410 ( .A(b[0]), .B(a[214]), .Z(n29639) );
  XNOR U30411 ( .A(b[1]), .B(n29639), .Z(n29641) );
  NANDN U30412 ( .A(b[0]), .B(a[213]), .Z(n29640) );
  NAND U30413 ( .A(n29641), .B(n29640), .Z(n29725) );
  NAND U30414 ( .A(n194), .B(n29642), .Z(n29644) );
  XOR U30415 ( .A(b[29]), .B(a[186]), .Z(n29798) );
  NAND U30416 ( .A(n38456), .B(n29798), .Z(n29643) );
  AND U30417 ( .A(n29644), .B(n29643), .Z(n29723) );
  AND U30418 ( .A(b[31]), .B(a[182]), .Z(n29722) );
  XNOR U30419 ( .A(n29723), .B(n29722), .Z(n29724) );
  XNOR U30420 ( .A(n29725), .B(n29724), .Z(n29765) );
  NAND U30421 ( .A(n38185), .B(n29645), .Z(n29647) );
  XOR U30422 ( .A(b[23]), .B(a[192]), .Z(n29804) );
  NAND U30423 ( .A(n38132), .B(n29804), .Z(n29646) );
  AND U30424 ( .A(n29647), .B(n29646), .Z(n29794) );
  NAND U30425 ( .A(n184), .B(n29648), .Z(n29650) );
  XOR U30426 ( .A(b[7]), .B(a[208]), .Z(n29807) );
  NAND U30427 ( .A(n36592), .B(n29807), .Z(n29649) );
  AND U30428 ( .A(n29650), .B(n29649), .Z(n29793) );
  NAND U30429 ( .A(n38289), .B(n29651), .Z(n29653) );
  XOR U30430 ( .A(b[25]), .B(a[190]), .Z(n29810) );
  NAND U30431 ( .A(n38247), .B(n29810), .Z(n29652) );
  NAND U30432 ( .A(n29653), .B(n29652), .Z(n29792) );
  XOR U30433 ( .A(n29793), .B(n29792), .Z(n29795) );
  XOR U30434 ( .A(n29794), .B(n29795), .Z(n29764) );
  XOR U30435 ( .A(n29765), .B(n29764), .Z(n29767) );
  NAND U30436 ( .A(n187), .B(n29654), .Z(n29656) );
  XOR U30437 ( .A(b[13]), .B(a[202]), .Z(n29813) );
  NAND U30438 ( .A(n37295), .B(n29813), .Z(n29655) );
  AND U30439 ( .A(n29656), .B(n29655), .Z(n29759) );
  NAND U30440 ( .A(n186), .B(n29657), .Z(n29659) );
  XOR U30441 ( .A(b[11]), .B(a[204]), .Z(n29816) );
  NAND U30442 ( .A(n37097), .B(n29816), .Z(n29658) );
  NAND U30443 ( .A(n29659), .B(n29658), .Z(n29758) );
  XNOR U30444 ( .A(n29759), .B(n29758), .Z(n29761) );
  NAND U30445 ( .A(n188), .B(n29660), .Z(n29662) );
  XOR U30446 ( .A(b[15]), .B(a[200]), .Z(n29819) );
  NAND U30447 ( .A(n37382), .B(n29819), .Z(n29661) );
  AND U30448 ( .A(n29662), .B(n29661), .Z(n29755) );
  NAND U30449 ( .A(n38064), .B(n29663), .Z(n29665) );
  XOR U30450 ( .A(b[21]), .B(a[194]), .Z(n29822) );
  NAND U30451 ( .A(n37993), .B(n29822), .Z(n29664) );
  AND U30452 ( .A(n29665), .B(n29664), .Z(n29753) );
  NAND U30453 ( .A(n185), .B(n29666), .Z(n29668) );
  XOR U30454 ( .A(b[9]), .B(a[206]), .Z(n29825) );
  NAND U30455 ( .A(n36805), .B(n29825), .Z(n29667) );
  NAND U30456 ( .A(n29668), .B(n29667), .Z(n29752) );
  XNOR U30457 ( .A(n29753), .B(n29752), .Z(n29754) );
  XNOR U30458 ( .A(n29755), .B(n29754), .Z(n29760) );
  XOR U30459 ( .A(n29761), .B(n29760), .Z(n29766) );
  XNOR U30460 ( .A(n29767), .B(n29766), .Z(n29778) );
  XNOR U30461 ( .A(n29779), .B(n29778), .Z(n29710) );
  XNOR U30462 ( .A(n29711), .B(n29710), .Z(n29712) );
  XOR U30463 ( .A(n29713), .B(n29712), .Z(n29829) );
  XOR U30464 ( .A(n29828), .B(n29829), .Z(n29831) );
  XOR U30465 ( .A(n29830), .B(n29831), .Z(n29707) );
  NANDN U30466 ( .A(n29670), .B(n29669), .Z(n29674) );
  NAND U30467 ( .A(n29672), .B(n29671), .Z(n29673) );
  AND U30468 ( .A(n29674), .B(n29673), .Z(n29705) );
  NANDN U30469 ( .A(n29676), .B(n29675), .Z(n29680) );
  NANDN U30470 ( .A(n29678), .B(n29677), .Z(n29679) );
  AND U30471 ( .A(n29680), .B(n29679), .Z(n29704) );
  XNOR U30472 ( .A(n29705), .B(n29704), .Z(n29706) );
  XNOR U30473 ( .A(n29707), .B(n29706), .Z(n29698) );
  NANDN U30474 ( .A(n29682), .B(n29681), .Z(n29686) );
  OR U30475 ( .A(n29684), .B(n29683), .Z(n29685) );
  NAND U30476 ( .A(n29686), .B(n29685), .Z(n29699) );
  XNOR U30477 ( .A(n29698), .B(n29699), .Z(n29700) );
  XNOR U30478 ( .A(n29701), .B(n29700), .Z(n29692) );
  XNOR U30479 ( .A(n29693), .B(n29692), .Z(n29694) );
  XNOR U30480 ( .A(n29695), .B(n29694), .Z(n29834) );
  XNOR U30481 ( .A(sreg[438]), .B(n29834), .Z(n29836) );
  NANDN U30482 ( .A(sreg[437]), .B(n29687), .Z(n29691) );
  NAND U30483 ( .A(n29689), .B(n29688), .Z(n29690) );
  NAND U30484 ( .A(n29691), .B(n29690), .Z(n29835) );
  XNOR U30485 ( .A(n29836), .B(n29835), .Z(c[438]) );
  NANDN U30486 ( .A(n29693), .B(n29692), .Z(n29697) );
  NANDN U30487 ( .A(n29695), .B(n29694), .Z(n29696) );
  AND U30488 ( .A(n29697), .B(n29696), .Z(n29842) );
  NANDN U30489 ( .A(n29699), .B(n29698), .Z(n29703) );
  NANDN U30490 ( .A(n29701), .B(n29700), .Z(n29702) );
  AND U30491 ( .A(n29703), .B(n29702), .Z(n29840) );
  NANDN U30492 ( .A(n29705), .B(n29704), .Z(n29709) );
  NANDN U30493 ( .A(n29707), .B(n29706), .Z(n29708) );
  AND U30494 ( .A(n29709), .B(n29708), .Z(n29848) );
  NANDN U30495 ( .A(n29711), .B(n29710), .Z(n29715) );
  NANDN U30496 ( .A(n29713), .B(n29712), .Z(n29714) );
  AND U30497 ( .A(n29715), .B(n29714), .Z(n29852) );
  NANDN U30498 ( .A(n29717), .B(n29716), .Z(n29721) );
  NAND U30499 ( .A(n29719), .B(n29718), .Z(n29720) );
  AND U30500 ( .A(n29721), .B(n29720), .Z(n29851) );
  XNOR U30501 ( .A(n29852), .B(n29851), .Z(n29854) );
  NANDN U30502 ( .A(n29723), .B(n29722), .Z(n29727) );
  NANDN U30503 ( .A(n29725), .B(n29724), .Z(n29726) );
  AND U30504 ( .A(n29727), .B(n29726), .Z(n29919) );
  NAND U30505 ( .A(n38385), .B(n29728), .Z(n29730) );
  XOR U30506 ( .A(b[27]), .B(a[189]), .Z(n29863) );
  NAND U30507 ( .A(n38343), .B(n29863), .Z(n29729) );
  AND U30508 ( .A(n29730), .B(n29729), .Z(n29926) );
  NAND U30509 ( .A(n183), .B(n29731), .Z(n29733) );
  XOR U30510 ( .A(b[5]), .B(a[211]), .Z(n29866) );
  NAND U30511 ( .A(n36296), .B(n29866), .Z(n29732) );
  AND U30512 ( .A(n29733), .B(n29732), .Z(n29924) );
  NAND U30513 ( .A(n190), .B(n29734), .Z(n29736) );
  XOR U30514 ( .A(b[19]), .B(a[197]), .Z(n29869) );
  NAND U30515 ( .A(n37821), .B(n29869), .Z(n29735) );
  NAND U30516 ( .A(n29736), .B(n29735), .Z(n29923) );
  XNOR U30517 ( .A(n29924), .B(n29923), .Z(n29925) );
  XNOR U30518 ( .A(n29926), .B(n29925), .Z(n29917) );
  NAND U30519 ( .A(n38470), .B(n29737), .Z(n29739) );
  XOR U30520 ( .A(b[31]), .B(a[185]), .Z(n29872) );
  NAND U30521 ( .A(n38453), .B(n29872), .Z(n29738) );
  AND U30522 ( .A(n29739), .B(n29738), .Z(n29884) );
  NAND U30523 ( .A(n181), .B(n29740), .Z(n29742) );
  XOR U30524 ( .A(b[3]), .B(a[213]), .Z(n29875) );
  NAND U30525 ( .A(n182), .B(n29875), .Z(n29741) );
  AND U30526 ( .A(n29742), .B(n29741), .Z(n29882) );
  NAND U30527 ( .A(n189), .B(n29743), .Z(n29745) );
  XOR U30528 ( .A(b[17]), .B(a[199]), .Z(n29878) );
  NAND U30529 ( .A(n37652), .B(n29878), .Z(n29744) );
  NAND U30530 ( .A(n29745), .B(n29744), .Z(n29881) );
  XNOR U30531 ( .A(n29882), .B(n29881), .Z(n29883) );
  XOR U30532 ( .A(n29884), .B(n29883), .Z(n29918) );
  XOR U30533 ( .A(n29917), .B(n29918), .Z(n29920) );
  XOR U30534 ( .A(n29919), .B(n29920), .Z(n29966) );
  NANDN U30535 ( .A(n29747), .B(n29746), .Z(n29751) );
  NANDN U30536 ( .A(n29749), .B(n29748), .Z(n29750) );
  AND U30537 ( .A(n29751), .B(n29750), .Z(n29905) );
  NANDN U30538 ( .A(n29753), .B(n29752), .Z(n29757) );
  NANDN U30539 ( .A(n29755), .B(n29754), .Z(n29756) );
  NAND U30540 ( .A(n29757), .B(n29756), .Z(n29906) );
  XNOR U30541 ( .A(n29905), .B(n29906), .Z(n29907) );
  NANDN U30542 ( .A(n29759), .B(n29758), .Z(n29763) );
  NAND U30543 ( .A(n29761), .B(n29760), .Z(n29762) );
  NAND U30544 ( .A(n29763), .B(n29762), .Z(n29908) );
  XNOR U30545 ( .A(n29907), .B(n29908), .Z(n29965) );
  XNOR U30546 ( .A(n29966), .B(n29965), .Z(n29968) );
  NAND U30547 ( .A(n29765), .B(n29764), .Z(n29769) );
  NAND U30548 ( .A(n29767), .B(n29766), .Z(n29768) );
  AND U30549 ( .A(n29769), .B(n29768), .Z(n29967) );
  XOR U30550 ( .A(n29968), .B(n29967), .Z(n29980) );
  NANDN U30551 ( .A(n29771), .B(n29770), .Z(n29775) );
  NANDN U30552 ( .A(n29773), .B(n29772), .Z(n29774) );
  AND U30553 ( .A(n29775), .B(n29774), .Z(n29977) );
  NANDN U30554 ( .A(n29781), .B(n29780), .Z(n29785) );
  OR U30555 ( .A(n29783), .B(n29782), .Z(n29784) );
  AND U30556 ( .A(n29785), .B(n29784), .Z(n29972) );
  NANDN U30557 ( .A(n29787), .B(n29786), .Z(n29791) );
  NANDN U30558 ( .A(n29789), .B(n29788), .Z(n29790) );
  AND U30559 ( .A(n29791), .B(n29790), .Z(n29912) );
  NANDN U30560 ( .A(n29793), .B(n29792), .Z(n29797) );
  OR U30561 ( .A(n29795), .B(n29794), .Z(n29796) );
  NAND U30562 ( .A(n29797), .B(n29796), .Z(n29911) );
  XNOR U30563 ( .A(n29912), .B(n29911), .Z(n29913) );
  NAND U30564 ( .A(n194), .B(n29798), .Z(n29800) );
  XOR U30565 ( .A(b[29]), .B(a[187]), .Z(n29938) );
  NAND U30566 ( .A(n38456), .B(n29938), .Z(n29799) );
  AND U30567 ( .A(n29800), .B(n29799), .Z(n29858) );
  AND U30568 ( .A(b[31]), .B(a[183]), .Z(n29857) );
  XNOR U30569 ( .A(n29858), .B(n29857), .Z(n29859) );
  NAND U30570 ( .A(b[0]), .B(a[215]), .Z(n29801) );
  XNOR U30571 ( .A(b[1]), .B(n29801), .Z(n29803) );
  NANDN U30572 ( .A(b[0]), .B(a[214]), .Z(n29802) );
  NAND U30573 ( .A(n29803), .B(n29802), .Z(n29860) );
  XNOR U30574 ( .A(n29859), .B(n29860), .Z(n29899) );
  NAND U30575 ( .A(n38185), .B(n29804), .Z(n29806) );
  XOR U30576 ( .A(b[23]), .B(a[193]), .Z(n29941) );
  NAND U30577 ( .A(n38132), .B(n29941), .Z(n29805) );
  AND U30578 ( .A(n29806), .B(n29805), .Z(n29932) );
  NAND U30579 ( .A(n184), .B(n29807), .Z(n29809) );
  XOR U30580 ( .A(b[7]), .B(a[209]), .Z(n29944) );
  NAND U30581 ( .A(n36592), .B(n29944), .Z(n29808) );
  AND U30582 ( .A(n29809), .B(n29808), .Z(n29930) );
  NAND U30583 ( .A(n38289), .B(n29810), .Z(n29812) );
  XOR U30584 ( .A(b[25]), .B(a[191]), .Z(n29947) );
  NAND U30585 ( .A(n38247), .B(n29947), .Z(n29811) );
  NAND U30586 ( .A(n29812), .B(n29811), .Z(n29929) );
  XNOR U30587 ( .A(n29930), .B(n29929), .Z(n29931) );
  XOR U30588 ( .A(n29932), .B(n29931), .Z(n29900) );
  XNOR U30589 ( .A(n29899), .B(n29900), .Z(n29901) );
  NAND U30590 ( .A(n187), .B(n29813), .Z(n29815) );
  XOR U30591 ( .A(b[13]), .B(a[203]), .Z(n29950) );
  NAND U30592 ( .A(n37295), .B(n29950), .Z(n29814) );
  AND U30593 ( .A(n29815), .B(n29814), .Z(n29894) );
  NAND U30594 ( .A(n186), .B(n29816), .Z(n29818) );
  XOR U30595 ( .A(b[11]), .B(a[205]), .Z(n29953) );
  NAND U30596 ( .A(n37097), .B(n29953), .Z(n29817) );
  NAND U30597 ( .A(n29818), .B(n29817), .Z(n29893) );
  XNOR U30598 ( .A(n29894), .B(n29893), .Z(n29895) );
  NAND U30599 ( .A(n188), .B(n29819), .Z(n29821) );
  XOR U30600 ( .A(b[15]), .B(a[201]), .Z(n29956) );
  NAND U30601 ( .A(n37382), .B(n29956), .Z(n29820) );
  AND U30602 ( .A(n29821), .B(n29820), .Z(n29890) );
  NAND U30603 ( .A(n38064), .B(n29822), .Z(n29824) );
  XOR U30604 ( .A(b[21]), .B(a[195]), .Z(n29959) );
  NAND U30605 ( .A(n37993), .B(n29959), .Z(n29823) );
  AND U30606 ( .A(n29824), .B(n29823), .Z(n29888) );
  NAND U30607 ( .A(n185), .B(n29825), .Z(n29827) );
  XOR U30608 ( .A(b[9]), .B(a[207]), .Z(n29962) );
  NAND U30609 ( .A(n36805), .B(n29962), .Z(n29826) );
  NAND U30610 ( .A(n29827), .B(n29826), .Z(n29887) );
  XNOR U30611 ( .A(n29888), .B(n29887), .Z(n29889) );
  XOR U30612 ( .A(n29890), .B(n29889), .Z(n29896) );
  XOR U30613 ( .A(n29895), .B(n29896), .Z(n29902) );
  XOR U30614 ( .A(n29901), .B(n29902), .Z(n29914) );
  XNOR U30615 ( .A(n29913), .B(n29914), .Z(n29971) );
  XNOR U30616 ( .A(n29972), .B(n29971), .Z(n29973) );
  XOR U30617 ( .A(n29974), .B(n29973), .Z(n29978) );
  XNOR U30618 ( .A(n29977), .B(n29978), .Z(n29979) );
  XNOR U30619 ( .A(n29980), .B(n29979), .Z(n29853) );
  XOR U30620 ( .A(n29854), .B(n29853), .Z(n29846) );
  NANDN U30621 ( .A(n29829), .B(n29828), .Z(n29833) );
  OR U30622 ( .A(n29831), .B(n29830), .Z(n29832) );
  AND U30623 ( .A(n29833), .B(n29832), .Z(n29845) );
  XNOR U30624 ( .A(n29846), .B(n29845), .Z(n29847) );
  XNOR U30625 ( .A(n29848), .B(n29847), .Z(n29839) );
  XNOR U30626 ( .A(n29840), .B(n29839), .Z(n29841) );
  XNOR U30627 ( .A(n29842), .B(n29841), .Z(n29983) );
  XNOR U30628 ( .A(sreg[439]), .B(n29983), .Z(n29985) );
  NANDN U30629 ( .A(sreg[438]), .B(n29834), .Z(n29838) );
  NAND U30630 ( .A(n29836), .B(n29835), .Z(n29837) );
  NAND U30631 ( .A(n29838), .B(n29837), .Z(n29984) );
  XNOR U30632 ( .A(n29985), .B(n29984), .Z(c[439]) );
  NANDN U30633 ( .A(n29840), .B(n29839), .Z(n29844) );
  NANDN U30634 ( .A(n29842), .B(n29841), .Z(n29843) );
  AND U30635 ( .A(n29844), .B(n29843), .Z(n29991) );
  NANDN U30636 ( .A(n29846), .B(n29845), .Z(n29850) );
  NANDN U30637 ( .A(n29848), .B(n29847), .Z(n29849) );
  AND U30638 ( .A(n29850), .B(n29849), .Z(n29989) );
  NANDN U30639 ( .A(n29852), .B(n29851), .Z(n29856) );
  NAND U30640 ( .A(n29854), .B(n29853), .Z(n29855) );
  AND U30641 ( .A(n29856), .B(n29855), .Z(n29996) );
  NANDN U30642 ( .A(n29858), .B(n29857), .Z(n29862) );
  NANDN U30643 ( .A(n29860), .B(n29859), .Z(n29861) );
  AND U30644 ( .A(n29862), .B(n29861), .Z(n30080) );
  NAND U30645 ( .A(n38385), .B(n29863), .Z(n29865) );
  XOR U30646 ( .A(b[27]), .B(a[190]), .Z(n30024) );
  NAND U30647 ( .A(n38343), .B(n30024), .Z(n29864) );
  AND U30648 ( .A(n29865), .B(n29864), .Z(n30087) );
  NAND U30649 ( .A(n183), .B(n29866), .Z(n29868) );
  XOR U30650 ( .A(b[5]), .B(a[212]), .Z(n30027) );
  NAND U30651 ( .A(n36296), .B(n30027), .Z(n29867) );
  AND U30652 ( .A(n29868), .B(n29867), .Z(n30085) );
  NAND U30653 ( .A(n190), .B(n29869), .Z(n29871) );
  XOR U30654 ( .A(b[19]), .B(a[198]), .Z(n30030) );
  NAND U30655 ( .A(n37821), .B(n30030), .Z(n29870) );
  NAND U30656 ( .A(n29871), .B(n29870), .Z(n30084) );
  XNOR U30657 ( .A(n30085), .B(n30084), .Z(n30086) );
  XNOR U30658 ( .A(n30087), .B(n30086), .Z(n30078) );
  NAND U30659 ( .A(n38470), .B(n29872), .Z(n29874) );
  XOR U30660 ( .A(b[31]), .B(a[186]), .Z(n30033) );
  NAND U30661 ( .A(n38453), .B(n30033), .Z(n29873) );
  AND U30662 ( .A(n29874), .B(n29873), .Z(n30045) );
  NAND U30663 ( .A(n181), .B(n29875), .Z(n29877) );
  XOR U30664 ( .A(b[3]), .B(a[214]), .Z(n30036) );
  NAND U30665 ( .A(n182), .B(n30036), .Z(n29876) );
  AND U30666 ( .A(n29877), .B(n29876), .Z(n30043) );
  NAND U30667 ( .A(n189), .B(n29878), .Z(n29880) );
  XOR U30668 ( .A(b[17]), .B(a[200]), .Z(n30039) );
  NAND U30669 ( .A(n37652), .B(n30039), .Z(n29879) );
  NAND U30670 ( .A(n29880), .B(n29879), .Z(n30042) );
  XNOR U30671 ( .A(n30043), .B(n30042), .Z(n30044) );
  XOR U30672 ( .A(n30045), .B(n30044), .Z(n30079) );
  XOR U30673 ( .A(n30078), .B(n30079), .Z(n30081) );
  XOR U30674 ( .A(n30080), .B(n30081), .Z(n30013) );
  NANDN U30675 ( .A(n29882), .B(n29881), .Z(n29886) );
  NANDN U30676 ( .A(n29884), .B(n29883), .Z(n29885) );
  AND U30677 ( .A(n29886), .B(n29885), .Z(n30066) );
  NANDN U30678 ( .A(n29888), .B(n29887), .Z(n29892) );
  NANDN U30679 ( .A(n29890), .B(n29889), .Z(n29891) );
  NAND U30680 ( .A(n29892), .B(n29891), .Z(n30067) );
  XNOR U30681 ( .A(n30066), .B(n30067), .Z(n30068) );
  NANDN U30682 ( .A(n29894), .B(n29893), .Z(n29898) );
  NANDN U30683 ( .A(n29896), .B(n29895), .Z(n29897) );
  NAND U30684 ( .A(n29898), .B(n29897), .Z(n30069) );
  XNOR U30685 ( .A(n30068), .B(n30069), .Z(n30012) );
  XNOR U30686 ( .A(n30013), .B(n30012), .Z(n30015) );
  NANDN U30687 ( .A(n29900), .B(n29899), .Z(n29904) );
  NANDN U30688 ( .A(n29902), .B(n29901), .Z(n29903) );
  AND U30689 ( .A(n29904), .B(n29903), .Z(n30014) );
  XOR U30690 ( .A(n30015), .B(n30014), .Z(n30128) );
  NANDN U30691 ( .A(n29906), .B(n29905), .Z(n29910) );
  NANDN U30692 ( .A(n29908), .B(n29907), .Z(n29909) );
  AND U30693 ( .A(n29910), .B(n29909), .Z(n30126) );
  NANDN U30694 ( .A(n29912), .B(n29911), .Z(n29916) );
  NANDN U30695 ( .A(n29914), .B(n29913), .Z(n29915) );
  AND U30696 ( .A(n29916), .B(n29915), .Z(n30009) );
  NANDN U30697 ( .A(n29918), .B(n29917), .Z(n29922) );
  OR U30698 ( .A(n29920), .B(n29919), .Z(n29921) );
  AND U30699 ( .A(n29922), .B(n29921), .Z(n30007) );
  NANDN U30700 ( .A(n29924), .B(n29923), .Z(n29928) );
  NANDN U30701 ( .A(n29926), .B(n29925), .Z(n29927) );
  AND U30702 ( .A(n29928), .B(n29927), .Z(n30073) );
  NANDN U30703 ( .A(n29930), .B(n29929), .Z(n29934) );
  NANDN U30704 ( .A(n29932), .B(n29931), .Z(n29933) );
  NAND U30705 ( .A(n29934), .B(n29933), .Z(n30072) );
  XNOR U30706 ( .A(n30073), .B(n30072), .Z(n30074) );
  NAND U30707 ( .A(b[0]), .B(a[216]), .Z(n29935) );
  XNOR U30708 ( .A(b[1]), .B(n29935), .Z(n29937) );
  NANDN U30709 ( .A(b[0]), .B(a[215]), .Z(n29936) );
  NAND U30710 ( .A(n29937), .B(n29936), .Z(n30021) );
  NAND U30711 ( .A(n194), .B(n29938), .Z(n29940) );
  XOR U30712 ( .A(b[29]), .B(a[188]), .Z(n30099) );
  NAND U30713 ( .A(n38456), .B(n30099), .Z(n29939) );
  AND U30714 ( .A(n29940), .B(n29939), .Z(n30019) );
  AND U30715 ( .A(b[31]), .B(a[184]), .Z(n30018) );
  XNOR U30716 ( .A(n30019), .B(n30018), .Z(n30020) );
  XNOR U30717 ( .A(n30021), .B(n30020), .Z(n30060) );
  NAND U30718 ( .A(n38185), .B(n29941), .Z(n29943) );
  XOR U30719 ( .A(b[23]), .B(a[194]), .Z(n30102) );
  NAND U30720 ( .A(n38132), .B(n30102), .Z(n29942) );
  AND U30721 ( .A(n29943), .B(n29942), .Z(n30093) );
  NAND U30722 ( .A(n184), .B(n29944), .Z(n29946) );
  XOR U30723 ( .A(b[7]), .B(a[210]), .Z(n30105) );
  NAND U30724 ( .A(n36592), .B(n30105), .Z(n29945) );
  AND U30725 ( .A(n29946), .B(n29945), .Z(n30091) );
  NAND U30726 ( .A(n38289), .B(n29947), .Z(n29949) );
  XOR U30727 ( .A(b[25]), .B(a[192]), .Z(n30108) );
  NAND U30728 ( .A(n38247), .B(n30108), .Z(n29948) );
  NAND U30729 ( .A(n29949), .B(n29948), .Z(n30090) );
  XNOR U30730 ( .A(n30091), .B(n30090), .Z(n30092) );
  XOR U30731 ( .A(n30093), .B(n30092), .Z(n30061) );
  XNOR U30732 ( .A(n30060), .B(n30061), .Z(n30062) );
  NAND U30733 ( .A(n187), .B(n29950), .Z(n29952) );
  XOR U30734 ( .A(b[13]), .B(a[204]), .Z(n30111) );
  NAND U30735 ( .A(n37295), .B(n30111), .Z(n29951) );
  AND U30736 ( .A(n29952), .B(n29951), .Z(n30055) );
  NAND U30737 ( .A(n186), .B(n29953), .Z(n29955) );
  XOR U30738 ( .A(b[11]), .B(a[206]), .Z(n30114) );
  NAND U30739 ( .A(n37097), .B(n30114), .Z(n29954) );
  NAND U30740 ( .A(n29955), .B(n29954), .Z(n30054) );
  XNOR U30741 ( .A(n30055), .B(n30054), .Z(n30056) );
  NAND U30742 ( .A(n188), .B(n29956), .Z(n29958) );
  XOR U30743 ( .A(b[15]), .B(a[202]), .Z(n30117) );
  NAND U30744 ( .A(n37382), .B(n30117), .Z(n29957) );
  AND U30745 ( .A(n29958), .B(n29957), .Z(n30051) );
  NAND U30746 ( .A(n38064), .B(n29959), .Z(n29961) );
  XOR U30747 ( .A(b[21]), .B(a[196]), .Z(n30120) );
  NAND U30748 ( .A(n37993), .B(n30120), .Z(n29960) );
  AND U30749 ( .A(n29961), .B(n29960), .Z(n30049) );
  NAND U30750 ( .A(n185), .B(n29962), .Z(n29964) );
  XOR U30751 ( .A(b[9]), .B(a[208]), .Z(n30123) );
  NAND U30752 ( .A(n36805), .B(n30123), .Z(n29963) );
  NAND U30753 ( .A(n29964), .B(n29963), .Z(n30048) );
  XNOR U30754 ( .A(n30049), .B(n30048), .Z(n30050) );
  XOR U30755 ( .A(n30051), .B(n30050), .Z(n30057) );
  XOR U30756 ( .A(n30056), .B(n30057), .Z(n30063) );
  XOR U30757 ( .A(n30062), .B(n30063), .Z(n30075) );
  XNOR U30758 ( .A(n30074), .B(n30075), .Z(n30006) );
  XNOR U30759 ( .A(n30007), .B(n30006), .Z(n30008) );
  XOR U30760 ( .A(n30009), .B(n30008), .Z(n30127) );
  XOR U30761 ( .A(n30126), .B(n30127), .Z(n30129) );
  XOR U30762 ( .A(n30128), .B(n30129), .Z(n30003) );
  NANDN U30763 ( .A(n29966), .B(n29965), .Z(n29970) );
  NAND U30764 ( .A(n29968), .B(n29967), .Z(n29969) );
  AND U30765 ( .A(n29970), .B(n29969), .Z(n30001) );
  NANDN U30766 ( .A(n29972), .B(n29971), .Z(n29976) );
  NANDN U30767 ( .A(n29974), .B(n29973), .Z(n29975) );
  AND U30768 ( .A(n29976), .B(n29975), .Z(n30000) );
  XNOR U30769 ( .A(n30001), .B(n30000), .Z(n30002) );
  XNOR U30770 ( .A(n30003), .B(n30002), .Z(n29994) );
  NANDN U30771 ( .A(n29978), .B(n29977), .Z(n29982) );
  NANDN U30772 ( .A(n29980), .B(n29979), .Z(n29981) );
  NAND U30773 ( .A(n29982), .B(n29981), .Z(n29995) );
  XOR U30774 ( .A(n29994), .B(n29995), .Z(n29997) );
  XNOR U30775 ( .A(n29996), .B(n29997), .Z(n29988) );
  XNOR U30776 ( .A(n29989), .B(n29988), .Z(n29990) );
  XNOR U30777 ( .A(n29991), .B(n29990), .Z(n30132) );
  XNOR U30778 ( .A(sreg[440]), .B(n30132), .Z(n30134) );
  NANDN U30779 ( .A(sreg[439]), .B(n29983), .Z(n29987) );
  NAND U30780 ( .A(n29985), .B(n29984), .Z(n29986) );
  NAND U30781 ( .A(n29987), .B(n29986), .Z(n30133) );
  XNOR U30782 ( .A(n30134), .B(n30133), .Z(c[440]) );
  NANDN U30783 ( .A(n29989), .B(n29988), .Z(n29993) );
  NANDN U30784 ( .A(n29991), .B(n29990), .Z(n29992) );
  AND U30785 ( .A(n29993), .B(n29992), .Z(n30140) );
  NANDN U30786 ( .A(n29995), .B(n29994), .Z(n29999) );
  NANDN U30787 ( .A(n29997), .B(n29996), .Z(n29998) );
  AND U30788 ( .A(n29999), .B(n29998), .Z(n30138) );
  NANDN U30789 ( .A(n30001), .B(n30000), .Z(n30005) );
  NANDN U30790 ( .A(n30003), .B(n30002), .Z(n30004) );
  AND U30791 ( .A(n30005), .B(n30004), .Z(n30146) );
  NANDN U30792 ( .A(n30007), .B(n30006), .Z(n30011) );
  NANDN U30793 ( .A(n30009), .B(n30008), .Z(n30010) );
  AND U30794 ( .A(n30011), .B(n30010), .Z(n30150) );
  NANDN U30795 ( .A(n30013), .B(n30012), .Z(n30017) );
  NAND U30796 ( .A(n30015), .B(n30014), .Z(n30016) );
  AND U30797 ( .A(n30017), .B(n30016), .Z(n30149) );
  XNOR U30798 ( .A(n30150), .B(n30149), .Z(n30152) );
  NANDN U30799 ( .A(n30019), .B(n30018), .Z(n30023) );
  NANDN U30800 ( .A(n30021), .B(n30020), .Z(n30022) );
  AND U30801 ( .A(n30023), .B(n30022), .Z(n30229) );
  NAND U30802 ( .A(n38385), .B(n30024), .Z(n30026) );
  XOR U30803 ( .A(b[27]), .B(a[191]), .Z(n30173) );
  NAND U30804 ( .A(n38343), .B(n30173), .Z(n30025) );
  AND U30805 ( .A(n30026), .B(n30025), .Z(n30236) );
  NAND U30806 ( .A(n183), .B(n30027), .Z(n30029) );
  XOR U30807 ( .A(b[5]), .B(a[213]), .Z(n30176) );
  NAND U30808 ( .A(n36296), .B(n30176), .Z(n30028) );
  AND U30809 ( .A(n30029), .B(n30028), .Z(n30234) );
  NAND U30810 ( .A(n190), .B(n30030), .Z(n30032) );
  XOR U30811 ( .A(b[19]), .B(a[199]), .Z(n30179) );
  NAND U30812 ( .A(n37821), .B(n30179), .Z(n30031) );
  NAND U30813 ( .A(n30032), .B(n30031), .Z(n30233) );
  XNOR U30814 ( .A(n30234), .B(n30233), .Z(n30235) );
  XNOR U30815 ( .A(n30236), .B(n30235), .Z(n30227) );
  NAND U30816 ( .A(n38470), .B(n30033), .Z(n30035) );
  XOR U30817 ( .A(b[31]), .B(a[187]), .Z(n30182) );
  NAND U30818 ( .A(n38453), .B(n30182), .Z(n30034) );
  AND U30819 ( .A(n30035), .B(n30034), .Z(n30194) );
  NAND U30820 ( .A(n181), .B(n30036), .Z(n30038) );
  XOR U30821 ( .A(b[3]), .B(a[215]), .Z(n30185) );
  NAND U30822 ( .A(n182), .B(n30185), .Z(n30037) );
  AND U30823 ( .A(n30038), .B(n30037), .Z(n30192) );
  NAND U30824 ( .A(n189), .B(n30039), .Z(n30041) );
  XOR U30825 ( .A(b[17]), .B(a[201]), .Z(n30188) );
  NAND U30826 ( .A(n37652), .B(n30188), .Z(n30040) );
  NAND U30827 ( .A(n30041), .B(n30040), .Z(n30191) );
  XNOR U30828 ( .A(n30192), .B(n30191), .Z(n30193) );
  XOR U30829 ( .A(n30194), .B(n30193), .Z(n30228) );
  XOR U30830 ( .A(n30227), .B(n30228), .Z(n30230) );
  XOR U30831 ( .A(n30229), .B(n30230), .Z(n30162) );
  NANDN U30832 ( .A(n30043), .B(n30042), .Z(n30047) );
  NANDN U30833 ( .A(n30045), .B(n30044), .Z(n30046) );
  AND U30834 ( .A(n30047), .B(n30046), .Z(n30215) );
  NANDN U30835 ( .A(n30049), .B(n30048), .Z(n30053) );
  NANDN U30836 ( .A(n30051), .B(n30050), .Z(n30052) );
  NAND U30837 ( .A(n30053), .B(n30052), .Z(n30216) );
  XNOR U30838 ( .A(n30215), .B(n30216), .Z(n30217) );
  NANDN U30839 ( .A(n30055), .B(n30054), .Z(n30059) );
  NANDN U30840 ( .A(n30057), .B(n30056), .Z(n30058) );
  NAND U30841 ( .A(n30059), .B(n30058), .Z(n30218) );
  XNOR U30842 ( .A(n30217), .B(n30218), .Z(n30161) );
  XNOR U30843 ( .A(n30162), .B(n30161), .Z(n30164) );
  NANDN U30844 ( .A(n30061), .B(n30060), .Z(n30065) );
  NANDN U30845 ( .A(n30063), .B(n30062), .Z(n30064) );
  AND U30846 ( .A(n30065), .B(n30064), .Z(n30163) );
  XOR U30847 ( .A(n30164), .B(n30163), .Z(n30278) );
  NANDN U30848 ( .A(n30067), .B(n30066), .Z(n30071) );
  NANDN U30849 ( .A(n30069), .B(n30068), .Z(n30070) );
  AND U30850 ( .A(n30071), .B(n30070), .Z(n30275) );
  NANDN U30851 ( .A(n30073), .B(n30072), .Z(n30077) );
  NANDN U30852 ( .A(n30075), .B(n30074), .Z(n30076) );
  AND U30853 ( .A(n30077), .B(n30076), .Z(n30158) );
  NANDN U30854 ( .A(n30079), .B(n30078), .Z(n30083) );
  OR U30855 ( .A(n30081), .B(n30080), .Z(n30082) );
  AND U30856 ( .A(n30083), .B(n30082), .Z(n30156) );
  NANDN U30857 ( .A(n30085), .B(n30084), .Z(n30089) );
  NANDN U30858 ( .A(n30087), .B(n30086), .Z(n30088) );
  AND U30859 ( .A(n30089), .B(n30088), .Z(n30222) );
  NANDN U30860 ( .A(n30091), .B(n30090), .Z(n30095) );
  NANDN U30861 ( .A(n30093), .B(n30092), .Z(n30094) );
  NAND U30862 ( .A(n30095), .B(n30094), .Z(n30221) );
  XNOR U30863 ( .A(n30222), .B(n30221), .Z(n30223) );
  NAND U30864 ( .A(b[0]), .B(a[217]), .Z(n30096) );
  XNOR U30865 ( .A(b[1]), .B(n30096), .Z(n30098) );
  NANDN U30866 ( .A(b[0]), .B(a[216]), .Z(n30097) );
  NAND U30867 ( .A(n30098), .B(n30097), .Z(n30170) );
  NAND U30868 ( .A(n194), .B(n30099), .Z(n30101) );
  XOR U30869 ( .A(b[29]), .B(a[189]), .Z(n30248) );
  NAND U30870 ( .A(n38456), .B(n30248), .Z(n30100) );
  AND U30871 ( .A(n30101), .B(n30100), .Z(n30168) );
  AND U30872 ( .A(b[31]), .B(a[185]), .Z(n30167) );
  XNOR U30873 ( .A(n30168), .B(n30167), .Z(n30169) );
  XNOR U30874 ( .A(n30170), .B(n30169), .Z(n30209) );
  NAND U30875 ( .A(n38185), .B(n30102), .Z(n30104) );
  XOR U30876 ( .A(b[23]), .B(a[195]), .Z(n30251) );
  NAND U30877 ( .A(n38132), .B(n30251), .Z(n30103) );
  AND U30878 ( .A(n30104), .B(n30103), .Z(n30242) );
  NAND U30879 ( .A(n184), .B(n30105), .Z(n30107) );
  XOR U30880 ( .A(b[7]), .B(a[211]), .Z(n30254) );
  NAND U30881 ( .A(n36592), .B(n30254), .Z(n30106) );
  AND U30882 ( .A(n30107), .B(n30106), .Z(n30240) );
  NAND U30883 ( .A(n38289), .B(n30108), .Z(n30110) );
  XOR U30884 ( .A(b[25]), .B(a[193]), .Z(n30257) );
  NAND U30885 ( .A(n38247), .B(n30257), .Z(n30109) );
  NAND U30886 ( .A(n30110), .B(n30109), .Z(n30239) );
  XNOR U30887 ( .A(n30240), .B(n30239), .Z(n30241) );
  XOR U30888 ( .A(n30242), .B(n30241), .Z(n30210) );
  XNOR U30889 ( .A(n30209), .B(n30210), .Z(n30211) );
  NAND U30890 ( .A(n187), .B(n30111), .Z(n30113) );
  XOR U30891 ( .A(b[13]), .B(a[205]), .Z(n30260) );
  NAND U30892 ( .A(n37295), .B(n30260), .Z(n30112) );
  AND U30893 ( .A(n30113), .B(n30112), .Z(n30204) );
  NAND U30894 ( .A(n186), .B(n30114), .Z(n30116) );
  XOR U30895 ( .A(b[11]), .B(a[207]), .Z(n30263) );
  NAND U30896 ( .A(n37097), .B(n30263), .Z(n30115) );
  NAND U30897 ( .A(n30116), .B(n30115), .Z(n30203) );
  XNOR U30898 ( .A(n30204), .B(n30203), .Z(n30205) );
  NAND U30899 ( .A(n188), .B(n30117), .Z(n30119) );
  XOR U30900 ( .A(b[15]), .B(a[203]), .Z(n30266) );
  NAND U30901 ( .A(n37382), .B(n30266), .Z(n30118) );
  AND U30902 ( .A(n30119), .B(n30118), .Z(n30200) );
  NAND U30903 ( .A(n38064), .B(n30120), .Z(n30122) );
  XOR U30904 ( .A(b[21]), .B(a[197]), .Z(n30269) );
  NAND U30905 ( .A(n37993), .B(n30269), .Z(n30121) );
  AND U30906 ( .A(n30122), .B(n30121), .Z(n30198) );
  NAND U30907 ( .A(n185), .B(n30123), .Z(n30125) );
  XOR U30908 ( .A(b[9]), .B(a[209]), .Z(n30272) );
  NAND U30909 ( .A(n36805), .B(n30272), .Z(n30124) );
  NAND U30910 ( .A(n30125), .B(n30124), .Z(n30197) );
  XNOR U30911 ( .A(n30198), .B(n30197), .Z(n30199) );
  XOR U30912 ( .A(n30200), .B(n30199), .Z(n30206) );
  XOR U30913 ( .A(n30205), .B(n30206), .Z(n30212) );
  XOR U30914 ( .A(n30211), .B(n30212), .Z(n30224) );
  XNOR U30915 ( .A(n30223), .B(n30224), .Z(n30155) );
  XNOR U30916 ( .A(n30156), .B(n30155), .Z(n30157) );
  XOR U30917 ( .A(n30158), .B(n30157), .Z(n30276) );
  XNOR U30918 ( .A(n30275), .B(n30276), .Z(n30277) );
  XNOR U30919 ( .A(n30278), .B(n30277), .Z(n30151) );
  XOR U30920 ( .A(n30152), .B(n30151), .Z(n30144) );
  NANDN U30921 ( .A(n30127), .B(n30126), .Z(n30131) );
  OR U30922 ( .A(n30129), .B(n30128), .Z(n30130) );
  AND U30923 ( .A(n30131), .B(n30130), .Z(n30143) );
  XNOR U30924 ( .A(n30144), .B(n30143), .Z(n30145) );
  XNOR U30925 ( .A(n30146), .B(n30145), .Z(n30137) );
  XNOR U30926 ( .A(n30138), .B(n30137), .Z(n30139) );
  XNOR U30927 ( .A(n30140), .B(n30139), .Z(n30281) );
  XNOR U30928 ( .A(sreg[441]), .B(n30281), .Z(n30283) );
  NANDN U30929 ( .A(sreg[440]), .B(n30132), .Z(n30136) );
  NAND U30930 ( .A(n30134), .B(n30133), .Z(n30135) );
  NAND U30931 ( .A(n30136), .B(n30135), .Z(n30282) );
  XNOR U30932 ( .A(n30283), .B(n30282), .Z(c[441]) );
  NANDN U30933 ( .A(n30138), .B(n30137), .Z(n30142) );
  NANDN U30934 ( .A(n30140), .B(n30139), .Z(n30141) );
  AND U30935 ( .A(n30142), .B(n30141), .Z(n30289) );
  NANDN U30936 ( .A(n30144), .B(n30143), .Z(n30148) );
  NANDN U30937 ( .A(n30146), .B(n30145), .Z(n30147) );
  AND U30938 ( .A(n30148), .B(n30147), .Z(n30287) );
  NANDN U30939 ( .A(n30150), .B(n30149), .Z(n30154) );
  NAND U30940 ( .A(n30152), .B(n30151), .Z(n30153) );
  AND U30941 ( .A(n30154), .B(n30153), .Z(n30294) );
  NANDN U30942 ( .A(n30156), .B(n30155), .Z(n30160) );
  NANDN U30943 ( .A(n30158), .B(n30157), .Z(n30159) );
  AND U30944 ( .A(n30160), .B(n30159), .Z(n30425) );
  NANDN U30945 ( .A(n30162), .B(n30161), .Z(n30166) );
  NAND U30946 ( .A(n30164), .B(n30163), .Z(n30165) );
  AND U30947 ( .A(n30166), .B(n30165), .Z(n30424) );
  XNOR U30948 ( .A(n30425), .B(n30424), .Z(n30427) );
  NANDN U30949 ( .A(n30168), .B(n30167), .Z(n30172) );
  NANDN U30950 ( .A(n30170), .B(n30169), .Z(n30171) );
  AND U30951 ( .A(n30172), .B(n30171), .Z(n30372) );
  NAND U30952 ( .A(n38385), .B(n30173), .Z(n30175) );
  XOR U30953 ( .A(b[27]), .B(a[192]), .Z(n30316) );
  NAND U30954 ( .A(n38343), .B(n30316), .Z(n30174) );
  AND U30955 ( .A(n30175), .B(n30174), .Z(n30379) );
  NAND U30956 ( .A(n183), .B(n30176), .Z(n30178) );
  XOR U30957 ( .A(b[5]), .B(a[214]), .Z(n30319) );
  NAND U30958 ( .A(n36296), .B(n30319), .Z(n30177) );
  AND U30959 ( .A(n30178), .B(n30177), .Z(n30377) );
  NAND U30960 ( .A(n190), .B(n30179), .Z(n30181) );
  XOR U30961 ( .A(b[19]), .B(a[200]), .Z(n30322) );
  NAND U30962 ( .A(n37821), .B(n30322), .Z(n30180) );
  NAND U30963 ( .A(n30181), .B(n30180), .Z(n30376) );
  XNOR U30964 ( .A(n30377), .B(n30376), .Z(n30378) );
  XNOR U30965 ( .A(n30379), .B(n30378), .Z(n30370) );
  NAND U30966 ( .A(n38470), .B(n30182), .Z(n30184) );
  XOR U30967 ( .A(b[31]), .B(a[188]), .Z(n30325) );
  NAND U30968 ( .A(n38453), .B(n30325), .Z(n30183) );
  AND U30969 ( .A(n30184), .B(n30183), .Z(n30337) );
  NAND U30970 ( .A(n181), .B(n30185), .Z(n30187) );
  XOR U30971 ( .A(b[3]), .B(a[216]), .Z(n30328) );
  NAND U30972 ( .A(n182), .B(n30328), .Z(n30186) );
  AND U30973 ( .A(n30187), .B(n30186), .Z(n30335) );
  NAND U30974 ( .A(n189), .B(n30188), .Z(n30190) );
  XOR U30975 ( .A(b[17]), .B(a[202]), .Z(n30331) );
  NAND U30976 ( .A(n37652), .B(n30331), .Z(n30189) );
  NAND U30977 ( .A(n30190), .B(n30189), .Z(n30334) );
  XNOR U30978 ( .A(n30335), .B(n30334), .Z(n30336) );
  XOR U30979 ( .A(n30337), .B(n30336), .Z(n30371) );
  XOR U30980 ( .A(n30370), .B(n30371), .Z(n30373) );
  XOR U30981 ( .A(n30372), .B(n30373), .Z(n30305) );
  NANDN U30982 ( .A(n30192), .B(n30191), .Z(n30196) );
  NANDN U30983 ( .A(n30194), .B(n30193), .Z(n30195) );
  AND U30984 ( .A(n30196), .B(n30195), .Z(n30358) );
  NANDN U30985 ( .A(n30198), .B(n30197), .Z(n30202) );
  NANDN U30986 ( .A(n30200), .B(n30199), .Z(n30201) );
  NAND U30987 ( .A(n30202), .B(n30201), .Z(n30359) );
  XNOR U30988 ( .A(n30358), .B(n30359), .Z(n30360) );
  NANDN U30989 ( .A(n30204), .B(n30203), .Z(n30208) );
  NANDN U30990 ( .A(n30206), .B(n30205), .Z(n30207) );
  NAND U30991 ( .A(n30208), .B(n30207), .Z(n30361) );
  XNOR U30992 ( .A(n30360), .B(n30361), .Z(n30304) );
  XNOR U30993 ( .A(n30305), .B(n30304), .Z(n30307) );
  NANDN U30994 ( .A(n30210), .B(n30209), .Z(n30214) );
  NANDN U30995 ( .A(n30212), .B(n30211), .Z(n30213) );
  AND U30996 ( .A(n30214), .B(n30213), .Z(n30306) );
  XOR U30997 ( .A(n30307), .B(n30306), .Z(n30421) );
  NANDN U30998 ( .A(n30216), .B(n30215), .Z(n30220) );
  NANDN U30999 ( .A(n30218), .B(n30217), .Z(n30219) );
  AND U31000 ( .A(n30220), .B(n30219), .Z(n30418) );
  NANDN U31001 ( .A(n30222), .B(n30221), .Z(n30226) );
  NANDN U31002 ( .A(n30224), .B(n30223), .Z(n30225) );
  AND U31003 ( .A(n30226), .B(n30225), .Z(n30301) );
  NANDN U31004 ( .A(n30228), .B(n30227), .Z(n30232) );
  OR U31005 ( .A(n30230), .B(n30229), .Z(n30231) );
  AND U31006 ( .A(n30232), .B(n30231), .Z(n30299) );
  NANDN U31007 ( .A(n30234), .B(n30233), .Z(n30238) );
  NANDN U31008 ( .A(n30236), .B(n30235), .Z(n30237) );
  AND U31009 ( .A(n30238), .B(n30237), .Z(n30365) );
  NANDN U31010 ( .A(n30240), .B(n30239), .Z(n30244) );
  NANDN U31011 ( .A(n30242), .B(n30241), .Z(n30243) );
  NAND U31012 ( .A(n30244), .B(n30243), .Z(n30364) );
  XNOR U31013 ( .A(n30365), .B(n30364), .Z(n30366) );
  NAND U31014 ( .A(b[0]), .B(a[218]), .Z(n30245) );
  XNOR U31015 ( .A(b[1]), .B(n30245), .Z(n30247) );
  NANDN U31016 ( .A(b[0]), .B(a[217]), .Z(n30246) );
  NAND U31017 ( .A(n30247), .B(n30246), .Z(n30313) );
  NAND U31018 ( .A(n194), .B(n30248), .Z(n30250) );
  XOR U31019 ( .A(b[29]), .B(a[190]), .Z(n30391) );
  NAND U31020 ( .A(n38456), .B(n30391), .Z(n30249) );
  AND U31021 ( .A(n30250), .B(n30249), .Z(n30311) );
  AND U31022 ( .A(b[31]), .B(a[186]), .Z(n30310) );
  XNOR U31023 ( .A(n30311), .B(n30310), .Z(n30312) );
  XNOR U31024 ( .A(n30313), .B(n30312), .Z(n30352) );
  NAND U31025 ( .A(n38185), .B(n30251), .Z(n30253) );
  XOR U31026 ( .A(b[23]), .B(a[196]), .Z(n30394) );
  NAND U31027 ( .A(n38132), .B(n30394), .Z(n30252) );
  AND U31028 ( .A(n30253), .B(n30252), .Z(n30385) );
  NAND U31029 ( .A(n184), .B(n30254), .Z(n30256) );
  XOR U31030 ( .A(b[7]), .B(a[212]), .Z(n30397) );
  NAND U31031 ( .A(n36592), .B(n30397), .Z(n30255) );
  AND U31032 ( .A(n30256), .B(n30255), .Z(n30383) );
  NAND U31033 ( .A(n38289), .B(n30257), .Z(n30259) );
  XOR U31034 ( .A(b[25]), .B(a[194]), .Z(n30400) );
  NAND U31035 ( .A(n38247), .B(n30400), .Z(n30258) );
  NAND U31036 ( .A(n30259), .B(n30258), .Z(n30382) );
  XNOR U31037 ( .A(n30383), .B(n30382), .Z(n30384) );
  XOR U31038 ( .A(n30385), .B(n30384), .Z(n30353) );
  XNOR U31039 ( .A(n30352), .B(n30353), .Z(n30354) );
  NAND U31040 ( .A(n187), .B(n30260), .Z(n30262) );
  XOR U31041 ( .A(b[13]), .B(a[206]), .Z(n30403) );
  NAND U31042 ( .A(n37295), .B(n30403), .Z(n30261) );
  AND U31043 ( .A(n30262), .B(n30261), .Z(n30347) );
  NAND U31044 ( .A(n186), .B(n30263), .Z(n30265) );
  XOR U31045 ( .A(b[11]), .B(a[208]), .Z(n30406) );
  NAND U31046 ( .A(n37097), .B(n30406), .Z(n30264) );
  NAND U31047 ( .A(n30265), .B(n30264), .Z(n30346) );
  XNOR U31048 ( .A(n30347), .B(n30346), .Z(n30348) );
  NAND U31049 ( .A(n188), .B(n30266), .Z(n30268) );
  XOR U31050 ( .A(b[15]), .B(a[204]), .Z(n30409) );
  NAND U31051 ( .A(n37382), .B(n30409), .Z(n30267) );
  AND U31052 ( .A(n30268), .B(n30267), .Z(n30343) );
  NAND U31053 ( .A(n38064), .B(n30269), .Z(n30271) );
  XOR U31054 ( .A(b[21]), .B(a[198]), .Z(n30412) );
  NAND U31055 ( .A(n37993), .B(n30412), .Z(n30270) );
  AND U31056 ( .A(n30271), .B(n30270), .Z(n30341) );
  NAND U31057 ( .A(n185), .B(n30272), .Z(n30274) );
  XOR U31058 ( .A(b[9]), .B(a[210]), .Z(n30415) );
  NAND U31059 ( .A(n36805), .B(n30415), .Z(n30273) );
  NAND U31060 ( .A(n30274), .B(n30273), .Z(n30340) );
  XNOR U31061 ( .A(n30341), .B(n30340), .Z(n30342) );
  XOR U31062 ( .A(n30343), .B(n30342), .Z(n30349) );
  XOR U31063 ( .A(n30348), .B(n30349), .Z(n30355) );
  XOR U31064 ( .A(n30354), .B(n30355), .Z(n30367) );
  XNOR U31065 ( .A(n30366), .B(n30367), .Z(n30298) );
  XNOR U31066 ( .A(n30299), .B(n30298), .Z(n30300) );
  XOR U31067 ( .A(n30301), .B(n30300), .Z(n30419) );
  XNOR U31068 ( .A(n30418), .B(n30419), .Z(n30420) );
  XNOR U31069 ( .A(n30421), .B(n30420), .Z(n30426) );
  XOR U31070 ( .A(n30427), .B(n30426), .Z(n30293) );
  NANDN U31071 ( .A(n30276), .B(n30275), .Z(n30280) );
  NANDN U31072 ( .A(n30278), .B(n30277), .Z(n30279) );
  AND U31073 ( .A(n30280), .B(n30279), .Z(n30292) );
  XOR U31074 ( .A(n30293), .B(n30292), .Z(n30295) );
  XNOR U31075 ( .A(n30294), .B(n30295), .Z(n30286) );
  XNOR U31076 ( .A(n30287), .B(n30286), .Z(n30288) );
  XNOR U31077 ( .A(n30289), .B(n30288), .Z(n30430) );
  XNOR U31078 ( .A(sreg[442]), .B(n30430), .Z(n30432) );
  NANDN U31079 ( .A(sreg[441]), .B(n30281), .Z(n30285) );
  NAND U31080 ( .A(n30283), .B(n30282), .Z(n30284) );
  NAND U31081 ( .A(n30285), .B(n30284), .Z(n30431) );
  XNOR U31082 ( .A(n30432), .B(n30431), .Z(c[442]) );
  NANDN U31083 ( .A(n30287), .B(n30286), .Z(n30291) );
  NANDN U31084 ( .A(n30289), .B(n30288), .Z(n30290) );
  AND U31085 ( .A(n30291), .B(n30290), .Z(n30438) );
  NANDN U31086 ( .A(n30293), .B(n30292), .Z(n30297) );
  NANDN U31087 ( .A(n30295), .B(n30294), .Z(n30296) );
  AND U31088 ( .A(n30297), .B(n30296), .Z(n30436) );
  NANDN U31089 ( .A(n30299), .B(n30298), .Z(n30303) );
  NANDN U31090 ( .A(n30301), .B(n30300), .Z(n30302) );
  AND U31091 ( .A(n30303), .B(n30302), .Z(n30448) );
  NANDN U31092 ( .A(n30305), .B(n30304), .Z(n30309) );
  NAND U31093 ( .A(n30307), .B(n30306), .Z(n30308) );
  AND U31094 ( .A(n30309), .B(n30308), .Z(n30447) );
  XNOR U31095 ( .A(n30448), .B(n30447), .Z(n30450) );
  NANDN U31096 ( .A(n30311), .B(n30310), .Z(n30315) );
  NANDN U31097 ( .A(n30313), .B(n30312), .Z(n30314) );
  AND U31098 ( .A(n30315), .B(n30314), .Z(n30527) );
  NAND U31099 ( .A(n38385), .B(n30316), .Z(n30318) );
  XOR U31100 ( .A(b[27]), .B(a[193]), .Z(n30471) );
  NAND U31101 ( .A(n38343), .B(n30471), .Z(n30317) );
  AND U31102 ( .A(n30318), .B(n30317), .Z(n30534) );
  NAND U31103 ( .A(n183), .B(n30319), .Z(n30321) );
  XOR U31104 ( .A(b[5]), .B(a[215]), .Z(n30474) );
  NAND U31105 ( .A(n36296), .B(n30474), .Z(n30320) );
  AND U31106 ( .A(n30321), .B(n30320), .Z(n30532) );
  NAND U31107 ( .A(n190), .B(n30322), .Z(n30324) );
  XOR U31108 ( .A(b[19]), .B(a[201]), .Z(n30477) );
  NAND U31109 ( .A(n37821), .B(n30477), .Z(n30323) );
  NAND U31110 ( .A(n30324), .B(n30323), .Z(n30531) );
  XNOR U31111 ( .A(n30532), .B(n30531), .Z(n30533) );
  XNOR U31112 ( .A(n30534), .B(n30533), .Z(n30525) );
  NAND U31113 ( .A(n38470), .B(n30325), .Z(n30327) );
  XOR U31114 ( .A(b[31]), .B(a[189]), .Z(n30480) );
  NAND U31115 ( .A(n38453), .B(n30480), .Z(n30326) );
  AND U31116 ( .A(n30327), .B(n30326), .Z(n30492) );
  NAND U31117 ( .A(n181), .B(n30328), .Z(n30330) );
  XOR U31118 ( .A(b[3]), .B(a[217]), .Z(n30483) );
  NAND U31119 ( .A(n182), .B(n30483), .Z(n30329) );
  AND U31120 ( .A(n30330), .B(n30329), .Z(n30490) );
  NAND U31121 ( .A(n189), .B(n30331), .Z(n30333) );
  XOR U31122 ( .A(b[17]), .B(a[203]), .Z(n30486) );
  NAND U31123 ( .A(n37652), .B(n30486), .Z(n30332) );
  NAND U31124 ( .A(n30333), .B(n30332), .Z(n30489) );
  XNOR U31125 ( .A(n30490), .B(n30489), .Z(n30491) );
  XOR U31126 ( .A(n30492), .B(n30491), .Z(n30526) );
  XOR U31127 ( .A(n30525), .B(n30526), .Z(n30528) );
  XOR U31128 ( .A(n30527), .B(n30528), .Z(n30460) );
  NANDN U31129 ( .A(n30335), .B(n30334), .Z(n30339) );
  NANDN U31130 ( .A(n30337), .B(n30336), .Z(n30338) );
  AND U31131 ( .A(n30339), .B(n30338), .Z(n30513) );
  NANDN U31132 ( .A(n30341), .B(n30340), .Z(n30345) );
  NANDN U31133 ( .A(n30343), .B(n30342), .Z(n30344) );
  NAND U31134 ( .A(n30345), .B(n30344), .Z(n30514) );
  XNOR U31135 ( .A(n30513), .B(n30514), .Z(n30515) );
  NANDN U31136 ( .A(n30347), .B(n30346), .Z(n30351) );
  NANDN U31137 ( .A(n30349), .B(n30348), .Z(n30350) );
  NAND U31138 ( .A(n30351), .B(n30350), .Z(n30516) );
  XNOR U31139 ( .A(n30515), .B(n30516), .Z(n30459) );
  XNOR U31140 ( .A(n30460), .B(n30459), .Z(n30462) );
  NANDN U31141 ( .A(n30353), .B(n30352), .Z(n30357) );
  NANDN U31142 ( .A(n30355), .B(n30354), .Z(n30356) );
  AND U31143 ( .A(n30357), .B(n30356), .Z(n30461) );
  XOR U31144 ( .A(n30462), .B(n30461), .Z(n30576) );
  NANDN U31145 ( .A(n30359), .B(n30358), .Z(n30363) );
  NANDN U31146 ( .A(n30361), .B(n30360), .Z(n30362) );
  AND U31147 ( .A(n30363), .B(n30362), .Z(n30573) );
  NANDN U31148 ( .A(n30365), .B(n30364), .Z(n30369) );
  NANDN U31149 ( .A(n30367), .B(n30366), .Z(n30368) );
  AND U31150 ( .A(n30369), .B(n30368), .Z(n30456) );
  NANDN U31151 ( .A(n30371), .B(n30370), .Z(n30375) );
  OR U31152 ( .A(n30373), .B(n30372), .Z(n30374) );
  AND U31153 ( .A(n30375), .B(n30374), .Z(n30454) );
  NANDN U31154 ( .A(n30377), .B(n30376), .Z(n30381) );
  NANDN U31155 ( .A(n30379), .B(n30378), .Z(n30380) );
  AND U31156 ( .A(n30381), .B(n30380), .Z(n30520) );
  NANDN U31157 ( .A(n30383), .B(n30382), .Z(n30387) );
  NANDN U31158 ( .A(n30385), .B(n30384), .Z(n30386) );
  NAND U31159 ( .A(n30387), .B(n30386), .Z(n30519) );
  XNOR U31160 ( .A(n30520), .B(n30519), .Z(n30521) );
  NAND U31161 ( .A(b[0]), .B(a[219]), .Z(n30388) );
  XNOR U31162 ( .A(b[1]), .B(n30388), .Z(n30390) );
  NANDN U31163 ( .A(b[0]), .B(a[218]), .Z(n30389) );
  NAND U31164 ( .A(n30390), .B(n30389), .Z(n30468) );
  NAND U31165 ( .A(n194), .B(n30391), .Z(n30393) );
  XOR U31166 ( .A(b[29]), .B(a[191]), .Z(n30546) );
  NAND U31167 ( .A(n38456), .B(n30546), .Z(n30392) );
  AND U31168 ( .A(n30393), .B(n30392), .Z(n30466) );
  AND U31169 ( .A(b[31]), .B(a[187]), .Z(n30465) );
  XNOR U31170 ( .A(n30466), .B(n30465), .Z(n30467) );
  XNOR U31171 ( .A(n30468), .B(n30467), .Z(n30507) );
  NAND U31172 ( .A(n38185), .B(n30394), .Z(n30396) );
  XOR U31173 ( .A(b[23]), .B(a[197]), .Z(n30549) );
  NAND U31174 ( .A(n38132), .B(n30549), .Z(n30395) );
  AND U31175 ( .A(n30396), .B(n30395), .Z(n30540) );
  NAND U31176 ( .A(n184), .B(n30397), .Z(n30399) );
  XOR U31177 ( .A(b[7]), .B(a[213]), .Z(n30552) );
  NAND U31178 ( .A(n36592), .B(n30552), .Z(n30398) );
  AND U31179 ( .A(n30399), .B(n30398), .Z(n30538) );
  NAND U31180 ( .A(n38289), .B(n30400), .Z(n30402) );
  XOR U31181 ( .A(b[25]), .B(a[195]), .Z(n30555) );
  NAND U31182 ( .A(n38247), .B(n30555), .Z(n30401) );
  NAND U31183 ( .A(n30402), .B(n30401), .Z(n30537) );
  XNOR U31184 ( .A(n30538), .B(n30537), .Z(n30539) );
  XOR U31185 ( .A(n30540), .B(n30539), .Z(n30508) );
  XNOR U31186 ( .A(n30507), .B(n30508), .Z(n30509) );
  NAND U31187 ( .A(n187), .B(n30403), .Z(n30405) );
  XOR U31188 ( .A(b[13]), .B(a[207]), .Z(n30558) );
  NAND U31189 ( .A(n37295), .B(n30558), .Z(n30404) );
  AND U31190 ( .A(n30405), .B(n30404), .Z(n30502) );
  NAND U31191 ( .A(n186), .B(n30406), .Z(n30408) );
  XOR U31192 ( .A(b[11]), .B(a[209]), .Z(n30561) );
  NAND U31193 ( .A(n37097), .B(n30561), .Z(n30407) );
  NAND U31194 ( .A(n30408), .B(n30407), .Z(n30501) );
  XNOR U31195 ( .A(n30502), .B(n30501), .Z(n30503) );
  NAND U31196 ( .A(n188), .B(n30409), .Z(n30411) );
  XOR U31197 ( .A(b[15]), .B(a[205]), .Z(n30564) );
  NAND U31198 ( .A(n37382), .B(n30564), .Z(n30410) );
  AND U31199 ( .A(n30411), .B(n30410), .Z(n30498) );
  NAND U31200 ( .A(n38064), .B(n30412), .Z(n30414) );
  XOR U31201 ( .A(b[21]), .B(a[199]), .Z(n30567) );
  NAND U31202 ( .A(n37993), .B(n30567), .Z(n30413) );
  AND U31203 ( .A(n30414), .B(n30413), .Z(n30496) );
  NAND U31204 ( .A(n185), .B(n30415), .Z(n30417) );
  XOR U31205 ( .A(b[9]), .B(a[211]), .Z(n30570) );
  NAND U31206 ( .A(n36805), .B(n30570), .Z(n30416) );
  NAND U31207 ( .A(n30417), .B(n30416), .Z(n30495) );
  XNOR U31208 ( .A(n30496), .B(n30495), .Z(n30497) );
  XOR U31209 ( .A(n30498), .B(n30497), .Z(n30504) );
  XOR U31210 ( .A(n30503), .B(n30504), .Z(n30510) );
  XOR U31211 ( .A(n30509), .B(n30510), .Z(n30522) );
  XNOR U31212 ( .A(n30521), .B(n30522), .Z(n30453) );
  XNOR U31213 ( .A(n30454), .B(n30453), .Z(n30455) );
  XOR U31214 ( .A(n30456), .B(n30455), .Z(n30574) );
  XNOR U31215 ( .A(n30573), .B(n30574), .Z(n30575) );
  XNOR U31216 ( .A(n30576), .B(n30575), .Z(n30449) );
  XOR U31217 ( .A(n30450), .B(n30449), .Z(n30442) );
  NANDN U31218 ( .A(n30419), .B(n30418), .Z(n30423) );
  NANDN U31219 ( .A(n30421), .B(n30420), .Z(n30422) );
  AND U31220 ( .A(n30423), .B(n30422), .Z(n30441) );
  XNOR U31221 ( .A(n30442), .B(n30441), .Z(n30443) );
  NANDN U31222 ( .A(n30425), .B(n30424), .Z(n30429) );
  NAND U31223 ( .A(n30427), .B(n30426), .Z(n30428) );
  NAND U31224 ( .A(n30429), .B(n30428), .Z(n30444) );
  XNOR U31225 ( .A(n30443), .B(n30444), .Z(n30435) );
  XNOR U31226 ( .A(n30436), .B(n30435), .Z(n30437) );
  XNOR U31227 ( .A(n30438), .B(n30437), .Z(n30579) );
  XNOR U31228 ( .A(sreg[443]), .B(n30579), .Z(n30581) );
  NANDN U31229 ( .A(sreg[442]), .B(n30430), .Z(n30434) );
  NAND U31230 ( .A(n30432), .B(n30431), .Z(n30433) );
  NAND U31231 ( .A(n30434), .B(n30433), .Z(n30580) );
  XNOR U31232 ( .A(n30581), .B(n30580), .Z(c[443]) );
  NANDN U31233 ( .A(n30436), .B(n30435), .Z(n30440) );
  NANDN U31234 ( .A(n30438), .B(n30437), .Z(n30439) );
  AND U31235 ( .A(n30440), .B(n30439), .Z(n30587) );
  NANDN U31236 ( .A(n30442), .B(n30441), .Z(n30446) );
  NANDN U31237 ( .A(n30444), .B(n30443), .Z(n30445) );
  AND U31238 ( .A(n30446), .B(n30445), .Z(n30585) );
  NANDN U31239 ( .A(n30448), .B(n30447), .Z(n30452) );
  NAND U31240 ( .A(n30450), .B(n30449), .Z(n30451) );
  AND U31241 ( .A(n30452), .B(n30451), .Z(n30592) );
  NANDN U31242 ( .A(n30454), .B(n30453), .Z(n30458) );
  NANDN U31243 ( .A(n30456), .B(n30455), .Z(n30457) );
  AND U31244 ( .A(n30458), .B(n30457), .Z(n30597) );
  NANDN U31245 ( .A(n30460), .B(n30459), .Z(n30464) );
  NAND U31246 ( .A(n30462), .B(n30461), .Z(n30463) );
  AND U31247 ( .A(n30464), .B(n30463), .Z(n30596) );
  XNOR U31248 ( .A(n30597), .B(n30596), .Z(n30599) );
  NANDN U31249 ( .A(n30466), .B(n30465), .Z(n30470) );
  NANDN U31250 ( .A(n30468), .B(n30467), .Z(n30469) );
  AND U31251 ( .A(n30470), .B(n30469), .Z(n30674) );
  NAND U31252 ( .A(n38385), .B(n30471), .Z(n30473) );
  XOR U31253 ( .A(b[27]), .B(a[194]), .Z(n30620) );
  NAND U31254 ( .A(n38343), .B(n30620), .Z(n30472) );
  AND U31255 ( .A(n30473), .B(n30472), .Z(n30681) );
  NAND U31256 ( .A(n183), .B(n30474), .Z(n30476) );
  XOR U31257 ( .A(b[5]), .B(a[216]), .Z(n30623) );
  NAND U31258 ( .A(n36296), .B(n30623), .Z(n30475) );
  AND U31259 ( .A(n30476), .B(n30475), .Z(n30679) );
  NAND U31260 ( .A(n190), .B(n30477), .Z(n30479) );
  XOR U31261 ( .A(b[19]), .B(a[202]), .Z(n30626) );
  NAND U31262 ( .A(n37821), .B(n30626), .Z(n30478) );
  NAND U31263 ( .A(n30479), .B(n30478), .Z(n30678) );
  XNOR U31264 ( .A(n30679), .B(n30678), .Z(n30680) );
  XNOR U31265 ( .A(n30681), .B(n30680), .Z(n30672) );
  NAND U31266 ( .A(n38470), .B(n30480), .Z(n30482) );
  XOR U31267 ( .A(b[31]), .B(a[190]), .Z(n30629) );
  NAND U31268 ( .A(n38453), .B(n30629), .Z(n30481) );
  AND U31269 ( .A(n30482), .B(n30481), .Z(n30641) );
  NAND U31270 ( .A(n181), .B(n30483), .Z(n30485) );
  XOR U31271 ( .A(b[3]), .B(a[218]), .Z(n30632) );
  NAND U31272 ( .A(n182), .B(n30632), .Z(n30484) );
  AND U31273 ( .A(n30485), .B(n30484), .Z(n30639) );
  NAND U31274 ( .A(n189), .B(n30486), .Z(n30488) );
  XOR U31275 ( .A(b[17]), .B(a[204]), .Z(n30635) );
  NAND U31276 ( .A(n37652), .B(n30635), .Z(n30487) );
  NAND U31277 ( .A(n30488), .B(n30487), .Z(n30638) );
  XNOR U31278 ( .A(n30639), .B(n30638), .Z(n30640) );
  XOR U31279 ( .A(n30641), .B(n30640), .Z(n30673) );
  XOR U31280 ( .A(n30672), .B(n30673), .Z(n30675) );
  XOR U31281 ( .A(n30674), .B(n30675), .Z(n30609) );
  NANDN U31282 ( .A(n30490), .B(n30489), .Z(n30494) );
  NANDN U31283 ( .A(n30492), .B(n30491), .Z(n30493) );
  AND U31284 ( .A(n30494), .B(n30493), .Z(n30662) );
  NANDN U31285 ( .A(n30496), .B(n30495), .Z(n30500) );
  NANDN U31286 ( .A(n30498), .B(n30497), .Z(n30499) );
  NAND U31287 ( .A(n30500), .B(n30499), .Z(n30663) );
  XNOR U31288 ( .A(n30662), .B(n30663), .Z(n30664) );
  NANDN U31289 ( .A(n30502), .B(n30501), .Z(n30506) );
  NANDN U31290 ( .A(n30504), .B(n30503), .Z(n30505) );
  NAND U31291 ( .A(n30506), .B(n30505), .Z(n30665) );
  XNOR U31292 ( .A(n30664), .B(n30665), .Z(n30608) );
  XNOR U31293 ( .A(n30609), .B(n30608), .Z(n30611) );
  NANDN U31294 ( .A(n30508), .B(n30507), .Z(n30512) );
  NANDN U31295 ( .A(n30510), .B(n30509), .Z(n30511) );
  AND U31296 ( .A(n30512), .B(n30511), .Z(n30610) );
  XOR U31297 ( .A(n30611), .B(n30610), .Z(n30723) );
  NANDN U31298 ( .A(n30514), .B(n30513), .Z(n30518) );
  NANDN U31299 ( .A(n30516), .B(n30515), .Z(n30517) );
  AND U31300 ( .A(n30518), .B(n30517), .Z(n30720) );
  NANDN U31301 ( .A(n30520), .B(n30519), .Z(n30524) );
  NANDN U31302 ( .A(n30522), .B(n30521), .Z(n30523) );
  AND U31303 ( .A(n30524), .B(n30523), .Z(n30605) );
  NANDN U31304 ( .A(n30526), .B(n30525), .Z(n30530) );
  OR U31305 ( .A(n30528), .B(n30527), .Z(n30529) );
  AND U31306 ( .A(n30530), .B(n30529), .Z(n30603) );
  NANDN U31307 ( .A(n30532), .B(n30531), .Z(n30536) );
  NANDN U31308 ( .A(n30534), .B(n30533), .Z(n30535) );
  AND U31309 ( .A(n30536), .B(n30535), .Z(n30669) );
  NANDN U31310 ( .A(n30538), .B(n30537), .Z(n30542) );
  NANDN U31311 ( .A(n30540), .B(n30539), .Z(n30541) );
  NAND U31312 ( .A(n30542), .B(n30541), .Z(n30668) );
  XNOR U31313 ( .A(n30669), .B(n30668), .Z(n30671) );
  NAND U31314 ( .A(b[0]), .B(a[220]), .Z(n30543) );
  XNOR U31315 ( .A(b[1]), .B(n30543), .Z(n30545) );
  NANDN U31316 ( .A(b[0]), .B(a[219]), .Z(n30544) );
  NAND U31317 ( .A(n30545), .B(n30544), .Z(n30617) );
  NAND U31318 ( .A(n194), .B(n30546), .Z(n30548) );
  XOR U31319 ( .A(b[29]), .B(a[192]), .Z(n30693) );
  NAND U31320 ( .A(n38456), .B(n30693), .Z(n30547) );
  AND U31321 ( .A(n30548), .B(n30547), .Z(n30615) );
  AND U31322 ( .A(b[31]), .B(a[188]), .Z(n30614) );
  XNOR U31323 ( .A(n30615), .B(n30614), .Z(n30616) );
  XNOR U31324 ( .A(n30617), .B(n30616), .Z(n30657) );
  NAND U31325 ( .A(n38185), .B(n30549), .Z(n30551) );
  XOR U31326 ( .A(b[23]), .B(a[198]), .Z(n30696) );
  NAND U31327 ( .A(n38132), .B(n30696), .Z(n30550) );
  AND U31328 ( .A(n30551), .B(n30550), .Z(n30686) );
  NAND U31329 ( .A(n184), .B(n30552), .Z(n30554) );
  XOR U31330 ( .A(b[7]), .B(a[214]), .Z(n30699) );
  NAND U31331 ( .A(n36592), .B(n30699), .Z(n30553) );
  AND U31332 ( .A(n30554), .B(n30553), .Z(n30685) );
  NAND U31333 ( .A(n38289), .B(n30555), .Z(n30557) );
  XOR U31334 ( .A(b[25]), .B(a[196]), .Z(n30702) );
  NAND U31335 ( .A(n38247), .B(n30702), .Z(n30556) );
  NAND U31336 ( .A(n30557), .B(n30556), .Z(n30684) );
  XOR U31337 ( .A(n30685), .B(n30684), .Z(n30687) );
  XOR U31338 ( .A(n30686), .B(n30687), .Z(n30656) );
  XOR U31339 ( .A(n30657), .B(n30656), .Z(n30659) );
  NAND U31340 ( .A(n187), .B(n30558), .Z(n30560) );
  XOR U31341 ( .A(b[13]), .B(a[208]), .Z(n30705) );
  NAND U31342 ( .A(n37295), .B(n30705), .Z(n30559) );
  AND U31343 ( .A(n30560), .B(n30559), .Z(n30651) );
  NAND U31344 ( .A(n186), .B(n30561), .Z(n30563) );
  XOR U31345 ( .A(b[11]), .B(a[210]), .Z(n30708) );
  NAND U31346 ( .A(n37097), .B(n30708), .Z(n30562) );
  NAND U31347 ( .A(n30563), .B(n30562), .Z(n30650) );
  XNOR U31348 ( .A(n30651), .B(n30650), .Z(n30653) );
  NAND U31349 ( .A(n188), .B(n30564), .Z(n30566) );
  XOR U31350 ( .A(b[15]), .B(a[206]), .Z(n30711) );
  NAND U31351 ( .A(n37382), .B(n30711), .Z(n30565) );
  AND U31352 ( .A(n30566), .B(n30565), .Z(n30647) );
  NAND U31353 ( .A(n38064), .B(n30567), .Z(n30569) );
  XOR U31354 ( .A(b[21]), .B(a[200]), .Z(n30714) );
  NAND U31355 ( .A(n37993), .B(n30714), .Z(n30568) );
  AND U31356 ( .A(n30569), .B(n30568), .Z(n30645) );
  NAND U31357 ( .A(n185), .B(n30570), .Z(n30572) );
  XOR U31358 ( .A(b[9]), .B(a[212]), .Z(n30717) );
  NAND U31359 ( .A(n36805), .B(n30717), .Z(n30571) );
  NAND U31360 ( .A(n30572), .B(n30571), .Z(n30644) );
  XNOR U31361 ( .A(n30645), .B(n30644), .Z(n30646) );
  XNOR U31362 ( .A(n30647), .B(n30646), .Z(n30652) );
  XOR U31363 ( .A(n30653), .B(n30652), .Z(n30658) );
  XNOR U31364 ( .A(n30659), .B(n30658), .Z(n30670) );
  XNOR U31365 ( .A(n30671), .B(n30670), .Z(n30602) );
  XNOR U31366 ( .A(n30603), .B(n30602), .Z(n30604) );
  XOR U31367 ( .A(n30605), .B(n30604), .Z(n30721) );
  XNOR U31368 ( .A(n30720), .B(n30721), .Z(n30722) );
  XNOR U31369 ( .A(n30723), .B(n30722), .Z(n30598) );
  XOR U31370 ( .A(n30599), .B(n30598), .Z(n30591) );
  NANDN U31371 ( .A(n30574), .B(n30573), .Z(n30578) );
  NANDN U31372 ( .A(n30576), .B(n30575), .Z(n30577) );
  AND U31373 ( .A(n30578), .B(n30577), .Z(n30590) );
  XOR U31374 ( .A(n30591), .B(n30590), .Z(n30593) );
  XNOR U31375 ( .A(n30592), .B(n30593), .Z(n30584) );
  XNOR U31376 ( .A(n30585), .B(n30584), .Z(n30586) );
  XNOR U31377 ( .A(n30587), .B(n30586), .Z(n30726) );
  XNOR U31378 ( .A(sreg[444]), .B(n30726), .Z(n30728) );
  NANDN U31379 ( .A(sreg[443]), .B(n30579), .Z(n30583) );
  NAND U31380 ( .A(n30581), .B(n30580), .Z(n30582) );
  NAND U31381 ( .A(n30583), .B(n30582), .Z(n30727) );
  XNOR U31382 ( .A(n30728), .B(n30727), .Z(c[444]) );
  NANDN U31383 ( .A(n30585), .B(n30584), .Z(n30589) );
  NANDN U31384 ( .A(n30587), .B(n30586), .Z(n30588) );
  AND U31385 ( .A(n30589), .B(n30588), .Z(n30734) );
  NANDN U31386 ( .A(n30591), .B(n30590), .Z(n30595) );
  NANDN U31387 ( .A(n30593), .B(n30592), .Z(n30594) );
  AND U31388 ( .A(n30595), .B(n30594), .Z(n30732) );
  NANDN U31389 ( .A(n30597), .B(n30596), .Z(n30601) );
  NAND U31390 ( .A(n30599), .B(n30598), .Z(n30600) );
  AND U31391 ( .A(n30601), .B(n30600), .Z(n30739) );
  NANDN U31392 ( .A(n30603), .B(n30602), .Z(n30607) );
  NANDN U31393 ( .A(n30605), .B(n30604), .Z(n30606) );
  AND U31394 ( .A(n30607), .B(n30606), .Z(n30744) );
  NANDN U31395 ( .A(n30609), .B(n30608), .Z(n30613) );
  NAND U31396 ( .A(n30611), .B(n30610), .Z(n30612) );
  AND U31397 ( .A(n30613), .B(n30612), .Z(n30743) );
  XNOR U31398 ( .A(n30744), .B(n30743), .Z(n30746) );
  NANDN U31399 ( .A(n30615), .B(n30614), .Z(n30619) );
  NANDN U31400 ( .A(n30617), .B(n30616), .Z(n30618) );
  AND U31401 ( .A(n30619), .B(n30618), .Z(n30809) );
  NAND U31402 ( .A(n38385), .B(n30620), .Z(n30622) );
  XOR U31403 ( .A(b[27]), .B(a[195]), .Z(n30755) );
  NAND U31404 ( .A(n38343), .B(n30755), .Z(n30621) );
  AND U31405 ( .A(n30622), .B(n30621), .Z(n30816) );
  NAND U31406 ( .A(n183), .B(n30623), .Z(n30625) );
  XOR U31407 ( .A(b[5]), .B(a[217]), .Z(n30758) );
  NAND U31408 ( .A(n36296), .B(n30758), .Z(n30624) );
  AND U31409 ( .A(n30625), .B(n30624), .Z(n30814) );
  NAND U31410 ( .A(n190), .B(n30626), .Z(n30628) );
  XOR U31411 ( .A(b[19]), .B(a[203]), .Z(n30761) );
  NAND U31412 ( .A(n37821), .B(n30761), .Z(n30627) );
  NAND U31413 ( .A(n30628), .B(n30627), .Z(n30813) );
  XNOR U31414 ( .A(n30814), .B(n30813), .Z(n30815) );
  XNOR U31415 ( .A(n30816), .B(n30815), .Z(n30807) );
  NAND U31416 ( .A(n38470), .B(n30629), .Z(n30631) );
  XOR U31417 ( .A(b[31]), .B(a[191]), .Z(n30764) );
  NAND U31418 ( .A(n38453), .B(n30764), .Z(n30630) );
  AND U31419 ( .A(n30631), .B(n30630), .Z(n30776) );
  NAND U31420 ( .A(n181), .B(n30632), .Z(n30634) );
  XOR U31421 ( .A(b[3]), .B(a[219]), .Z(n30767) );
  NAND U31422 ( .A(n182), .B(n30767), .Z(n30633) );
  AND U31423 ( .A(n30634), .B(n30633), .Z(n30774) );
  NAND U31424 ( .A(n189), .B(n30635), .Z(n30637) );
  XOR U31425 ( .A(b[17]), .B(a[205]), .Z(n30770) );
  NAND U31426 ( .A(n37652), .B(n30770), .Z(n30636) );
  NAND U31427 ( .A(n30637), .B(n30636), .Z(n30773) );
  XNOR U31428 ( .A(n30774), .B(n30773), .Z(n30775) );
  XOR U31429 ( .A(n30776), .B(n30775), .Z(n30808) );
  XOR U31430 ( .A(n30807), .B(n30808), .Z(n30810) );
  XOR U31431 ( .A(n30809), .B(n30810), .Z(n30856) );
  NANDN U31432 ( .A(n30639), .B(n30638), .Z(n30643) );
  NANDN U31433 ( .A(n30641), .B(n30640), .Z(n30642) );
  AND U31434 ( .A(n30643), .B(n30642), .Z(n30797) );
  NANDN U31435 ( .A(n30645), .B(n30644), .Z(n30649) );
  NANDN U31436 ( .A(n30647), .B(n30646), .Z(n30648) );
  NAND U31437 ( .A(n30649), .B(n30648), .Z(n30798) );
  XNOR U31438 ( .A(n30797), .B(n30798), .Z(n30799) );
  NANDN U31439 ( .A(n30651), .B(n30650), .Z(n30655) );
  NAND U31440 ( .A(n30653), .B(n30652), .Z(n30654) );
  NAND U31441 ( .A(n30655), .B(n30654), .Z(n30800) );
  XNOR U31442 ( .A(n30799), .B(n30800), .Z(n30855) );
  XNOR U31443 ( .A(n30856), .B(n30855), .Z(n30858) );
  NAND U31444 ( .A(n30657), .B(n30656), .Z(n30661) );
  NAND U31445 ( .A(n30659), .B(n30658), .Z(n30660) );
  AND U31446 ( .A(n30661), .B(n30660), .Z(n30857) );
  XOR U31447 ( .A(n30858), .B(n30857), .Z(n30870) );
  NANDN U31448 ( .A(n30663), .B(n30662), .Z(n30667) );
  NANDN U31449 ( .A(n30665), .B(n30664), .Z(n30666) );
  AND U31450 ( .A(n30667), .B(n30666), .Z(n30867) );
  NANDN U31451 ( .A(n30673), .B(n30672), .Z(n30677) );
  OR U31452 ( .A(n30675), .B(n30674), .Z(n30676) );
  AND U31453 ( .A(n30677), .B(n30676), .Z(n30862) );
  NANDN U31454 ( .A(n30679), .B(n30678), .Z(n30683) );
  NANDN U31455 ( .A(n30681), .B(n30680), .Z(n30682) );
  AND U31456 ( .A(n30683), .B(n30682), .Z(n30804) );
  NANDN U31457 ( .A(n30685), .B(n30684), .Z(n30689) );
  OR U31458 ( .A(n30687), .B(n30686), .Z(n30688) );
  NAND U31459 ( .A(n30689), .B(n30688), .Z(n30803) );
  XNOR U31460 ( .A(n30804), .B(n30803), .Z(n30806) );
  NAND U31461 ( .A(b[0]), .B(a[221]), .Z(n30690) );
  XNOR U31462 ( .A(b[1]), .B(n30690), .Z(n30692) );
  NANDN U31463 ( .A(b[0]), .B(a[220]), .Z(n30691) );
  NAND U31464 ( .A(n30692), .B(n30691), .Z(n30752) );
  NAND U31465 ( .A(n194), .B(n30693), .Z(n30695) );
  XOR U31466 ( .A(b[29]), .B(a[193]), .Z(n30825) );
  NAND U31467 ( .A(n38456), .B(n30825), .Z(n30694) );
  AND U31468 ( .A(n30695), .B(n30694), .Z(n30750) );
  AND U31469 ( .A(b[31]), .B(a[189]), .Z(n30749) );
  XNOR U31470 ( .A(n30750), .B(n30749), .Z(n30751) );
  XNOR U31471 ( .A(n30752), .B(n30751), .Z(n30792) );
  NAND U31472 ( .A(n38185), .B(n30696), .Z(n30698) );
  XOR U31473 ( .A(b[23]), .B(a[199]), .Z(n30831) );
  NAND U31474 ( .A(n38132), .B(n30831), .Z(n30697) );
  AND U31475 ( .A(n30698), .B(n30697), .Z(n30821) );
  NAND U31476 ( .A(n184), .B(n30699), .Z(n30701) );
  XOR U31477 ( .A(b[7]), .B(a[215]), .Z(n30834) );
  NAND U31478 ( .A(n36592), .B(n30834), .Z(n30700) );
  AND U31479 ( .A(n30701), .B(n30700), .Z(n30820) );
  NAND U31480 ( .A(n38289), .B(n30702), .Z(n30704) );
  XOR U31481 ( .A(b[25]), .B(a[197]), .Z(n30837) );
  NAND U31482 ( .A(n38247), .B(n30837), .Z(n30703) );
  NAND U31483 ( .A(n30704), .B(n30703), .Z(n30819) );
  XOR U31484 ( .A(n30820), .B(n30819), .Z(n30822) );
  XOR U31485 ( .A(n30821), .B(n30822), .Z(n30791) );
  XOR U31486 ( .A(n30792), .B(n30791), .Z(n30794) );
  NAND U31487 ( .A(n187), .B(n30705), .Z(n30707) );
  XOR U31488 ( .A(b[13]), .B(a[209]), .Z(n30840) );
  NAND U31489 ( .A(n37295), .B(n30840), .Z(n30706) );
  AND U31490 ( .A(n30707), .B(n30706), .Z(n30786) );
  NAND U31491 ( .A(n186), .B(n30708), .Z(n30710) );
  XOR U31492 ( .A(b[11]), .B(a[211]), .Z(n30843) );
  NAND U31493 ( .A(n37097), .B(n30843), .Z(n30709) );
  NAND U31494 ( .A(n30710), .B(n30709), .Z(n30785) );
  XNOR U31495 ( .A(n30786), .B(n30785), .Z(n30788) );
  NAND U31496 ( .A(n188), .B(n30711), .Z(n30713) );
  XOR U31497 ( .A(b[15]), .B(a[207]), .Z(n30846) );
  NAND U31498 ( .A(n37382), .B(n30846), .Z(n30712) );
  AND U31499 ( .A(n30713), .B(n30712), .Z(n30782) );
  NAND U31500 ( .A(n38064), .B(n30714), .Z(n30716) );
  XOR U31501 ( .A(b[21]), .B(a[201]), .Z(n30849) );
  NAND U31502 ( .A(n37993), .B(n30849), .Z(n30715) );
  AND U31503 ( .A(n30716), .B(n30715), .Z(n30780) );
  NAND U31504 ( .A(n185), .B(n30717), .Z(n30719) );
  XOR U31505 ( .A(b[9]), .B(a[213]), .Z(n30852) );
  NAND U31506 ( .A(n36805), .B(n30852), .Z(n30718) );
  NAND U31507 ( .A(n30719), .B(n30718), .Z(n30779) );
  XNOR U31508 ( .A(n30780), .B(n30779), .Z(n30781) );
  XNOR U31509 ( .A(n30782), .B(n30781), .Z(n30787) );
  XOR U31510 ( .A(n30788), .B(n30787), .Z(n30793) );
  XNOR U31511 ( .A(n30794), .B(n30793), .Z(n30805) );
  XNOR U31512 ( .A(n30806), .B(n30805), .Z(n30861) );
  XNOR U31513 ( .A(n30862), .B(n30861), .Z(n30863) );
  XOR U31514 ( .A(n30864), .B(n30863), .Z(n30868) );
  XNOR U31515 ( .A(n30867), .B(n30868), .Z(n30869) );
  XNOR U31516 ( .A(n30870), .B(n30869), .Z(n30745) );
  XOR U31517 ( .A(n30746), .B(n30745), .Z(n30738) );
  NANDN U31518 ( .A(n30721), .B(n30720), .Z(n30725) );
  NANDN U31519 ( .A(n30723), .B(n30722), .Z(n30724) );
  AND U31520 ( .A(n30725), .B(n30724), .Z(n30737) );
  XOR U31521 ( .A(n30738), .B(n30737), .Z(n30740) );
  XNOR U31522 ( .A(n30739), .B(n30740), .Z(n30731) );
  XNOR U31523 ( .A(n30732), .B(n30731), .Z(n30733) );
  XNOR U31524 ( .A(n30734), .B(n30733), .Z(n30873) );
  XNOR U31525 ( .A(sreg[445]), .B(n30873), .Z(n30875) );
  NANDN U31526 ( .A(sreg[444]), .B(n30726), .Z(n30730) );
  NAND U31527 ( .A(n30728), .B(n30727), .Z(n30729) );
  NAND U31528 ( .A(n30730), .B(n30729), .Z(n30874) );
  XNOR U31529 ( .A(n30875), .B(n30874), .Z(c[445]) );
  NANDN U31530 ( .A(n30732), .B(n30731), .Z(n30736) );
  NANDN U31531 ( .A(n30734), .B(n30733), .Z(n30735) );
  AND U31532 ( .A(n30736), .B(n30735), .Z(n30881) );
  NANDN U31533 ( .A(n30738), .B(n30737), .Z(n30742) );
  NANDN U31534 ( .A(n30740), .B(n30739), .Z(n30741) );
  AND U31535 ( .A(n30742), .B(n30741), .Z(n30879) );
  NANDN U31536 ( .A(n30744), .B(n30743), .Z(n30748) );
  NAND U31537 ( .A(n30746), .B(n30745), .Z(n30747) );
  AND U31538 ( .A(n30748), .B(n30747), .Z(n30886) );
  NANDN U31539 ( .A(n30750), .B(n30749), .Z(n30754) );
  NANDN U31540 ( .A(n30752), .B(n30751), .Z(n30753) );
  AND U31541 ( .A(n30754), .B(n30753), .Z(n30956) );
  NAND U31542 ( .A(n38385), .B(n30755), .Z(n30757) );
  XOR U31543 ( .A(b[27]), .B(a[196]), .Z(n30902) );
  NAND U31544 ( .A(n38343), .B(n30902), .Z(n30756) );
  AND U31545 ( .A(n30757), .B(n30756), .Z(n30963) );
  NAND U31546 ( .A(n183), .B(n30758), .Z(n30760) );
  XOR U31547 ( .A(b[5]), .B(a[218]), .Z(n30905) );
  NAND U31548 ( .A(n36296), .B(n30905), .Z(n30759) );
  AND U31549 ( .A(n30760), .B(n30759), .Z(n30961) );
  NAND U31550 ( .A(n190), .B(n30761), .Z(n30763) );
  XOR U31551 ( .A(b[19]), .B(a[204]), .Z(n30908) );
  NAND U31552 ( .A(n37821), .B(n30908), .Z(n30762) );
  NAND U31553 ( .A(n30763), .B(n30762), .Z(n30960) );
  XNOR U31554 ( .A(n30961), .B(n30960), .Z(n30962) );
  XNOR U31555 ( .A(n30963), .B(n30962), .Z(n30954) );
  NAND U31556 ( .A(n38470), .B(n30764), .Z(n30766) );
  XOR U31557 ( .A(b[31]), .B(a[192]), .Z(n30911) );
  NAND U31558 ( .A(n38453), .B(n30911), .Z(n30765) );
  AND U31559 ( .A(n30766), .B(n30765), .Z(n30923) );
  NAND U31560 ( .A(n181), .B(n30767), .Z(n30769) );
  XOR U31561 ( .A(b[3]), .B(a[220]), .Z(n30914) );
  NAND U31562 ( .A(n182), .B(n30914), .Z(n30768) );
  AND U31563 ( .A(n30769), .B(n30768), .Z(n30921) );
  NAND U31564 ( .A(n189), .B(n30770), .Z(n30772) );
  XOR U31565 ( .A(b[17]), .B(a[206]), .Z(n30917) );
  NAND U31566 ( .A(n37652), .B(n30917), .Z(n30771) );
  NAND U31567 ( .A(n30772), .B(n30771), .Z(n30920) );
  XNOR U31568 ( .A(n30921), .B(n30920), .Z(n30922) );
  XOR U31569 ( .A(n30923), .B(n30922), .Z(n30955) );
  XOR U31570 ( .A(n30954), .B(n30955), .Z(n30957) );
  XOR U31571 ( .A(n30956), .B(n30957), .Z(n31003) );
  NANDN U31572 ( .A(n30774), .B(n30773), .Z(n30778) );
  NANDN U31573 ( .A(n30776), .B(n30775), .Z(n30777) );
  AND U31574 ( .A(n30778), .B(n30777), .Z(n30944) );
  NANDN U31575 ( .A(n30780), .B(n30779), .Z(n30784) );
  NANDN U31576 ( .A(n30782), .B(n30781), .Z(n30783) );
  NAND U31577 ( .A(n30784), .B(n30783), .Z(n30945) );
  XNOR U31578 ( .A(n30944), .B(n30945), .Z(n30946) );
  NANDN U31579 ( .A(n30786), .B(n30785), .Z(n30790) );
  NAND U31580 ( .A(n30788), .B(n30787), .Z(n30789) );
  NAND U31581 ( .A(n30790), .B(n30789), .Z(n30947) );
  XNOR U31582 ( .A(n30946), .B(n30947), .Z(n31002) );
  XNOR U31583 ( .A(n31003), .B(n31002), .Z(n31005) );
  NAND U31584 ( .A(n30792), .B(n30791), .Z(n30796) );
  NAND U31585 ( .A(n30794), .B(n30793), .Z(n30795) );
  AND U31586 ( .A(n30796), .B(n30795), .Z(n31004) );
  XOR U31587 ( .A(n31005), .B(n31004), .Z(n31016) );
  NANDN U31588 ( .A(n30798), .B(n30797), .Z(n30802) );
  NANDN U31589 ( .A(n30800), .B(n30799), .Z(n30801) );
  AND U31590 ( .A(n30802), .B(n30801), .Z(n31014) );
  NANDN U31591 ( .A(n30808), .B(n30807), .Z(n30812) );
  OR U31592 ( .A(n30810), .B(n30809), .Z(n30811) );
  AND U31593 ( .A(n30812), .B(n30811), .Z(n31009) );
  NANDN U31594 ( .A(n30814), .B(n30813), .Z(n30818) );
  NANDN U31595 ( .A(n30816), .B(n30815), .Z(n30817) );
  AND U31596 ( .A(n30818), .B(n30817), .Z(n30951) );
  NANDN U31597 ( .A(n30820), .B(n30819), .Z(n30824) );
  OR U31598 ( .A(n30822), .B(n30821), .Z(n30823) );
  NAND U31599 ( .A(n30824), .B(n30823), .Z(n30950) );
  XNOR U31600 ( .A(n30951), .B(n30950), .Z(n30953) );
  NAND U31601 ( .A(n194), .B(n30825), .Z(n30827) );
  XOR U31602 ( .A(b[29]), .B(a[194]), .Z(n30975) );
  NAND U31603 ( .A(n38456), .B(n30975), .Z(n30826) );
  AND U31604 ( .A(n30827), .B(n30826), .Z(n30897) );
  AND U31605 ( .A(b[31]), .B(a[190]), .Z(n30896) );
  XNOR U31606 ( .A(n30897), .B(n30896), .Z(n30898) );
  NAND U31607 ( .A(b[0]), .B(a[222]), .Z(n30828) );
  XNOR U31608 ( .A(b[1]), .B(n30828), .Z(n30830) );
  NANDN U31609 ( .A(b[0]), .B(a[221]), .Z(n30829) );
  NAND U31610 ( .A(n30830), .B(n30829), .Z(n30899) );
  XNOR U31611 ( .A(n30898), .B(n30899), .Z(n30939) );
  NAND U31612 ( .A(n38185), .B(n30831), .Z(n30833) );
  XOR U31613 ( .A(b[23]), .B(a[200]), .Z(n30978) );
  NAND U31614 ( .A(n38132), .B(n30978), .Z(n30832) );
  AND U31615 ( .A(n30833), .B(n30832), .Z(n30968) );
  NAND U31616 ( .A(n184), .B(n30834), .Z(n30836) );
  XOR U31617 ( .A(b[7]), .B(a[216]), .Z(n30981) );
  NAND U31618 ( .A(n36592), .B(n30981), .Z(n30835) );
  AND U31619 ( .A(n30836), .B(n30835), .Z(n30967) );
  NAND U31620 ( .A(n38289), .B(n30837), .Z(n30839) );
  XOR U31621 ( .A(b[25]), .B(a[198]), .Z(n30984) );
  NAND U31622 ( .A(n38247), .B(n30984), .Z(n30838) );
  NAND U31623 ( .A(n30839), .B(n30838), .Z(n30966) );
  XOR U31624 ( .A(n30967), .B(n30966), .Z(n30969) );
  XOR U31625 ( .A(n30968), .B(n30969), .Z(n30938) );
  XOR U31626 ( .A(n30939), .B(n30938), .Z(n30941) );
  NAND U31627 ( .A(n187), .B(n30840), .Z(n30842) );
  XOR U31628 ( .A(b[13]), .B(a[210]), .Z(n30987) );
  NAND U31629 ( .A(n37295), .B(n30987), .Z(n30841) );
  AND U31630 ( .A(n30842), .B(n30841), .Z(n30933) );
  NAND U31631 ( .A(n186), .B(n30843), .Z(n30845) );
  XOR U31632 ( .A(b[11]), .B(a[212]), .Z(n30990) );
  NAND U31633 ( .A(n37097), .B(n30990), .Z(n30844) );
  NAND U31634 ( .A(n30845), .B(n30844), .Z(n30932) );
  XNOR U31635 ( .A(n30933), .B(n30932), .Z(n30935) );
  NAND U31636 ( .A(n188), .B(n30846), .Z(n30848) );
  XOR U31637 ( .A(b[15]), .B(a[208]), .Z(n30993) );
  NAND U31638 ( .A(n37382), .B(n30993), .Z(n30847) );
  AND U31639 ( .A(n30848), .B(n30847), .Z(n30929) );
  NAND U31640 ( .A(n38064), .B(n30849), .Z(n30851) );
  XOR U31641 ( .A(b[21]), .B(a[202]), .Z(n30996) );
  NAND U31642 ( .A(n37993), .B(n30996), .Z(n30850) );
  AND U31643 ( .A(n30851), .B(n30850), .Z(n30927) );
  NAND U31644 ( .A(n185), .B(n30852), .Z(n30854) );
  XOR U31645 ( .A(b[9]), .B(a[214]), .Z(n30999) );
  NAND U31646 ( .A(n36805), .B(n30999), .Z(n30853) );
  NAND U31647 ( .A(n30854), .B(n30853), .Z(n30926) );
  XNOR U31648 ( .A(n30927), .B(n30926), .Z(n30928) );
  XNOR U31649 ( .A(n30929), .B(n30928), .Z(n30934) );
  XOR U31650 ( .A(n30935), .B(n30934), .Z(n30940) );
  XNOR U31651 ( .A(n30941), .B(n30940), .Z(n30952) );
  XNOR U31652 ( .A(n30953), .B(n30952), .Z(n31008) );
  XNOR U31653 ( .A(n31009), .B(n31008), .Z(n31010) );
  XOR U31654 ( .A(n31011), .B(n31010), .Z(n31015) );
  XOR U31655 ( .A(n31014), .B(n31015), .Z(n31017) );
  XOR U31656 ( .A(n31016), .B(n31017), .Z(n30893) );
  NANDN U31657 ( .A(n30856), .B(n30855), .Z(n30860) );
  NAND U31658 ( .A(n30858), .B(n30857), .Z(n30859) );
  AND U31659 ( .A(n30860), .B(n30859), .Z(n30891) );
  NANDN U31660 ( .A(n30862), .B(n30861), .Z(n30866) );
  NANDN U31661 ( .A(n30864), .B(n30863), .Z(n30865) );
  AND U31662 ( .A(n30866), .B(n30865), .Z(n30890) );
  XNOR U31663 ( .A(n30891), .B(n30890), .Z(n30892) );
  XNOR U31664 ( .A(n30893), .B(n30892), .Z(n30884) );
  NANDN U31665 ( .A(n30868), .B(n30867), .Z(n30872) );
  NANDN U31666 ( .A(n30870), .B(n30869), .Z(n30871) );
  NAND U31667 ( .A(n30872), .B(n30871), .Z(n30885) );
  XOR U31668 ( .A(n30884), .B(n30885), .Z(n30887) );
  XNOR U31669 ( .A(n30886), .B(n30887), .Z(n30878) );
  XNOR U31670 ( .A(n30879), .B(n30878), .Z(n30880) );
  XNOR U31671 ( .A(n30881), .B(n30880), .Z(n31020) );
  XNOR U31672 ( .A(sreg[446]), .B(n31020), .Z(n31022) );
  NANDN U31673 ( .A(sreg[445]), .B(n30873), .Z(n30877) );
  NAND U31674 ( .A(n30875), .B(n30874), .Z(n30876) );
  NAND U31675 ( .A(n30877), .B(n30876), .Z(n31021) );
  XNOR U31676 ( .A(n31022), .B(n31021), .Z(c[446]) );
  NANDN U31677 ( .A(n30879), .B(n30878), .Z(n30883) );
  NANDN U31678 ( .A(n30881), .B(n30880), .Z(n30882) );
  AND U31679 ( .A(n30883), .B(n30882), .Z(n31028) );
  NANDN U31680 ( .A(n30885), .B(n30884), .Z(n30889) );
  NANDN U31681 ( .A(n30887), .B(n30886), .Z(n30888) );
  AND U31682 ( .A(n30889), .B(n30888), .Z(n31026) );
  NANDN U31683 ( .A(n30891), .B(n30890), .Z(n30895) );
  NANDN U31684 ( .A(n30893), .B(n30892), .Z(n30894) );
  AND U31685 ( .A(n30895), .B(n30894), .Z(n31034) );
  NANDN U31686 ( .A(n30897), .B(n30896), .Z(n30901) );
  NANDN U31687 ( .A(n30899), .B(n30898), .Z(n30900) );
  AND U31688 ( .A(n30901), .B(n30900), .Z(n31103) );
  NAND U31689 ( .A(n38385), .B(n30902), .Z(n30904) );
  XOR U31690 ( .A(b[27]), .B(a[197]), .Z(n31049) );
  NAND U31691 ( .A(n38343), .B(n31049), .Z(n30903) );
  AND U31692 ( .A(n30904), .B(n30903), .Z(n31110) );
  NAND U31693 ( .A(n183), .B(n30905), .Z(n30907) );
  XOR U31694 ( .A(b[5]), .B(a[219]), .Z(n31052) );
  NAND U31695 ( .A(n36296), .B(n31052), .Z(n30906) );
  AND U31696 ( .A(n30907), .B(n30906), .Z(n31108) );
  NAND U31697 ( .A(n190), .B(n30908), .Z(n30910) );
  XOR U31698 ( .A(b[19]), .B(a[205]), .Z(n31055) );
  NAND U31699 ( .A(n37821), .B(n31055), .Z(n30909) );
  NAND U31700 ( .A(n30910), .B(n30909), .Z(n31107) );
  XNOR U31701 ( .A(n31108), .B(n31107), .Z(n31109) );
  XNOR U31702 ( .A(n31110), .B(n31109), .Z(n31101) );
  NAND U31703 ( .A(n38470), .B(n30911), .Z(n30913) );
  XOR U31704 ( .A(b[31]), .B(a[193]), .Z(n31058) );
  NAND U31705 ( .A(n38453), .B(n31058), .Z(n30912) );
  AND U31706 ( .A(n30913), .B(n30912), .Z(n31070) );
  NAND U31707 ( .A(n181), .B(n30914), .Z(n30916) );
  XOR U31708 ( .A(b[3]), .B(a[221]), .Z(n31061) );
  NAND U31709 ( .A(n182), .B(n31061), .Z(n30915) );
  AND U31710 ( .A(n30916), .B(n30915), .Z(n31068) );
  NAND U31711 ( .A(n189), .B(n30917), .Z(n30919) );
  XOR U31712 ( .A(b[17]), .B(a[207]), .Z(n31064) );
  NAND U31713 ( .A(n37652), .B(n31064), .Z(n30918) );
  NAND U31714 ( .A(n30919), .B(n30918), .Z(n31067) );
  XNOR U31715 ( .A(n31068), .B(n31067), .Z(n31069) );
  XOR U31716 ( .A(n31070), .B(n31069), .Z(n31102) );
  XOR U31717 ( .A(n31101), .B(n31102), .Z(n31104) );
  XOR U31718 ( .A(n31103), .B(n31104), .Z(n31150) );
  NANDN U31719 ( .A(n30921), .B(n30920), .Z(n30925) );
  NANDN U31720 ( .A(n30923), .B(n30922), .Z(n30924) );
  AND U31721 ( .A(n30925), .B(n30924), .Z(n31091) );
  NANDN U31722 ( .A(n30927), .B(n30926), .Z(n30931) );
  NANDN U31723 ( .A(n30929), .B(n30928), .Z(n30930) );
  NAND U31724 ( .A(n30931), .B(n30930), .Z(n31092) );
  XNOR U31725 ( .A(n31091), .B(n31092), .Z(n31093) );
  NANDN U31726 ( .A(n30933), .B(n30932), .Z(n30937) );
  NAND U31727 ( .A(n30935), .B(n30934), .Z(n30936) );
  NAND U31728 ( .A(n30937), .B(n30936), .Z(n31094) );
  XNOR U31729 ( .A(n31093), .B(n31094), .Z(n31149) );
  XNOR U31730 ( .A(n31150), .B(n31149), .Z(n31152) );
  NAND U31731 ( .A(n30939), .B(n30938), .Z(n30943) );
  NAND U31732 ( .A(n30941), .B(n30940), .Z(n30942) );
  AND U31733 ( .A(n30943), .B(n30942), .Z(n31151) );
  XOR U31734 ( .A(n31152), .B(n31151), .Z(n31163) );
  NANDN U31735 ( .A(n30945), .B(n30944), .Z(n30949) );
  NANDN U31736 ( .A(n30947), .B(n30946), .Z(n30948) );
  AND U31737 ( .A(n30949), .B(n30948), .Z(n31161) );
  NANDN U31738 ( .A(n30955), .B(n30954), .Z(n30959) );
  OR U31739 ( .A(n30957), .B(n30956), .Z(n30958) );
  AND U31740 ( .A(n30959), .B(n30958), .Z(n31156) );
  NANDN U31741 ( .A(n30961), .B(n30960), .Z(n30965) );
  NANDN U31742 ( .A(n30963), .B(n30962), .Z(n30964) );
  AND U31743 ( .A(n30965), .B(n30964), .Z(n31098) );
  NANDN U31744 ( .A(n30967), .B(n30966), .Z(n30971) );
  OR U31745 ( .A(n30969), .B(n30968), .Z(n30970) );
  NAND U31746 ( .A(n30971), .B(n30970), .Z(n31097) );
  XNOR U31747 ( .A(n31098), .B(n31097), .Z(n31100) );
  NAND U31748 ( .A(b[0]), .B(a[223]), .Z(n30972) );
  XNOR U31749 ( .A(b[1]), .B(n30972), .Z(n30974) );
  NANDN U31750 ( .A(b[0]), .B(a[222]), .Z(n30973) );
  NAND U31751 ( .A(n30974), .B(n30973), .Z(n31046) );
  NAND U31752 ( .A(n194), .B(n30975), .Z(n30977) );
  XOR U31753 ( .A(b[29]), .B(a[195]), .Z(n31122) );
  NAND U31754 ( .A(n38456), .B(n31122), .Z(n30976) );
  AND U31755 ( .A(n30977), .B(n30976), .Z(n31044) );
  AND U31756 ( .A(b[31]), .B(a[191]), .Z(n31043) );
  XNOR U31757 ( .A(n31044), .B(n31043), .Z(n31045) );
  XNOR U31758 ( .A(n31046), .B(n31045), .Z(n31086) );
  NAND U31759 ( .A(n38185), .B(n30978), .Z(n30980) );
  XOR U31760 ( .A(b[23]), .B(a[201]), .Z(n31125) );
  NAND U31761 ( .A(n38132), .B(n31125), .Z(n30979) );
  AND U31762 ( .A(n30980), .B(n30979), .Z(n31115) );
  NAND U31763 ( .A(n184), .B(n30981), .Z(n30983) );
  XOR U31764 ( .A(b[7]), .B(a[217]), .Z(n31128) );
  NAND U31765 ( .A(n36592), .B(n31128), .Z(n30982) );
  AND U31766 ( .A(n30983), .B(n30982), .Z(n31114) );
  NAND U31767 ( .A(n38289), .B(n30984), .Z(n30986) );
  XOR U31768 ( .A(b[25]), .B(a[199]), .Z(n31131) );
  NAND U31769 ( .A(n38247), .B(n31131), .Z(n30985) );
  NAND U31770 ( .A(n30986), .B(n30985), .Z(n31113) );
  XOR U31771 ( .A(n31114), .B(n31113), .Z(n31116) );
  XOR U31772 ( .A(n31115), .B(n31116), .Z(n31085) );
  XOR U31773 ( .A(n31086), .B(n31085), .Z(n31088) );
  NAND U31774 ( .A(n187), .B(n30987), .Z(n30989) );
  XOR U31775 ( .A(b[13]), .B(a[211]), .Z(n31134) );
  NAND U31776 ( .A(n37295), .B(n31134), .Z(n30988) );
  AND U31777 ( .A(n30989), .B(n30988), .Z(n31080) );
  NAND U31778 ( .A(n186), .B(n30990), .Z(n30992) );
  XOR U31779 ( .A(b[11]), .B(a[213]), .Z(n31137) );
  NAND U31780 ( .A(n37097), .B(n31137), .Z(n30991) );
  NAND U31781 ( .A(n30992), .B(n30991), .Z(n31079) );
  XNOR U31782 ( .A(n31080), .B(n31079), .Z(n31082) );
  NAND U31783 ( .A(n188), .B(n30993), .Z(n30995) );
  XOR U31784 ( .A(b[15]), .B(a[209]), .Z(n31140) );
  NAND U31785 ( .A(n37382), .B(n31140), .Z(n30994) );
  AND U31786 ( .A(n30995), .B(n30994), .Z(n31076) );
  NAND U31787 ( .A(n38064), .B(n30996), .Z(n30998) );
  XOR U31788 ( .A(b[21]), .B(a[203]), .Z(n31143) );
  NAND U31789 ( .A(n37993), .B(n31143), .Z(n30997) );
  AND U31790 ( .A(n30998), .B(n30997), .Z(n31074) );
  NAND U31791 ( .A(n185), .B(n30999), .Z(n31001) );
  XOR U31792 ( .A(b[9]), .B(a[215]), .Z(n31146) );
  NAND U31793 ( .A(n36805), .B(n31146), .Z(n31000) );
  NAND U31794 ( .A(n31001), .B(n31000), .Z(n31073) );
  XNOR U31795 ( .A(n31074), .B(n31073), .Z(n31075) );
  XNOR U31796 ( .A(n31076), .B(n31075), .Z(n31081) );
  XOR U31797 ( .A(n31082), .B(n31081), .Z(n31087) );
  XNOR U31798 ( .A(n31088), .B(n31087), .Z(n31099) );
  XNOR U31799 ( .A(n31100), .B(n31099), .Z(n31155) );
  XNOR U31800 ( .A(n31156), .B(n31155), .Z(n31157) );
  XOR U31801 ( .A(n31158), .B(n31157), .Z(n31162) );
  XOR U31802 ( .A(n31161), .B(n31162), .Z(n31164) );
  XOR U31803 ( .A(n31163), .B(n31164), .Z(n31040) );
  NANDN U31804 ( .A(n31003), .B(n31002), .Z(n31007) );
  NAND U31805 ( .A(n31005), .B(n31004), .Z(n31006) );
  AND U31806 ( .A(n31007), .B(n31006), .Z(n31038) );
  NANDN U31807 ( .A(n31009), .B(n31008), .Z(n31013) );
  NANDN U31808 ( .A(n31011), .B(n31010), .Z(n31012) );
  AND U31809 ( .A(n31013), .B(n31012), .Z(n31037) );
  XNOR U31810 ( .A(n31038), .B(n31037), .Z(n31039) );
  XNOR U31811 ( .A(n31040), .B(n31039), .Z(n31031) );
  NANDN U31812 ( .A(n31015), .B(n31014), .Z(n31019) );
  OR U31813 ( .A(n31017), .B(n31016), .Z(n31018) );
  NAND U31814 ( .A(n31019), .B(n31018), .Z(n31032) );
  XNOR U31815 ( .A(n31031), .B(n31032), .Z(n31033) );
  XNOR U31816 ( .A(n31034), .B(n31033), .Z(n31025) );
  XNOR U31817 ( .A(n31026), .B(n31025), .Z(n31027) );
  XNOR U31818 ( .A(n31028), .B(n31027), .Z(n31167) );
  XNOR U31819 ( .A(sreg[447]), .B(n31167), .Z(n31169) );
  NANDN U31820 ( .A(sreg[446]), .B(n31020), .Z(n31024) );
  NAND U31821 ( .A(n31022), .B(n31021), .Z(n31023) );
  NAND U31822 ( .A(n31024), .B(n31023), .Z(n31168) );
  XNOR U31823 ( .A(n31169), .B(n31168), .Z(c[447]) );
  NANDN U31824 ( .A(n31026), .B(n31025), .Z(n31030) );
  NANDN U31825 ( .A(n31028), .B(n31027), .Z(n31029) );
  AND U31826 ( .A(n31030), .B(n31029), .Z(n31175) );
  NANDN U31827 ( .A(n31032), .B(n31031), .Z(n31036) );
  NANDN U31828 ( .A(n31034), .B(n31033), .Z(n31035) );
  AND U31829 ( .A(n31036), .B(n31035), .Z(n31173) );
  NANDN U31830 ( .A(n31038), .B(n31037), .Z(n31042) );
  NANDN U31831 ( .A(n31040), .B(n31039), .Z(n31041) );
  AND U31832 ( .A(n31042), .B(n31041), .Z(n31181) );
  NANDN U31833 ( .A(n31044), .B(n31043), .Z(n31048) );
  NANDN U31834 ( .A(n31046), .B(n31045), .Z(n31047) );
  AND U31835 ( .A(n31048), .B(n31047), .Z(n31252) );
  NAND U31836 ( .A(n38385), .B(n31049), .Z(n31051) );
  XOR U31837 ( .A(b[27]), .B(a[198]), .Z(n31196) );
  NAND U31838 ( .A(n38343), .B(n31196), .Z(n31050) );
  AND U31839 ( .A(n31051), .B(n31050), .Z(n31259) );
  NAND U31840 ( .A(n183), .B(n31052), .Z(n31054) );
  XOR U31841 ( .A(b[5]), .B(a[220]), .Z(n31199) );
  NAND U31842 ( .A(n36296), .B(n31199), .Z(n31053) );
  AND U31843 ( .A(n31054), .B(n31053), .Z(n31257) );
  NAND U31844 ( .A(n190), .B(n31055), .Z(n31057) );
  XOR U31845 ( .A(b[19]), .B(a[206]), .Z(n31202) );
  NAND U31846 ( .A(n37821), .B(n31202), .Z(n31056) );
  NAND U31847 ( .A(n31057), .B(n31056), .Z(n31256) );
  XNOR U31848 ( .A(n31257), .B(n31256), .Z(n31258) );
  XNOR U31849 ( .A(n31259), .B(n31258), .Z(n31250) );
  NAND U31850 ( .A(n38470), .B(n31058), .Z(n31060) );
  XOR U31851 ( .A(b[31]), .B(a[194]), .Z(n31205) );
  NAND U31852 ( .A(n38453), .B(n31205), .Z(n31059) );
  AND U31853 ( .A(n31060), .B(n31059), .Z(n31217) );
  NAND U31854 ( .A(n181), .B(n31061), .Z(n31063) );
  XOR U31855 ( .A(b[3]), .B(a[222]), .Z(n31208) );
  NAND U31856 ( .A(n182), .B(n31208), .Z(n31062) );
  AND U31857 ( .A(n31063), .B(n31062), .Z(n31215) );
  NAND U31858 ( .A(n189), .B(n31064), .Z(n31066) );
  XOR U31859 ( .A(b[17]), .B(a[208]), .Z(n31211) );
  NAND U31860 ( .A(n37652), .B(n31211), .Z(n31065) );
  NAND U31861 ( .A(n31066), .B(n31065), .Z(n31214) );
  XNOR U31862 ( .A(n31215), .B(n31214), .Z(n31216) );
  XOR U31863 ( .A(n31217), .B(n31216), .Z(n31251) );
  XOR U31864 ( .A(n31250), .B(n31251), .Z(n31253) );
  XOR U31865 ( .A(n31252), .B(n31253), .Z(n31299) );
  NANDN U31866 ( .A(n31068), .B(n31067), .Z(n31072) );
  NANDN U31867 ( .A(n31070), .B(n31069), .Z(n31071) );
  AND U31868 ( .A(n31072), .B(n31071), .Z(n31238) );
  NANDN U31869 ( .A(n31074), .B(n31073), .Z(n31078) );
  NANDN U31870 ( .A(n31076), .B(n31075), .Z(n31077) );
  NAND U31871 ( .A(n31078), .B(n31077), .Z(n31239) );
  XNOR U31872 ( .A(n31238), .B(n31239), .Z(n31240) );
  NANDN U31873 ( .A(n31080), .B(n31079), .Z(n31084) );
  NAND U31874 ( .A(n31082), .B(n31081), .Z(n31083) );
  NAND U31875 ( .A(n31084), .B(n31083), .Z(n31241) );
  XNOR U31876 ( .A(n31240), .B(n31241), .Z(n31298) );
  XNOR U31877 ( .A(n31299), .B(n31298), .Z(n31301) );
  NAND U31878 ( .A(n31086), .B(n31085), .Z(n31090) );
  NAND U31879 ( .A(n31088), .B(n31087), .Z(n31089) );
  AND U31880 ( .A(n31090), .B(n31089), .Z(n31300) );
  XOR U31881 ( .A(n31301), .B(n31300), .Z(n31312) );
  NANDN U31882 ( .A(n31092), .B(n31091), .Z(n31096) );
  NANDN U31883 ( .A(n31094), .B(n31093), .Z(n31095) );
  AND U31884 ( .A(n31096), .B(n31095), .Z(n31310) );
  NANDN U31885 ( .A(n31102), .B(n31101), .Z(n31106) );
  OR U31886 ( .A(n31104), .B(n31103), .Z(n31105) );
  AND U31887 ( .A(n31106), .B(n31105), .Z(n31305) );
  NANDN U31888 ( .A(n31108), .B(n31107), .Z(n31112) );
  NANDN U31889 ( .A(n31110), .B(n31109), .Z(n31111) );
  AND U31890 ( .A(n31112), .B(n31111), .Z(n31245) );
  NANDN U31891 ( .A(n31114), .B(n31113), .Z(n31118) );
  OR U31892 ( .A(n31116), .B(n31115), .Z(n31117) );
  NAND U31893 ( .A(n31118), .B(n31117), .Z(n31244) );
  XNOR U31894 ( .A(n31245), .B(n31244), .Z(n31246) );
  NAND U31895 ( .A(b[0]), .B(a[224]), .Z(n31119) );
  XNOR U31896 ( .A(b[1]), .B(n31119), .Z(n31121) );
  NANDN U31897 ( .A(b[0]), .B(a[223]), .Z(n31120) );
  NAND U31898 ( .A(n31121), .B(n31120), .Z(n31193) );
  NAND U31899 ( .A(n194), .B(n31122), .Z(n31124) );
  XOR U31900 ( .A(b[29]), .B(a[196]), .Z(n31271) );
  NAND U31901 ( .A(n38456), .B(n31271), .Z(n31123) );
  AND U31902 ( .A(n31124), .B(n31123), .Z(n31191) );
  AND U31903 ( .A(b[31]), .B(a[192]), .Z(n31190) );
  XNOR U31904 ( .A(n31191), .B(n31190), .Z(n31192) );
  XNOR U31905 ( .A(n31193), .B(n31192), .Z(n31232) );
  NAND U31906 ( .A(n38185), .B(n31125), .Z(n31127) );
  XOR U31907 ( .A(b[23]), .B(a[202]), .Z(n31274) );
  NAND U31908 ( .A(n38132), .B(n31274), .Z(n31126) );
  AND U31909 ( .A(n31127), .B(n31126), .Z(n31265) );
  NAND U31910 ( .A(n184), .B(n31128), .Z(n31130) );
  XOR U31911 ( .A(b[7]), .B(a[218]), .Z(n31277) );
  NAND U31912 ( .A(n36592), .B(n31277), .Z(n31129) );
  AND U31913 ( .A(n31130), .B(n31129), .Z(n31263) );
  NAND U31914 ( .A(n38289), .B(n31131), .Z(n31133) );
  XOR U31915 ( .A(b[25]), .B(a[200]), .Z(n31280) );
  NAND U31916 ( .A(n38247), .B(n31280), .Z(n31132) );
  NAND U31917 ( .A(n31133), .B(n31132), .Z(n31262) );
  XNOR U31918 ( .A(n31263), .B(n31262), .Z(n31264) );
  XOR U31919 ( .A(n31265), .B(n31264), .Z(n31233) );
  XNOR U31920 ( .A(n31232), .B(n31233), .Z(n31234) );
  NAND U31921 ( .A(n187), .B(n31134), .Z(n31136) );
  XOR U31922 ( .A(b[13]), .B(a[212]), .Z(n31283) );
  NAND U31923 ( .A(n37295), .B(n31283), .Z(n31135) );
  AND U31924 ( .A(n31136), .B(n31135), .Z(n31227) );
  NAND U31925 ( .A(n186), .B(n31137), .Z(n31139) );
  XOR U31926 ( .A(b[11]), .B(a[214]), .Z(n31286) );
  NAND U31927 ( .A(n37097), .B(n31286), .Z(n31138) );
  NAND U31928 ( .A(n31139), .B(n31138), .Z(n31226) );
  XNOR U31929 ( .A(n31227), .B(n31226), .Z(n31228) );
  NAND U31930 ( .A(n188), .B(n31140), .Z(n31142) );
  XOR U31931 ( .A(b[15]), .B(a[210]), .Z(n31289) );
  NAND U31932 ( .A(n37382), .B(n31289), .Z(n31141) );
  AND U31933 ( .A(n31142), .B(n31141), .Z(n31223) );
  NAND U31934 ( .A(n38064), .B(n31143), .Z(n31145) );
  XOR U31935 ( .A(b[21]), .B(a[204]), .Z(n31292) );
  NAND U31936 ( .A(n37993), .B(n31292), .Z(n31144) );
  AND U31937 ( .A(n31145), .B(n31144), .Z(n31221) );
  NAND U31938 ( .A(n185), .B(n31146), .Z(n31148) );
  XOR U31939 ( .A(b[9]), .B(a[216]), .Z(n31295) );
  NAND U31940 ( .A(n36805), .B(n31295), .Z(n31147) );
  NAND U31941 ( .A(n31148), .B(n31147), .Z(n31220) );
  XNOR U31942 ( .A(n31221), .B(n31220), .Z(n31222) );
  XOR U31943 ( .A(n31223), .B(n31222), .Z(n31229) );
  XOR U31944 ( .A(n31228), .B(n31229), .Z(n31235) );
  XOR U31945 ( .A(n31234), .B(n31235), .Z(n31247) );
  XNOR U31946 ( .A(n31246), .B(n31247), .Z(n31304) );
  XNOR U31947 ( .A(n31305), .B(n31304), .Z(n31306) );
  XOR U31948 ( .A(n31307), .B(n31306), .Z(n31311) );
  XOR U31949 ( .A(n31310), .B(n31311), .Z(n31313) );
  XOR U31950 ( .A(n31312), .B(n31313), .Z(n31187) );
  NANDN U31951 ( .A(n31150), .B(n31149), .Z(n31154) );
  NAND U31952 ( .A(n31152), .B(n31151), .Z(n31153) );
  AND U31953 ( .A(n31154), .B(n31153), .Z(n31185) );
  NANDN U31954 ( .A(n31156), .B(n31155), .Z(n31160) );
  NANDN U31955 ( .A(n31158), .B(n31157), .Z(n31159) );
  AND U31956 ( .A(n31160), .B(n31159), .Z(n31184) );
  XNOR U31957 ( .A(n31185), .B(n31184), .Z(n31186) );
  XNOR U31958 ( .A(n31187), .B(n31186), .Z(n31178) );
  NANDN U31959 ( .A(n31162), .B(n31161), .Z(n31166) );
  OR U31960 ( .A(n31164), .B(n31163), .Z(n31165) );
  NAND U31961 ( .A(n31166), .B(n31165), .Z(n31179) );
  XNOR U31962 ( .A(n31178), .B(n31179), .Z(n31180) );
  XNOR U31963 ( .A(n31181), .B(n31180), .Z(n31172) );
  XNOR U31964 ( .A(n31173), .B(n31172), .Z(n31174) );
  XNOR U31965 ( .A(n31175), .B(n31174), .Z(n31316) );
  XNOR U31966 ( .A(sreg[448]), .B(n31316), .Z(n31318) );
  NANDN U31967 ( .A(sreg[447]), .B(n31167), .Z(n31171) );
  NAND U31968 ( .A(n31169), .B(n31168), .Z(n31170) );
  NAND U31969 ( .A(n31171), .B(n31170), .Z(n31317) );
  XNOR U31970 ( .A(n31318), .B(n31317), .Z(c[448]) );
  NANDN U31971 ( .A(n31173), .B(n31172), .Z(n31177) );
  NANDN U31972 ( .A(n31175), .B(n31174), .Z(n31176) );
  AND U31973 ( .A(n31177), .B(n31176), .Z(n31324) );
  NANDN U31974 ( .A(n31179), .B(n31178), .Z(n31183) );
  NANDN U31975 ( .A(n31181), .B(n31180), .Z(n31182) );
  AND U31976 ( .A(n31183), .B(n31182), .Z(n31322) );
  NANDN U31977 ( .A(n31185), .B(n31184), .Z(n31189) );
  NANDN U31978 ( .A(n31187), .B(n31186), .Z(n31188) );
  AND U31979 ( .A(n31189), .B(n31188), .Z(n31330) );
  NANDN U31980 ( .A(n31191), .B(n31190), .Z(n31195) );
  NANDN U31981 ( .A(n31193), .B(n31192), .Z(n31194) );
  AND U31982 ( .A(n31195), .B(n31194), .Z(n31413) );
  NAND U31983 ( .A(n38385), .B(n31196), .Z(n31198) );
  XOR U31984 ( .A(b[27]), .B(a[199]), .Z(n31357) );
  NAND U31985 ( .A(n38343), .B(n31357), .Z(n31197) );
  AND U31986 ( .A(n31198), .B(n31197), .Z(n31420) );
  NAND U31987 ( .A(n183), .B(n31199), .Z(n31201) );
  XOR U31988 ( .A(b[5]), .B(a[221]), .Z(n31360) );
  NAND U31989 ( .A(n36296), .B(n31360), .Z(n31200) );
  AND U31990 ( .A(n31201), .B(n31200), .Z(n31418) );
  NAND U31991 ( .A(n190), .B(n31202), .Z(n31204) );
  XOR U31992 ( .A(b[19]), .B(a[207]), .Z(n31363) );
  NAND U31993 ( .A(n37821), .B(n31363), .Z(n31203) );
  NAND U31994 ( .A(n31204), .B(n31203), .Z(n31417) );
  XNOR U31995 ( .A(n31418), .B(n31417), .Z(n31419) );
  XNOR U31996 ( .A(n31420), .B(n31419), .Z(n31411) );
  NAND U31997 ( .A(n38470), .B(n31205), .Z(n31207) );
  XOR U31998 ( .A(b[31]), .B(a[195]), .Z(n31366) );
  NAND U31999 ( .A(n38453), .B(n31366), .Z(n31206) );
  AND U32000 ( .A(n31207), .B(n31206), .Z(n31378) );
  NAND U32001 ( .A(n181), .B(n31208), .Z(n31210) );
  XOR U32002 ( .A(b[3]), .B(a[223]), .Z(n31369) );
  NAND U32003 ( .A(n182), .B(n31369), .Z(n31209) );
  AND U32004 ( .A(n31210), .B(n31209), .Z(n31376) );
  NAND U32005 ( .A(n189), .B(n31211), .Z(n31213) );
  XOR U32006 ( .A(b[17]), .B(a[209]), .Z(n31372) );
  NAND U32007 ( .A(n37652), .B(n31372), .Z(n31212) );
  NAND U32008 ( .A(n31213), .B(n31212), .Z(n31375) );
  XNOR U32009 ( .A(n31376), .B(n31375), .Z(n31377) );
  XOR U32010 ( .A(n31378), .B(n31377), .Z(n31412) );
  XOR U32011 ( .A(n31411), .B(n31412), .Z(n31414) );
  XOR U32012 ( .A(n31413), .B(n31414), .Z(n31346) );
  NANDN U32013 ( .A(n31215), .B(n31214), .Z(n31219) );
  NANDN U32014 ( .A(n31217), .B(n31216), .Z(n31218) );
  AND U32015 ( .A(n31219), .B(n31218), .Z(n31399) );
  NANDN U32016 ( .A(n31221), .B(n31220), .Z(n31225) );
  NANDN U32017 ( .A(n31223), .B(n31222), .Z(n31224) );
  NAND U32018 ( .A(n31225), .B(n31224), .Z(n31400) );
  XNOR U32019 ( .A(n31399), .B(n31400), .Z(n31401) );
  NANDN U32020 ( .A(n31227), .B(n31226), .Z(n31231) );
  NANDN U32021 ( .A(n31229), .B(n31228), .Z(n31230) );
  NAND U32022 ( .A(n31231), .B(n31230), .Z(n31402) );
  XNOR U32023 ( .A(n31401), .B(n31402), .Z(n31345) );
  XNOR U32024 ( .A(n31346), .B(n31345), .Z(n31348) );
  NANDN U32025 ( .A(n31233), .B(n31232), .Z(n31237) );
  NANDN U32026 ( .A(n31235), .B(n31234), .Z(n31236) );
  AND U32027 ( .A(n31237), .B(n31236), .Z(n31347) );
  XOR U32028 ( .A(n31348), .B(n31347), .Z(n31461) );
  NANDN U32029 ( .A(n31239), .B(n31238), .Z(n31243) );
  NANDN U32030 ( .A(n31241), .B(n31240), .Z(n31242) );
  AND U32031 ( .A(n31243), .B(n31242), .Z(n31459) );
  NANDN U32032 ( .A(n31245), .B(n31244), .Z(n31249) );
  NANDN U32033 ( .A(n31247), .B(n31246), .Z(n31248) );
  AND U32034 ( .A(n31249), .B(n31248), .Z(n31342) );
  NANDN U32035 ( .A(n31251), .B(n31250), .Z(n31255) );
  OR U32036 ( .A(n31253), .B(n31252), .Z(n31254) );
  AND U32037 ( .A(n31255), .B(n31254), .Z(n31340) );
  NANDN U32038 ( .A(n31257), .B(n31256), .Z(n31261) );
  NANDN U32039 ( .A(n31259), .B(n31258), .Z(n31260) );
  AND U32040 ( .A(n31261), .B(n31260), .Z(n31406) );
  NANDN U32041 ( .A(n31263), .B(n31262), .Z(n31267) );
  NANDN U32042 ( .A(n31265), .B(n31264), .Z(n31266) );
  NAND U32043 ( .A(n31267), .B(n31266), .Z(n31405) );
  XNOR U32044 ( .A(n31406), .B(n31405), .Z(n31407) );
  NAND U32045 ( .A(b[0]), .B(a[225]), .Z(n31268) );
  XNOR U32046 ( .A(b[1]), .B(n31268), .Z(n31270) );
  NANDN U32047 ( .A(b[0]), .B(a[224]), .Z(n31269) );
  NAND U32048 ( .A(n31270), .B(n31269), .Z(n31354) );
  NAND U32049 ( .A(n194), .B(n31271), .Z(n31273) );
  XOR U32050 ( .A(b[29]), .B(a[197]), .Z(n31432) );
  NAND U32051 ( .A(n38456), .B(n31432), .Z(n31272) );
  AND U32052 ( .A(n31273), .B(n31272), .Z(n31352) );
  AND U32053 ( .A(b[31]), .B(a[193]), .Z(n31351) );
  XNOR U32054 ( .A(n31352), .B(n31351), .Z(n31353) );
  XNOR U32055 ( .A(n31354), .B(n31353), .Z(n31393) );
  NAND U32056 ( .A(n38185), .B(n31274), .Z(n31276) );
  XOR U32057 ( .A(b[23]), .B(a[203]), .Z(n31435) );
  NAND U32058 ( .A(n38132), .B(n31435), .Z(n31275) );
  AND U32059 ( .A(n31276), .B(n31275), .Z(n31426) );
  NAND U32060 ( .A(n184), .B(n31277), .Z(n31279) );
  XOR U32061 ( .A(b[7]), .B(a[219]), .Z(n31438) );
  NAND U32062 ( .A(n36592), .B(n31438), .Z(n31278) );
  AND U32063 ( .A(n31279), .B(n31278), .Z(n31424) );
  NAND U32064 ( .A(n38289), .B(n31280), .Z(n31282) );
  XOR U32065 ( .A(b[25]), .B(a[201]), .Z(n31441) );
  NAND U32066 ( .A(n38247), .B(n31441), .Z(n31281) );
  NAND U32067 ( .A(n31282), .B(n31281), .Z(n31423) );
  XNOR U32068 ( .A(n31424), .B(n31423), .Z(n31425) );
  XOR U32069 ( .A(n31426), .B(n31425), .Z(n31394) );
  XNOR U32070 ( .A(n31393), .B(n31394), .Z(n31395) );
  NAND U32071 ( .A(n187), .B(n31283), .Z(n31285) );
  XOR U32072 ( .A(b[13]), .B(a[213]), .Z(n31444) );
  NAND U32073 ( .A(n37295), .B(n31444), .Z(n31284) );
  AND U32074 ( .A(n31285), .B(n31284), .Z(n31388) );
  NAND U32075 ( .A(n186), .B(n31286), .Z(n31288) );
  XOR U32076 ( .A(b[11]), .B(a[215]), .Z(n31447) );
  NAND U32077 ( .A(n37097), .B(n31447), .Z(n31287) );
  NAND U32078 ( .A(n31288), .B(n31287), .Z(n31387) );
  XNOR U32079 ( .A(n31388), .B(n31387), .Z(n31389) );
  NAND U32080 ( .A(n188), .B(n31289), .Z(n31291) );
  XOR U32081 ( .A(b[15]), .B(a[211]), .Z(n31450) );
  NAND U32082 ( .A(n37382), .B(n31450), .Z(n31290) );
  AND U32083 ( .A(n31291), .B(n31290), .Z(n31384) );
  NAND U32084 ( .A(n38064), .B(n31292), .Z(n31294) );
  XOR U32085 ( .A(b[21]), .B(a[205]), .Z(n31453) );
  NAND U32086 ( .A(n37993), .B(n31453), .Z(n31293) );
  AND U32087 ( .A(n31294), .B(n31293), .Z(n31382) );
  NAND U32088 ( .A(n185), .B(n31295), .Z(n31297) );
  XOR U32089 ( .A(b[9]), .B(a[217]), .Z(n31456) );
  NAND U32090 ( .A(n36805), .B(n31456), .Z(n31296) );
  NAND U32091 ( .A(n31297), .B(n31296), .Z(n31381) );
  XNOR U32092 ( .A(n31382), .B(n31381), .Z(n31383) );
  XOR U32093 ( .A(n31384), .B(n31383), .Z(n31390) );
  XOR U32094 ( .A(n31389), .B(n31390), .Z(n31396) );
  XOR U32095 ( .A(n31395), .B(n31396), .Z(n31408) );
  XNOR U32096 ( .A(n31407), .B(n31408), .Z(n31339) );
  XNOR U32097 ( .A(n31340), .B(n31339), .Z(n31341) );
  XOR U32098 ( .A(n31342), .B(n31341), .Z(n31460) );
  XOR U32099 ( .A(n31459), .B(n31460), .Z(n31462) );
  XOR U32100 ( .A(n31461), .B(n31462), .Z(n31336) );
  NANDN U32101 ( .A(n31299), .B(n31298), .Z(n31303) );
  NAND U32102 ( .A(n31301), .B(n31300), .Z(n31302) );
  AND U32103 ( .A(n31303), .B(n31302), .Z(n31334) );
  NANDN U32104 ( .A(n31305), .B(n31304), .Z(n31309) );
  NANDN U32105 ( .A(n31307), .B(n31306), .Z(n31308) );
  AND U32106 ( .A(n31309), .B(n31308), .Z(n31333) );
  XNOR U32107 ( .A(n31334), .B(n31333), .Z(n31335) );
  XNOR U32108 ( .A(n31336), .B(n31335), .Z(n31327) );
  NANDN U32109 ( .A(n31311), .B(n31310), .Z(n31315) );
  OR U32110 ( .A(n31313), .B(n31312), .Z(n31314) );
  NAND U32111 ( .A(n31315), .B(n31314), .Z(n31328) );
  XNOR U32112 ( .A(n31327), .B(n31328), .Z(n31329) );
  XNOR U32113 ( .A(n31330), .B(n31329), .Z(n31321) );
  XNOR U32114 ( .A(n31322), .B(n31321), .Z(n31323) );
  XNOR U32115 ( .A(n31324), .B(n31323), .Z(n31465) );
  XNOR U32116 ( .A(sreg[449]), .B(n31465), .Z(n31467) );
  NANDN U32117 ( .A(sreg[448]), .B(n31316), .Z(n31320) );
  NAND U32118 ( .A(n31318), .B(n31317), .Z(n31319) );
  NAND U32119 ( .A(n31320), .B(n31319), .Z(n31466) );
  XNOR U32120 ( .A(n31467), .B(n31466), .Z(c[449]) );
  NANDN U32121 ( .A(n31322), .B(n31321), .Z(n31326) );
  NANDN U32122 ( .A(n31324), .B(n31323), .Z(n31325) );
  AND U32123 ( .A(n31326), .B(n31325), .Z(n31473) );
  NANDN U32124 ( .A(n31328), .B(n31327), .Z(n31332) );
  NANDN U32125 ( .A(n31330), .B(n31329), .Z(n31331) );
  AND U32126 ( .A(n31332), .B(n31331), .Z(n31471) );
  NANDN U32127 ( .A(n31334), .B(n31333), .Z(n31338) );
  NANDN U32128 ( .A(n31336), .B(n31335), .Z(n31337) );
  AND U32129 ( .A(n31338), .B(n31337), .Z(n31479) );
  NANDN U32130 ( .A(n31340), .B(n31339), .Z(n31344) );
  NANDN U32131 ( .A(n31342), .B(n31341), .Z(n31343) );
  AND U32132 ( .A(n31344), .B(n31343), .Z(n31483) );
  NANDN U32133 ( .A(n31346), .B(n31345), .Z(n31350) );
  NAND U32134 ( .A(n31348), .B(n31347), .Z(n31349) );
  AND U32135 ( .A(n31350), .B(n31349), .Z(n31482) );
  XNOR U32136 ( .A(n31483), .B(n31482), .Z(n31485) );
  NANDN U32137 ( .A(n31352), .B(n31351), .Z(n31356) );
  NANDN U32138 ( .A(n31354), .B(n31353), .Z(n31355) );
  AND U32139 ( .A(n31356), .B(n31355), .Z(n31562) );
  NAND U32140 ( .A(n38385), .B(n31357), .Z(n31359) );
  XOR U32141 ( .A(b[27]), .B(a[200]), .Z(n31506) );
  NAND U32142 ( .A(n38343), .B(n31506), .Z(n31358) );
  AND U32143 ( .A(n31359), .B(n31358), .Z(n31569) );
  NAND U32144 ( .A(n183), .B(n31360), .Z(n31362) );
  XOR U32145 ( .A(b[5]), .B(a[222]), .Z(n31509) );
  NAND U32146 ( .A(n36296), .B(n31509), .Z(n31361) );
  AND U32147 ( .A(n31362), .B(n31361), .Z(n31567) );
  NAND U32148 ( .A(n190), .B(n31363), .Z(n31365) );
  XOR U32149 ( .A(b[19]), .B(a[208]), .Z(n31512) );
  NAND U32150 ( .A(n37821), .B(n31512), .Z(n31364) );
  NAND U32151 ( .A(n31365), .B(n31364), .Z(n31566) );
  XNOR U32152 ( .A(n31567), .B(n31566), .Z(n31568) );
  XNOR U32153 ( .A(n31569), .B(n31568), .Z(n31560) );
  NAND U32154 ( .A(n38470), .B(n31366), .Z(n31368) );
  XOR U32155 ( .A(b[31]), .B(a[196]), .Z(n31515) );
  NAND U32156 ( .A(n38453), .B(n31515), .Z(n31367) );
  AND U32157 ( .A(n31368), .B(n31367), .Z(n31527) );
  NAND U32158 ( .A(n181), .B(n31369), .Z(n31371) );
  XOR U32159 ( .A(b[3]), .B(a[224]), .Z(n31518) );
  NAND U32160 ( .A(n182), .B(n31518), .Z(n31370) );
  AND U32161 ( .A(n31371), .B(n31370), .Z(n31525) );
  NAND U32162 ( .A(n189), .B(n31372), .Z(n31374) );
  XOR U32163 ( .A(b[17]), .B(a[210]), .Z(n31521) );
  NAND U32164 ( .A(n37652), .B(n31521), .Z(n31373) );
  NAND U32165 ( .A(n31374), .B(n31373), .Z(n31524) );
  XNOR U32166 ( .A(n31525), .B(n31524), .Z(n31526) );
  XOR U32167 ( .A(n31527), .B(n31526), .Z(n31561) );
  XOR U32168 ( .A(n31560), .B(n31561), .Z(n31563) );
  XOR U32169 ( .A(n31562), .B(n31563), .Z(n31495) );
  NANDN U32170 ( .A(n31376), .B(n31375), .Z(n31380) );
  NANDN U32171 ( .A(n31378), .B(n31377), .Z(n31379) );
  AND U32172 ( .A(n31380), .B(n31379), .Z(n31548) );
  NANDN U32173 ( .A(n31382), .B(n31381), .Z(n31386) );
  NANDN U32174 ( .A(n31384), .B(n31383), .Z(n31385) );
  NAND U32175 ( .A(n31386), .B(n31385), .Z(n31549) );
  XNOR U32176 ( .A(n31548), .B(n31549), .Z(n31550) );
  NANDN U32177 ( .A(n31388), .B(n31387), .Z(n31392) );
  NANDN U32178 ( .A(n31390), .B(n31389), .Z(n31391) );
  NAND U32179 ( .A(n31392), .B(n31391), .Z(n31551) );
  XNOR U32180 ( .A(n31550), .B(n31551), .Z(n31494) );
  XNOR U32181 ( .A(n31495), .B(n31494), .Z(n31497) );
  NANDN U32182 ( .A(n31394), .B(n31393), .Z(n31398) );
  NANDN U32183 ( .A(n31396), .B(n31395), .Z(n31397) );
  AND U32184 ( .A(n31398), .B(n31397), .Z(n31496) );
  XOR U32185 ( .A(n31497), .B(n31496), .Z(n31611) );
  NANDN U32186 ( .A(n31400), .B(n31399), .Z(n31404) );
  NANDN U32187 ( .A(n31402), .B(n31401), .Z(n31403) );
  AND U32188 ( .A(n31404), .B(n31403), .Z(n31608) );
  NANDN U32189 ( .A(n31406), .B(n31405), .Z(n31410) );
  NANDN U32190 ( .A(n31408), .B(n31407), .Z(n31409) );
  AND U32191 ( .A(n31410), .B(n31409), .Z(n31491) );
  NANDN U32192 ( .A(n31412), .B(n31411), .Z(n31416) );
  OR U32193 ( .A(n31414), .B(n31413), .Z(n31415) );
  AND U32194 ( .A(n31416), .B(n31415), .Z(n31489) );
  NANDN U32195 ( .A(n31418), .B(n31417), .Z(n31422) );
  NANDN U32196 ( .A(n31420), .B(n31419), .Z(n31421) );
  AND U32197 ( .A(n31422), .B(n31421), .Z(n31555) );
  NANDN U32198 ( .A(n31424), .B(n31423), .Z(n31428) );
  NANDN U32199 ( .A(n31426), .B(n31425), .Z(n31427) );
  NAND U32200 ( .A(n31428), .B(n31427), .Z(n31554) );
  XNOR U32201 ( .A(n31555), .B(n31554), .Z(n31556) );
  NAND U32202 ( .A(b[0]), .B(a[226]), .Z(n31429) );
  XNOR U32203 ( .A(b[1]), .B(n31429), .Z(n31431) );
  NANDN U32204 ( .A(b[0]), .B(a[225]), .Z(n31430) );
  NAND U32205 ( .A(n31431), .B(n31430), .Z(n31503) );
  NAND U32206 ( .A(n194), .B(n31432), .Z(n31434) );
  XOR U32207 ( .A(b[29]), .B(a[198]), .Z(n31581) );
  NAND U32208 ( .A(n38456), .B(n31581), .Z(n31433) );
  AND U32209 ( .A(n31434), .B(n31433), .Z(n31501) );
  AND U32210 ( .A(b[31]), .B(a[194]), .Z(n31500) );
  XNOR U32211 ( .A(n31501), .B(n31500), .Z(n31502) );
  XNOR U32212 ( .A(n31503), .B(n31502), .Z(n31542) );
  NAND U32213 ( .A(n38185), .B(n31435), .Z(n31437) );
  XOR U32214 ( .A(b[23]), .B(a[204]), .Z(n31584) );
  NAND U32215 ( .A(n38132), .B(n31584), .Z(n31436) );
  AND U32216 ( .A(n31437), .B(n31436), .Z(n31575) );
  NAND U32217 ( .A(n184), .B(n31438), .Z(n31440) );
  XOR U32218 ( .A(b[7]), .B(a[220]), .Z(n31587) );
  NAND U32219 ( .A(n36592), .B(n31587), .Z(n31439) );
  AND U32220 ( .A(n31440), .B(n31439), .Z(n31573) );
  NAND U32221 ( .A(n38289), .B(n31441), .Z(n31443) );
  XOR U32222 ( .A(b[25]), .B(a[202]), .Z(n31590) );
  NAND U32223 ( .A(n38247), .B(n31590), .Z(n31442) );
  NAND U32224 ( .A(n31443), .B(n31442), .Z(n31572) );
  XNOR U32225 ( .A(n31573), .B(n31572), .Z(n31574) );
  XOR U32226 ( .A(n31575), .B(n31574), .Z(n31543) );
  XNOR U32227 ( .A(n31542), .B(n31543), .Z(n31544) );
  NAND U32228 ( .A(n187), .B(n31444), .Z(n31446) );
  XOR U32229 ( .A(b[13]), .B(a[214]), .Z(n31593) );
  NAND U32230 ( .A(n37295), .B(n31593), .Z(n31445) );
  AND U32231 ( .A(n31446), .B(n31445), .Z(n31537) );
  NAND U32232 ( .A(n186), .B(n31447), .Z(n31449) );
  XOR U32233 ( .A(b[11]), .B(a[216]), .Z(n31596) );
  NAND U32234 ( .A(n37097), .B(n31596), .Z(n31448) );
  NAND U32235 ( .A(n31449), .B(n31448), .Z(n31536) );
  XNOR U32236 ( .A(n31537), .B(n31536), .Z(n31538) );
  NAND U32237 ( .A(n188), .B(n31450), .Z(n31452) );
  XOR U32238 ( .A(b[15]), .B(a[212]), .Z(n31599) );
  NAND U32239 ( .A(n37382), .B(n31599), .Z(n31451) );
  AND U32240 ( .A(n31452), .B(n31451), .Z(n31533) );
  NAND U32241 ( .A(n38064), .B(n31453), .Z(n31455) );
  XOR U32242 ( .A(b[21]), .B(a[206]), .Z(n31602) );
  NAND U32243 ( .A(n37993), .B(n31602), .Z(n31454) );
  AND U32244 ( .A(n31455), .B(n31454), .Z(n31531) );
  NAND U32245 ( .A(n185), .B(n31456), .Z(n31458) );
  XOR U32246 ( .A(b[9]), .B(a[218]), .Z(n31605) );
  NAND U32247 ( .A(n36805), .B(n31605), .Z(n31457) );
  NAND U32248 ( .A(n31458), .B(n31457), .Z(n31530) );
  XNOR U32249 ( .A(n31531), .B(n31530), .Z(n31532) );
  XOR U32250 ( .A(n31533), .B(n31532), .Z(n31539) );
  XOR U32251 ( .A(n31538), .B(n31539), .Z(n31545) );
  XOR U32252 ( .A(n31544), .B(n31545), .Z(n31557) );
  XNOR U32253 ( .A(n31556), .B(n31557), .Z(n31488) );
  XNOR U32254 ( .A(n31489), .B(n31488), .Z(n31490) );
  XOR U32255 ( .A(n31491), .B(n31490), .Z(n31609) );
  XNOR U32256 ( .A(n31608), .B(n31609), .Z(n31610) );
  XNOR U32257 ( .A(n31611), .B(n31610), .Z(n31484) );
  XOR U32258 ( .A(n31485), .B(n31484), .Z(n31477) );
  NANDN U32259 ( .A(n31460), .B(n31459), .Z(n31464) );
  OR U32260 ( .A(n31462), .B(n31461), .Z(n31463) );
  AND U32261 ( .A(n31464), .B(n31463), .Z(n31476) );
  XNOR U32262 ( .A(n31477), .B(n31476), .Z(n31478) );
  XNOR U32263 ( .A(n31479), .B(n31478), .Z(n31470) );
  XNOR U32264 ( .A(n31471), .B(n31470), .Z(n31472) );
  XNOR U32265 ( .A(n31473), .B(n31472), .Z(n31614) );
  XNOR U32266 ( .A(sreg[450]), .B(n31614), .Z(n31616) );
  NANDN U32267 ( .A(sreg[449]), .B(n31465), .Z(n31469) );
  NAND U32268 ( .A(n31467), .B(n31466), .Z(n31468) );
  NAND U32269 ( .A(n31469), .B(n31468), .Z(n31615) );
  XNOR U32270 ( .A(n31616), .B(n31615), .Z(c[450]) );
  NANDN U32271 ( .A(n31471), .B(n31470), .Z(n31475) );
  NANDN U32272 ( .A(n31473), .B(n31472), .Z(n31474) );
  AND U32273 ( .A(n31475), .B(n31474), .Z(n31622) );
  NANDN U32274 ( .A(n31477), .B(n31476), .Z(n31481) );
  NANDN U32275 ( .A(n31479), .B(n31478), .Z(n31480) );
  AND U32276 ( .A(n31481), .B(n31480), .Z(n31620) );
  NANDN U32277 ( .A(n31483), .B(n31482), .Z(n31487) );
  NAND U32278 ( .A(n31485), .B(n31484), .Z(n31486) );
  AND U32279 ( .A(n31487), .B(n31486), .Z(n31627) );
  NANDN U32280 ( .A(n31489), .B(n31488), .Z(n31493) );
  NANDN U32281 ( .A(n31491), .B(n31490), .Z(n31492) );
  AND U32282 ( .A(n31493), .B(n31492), .Z(n31632) );
  NANDN U32283 ( .A(n31495), .B(n31494), .Z(n31499) );
  NAND U32284 ( .A(n31497), .B(n31496), .Z(n31498) );
  AND U32285 ( .A(n31499), .B(n31498), .Z(n31631) );
  XNOR U32286 ( .A(n31632), .B(n31631), .Z(n31634) );
  NANDN U32287 ( .A(n31501), .B(n31500), .Z(n31505) );
  NANDN U32288 ( .A(n31503), .B(n31502), .Z(n31504) );
  AND U32289 ( .A(n31505), .B(n31504), .Z(n31711) );
  NAND U32290 ( .A(n38385), .B(n31506), .Z(n31508) );
  XOR U32291 ( .A(b[27]), .B(a[201]), .Z(n31655) );
  NAND U32292 ( .A(n38343), .B(n31655), .Z(n31507) );
  AND U32293 ( .A(n31508), .B(n31507), .Z(n31718) );
  NAND U32294 ( .A(n183), .B(n31509), .Z(n31511) );
  XOR U32295 ( .A(b[5]), .B(a[223]), .Z(n31658) );
  NAND U32296 ( .A(n36296), .B(n31658), .Z(n31510) );
  AND U32297 ( .A(n31511), .B(n31510), .Z(n31716) );
  NAND U32298 ( .A(n190), .B(n31512), .Z(n31514) );
  XOR U32299 ( .A(b[19]), .B(a[209]), .Z(n31661) );
  NAND U32300 ( .A(n37821), .B(n31661), .Z(n31513) );
  NAND U32301 ( .A(n31514), .B(n31513), .Z(n31715) );
  XNOR U32302 ( .A(n31716), .B(n31715), .Z(n31717) );
  XNOR U32303 ( .A(n31718), .B(n31717), .Z(n31709) );
  NAND U32304 ( .A(n38470), .B(n31515), .Z(n31517) );
  XOR U32305 ( .A(b[31]), .B(a[197]), .Z(n31664) );
  NAND U32306 ( .A(n38453), .B(n31664), .Z(n31516) );
  AND U32307 ( .A(n31517), .B(n31516), .Z(n31676) );
  NAND U32308 ( .A(n181), .B(n31518), .Z(n31520) );
  XOR U32309 ( .A(b[3]), .B(a[225]), .Z(n31667) );
  NAND U32310 ( .A(n182), .B(n31667), .Z(n31519) );
  AND U32311 ( .A(n31520), .B(n31519), .Z(n31674) );
  NAND U32312 ( .A(n189), .B(n31521), .Z(n31523) );
  XOR U32313 ( .A(b[17]), .B(a[211]), .Z(n31670) );
  NAND U32314 ( .A(n37652), .B(n31670), .Z(n31522) );
  NAND U32315 ( .A(n31523), .B(n31522), .Z(n31673) );
  XNOR U32316 ( .A(n31674), .B(n31673), .Z(n31675) );
  XOR U32317 ( .A(n31676), .B(n31675), .Z(n31710) );
  XOR U32318 ( .A(n31709), .B(n31710), .Z(n31712) );
  XOR U32319 ( .A(n31711), .B(n31712), .Z(n31644) );
  NANDN U32320 ( .A(n31525), .B(n31524), .Z(n31529) );
  NANDN U32321 ( .A(n31527), .B(n31526), .Z(n31528) );
  AND U32322 ( .A(n31529), .B(n31528), .Z(n31697) );
  NANDN U32323 ( .A(n31531), .B(n31530), .Z(n31535) );
  NANDN U32324 ( .A(n31533), .B(n31532), .Z(n31534) );
  NAND U32325 ( .A(n31535), .B(n31534), .Z(n31698) );
  XNOR U32326 ( .A(n31697), .B(n31698), .Z(n31699) );
  NANDN U32327 ( .A(n31537), .B(n31536), .Z(n31541) );
  NANDN U32328 ( .A(n31539), .B(n31538), .Z(n31540) );
  NAND U32329 ( .A(n31541), .B(n31540), .Z(n31700) );
  XNOR U32330 ( .A(n31699), .B(n31700), .Z(n31643) );
  XNOR U32331 ( .A(n31644), .B(n31643), .Z(n31646) );
  NANDN U32332 ( .A(n31543), .B(n31542), .Z(n31547) );
  NANDN U32333 ( .A(n31545), .B(n31544), .Z(n31546) );
  AND U32334 ( .A(n31547), .B(n31546), .Z(n31645) );
  XOR U32335 ( .A(n31646), .B(n31645), .Z(n31760) );
  NANDN U32336 ( .A(n31549), .B(n31548), .Z(n31553) );
  NANDN U32337 ( .A(n31551), .B(n31550), .Z(n31552) );
  AND U32338 ( .A(n31553), .B(n31552), .Z(n31757) );
  NANDN U32339 ( .A(n31555), .B(n31554), .Z(n31559) );
  NANDN U32340 ( .A(n31557), .B(n31556), .Z(n31558) );
  AND U32341 ( .A(n31559), .B(n31558), .Z(n31640) );
  NANDN U32342 ( .A(n31561), .B(n31560), .Z(n31565) );
  OR U32343 ( .A(n31563), .B(n31562), .Z(n31564) );
  AND U32344 ( .A(n31565), .B(n31564), .Z(n31638) );
  NANDN U32345 ( .A(n31567), .B(n31566), .Z(n31571) );
  NANDN U32346 ( .A(n31569), .B(n31568), .Z(n31570) );
  AND U32347 ( .A(n31571), .B(n31570), .Z(n31704) );
  NANDN U32348 ( .A(n31573), .B(n31572), .Z(n31577) );
  NANDN U32349 ( .A(n31575), .B(n31574), .Z(n31576) );
  NAND U32350 ( .A(n31577), .B(n31576), .Z(n31703) );
  XNOR U32351 ( .A(n31704), .B(n31703), .Z(n31705) );
  NAND U32352 ( .A(b[0]), .B(a[227]), .Z(n31578) );
  XNOR U32353 ( .A(b[1]), .B(n31578), .Z(n31580) );
  NANDN U32354 ( .A(b[0]), .B(a[226]), .Z(n31579) );
  NAND U32355 ( .A(n31580), .B(n31579), .Z(n31652) );
  NAND U32356 ( .A(n194), .B(n31581), .Z(n31583) );
  XOR U32357 ( .A(b[29]), .B(a[199]), .Z(n31727) );
  NAND U32358 ( .A(n38456), .B(n31727), .Z(n31582) );
  AND U32359 ( .A(n31583), .B(n31582), .Z(n31650) );
  AND U32360 ( .A(b[31]), .B(a[195]), .Z(n31649) );
  XNOR U32361 ( .A(n31650), .B(n31649), .Z(n31651) );
  XNOR U32362 ( .A(n31652), .B(n31651), .Z(n31691) );
  NAND U32363 ( .A(n38185), .B(n31584), .Z(n31586) );
  XOR U32364 ( .A(b[23]), .B(a[205]), .Z(n31733) );
  NAND U32365 ( .A(n38132), .B(n31733), .Z(n31585) );
  AND U32366 ( .A(n31586), .B(n31585), .Z(n31724) );
  NAND U32367 ( .A(n184), .B(n31587), .Z(n31589) );
  XOR U32368 ( .A(b[7]), .B(a[221]), .Z(n31736) );
  NAND U32369 ( .A(n36592), .B(n31736), .Z(n31588) );
  AND U32370 ( .A(n31589), .B(n31588), .Z(n31722) );
  NAND U32371 ( .A(n38289), .B(n31590), .Z(n31592) );
  XOR U32372 ( .A(b[25]), .B(a[203]), .Z(n31739) );
  NAND U32373 ( .A(n38247), .B(n31739), .Z(n31591) );
  NAND U32374 ( .A(n31592), .B(n31591), .Z(n31721) );
  XNOR U32375 ( .A(n31722), .B(n31721), .Z(n31723) );
  XOR U32376 ( .A(n31724), .B(n31723), .Z(n31692) );
  XNOR U32377 ( .A(n31691), .B(n31692), .Z(n31693) );
  NAND U32378 ( .A(n187), .B(n31593), .Z(n31595) );
  XOR U32379 ( .A(b[13]), .B(a[215]), .Z(n31742) );
  NAND U32380 ( .A(n37295), .B(n31742), .Z(n31594) );
  AND U32381 ( .A(n31595), .B(n31594), .Z(n31686) );
  NAND U32382 ( .A(n186), .B(n31596), .Z(n31598) );
  XOR U32383 ( .A(b[11]), .B(a[217]), .Z(n31745) );
  NAND U32384 ( .A(n37097), .B(n31745), .Z(n31597) );
  NAND U32385 ( .A(n31598), .B(n31597), .Z(n31685) );
  XNOR U32386 ( .A(n31686), .B(n31685), .Z(n31687) );
  NAND U32387 ( .A(n188), .B(n31599), .Z(n31601) );
  XOR U32388 ( .A(b[15]), .B(a[213]), .Z(n31748) );
  NAND U32389 ( .A(n37382), .B(n31748), .Z(n31600) );
  AND U32390 ( .A(n31601), .B(n31600), .Z(n31682) );
  NAND U32391 ( .A(n38064), .B(n31602), .Z(n31604) );
  XOR U32392 ( .A(b[21]), .B(a[207]), .Z(n31751) );
  NAND U32393 ( .A(n37993), .B(n31751), .Z(n31603) );
  AND U32394 ( .A(n31604), .B(n31603), .Z(n31680) );
  NAND U32395 ( .A(n185), .B(n31605), .Z(n31607) );
  XOR U32396 ( .A(b[9]), .B(a[219]), .Z(n31754) );
  NAND U32397 ( .A(n36805), .B(n31754), .Z(n31606) );
  NAND U32398 ( .A(n31607), .B(n31606), .Z(n31679) );
  XNOR U32399 ( .A(n31680), .B(n31679), .Z(n31681) );
  XOR U32400 ( .A(n31682), .B(n31681), .Z(n31688) );
  XOR U32401 ( .A(n31687), .B(n31688), .Z(n31694) );
  XOR U32402 ( .A(n31693), .B(n31694), .Z(n31706) );
  XNOR U32403 ( .A(n31705), .B(n31706), .Z(n31637) );
  XNOR U32404 ( .A(n31638), .B(n31637), .Z(n31639) );
  XOR U32405 ( .A(n31640), .B(n31639), .Z(n31758) );
  XNOR U32406 ( .A(n31757), .B(n31758), .Z(n31759) );
  XNOR U32407 ( .A(n31760), .B(n31759), .Z(n31633) );
  XOR U32408 ( .A(n31634), .B(n31633), .Z(n31626) );
  NANDN U32409 ( .A(n31609), .B(n31608), .Z(n31613) );
  NANDN U32410 ( .A(n31611), .B(n31610), .Z(n31612) );
  AND U32411 ( .A(n31613), .B(n31612), .Z(n31625) );
  XOR U32412 ( .A(n31626), .B(n31625), .Z(n31628) );
  XNOR U32413 ( .A(n31627), .B(n31628), .Z(n31619) );
  XNOR U32414 ( .A(n31620), .B(n31619), .Z(n31621) );
  XNOR U32415 ( .A(n31622), .B(n31621), .Z(n31763) );
  XNOR U32416 ( .A(sreg[451]), .B(n31763), .Z(n31765) );
  NANDN U32417 ( .A(sreg[450]), .B(n31614), .Z(n31618) );
  NAND U32418 ( .A(n31616), .B(n31615), .Z(n31617) );
  NAND U32419 ( .A(n31618), .B(n31617), .Z(n31764) );
  XNOR U32420 ( .A(n31765), .B(n31764), .Z(c[451]) );
  NANDN U32421 ( .A(n31620), .B(n31619), .Z(n31624) );
  NANDN U32422 ( .A(n31622), .B(n31621), .Z(n31623) );
  AND U32423 ( .A(n31624), .B(n31623), .Z(n31775) );
  NANDN U32424 ( .A(n31626), .B(n31625), .Z(n31630) );
  NANDN U32425 ( .A(n31628), .B(n31627), .Z(n31629) );
  AND U32426 ( .A(n31630), .B(n31629), .Z(n31774) );
  NANDN U32427 ( .A(n31632), .B(n31631), .Z(n31636) );
  NAND U32428 ( .A(n31634), .B(n31633), .Z(n31635) );
  AND U32429 ( .A(n31636), .B(n31635), .Z(n31781) );
  NANDN U32430 ( .A(n31638), .B(n31637), .Z(n31642) );
  NANDN U32431 ( .A(n31640), .B(n31639), .Z(n31641) );
  AND U32432 ( .A(n31642), .B(n31641), .Z(n31910) );
  NANDN U32433 ( .A(n31644), .B(n31643), .Z(n31648) );
  NAND U32434 ( .A(n31646), .B(n31645), .Z(n31647) );
  AND U32435 ( .A(n31648), .B(n31647), .Z(n31909) );
  XNOR U32436 ( .A(n31910), .B(n31909), .Z(n31912) );
  NANDN U32437 ( .A(n31650), .B(n31649), .Z(n31654) );
  NANDN U32438 ( .A(n31652), .B(n31651), .Z(n31653) );
  AND U32439 ( .A(n31654), .B(n31653), .Z(n31857) );
  NAND U32440 ( .A(n38385), .B(n31655), .Z(n31657) );
  XOR U32441 ( .A(b[27]), .B(a[202]), .Z(n31803) );
  NAND U32442 ( .A(n38343), .B(n31803), .Z(n31656) );
  AND U32443 ( .A(n31657), .B(n31656), .Z(n31864) );
  NAND U32444 ( .A(n183), .B(n31658), .Z(n31660) );
  XOR U32445 ( .A(b[5]), .B(a[224]), .Z(n31806) );
  NAND U32446 ( .A(n36296), .B(n31806), .Z(n31659) );
  AND U32447 ( .A(n31660), .B(n31659), .Z(n31862) );
  NAND U32448 ( .A(n190), .B(n31661), .Z(n31663) );
  XOR U32449 ( .A(b[19]), .B(a[210]), .Z(n31809) );
  NAND U32450 ( .A(n37821), .B(n31809), .Z(n31662) );
  NAND U32451 ( .A(n31663), .B(n31662), .Z(n31861) );
  XNOR U32452 ( .A(n31862), .B(n31861), .Z(n31863) );
  XNOR U32453 ( .A(n31864), .B(n31863), .Z(n31855) );
  NAND U32454 ( .A(n38470), .B(n31664), .Z(n31666) );
  XOR U32455 ( .A(b[31]), .B(a[198]), .Z(n31812) );
  NAND U32456 ( .A(n38453), .B(n31812), .Z(n31665) );
  AND U32457 ( .A(n31666), .B(n31665), .Z(n31824) );
  NAND U32458 ( .A(n181), .B(n31667), .Z(n31669) );
  XOR U32459 ( .A(b[3]), .B(a[226]), .Z(n31815) );
  NAND U32460 ( .A(n182), .B(n31815), .Z(n31668) );
  AND U32461 ( .A(n31669), .B(n31668), .Z(n31822) );
  NAND U32462 ( .A(n189), .B(n31670), .Z(n31672) );
  XOR U32463 ( .A(b[17]), .B(a[212]), .Z(n31818) );
  NAND U32464 ( .A(n37652), .B(n31818), .Z(n31671) );
  NAND U32465 ( .A(n31672), .B(n31671), .Z(n31821) );
  XNOR U32466 ( .A(n31822), .B(n31821), .Z(n31823) );
  XOR U32467 ( .A(n31824), .B(n31823), .Z(n31856) );
  XOR U32468 ( .A(n31855), .B(n31856), .Z(n31858) );
  XOR U32469 ( .A(n31857), .B(n31858), .Z(n31792) );
  NANDN U32470 ( .A(n31674), .B(n31673), .Z(n31678) );
  NANDN U32471 ( .A(n31676), .B(n31675), .Z(n31677) );
  AND U32472 ( .A(n31678), .B(n31677), .Z(n31845) );
  NANDN U32473 ( .A(n31680), .B(n31679), .Z(n31684) );
  NANDN U32474 ( .A(n31682), .B(n31681), .Z(n31683) );
  NAND U32475 ( .A(n31684), .B(n31683), .Z(n31846) );
  XNOR U32476 ( .A(n31845), .B(n31846), .Z(n31847) );
  NANDN U32477 ( .A(n31686), .B(n31685), .Z(n31690) );
  NANDN U32478 ( .A(n31688), .B(n31687), .Z(n31689) );
  NAND U32479 ( .A(n31690), .B(n31689), .Z(n31848) );
  XNOR U32480 ( .A(n31847), .B(n31848), .Z(n31791) );
  XNOR U32481 ( .A(n31792), .B(n31791), .Z(n31794) );
  NANDN U32482 ( .A(n31692), .B(n31691), .Z(n31696) );
  NANDN U32483 ( .A(n31694), .B(n31693), .Z(n31695) );
  AND U32484 ( .A(n31696), .B(n31695), .Z(n31793) );
  XOR U32485 ( .A(n31794), .B(n31793), .Z(n31906) );
  NANDN U32486 ( .A(n31698), .B(n31697), .Z(n31702) );
  NANDN U32487 ( .A(n31700), .B(n31699), .Z(n31701) );
  AND U32488 ( .A(n31702), .B(n31701), .Z(n31903) );
  NANDN U32489 ( .A(n31704), .B(n31703), .Z(n31708) );
  NANDN U32490 ( .A(n31706), .B(n31705), .Z(n31707) );
  AND U32491 ( .A(n31708), .B(n31707), .Z(n31788) );
  NANDN U32492 ( .A(n31710), .B(n31709), .Z(n31714) );
  OR U32493 ( .A(n31712), .B(n31711), .Z(n31713) );
  AND U32494 ( .A(n31714), .B(n31713), .Z(n31786) );
  NANDN U32495 ( .A(n31716), .B(n31715), .Z(n31720) );
  NANDN U32496 ( .A(n31718), .B(n31717), .Z(n31719) );
  AND U32497 ( .A(n31720), .B(n31719), .Z(n31852) );
  NANDN U32498 ( .A(n31722), .B(n31721), .Z(n31726) );
  NANDN U32499 ( .A(n31724), .B(n31723), .Z(n31725) );
  NAND U32500 ( .A(n31726), .B(n31725), .Z(n31851) );
  XNOR U32501 ( .A(n31852), .B(n31851), .Z(n31854) );
  NAND U32502 ( .A(n194), .B(n31727), .Z(n31729) );
  XOR U32503 ( .A(b[29]), .B(a[200]), .Z(n31876) );
  NAND U32504 ( .A(n38456), .B(n31876), .Z(n31728) );
  AND U32505 ( .A(n31729), .B(n31728), .Z(n31798) );
  AND U32506 ( .A(b[31]), .B(a[196]), .Z(n31797) );
  XNOR U32507 ( .A(n31798), .B(n31797), .Z(n31799) );
  NAND U32508 ( .A(b[0]), .B(a[228]), .Z(n31730) );
  XNOR U32509 ( .A(b[1]), .B(n31730), .Z(n31732) );
  NANDN U32510 ( .A(b[0]), .B(a[227]), .Z(n31731) );
  NAND U32511 ( .A(n31732), .B(n31731), .Z(n31800) );
  XNOR U32512 ( .A(n31799), .B(n31800), .Z(n31840) );
  NAND U32513 ( .A(n38185), .B(n31733), .Z(n31735) );
  XOR U32514 ( .A(b[23]), .B(a[206]), .Z(n31879) );
  NAND U32515 ( .A(n38132), .B(n31879), .Z(n31734) );
  AND U32516 ( .A(n31735), .B(n31734), .Z(n31869) );
  NAND U32517 ( .A(n184), .B(n31736), .Z(n31738) );
  XOR U32518 ( .A(b[7]), .B(a[222]), .Z(n31882) );
  NAND U32519 ( .A(n36592), .B(n31882), .Z(n31737) );
  AND U32520 ( .A(n31738), .B(n31737), .Z(n31868) );
  NAND U32521 ( .A(n38289), .B(n31739), .Z(n31741) );
  XOR U32522 ( .A(b[25]), .B(a[204]), .Z(n31885) );
  NAND U32523 ( .A(n38247), .B(n31885), .Z(n31740) );
  NAND U32524 ( .A(n31741), .B(n31740), .Z(n31867) );
  XOR U32525 ( .A(n31868), .B(n31867), .Z(n31870) );
  XOR U32526 ( .A(n31869), .B(n31870), .Z(n31839) );
  XOR U32527 ( .A(n31840), .B(n31839), .Z(n31842) );
  NAND U32528 ( .A(n187), .B(n31742), .Z(n31744) );
  XOR U32529 ( .A(b[13]), .B(a[216]), .Z(n31888) );
  NAND U32530 ( .A(n37295), .B(n31888), .Z(n31743) );
  AND U32531 ( .A(n31744), .B(n31743), .Z(n31834) );
  NAND U32532 ( .A(n186), .B(n31745), .Z(n31747) );
  XOR U32533 ( .A(b[11]), .B(a[218]), .Z(n31891) );
  NAND U32534 ( .A(n37097), .B(n31891), .Z(n31746) );
  NAND U32535 ( .A(n31747), .B(n31746), .Z(n31833) );
  XNOR U32536 ( .A(n31834), .B(n31833), .Z(n31836) );
  NAND U32537 ( .A(n188), .B(n31748), .Z(n31750) );
  XOR U32538 ( .A(b[15]), .B(a[214]), .Z(n31894) );
  NAND U32539 ( .A(n37382), .B(n31894), .Z(n31749) );
  AND U32540 ( .A(n31750), .B(n31749), .Z(n31830) );
  NAND U32541 ( .A(n38064), .B(n31751), .Z(n31753) );
  XOR U32542 ( .A(b[21]), .B(a[208]), .Z(n31897) );
  NAND U32543 ( .A(n37993), .B(n31897), .Z(n31752) );
  AND U32544 ( .A(n31753), .B(n31752), .Z(n31828) );
  NAND U32545 ( .A(n185), .B(n31754), .Z(n31756) );
  XOR U32546 ( .A(b[9]), .B(a[220]), .Z(n31900) );
  NAND U32547 ( .A(n36805), .B(n31900), .Z(n31755) );
  NAND U32548 ( .A(n31756), .B(n31755), .Z(n31827) );
  XNOR U32549 ( .A(n31828), .B(n31827), .Z(n31829) );
  XNOR U32550 ( .A(n31830), .B(n31829), .Z(n31835) );
  XOR U32551 ( .A(n31836), .B(n31835), .Z(n31841) );
  XNOR U32552 ( .A(n31842), .B(n31841), .Z(n31853) );
  XNOR U32553 ( .A(n31854), .B(n31853), .Z(n31785) );
  XNOR U32554 ( .A(n31786), .B(n31785), .Z(n31787) );
  XOR U32555 ( .A(n31788), .B(n31787), .Z(n31904) );
  XNOR U32556 ( .A(n31903), .B(n31904), .Z(n31905) );
  XNOR U32557 ( .A(n31906), .B(n31905), .Z(n31911) );
  XOR U32558 ( .A(n31912), .B(n31911), .Z(n31780) );
  NANDN U32559 ( .A(n31758), .B(n31757), .Z(n31762) );
  NANDN U32560 ( .A(n31760), .B(n31759), .Z(n31761) );
  AND U32561 ( .A(n31762), .B(n31761), .Z(n31779) );
  XOR U32562 ( .A(n31780), .B(n31779), .Z(n31782) );
  XNOR U32563 ( .A(n31781), .B(n31782), .Z(n31773) );
  XOR U32564 ( .A(n31774), .B(n31773), .Z(n31776) );
  XOR U32565 ( .A(n31775), .B(n31776), .Z(n31768) );
  XNOR U32566 ( .A(n31768), .B(sreg[452]), .Z(n31770) );
  NANDN U32567 ( .A(sreg[451]), .B(n31763), .Z(n31767) );
  NAND U32568 ( .A(n31765), .B(n31764), .Z(n31766) );
  AND U32569 ( .A(n31767), .B(n31766), .Z(n31769) );
  XOR U32570 ( .A(n31770), .B(n31769), .Z(c[452]) );
  NANDN U32571 ( .A(n31768), .B(sreg[452]), .Z(n31772) );
  NAND U32572 ( .A(n31770), .B(n31769), .Z(n31771) );
  AND U32573 ( .A(n31772), .B(n31771), .Z(n32061) );
  NANDN U32574 ( .A(n31774), .B(n31773), .Z(n31778) );
  OR U32575 ( .A(n31776), .B(n31775), .Z(n31777) );
  AND U32576 ( .A(n31778), .B(n31777), .Z(n31918) );
  NANDN U32577 ( .A(n31780), .B(n31779), .Z(n31784) );
  NANDN U32578 ( .A(n31782), .B(n31781), .Z(n31783) );
  AND U32579 ( .A(n31784), .B(n31783), .Z(n31916) );
  NANDN U32580 ( .A(n31786), .B(n31785), .Z(n31790) );
  NANDN U32581 ( .A(n31788), .B(n31787), .Z(n31789) );
  AND U32582 ( .A(n31790), .B(n31789), .Z(n32054) );
  NANDN U32583 ( .A(n31792), .B(n31791), .Z(n31796) );
  NAND U32584 ( .A(n31794), .B(n31793), .Z(n31795) );
  AND U32585 ( .A(n31796), .B(n31795), .Z(n32053) );
  XNOR U32586 ( .A(n32054), .B(n32053), .Z(n32056) );
  NANDN U32587 ( .A(n31798), .B(n31797), .Z(n31802) );
  NANDN U32588 ( .A(n31800), .B(n31799), .Z(n31801) );
  AND U32589 ( .A(n31802), .B(n31801), .Z(n31989) );
  NAND U32590 ( .A(n38385), .B(n31803), .Z(n31805) );
  XOR U32591 ( .A(b[27]), .B(a[203]), .Z(n31933) );
  NAND U32592 ( .A(n38343), .B(n31933), .Z(n31804) );
  AND U32593 ( .A(n31805), .B(n31804), .Z(n31996) );
  NAND U32594 ( .A(n183), .B(n31806), .Z(n31808) );
  XOR U32595 ( .A(b[5]), .B(a[225]), .Z(n31936) );
  NAND U32596 ( .A(n36296), .B(n31936), .Z(n31807) );
  AND U32597 ( .A(n31808), .B(n31807), .Z(n31994) );
  NAND U32598 ( .A(n190), .B(n31809), .Z(n31811) );
  XOR U32599 ( .A(b[19]), .B(a[211]), .Z(n31939) );
  NAND U32600 ( .A(n37821), .B(n31939), .Z(n31810) );
  NAND U32601 ( .A(n31811), .B(n31810), .Z(n31993) );
  XNOR U32602 ( .A(n31994), .B(n31993), .Z(n31995) );
  XNOR U32603 ( .A(n31996), .B(n31995), .Z(n31987) );
  NAND U32604 ( .A(n38470), .B(n31812), .Z(n31814) );
  XOR U32605 ( .A(b[31]), .B(a[199]), .Z(n31942) );
  NAND U32606 ( .A(n38453), .B(n31942), .Z(n31813) );
  AND U32607 ( .A(n31814), .B(n31813), .Z(n31954) );
  NAND U32608 ( .A(n181), .B(n31815), .Z(n31817) );
  XOR U32609 ( .A(b[3]), .B(a[227]), .Z(n31945) );
  NAND U32610 ( .A(n182), .B(n31945), .Z(n31816) );
  AND U32611 ( .A(n31817), .B(n31816), .Z(n31952) );
  NAND U32612 ( .A(n189), .B(n31818), .Z(n31820) );
  XOR U32613 ( .A(b[17]), .B(a[213]), .Z(n31948) );
  NAND U32614 ( .A(n37652), .B(n31948), .Z(n31819) );
  NAND U32615 ( .A(n31820), .B(n31819), .Z(n31951) );
  XNOR U32616 ( .A(n31952), .B(n31951), .Z(n31953) );
  XOR U32617 ( .A(n31954), .B(n31953), .Z(n31988) );
  XOR U32618 ( .A(n31987), .B(n31988), .Z(n31990) );
  XOR U32619 ( .A(n31989), .B(n31990), .Z(n32036) );
  NANDN U32620 ( .A(n31822), .B(n31821), .Z(n31826) );
  NANDN U32621 ( .A(n31824), .B(n31823), .Z(n31825) );
  AND U32622 ( .A(n31826), .B(n31825), .Z(n31975) );
  NANDN U32623 ( .A(n31828), .B(n31827), .Z(n31832) );
  NANDN U32624 ( .A(n31830), .B(n31829), .Z(n31831) );
  NAND U32625 ( .A(n31832), .B(n31831), .Z(n31976) );
  XNOR U32626 ( .A(n31975), .B(n31976), .Z(n31977) );
  NANDN U32627 ( .A(n31834), .B(n31833), .Z(n31838) );
  NAND U32628 ( .A(n31836), .B(n31835), .Z(n31837) );
  NAND U32629 ( .A(n31838), .B(n31837), .Z(n31978) );
  XNOR U32630 ( .A(n31977), .B(n31978), .Z(n32035) );
  XNOR U32631 ( .A(n32036), .B(n32035), .Z(n32038) );
  NAND U32632 ( .A(n31840), .B(n31839), .Z(n31844) );
  NAND U32633 ( .A(n31842), .B(n31841), .Z(n31843) );
  AND U32634 ( .A(n31844), .B(n31843), .Z(n32037) );
  XOR U32635 ( .A(n32038), .B(n32037), .Z(n32050) );
  NANDN U32636 ( .A(n31846), .B(n31845), .Z(n31850) );
  NANDN U32637 ( .A(n31848), .B(n31847), .Z(n31849) );
  AND U32638 ( .A(n31850), .B(n31849), .Z(n32047) );
  NANDN U32639 ( .A(n31856), .B(n31855), .Z(n31860) );
  OR U32640 ( .A(n31858), .B(n31857), .Z(n31859) );
  AND U32641 ( .A(n31860), .B(n31859), .Z(n32042) );
  NANDN U32642 ( .A(n31862), .B(n31861), .Z(n31866) );
  NANDN U32643 ( .A(n31864), .B(n31863), .Z(n31865) );
  AND U32644 ( .A(n31866), .B(n31865), .Z(n31982) );
  NANDN U32645 ( .A(n31868), .B(n31867), .Z(n31872) );
  OR U32646 ( .A(n31870), .B(n31869), .Z(n31871) );
  NAND U32647 ( .A(n31872), .B(n31871), .Z(n31981) );
  XNOR U32648 ( .A(n31982), .B(n31981), .Z(n31983) );
  NAND U32649 ( .A(b[0]), .B(a[229]), .Z(n31873) );
  XNOR U32650 ( .A(b[1]), .B(n31873), .Z(n31875) );
  NANDN U32651 ( .A(b[0]), .B(a[228]), .Z(n31874) );
  NAND U32652 ( .A(n31875), .B(n31874), .Z(n31930) );
  NAND U32653 ( .A(n194), .B(n31876), .Z(n31878) );
  XOR U32654 ( .A(b[29]), .B(a[201]), .Z(n32008) );
  NAND U32655 ( .A(n38456), .B(n32008), .Z(n31877) );
  AND U32656 ( .A(n31878), .B(n31877), .Z(n31928) );
  AND U32657 ( .A(b[31]), .B(a[197]), .Z(n31927) );
  XNOR U32658 ( .A(n31928), .B(n31927), .Z(n31929) );
  XNOR U32659 ( .A(n31930), .B(n31929), .Z(n31969) );
  NAND U32660 ( .A(n38185), .B(n31879), .Z(n31881) );
  XOR U32661 ( .A(b[23]), .B(a[207]), .Z(n32011) );
  NAND U32662 ( .A(n38132), .B(n32011), .Z(n31880) );
  AND U32663 ( .A(n31881), .B(n31880), .Z(n32002) );
  NAND U32664 ( .A(n184), .B(n31882), .Z(n31884) );
  XOR U32665 ( .A(b[7]), .B(a[223]), .Z(n32014) );
  NAND U32666 ( .A(n36592), .B(n32014), .Z(n31883) );
  AND U32667 ( .A(n31884), .B(n31883), .Z(n32000) );
  NAND U32668 ( .A(n38289), .B(n31885), .Z(n31887) );
  XOR U32669 ( .A(b[25]), .B(a[205]), .Z(n32017) );
  NAND U32670 ( .A(n38247), .B(n32017), .Z(n31886) );
  NAND U32671 ( .A(n31887), .B(n31886), .Z(n31999) );
  XNOR U32672 ( .A(n32000), .B(n31999), .Z(n32001) );
  XOR U32673 ( .A(n32002), .B(n32001), .Z(n31970) );
  XNOR U32674 ( .A(n31969), .B(n31970), .Z(n31971) );
  NAND U32675 ( .A(n187), .B(n31888), .Z(n31890) );
  XOR U32676 ( .A(b[13]), .B(a[217]), .Z(n32020) );
  NAND U32677 ( .A(n37295), .B(n32020), .Z(n31889) );
  AND U32678 ( .A(n31890), .B(n31889), .Z(n31964) );
  NAND U32679 ( .A(n186), .B(n31891), .Z(n31893) );
  XOR U32680 ( .A(b[11]), .B(a[219]), .Z(n32023) );
  NAND U32681 ( .A(n37097), .B(n32023), .Z(n31892) );
  NAND U32682 ( .A(n31893), .B(n31892), .Z(n31963) );
  XNOR U32683 ( .A(n31964), .B(n31963), .Z(n31965) );
  NAND U32684 ( .A(n188), .B(n31894), .Z(n31896) );
  XOR U32685 ( .A(b[15]), .B(a[215]), .Z(n32026) );
  NAND U32686 ( .A(n37382), .B(n32026), .Z(n31895) );
  AND U32687 ( .A(n31896), .B(n31895), .Z(n31960) );
  NAND U32688 ( .A(n38064), .B(n31897), .Z(n31899) );
  XOR U32689 ( .A(b[21]), .B(a[209]), .Z(n32029) );
  NAND U32690 ( .A(n37993), .B(n32029), .Z(n31898) );
  AND U32691 ( .A(n31899), .B(n31898), .Z(n31958) );
  NAND U32692 ( .A(n185), .B(n31900), .Z(n31902) );
  XOR U32693 ( .A(b[9]), .B(a[221]), .Z(n32032) );
  NAND U32694 ( .A(n36805), .B(n32032), .Z(n31901) );
  NAND U32695 ( .A(n31902), .B(n31901), .Z(n31957) );
  XNOR U32696 ( .A(n31958), .B(n31957), .Z(n31959) );
  XOR U32697 ( .A(n31960), .B(n31959), .Z(n31966) );
  XOR U32698 ( .A(n31965), .B(n31966), .Z(n31972) );
  XOR U32699 ( .A(n31971), .B(n31972), .Z(n31984) );
  XNOR U32700 ( .A(n31983), .B(n31984), .Z(n32041) );
  XNOR U32701 ( .A(n32042), .B(n32041), .Z(n32043) );
  XOR U32702 ( .A(n32044), .B(n32043), .Z(n32048) );
  XNOR U32703 ( .A(n32047), .B(n32048), .Z(n32049) );
  XNOR U32704 ( .A(n32050), .B(n32049), .Z(n32055) );
  XOR U32705 ( .A(n32056), .B(n32055), .Z(n31922) );
  NANDN U32706 ( .A(n31904), .B(n31903), .Z(n31908) );
  NANDN U32707 ( .A(n31906), .B(n31905), .Z(n31907) );
  AND U32708 ( .A(n31908), .B(n31907), .Z(n31921) );
  XNOR U32709 ( .A(n31922), .B(n31921), .Z(n31923) );
  NANDN U32710 ( .A(n31910), .B(n31909), .Z(n31914) );
  NAND U32711 ( .A(n31912), .B(n31911), .Z(n31913) );
  NAND U32712 ( .A(n31914), .B(n31913), .Z(n31924) );
  XNOR U32713 ( .A(n31923), .B(n31924), .Z(n31915) );
  XNOR U32714 ( .A(n31916), .B(n31915), .Z(n31917) );
  XNOR U32715 ( .A(n31918), .B(n31917), .Z(n32059) );
  XNOR U32716 ( .A(sreg[453]), .B(n32059), .Z(n32060) );
  XNOR U32717 ( .A(n32061), .B(n32060), .Z(c[453]) );
  NANDN U32718 ( .A(n31916), .B(n31915), .Z(n31920) );
  NANDN U32719 ( .A(n31918), .B(n31917), .Z(n31919) );
  AND U32720 ( .A(n31920), .B(n31919), .Z(n32067) );
  NANDN U32721 ( .A(n31922), .B(n31921), .Z(n31926) );
  NANDN U32722 ( .A(n31924), .B(n31923), .Z(n31925) );
  AND U32723 ( .A(n31926), .B(n31925), .Z(n32065) );
  NANDN U32724 ( .A(n31928), .B(n31927), .Z(n31932) );
  NANDN U32725 ( .A(n31930), .B(n31929), .Z(n31931) );
  AND U32726 ( .A(n31932), .B(n31931), .Z(n32156) );
  NAND U32727 ( .A(n38385), .B(n31933), .Z(n31935) );
  XOR U32728 ( .A(b[27]), .B(a[204]), .Z(n32100) );
  NAND U32729 ( .A(n38343), .B(n32100), .Z(n31934) );
  AND U32730 ( .A(n31935), .B(n31934), .Z(n32163) );
  NAND U32731 ( .A(n183), .B(n31936), .Z(n31938) );
  XOR U32732 ( .A(b[5]), .B(a[226]), .Z(n32103) );
  NAND U32733 ( .A(n36296), .B(n32103), .Z(n31937) );
  AND U32734 ( .A(n31938), .B(n31937), .Z(n32161) );
  NAND U32735 ( .A(n190), .B(n31939), .Z(n31941) );
  XOR U32736 ( .A(b[19]), .B(a[212]), .Z(n32106) );
  NAND U32737 ( .A(n37821), .B(n32106), .Z(n31940) );
  NAND U32738 ( .A(n31941), .B(n31940), .Z(n32160) );
  XNOR U32739 ( .A(n32161), .B(n32160), .Z(n32162) );
  XNOR U32740 ( .A(n32163), .B(n32162), .Z(n32154) );
  NAND U32741 ( .A(n38470), .B(n31942), .Z(n31944) );
  XOR U32742 ( .A(b[31]), .B(a[200]), .Z(n32109) );
  NAND U32743 ( .A(n38453), .B(n32109), .Z(n31943) );
  AND U32744 ( .A(n31944), .B(n31943), .Z(n32121) );
  NAND U32745 ( .A(n181), .B(n31945), .Z(n31947) );
  XOR U32746 ( .A(b[3]), .B(a[228]), .Z(n32112) );
  NAND U32747 ( .A(n182), .B(n32112), .Z(n31946) );
  AND U32748 ( .A(n31947), .B(n31946), .Z(n32119) );
  NAND U32749 ( .A(n189), .B(n31948), .Z(n31950) );
  XOR U32750 ( .A(b[17]), .B(a[214]), .Z(n32115) );
  NAND U32751 ( .A(n37652), .B(n32115), .Z(n31949) );
  NAND U32752 ( .A(n31950), .B(n31949), .Z(n32118) );
  XNOR U32753 ( .A(n32119), .B(n32118), .Z(n32120) );
  XOR U32754 ( .A(n32121), .B(n32120), .Z(n32155) );
  XOR U32755 ( .A(n32154), .B(n32155), .Z(n32157) );
  XOR U32756 ( .A(n32156), .B(n32157), .Z(n32089) );
  NANDN U32757 ( .A(n31952), .B(n31951), .Z(n31956) );
  NANDN U32758 ( .A(n31954), .B(n31953), .Z(n31955) );
  AND U32759 ( .A(n31956), .B(n31955), .Z(n32142) );
  NANDN U32760 ( .A(n31958), .B(n31957), .Z(n31962) );
  NANDN U32761 ( .A(n31960), .B(n31959), .Z(n31961) );
  NAND U32762 ( .A(n31962), .B(n31961), .Z(n32143) );
  XNOR U32763 ( .A(n32142), .B(n32143), .Z(n32144) );
  NANDN U32764 ( .A(n31964), .B(n31963), .Z(n31968) );
  NANDN U32765 ( .A(n31966), .B(n31965), .Z(n31967) );
  NAND U32766 ( .A(n31968), .B(n31967), .Z(n32145) );
  XNOR U32767 ( .A(n32144), .B(n32145), .Z(n32088) );
  XNOR U32768 ( .A(n32089), .B(n32088), .Z(n32091) );
  NANDN U32769 ( .A(n31970), .B(n31969), .Z(n31974) );
  NANDN U32770 ( .A(n31972), .B(n31971), .Z(n31973) );
  AND U32771 ( .A(n31974), .B(n31973), .Z(n32090) );
  XOR U32772 ( .A(n32091), .B(n32090), .Z(n32204) );
  NANDN U32773 ( .A(n31976), .B(n31975), .Z(n31980) );
  NANDN U32774 ( .A(n31978), .B(n31977), .Z(n31979) );
  AND U32775 ( .A(n31980), .B(n31979), .Z(n32202) );
  NANDN U32776 ( .A(n31982), .B(n31981), .Z(n31986) );
  NANDN U32777 ( .A(n31984), .B(n31983), .Z(n31985) );
  AND U32778 ( .A(n31986), .B(n31985), .Z(n32085) );
  NANDN U32779 ( .A(n31988), .B(n31987), .Z(n31992) );
  OR U32780 ( .A(n31990), .B(n31989), .Z(n31991) );
  AND U32781 ( .A(n31992), .B(n31991), .Z(n32083) );
  NANDN U32782 ( .A(n31994), .B(n31993), .Z(n31998) );
  NANDN U32783 ( .A(n31996), .B(n31995), .Z(n31997) );
  AND U32784 ( .A(n31998), .B(n31997), .Z(n32149) );
  NANDN U32785 ( .A(n32000), .B(n31999), .Z(n32004) );
  NANDN U32786 ( .A(n32002), .B(n32001), .Z(n32003) );
  NAND U32787 ( .A(n32004), .B(n32003), .Z(n32148) );
  XNOR U32788 ( .A(n32149), .B(n32148), .Z(n32150) );
  NAND U32789 ( .A(b[0]), .B(a[230]), .Z(n32005) );
  XNOR U32790 ( .A(b[1]), .B(n32005), .Z(n32007) );
  NANDN U32791 ( .A(b[0]), .B(a[229]), .Z(n32006) );
  NAND U32792 ( .A(n32007), .B(n32006), .Z(n32097) );
  NAND U32793 ( .A(n194), .B(n32008), .Z(n32010) );
  XOR U32794 ( .A(b[29]), .B(a[202]), .Z(n32175) );
  NAND U32795 ( .A(n38456), .B(n32175), .Z(n32009) );
  AND U32796 ( .A(n32010), .B(n32009), .Z(n32095) );
  AND U32797 ( .A(b[31]), .B(a[198]), .Z(n32094) );
  XNOR U32798 ( .A(n32095), .B(n32094), .Z(n32096) );
  XNOR U32799 ( .A(n32097), .B(n32096), .Z(n32136) );
  NAND U32800 ( .A(n38185), .B(n32011), .Z(n32013) );
  XOR U32801 ( .A(b[23]), .B(a[208]), .Z(n32178) );
  NAND U32802 ( .A(n38132), .B(n32178), .Z(n32012) );
  AND U32803 ( .A(n32013), .B(n32012), .Z(n32169) );
  NAND U32804 ( .A(n184), .B(n32014), .Z(n32016) );
  XOR U32805 ( .A(b[7]), .B(a[224]), .Z(n32181) );
  NAND U32806 ( .A(n36592), .B(n32181), .Z(n32015) );
  AND U32807 ( .A(n32016), .B(n32015), .Z(n32167) );
  NAND U32808 ( .A(n38289), .B(n32017), .Z(n32019) );
  XOR U32809 ( .A(b[25]), .B(a[206]), .Z(n32184) );
  NAND U32810 ( .A(n38247), .B(n32184), .Z(n32018) );
  NAND U32811 ( .A(n32019), .B(n32018), .Z(n32166) );
  XNOR U32812 ( .A(n32167), .B(n32166), .Z(n32168) );
  XOR U32813 ( .A(n32169), .B(n32168), .Z(n32137) );
  XNOR U32814 ( .A(n32136), .B(n32137), .Z(n32138) );
  NAND U32815 ( .A(n187), .B(n32020), .Z(n32022) );
  XOR U32816 ( .A(b[13]), .B(a[218]), .Z(n32187) );
  NAND U32817 ( .A(n37295), .B(n32187), .Z(n32021) );
  AND U32818 ( .A(n32022), .B(n32021), .Z(n32131) );
  NAND U32819 ( .A(n186), .B(n32023), .Z(n32025) );
  XOR U32820 ( .A(b[11]), .B(a[220]), .Z(n32190) );
  NAND U32821 ( .A(n37097), .B(n32190), .Z(n32024) );
  NAND U32822 ( .A(n32025), .B(n32024), .Z(n32130) );
  XNOR U32823 ( .A(n32131), .B(n32130), .Z(n32132) );
  NAND U32824 ( .A(n188), .B(n32026), .Z(n32028) );
  XOR U32825 ( .A(b[15]), .B(a[216]), .Z(n32193) );
  NAND U32826 ( .A(n37382), .B(n32193), .Z(n32027) );
  AND U32827 ( .A(n32028), .B(n32027), .Z(n32127) );
  NAND U32828 ( .A(n38064), .B(n32029), .Z(n32031) );
  XOR U32829 ( .A(b[21]), .B(a[210]), .Z(n32196) );
  NAND U32830 ( .A(n37993), .B(n32196), .Z(n32030) );
  AND U32831 ( .A(n32031), .B(n32030), .Z(n32125) );
  NAND U32832 ( .A(n185), .B(n32032), .Z(n32034) );
  XOR U32833 ( .A(b[9]), .B(a[222]), .Z(n32199) );
  NAND U32834 ( .A(n36805), .B(n32199), .Z(n32033) );
  NAND U32835 ( .A(n32034), .B(n32033), .Z(n32124) );
  XNOR U32836 ( .A(n32125), .B(n32124), .Z(n32126) );
  XOR U32837 ( .A(n32127), .B(n32126), .Z(n32133) );
  XOR U32838 ( .A(n32132), .B(n32133), .Z(n32139) );
  XOR U32839 ( .A(n32138), .B(n32139), .Z(n32151) );
  XNOR U32840 ( .A(n32150), .B(n32151), .Z(n32082) );
  XNOR U32841 ( .A(n32083), .B(n32082), .Z(n32084) );
  XOR U32842 ( .A(n32085), .B(n32084), .Z(n32203) );
  XOR U32843 ( .A(n32202), .B(n32203), .Z(n32205) );
  XOR U32844 ( .A(n32204), .B(n32205), .Z(n32079) );
  NANDN U32845 ( .A(n32036), .B(n32035), .Z(n32040) );
  NAND U32846 ( .A(n32038), .B(n32037), .Z(n32039) );
  AND U32847 ( .A(n32040), .B(n32039), .Z(n32077) );
  NANDN U32848 ( .A(n32042), .B(n32041), .Z(n32046) );
  NANDN U32849 ( .A(n32044), .B(n32043), .Z(n32045) );
  AND U32850 ( .A(n32046), .B(n32045), .Z(n32076) );
  XNOR U32851 ( .A(n32077), .B(n32076), .Z(n32078) );
  XNOR U32852 ( .A(n32079), .B(n32078), .Z(n32070) );
  NANDN U32853 ( .A(n32048), .B(n32047), .Z(n32052) );
  NANDN U32854 ( .A(n32050), .B(n32049), .Z(n32051) );
  NAND U32855 ( .A(n32052), .B(n32051), .Z(n32071) );
  XNOR U32856 ( .A(n32070), .B(n32071), .Z(n32072) );
  NANDN U32857 ( .A(n32054), .B(n32053), .Z(n32058) );
  NAND U32858 ( .A(n32056), .B(n32055), .Z(n32057) );
  NAND U32859 ( .A(n32058), .B(n32057), .Z(n32073) );
  XNOR U32860 ( .A(n32072), .B(n32073), .Z(n32064) );
  XNOR U32861 ( .A(n32065), .B(n32064), .Z(n32066) );
  XNOR U32862 ( .A(n32067), .B(n32066), .Z(n32208) );
  XNOR U32863 ( .A(sreg[454]), .B(n32208), .Z(n32210) );
  NANDN U32864 ( .A(sreg[453]), .B(n32059), .Z(n32063) );
  NAND U32865 ( .A(n32061), .B(n32060), .Z(n32062) );
  NAND U32866 ( .A(n32063), .B(n32062), .Z(n32209) );
  XNOR U32867 ( .A(n32210), .B(n32209), .Z(c[454]) );
  NANDN U32868 ( .A(n32065), .B(n32064), .Z(n32069) );
  NANDN U32869 ( .A(n32067), .B(n32066), .Z(n32068) );
  AND U32870 ( .A(n32069), .B(n32068), .Z(n32216) );
  NANDN U32871 ( .A(n32071), .B(n32070), .Z(n32075) );
  NANDN U32872 ( .A(n32073), .B(n32072), .Z(n32074) );
  AND U32873 ( .A(n32075), .B(n32074), .Z(n32214) );
  NANDN U32874 ( .A(n32077), .B(n32076), .Z(n32081) );
  NANDN U32875 ( .A(n32079), .B(n32078), .Z(n32080) );
  AND U32876 ( .A(n32081), .B(n32080), .Z(n32222) );
  NANDN U32877 ( .A(n32083), .B(n32082), .Z(n32087) );
  NANDN U32878 ( .A(n32085), .B(n32084), .Z(n32086) );
  AND U32879 ( .A(n32087), .B(n32086), .Z(n32226) );
  NANDN U32880 ( .A(n32089), .B(n32088), .Z(n32093) );
  NAND U32881 ( .A(n32091), .B(n32090), .Z(n32092) );
  AND U32882 ( .A(n32093), .B(n32092), .Z(n32225) );
  XNOR U32883 ( .A(n32226), .B(n32225), .Z(n32228) );
  NANDN U32884 ( .A(n32095), .B(n32094), .Z(n32099) );
  NANDN U32885 ( .A(n32097), .B(n32096), .Z(n32098) );
  AND U32886 ( .A(n32099), .B(n32098), .Z(n32305) );
  NAND U32887 ( .A(n38385), .B(n32100), .Z(n32102) );
  XOR U32888 ( .A(b[27]), .B(a[205]), .Z(n32249) );
  NAND U32889 ( .A(n38343), .B(n32249), .Z(n32101) );
  AND U32890 ( .A(n32102), .B(n32101), .Z(n32312) );
  NAND U32891 ( .A(n183), .B(n32103), .Z(n32105) );
  XOR U32892 ( .A(b[5]), .B(a[227]), .Z(n32252) );
  NAND U32893 ( .A(n36296), .B(n32252), .Z(n32104) );
  AND U32894 ( .A(n32105), .B(n32104), .Z(n32310) );
  NAND U32895 ( .A(n190), .B(n32106), .Z(n32108) );
  XOR U32896 ( .A(b[19]), .B(a[213]), .Z(n32255) );
  NAND U32897 ( .A(n37821), .B(n32255), .Z(n32107) );
  NAND U32898 ( .A(n32108), .B(n32107), .Z(n32309) );
  XNOR U32899 ( .A(n32310), .B(n32309), .Z(n32311) );
  XNOR U32900 ( .A(n32312), .B(n32311), .Z(n32303) );
  NAND U32901 ( .A(n38470), .B(n32109), .Z(n32111) );
  XOR U32902 ( .A(b[31]), .B(a[201]), .Z(n32258) );
  NAND U32903 ( .A(n38453), .B(n32258), .Z(n32110) );
  AND U32904 ( .A(n32111), .B(n32110), .Z(n32270) );
  NAND U32905 ( .A(n181), .B(n32112), .Z(n32114) );
  XOR U32906 ( .A(b[3]), .B(a[229]), .Z(n32261) );
  NAND U32907 ( .A(n182), .B(n32261), .Z(n32113) );
  AND U32908 ( .A(n32114), .B(n32113), .Z(n32268) );
  NAND U32909 ( .A(n189), .B(n32115), .Z(n32117) );
  XOR U32910 ( .A(b[17]), .B(a[215]), .Z(n32264) );
  NAND U32911 ( .A(n37652), .B(n32264), .Z(n32116) );
  NAND U32912 ( .A(n32117), .B(n32116), .Z(n32267) );
  XNOR U32913 ( .A(n32268), .B(n32267), .Z(n32269) );
  XOR U32914 ( .A(n32270), .B(n32269), .Z(n32304) );
  XOR U32915 ( .A(n32303), .B(n32304), .Z(n32306) );
  XOR U32916 ( .A(n32305), .B(n32306), .Z(n32238) );
  NANDN U32917 ( .A(n32119), .B(n32118), .Z(n32123) );
  NANDN U32918 ( .A(n32121), .B(n32120), .Z(n32122) );
  AND U32919 ( .A(n32123), .B(n32122), .Z(n32291) );
  NANDN U32920 ( .A(n32125), .B(n32124), .Z(n32129) );
  NANDN U32921 ( .A(n32127), .B(n32126), .Z(n32128) );
  NAND U32922 ( .A(n32129), .B(n32128), .Z(n32292) );
  XNOR U32923 ( .A(n32291), .B(n32292), .Z(n32293) );
  NANDN U32924 ( .A(n32131), .B(n32130), .Z(n32135) );
  NANDN U32925 ( .A(n32133), .B(n32132), .Z(n32134) );
  NAND U32926 ( .A(n32135), .B(n32134), .Z(n32294) );
  XNOR U32927 ( .A(n32293), .B(n32294), .Z(n32237) );
  XNOR U32928 ( .A(n32238), .B(n32237), .Z(n32240) );
  NANDN U32929 ( .A(n32137), .B(n32136), .Z(n32141) );
  NANDN U32930 ( .A(n32139), .B(n32138), .Z(n32140) );
  AND U32931 ( .A(n32141), .B(n32140), .Z(n32239) );
  XOR U32932 ( .A(n32240), .B(n32239), .Z(n32354) );
  NANDN U32933 ( .A(n32143), .B(n32142), .Z(n32147) );
  NANDN U32934 ( .A(n32145), .B(n32144), .Z(n32146) );
  AND U32935 ( .A(n32147), .B(n32146), .Z(n32351) );
  NANDN U32936 ( .A(n32149), .B(n32148), .Z(n32153) );
  NANDN U32937 ( .A(n32151), .B(n32150), .Z(n32152) );
  AND U32938 ( .A(n32153), .B(n32152), .Z(n32234) );
  NANDN U32939 ( .A(n32155), .B(n32154), .Z(n32159) );
  OR U32940 ( .A(n32157), .B(n32156), .Z(n32158) );
  AND U32941 ( .A(n32159), .B(n32158), .Z(n32232) );
  NANDN U32942 ( .A(n32161), .B(n32160), .Z(n32165) );
  NANDN U32943 ( .A(n32163), .B(n32162), .Z(n32164) );
  AND U32944 ( .A(n32165), .B(n32164), .Z(n32298) );
  NANDN U32945 ( .A(n32167), .B(n32166), .Z(n32171) );
  NANDN U32946 ( .A(n32169), .B(n32168), .Z(n32170) );
  NAND U32947 ( .A(n32171), .B(n32170), .Z(n32297) );
  XNOR U32948 ( .A(n32298), .B(n32297), .Z(n32299) );
  NAND U32949 ( .A(b[0]), .B(a[231]), .Z(n32172) );
  XNOR U32950 ( .A(b[1]), .B(n32172), .Z(n32174) );
  NANDN U32951 ( .A(b[0]), .B(a[230]), .Z(n32173) );
  NAND U32952 ( .A(n32174), .B(n32173), .Z(n32246) );
  NAND U32953 ( .A(n194), .B(n32175), .Z(n32177) );
  XOR U32954 ( .A(b[29]), .B(a[203]), .Z(n32324) );
  NAND U32955 ( .A(n38456), .B(n32324), .Z(n32176) );
  AND U32956 ( .A(n32177), .B(n32176), .Z(n32244) );
  AND U32957 ( .A(b[31]), .B(a[199]), .Z(n32243) );
  XNOR U32958 ( .A(n32244), .B(n32243), .Z(n32245) );
  XNOR U32959 ( .A(n32246), .B(n32245), .Z(n32285) );
  NAND U32960 ( .A(n38185), .B(n32178), .Z(n32180) );
  XOR U32961 ( .A(b[23]), .B(a[209]), .Z(n32327) );
  NAND U32962 ( .A(n38132), .B(n32327), .Z(n32179) );
  AND U32963 ( .A(n32180), .B(n32179), .Z(n32318) );
  NAND U32964 ( .A(n184), .B(n32181), .Z(n32183) );
  XOR U32965 ( .A(b[7]), .B(a[225]), .Z(n32330) );
  NAND U32966 ( .A(n36592), .B(n32330), .Z(n32182) );
  AND U32967 ( .A(n32183), .B(n32182), .Z(n32316) );
  NAND U32968 ( .A(n38289), .B(n32184), .Z(n32186) );
  XOR U32969 ( .A(b[25]), .B(a[207]), .Z(n32333) );
  NAND U32970 ( .A(n38247), .B(n32333), .Z(n32185) );
  NAND U32971 ( .A(n32186), .B(n32185), .Z(n32315) );
  XNOR U32972 ( .A(n32316), .B(n32315), .Z(n32317) );
  XOR U32973 ( .A(n32318), .B(n32317), .Z(n32286) );
  XNOR U32974 ( .A(n32285), .B(n32286), .Z(n32287) );
  NAND U32975 ( .A(n187), .B(n32187), .Z(n32189) );
  XOR U32976 ( .A(b[13]), .B(a[219]), .Z(n32336) );
  NAND U32977 ( .A(n37295), .B(n32336), .Z(n32188) );
  AND U32978 ( .A(n32189), .B(n32188), .Z(n32280) );
  NAND U32979 ( .A(n186), .B(n32190), .Z(n32192) );
  XOR U32980 ( .A(b[11]), .B(a[221]), .Z(n32339) );
  NAND U32981 ( .A(n37097), .B(n32339), .Z(n32191) );
  NAND U32982 ( .A(n32192), .B(n32191), .Z(n32279) );
  XNOR U32983 ( .A(n32280), .B(n32279), .Z(n32281) );
  NAND U32984 ( .A(n188), .B(n32193), .Z(n32195) );
  XOR U32985 ( .A(b[15]), .B(a[217]), .Z(n32342) );
  NAND U32986 ( .A(n37382), .B(n32342), .Z(n32194) );
  AND U32987 ( .A(n32195), .B(n32194), .Z(n32276) );
  NAND U32988 ( .A(n38064), .B(n32196), .Z(n32198) );
  XOR U32989 ( .A(b[21]), .B(a[211]), .Z(n32345) );
  NAND U32990 ( .A(n37993), .B(n32345), .Z(n32197) );
  AND U32991 ( .A(n32198), .B(n32197), .Z(n32274) );
  NAND U32992 ( .A(n185), .B(n32199), .Z(n32201) );
  XOR U32993 ( .A(b[9]), .B(a[223]), .Z(n32348) );
  NAND U32994 ( .A(n36805), .B(n32348), .Z(n32200) );
  NAND U32995 ( .A(n32201), .B(n32200), .Z(n32273) );
  XNOR U32996 ( .A(n32274), .B(n32273), .Z(n32275) );
  XOR U32997 ( .A(n32276), .B(n32275), .Z(n32282) );
  XOR U32998 ( .A(n32281), .B(n32282), .Z(n32288) );
  XOR U32999 ( .A(n32287), .B(n32288), .Z(n32300) );
  XNOR U33000 ( .A(n32299), .B(n32300), .Z(n32231) );
  XNOR U33001 ( .A(n32232), .B(n32231), .Z(n32233) );
  XOR U33002 ( .A(n32234), .B(n32233), .Z(n32352) );
  XNOR U33003 ( .A(n32351), .B(n32352), .Z(n32353) );
  XNOR U33004 ( .A(n32354), .B(n32353), .Z(n32227) );
  XOR U33005 ( .A(n32228), .B(n32227), .Z(n32220) );
  NANDN U33006 ( .A(n32203), .B(n32202), .Z(n32207) );
  OR U33007 ( .A(n32205), .B(n32204), .Z(n32206) );
  AND U33008 ( .A(n32207), .B(n32206), .Z(n32219) );
  XNOR U33009 ( .A(n32220), .B(n32219), .Z(n32221) );
  XNOR U33010 ( .A(n32222), .B(n32221), .Z(n32213) );
  XNOR U33011 ( .A(n32214), .B(n32213), .Z(n32215) );
  XNOR U33012 ( .A(n32216), .B(n32215), .Z(n32357) );
  XNOR U33013 ( .A(sreg[455]), .B(n32357), .Z(n32359) );
  NANDN U33014 ( .A(sreg[454]), .B(n32208), .Z(n32212) );
  NAND U33015 ( .A(n32210), .B(n32209), .Z(n32211) );
  NAND U33016 ( .A(n32212), .B(n32211), .Z(n32358) );
  XNOR U33017 ( .A(n32359), .B(n32358), .Z(c[455]) );
  NANDN U33018 ( .A(n32214), .B(n32213), .Z(n32218) );
  NANDN U33019 ( .A(n32216), .B(n32215), .Z(n32217) );
  AND U33020 ( .A(n32218), .B(n32217), .Z(n32365) );
  NANDN U33021 ( .A(n32220), .B(n32219), .Z(n32224) );
  NANDN U33022 ( .A(n32222), .B(n32221), .Z(n32223) );
  AND U33023 ( .A(n32224), .B(n32223), .Z(n32363) );
  NANDN U33024 ( .A(n32226), .B(n32225), .Z(n32230) );
  NAND U33025 ( .A(n32228), .B(n32227), .Z(n32229) );
  AND U33026 ( .A(n32230), .B(n32229), .Z(n32370) );
  NANDN U33027 ( .A(n32232), .B(n32231), .Z(n32236) );
  NANDN U33028 ( .A(n32234), .B(n32233), .Z(n32235) );
  AND U33029 ( .A(n32236), .B(n32235), .Z(n32375) );
  NANDN U33030 ( .A(n32238), .B(n32237), .Z(n32242) );
  NAND U33031 ( .A(n32240), .B(n32239), .Z(n32241) );
  AND U33032 ( .A(n32242), .B(n32241), .Z(n32374) );
  XNOR U33033 ( .A(n32375), .B(n32374), .Z(n32377) );
  NANDN U33034 ( .A(n32244), .B(n32243), .Z(n32248) );
  NANDN U33035 ( .A(n32246), .B(n32245), .Z(n32247) );
  AND U33036 ( .A(n32248), .B(n32247), .Z(n32454) );
  NAND U33037 ( .A(n38385), .B(n32249), .Z(n32251) );
  XOR U33038 ( .A(b[27]), .B(a[206]), .Z(n32398) );
  NAND U33039 ( .A(n38343), .B(n32398), .Z(n32250) );
  AND U33040 ( .A(n32251), .B(n32250), .Z(n32461) );
  NAND U33041 ( .A(n183), .B(n32252), .Z(n32254) );
  XOR U33042 ( .A(b[5]), .B(a[228]), .Z(n32401) );
  NAND U33043 ( .A(n36296), .B(n32401), .Z(n32253) );
  AND U33044 ( .A(n32254), .B(n32253), .Z(n32459) );
  NAND U33045 ( .A(n190), .B(n32255), .Z(n32257) );
  XOR U33046 ( .A(b[19]), .B(a[214]), .Z(n32404) );
  NAND U33047 ( .A(n37821), .B(n32404), .Z(n32256) );
  NAND U33048 ( .A(n32257), .B(n32256), .Z(n32458) );
  XNOR U33049 ( .A(n32459), .B(n32458), .Z(n32460) );
  XNOR U33050 ( .A(n32461), .B(n32460), .Z(n32452) );
  NAND U33051 ( .A(n38470), .B(n32258), .Z(n32260) );
  XOR U33052 ( .A(b[31]), .B(a[202]), .Z(n32407) );
  NAND U33053 ( .A(n38453), .B(n32407), .Z(n32259) );
  AND U33054 ( .A(n32260), .B(n32259), .Z(n32419) );
  NAND U33055 ( .A(n181), .B(n32261), .Z(n32263) );
  XOR U33056 ( .A(a[230]), .B(b[3]), .Z(n32410) );
  NAND U33057 ( .A(n182), .B(n32410), .Z(n32262) );
  AND U33058 ( .A(n32263), .B(n32262), .Z(n32417) );
  NAND U33059 ( .A(n189), .B(n32264), .Z(n32266) );
  XOR U33060 ( .A(b[17]), .B(a[216]), .Z(n32413) );
  NAND U33061 ( .A(n37652), .B(n32413), .Z(n32265) );
  NAND U33062 ( .A(n32266), .B(n32265), .Z(n32416) );
  XNOR U33063 ( .A(n32417), .B(n32416), .Z(n32418) );
  XOR U33064 ( .A(n32419), .B(n32418), .Z(n32453) );
  XOR U33065 ( .A(n32452), .B(n32453), .Z(n32455) );
  XOR U33066 ( .A(n32454), .B(n32455), .Z(n32387) );
  NANDN U33067 ( .A(n32268), .B(n32267), .Z(n32272) );
  NANDN U33068 ( .A(n32270), .B(n32269), .Z(n32271) );
  AND U33069 ( .A(n32272), .B(n32271), .Z(n32440) );
  NANDN U33070 ( .A(n32274), .B(n32273), .Z(n32278) );
  NANDN U33071 ( .A(n32276), .B(n32275), .Z(n32277) );
  NAND U33072 ( .A(n32278), .B(n32277), .Z(n32441) );
  XNOR U33073 ( .A(n32440), .B(n32441), .Z(n32442) );
  NANDN U33074 ( .A(n32280), .B(n32279), .Z(n32284) );
  NANDN U33075 ( .A(n32282), .B(n32281), .Z(n32283) );
  NAND U33076 ( .A(n32284), .B(n32283), .Z(n32443) );
  XNOR U33077 ( .A(n32442), .B(n32443), .Z(n32386) );
  XNOR U33078 ( .A(n32387), .B(n32386), .Z(n32389) );
  NANDN U33079 ( .A(n32286), .B(n32285), .Z(n32290) );
  NANDN U33080 ( .A(n32288), .B(n32287), .Z(n32289) );
  AND U33081 ( .A(n32290), .B(n32289), .Z(n32388) );
  XOR U33082 ( .A(n32389), .B(n32388), .Z(n32500) );
  NANDN U33083 ( .A(n32292), .B(n32291), .Z(n32296) );
  NANDN U33084 ( .A(n32294), .B(n32293), .Z(n32295) );
  AND U33085 ( .A(n32296), .B(n32295), .Z(n32497) );
  NANDN U33086 ( .A(n32298), .B(n32297), .Z(n32302) );
  NANDN U33087 ( .A(n32300), .B(n32299), .Z(n32301) );
  AND U33088 ( .A(n32302), .B(n32301), .Z(n32383) );
  NANDN U33089 ( .A(n32304), .B(n32303), .Z(n32308) );
  OR U33090 ( .A(n32306), .B(n32305), .Z(n32307) );
  AND U33091 ( .A(n32308), .B(n32307), .Z(n32381) );
  NANDN U33092 ( .A(n32310), .B(n32309), .Z(n32314) );
  NANDN U33093 ( .A(n32312), .B(n32311), .Z(n32313) );
  AND U33094 ( .A(n32314), .B(n32313), .Z(n32447) );
  NANDN U33095 ( .A(n32316), .B(n32315), .Z(n32320) );
  NANDN U33096 ( .A(n32318), .B(n32317), .Z(n32319) );
  NAND U33097 ( .A(n32320), .B(n32319), .Z(n32446) );
  XNOR U33098 ( .A(n32447), .B(n32446), .Z(n32448) );
  NAND U33099 ( .A(b[0]), .B(a[232]), .Z(n32321) );
  XNOR U33100 ( .A(b[1]), .B(n32321), .Z(n32323) );
  NANDN U33101 ( .A(b[0]), .B(a[231]), .Z(n32322) );
  NAND U33102 ( .A(n32323), .B(n32322), .Z(n32395) );
  NAND U33103 ( .A(n194), .B(n32324), .Z(n32326) );
  XOR U33104 ( .A(b[29]), .B(a[204]), .Z(n32470) );
  NAND U33105 ( .A(n38456), .B(n32470), .Z(n32325) );
  AND U33106 ( .A(n32326), .B(n32325), .Z(n32393) );
  AND U33107 ( .A(b[31]), .B(a[200]), .Z(n32392) );
  XNOR U33108 ( .A(n32393), .B(n32392), .Z(n32394) );
  XNOR U33109 ( .A(n32395), .B(n32394), .Z(n32434) );
  NAND U33110 ( .A(n38185), .B(n32327), .Z(n32329) );
  XOR U33111 ( .A(b[23]), .B(a[210]), .Z(n32473) );
  NAND U33112 ( .A(n38132), .B(n32473), .Z(n32328) );
  AND U33113 ( .A(n32329), .B(n32328), .Z(n32467) );
  NAND U33114 ( .A(n184), .B(n32330), .Z(n32332) );
  XOR U33115 ( .A(b[7]), .B(a[226]), .Z(n32476) );
  NAND U33116 ( .A(n36592), .B(n32476), .Z(n32331) );
  AND U33117 ( .A(n32332), .B(n32331), .Z(n32465) );
  NAND U33118 ( .A(n38289), .B(n32333), .Z(n32335) );
  XOR U33119 ( .A(b[25]), .B(a[208]), .Z(n32479) );
  NAND U33120 ( .A(n38247), .B(n32479), .Z(n32334) );
  NAND U33121 ( .A(n32335), .B(n32334), .Z(n32464) );
  XNOR U33122 ( .A(n32465), .B(n32464), .Z(n32466) );
  XOR U33123 ( .A(n32467), .B(n32466), .Z(n32435) );
  XNOR U33124 ( .A(n32434), .B(n32435), .Z(n32436) );
  NAND U33125 ( .A(n187), .B(n32336), .Z(n32338) );
  XOR U33126 ( .A(b[13]), .B(a[220]), .Z(n32482) );
  NAND U33127 ( .A(n37295), .B(n32482), .Z(n32337) );
  AND U33128 ( .A(n32338), .B(n32337), .Z(n32429) );
  NAND U33129 ( .A(n186), .B(n32339), .Z(n32341) );
  XOR U33130 ( .A(b[11]), .B(a[222]), .Z(n32485) );
  NAND U33131 ( .A(n37097), .B(n32485), .Z(n32340) );
  NAND U33132 ( .A(n32341), .B(n32340), .Z(n32428) );
  XNOR U33133 ( .A(n32429), .B(n32428), .Z(n32430) );
  NAND U33134 ( .A(n188), .B(n32342), .Z(n32344) );
  XOR U33135 ( .A(b[15]), .B(a[218]), .Z(n32488) );
  NAND U33136 ( .A(n37382), .B(n32488), .Z(n32343) );
  AND U33137 ( .A(n32344), .B(n32343), .Z(n32425) );
  NAND U33138 ( .A(n38064), .B(n32345), .Z(n32347) );
  XOR U33139 ( .A(b[21]), .B(a[212]), .Z(n32491) );
  NAND U33140 ( .A(n37993), .B(n32491), .Z(n32346) );
  AND U33141 ( .A(n32347), .B(n32346), .Z(n32423) );
  NAND U33142 ( .A(n185), .B(n32348), .Z(n32350) );
  XOR U33143 ( .A(b[9]), .B(a[224]), .Z(n32494) );
  NAND U33144 ( .A(n36805), .B(n32494), .Z(n32349) );
  NAND U33145 ( .A(n32350), .B(n32349), .Z(n32422) );
  XNOR U33146 ( .A(n32423), .B(n32422), .Z(n32424) );
  XOR U33147 ( .A(n32425), .B(n32424), .Z(n32431) );
  XOR U33148 ( .A(n32430), .B(n32431), .Z(n32437) );
  XOR U33149 ( .A(n32436), .B(n32437), .Z(n32449) );
  XNOR U33150 ( .A(n32448), .B(n32449), .Z(n32380) );
  XNOR U33151 ( .A(n32381), .B(n32380), .Z(n32382) );
  XOR U33152 ( .A(n32383), .B(n32382), .Z(n32498) );
  XNOR U33153 ( .A(n32497), .B(n32498), .Z(n32499) );
  XNOR U33154 ( .A(n32500), .B(n32499), .Z(n32376) );
  XOR U33155 ( .A(n32377), .B(n32376), .Z(n32369) );
  NANDN U33156 ( .A(n32352), .B(n32351), .Z(n32356) );
  NANDN U33157 ( .A(n32354), .B(n32353), .Z(n32355) );
  AND U33158 ( .A(n32356), .B(n32355), .Z(n32368) );
  XOR U33159 ( .A(n32369), .B(n32368), .Z(n32371) );
  XNOR U33160 ( .A(n32370), .B(n32371), .Z(n32362) );
  XNOR U33161 ( .A(n32363), .B(n32362), .Z(n32364) );
  XNOR U33162 ( .A(n32365), .B(n32364), .Z(n32503) );
  XNOR U33163 ( .A(sreg[456]), .B(n32503), .Z(n32505) );
  NANDN U33164 ( .A(sreg[455]), .B(n32357), .Z(n32361) );
  NAND U33165 ( .A(n32359), .B(n32358), .Z(n32360) );
  NAND U33166 ( .A(n32361), .B(n32360), .Z(n32504) );
  XNOR U33167 ( .A(n32505), .B(n32504), .Z(c[456]) );
  NANDN U33168 ( .A(n32363), .B(n32362), .Z(n32367) );
  NANDN U33169 ( .A(n32365), .B(n32364), .Z(n32366) );
  AND U33170 ( .A(n32367), .B(n32366), .Z(n32511) );
  NANDN U33171 ( .A(n32369), .B(n32368), .Z(n32373) );
  NANDN U33172 ( .A(n32371), .B(n32370), .Z(n32372) );
  AND U33173 ( .A(n32373), .B(n32372), .Z(n32509) );
  NANDN U33174 ( .A(n32375), .B(n32374), .Z(n32379) );
  NAND U33175 ( .A(n32377), .B(n32376), .Z(n32378) );
  AND U33176 ( .A(n32379), .B(n32378), .Z(n32516) );
  NANDN U33177 ( .A(n32381), .B(n32380), .Z(n32385) );
  NANDN U33178 ( .A(n32383), .B(n32382), .Z(n32384) );
  AND U33179 ( .A(n32385), .B(n32384), .Z(n32521) );
  NANDN U33180 ( .A(n32387), .B(n32386), .Z(n32391) );
  NAND U33181 ( .A(n32389), .B(n32388), .Z(n32390) );
  AND U33182 ( .A(n32391), .B(n32390), .Z(n32520) );
  XNOR U33183 ( .A(n32521), .B(n32520), .Z(n32523) );
  NANDN U33184 ( .A(n32393), .B(n32392), .Z(n32397) );
  NANDN U33185 ( .A(n32395), .B(n32394), .Z(n32396) );
  AND U33186 ( .A(n32397), .B(n32396), .Z(n32598) );
  NAND U33187 ( .A(n38385), .B(n32398), .Z(n32400) );
  XOR U33188 ( .A(b[27]), .B(a[207]), .Z(n32544) );
  NAND U33189 ( .A(n38343), .B(n32544), .Z(n32399) );
  AND U33190 ( .A(n32400), .B(n32399), .Z(n32605) );
  NAND U33191 ( .A(n183), .B(n32401), .Z(n32403) );
  XOR U33192 ( .A(b[5]), .B(a[229]), .Z(n32547) );
  NAND U33193 ( .A(n36296), .B(n32547), .Z(n32402) );
  AND U33194 ( .A(n32403), .B(n32402), .Z(n32603) );
  NAND U33195 ( .A(n190), .B(n32404), .Z(n32406) );
  XOR U33196 ( .A(b[19]), .B(a[215]), .Z(n32550) );
  NAND U33197 ( .A(n37821), .B(n32550), .Z(n32405) );
  NAND U33198 ( .A(n32406), .B(n32405), .Z(n32602) );
  XNOR U33199 ( .A(n32603), .B(n32602), .Z(n32604) );
  XNOR U33200 ( .A(n32605), .B(n32604), .Z(n32596) );
  NAND U33201 ( .A(n38470), .B(n32407), .Z(n32409) );
  XOR U33202 ( .A(b[31]), .B(a[203]), .Z(n32553) );
  NAND U33203 ( .A(n38453), .B(n32553), .Z(n32408) );
  AND U33204 ( .A(n32409), .B(n32408), .Z(n32565) );
  NAND U33205 ( .A(n181), .B(n32410), .Z(n32412) );
  XOR U33206 ( .A(a[231]), .B(b[3]), .Z(n32556) );
  NAND U33207 ( .A(n182), .B(n32556), .Z(n32411) );
  AND U33208 ( .A(n32412), .B(n32411), .Z(n32563) );
  NAND U33209 ( .A(n189), .B(n32413), .Z(n32415) );
  XOR U33210 ( .A(b[17]), .B(a[217]), .Z(n32559) );
  NAND U33211 ( .A(n37652), .B(n32559), .Z(n32414) );
  NAND U33212 ( .A(n32415), .B(n32414), .Z(n32562) );
  XNOR U33213 ( .A(n32563), .B(n32562), .Z(n32564) );
  XOR U33214 ( .A(n32565), .B(n32564), .Z(n32597) );
  XOR U33215 ( .A(n32596), .B(n32597), .Z(n32599) );
  XOR U33216 ( .A(n32598), .B(n32599), .Z(n32533) );
  NANDN U33217 ( .A(n32417), .B(n32416), .Z(n32421) );
  NANDN U33218 ( .A(n32419), .B(n32418), .Z(n32420) );
  AND U33219 ( .A(n32421), .B(n32420), .Z(n32586) );
  NANDN U33220 ( .A(n32423), .B(n32422), .Z(n32427) );
  NANDN U33221 ( .A(n32425), .B(n32424), .Z(n32426) );
  NAND U33222 ( .A(n32427), .B(n32426), .Z(n32587) );
  XNOR U33223 ( .A(n32586), .B(n32587), .Z(n32588) );
  NANDN U33224 ( .A(n32429), .B(n32428), .Z(n32433) );
  NANDN U33225 ( .A(n32431), .B(n32430), .Z(n32432) );
  NAND U33226 ( .A(n32433), .B(n32432), .Z(n32589) );
  XNOR U33227 ( .A(n32588), .B(n32589), .Z(n32532) );
  XNOR U33228 ( .A(n32533), .B(n32532), .Z(n32535) );
  NANDN U33229 ( .A(n32435), .B(n32434), .Z(n32439) );
  NANDN U33230 ( .A(n32437), .B(n32436), .Z(n32438) );
  AND U33231 ( .A(n32439), .B(n32438), .Z(n32534) );
  XOR U33232 ( .A(n32535), .B(n32534), .Z(n32647) );
  NANDN U33233 ( .A(n32441), .B(n32440), .Z(n32445) );
  NANDN U33234 ( .A(n32443), .B(n32442), .Z(n32444) );
  AND U33235 ( .A(n32445), .B(n32444), .Z(n32644) );
  NANDN U33236 ( .A(n32447), .B(n32446), .Z(n32451) );
  NANDN U33237 ( .A(n32449), .B(n32448), .Z(n32450) );
  AND U33238 ( .A(n32451), .B(n32450), .Z(n32529) );
  NANDN U33239 ( .A(n32453), .B(n32452), .Z(n32457) );
  OR U33240 ( .A(n32455), .B(n32454), .Z(n32456) );
  AND U33241 ( .A(n32457), .B(n32456), .Z(n32527) );
  NANDN U33242 ( .A(n32459), .B(n32458), .Z(n32463) );
  NANDN U33243 ( .A(n32461), .B(n32460), .Z(n32462) );
  AND U33244 ( .A(n32463), .B(n32462), .Z(n32593) );
  NANDN U33245 ( .A(n32465), .B(n32464), .Z(n32469) );
  NANDN U33246 ( .A(n32467), .B(n32466), .Z(n32468) );
  NAND U33247 ( .A(n32469), .B(n32468), .Z(n32592) );
  XNOR U33248 ( .A(n32593), .B(n32592), .Z(n32595) );
  NAND U33249 ( .A(n194), .B(n32470), .Z(n32472) );
  XOR U33250 ( .A(b[29]), .B(a[205]), .Z(n32617) );
  NAND U33251 ( .A(n38456), .B(n32617), .Z(n32471) );
  AND U33252 ( .A(n32472), .B(n32471), .Z(n32539) );
  AND U33253 ( .A(b[31]), .B(a[201]), .Z(n32538) );
  XOR U33254 ( .A(n32539), .B(n32538), .Z(n32541) );
  XNOR U33255 ( .A(n32540), .B(n32541), .Z(n32581) );
  NAND U33256 ( .A(n38185), .B(n32473), .Z(n32475) );
  XOR U33257 ( .A(b[23]), .B(a[211]), .Z(n32620) );
  NAND U33258 ( .A(n38132), .B(n32620), .Z(n32474) );
  AND U33259 ( .A(n32475), .B(n32474), .Z(n32610) );
  NAND U33260 ( .A(n184), .B(n32476), .Z(n32478) );
  XOR U33261 ( .A(b[7]), .B(a[227]), .Z(n32623) );
  NAND U33262 ( .A(n36592), .B(n32623), .Z(n32477) );
  AND U33263 ( .A(n32478), .B(n32477), .Z(n32609) );
  NAND U33264 ( .A(n38289), .B(n32479), .Z(n32481) );
  XOR U33265 ( .A(b[25]), .B(a[209]), .Z(n32626) );
  NAND U33266 ( .A(n38247), .B(n32626), .Z(n32480) );
  NAND U33267 ( .A(n32481), .B(n32480), .Z(n32608) );
  XOR U33268 ( .A(n32609), .B(n32608), .Z(n32611) );
  XOR U33269 ( .A(n32610), .B(n32611), .Z(n32580) );
  XOR U33270 ( .A(n32581), .B(n32580), .Z(n32583) );
  NAND U33271 ( .A(n187), .B(n32482), .Z(n32484) );
  XOR U33272 ( .A(b[13]), .B(a[221]), .Z(n32629) );
  NAND U33273 ( .A(n37295), .B(n32629), .Z(n32483) );
  AND U33274 ( .A(n32484), .B(n32483), .Z(n32575) );
  NAND U33275 ( .A(n186), .B(n32485), .Z(n32487) );
  XOR U33276 ( .A(b[11]), .B(a[223]), .Z(n32632) );
  NAND U33277 ( .A(n37097), .B(n32632), .Z(n32486) );
  NAND U33278 ( .A(n32487), .B(n32486), .Z(n32574) );
  XNOR U33279 ( .A(n32575), .B(n32574), .Z(n32577) );
  NAND U33280 ( .A(n188), .B(n32488), .Z(n32490) );
  XOR U33281 ( .A(b[15]), .B(a[219]), .Z(n32635) );
  NAND U33282 ( .A(n37382), .B(n32635), .Z(n32489) );
  AND U33283 ( .A(n32490), .B(n32489), .Z(n32571) );
  NAND U33284 ( .A(n38064), .B(n32491), .Z(n32493) );
  XOR U33285 ( .A(b[21]), .B(a[213]), .Z(n32638) );
  NAND U33286 ( .A(n37993), .B(n32638), .Z(n32492) );
  AND U33287 ( .A(n32493), .B(n32492), .Z(n32569) );
  NAND U33288 ( .A(n185), .B(n32494), .Z(n32496) );
  XOR U33289 ( .A(b[9]), .B(a[225]), .Z(n32641) );
  NAND U33290 ( .A(n36805), .B(n32641), .Z(n32495) );
  NAND U33291 ( .A(n32496), .B(n32495), .Z(n32568) );
  XNOR U33292 ( .A(n32569), .B(n32568), .Z(n32570) );
  XNOR U33293 ( .A(n32571), .B(n32570), .Z(n32576) );
  XOR U33294 ( .A(n32577), .B(n32576), .Z(n32582) );
  XNOR U33295 ( .A(n32583), .B(n32582), .Z(n32594) );
  XNOR U33296 ( .A(n32595), .B(n32594), .Z(n32526) );
  XNOR U33297 ( .A(n32527), .B(n32526), .Z(n32528) );
  XOR U33298 ( .A(n32529), .B(n32528), .Z(n32645) );
  XNOR U33299 ( .A(n32644), .B(n32645), .Z(n32646) );
  XNOR U33300 ( .A(n32647), .B(n32646), .Z(n32522) );
  XOR U33301 ( .A(n32523), .B(n32522), .Z(n32515) );
  NANDN U33302 ( .A(n32498), .B(n32497), .Z(n32502) );
  NANDN U33303 ( .A(n32500), .B(n32499), .Z(n32501) );
  AND U33304 ( .A(n32502), .B(n32501), .Z(n32514) );
  XOR U33305 ( .A(n32515), .B(n32514), .Z(n32517) );
  XNOR U33306 ( .A(n32516), .B(n32517), .Z(n32508) );
  XNOR U33307 ( .A(n32509), .B(n32508), .Z(n32510) );
  XNOR U33308 ( .A(n32511), .B(n32510), .Z(n32650) );
  XNOR U33309 ( .A(sreg[457]), .B(n32650), .Z(n32652) );
  NANDN U33310 ( .A(sreg[456]), .B(n32503), .Z(n32507) );
  NAND U33311 ( .A(n32505), .B(n32504), .Z(n32506) );
  NAND U33312 ( .A(n32507), .B(n32506), .Z(n32651) );
  XNOR U33313 ( .A(n32652), .B(n32651), .Z(c[457]) );
  NANDN U33314 ( .A(n32509), .B(n32508), .Z(n32513) );
  NANDN U33315 ( .A(n32511), .B(n32510), .Z(n32512) );
  AND U33316 ( .A(n32513), .B(n32512), .Z(n32658) );
  NANDN U33317 ( .A(n32515), .B(n32514), .Z(n32519) );
  NANDN U33318 ( .A(n32517), .B(n32516), .Z(n32518) );
  AND U33319 ( .A(n32519), .B(n32518), .Z(n32656) );
  NANDN U33320 ( .A(n32521), .B(n32520), .Z(n32525) );
  NAND U33321 ( .A(n32523), .B(n32522), .Z(n32524) );
  AND U33322 ( .A(n32525), .B(n32524), .Z(n32663) );
  NANDN U33323 ( .A(n32527), .B(n32526), .Z(n32531) );
  NANDN U33324 ( .A(n32529), .B(n32528), .Z(n32530) );
  AND U33325 ( .A(n32531), .B(n32530), .Z(n32794) );
  NANDN U33326 ( .A(n32533), .B(n32532), .Z(n32537) );
  NAND U33327 ( .A(n32535), .B(n32534), .Z(n32536) );
  AND U33328 ( .A(n32537), .B(n32536), .Z(n32793) );
  XNOR U33329 ( .A(n32794), .B(n32793), .Z(n32796) );
  NANDN U33330 ( .A(n32539), .B(n32538), .Z(n32543) );
  NANDN U33331 ( .A(n32541), .B(n32540), .Z(n32542) );
  AND U33332 ( .A(n32543), .B(n32542), .Z(n32729) );
  NAND U33333 ( .A(n38385), .B(n32544), .Z(n32546) );
  XOR U33334 ( .A(b[27]), .B(a[208]), .Z(n32673) );
  NAND U33335 ( .A(n38343), .B(n32673), .Z(n32545) );
  AND U33336 ( .A(n32546), .B(n32545), .Z(n32736) );
  NAND U33337 ( .A(n183), .B(n32547), .Z(n32549) );
  XOR U33338 ( .A(b[5]), .B(a[230]), .Z(n32676) );
  NAND U33339 ( .A(n36296), .B(n32676), .Z(n32548) );
  AND U33340 ( .A(n32549), .B(n32548), .Z(n32734) );
  NAND U33341 ( .A(n190), .B(n32550), .Z(n32552) );
  XOR U33342 ( .A(b[19]), .B(a[216]), .Z(n32679) );
  NAND U33343 ( .A(n37821), .B(n32679), .Z(n32551) );
  NAND U33344 ( .A(n32552), .B(n32551), .Z(n32733) );
  XNOR U33345 ( .A(n32734), .B(n32733), .Z(n32735) );
  XNOR U33346 ( .A(n32736), .B(n32735), .Z(n32727) );
  NAND U33347 ( .A(n38470), .B(n32553), .Z(n32555) );
  XOR U33348 ( .A(b[31]), .B(a[204]), .Z(n32682) );
  NAND U33349 ( .A(n38453), .B(n32682), .Z(n32554) );
  AND U33350 ( .A(n32555), .B(n32554), .Z(n32694) );
  NAND U33351 ( .A(n181), .B(n32556), .Z(n32558) );
  XOR U33352 ( .A(a[232]), .B(b[3]), .Z(n32685) );
  NAND U33353 ( .A(n182), .B(n32685), .Z(n32557) );
  AND U33354 ( .A(n32558), .B(n32557), .Z(n32692) );
  NAND U33355 ( .A(n189), .B(n32559), .Z(n32561) );
  XOR U33356 ( .A(b[17]), .B(a[218]), .Z(n32688) );
  NAND U33357 ( .A(n37652), .B(n32688), .Z(n32560) );
  NAND U33358 ( .A(n32561), .B(n32560), .Z(n32691) );
  XNOR U33359 ( .A(n32692), .B(n32691), .Z(n32693) );
  XOR U33360 ( .A(n32694), .B(n32693), .Z(n32728) );
  XOR U33361 ( .A(n32727), .B(n32728), .Z(n32730) );
  XOR U33362 ( .A(n32729), .B(n32730), .Z(n32776) );
  NANDN U33363 ( .A(n32563), .B(n32562), .Z(n32567) );
  NANDN U33364 ( .A(n32565), .B(n32564), .Z(n32566) );
  AND U33365 ( .A(n32567), .B(n32566), .Z(n32715) );
  NANDN U33366 ( .A(n32569), .B(n32568), .Z(n32573) );
  NANDN U33367 ( .A(n32571), .B(n32570), .Z(n32572) );
  NAND U33368 ( .A(n32573), .B(n32572), .Z(n32716) );
  XNOR U33369 ( .A(n32715), .B(n32716), .Z(n32717) );
  NANDN U33370 ( .A(n32575), .B(n32574), .Z(n32579) );
  NAND U33371 ( .A(n32577), .B(n32576), .Z(n32578) );
  NAND U33372 ( .A(n32579), .B(n32578), .Z(n32718) );
  XNOR U33373 ( .A(n32717), .B(n32718), .Z(n32775) );
  XNOR U33374 ( .A(n32776), .B(n32775), .Z(n32778) );
  NAND U33375 ( .A(n32581), .B(n32580), .Z(n32585) );
  NAND U33376 ( .A(n32583), .B(n32582), .Z(n32584) );
  AND U33377 ( .A(n32585), .B(n32584), .Z(n32777) );
  XOR U33378 ( .A(n32778), .B(n32777), .Z(n32790) );
  NANDN U33379 ( .A(n32587), .B(n32586), .Z(n32591) );
  NANDN U33380 ( .A(n32589), .B(n32588), .Z(n32590) );
  AND U33381 ( .A(n32591), .B(n32590), .Z(n32787) );
  NANDN U33382 ( .A(n32597), .B(n32596), .Z(n32601) );
  OR U33383 ( .A(n32599), .B(n32598), .Z(n32600) );
  AND U33384 ( .A(n32601), .B(n32600), .Z(n32782) );
  NANDN U33385 ( .A(n32603), .B(n32602), .Z(n32607) );
  NANDN U33386 ( .A(n32605), .B(n32604), .Z(n32606) );
  AND U33387 ( .A(n32607), .B(n32606), .Z(n32722) );
  NANDN U33388 ( .A(n32609), .B(n32608), .Z(n32613) );
  OR U33389 ( .A(n32611), .B(n32610), .Z(n32612) );
  NAND U33390 ( .A(n32613), .B(n32612), .Z(n32721) );
  XNOR U33391 ( .A(n32722), .B(n32721), .Z(n32723) );
  NAND U33392 ( .A(b[0]), .B(a[234]), .Z(n32614) );
  XNOR U33393 ( .A(b[1]), .B(n32614), .Z(n32616) );
  NANDN U33394 ( .A(b[0]), .B(a[233]), .Z(n32615) );
  NAND U33395 ( .A(n32616), .B(n32615), .Z(n32670) );
  NAND U33396 ( .A(n194), .B(n32617), .Z(n32619) );
  XOR U33397 ( .A(b[29]), .B(a[206]), .Z(n32748) );
  NAND U33398 ( .A(n38456), .B(n32748), .Z(n32618) );
  AND U33399 ( .A(n32619), .B(n32618), .Z(n32668) );
  AND U33400 ( .A(b[31]), .B(a[202]), .Z(n32667) );
  XNOR U33401 ( .A(n32668), .B(n32667), .Z(n32669) );
  XNOR U33402 ( .A(n32670), .B(n32669), .Z(n32709) );
  NAND U33403 ( .A(n38185), .B(n32620), .Z(n32622) );
  XOR U33404 ( .A(b[23]), .B(a[212]), .Z(n32751) );
  NAND U33405 ( .A(n38132), .B(n32751), .Z(n32621) );
  AND U33406 ( .A(n32622), .B(n32621), .Z(n32742) );
  NAND U33407 ( .A(n184), .B(n32623), .Z(n32625) );
  XOR U33408 ( .A(b[7]), .B(a[228]), .Z(n32754) );
  NAND U33409 ( .A(n36592), .B(n32754), .Z(n32624) );
  AND U33410 ( .A(n32625), .B(n32624), .Z(n32740) );
  NAND U33411 ( .A(n38289), .B(n32626), .Z(n32628) );
  XOR U33412 ( .A(b[25]), .B(a[210]), .Z(n32757) );
  NAND U33413 ( .A(n38247), .B(n32757), .Z(n32627) );
  NAND U33414 ( .A(n32628), .B(n32627), .Z(n32739) );
  XNOR U33415 ( .A(n32740), .B(n32739), .Z(n32741) );
  XOR U33416 ( .A(n32742), .B(n32741), .Z(n32710) );
  XNOR U33417 ( .A(n32709), .B(n32710), .Z(n32711) );
  NAND U33418 ( .A(n187), .B(n32629), .Z(n32631) );
  XOR U33419 ( .A(b[13]), .B(a[222]), .Z(n32760) );
  NAND U33420 ( .A(n37295), .B(n32760), .Z(n32630) );
  AND U33421 ( .A(n32631), .B(n32630), .Z(n32704) );
  NAND U33422 ( .A(n186), .B(n32632), .Z(n32634) );
  XOR U33423 ( .A(b[11]), .B(a[224]), .Z(n32763) );
  NAND U33424 ( .A(n37097), .B(n32763), .Z(n32633) );
  NAND U33425 ( .A(n32634), .B(n32633), .Z(n32703) );
  XNOR U33426 ( .A(n32704), .B(n32703), .Z(n32705) );
  NAND U33427 ( .A(n188), .B(n32635), .Z(n32637) );
  XOR U33428 ( .A(b[15]), .B(a[220]), .Z(n32766) );
  NAND U33429 ( .A(n37382), .B(n32766), .Z(n32636) );
  AND U33430 ( .A(n32637), .B(n32636), .Z(n32700) );
  NAND U33431 ( .A(n38064), .B(n32638), .Z(n32640) );
  XOR U33432 ( .A(b[21]), .B(a[214]), .Z(n32769) );
  NAND U33433 ( .A(n37993), .B(n32769), .Z(n32639) );
  AND U33434 ( .A(n32640), .B(n32639), .Z(n32698) );
  NAND U33435 ( .A(n185), .B(n32641), .Z(n32643) );
  XOR U33436 ( .A(b[9]), .B(a[226]), .Z(n32772) );
  NAND U33437 ( .A(n36805), .B(n32772), .Z(n32642) );
  NAND U33438 ( .A(n32643), .B(n32642), .Z(n32697) );
  XNOR U33439 ( .A(n32698), .B(n32697), .Z(n32699) );
  XOR U33440 ( .A(n32700), .B(n32699), .Z(n32706) );
  XOR U33441 ( .A(n32705), .B(n32706), .Z(n32712) );
  XOR U33442 ( .A(n32711), .B(n32712), .Z(n32724) );
  XNOR U33443 ( .A(n32723), .B(n32724), .Z(n32781) );
  XNOR U33444 ( .A(n32782), .B(n32781), .Z(n32783) );
  XOR U33445 ( .A(n32784), .B(n32783), .Z(n32788) );
  XNOR U33446 ( .A(n32787), .B(n32788), .Z(n32789) );
  XNOR U33447 ( .A(n32790), .B(n32789), .Z(n32795) );
  XOR U33448 ( .A(n32796), .B(n32795), .Z(n32662) );
  NANDN U33449 ( .A(n32645), .B(n32644), .Z(n32649) );
  NANDN U33450 ( .A(n32647), .B(n32646), .Z(n32648) );
  AND U33451 ( .A(n32649), .B(n32648), .Z(n32661) );
  XOR U33452 ( .A(n32662), .B(n32661), .Z(n32664) );
  XNOR U33453 ( .A(n32663), .B(n32664), .Z(n32655) );
  XNOR U33454 ( .A(n32656), .B(n32655), .Z(n32657) );
  XNOR U33455 ( .A(n32658), .B(n32657), .Z(n32799) );
  XNOR U33456 ( .A(sreg[458]), .B(n32799), .Z(n32801) );
  NANDN U33457 ( .A(sreg[457]), .B(n32650), .Z(n32654) );
  NAND U33458 ( .A(n32652), .B(n32651), .Z(n32653) );
  NAND U33459 ( .A(n32654), .B(n32653), .Z(n32800) );
  XNOR U33460 ( .A(n32801), .B(n32800), .Z(c[458]) );
  NANDN U33461 ( .A(n32656), .B(n32655), .Z(n32660) );
  NANDN U33462 ( .A(n32658), .B(n32657), .Z(n32659) );
  AND U33463 ( .A(n32660), .B(n32659), .Z(n32807) );
  NANDN U33464 ( .A(n32662), .B(n32661), .Z(n32666) );
  NANDN U33465 ( .A(n32664), .B(n32663), .Z(n32665) );
  AND U33466 ( .A(n32666), .B(n32665), .Z(n32805) );
  NANDN U33467 ( .A(n32668), .B(n32667), .Z(n32672) );
  NANDN U33468 ( .A(n32670), .B(n32669), .Z(n32671) );
  AND U33469 ( .A(n32672), .B(n32671), .Z(n32896) );
  NAND U33470 ( .A(n38385), .B(n32673), .Z(n32675) );
  XOR U33471 ( .A(b[27]), .B(a[209]), .Z(n32840) );
  NAND U33472 ( .A(n38343), .B(n32840), .Z(n32674) );
  AND U33473 ( .A(n32675), .B(n32674), .Z(n32903) );
  NAND U33474 ( .A(n183), .B(n32676), .Z(n32678) );
  XOR U33475 ( .A(b[5]), .B(a[231]), .Z(n32843) );
  NAND U33476 ( .A(n36296), .B(n32843), .Z(n32677) );
  AND U33477 ( .A(n32678), .B(n32677), .Z(n32901) );
  NAND U33478 ( .A(n190), .B(n32679), .Z(n32681) );
  XOR U33479 ( .A(b[19]), .B(a[217]), .Z(n32846) );
  NAND U33480 ( .A(n37821), .B(n32846), .Z(n32680) );
  NAND U33481 ( .A(n32681), .B(n32680), .Z(n32900) );
  XNOR U33482 ( .A(n32901), .B(n32900), .Z(n32902) );
  XNOR U33483 ( .A(n32903), .B(n32902), .Z(n32894) );
  NAND U33484 ( .A(n38470), .B(n32682), .Z(n32684) );
  XOR U33485 ( .A(b[31]), .B(a[205]), .Z(n32849) );
  NAND U33486 ( .A(n38453), .B(n32849), .Z(n32683) );
  AND U33487 ( .A(n32684), .B(n32683), .Z(n32861) );
  NAND U33488 ( .A(n181), .B(n32685), .Z(n32687) );
  XOR U33489 ( .A(a[233]), .B(b[3]), .Z(n32852) );
  NAND U33490 ( .A(n182), .B(n32852), .Z(n32686) );
  AND U33491 ( .A(n32687), .B(n32686), .Z(n32859) );
  NAND U33492 ( .A(n189), .B(n32688), .Z(n32690) );
  XOR U33493 ( .A(b[17]), .B(a[219]), .Z(n32855) );
  NAND U33494 ( .A(n37652), .B(n32855), .Z(n32689) );
  NAND U33495 ( .A(n32690), .B(n32689), .Z(n32858) );
  XNOR U33496 ( .A(n32859), .B(n32858), .Z(n32860) );
  XOR U33497 ( .A(n32861), .B(n32860), .Z(n32895) );
  XOR U33498 ( .A(n32894), .B(n32895), .Z(n32897) );
  XOR U33499 ( .A(n32896), .B(n32897), .Z(n32829) );
  NANDN U33500 ( .A(n32692), .B(n32691), .Z(n32696) );
  NANDN U33501 ( .A(n32694), .B(n32693), .Z(n32695) );
  AND U33502 ( .A(n32696), .B(n32695), .Z(n32882) );
  NANDN U33503 ( .A(n32698), .B(n32697), .Z(n32702) );
  NANDN U33504 ( .A(n32700), .B(n32699), .Z(n32701) );
  NAND U33505 ( .A(n32702), .B(n32701), .Z(n32883) );
  XNOR U33506 ( .A(n32882), .B(n32883), .Z(n32884) );
  NANDN U33507 ( .A(n32704), .B(n32703), .Z(n32708) );
  NANDN U33508 ( .A(n32706), .B(n32705), .Z(n32707) );
  NAND U33509 ( .A(n32708), .B(n32707), .Z(n32885) );
  XNOR U33510 ( .A(n32884), .B(n32885), .Z(n32828) );
  XNOR U33511 ( .A(n32829), .B(n32828), .Z(n32831) );
  NANDN U33512 ( .A(n32710), .B(n32709), .Z(n32714) );
  NANDN U33513 ( .A(n32712), .B(n32711), .Z(n32713) );
  AND U33514 ( .A(n32714), .B(n32713), .Z(n32830) );
  XOR U33515 ( .A(n32831), .B(n32830), .Z(n32944) );
  NANDN U33516 ( .A(n32716), .B(n32715), .Z(n32720) );
  NANDN U33517 ( .A(n32718), .B(n32717), .Z(n32719) );
  AND U33518 ( .A(n32720), .B(n32719), .Z(n32942) );
  NANDN U33519 ( .A(n32722), .B(n32721), .Z(n32726) );
  NANDN U33520 ( .A(n32724), .B(n32723), .Z(n32725) );
  AND U33521 ( .A(n32726), .B(n32725), .Z(n32825) );
  NANDN U33522 ( .A(n32728), .B(n32727), .Z(n32732) );
  OR U33523 ( .A(n32730), .B(n32729), .Z(n32731) );
  AND U33524 ( .A(n32732), .B(n32731), .Z(n32823) );
  NANDN U33525 ( .A(n32734), .B(n32733), .Z(n32738) );
  NANDN U33526 ( .A(n32736), .B(n32735), .Z(n32737) );
  AND U33527 ( .A(n32738), .B(n32737), .Z(n32889) );
  NANDN U33528 ( .A(n32740), .B(n32739), .Z(n32744) );
  NANDN U33529 ( .A(n32742), .B(n32741), .Z(n32743) );
  NAND U33530 ( .A(n32744), .B(n32743), .Z(n32888) );
  XNOR U33531 ( .A(n32889), .B(n32888), .Z(n32890) );
  NAND U33532 ( .A(b[0]), .B(a[235]), .Z(n32745) );
  XNOR U33533 ( .A(b[1]), .B(n32745), .Z(n32747) );
  NANDN U33534 ( .A(b[0]), .B(a[234]), .Z(n32746) );
  NAND U33535 ( .A(n32747), .B(n32746), .Z(n32837) );
  NAND U33536 ( .A(n194), .B(n32748), .Z(n32750) );
  XOR U33537 ( .A(b[29]), .B(a[207]), .Z(n32915) );
  NAND U33538 ( .A(n38456), .B(n32915), .Z(n32749) );
  AND U33539 ( .A(n32750), .B(n32749), .Z(n32835) );
  AND U33540 ( .A(b[31]), .B(a[203]), .Z(n32834) );
  XNOR U33541 ( .A(n32835), .B(n32834), .Z(n32836) );
  XNOR U33542 ( .A(n32837), .B(n32836), .Z(n32876) );
  NAND U33543 ( .A(n38185), .B(n32751), .Z(n32753) );
  XOR U33544 ( .A(b[23]), .B(a[213]), .Z(n32918) );
  NAND U33545 ( .A(n38132), .B(n32918), .Z(n32752) );
  AND U33546 ( .A(n32753), .B(n32752), .Z(n32909) );
  NAND U33547 ( .A(n184), .B(n32754), .Z(n32756) );
  XOR U33548 ( .A(b[7]), .B(a[229]), .Z(n32921) );
  NAND U33549 ( .A(n36592), .B(n32921), .Z(n32755) );
  AND U33550 ( .A(n32756), .B(n32755), .Z(n32907) );
  NAND U33551 ( .A(n38289), .B(n32757), .Z(n32759) );
  XOR U33552 ( .A(b[25]), .B(a[211]), .Z(n32924) );
  NAND U33553 ( .A(n38247), .B(n32924), .Z(n32758) );
  NAND U33554 ( .A(n32759), .B(n32758), .Z(n32906) );
  XNOR U33555 ( .A(n32907), .B(n32906), .Z(n32908) );
  XOR U33556 ( .A(n32909), .B(n32908), .Z(n32877) );
  XNOR U33557 ( .A(n32876), .B(n32877), .Z(n32878) );
  NAND U33558 ( .A(n187), .B(n32760), .Z(n32762) );
  XOR U33559 ( .A(b[13]), .B(a[223]), .Z(n32927) );
  NAND U33560 ( .A(n37295), .B(n32927), .Z(n32761) );
  AND U33561 ( .A(n32762), .B(n32761), .Z(n32871) );
  NAND U33562 ( .A(n186), .B(n32763), .Z(n32765) );
  XOR U33563 ( .A(b[11]), .B(a[225]), .Z(n32930) );
  NAND U33564 ( .A(n37097), .B(n32930), .Z(n32764) );
  NAND U33565 ( .A(n32765), .B(n32764), .Z(n32870) );
  XNOR U33566 ( .A(n32871), .B(n32870), .Z(n32872) );
  NAND U33567 ( .A(n188), .B(n32766), .Z(n32768) );
  XOR U33568 ( .A(b[15]), .B(a[221]), .Z(n32933) );
  NAND U33569 ( .A(n37382), .B(n32933), .Z(n32767) );
  AND U33570 ( .A(n32768), .B(n32767), .Z(n32867) );
  NAND U33571 ( .A(n38064), .B(n32769), .Z(n32771) );
  XOR U33572 ( .A(b[21]), .B(a[215]), .Z(n32936) );
  NAND U33573 ( .A(n37993), .B(n32936), .Z(n32770) );
  AND U33574 ( .A(n32771), .B(n32770), .Z(n32865) );
  NAND U33575 ( .A(n185), .B(n32772), .Z(n32774) );
  XOR U33576 ( .A(b[9]), .B(a[227]), .Z(n32939) );
  NAND U33577 ( .A(n36805), .B(n32939), .Z(n32773) );
  NAND U33578 ( .A(n32774), .B(n32773), .Z(n32864) );
  XNOR U33579 ( .A(n32865), .B(n32864), .Z(n32866) );
  XOR U33580 ( .A(n32867), .B(n32866), .Z(n32873) );
  XOR U33581 ( .A(n32872), .B(n32873), .Z(n32879) );
  XOR U33582 ( .A(n32878), .B(n32879), .Z(n32891) );
  XNOR U33583 ( .A(n32890), .B(n32891), .Z(n32822) );
  XNOR U33584 ( .A(n32823), .B(n32822), .Z(n32824) );
  XOR U33585 ( .A(n32825), .B(n32824), .Z(n32943) );
  XOR U33586 ( .A(n32942), .B(n32943), .Z(n32945) );
  XOR U33587 ( .A(n32944), .B(n32945), .Z(n32819) );
  NANDN U33588 ( .A(n32776), .B(n32775), .Z(n32780) );
  NAND U33589 ( .A(n32778), .B(n32777), .Z(n32779) );
  AND U33590 ( .A(n32780), .B(n32779), .Z(n32817) );
  NANDN U33591 ( .A(n32782), .B(n32781), .Z(n32786) );
  NANDN U33592 ( .A(n32784), .B(n32783), .Z(n32785) );
  AND U33593 ( .A(n32786), .B(n32785), .Z(n32816) );
  XNOR U33594 ( .A(n32817), .B(n32816), .Z(n32818) );
  XNOR U33595 ( .A(n32819), .B(n32818), .Z(n32810) );
  NANDN U33596 ( .A(n32788), .B(n32787), .Z(n32792) );
  NANDN U33597 ( .A(n32790), .B(n32789), .Z(n32791) );
  NAND U33598 ( .A(n32792), .B(n32791), .Z(n32811) );
  XNOR U33599 ( .A(n32810), .B(n32811), .Z(n32812) );
  NANDN U33600 ( .A(n32794), .B(n32793), .Z(n32798) );
  NAND U33601 ( .A(n32796), .B(n32795), .Z(n32797) );
  NAND U33602 ( .A(n32798), .B(n32797), .Z(n32813) );
  XNOR U33603 ( .A(n32812), .B(n32813), .Z(n32804) );
  XNOR U33604 ( .A(n32805), .B(n32804), .Z(n32806) );
  XNOR U33605 ( .A(n32807), .B(n32806), .Z(n32948) );
  XNOR U33606 ( .A(sreg[459]), .B(n32948), .Z(n32950) );
  NANDN U33607 ( .A(sreg[458]), .B(n32799), .Z(n32803) );
  NAND U33608 ( .A(n32801), .B(n32800), .Z(n32802) );
  NAND U33609 ( .A(n32803), .B(n32802), .Z(n32949) );
  XNOR U33610 ( .A(n32950), .B(n32949), .Z(c[459]) );
  NANDN U33611 ( .A(n32805), .B(n32804), .Z(n32809) );
  NANDN U33612 ( .A(n32807), .B(n32806), .Z(n32808) );
  AND U33613 ( .A(n32809), .B(n32808), .Z(n32956) );
  NANDN U33614 ( .A(n32811), .B(n32810), .Z(n32815) );
  NANDN U33615 ( .A(n32813), .B(n32812), .Z(n32814) );
  AND U33616 ( .A(n32815), .B(n32814), .Z(n32954) );
  NANDN U33617 ( .A(n32817), .B(n32816), .Z(n32821) );
  NANDN U33618 ( .A(n32819), .B(n32818), .Z(n32820) );
  AND U33619 ( .A(n32821), .B(n32820), .Z(n32962) );
  NANDN U33620 ( .A(n32823), .B(n32822), .Z(n32827) );
  NANDN U33621 ( .A(n32825), .B(n32824), .Z(n32826) );
  AND U33622 ( .A(n32827), .B(n32826), .Z(n32966) );
  NANDN U33623 ( .A(n32829), .B(n32828), .Z(n32833) );
  NAND U33624 ( .A(n32831), .B(n32830), .Z(n32832) );
  AND U33625 ( .A(n32833), .B(n32832), .Z(n32965) );
  XNOR U33626 ( .A(n32966), .B(n32965), .Z(n32968) );
  NANDN U33627 ( .A(n32835), .B(n32834), .Z(n32839) );
  NANDN U33628 ( .A(n32837), .B(n32836), .Z(n32838) );
  AND U33629 ( .A(n32839), .B(n32838), .Z(n33045) );
  NAND U33630 ( .A(n38385), .B(n32840), .Z(n32842) );
  XOR U33631 ( .A(b[27]), .B(a[210]), .Z(n32989) );
  NAND U33632 ( .A(n38343), .B(n32989), .Z(n32841) );
  AND U33633 ( .A(n32842), .B(n32841), .Z(n33052) );
  NAND U33634 ( .A(n183), .B(n32843), .Z(n32845) );
  XOR U33635 ( .A(a[232]), .B(b[5]), .Z(n32992) );
  NAND U33636 ( .A(n36296), .B(n32992), .Z(n32844) );
  AND U33637 ( .A(n32845), .B(n32844), .Z(n33050) );
  NAND U33638 ( .A(n190), .B(n32846), .Z(n32848) );
  XOR U33639 ( .A(b[19]), .B(a[218]), .Z(n32995) );
  NAND U33640 ( .A(n37821), .B(n32995), .Z(n32847) );
  NAND U33641 ( .A(n32848), .B(n32847), .Z(n33049) );
  XNOR U33642 ( .A(n33050), .B(n33049), .Z(n33051) );
  XNOR U33643 ( .A(n33052), .B(n33051), .Z(n33043) );
  NAND U33644 ( .A(n38470), .B(n32849), .Z(n32851) );
  XOR U33645 ( .A(b[31]), .B(a[206]), .Z(n32998) );
  NAND U33646 ( .A(n38453), .B(n32998), .Z(n32850) );
  AND U33647 ( .A(n32851), .B(n32850), .Z(n33010) );
  NAND U33648 ( .A(n181), .B(n32852), .Z(n32854) );
  XOR U33649 ( .A(a[234]), .B(b[3]), .Z(n33001) );
  NAND U33650 ( .A(n182), .B(n33001), .Z(n32853) );
  AND U33651 ( .A(n32854), .B(n32853), .Z(n33008) );
  NAND U33652 ( .A(n189), .B(n32855), .Z(n32857) );
  XOR U33653 ( .A(b[17]), .B(a[220]), .Z(n33004) );
  NAND U33654 ( .A(n37652), .B(n33004), .Z(n32856) );
  NAND U33655 ( .A(n32857), .B(n32856), .Z(n33007) );
  XNOR U33656 ( .A(n33008), .B(n33007), .Z(n33009) );
  XOR U33657 ( .A(n33010), .B(n33009), .Z(n33044) );
  XOR U33658 ( .A(n33043), .B(n33044), .Z(n33046) );
  XOR U33659 ( .A(n33045), .B(n33046), .Z(n32978) );
  NANDN U33660 ( .A(n32859), .B(n32858), .Z(n32863) );
  NANDN U33661 ( .A(n32861), .B(n32860), .Z(n32862) );
  AND U33662 ( .A(n32863), .B(n32862), .Z(n33031) );
  NANDN U33663 ( .A(n32865), .B(n32864), .Z(n32869) );
  NANDN U33664 ( .A(n32867), .B(n32866), .Z(n32868) );
  NAND U33665 ( .A(n32869), .B(n32868), .Z(n33032) );
  XNOR U33666 ( .A(n33031), .B(n33032), .Z(n33033) );
  NANDN U33667 ( .A(n32871), .B(n32870), .Z(n32875) );
  NANDN U33668 ( .A(n32873), .B(n32872), .Z(n32874) );
  NAND U33669 ( .A(n32875), .B(n32874), .Z(n33034) );
  XNOR U33670 ( .A(n33033), .B(n33034), .Z(n32977) );
  XNOR U33671 ( .A(n32978), .B(n32977), .Z(n32980) );
  NANDN U33672 ( .A(n32877), .B(n32876), .Z(n32881) );
  NANDN U33673 ( .A(n32879), .B(n32878), .Z(n32880) );
  AND U33674 ( .A(n32881), .B(n32880), .Z(n32979) );
  XOR U33675 ( .A(n32980), .B(n32979), .Z(n33094) );
  NANDN U33676 ( .A(n32883), .B(n32882), .Z(n32887) );
  NANDN U33677 ( .A(n32885), .B(n32884), .Z(n32886) );
  AND U33678 ( .A(n32887), .B(n32886), .Z(n33091) );
  NANDN U33679 ( .A(n32889), .B(n32888), .Z(n32893) );
  NANDN U33680 ( .A(n32891), .B(n32890), .Z(n32892) );
  AND U33681 ( .A(n32893), .B(n32892), .Z(n32974) );
  NANDN U33682 ( .A(n32895), .B(n32894), .Z(n32899) );
  OR U33683 ( .A(n32897), .B(n32896), .Z(n32898) );
  AND U33684 ( .A(n32899), .B(n32898), .Z(n32972) );
  NANDN U33685 ( .A(n32901), .B(n32900), .Z(n32905) );
  NANDN U33686 ( .A(n32903), .B(n32902), .Z(n32904) );
  AND U33687 ( .A(n32905), .B(n32904), .Z(n33038) );
  NANDN U33688 ( .A(n32907), .B(n32906), .Z(n32911) );
  NANDN U33689 ( .A(n32909), .B(n32908), .Z(n32910) );
  NAND U33690 ( .A(n32911), .B(n32910), .Z(n33037) );
  XNOR U33691 ( .A(n33038), .B(n33037), .Z(n33039) );
  NAND U33692 ( .A(b[0]), .B(a[236]), .Z(n32912) );
  XNOR U33693 ( .A(b[1]), .B(n32912), .Z(n32914) );
  NANDN U33694 ( .A(b[0]), .B(a[235]), .Z(n32913) );
  NAND U33695 ( .A(n32914), .B(n32913), .Z(n32986) );
  NAND U33696 ( .A(n194), .B(n32915), .Z(n32917) );
  XOR U33697 ( .A(b[29]), .B(a[208]), .Z(n33061) );
  NAND U33698 ( .A(n38456), .B(n33061), .Z(n32916) );
  AND U33699 ( .A(n32917), .B(n32916), .Z(n32984) );
  AND U33700 ( .A(b[31]), .B(a[204]), .Z(n32983) );
  XNOR U33701 ( .A(n32984), .B(n32983), .Z(n32985) );
  XNOR U33702 ( .A(n32986), .B(n32985), .Z(n33025) );
  NAND U33703 ( .A(n38185), .B(n32918), .Z(n32920) );
  XOR U33704 ( .A(b[23]), .B(a[214]), .Z(n33067) );
  NAND U33705 ( .A(n38132), .B(n33067), .Z(n32919) );
  AND U33706 ( .A(n32920), .B(n32919), .Z(n33058) );
  NAND U33707 ( .A(n184), .B(n32921), .Z(n32923) );
  XOR U33708 ( .A(b[7]), .B(a[230]), .Z(n33070) );
  NAND U33709 ( .A(n36592), .B(n33070), .Z(n32922) );
  AND U33710 ( .A(n32923), .B(n32922), .Z(n33056) );
  NAND U33711 ( .A(n38289), .B(n32924), .Z(n32926) );
  XOR U33712 ( .A(b[25]), .B(a[212]), .Z(n33073) );
  NAND U33713 ( .A(n38247), .B(n33073), .Z(n32925) );
  NAND U33714 ( .A(n32926), .B(n32925), .Z(n33055) );
  XNOR U33715 ( .A(n33056), .B(n33055), .Z(n33057) );
  XOR U33716 ( .A(n33058), .B(n33057), .Z(n33026) );
  XNOR U33717 ( .A(n33025), .B(n33026), .Z(n33027) );
  NAND U33718 ( .A(n187), .B(n32927), .Z(n32929) );
  XOR U33719 ( .A(b[13]), .B(a[224]), .Z(n33076) );
  NAND U33720 ( .A(n37295), .B(n33076), .Z(n32928) );
  AND U33721 ( .A(n32929), .B(n32928), .Z(n33020) );
  NAND U33722 ( .A(n186), .B(n32930), .Z(n32932) );
  XOR U33723 ( .A(b[11]), .B(a[226]), .Z(n33079) );
  NAND U33724 ( .A(n37097), .B(n33079), .Z(n32931) );
  NAND U33725 ( .A(n32932), .B(n32931), .Z(n33019) );
  XNOR U33726 ( .A(n33020), .B(n33019), .Z(n33021) );
  NAND U33727 ( .A(n188), .B(n32933), .Z(n32935) );
  XOR U33728 ( .A(b[15]), .B(a[222]), .Z(n33082) );
  NAND U33729 ( .A(n37382), .B(n33082), .Z(n32934) );
  AND U33730 ( .A(n32935), .B(n32934), .Z(n33016) );
  NAND U33731 ( .A(n38064), .B(n32936), .Z(n32938) );
  XOR U33732 ( .A(b[21]), .B(a[216]), .Z(n33085) );
  NAND U33733 ( .A(n37993), .B(n33085), .Z(n32937) );
  AND U33734 ( .A(n32938), .B(n32937), .Z(n33014) );
  NAND U33735 ( .A(n185), .B(n32939), .Z(n32941) );
  XOR U33736 ( .A(b[9]), .B(a[228]), .Z(n33088) );
  NAND U33737 ( .A(n36805), .B(n33088), .Z(n32940) );
  NAND U33738 ( .A(n32941), .B(n32940), .Z(n33013) );
  XNOR U33739 ( .A(n33014), .B(n33013), .Z(n33015) );
  XOR U33740 ( .A(n33016), .B(n33015), .Z(n33022) );
  XOR U33741 ( .A(n33021), .B(n33022), .Z(n33028) );
  XOR U33742 ( .A(n33027), .B(n33028), .Z(n33040) );
  XNOR U33743 ( .A(n33039), .B(n33040), .Z(n32971) );
  XNOR U33744 ( .A(n32972), .B(n32971), .Z(n32973) );
  XOR U33745 ( .A(n32974), .B(n32973), .Z(n33092) );
  XNOR U33746 ( .A(n33091), .B(n33092), .Z(n33093) );
  XNOR U33747 ( .A(n33094), .B(n33093), .Z(n32967) );
  XOR U33748 ( .A(n32968), .B(n32967), .Z(n32960) );
  NANDN U33749 ( .A(n32943), .B(n32942), .Z(n32947) );
  OR U33750 ( .A(n32945), .B(n32944), .Z(n32946) );
  AND U33751 ( .A(n32947), .B(n32946), .Z(n32959) );
  XNOR U33752 ( .A(n32960), .B(n32959), .Z(n32961) );
  XNOR U33753 ( .A(n32962), .B(n32961), .Z(n32953) );
  XNOR U33754 ( .A(n32954), .B(n32953), .Z(n32955) );
  XNOR U33755 ( .A(n32956), .B(n32955), .Z(n33097) );
  XNOR U33756 ( .A(sreg[460]), .B(n33097), .Z(n33099) );
  NANDN U33757 ( .A(sreg[459]), .B(n32948), .Z(n32952) );
  NAND U33758 ( .A(n32950), .B(n32949), .Z(n32951) );
  NAND U33759 ( .A(n32952), .B(n32951), .Z(n33098) );
  XNOR U33760 ( .A(n33099), .B(n33098), .Z(c[460]) );
  NANDN U33761 ( .A(n32954), .B(n32953), .Z(n32958) );
  NANDN U33762 ( .A(n32956), .B(n32955), .Z(n32957) );
  AND U33763 ( .A(n32958), .B(n32957), .Z(n33105) );
  NANDN U33764 ( .A(n32960), .B(n32959), .Z(n32964) );
  NANDN U33765 ( .A(n32962), .B(n32961), .Z(n32963) );
  AND U33766 ( .A(n32964), .B(n32963), .Z(n33103) );
  NANDN U33767 ( .A(n32966), .B(n32965), .Z(n32970) );
  NAND U33768 ( .A(n32968), .B(n32967), .Z(n32969) );
  AND U33769 ( .A(n32970), .B(n32969), .Z(n33110) );
  NANDN U33770 ( .A(n32972), .B(n32971), .Z(n32976) );
  NANDN U33771 ( .A(n32974), .B(n32973), .Z(n32975) );
  AND U33772 ( .A(n32976), .B(n32975), .Z(n33115) );
  NANDN U33773 ( .A(n32978), .B(n32977), .Z(n32982) );
  NAND U33774 ( .A(n32980), .B(n32979), .Z(n32981) );
  AND U33775 ( .A(n32982), .B(n32981), .Z(n33114) );
  XNOR U33776 ( .A(n33115), .B(n33114), .Z(n33117) );
  NANDN U33777 ( .A(n32984), .B(n32983), .Z(n32988) );
  NANDN U33778 ( .A(n32986), .B(n32985), .Z(n32987) );
  AND U33779 ( .A(n32988), .B(n32987), .Z(n33194) );
  NAND U33780 ( .A(n38385), .B(n32989), .Z(n32991) );
  XOR U33781 ( .A(b[27]), .B(a[211]), .Z(n33138) );
  NAND U33782 ( .A(n38343), .B(n33138), .Z(n32990) );
  AND U33783 ( .A(n32991), .B(n32990), .Z(n33201) );
  NAND U33784 ( .A(n183), .B(n32992), .Z(n32994) );
  XOR U33785 ( .A(a[233]), .B(b[5]), .Z(n33141) );
  NAND U33786 ( .A(n36296), .B(n33141), .Z(n32993) );
  AND U33787 ( .A(n32994), .B(n32993), .Z(n33199) );
  NAND U33788 ( .A(n190), .B(n32995), .Z(n32997) );
  XOR U33789 ( .A(b[19]), .B(a[219]), .Z(n33144) );
  NAND U33790 ( .A(n37821), .B(n33144), .Z(n32996) );
  NAND U33791 ( .A(n32997), .B(n32996), .Z(n33198) );
  XNOR U33792 ( .A(n33199), .B(n33198), .Z(n33200) );
  XNOR U33793 ( .A(n33201), .B(n33200), .Z(n33192) );
  NAND U33794 ( .A(n38470), .B(n32998), .Z(n33000) );
  XOR U33795 ( .A(b[31]), .B(a[207]), .Z(n33147) );
  NAND U33796 ( .A(n38453), .B(n33147), .Z(n32999) );
  AND U33797 ( .A(n33000), .B(n32999), .Z(n33159) );
  NAND U33798 ( .A(n181), .B(n33001), .Z(n33003) );
  XOR U33799 ( .A(a[235]), .B(b[3]), .Z(n33150) );
  NAND U33800 ( .A(n182), .B(n33150), .Z(n33002) );
  AND U33801 ( .A(n33003), .B(n33002), .Z(n33157) );
  NAND U33802 ( .A(n189), .B(n33004), .Z(n33006) );
  XOR U33803 ( .A(b[17]), .B(a[221]), .Z(n33153) );
  NAND U33804 ( .A(n37652), .B(n33153), .Z(n33005) );
  NAND U33805 ( .A(n33006), .B(n33005), .Z(n33156) );
  XNOR U33806 ( .A(n33157), .B(n33156), .Z(n33158) );
  XOR U33807 ( .A(n33159), .B(n33158), .Z(n33193) );
  XOR U33808 ( .A(n33192), .B(n33193), .Z(n33195) );
  XOR U33809 ( .A(n33194), .B(n33195), .Z(n33127) );
  NANDN U33810 ( .A(n33008), .B(n33007), .Z(n33012) );
  NANDN U33811 ( .A(n33010), .B(n33009), .Z(n33011) );
  AND U33812 ( .A(n33012), .B(n33011), .Z(n33180) );
  NANDN U33813 ( .A(n33014), .B(n33013), .Z(n33018) );
  NANDN U33814 ( .A(n33016), .B(n33015), .Z(n33017) );
  NAND U33815 ( .A(n33018), .B(n33017), .Z(n33181) );
  XNOR U33816 ( .A(n33180), .B(n33181), .Z(n33182) );
  NANDN U33817 ( .A(n33020), .B(n33019), .Z(n33024) );
  NANDN U33818 ( .A(n33022), .B(n33021), .Z(n33023) );
  NAND U33819 ( .A(n33024), .B(n33023), .Z(n33183) );
  XNOR U33820 ( .A(n33182), .B(n33183), .Z(n33126) );
  XNOR U33821 ( .A(n33127), .B(n33126), .Z(n33129) );
  NANDN U33822 ( .A(n33026), .B(n33025), .Z(n33030) );
  NANDN U33823 ( .A(n33028), .B(n33027), .Z(n33029) );
  AND U33824 ( .A(n33030), .B(n33029), .Z(n33128) );
  XOR U33825 ( .A(n33129), .B(n33128), .Z(n33243) );
  NANDN U33826 ( .A(n33032), .B(n33031), .Z(n33036) );
  NANDN U33827 ( .A(n33034), .B(n33033), .Z(n33035) );
  AND U33828 ( .A(n33036), .B(n33035), .Z(n33240) );
  NANDN U33829 ( .A(n33038), .B(n33037), .Z(n33042) );
  NANDN U33830 ( .A(n33040), .B(n33039), .Z(n33041) );
  AND U33831 ( .A(n33042), .B(n33041), .Z(n33123) );
  NANDN U33832 ( .A(n33044), .B(n33043), .Z(n33048) );
  OR U33833 ( .A(n33046), .B(n33045), .Z(n33047) );
  AND U33834 ( .A(n33048), .B(n33047), .Z(n33121) );
  NANDN U33835 ( .A(n33050), .B(n33049), .Z(n33054) );
  NANDN U33836 ( .A(n33052), .B(n33051), .Z(n33053) );
  AND U33837 ( .A(n33054), .B(n33053), .Z(n33187) );
  NANDN U33838 ( .A(n33056), .B(n33055), .Z(n33060) );
  NANDN U33839 ( .A(n33058), .B(n33057), .Z(n33059) );
  NAND U33840 ( .A(n33060), .B(n33059), .Z(n33186) );
  XNOR U33841 ( .A(n33187), .B(n33186), .Z(n33188) );
  NAND U33842 ( .A(n194), .B(n33061), .Z(n33063) );
  XOR U33843 ( .A(b[29]), .B(a[209]), .Z(n33213) );
  NAND U33844 ( .A(n38456), .B(n33213), .Z(n33062) );
  AND U33845 ( .A(n33063), .B(n33062), .Z(n33133) );
  AND U33846 ( .A(b[31]), .B(a[205]), .Z(n33132) );
  XNOR U33847 ( .A(n33133), .B(n33132), .Z(n33134) );
  NAND U33848 ( .A(b[0]), .B(a[237]), .Z(n33064) );
  XNOR U33849 ( .A(b[1]), .B(n33064), .Z(n33066) );
  NANDN U33850 ( .A(b[0]), .B(a[236]), .Z(n33065) );
  NAND U33851 ( .A(n33066), .B(n33065), .Z(n33135) );
  XNOR U33852 ( .A(n33134), .B(n33135), .Z(n33174) );
  NAND U33853 ( .A(n38185), .B(n33067), .Z(n33069) );
  XOR U33854 ( .A(b[23]), .B(a[215]), .Z(n33216) );
  NAND U33855 ( .A(n38132), .B(n33216), .Z(n33068) );
  AND U33856 ( .A(n33069), .B(n33068), .Z(n33207) );
  NAND U33857 ( .A(n184), .B(n33070), .Z(n33072) );
  XOR U33858 ( .A(b[7]), .B(a[231]), .Z(n33219) );
  NAND U33859 ( .A(n36592), .B(n33219), .Z(n33071) );
  AND U33860 ( .A(n33072), .B(n33071), .Z(n33205) );
  NAND U33861 ( .A(n38289), .B(n33073), .Z(n33075) );
  XOR U33862 ( .A(b[25]), .B(a[213]), .Z(n33222) );
  NAND U33863 ( .A(n38247), .B(n33222), .Z(n33074) );
  NAND U33864 ( .A(n33075), .B(n33074), .Z(n33204) );
  XNOR U33865 ( .A(n33205), .B(n33204), .Z(n33206) );
  XOR U33866 ( .A(n33207), .B(n33206), .Z(n33175) );
  XNOR U33867 ( .A(n33174), .B(n33175), .Z(n33176) );
  NAND U33868 ( .A(n187), .B(n33076), .Z(n33078) );
  XOR U33869 ( .A(b[13]), .B(a[225]), .Z(n33225) );
  NAND U33870 ( .A(n37295), .B(n33225), .Z(n33077) );
  AND U33871 ( .A(n33078), .B(n33077), .Z(n33169) );
  NAND U33872 ( .A(n186), .B(n33079), .Z(n33081) );
  XOR U33873 ( .A(b[11]), .B(a[227]), .Z(n33228) );
  NAND U33874 ( .A(n37097), .B(n33228), .Z(n33080) );
  NAND U33875 ( .A(n33081), .B(n33080), .Z(n33168) );
  XNOR U33876 ( .A(n33169), .B(n33168), .Z(n33170) );
  NAND U33877 ( .A(n188), .B(n33082), .Z(n33084) );
  XOR U33878 ( .A(b[15]), .B(a[223]), .Z(n33231) );
  NAND U33879 ( .A(n37382), .B(n33231), .Z(n33083) );
  AND U33880 ( .A(n33084), .B(n33083), .Z(n33165) );
  NAND U33881 ( .A(n38064), .B(n33085), .Z(n33087) );
  XOR U33882 ( .A(b[21]), .B(a[217]), .Z(n33234) );
  NAND U33883 ( .A(n37993), .B(n33234), .Z(n33086) );
  AND U33884 ( .A(n33087), .B(n33086), .Z(n33163) );
  NAND U33885 ( .A(n185), .B(n33088), .Z(n33090) );
  XOR U33886 ( .A(b[9]), .B(a[229]), .Z(n33237) );
  NAND U33887 ( .A(n36805), .B(n33237), .Z(n33089) );
  NAND U33888 ( .A(n33090), .B(n33089), .Z(n33162) );
  XNOR U33889 ( .A(n33163), .B(n33162), .Z(n33164) );
  XOR U33890 ( .A(n33165), .B(n33164), .Z(n33171) );
  XOR U33891 ( .A(n33170), .B(n33171), .Z(n33177) );
  XOR U33892 ( .A(n33176), .B(n33177), .Z(n33189) );
  XNOR U33893 ( .A(n33188), .B(n33189), .Z(n33120) );
  XNOR U33894 ( .A(n33121), .B(n33120), .Z(n33122) );
  XOR U33895 ( .A(n33123), .B(n33122), .Z(n33241) );
  XNOR U33896 ( .A(n33240), .B(n33241), .Z(n33242) );
  XNOR U33897 ( .A(n33243), .B(n33242), .Z(n33116) );
  XOR U33898 ( .A(n33117), .B(n33116), .Z(n33109) );
  NANDN U33899 ( .A(n33092), .B(n33091), .Z(n33096) );
  NANDN U33900 ( .A(n33094), .B(n33093), .Z(n33095) );
  AND U33901 ( .A(n33096), .B(n33095), .Z(n33108) );
  XOR U33902 ( .A(n33109), .B(n33108), .Z(n33111) );
  XNOR U33903 ( .A(n33110), .B(n33111), .Z(n33102) );
  XNOR U33904 ( .A(n33103), .B(n33102), .Z(n33104) );
  XNOR U33905 ( .A(n33105), .B(n33104), .Z(n33246) );
  XNOR U33906 ( .A(sreg[461]), .B(n33246), .Z(n33248) );
  NANDN U33907 ( .A(sreg[460]), .B(n33097), .Z(n33101) );
  NAND U33908 ( .A(n33099), .B(n33098), .Z(n33100) );
  NAND U33909 ( .A(n33101), .B(n33100), .Z(n33247) );
  XNOR U33910 ( .A(n33248), .B(n33247), .Z(c[461]) );
  NANDN U33911 ( .A(n33103), .B(n33102), .Z(n33107) );
  NANDN U33912 ( .A(n33105), .B(n33104), .Z(n33106) );
  AND U33913 ( .A(n33107), .B(n33106), .Z(n33254) );
  NANDN U33914 ( .A(n33109), .B(n33108), .Z(n33113) );
  NANDN U33915 ( .A(n33111), .B(n33110), .Z(n33112) );
  AND U33916 ( .A(n33113), .B(n33112), .Z(n33252) );
  NANDN U33917 ( .A(n33115), .B(n33114), .Z(n33119) );
  NAND U33918 ( .A(n33117), .B(n33116), .Z(n33118) );
  AND U33919 ( .A(n33119), .B(n33118), .Z(n33259) );
  NANDN U33920 ( .A(n33121), .B(n33120), .Z(n33125) );
  NANDN U33921 ( .A(n33123), .B(n33122), .Z(n33124) );
  AND U33922 ( .A(n33125), .B(n33124), .Z(n33264) );
  NANDN U33923 ( .A(n33127), .B(n33126), .Z(n33131) );
  NAND U33924 ( .A(n33129), .B(n33128), .Z(n33130) );
  AND U33925 ( .A(n33131), .B(n33130), .Z(n33263) );
  XNOR U33926 ( .A(n33264), .B(n33263), .Z(n33266) );
  NANDN U33927 ( .A(n33133), .B(n33132), .Z(n33137) );
  NANDN U33928 ( .A(n33135), .B(n33134), .Z(n33136) );
  AND U33929 ( .A(n33137), .B(n33136), .Z(n33343) );
  NAND U33930 ( .A(n38385), .B(n33138), .Z(n33140) );
  XOR U33931 ( .A(b[27]), .B(a[212]), .Z(n33287) );
  NAND U33932 ( .A(n38343), .B(n33287), .Z(n33139) );
  AND U33933 ( .A(n33140), .B(n33139), .Z(n33350) );
  NAND U33934 ( .A(n183), .B(n33141), .Z(n33143) );
  XOR U33935 ( .A(a[234]), .B(b[5]), .Z(n33290) );
  NAND U33936 ( .A(n36296), .B(n33290), .Z(n33142) );
  AND U33937 ( .A(n33143), .B(n33142), .Z(n33348) );
  NAND U33938 ( .A(n190), .B(n33144), .Z(n33146) );
  XOR U33939 ( .A(b[19]), .B(a[220]), .Z(n33293) );
  NAND U33940 ( .A(n37821), .B(n33293), .Z(n33145) );
  NAND U33941 ( .A(n33146), .B(n33145), .Z(n33347) );
  XNOR U33942 ( .A(n33348), .B(n33347), .Z(n33349) );
  XNOR U33943 ( .A(n33350), .B(n33349), .Z(n33341) );
  NAND U33944 ( .A(n38470), .B(n33147), .Z(n33149) );
  XOR U33945 ( .A(b[31]), .B(a[208]), .Z(n33296) );
  NAND U33946 ( .A(n38453), .B(n33296), .Z(n33148) );
  AND U33947 ( .A(n33149), .B(n33148), .Z(n33308) );
  NAND U33948 ( .A(n181), .B(n33150), .Z(n33152) );
  XOR U33949 ( .A(a[236]), .B(b[3]), .Z(n33299) );
  NAND U33950 ( .A(n182), .B(n33299), .Z(n33151) );
  AND U33951 ( .A(n33152), .B(n33151), .Z(n33306) );
  NAND U33952 ( .A(n189), .B(n33153), .Z(n33155) );
  XOR U33953 ( .A(b[17]), .B(a[222]), .Z(n33302) );
  NAND U33954 ( .A(n37652), .B(n33302), .Z(n33154) );
  NAND U33955 ( .A(n33155), .B(n33154), .Z(n33305) );
  XNOR U33956 ( .A(n33306), .B(n33305), .Z(n33307) );
  XOR U33957 ( .A(n33308), .B(n33307), .Z(n33342) );
  XOR U33958 ( .A(n33341), .B(n33342), .Z(n33344) );
  XOR U33959 ( .A(n33343), .B(n33344), .Z(n33276) );
  NANDN U33960 ( .A(n33157), .B(n33156), .Z(n33161) );
  NANDN U33961 ( .A(n33159), .B(n33158), .Z(n33160) );
  AND U33962 ( .A(n33161), .B(n33160), .Z(n33329) );
  NANDN U33963 ( .A(n33163), .B(n33162), .Z(n33167) );
  NANDN U33964 ( .A(n33165), .B(n33164), .Z(n33166) );
  NAND U33965 ( .A(n33167), .B(n33166), .Z(n33330) );
  XNOR U33966 ( .A(n33329), .B(n33330), .Z(n33331) );
  NANDN U33967 ( .A(n33169), .B(n33168), .Z(n33173) );
  NANDN U33968 ( .A(n33171), .B(n33170), .Z(n33172) );
  NAND U33969 ( .A(n33173), .B(n33172), .Z(n33332) );
  XNOR U33970 ( .A(n33331), .B(n33332), .Z(n33275) );
  XNOR U33971 ( .A(n33276), .B(n33275), .Z(n33278) );
  NANDN U33972 ( .A(n33175), .B(n33174), .Z(n33179) );
  NANDN U33973 ( .A(n33177), .B(n33176), .Z(n33178) );
  AND U33974 ( .A(n33179), .B(n33178), .Z(n33277) );
  XOR U33975 ( .A(n33278), .B(n33277), .Z(n33392) );
  NANDN U33976 ( .A(n33181), .B(n33180), .Z(n33185) );
  NANDN U33977 ( .A(n33183), .B(n33182), .Z(n33184) );
  AND U33978 ( .A(n33185), .B(n33184), .Z(n33389) );
  NANDN U33979 ( .A(n33187), .B(n33186), .Z(n33191) );
  NANDN U33980 ( .A(n33189), .B(n33188), .Z(n33190) );
  AND U33981 ( .A(n33191), .B(n33190), .Z(n33272) );
  NANDN U33982 ( .A(n33193), .B(n33192), .Z(n33197) );
  OR U33983 ( .A(n33195), .B(n33194), .Z(n33196) );
  AND U33984 ( .A(n33197), .B(n33196), .Z(n33270) );
  NANDN U33985 ( .A(n33199), .B(n33198), .Z(n33203) );
  NANDN U33986 ( .A(n33201), .B(n33200), .Z(n33202) );
  AND U33987 ( .A(n33203), .B(n33202), .Z(n33336) );
  NANDN U33988 ( .A(n33205), .B(n33204), .Z(n33209) );
  NANDN U33989 ( .A(n33207), .B(n33206), .Z(n33208) );
  NAND U33990 ( .A(n33209), .B(n33208), .Z(n33335) );
  XNOR U33991 ( .A(n33336), .B(n33335), .Z(n33337) );
  NAND U33992 ( .A(b[0]), .B(a[238]), .Z(n33210) );
  XNOR U33993 ( .A(b[1]), .B(n33210), .Z(n33212) );
  NANDN U33994 ( .A(b[0]), .B(a[237]), .Z(n33211) );
  NAND U33995 ( .A(n33212), .B(n33211), .Z(n33284) );
  NAND U33996 ( .A(n194), .B(n33213), .Z(n33215) );
  XOR U33997 ( .A(b[29]), .B(a[210]), .Z(n33362) );
  NAND U33998 ( .A(n38456), .B(n33362), .Z(n33214) );
  AND U33999 ( .A(n33215), .B(n33214), .Z(n33282) );
  AND U34000 ( .A(b[31]), .B(a[206]), .Z(n33281) );
  XNOR U34001 ( .A(n33282), .B(n33281), .Z(n33283) );
  XNOR U34002 ( .A(n33284), .B(n33283), .Z(n33323) );
  NAND U34003 ( .A(n38185), .B(n33216), .Z(n33218) );
  XOR U34004 ( .A(b[23]), .B(a[216]), .Z(n33365) );
  NAND U34005 ( .A(n38132), .B(n33365), .Z(n33217) );
  AND U34006 ( .A(n33218), .B(n33217), .Z(n33356) );
  NAND U34007 ( .A(n184), .B(n33219), .Z(n33221) );
  XOR U34008 ( .A(a[232]), .B(b[7]), .Z(n33368) );
  NAND U34009 ( .A(n36592), .B(n33368), .Z(n33220) );
  AND U34010 ( .A(n33221), .B(n33220), .Z(n33354) );
  NAND U34011 ( .A(n38289), .B(n33222), .Z(n33224) );
  XOR U34012 ( .A(b[25]), .B(a[214]), .Z(n33371) );
  NAND U34013 ( .A(n38247), .B(n33371), .Z(n33223) );
  NAND U34014 ( .A(n33224), .B(n33223), .Z(n33353) );
  XNOR U34015 ( .A(n33354), .B(n33353), .Z(n33355) );
  XOR U34016 ( .A(n33356), .B(n33355), .Z(n33324) );
  XNOR U34017 ( .A(n33323), .B(n33324), .Z(n33325) );
  NAND U34018 ( .A(n187), .B(n33225), .Z(n33227) );
  XOR U34019 ( .A(b[13]), .B(a[226]), .Z(n33374) );
  NAND U34020 ( .A(n37295), .B(n33374), .Z(n33226) );
  AND U34021 ( .A(n33227), .B(n33226), .Z(n33318) );
  NAND U34022 ( .A(n186), .B(n33228), .Z(n33230) );
  XOR U34023 ( .A(b[11]), .B(a[228]), .Z(n33377) );
  NAND U34024 ( .A(n37097), .B(n33377), .Z(n33229) );
  NAND U34025 ( .A(n33230), .B(n33229), .Z(n33317) );
  XNOR U34026 ( .A(n33318), .B(n33317), .Z(n33319) );
  NAND U34027 ( .A(n188), .B(n33231), .Z(n33233) );
  XOR U34028 ( .A(b[15]), .B(a[224]), .Z(n33380) );
  NAND U34029 ( .A(n37382), .B(n33380), .Z(n33232) );
  AND U34030 ( .A(n33233), .B(n33232), .Z(n33314) );
  NAND U34031 ( .A(n38064), .B(n33234), .Z(n33236) );
  XOR U34032 ( .A(b[21]), .B(a[218]), .Z(n33383) );
  NAND U34033 ( .A(n37993), .B(n33383), .Z(n33235) );
  AND U34034 ( .A(n33236), .B(n33235), .Z(n33312) );
  NAND U34035 ( .A(n185), .B(n33237), .Z(n33239) );
  XOR U34036 ( .A(b[9]), .B(a[230]), .Z(n33386) );
  NAND U34037 ( .A(n36805), .B(n33386), .Z(n33238) );
  NAND U34038 ( .A(n33239), .B(n33238), .Z(n33311) );
  XNOR U34039 ( .A(n33312), .B(n33311), .Z(n33313) );
  XOR U34040 ( .A(n33314), .B(n33313), .Z(n33320) );
  XOR U34041 ( .A(n33319), .B(n33320), .Z(n33326) );
  XOR U34042 ( .A(n33325), .B(n33326), .Z(n33338) );
  XNOR U34043 ( .A(n33337), .B(n33338), .Z(n33269) );
  XNOR U34044 ( .A(n33270), .B(n33269), .Z(n33271) );
  XOR U34045 ( .A(n33272), .B(n33271), .Z(n33390) );
  XNOR U34046 ( .A(n33389), .B(n33390), .Z(n33391) );
  XNOR U34047 ( .A(n33392), .B(n33391), .Z(n33265) );
  XOR U34048 ( .A(n33266), .B(n33265), .Z(n33258) );
  NANDN U34049 ( .A(n33241), .B(n33240), .Z(n33245) );
  NANDN U34050 ( .A(n33243), .B(n33242), .Z(n33244) );
  AND U34051 ( .A(n33245), .B(n33244), .Z(n33257) );
  XOR U34052 ( .A(n33258), .B(n33257), .Z(n33260) );
  XNOR U34053 ( .A(n33259), .B(n33260), .Z(n33251) );
  XNOR U34054 ( .A(n33252), .B(n33251), .Z(n33253) );
  XNOR U34055 ( .A(n33254), .B(n33253), .Z(n33395) );
  XNOR U34056 ( .A(sreg[462]), .B(n33395), .Z(n33397) );
  NANDN U34057 ( .A(sreg[461]), .B(n33246), .Z(n33250) );
  NAND U34058 ( .A(n33248), .B(n33247), .Z(n33249) );
  NAND U34059 ( .A(n33250), .B(n33249), .Z(n33396) );
  XNOR U34060 ( .A(n33397), .B(n33396), .Z(c[462]) );
  NANDN U34061 ( .A(n33252), .B(n33251), .Z(n33256) );
  NANDN U34062 ( .A(n33254), .B(n33253), .Z(n33255) );
  AND U34063 ( .A(n33256), .B(n33255), .Z(n33403) );
  NANDN U34064 ( .A(n33258), .B(n33257), .Z(n33262) );
  NANDN U34065 ( .A(n33260), .B(n33259), .Z(n33261) );
  AND U34066 ( .A(n33262), .B(n33261), .Z(n33401) );
  NANDN U34067 ( .A(n33264), .B(n33263), .Z(n33268) );
  NAND U34068 ( .A(n33266), .B(n33265), .Z(n33267) );
  AND U34069 ( .A(n33268), .B(n33267), .Z(n33408) );
  NANDN U34070 ( .A(n33270), .B(n33269), .Z(n33274) );
  NANDN U34071 ( .A(n33272), .B(n33271), .Z(n33273) );
  AND U34072 ( .A(n33274), .B(n33273), .Z(n33413) );
  NANDN U34073 ( .A(n33276), .B(n33275), .Z(n33280) );
  NAND U34074 ( .A(n33278), .B(n33277), .Z(n33279) );
  AND U34075 ( .A(n33280), .B(n33279), .Z(n33412) );
  XNOR U34076 ( .A(n33413), .B(n33412), .Z(n33415) );
  NANDN U34077 ( .A(n33282), .B(n33281), .Z(n33286) );
  NANDN U34078 ( .A(n33284), .B(n33283), .Z(n33285) );
  AND U34079 ( .A(n33286), .B(n33285), .Z(n33492) );
  NAND U34080 ( .A(n38385), .B(n33287), .Z(n33289) );
  XOR U34081 ( .A(b[27]), .B(a[213]), .Z(n33436) );
  NAND U34082 ( .A(n38343), .B(n33436), .Z(n33288) );
  AND U34083 ( .A(n33289), .B(n33288), .Z(n33499) );
  NAND U34084 ( .A(n183), .B(n33290), .Z(n33292) );
  XOR U34085 ( .A(a[235]), .B(b[5]), .Z(n33439) );
  NAND U34086 ( .A(n36296), .B(n33439), .Z(n33291) );
  AND U34087 ( .A(n33292), .B(n33291), .Z(n33497) );
  NAND U34088 ( .A(n190), .B(n33293), .Z(n33295) );
  XOR U34089 ( .A(b[19]), .B(a[221]), .Z(n33442) );
  NAND U34090 ( .A(n37821), .B(n33442), .Z(n33294) );
  NAND U34091 ( .A(n33295), .B(n33294), .Z(n33496) );
  XNOR U34092 ( .A(n33497), .B(n33496), .Z(n33498) );
  XNOR U34093 ( .A(n33499), .B(n33498), .Z(n33490) );
  NAND U34094 ( .A(n38470), .B(n33296), .Z(n33298) );
  XOR U34095 ( .A(b[31]), .B(a[209]), .Z(n33445) );
  NAND U34096 ( .A(n38453), .B(n33445), .Z(n33297) );
  AND U34097 ( .A(n33298), .B(n33297), .Z(n33457) );
  NAND U34098 ( .A(n181), .B(n33299), .Z(n33301) );
  XOR U34099 ( .A(a[237]), .B(b[3]), .Z(n33448) );
  NAND U34100 ( .A(n182), .B(n33448), .Z(n33300) );
  AND U34101 ( .A(n33301), .B(n33300), .Z(n33455) );
  NAND U34102 ( .A(n189), .B(n33302), .Z(n33304) );
  XOR U34103 ( .A(b[17]), .B(a[223]), .Z(n33451) );
  NAND U34104 ( .A(n37652), .B(n33451), .Z(n33303) );
  NAND U34105 ( .A(n33304), .B(n33303), .Z(n33454) );
  XNOR U34106 ( .A(n33455), .B(n33454), .Z(n33456) );
  XOR U34107 ( .A(n33457), .B(n33456), .Z(n33491) );
  XOR U34108 ( .A(n33490), .B(n33491), .Z(n33493) );
  XOR U34109 ( .A(n33492), .B(n33493), .Z(n33425) );
  NANDN U34110 ( .A(n33306), .B(n33305), .Z(n33310) );
  NANDN U34111 ( .A(n33308), .B(n33307), .Z(n33309) );
  AND U34112 ( .A(n33310), .B(n33309), .Z(n33478) );
  NANDN U34113 ( .A(n33312), .B(n33311), .Z(n33316) );
  NANDN U34114 ( .A(n33314), .B(n33313), .Z(n33315) );
  NAND U34115 ( .A(n33316), .B(n33315), .Z(n33479) );
  XNOR U34116 ( .A(n33478), .B(n33479), .Z(n33480) );
  NANDN U34117 ( .A(n33318), .B(n33317), .Z(n33322) );
  NANDN U34118 ( .A(n33320), .B(n33319), .Z(n33321) );
  NAND U34119 ( .A(n33322), .B(n33321), .Z(n33481) );
  XNOR U34120 ( .A(n33480), .B(n33481), .Z(n33424) );
  XNOR U34121 ( .A(n33425), .B(n33424), .Z(n33427) );
  NANDN U34122 ( .A(n33324), .B(n33323), .Z(n33328) );
  NANDN U34123 ( .A(n33326), .B(n33325), .Z(n33327) );
  AND U34124 ( .A(n33328), .B(n33327), .Z(n33426) );
  XOR U34125 ( .A(n33427), .B(n33426), .Z(n33541) );
  NANDN U34126 ( .A(n33330), .B(n33329), .Z(n33334) );
  NANDN U34127 ( .A(n33332), .B(n33331), .Z(n33333) );
  AND U34128 ( .A(n33334), .B(n33333), .Z(n33538) );
  NANDN U34129 ( .A(n33336), .B(n33335), .Z(n33340) );
  NANDN U34130 ( .A(n33338), .B(n33337), .Z(n33339) );
  AND U34131 ( .A(n33340), .B(n33339), .Z(n33421) );
  NANDN U34132 ( .A(n33342), .B(n33341), .Z(n33346) );
  OR U34133 ( .A(n33344), .B(n33343), .Z(n33345) );
  AND U34134 ( .A(n33346), .B(n33345), .Z(n33419) );
  NANDN U34135 ( .A(n33348), .B(n33347), .Z(n33352) );
  NANDN U34136 ( .A(n33350), .B(n33349), .Z(n33351) );
  AND U34137 ( .A(n33352), .B(n33351), .Z(n33485) );
  NANDN U34138 ( .A(n33354), .B(n33353), .Z(n33358) );
  NANDN U34139 ( .A(n33356), .B(n33355), .Z(n33357) );
  NAND U34140 ( .A(n33358), .B(n33357), .Z(n33484) );
  XNOR U34141 ( .A(n33485), .B(n33484), .Z(n33486) );
  NAND U34142 ( .A(b[0]), .B(a[239]), .Z(n33359) );
  XNOR U34143 ( .A(b[1]), .B(n33359), .Z(n33361) );
  NANDN U34144 ( .A(b[0]), .B(a[238]), .Z(n33360) );
  NAND U34145 ( .A(n33361), .B(n33360), .Z(n33433) );
  NAND U34146 ( .A(n194), .B(n33362), .Z(n33364) );
  XOR U34147 ( .A(b[29]), .B(a[211]), .Z(n33511) );
  NAND U34148 ( .A(n38456), .B(n33511), .Z(n33363) );
  AND U34149 ( .A(n33364), .B(n33363), .Z(n33431) );
  AND U34150 ( .A(b[31]), .B(a[207]), .Z(n33430) );
  XNOR U34151 ( .A(n33431), .B(n33430), .Z(n33432) );
  XNOR U34152 ( .A(n33433), .B(n33432), .Z(n33472) );
  NAND U34153 ( .A(n38185), .B(n33365), .Z(n33367) );
  XOR U34154 ( .A(b[23]), .B(a[217]), .Z(n33514) );
  NAND U34155 ( .A(n38132), .B(n33514), .Z(n33366) );
  AND U34156 ( .A(n33367), .B(n33366), .Z(n33505) );
  NAND U34157 ( .A(n184), .B(n33368), .Z(n33370) );
  XOR U34158 ( .A(b[7]), .B(a[233]), .Z(n33517) );
  NAND U34159 ( .A(n36592), .B(n33517), .Z(n33369) );
  AND U34160 ( .A(n33370), .B(n33369), .Z(n33503) );
  NAND U34161 ( .A(n38289), .B(n33371), .Z(n33373) );
  XOR U34162 ( .A(b[25]), .B(a[215]), .Z(n33520) );
  NAND U34163 ( .A(n38247), .B(n33520), .Z(n33372) );
  NAND U34164 ( .A(n33373), .B(n33372), .Z(n33502) );
  XNOR U34165 ( .A(n33503), .B(n33502), .Z(n33504) );
  XOR U34166 ( .A(n33505), .B(n33504), .Z(n33473) );
  XNOR U34167 ( .A(n33472), .B(n33473), .Z(n33474) );
  NAND U34168 ( .A(n187), .B(n33374), .Z(n33376) );
  XOR U34169 ( .A(b[13]), .B(a[227]), .Z(n33523) );
  NAND U34170 ( .A(n37295), .B(n33523), .Z(n33375) );
  AND U34171 ( .A(n33376), .B(n33375), .Z(n33467) );
  NAND U34172 ( .A(n186), .B(n33377), .Z(n33379) );
  XOR U34173 ( .A(b[11]), .B(a[229]), .Z(n33526) );
  NAND U34174 ( .A(n37097), .B(n33526), .Z(n33378) );
  NAND U34175 ( .A(n33379), .B(n33378), .Z(n33466) );
  XNOR U34176 ( .A(n33467), .B(n33466), .Z(n33468) );
  NAND U34177 ( .A(n188), .B(n33380), .Z(n33382) );
  XOR U34178 ( .A(b[15]), .B(a[225]), .Z(n33529) );
  NAND U34179 ( .A(n37382), .B(n33529), .Z(n33381) );
  AND U34180 ( .A(n33382), .B(n33381), .Z(n33463) );
  NAND U34181 ( .A(n38064), .B(n33383), .Z(n33385) );
  XOR U34182 ( .A(b[21]), .B(a[219]), .Z(n33532) );
  NAND U34183 ( .A(n37993), .B(n33532), .Z(n33384) );
  AND U34184 ( .A(n33385), .B(n33384), .Z(n33461) );
  NAND U34185 ( .A(n185), .B(n33386), .Z(n33388) );
  XOR U34186 ( .A(b[9]), .B(a[231]), .Z(n33535) );
  NAND U34187 ( .A(n36805), .B(n33535), .Z(n33387) );
  NAND U34188 ( .A(n33388), .B(n33387), .Z(n33460) );
  XNOR U34189 ( .A(n33461), .B(n33460), .Z(n33462) );
  XOR U34190 ( .A(n33463), .B(n33462), .Z(n33469) );
  XOR U34191 ( .A(n33468), .B(n33469), .Z(n33475) );
  XOR U34192 ( .A(n33474), .B(n33475), .Z(n33487) );
  XNOR U34193 ( .A(n33486), .B(n33487), .Z(n33418) );
  XNOR U34194 ( .A(n33419), .B(n33418), .Z(n33420) );
  XOR U34195 ( .A(n33421), .B(n33420), .Z(n33539) );
  XNOR U34196 ( .A(n33538), .B(n33539), .Z(n33540) );
  XNOR U34197 ( .A(n33541), .B(n33540), .Z(n33414) );
  XOR U34198 ( .A(n33415), .B(n33414), .Z(n33407) );
  NANDN U34199 ( .A(n33390), .B(n33389), .Z(n33394) );
  NANDN U34200 ( .A(n33392), .B(n33391), .Z(n33393) );
  AND U34201 ( .A(n33394), .B(n33393), .Z(n33406) );
  XOR U34202 ( .A(n33407), .B(n33406), .Z(n33409) );
  XNOR U34203 ( .A(n33408), .B(n33409), .Z(n33400) );
  XNOR U34204 ( .A(n33401), .B(n33400), .Z(n33402) );
  XNOR U34205 ( .A(n33403), .B(n33402), .Z(n33544) );
  XNOR U34206 ( .A(sreg[463]), .B(n33544), .Z(n33546) );
  NANDN U34207 ( .A(sreg[462]), .B(n33395), .Z(n33399) );
  NAND U34208 ( .A(n33397), .B(n33396), .Z(n33398) );
  NAND U34209 ( .A(n33399), .B(n33398), .Z(n33545) );
  XNOR U34210 ( .A(n33546), .B(n33545), .Z(c[463]) );
  NANDN U34211 ( .A(n33401), .B(n33400), .Z(n33405) );
  NANDN U34212 ( .A(n33403), .B(n33402), .Z(n33404) );
  AND U34213 ( .A(n33405), .B(n33404), .Z(n33552) );
  NANDN U34214 ( .A(n33407), .B(n33406), .Z(n33411) );
  NANDN U34215 ( .A(n33409), .B(n33408), .Z(n33410) );
  AND U34216 ( .A(n33411), .B(n33410), .Z(n33550) );
  NANDN U34217 ( .A(n33413), .B(n33412), .Z(n33417) );
  NAND U34218 ( .A(n33415), .B(n33414), .Z(n33416) );
  AND U34219 ( .A(n33417), .B(n33416), .Z(n33557) );
  NANDN U34220 ( .A(n33419), .B(n33418), .Z(n33423) );
  NANDN U34221 ( .A(n33421), .B(n33420), .Z(n33422) );
  AND U34222 ( .A(n33423), .B(n33422), .Z(n33562) );
  NANDN U34223 ( .A(n33425), .B(n33424), .Z(n33429) );
  NAND U34224 ( .A(n33427), .B(n33426), .Z(n33428) );
  AND U34225 ( .A(n33429), .B(n33428), .Z(n33561) );
  XNOR U34226 ( .A(n33562), .B(n33561), .Z(n33564) );
  NANDN U34227 ( .A(n33431), .B(n33430), .Z(n33435) );
  NANDN U34228 ( .A(n33433), .B(n33432), .Z(n33434) );
  AND U34229 ( .A(n33435), .B(n33434), .Z(n33641) );
  NAND U34230 ( .A(n38385), .B(n33436), .Z(n33438) );
  XOR U34231 ( .A(b[27]), .B(a[214]), .Z(n33585) );
  NAND U34232 ( .A(n38343), .B(n33585), .Z(n33437) );
  AND U34233 ( .A(n33438), .B(n33437), .Z(n33648) );
  NAND U34234 ( .A(n183), .B(n33439), .Z(n33441) );
  XOR U34235 ( .A(a[236]), .B(b[5]), .Z(n33588) );
  NAND U34236 ( .A(n36296), .B(n33588), .Z(n33440) );
  AND U34237 ( .A(n33441), .B(n33440), .Z(n33646) );
  NAND U34238 ( .A(n190), .B(n33442), .Z(n33444) );
  XOR U34239 ( .A(b[19]), .B(a[222]), .Z(n33591) );
  NAND U34240 ( .A(n37821), .B(n33591), .Z(n33443) );
  NAND U34241 ( .A(n33444), .B(n33443), .Z(n33645) );
  XNOR U34242 ( .A(n33646), .B(n33645), .Z(n33647) );
  XNOR U34243 ( .A(n33648), .B(n33647), .Z(n33639) );
  NAND U34244 ( .A(n38470), .B(n33445), .Z(n33447) );
  XOR U34245 ( .A(b[31]), .B(a[210]), .Z(n33594) );
  NAND U34246 ( .A(n38453), .B(n33594), .Z(n33446) );
  AND U34247 ( .A(n33447), .B(n33446), .Z(n33606) );
  NAND U34248 ( .A(n181), .B(n33448), .Z(n33450) );
  XOR U34249 ( .A(a[238]), .B(b[3]), .Z(n33597) );
  NAND U34250 ( .A(n182), .B(n33597), .Z(n33449) );
  AND U34251 ( .A(n33450), .B(n33449), .Z(n33604) );
  NAND U34252 ( .A(n189), .B(n33451), .Z(n33453) );
  XOR U34253 ( .A(b[17]), .B(a[224]), .Z(n33600) );
  NAND U34254 ( .A(n37652), .B(n33600), .Z(n33452) );
  NAND U34255 ( .A(n33453), .B(n33452), .Z(n33603) );
  XNOR U34256 ( .A(n33604), .B(n33603), .Z(n33605) );
  XOR U34257 ( .A(n33606), .B(n33605), .Z(n33640) );
  XOR U34258 ( .A(n33639), .B(n33640), .Z(n33642) );
  XOR U34259 ( .A(n33641), .B(n33642), .Z(n33574) );
  NANDN U34260 ( .A(n33455), .B(n33454), .Z(n33459) );
  NANDN U34261 ( .A(n33457), .B(n33456), .Z(n33458) );
  AND U34262 ( .A(n33459), .B(n33458), .Z(n33627) );
  NANDN U34263 ( .A(n33461), .B(n33460), .Z(n33465) );
  NANDN U34264 ( .A(n33463), .B(n33462), .Z(n33464) );
  NAND U34265 ( .A(n33465), .B(n33464), .Z(n33628) );
  XNOR U34266 ( .A(n33627), .B(n33628), .Z(n33629) );
  NANDN U34267 ( .A(n33467), .B(n33466), .Z(n33471) );
  NANDN U34268 ( .A(n33469), .B(n33468), .Z(n33470) );
  NAND U34269 ( .A(n33471), .B(n33470), .Z(n33630) );
  XNOR U34270 ( .A(n33629), .B(n33630), .Z(n33573) );
  XNOR U34271 ( .A(n33574), .B(n33573), .Z(n33576) );
  NANDN U34272 ( .A(n33473), .B(n33472), .Z(n33477) );
  NANDN U34273 ( .A(n33475), .B(n33474), .Z(n33476) );
  AND U34274 ( .A(n33477), .B(n33476), .Z(n33575) );
  XOR U34275 ( .A(n33576), .B(n33575), .Z(n33690) );
  NANDN U34276 ( .A(n33479), .B(n33478), .Z(n33483) );
  NANDN U34277 ( .A(n33481), .B(n33480), .Z(n33482) );
  AND U34278 ( .A(n33483), .B(n33482), .Z(n33687) );
  NANDN U34279 ( .A(n33485), .B(n33484), .Z(n33489) );
  NANDN U34280 ( .A(n33487), .B(n33486), .Z(n33488) );
  AND U34281 ( .A(n33489), .B(n33488), .Z(n33570) );
  NANDN U34282 ( .A(n33491), .B(n33490), .Z(n33495) );
  OR U34283 ( .A(n33493), .B(n33492), .Z(n33494) );
  AND U34284 ( .A(n33495), .B(n33494), .Z(n33568) );
  NANDN U34285 ( .A(n33497), .B(n33496), .Z(n33501) );
  NANDN U34286 ( .A(n33499), .B(n33498), .Z(n33500) );
  AND U34287 ( .A(n33501), .B(n33500), .Z(n33634) );
  NANDN U34288 ( .A(n33503), .B(n33502), .Z(n33507) );
  NANDN U34289 ( .A(n33505), .B(n33504), .Z(n33506) );
  NAND U34290 ( .A(n33507), .B(n33506), .Z(n33633) );
  XNOR U34291 ( .A(n33634), .B(n33633), .Z(n33635) );
  NAND U34292 ( .A(b[0]), .B(a[240]), .Z(n33508) );
  XNOR U34293 ( .A(b[1]), .B(n33508), .Z(n33510) );
  NANDN U34294 ( .A(b[0]), .B(a[239]), .Z(n33509) );
  NAND U34295 ( .A(n33510), .B(n33509), .Z(n33582) );
  NAND U34296 ( .A(n194), .B(n33511), .Z(n33513) );
  XOR U34297 ( .A(b[29]), .B(a[212]), .Z(n33660) );
  NAND U34298 ( .A(n38456), .B(n33660), .Z(n33512) );
  AND U34299 ( .A(n33513), .B(n33512), .Z(n33580) );
  AND U34300 ( .A(b[31]), .B(a[208]), .Z(n33579) );
  XNOR U34301 ( .A(n33580), .B(n33579), .Z(n33581) );
  XNOR U34302 ( .A(n33582), .B(n33581), .Z(n33621) );
  NAND U34303 ( .A(n38185), .B(n33514), .Z(n33516) );
  XOR U34304 ( .A(b[23]), .B(a[218]), .Z(n33663) );
  NAND U34305 ( .A(n38132), .B(n33663), .Z(n33515) );
  AND U34306 ( .A(n33516), .B(n33515), .Z(n33654) );
  NAND U34307 ( .A(n184), .B(n33517), .Z(n33519) );
  XOR U34308 ( .A(a[234]), .B(b[7]), .Z(n33666) );
  NAND U34309 ( .A(n36592), .B(n33666), .Z(n33518) );
  AND U34310 ( .A(n33519), .B(n33518), .Z(n33652) );
  NAND U34311 ( .A(n38289), .B(n33520), .Z(n33522) );
  XOR U34312 ( .A(b[25]), .B(a[216]), .Z(n33669) );
  NAND U34313 ( .A(n38247), .B(n33669), .Z(n33521) );
  NAND U34314 ( .A(n33522), .B(n33521), .Z(n33651) );
  XNOR U34315 ( .A(n33652), .B(n33651), .Z(n33653) );
  XOR U34316 ( .A(n33654), .B(n33653), .Z(n33622) );
  XNOR U34317 ( .A(n33621), .B(n33622), .Z(n33623) );
  NAND U34318 ( .A(n187), .B(n33523), .Z(n33525) );
  XOR U34319 ( .A(b[13]), .B(a[228]), .Z(n33672) );
  NAND U34320 ( .A(n37295), .B(n33672), .Z(n33524) );
  AND U34321 ( .A(n33525), .B(n33524), .Z(n33616) );
  NAND U34322 ( .A(n186), .B(n33526), .Z(n33528) );
  XOR U34323 ( .A(b[11]), .B(a[230]), .Z(n33675) );
  NAND U34324 ( .A(n37097), .B(n33675), .Z(n33527) );
  NAND U34325 ( .A(n33528), .B(n33527), .Z(n33615) );
  XNOR U34326 ( .A(n33616), .B(n33615), .Z(n33617) );
  NAND U34327 ( .A(n188), .B(n33529), .Z(n33531) );
  XOR U34328 ( .A(b[15]), .B(a[226]), .Z(n33678) );
  NAND U34329 ( .A(n37382), .B(n33678), .Z(n33530) );
  AND U34330 ( .A(n33531), .B(n33530), .Z(n33612) );
  NAND U34331 ( .A(n38064), .B(n33532), .Z(n33534) );
  XOR U34332 ( .A(b[21]), .B(a[220]), .Z(n33681) );
  NAND U34333 ( .A(n37993), .B(n33681), .Z(n33533) );
  AND U34334 ( .A(n33534), .B(n33533), .Z(n33610) );
  NAND U34335 ( .A(n185), .B(n33535), .Z(n33537) );
  XOR U34336 ( .A(b[9]), .B(a[232]), .Z(n33684) );
  NAND U34337 ( .A(n36805), .B(n33684), .Z(n33536) );
  NAND U34338 ( .A(n33537), .B(n33536), .Z(n33609) );
  XNOR U34339 ( .A(n33610), .B(n33609), .Z(n33611) );
  XOR U34340 ( .A(n33612), .B(n33611), .Z(n33618) );
  XOR U34341 ( .A(n33617), .B(n33618), .Z(n33624) );
  XOR U34342 ( .A(n33623), .B(n33624), .Z(n33636) );
  XNOR U34343 ( .A(n33635), .B(n33636), .Z(n33567) );
  XNOR U34344 ( .A(n33568), .B(n33567), .Z(n33569) );
  XOR U34345 ( .A(n33570), .B(n33569), .Z(n33688) );
  XNOR U34346 ( .A(n33687), .B(n33688), .Z(n33689) );
  XNOR U34347 ( .A(n33690), .B(n33689), .Z(n33563) );
  XOR U34348 ( .A(n33564), .B(n33563), .Z(n33556) );
  NANDN U34349 ( .A(n33539), .B(n33538), .Z(n33543) );
  NANDN U34350 ( .A(n33541), .B(n33540), .Z(n33542) );
  AND U34351 ( .A(n33543), .B(n33542), .Z(n33555) );
  XOR U34352 ( .A(n33556), .B(n33555), .Z(n33558) );
  XNOR U34353 ( .A(n33557), .B(n33558), .Z(n33549) );
  XNOR U34354 ( .A(n33550), .B(n33549), .Z(n33551) );
  XNOR U34355 ( .A(n33552), .B(n33551), .Z(n33693) );
  XNOR U34356 ( .A(sreg[464]), .B(n33693), .Z(n33695) );
  NANDN U34357 ( .A(sreg[463]), .B(n33544), .Z(n33548) );
  NAND U34358 ( .A(n33546), .B(n33545), .Z(n33547) );
  NAND U34359 ( .A(n33548), .B(n33547), .Z(n33694) );
  XNOR U34360 ( .A(n33695), .B(n33694), .Z(c[464]) );
  NANDN U34361 ( .A(n33550), .B(n33549), .Z(n33554) );
  NANDN U34362 ( .A(n33552), .B(n33551), .Z(n33553) );
  AND U34363 ( .A(n33554), .B(n33553), .Z(n33701) );
  NANDN U34364 ( .A(n33556), .B(n33555), .Z(n33560) );
  NANDN U34365 ( .A(n33558), .B(n33557), .Z(n33559) );
  AND U34366 ( .A(n33560), .B(n33559), .Z(n33699) );
  NANDN U34367 ( .A(n33562), .B(n33561), .Z(n33566) );
  NAND U34368 ( .A(n33564), .B(n33563), .Z(n33565) );
  AND U34369 ( .A(n33566), .B(n33565), .Z(n33706) );
  NANDN U34370 ( .A(n33568), .B(n33567), .Z(n33572) );
  NANDN U34371 ( .A(n33570), .B(n33569), .Z(n33571) );
  AND U34372 ( .A(n33572), .B(n33571), .Z(n33711) );
  NANDN U34373 ( .A(n33574), .B(n33573), .Z(n33578) );
  NAND U34374 ( .A(n33576), .B(n33575), .Z(n33577) );
  AND U34375 ( .A(n33578), .B(n33577), .Z(n33710) );
  XNOR U34376 ( .A(n33711), .B(n33710), .Z(n33713) );
  NANDN U34377 ( .A(n33580), .B(n33579), .Z(n33584) );
  NANDN U34378 ( .A(n33582), .B(n33581), .Z(n33583) );
  AND U34379 ( .A(n33584), .B(n33583), .Z(n33790) );
  NAND U34380 ( .A(n38385), .B(n33585), .Z(n33587) );
  XOR U34381 ( .A(b[27]), .B(a[215]), .Z(n33734) );
  NAND U34382 ( .A(n38343), .B(n33734), .Z(n33586) );
  AND U34383 ( .A(n33587), .B(n33586), .Z(n33797) );
  NAND U34384 ( .A(n183), .B(n33588), .Z(n33590) );
  XOR U34385 ( .A(a[237]), .B(b[5]), .Z(n33737) );
  NAND U34386 ( .A(n36296), .B(n33737), .Z(n33589) );
  AND U34387 ( .A(n33590), .B(n33589), .Z(n33795) );
  NAND U34388 ( .A(n190), .B(n33591), .Z(n33593) );
  XOR U34389 ( .A(b[19]), .B(a[223]), .Z(n33740) );
  NAND U34390 ( .A(n37821), .B(n33740), .Z(n33592) );
  NAND U34391 ( .A(n33593), .B(n33592), .Z(n33794) );
  XNOR U34392 ( .A(n33795), .B(n33794), .Z(n33796) );
  XNOR U34393 ( .A(n33797), .B(n33796), .Z(n33788) );
  NAND U34394 ( .A(n38470), .B(n33594), .Z(n33596) );
  XOR U34395 ( .A(b[31]), .B(a[211]), .Z(n33743) );
  NAND U34396 ( .A(n38453), .B(n33743), .Z(n33595) );
  AND U34397 ( .A(n33596), .B(n33595), .Z(n33755) );
  NAND U34398 ( .A(n181), .B(n33597), .Z(n33599) );
  XOR U34399 ( .A(a[239]), .B(b[3]), .Z(n33746) );
  NAND U34400 ( .A(n182), .B(n33746), .Z(n33598) );
  AND U34401 ( .A(n33599), .B(n33598), .Z(n33753) );
  NAND U34402 ( .A(n189), .B(n33600), .Z(n33602) );
  XOR U34403 ( .A(b[17]), .B(a[225]), .Z(n33749) );
  NAND U34404 ( .A(n37652), .B(n33749), .Z(n33601) );
  NAND U34405 ( .A(n33602), .B(n33601), .Z(n33752) );
  XNOR U34406 ( .A(n33753), .B(n33752), .Z(n33754) );
  XOR U34407 ( .A(n33755), .B(n33754), .Z(n33789) );
  XOR U34408 ( .A(n33788), .B(n33789), .Z(n33791) );
  XOR U34409 ( .A(n33790), .B(n33791), .Z(n33723) );
  NANDN U34410 ( .A(n33604), .B(n33603), .Z(n33608) );
  NANDN U34411 ( .A(n33606), .B(n33605), .Z(n33607) );
  AND U34412 ( .A(n33608), .B(n33607), .Z(n33776) );
  NANDN U34413 ( .A(n33610), .B(n33609), .Z(n33614) );
  NANDN U34414 ( .A(n33612), .B(n33611), .Z(n33613) );
  NAND U34415 ( .A(n33614), .B(n33613), .Z(n33777) );
  XNOR U34416 ( .A(n33776), .B(n33777), .Z(n33778) );
  NANDN U34417 ( .A(n33616), .B(n33615), .Z(n33620) );
  NANDN U34418 ( .A(n33618), .B(n33617), .Z(n33619) );
  NAND U34419 ( .A(n33620), .B(n33619), .Z(n33779) );
  XNOR U34420 ( .A(n33778), .B(n33779), .Z(n33722) );
  XNOR U34421 ( .A(n33723), .B(n33722), .Z(n33725) );
  NANDN U34422 ( .A(n33622), .B(n33621), .Z(n33626) );
  NANDN U34423 ( .A(n33624), .B(n33623), .Z(n33625) );
  AND U34424 ( .A(n33626), .B(n33625), .Z(n33724) );
  XOR U34425 ( .A(n33725), .B(n33724), .Z(n33839) );
  NANDN U34426 ( .A(n33628), .B(n33627), .Z(n33632) );
  NANDN U34427 ( .A(n33630), .B(n33629), .Z(n33631) );
  AND U34428 ( .A(n33632), .B(n33631), .Z(n33836) );
  NANDN U34429 ( .A(n33634), .B(n33633), .Z(n33638) );
  NANDN U34430 ( .A(n33636), .B(n33635), .Z(n33637) );
  AND U34431 ( .A(n33638), .B(n33637), .Z(n33719) );
  NANDN U34432 ( .A(n33640), .B(n33639), .Z(n33644) );
  OR U34433 ( .A(n33642), .B(n33641), .Z(n33643) );
  AND U34434 ( .A(n33644), .B(n33643), .Z(n33717) );
  NANDN U34435 ( .A(n33646), .B(n33645), .Z(n33650) );
  NANDN U34436 ( .A(n33648), .B(n33647), .Z(n33649) );
  AND U34437 ( .A(n33650), .B(n33649), .Z(n33783) );
  NANDN U34438 ( .A(n33652), .B(n33651), .Z(n33656) );
  NANDN U34439 ( .A(n33654), .B(n33653), .Z(n33655) );
  NAND U34440 ( .A(n33656), .B(n33655), .Z(n33782) );
  XNOR U34441 ( .A(n33783), .B(n33782), .Z(n33784) );
  NAND U34442 ( .A(b[0]), .B(a[241]), .Z(n33657) );
  XNOR U34443 ( .A(b[1]), .B(n33657), .Z(n33659) );
  NANDN U34444 ( .A(b[0]), .B(a[240]), .Z(n33658) );
  NAND U34445 ( .A(n33659), .B(n33658), .Z(n33731) );
  NAND U34446 ( .A(n194), .B(n33660), .Z(n33662) );
  XOR U34447 ( .A(b[29]), .B(a[213]), .Z(n33809) );
  NAND U34448 ( .A(n38456), .B(n33809), .Z(n33661) );
  AND U34449 ( .A(n33662), .B(n33661), .Z(n33729) );
  AND U34450 ( .A(b[31]), .B(a[209]), .Z(n33728) );
  XNOR U34451 ( .A(n33729), .B(n33728), .Z(n33730) );
  XNOR U34452 ( .A(n33731), .B(n33730), .Z(n33770) );
  NAND U34453 ( .A(n38185), .B(n33663), .Z(n33665) );
  XOR U34454 ( .A(b[23]), .B(a[219]), .Z(n33812) );
  NAND U34455 ( .A(n38132), .B(n33812), .Z(n33664) );
  AND U34456 ( .A(n33665), .B(n33664), .Z(n33803) );
  NAND U34457 ( .A(n184), .B(n33666), .Z(n33668) );
  XOR U34458 ( .A(a[235]), .B(b[7]), .Z(n33815) );
  NAND U34459 ( .A(n36592), .B(n33815), .Z(n33667) );
  AND U34460 ( .A(n33668), .B(n33667), .Z(n33801) );
  NAND U34461 ( .A(n38289), .B(n33669), .Z(n33671) );
  XOR U34462 ( .A(b[25]), .B(a[217]), .Z(n33818) );
  NAND U34463 ( .A(n38247), .B(n33818), .Z(n33670) );
  NAND U34464 ( .A(n33671), .B(n33670), .Z(n33800) );
  XNOR U34465 ( .A(n33801), .B(n33800), .Z(n33802) );
  XOR U34466 ( .A(n33803), .B(n33802), .Z(n33771) );
  XNOR U34467 ( .A(n33770), .B(n33771), .Z(n33772) );
  NAND U34468 ( .A(n187), .B(n33672), .Z(n33674) );
  XOR U34469 ( .A(b[13]), .B(a[229]), .Z(n33821) );
  NAND U34470 ( .A(n37295), .B(n33821), .Z(n33673) );
  AND U34471 ( .A(n33674), .B(n33673), .Z(n33765) );
  NAND U34472 ( .A(n186), .B(n33675), .Z(n33677) );
  XOR U34473 ( .A(b[11]), .B(a[231]), .Z(n33824) );
  NAND U34474 ( .A(n37097), .B(n33824), .Z(n33676) );
  NAND U34475 ( .A(n33677), .B(n33676), .Z(n33764) );
  XNOR U34476 ( .A(n33765), .B(n33764), .Z(n33766) );
  NAND U34477 ( .A(n188), .B(n33678), .Z(n33680) );
  XOR U34478 ( .A(b[15]), .B(a[227]), .Z(n33827) );
  NAND U34479 ( .A(n37382), .B(n33827), .Z(n33679) );
  AND U34480 ( .A(n33680), .B(n33679), .Z(n33761) );
  NAND U34481 ( .A(n38064), .B(n33681), .Z(n33683) );
  XOR U34482 ( .A(b[21]), .B(a[221]), .Z(n33830) );
  NAND U34483 ( .A(n37993), .B(n33830), .Z(n33682) );
  AND U34484 ( .A(n33683), .B(n33682), .Z(n33759) );
  NAND U34485 ( .A(n185), .B(n33684), .Z(n33686) );
  XOR U34486 ( .A(b[9]), .B(a[233]), .Z(n33833) );
  NAND U34487 ( .A(n36805), .B(n33833), .Z(n33685) );
  NAND U34488 ( .A(n33686), .B(n33685), .Z(n33758) );
  XNOR U34489 ( .A(n33759), .B(n33758), .Z(n33760) );
  XOR U34490 ( .A(n33761), .B(n33760), .Z(n33767) );
  XOR U34491 ( .A(n33766), .B(n33767), .Z(n33773) );
  XOR U34492 ( .A(n33772), .B(n33773), .Z(n33785) );
  XNOR U34493 ( .A(n33784), .B(n33785), .Z(n33716) );
  XNOR U34494 ( .A(n33717), .B(n33716), .Z(n33718) );
  XOR U34495 ( .A(n33719), .B(n33718), .Z(n33837) );
  XNOR U34496 ( .A(n33836), .B(n33837), .Z(n33838) );
  XNOR U34497 ( .A(n33839), .B(n33838), .Z(n33712) );
  XOR U34498 ( .A(n33713), .B(n33712), .Z(n33705) );
  NANDN U34499 ( .A(n33688), .B(n33687), .Z(n33692) );
  NANDN U34500 ( .A(n33690), .B(n33689), .Z(n33691) );
  AND U34501 ( .A(n33692), .B(n33691), .Z(n33704) );
  XOR U34502 ( .A(n33705), .B(n33704), .Z(n33707) );
  XNOR U34503 ( .A(n33706), .B(n33707), .Z(n33698) );
  XNOR U34504 ( .A(n33699), .B(n33698), .Z(n33700) );
  XNOR U34505 ( .A(n33701), .B(n33700), .Z(n33842) );
  XNOR U34506 ( .A(sreg[465]), .B(n33842), .Z(n33844) );
  NANDN U34507 ( .A(sreg[464]), .B(n33693), .Z(n33697) );
  NAND U34508 ( .A(n33695), .B(n33694), .Z(n33696) );
  NAND U34509 ( .A(n33697), .B(n33696), .Z(n33843) );
  XNOR U34510 ( .A(n33844), .B(n33843), .Z(c[465]) );
  NANDN U34511 ( .A(n33699), .B(n33698), .Z(n33703) );
  NANDN U34512 ( .A(n33701), .B(n33700), .Z(n33702) );
  AND U34513 ( .A(n33703), .B(n33702), .Z(n33850) );
  NANDN U34514 ( .A(n33705), .B(n33704), .Z(n33709) );
  NANDN U34515 ( .A(n33707), .B(n33706), .Z(n33708) );
  AND U34516 ( .A(n33709), .B(n33708), .Z(n33848) );
  NANDN U34517 ( .A(n33711), .B(n33710), .Z(n33715) );
  NAND U34518 ( .A(n33713), .B(n33712), .Z(n33714) );
  AND U34519 ( .A(n33715), .B(n33714), .Z(n33855) );
  NANDN U34520 ( .A(n33717), .B(n33716), .Z(n33721) );
  NANDN U34521 ( .A(n33719), .B(n33718), .Z(n33720) );
  AND U34522 ( .A(n33721), .B(n33720), .Z(n33860) );
  NANDN U34523 ( .A(n33723), .B(n33722), .Z(n33727) );
  NAND U34524 ( .A(n33725), .B(n33724), .Z(n33726) );
  AND U34525 ( .A(n33727), .B(n33726), .Z(n33859) );
  XNOR U34526 ( .A(n33860), .B(n33859), .Z(n33862) );
  NANDN U34527 ( .A(n33729), .B(n33728), .Z(n33733) );
  NANDN U34528 ( .A(n33731), .B(n33730), .Z(n33732) );
  AND U34529 ( .A(n33733), .B(n33732), .Z(n33937) );
  NAND U34530 ( .A(n38385), .B(n33734), .Z(n33736) );
  XOR U34531 ( .A(b[27]), .B(a[216]), .Z(n33883) );
  NAND U34532 ( .A(n38343), .B(n33883), .Z(n33735) );
  AND U34533 ( .A(n33736), .B(n33735), .Z(n33944) );
  NAND U34534 ( .A(n183), .B(n33737), .Z(n33739) );
  XOR U34535 ( .A(a[238]), .B(b[5]), .Z(n33886) );
  NAND U34536 ( .A(n36296), .B(n33886), .Z(n33738) );
  AND U34537 ( .A(n33739), .B(n33738), .Z(n33942) );
  NAND U34538 ( .A(n190), .B(n33740), .Z(n33742) );
  XOR U34539 ( .A(b[19]), .B(a[224]), .Z(n33889) );
  NAND U34540 ( .A(n37821), .B(n33889), .Z(n33741) );
  NAND U34541 ( .A(n33742), .B(n33741), .Z(n33941) );
  XNOR U34542 ( .A(n33942), .B(n33941), .Z(n33943) );
  XNOR U34543 ( .A(n33944), .B(n33943), .Z(n33935) );
  NAND U34544 ( .A(n38470), .B(n33743), .Z(n33745) );
  XOR U34545 ( .A(b[31]), .B(a[212]), .Z(n33892) );
  NAND U34546 ( .A(n38453), .B(n33892), .Z(n33744) );
  AND U34547 ( .A(n33745), .B(n33744), .Z(n33904) );
  NAND U34548 ( .A(n181), .B(n33746), .Z(n33748) );
  XOR U34549 ( .A(a[240]), .B(b[3]), .Z(n33895) );
  NAND U34550 ( .A(n182), .B(n33895), .Z(n33747) );
  AND U34551 ( .A(n33748), .B(n33747), .Z(n33902) );
  NAND U34552 ( .A(n189), .B(n33749), .Z(n33751) );
  XOR U34553 ( .A(b[17]), .B(a[226]), .Z(n33898) );
  NAND U34554 ( .A(n37652), .B(n33898), .Z(n33750) );
  NAND U34555 ( .A(n33751), .B(n33750), .Z(n33901) );
  XNOR U34556 ( .A(n33902), .B(n33901), .Z(n33903) );
  XOR U34557 ( .A(n33904), .B(n33903), .Z(n33936) );
  XOR U34558 ( .A(n33935), .B(n33936), .Z(n33938) );
  XOR U34559 ( .A(n33937), .B(n33938), .Z(n33872) );
  NANDN U34560 ( .A(n33753), .B(n33752), .Z(n33757) );
  NANDN U34561 ( .A(n33755), .B(n33754), .Z(n33756) );
  AND U34562 ( .A(n33757), .B(n33756), .Z(n33925) );
  NANDN U34563 ( .A(n33759), .B(n33758), .Z(n33763) );
  NANDN U34564 ( .A(n33761), .B(n33760), .Z(n33762) );
  NAND U34565 ( .A(n33763), .B(n33762), .Z(n33926) );
  XNOR U34566 ( .A(n33925), .B(n33926), .Z(n33927) );
  NANDN U34567 ( .A(n33765), .B(n33764), .Z(n33769) );
  NANDN U34568 ( .A(n33767), .B(n33766), .Z(n33768) );
  NAND U34569 ( .A(n33769), .B(n33768), .Z(n33928) );
  XNOR U34570 ( .A(n33927), .B(n33928), .Z(n33871) );
  XNOR U34571 ( .A(n33872), .B(n33871), .Z(n33874) );
  NANDN U34572 ( .A(n33771), .B(n33770), .Z(n33775) );
  NANDN U34573 ( .A(n33773), .B(n33772), .Z(n33774) );
  AND U34574 ( .A(n33775), .B(n33774), .Z(n33873) );
  XOR U34575 ( .A(n33874), .B(n33873), .Z(n33986) );
  NANDN U34576 ( .A(n33777), .B(n33776), .Z(n33781) );
  NANDN U34577 ( .A(n33779), .B(n33778), .Z(n33780) );
  AND U34578 ( .A(n33781), .B(n33780), .Z(n33983) );
  NANDN U34579 ( .A(n33783), .B(n33782), .Z(n33787) );
  NANDN U34580 ( .A(n33785), .B(n33784), .Z(n33786) );
  AND U34581 ( .A(n33787), .B(n33786), .Z(n33868) );
  NANDN U34582 ( .A(n33789), .B(n33788), .Z(n33793) );
  OR U34583 ( .A(n33791), .B(n33790), .Z(n33792) );
  AND U34584 ( .A(n33793), .B(n33792), .Z(n33866) );
  NANDN U34585 ( .A(n33795), .B(n33794), .Z(n33799) );
  NANDN U34586 ( .A(n33797), .B(n33796), .Z(n33798) );
  AND U34587 ( .A(n33799), .B(n33798), .Z(n33932) );
  NANDN U34588 ( .A(n33801), .B(n33800), .Z(n33805) );
  NANDN U34589 ( .A(n33803), .B(n33802), .Z(n33804) );
  NAND U34590 ( .A(n33805), .B(n33804), .Z(n33931) );
  XNOR U34591 ( .A(n33932), .B(n33931), .Z(n33934) );
  NAND U34592 ( .A(b[0]), .B(a[242]), .Z(n33806) );
  XNOR U34593 ( .A(b[1]), .B(n33806), .Z(n33808) );
  NANDN U34594 ( .A(b[0]), .B(a[241]), .Z(n33807) );
  NAND U34595 ( .A(n33808), .B(n33807), .Z(n33880) );
  NAND U34596 ( .A(n194), .B(n33809), .Z(n33811) );
  XOR U34597 ( .A(b[29]), .B(a[214]), .Z(n33956) );
  NAND U34598 ( .A(n38456), .B(n33956), .Z(n33810) );
  AND U34599 ( .A(n33811), .B(n33810), .Z(n33878) );
  AND U34600 ( .A(b[31]), .B(a[210]), .Z(n33877) );
  XNOR U34601 ( .A(n33878), .B(n33877), .Z(n33879) );
  XNOR U34602 ( .A(n33880), .B(n33879), .Z(n33920) );
  NAND U34603 ( .A(n38185), .B(n33812), .Z(n33814) );
  XOR U34604 ( .A(b[23]), .B(a[220]), .Z(n33959) );
  NAND U34605 ( .A(n38132), .B(n33959), .Z(n33813) );
  AND U34606 ( .A(n33814), .B(n33813), .Z(n33949) );
  NAND U34607 ( .A(n184), .B(n33815), .Z(n33817) );
  XOR U34608 ( .A(a[236]), .B(b[7]), .Z(n33962) );
  NAND U34609 ( .A(n36592), .B(n33962), .Z(n33816) );
  AND U34610 ( .A(n33817), .B(n33816), .Z(n33948) );
  NAND U34611 ( .A(n38289), .B(n33818), .Z(n33820) );
  XOR U34612 ( .A(b[25]), .B(a[218]), .Z(n33965) );
  NAND U34613 ( .A(n38247), .B(n33965), .Z(n33819) );
  NAND U34614 ( .A(n33820), .B(n33819), .Z(n33947) );
  XOR U34615 ( .A(n33948), .B(n33947), .Z(n33950) );
  XOR U34616 ( .A(n33949), .B(n33950), .Z(n33919) );
  XOR U34617 ( .A(n33920), .B(n33919), .Z(n33922) );
  NAND U34618 ( .A(n187), .B(n33821), .Z(n33823) );
  XOR U34619 ( .A(b[13]), .B(a[230]), .Z(n33968) );
  NAND U34620 ( .A(n37295), .B(n33968), .Z(n33822) );
  AND U34621 ( .A(n33823), .B(n33822), .Z(n33914) );
  NAND U34622 ( .A(n186), .B(n33824), .Z(n33826) );
  XOR U34623 ( .A(b[11]), .B(a[232]), .Z(n33971) );
  NAND U34624 ( .A(n37097), .B(n33971), .Z(n33825) );
  NAND U34625 ( .A(n33826), .B(n33825), .Z(n33913) );
  XNOR U34626 ( .A(n33914), .B(n33913), .Z(n33916) );
  NAND U34627 ( .A(n188), .B(n33827), .Z(n33829) );
  XOR U34628 ( .A(b[15]), .B(a[228]), .Z(n33974) );
  NAND U34629 ( .A(n37382), .B(n33974), .Z(n33828) );
  AND U34630 ( .A(n33829), .B(n33828), .Z(n33910) );
  NAND U34631 ( .A(n38064), .B(n33830), .Z(n33832) );
  XOR U34632 ( .A(b[21]), .B(a[222]), .Z(n33977) );
  NAND U34633 ( .A(n37993), .B(n33977), .Z(n33831) );
  AND U34634 ( .A(n33832), .B(n33831), .Z(n33908) );
  NAND U34635 ( .A(n185), .B(n33833), .Z(n33835) );
  XOR U34636 ( .A(b[9]), .B(a[234]), .Z(n33980) );
  NAND U34637 ( .A(n36805), .B(n33980), .Z(n33834) );
  NAND U34638 ( .A(n33835), .B(n33834), .Z(n33907) );
  XNOR U34639 ( .A(n33908), .B(n33907), .Z(n33909) );
  XNOR U34640 ( .A(n33910), .B(n33909), .Z(n33915) );
  XOR U34641 ( .A(n33916), .B(n33915), .Z(n33921) );
  XNOR U34642 ( .A(n33922), .B(n33921), .Z(n33933) );
  XNOR U34643 ( .A(n33934), .B(n33933), .Z(n33865) );
  XNOR U34644 ( .A(n33866), .B(n33865), .Z(n33867) );
  XOR U34645 ( .A(n33868), .B(n33867), .Z(n33984) );
  XNOR U34646 ( .A(n33983), .B(n33984), .Z(n33985) );
  XNOR U34647 ( .A(n33986), .B(n33985), .Z(n33861) );
  XOR U34648 ( .A(n33862), .B(n33861), .Z(n33854) );
  NANDN U34649 ( .A(n33837), .B(n33836), .Z(n33841) );
  NANDN U34650 ( .A(n33839), .B(n33838), .Z(n33840) );
  AND U34651 ( .A(n33841), .B(n33840), .Z(n33853) );
  XOR U34652 ( .A(n33854), .B(n33853), .Z(n33856) );
  XNOR U34653 ( .A(n33855), .B(n33856), .Z(n33847) );
  XNOR U34654 ( .A(n33848), .B(n33847), .Z(n33849) );
  XNOR U34655 ( .A(n33850), .B(n33849), .Z(n33989) );
  XNOR U34656 ( .A(sreg[466]), .B(n33989), .Z(n33991) );
  NANDN U34657 ( .A(sreg[465]), .B(n33842), .Z(n33846) );
  NAND U34658 ( .A(n33844), .B(n33843), .Z(n33845) );
  NAND U34659 ( .A(n33846), .B(n33845), .Z(n33990) );
  XNOR U34660 ( .A(n33991), .B(n33990), .Z(c[466]) );
  NANDN U34661 ( .A(n33848), .B(n33847), .Z(n33852) );
  NANDN U34662 ( .A(n33850), .B(n33849), .Z(n33851) );
  AND U34663 ( .A(n33852), .B(n33851), .Z(n33997) );
  NANDN U34664 ( .A(n33854), .B(n33853), .Z(n33858) );
  NANDN U34665 ( .A(n33856), .B(n33855), .Z(n33857) );
  AND U34666 ( .A(n33858), .B(n33857), .Z(n33995) );
  NANDN U34667 ( .A(n33860), .B(n33859), .Z(n33864) );
  NAND U34668 ( .A(n33862), .B(n33861), .Z(n33863) );
  AND U34669 ( .A(n33864), .B(n33863), .Z(n34002) );
  NANDN U34670 ( .A(n33866), .B(n33865), .Z(n33870) );
  NANDN U34671 ( .A(n33868), .B(n33867), .Z(n33869) );
  AND U34672 ( .A(n33870), .B(n33869), .Z(n34007) );
  NANDN U34673 ( .A(n33872), .B(n33871), .Z(n33876) );
  NAND U34674 ( .A(n33874), .B(n33873), .Z(n33875) );
  AND U34675 ( .A(n33876), .B(n33875), .Z(n34006) );
  XNOR U34676 ( .A(n34007), .B(n34006), .Z(n34009) );
  NANDN U34677 ( .A(n33878), .B(n33877), .Z(n33882) );
  NANDN U34678 ( .A(n33880), .B(n33879), .Z(n33881) );
  AND U34679 ( .A(n33882), .B(n33881), .Z(n34074) );
  NAND U34680 ( .A(n38385), .B(n33883), .Z(n33885) );
  XOR U34681 ( .A(b[27]), .B(a[217]), .Z(n34018) );
  NAND U34682 ( .A(n38343), .B(n34018), .Z(n33884) );
  AND U34683 ( .A(n33885), .B(n33884), .Z(n34081) );
  NAND U34684 ( .A(n183), .B(n33886), .Z(n33888) );
  XOR U34685 ( .A(a[239]), .B(b[5]), .Z(n34021) );
  NAND U34686 ( .A(n36296), .B(n34021), .Z(n33887) );
  AND U34687 ( .A(n33888), .B(n33887), .Z(n34079) );
  NAND U34688 ( .A(n190), .B(n33889), .Z(n33891) );
  XOR U34689 ( .A(b[19]), .B(a[225]), .Z(n34024) );
  NAND U34690 ( .A(n37821), .B(n34024), .Z(n33890) );
  NAND U34691 ( .A(n33891), .B(n33890), .Z(n34078) );
  XNOR U34692 ( .A(n34079), .B(n34078), .Z(n34080) );
  XNOR U34693 ( .A(n34081), .B(n34080), .Z(n34072) );
  NAND U34694 ( .A(n38470), .B(n33892), .Z(n33894) );
  XOR U34695 ( .A(b[31]), .B(a[213]), .Z(n34027) );
  NAND U34696 ( .A(n38453), .B(n34027), .Z(n33893) );
  AND U34697 ( .A(n33894), .B(n33893), .Z(n34039) );
  NAND U34698 ( .A(n181), .B(n33895), .Z(n33897) );
  XOR U34699 ( .A(a[241]), .B(b[3]), .Z(n34030) );
  NAND U34700 ( .A(n182), .B(n34030), .Z(n33896) );
  AND U34701 ( .A(n33897), .B(n33896), .Z(n34037) );
  NAND U34702 ( .A(n189), .B(n33898), .Z(n33900) );
  XOR U34703 ( .A(b[17]), .B(a[227]), .Z(n34033) );
  NAND U34704 ( .A(n37652), .B(n34033), .Z(n33899) );
  NAND U34705 ( .A(n33900), .B(n33899), .Z(n34036) );
  XNOR U34706 ( .A(n34037), .B(n34036), .Z(n34038) );
  XOR U34707 ( .A(n34039), .B(n34038), .Z(n34073) );
  XOR U34708 ( .A(n34072), .B(n34073), .Z(n34075) );
  XOR U34709 ( .A(n34074), .B(n34075), .Z(n34121) );
  NANDN U34710 ( .A(n33902), .B(n33901), .Z(n33906) );
  NANDN U34711 ( .A(n33904), .B(n33903), .Z(n33905) );
  AND U34712 ( .A(n33906), .B(n33905), .Z(n34060) );
  NANDN U34713 ( .A(n33908), .B(n33907), .Z(n33912) );
  NANDN U34714 ( .A(n33910), .B(n33909), .Z(n33911) );
  NAND U34715 ( .A(n33912), .B(n33911), .Z(n34061) );
  XNOR U34716 ( .A(n34060), .B(n34061), .Z(n34062) );
  NANDN U34717 ( .A(n33914), .B(n33913), .Z(n33918) );
  NAND U34718 ( .A(n33916), .B(n33915), .Z(n33917) );
  NAND U34719 ( .A(n33918), .B(n33917), .Z(n34063) );
  XNOR U34720 ( .A(n34062), .B(n34063), .Z(n34120) );
  XNOR U34721 ( .A(n34121), .B(n34120), .Z(n34123) );
  NAND U34722 ( .A(n33920), .B(n33919), .Z(n33924) );
  NAND U34723 ( .A(n33922), .B(n33921), .Z(n33923) );
  AND U34724 ( .A(n33924), .B(n33923), .Z(n34122) );
  XOR U34725 ( .A(n34123), .B(n34122), .Z(n34135) );
  NANDN U34726 ( .A(n33926), .B(n33925), .Z(n33930) );
  NANDN U34727 ( .A(n33928), .B(n33927), .Z(n33929) );
  AND U34728 ( .A(n33930), .B(n33929), .Z(n34132) );
  NANDN U34729 ( .A(n33936), .B(n33935), .Z(n33940) );
  OR U34730 ( .A(n33938), .B(n33937), .Z(n33939) );
  AND U34731 ( .A(n33940), .B(n33939), .Z(n34127) );
  NANDN U34732 ( .A(n33942), .B(n33941), .Z(n33946) );
  NANDN U34733 ( .A(n33944), .B(n33943), .Z(n33945) );
  AND U34734 ( .A(n33946), .B(n33945), .Z(n34067) );
  NANDN U34735 ( .A(n33948), .B(n33947), .Z(n33952) );
  OR U34736 ( .A(n33950), .B(n33949), .Z(n33951) );
  NAND U34737 ( .A(n33952), .B(n33951), .Z(n34066) );
  XNOR U34738 ( .A(n34067), .B(n34066), .Z(n34068) );
  NAND U34739 ( .A(b[0]), .B(a[243]), .Z(n33953) );
  XNOR U34740 ( .A(b[1]), .B(n33953), .Z(n33955) );
  NANDN U34741 ( .A(b[0]), .B(a[242]), .Z(n33954) );
  NAND U34742 ( .A(n33955), .B(n33954), .Z(n34015) );
  NAND U34743 ( .A(n194), .B(n33956), .Z(n33958) );
  XOR U34744 ( .A(b[29]), .B(a[215]), .Z(n34093) );
  NAND U34745 ( .A(n38456), .B(n34093), .Z(n33957) );
  AND U34746 ( .A(n33958), .B(n33957), .Z(n34013) );
  AND U34747 ( .A(b[31]), .B(a[211]), .Z(n34012) );
  XNOR U34748 ( .A(n34013), .B(n34012), .Z(n34014) );
  XNOR U34749 ( .A(n34015), .B(n34014), .Z(n34054) );
  NAND U34750 ( .A(n38185), .B(n33959), .Z(n33961) );
  XOR U34751 ( .A(b[23]), .B(a[221]), .Z(n34096) );
  NAND U34752 ( .A(n38132), .B(n34096), .Z(n33960) );
  AND U34753 ( .A(n33961), .B(n33960), .Z(n34087) );
  NAND U34754 ( .A(n184), .B(n33962), .Z(n33964) );
  XOR U34755 ( .A(a[237]), .B(b[7]), .Z(n34099) );
  NAND U34756 ( .A(n36592), .B(n34099), .Z(n33963) );
  AND U34757 ( .A(n33964), .B(n33963), .Z(n34085) );
  NAND U34758 ( .A(n38289), .B(n33965), .Z(n33967) );
  XOR U34759 ( .A(b[25]), .B(a[219]), .Z(n34102) );
  NAND U34760 ( .A(n38247), .B(n34102), .Z(n33966) );
  NAND U34761 ( .A(n33967), .B(n33966), .Z(n34084) );
  XNOR U34762 ( .A(n34085), .B(n34084), .Z(n34086) );
  XOR U34763 ( .A(n34087), .B(n34086), .Z(n34055) );
  XNOR U34764 ( .A(n34054), .B(n34055), .Z(n34056) );
  NAND U34765 ( .A(n187), .B(n33968), .Z(n33970) );
  XOR U34766 ( .A(b[13]), .B(a[231]), .Z(n34105) );
  NAND U34767 ( .A(n37295), .B(n34105), .Z(n33969) );
  AND U34768 ( .A(n33970), .B(n33969), .Z(n34049) );
  NAND U34769 ( .A(n186), .B(n33971), .Z(n33973) );
  XOR U34770 ( .A(b[11]), .B(a[233]), .Z(n34108) );
  NAND U34771 ( .A(n37097), .B(n34108), .Z(n33972) );
  NAND U34772 ( .A(n33973), .B(n33972), .Z(n34048) );
  XNOR U34773 ( .A(n34049), .B(n34048), .Z(n34050) );
  NAND U34774 ( .A(n188), .B(n33974), .Z(n33976) );
  XOR U34775 ( .A(b[15]), .B(a[229]), .Z(n34111) );
  NAND U34776 ( .A(n37382), .B(n34111), .Z(n33975) );
  AND U34777 ( .A(n33976), .B(n33975), .Z(n34045) );
  NAND U34778 ( .A(n38064), .B(n33977), .Z(n33979) );
  XOR U34779 ( .A(b[21]), .B(a[223]), .Z(n34114) );
  NAND U34780 ( .A(n37993), .B(n34114), .Z(n33978) );
  AND U34781 ( .A(n33979), .B(n33978), .Z(n34043) );
  NAND U34782 ( .A(n185), .B(n33980), .Z(n33982) );
  XOR U34783 ( .A(b[9]), .B(a[235]), .Z(n34117) );
  NAND U34784 ( .A(n36805), .B(n34117), .Z(n33981) );
  NAND U34785 ( .A(n33982), .B(n33981), .Z(n34042) );
  XNOR U34786 ( .A(n34043), .B(n34042), .Z(n34044) );
  XOR U34787 ( .A(n34045), .B(n34044), .Z(n34051) );
  XOR U34788 ( .A(n34050), .B(n34051), .Z(n34057) );
  XOR U34789 ( .A(n34056), .B(n34057), .Z(n34069) );
  XNOR U34790 ( .A(n34068), .B(n34069), .Z(n34126) );
  XNOR U34791 ( .A(n34127), .B(n34126), .Z(n34128) );
  XOR U34792 ( .A(n34129), .B(n34128), .Z(n34133) );
  XNOR U34793 ( .A(n34132), .B(n34133), .Z(n34134) );
  XNOR U34794 ( .A(n34135), .B(n34134), .Z(n34008) );
  XOR U34795 ( .A(n34009), .B(n34008), .Z(n34001) );
  NANDN U34796 ( .A(n33984), .B(n33983), .Z(n33988) );
  NANDN U34797 ( .A(n33986), .B(n33985), .Z(n33987) );
  AND U34798 ( .A(n33988), .B(n33987), .Z(n34000) );
  XOR U34799 ( .A(n34001), .B(n34000), .Z(n34003) );
  XNOR U34800 ( .A(n34002), .B(n34003), .Z(n33994) );
  XNOR U34801 ( .A(n33995), .B(n33994), .Z(n33996) );
  XNOR U34802 ( .A(n33997), .B(n33996), .Z(n34138) );
  XNOR U34803 ( .A(sreg[467]), .B(n34138), .Z(n34140) );
  NANDN U34804 ( .A(sreg[466]), .B(n33989), .Z(n33993) );
  NAND U34805 ( .A(n33991), .B(n33990), .Z(n33992) );
  NAND U34806 ( .A(n33993), .B(n33992), .Z(n34139) );
  XNOR U34807 ( .A(n34140), .B(n34139), .Z(c[467]) );
  NANDN U34808 ( .A(n33995), .B(n33994), .Z(n33999) );
  NANDN U34809 ( .A(n33997), .B(n33996), .Z(n33998) );
  AND U34810 ( .A(n33999), .B(n33998), .Z(n34146) );
  NANDN U34811 ( .A(n34001), .B(n34000), .Z(n34005) );
  NANDN U34812 ( .A(n34003), .B(n34002), .Z(n34004) );
  AND U34813 ( .A(n34005), .B(n34004), .Z(n34144) );
  NANDN U34814 ( .A(n34007), .B(n34006), .Z(n34011) );
  NAND U34815 ( .A(n34009), .B(n34008), .Z(n34010) );
  AND U34816 ( .A(n34011), .B(n34010), .Z(n34151) );
  NANDN U34817 ( .A(n34013), .B(n34012), .Z(n34017) );
  NANDN U34818 ( .A(n34015), .B(n34014), .Z(n34016) );
  AND U34819 ( .A(n34017), .B(n34016), .Z(n34235) );
  NAND U34820 ( .A(n38385), .B(n34018), .Z(n34020) );
  XOR U34821 ( .A(b[27]), .B(a[218]), .Z(n34179) );
  NAND U34822 ( .A(n38343), .B(n34179), .Z(n34019) );
  AND U34823 ( .A(n34020), .B(n34019), .Z(n34242) );
  NAND U34824 ( .A(n183), .B(n34021), .Z(n34023) );
  XOR U34825 ( .A(a[240]), .B(b[5]), .Z(n34182) );
  NAND U34826 ( .A(n36296), .B(n34182), .Z(n34022) );
  AND U34827 ( .A(n34023), .B(n34022), .Z(n34240) );
  NAND U34828 ( .A(n190), .B(n34024), .Z(n34026) );
  XOR U34829 ( .A(b[19]), .B(a[226]), .Z(n34185) );
  NAND U34830 ( .A(n37821), .B(n34185), .Z(n34025) );
  NAND U34831 ( .A(n34026), .B(n34025), .Z(n34239) );
  XNOR U34832 ( .A(n34240), .B(n34239), .Z(n34241) );
  XNOR U34833 ( .A(n34242), .B(n34241), .Z(n34233) );
  NAND U34834 ( .A(n38470), .B(n34027), .Z(n34029) );
  XOR U34835 ( .A(b[31]), .B(a[214]), .Z(n34188) );
  NAND U34836 ( .A(n38453), .B(n34188), .Z(n34028) );
  AND U34837 ( .A(n34029), .B(n34028), .Z(n34200) );
  NAND U34838 ( .A(n181), .B(n34030), .Z(n34032) );
  XOR U34839 ( .A(a[242]), .B(b[3]), .Z(n34191) );
  NAND U34840 ( .A(n182), .B(n34191), .Z(n34031) );
  AND U34841 ( .A(n34032), .B(n34031), .Z(n34198) );
  NAND U34842 ( .A(n189), .B(n34033), .Z(n34035) );
  XOR U34843 ( .A(b[17]), .B(a[228]), .Z(n34194) );
  NAND U34844 ( .A(n37652), .B(n34194), .Z(n34034) );
  NAND U34845 ( .A(n34035), .B(n34034), .Z(n34197) );
  XNOR U34846 ( .A(n34198), .B(n34197), .Z(n34199) );
  XOR U34847 ( .A(n34200), .B(n34199), .Z(n34234) );
  XOR U34848 ( .A(n34233), .B(n34234), .Z(n34236) );
  XOR U34849 ( .A(n34235), .B(n34236), .Z(n34168) );
  NANDN U34850 ( .A(n34037), .B(n34036), .Z(n34041) );
  NANDN U34851 ( .A(n34039), .B(n34038), .Z(n34040) );
  AND U34852 ( .A(n34041), .B(n34040), .Z(n34221) );
  NANDN U34853 ( .A(n34043), .B(n34042), .Z(n34047) );
  NANDN U34854 ( .A(n34045), .B(n34044), .Z(n34046) );
  NAND U34855 ( .A(n34047), .B(n34046), .Z(n34222) );
  XNOR U34856 ( .A(n34221), .B(n34222), .Z(n34223) );
  NANDN U34857 ( .A(n34049), .B(n34048), .Z(n34053) );
  NANDN U34858 ( .A(n34051), .B(n34050), .Z(n34052) );
  NAND U34859 ( .A(n34053), .B(n34052), .Z(n34224) );
  XNOR U34860 ( .A(n34223), .B(n34224), .Z(n34167) );
  XNOR U34861 ( .A(n34168), .B(n34167), .Z(n34170) );
  NANDN U34862 ( .A(n34055), .B(n34054), .Z(n34059) );
  NANDN U34863 ( .A(n34057), .B(n34056), .Z(n34058) );
  AND U34864 ( .A(n34059), .B(n34058), .Z(n34169) );
  XOR U34865 ( .A(n34170), .B(n34169), .Z(n34283) );
  NANDN U34866 ( .A(n34061), .B(n34060), .Z(n34065) );
  NANDN U34867 ( .A(n34063), .B(n34062), .Z(n34064) );
  AND U34868 ( .A(n34065), .B(n34064), .Z(n34281) );
  NANDN U34869 ( .A(n34067), .B(n34066), .Z(n34071) );
  NANDN U34870 ( .A(n34069), .B(n34068), .Z(n34070) );
  AND U34871 ( .A(n34071), .B(n34070), .Z(n34164) );
  NANDN U34872 ( .A(n34073), .B(n34072), .Z(n34077) );
  OR U34873 ( .A(n34075), .B(n34074), .Z(n34076) );
  AND U34874 ( .A(n34077), .B(n34076), .Z(n34162) );
  NANDN U34875 ( .A(n34079), .B(n34078), .Z(n34083) );
  NANDN U34876 ( .A(n34081), .B(n34080), .Z(n34082) );
  AND U34877 ( .A(n34083), .B(n34082), .Z(n34228) );
  NANDN U34878 ( .A(n34085), .B(n34084), .Z(n34089) );
  NANDN U34879 ( .A(n34087), .B(n34086), .Z(n34088) );
  NAND U34880 ( .A(n34089), .B(n34088), .Z(n34227) );
  XNOR U34881 ( .A(n34228), .B(n34227), .Z(n34229) );
  NAND U34882 ( .A(b[0]), .B(a[244]), .Z(n34090) );
  XNOR U34883 ( .A(b[1]), .B(n34090), .Z(n34092) );
  NANDN U34884 ( .A(b[0]), .B(a[243]), .Z(n34091) );
  NAND U34885 ( .A(n34092), .B(n34091), .Z(n34176) );
  NAND U34886 ( .A(n194), .B(n34093), .Z(n34095) );
  XOR U34887 ( .A(b[29]), .B(a[216]), .Z(n34254) );
  NAND U34888 ( .A(n38456), .B(n34254), .Z(n34094) );
  AND U34889 ( .A(n34095), .B(n34094), .Z(n34174) );
  AND U34890 ( .A(b[31]), .B(a[212]), .Z(n34173) );
  XNOR U34891 ( .A(n34174), .B(n34173), .Z(n34175) );
  XNOR U34892 ( .A(n34176), .B(n34175), .Z(n34215) );
  NAND U34893 ( .A(n38185), .B(n34096), .Z(n34098) );
  XOR U34894 ( .A(b[23]), .B(a[222]), .Z(n34257) );
  NAND U34895 ( .A(n38132), .B(n34257), .Z(n34097) );
  AND U34896 ( .A(n34098), .B(n34097), .Z(n34248) );
  NAND U34897 ( .A(n184), .B(n34099), .Z(n34101) );
  XOR U34898 ( .A(a[238]), .B(b[7]), .Z(n34260) );
  NAND U34899 ( .A(n36592), .B(n34260), .Z(n34100) );
  AND U34900 ( .A(n34101), .B(n34100), .Z(n34246) );
  NAND U34901 ( .A(n38289), .B(n34102), .Z(n34104) );
  XOR U34902 ( .A(b[25]), .B(a[220]), .Z(n34263) );
  NAND U34903 ( .A(n38247), .B(n34263), .Z(n34103) );
  NAND U34904 ( .A(n34104), .B(n34103), .Z(n34245) );
  XNOR U34905 ( .A(n34246), .B(n34245), .Z(n34247) );
  XOR U34906 ( .A(n34248), .B(n34247), .Z(n34216) );
  XNOR U34907 ( .A(n34215), .B(n34216), .Z(n34217) );
  NAND U34908 ( .A(n187), .B(n34105), .Z(n34107) );
  XOR U34909 ( .A(b[13]), .B(a[232]), .Z(n34266) );
  NAND U34910 ( .A(n37295), .B(n34266), .Z(n34106) );
  AND U34911 ( .A(n34107), .B(n34106), .Z(n34210) );
  NAND U34912 ( .A(n186), .B(n34108), .Z(n34110) );
  XOR U34913 ( .A(b[11]), .B(a[234]), .Z(n34269) );
  NAND U34914 ( .A(n37097), .B(n34269), .Z(n34109) );
  NAND U34915 ( .A(n34110), .B(n34109), .Z(n34209) );
  XNOR U34916 ( .A(n34210), .B(n34209), .Z(n34211) );
  NAND U34917 ( .A(n188), .B(n34111), .Z(n34113) );
  XOR U34918 ( .A(b[15]), .B(a[230]), .Z(n34272) );
  NAND U34919 ( .A(n37382), .B(n34272), .Z(n34112) );
  AND U34920 ( .A(n34113), .B(n34112), .Z(n34206) );
  NAND U34921 ( .A(n38064), .B(n34114), .Z(n34116) );
  XOR U34922 ( .A(b[21]), .B(a[224]), .Z(n34275) );
  NAND U34923 ( .A(n37993), .B(n34275), .Z(n34115) );
  AND U34924 ( .A(n34116), .B(n34115), .Z(n34204) );
  NAND U34925 ( .A(n185), .B(n34117), .Z(n34119) );
  XOR U34926 ( .A(a[236]), .B(b[9]), .Z(n34278) );
  NAND U34927 ( .A(n36805), .B(n34278), .Z(n34118) );
  NAND U34928 ( .A(n34119), .B(n34118), .Z(n34203) );
  XNOR U34929 ( .A(n34204), .B(n34203), .Z(n34205) );
  XOR U34930 ( .A(n34206), .B(n34205), .Z(n34212) );
  XOR U34931 ( .A(n34211), .B(n34212), .Z(n34218) );
  XOR U34932 ( .A(n34217), .B(n34218), .Z(n34230) );
  XNOR U34933 ( .A(n34229), .B(n34230), .Z(n34161) );
  XNOR U34934 ( .A(n34162), .B(n34161), .Z(n34163) );
  XOR U34935 ( .A(n34164), .B(n34163), .Z(n34282) );
  XOR U34936 ( .A(n34281), .B(n34282), .Z(n34284) );
  XOR U34937 ( .A(n34283), .B(n34284), .Z(n34158) );
  NANDN U34938 ( .A(n34121), .B(n34120), .Z(n34125) );
  NAND U34939 ( .A(n34123), .B(n34122), .Z(n34124) );
  AND U34940 ( .A(n34125), .B(n34124), .Z(n34156) );
  NANDN U34941 ( .A(n34127), .B(n34126), .Z(n34131) );
  NANDN U34942 ( .A(n34129), .B(n34128), .Z(n34130) );
  AND U34943 ( .A(n34131), .B(n34130), .Z(n34155) );
  XNOR U34944 ( .A(n34156), .B(n34155), .Z(n34157) );
  XNOR U34945 ( .A(n34158), .B(n34157), .Z(n34149) );
  NANDN U34946 ( .A(n34133), .B(n34132), .Z(n34137) );
  NANDN U34947 ( .A(n34135), .B(n34134), .Z(n34136) );
  NAND U34948 ( .A(n34137), .B(n34136), .Z(n34150) );
  XOR U34949 ( .A(n34149), .B(n34150), .Z(n34152) );
  XNOR U34950 ( .A(n34151), .B(n34152), .Z(n34143) );
  XNOR U34951 ( .A(n34144), .B(n34143), .Z(n34145) );
  XNOR U34952 ( .A(n34146), .B(n34145), .Z(n34287) );
  XNOR U34953 ( .A(sreg[468]), .B(n34287), .Z(n34289) );
  NANDN U34954 ( .A(sreg[467]), .B(n34138), .Z(n34142) );
  NAND U34955 ( .A(n34140), .B(n34139), .Z(n34141) );
  NAND U34956 ( .A(n34142), .B(n34141), .Z(n34288) );
  XNOR U34957 ( .A(n34289), .B(n34288), .Z(c[468]) );
  NANDN U34958 ( .A(n34144), .B(n34143), .Z(n34148) );
  NANDN U34959 ( .A(n34146), .B(n34145), .Z(n34147) );
  AND U34960 ( .A(n34148), .B(n34147), .Z(n34295) );
  NANDN U34961 ( .A(n34150), .B(n34149), .Z(n34154) );
  NANDN U34962 ( .A(n34152), .B(n34151), .Z(n34153) );
  AND U34963 ( .A(n34154), .B(n34153), .Z(n34293) );
  NANDN U34964 ( .A(n34156), .B(n34155), .Z(n34160) );
  NANDN U34965 ( .A(n34158), .B(n34157), .Z(n34159) );
  AND U34966 ( .A(n34160), .B(n34159), .Z(n34301) );
  NANDN U34967 ( .A(n34162), .B(n34161), .Z(n34166) );
  NANDN U34968 ( .A(n34164), .B(n34163), .Z(n34165) );
  AND U34969 ( .A(n34166), .B(n34165), .Z(n34305) );
  NANDN U34970 ( .A(n34168), .B(n34167), .Z(n34172) );
  NAND U34971 ( .A(n34170), .B(n34169), .Z(n34171) );
  AND U34972 ( .A(n34172), .B(n34171), .Z(n34304) );
  XNOR U34973 ( .A(n34305), .B(n34304), .Z(n34307) );
  NANDN U34974 ( .A(n34174), .B(n34173), .Z(n34178) );
  NANDN U34975 ( .A(n34176), .B(n34175), .Z(n34177) );
  AND U34976 ( .A(n34178), .B(n34177), .Z(n34384) );
  NAND U34977 ( .A(n38385), .B(n34179), .Z(n34181) );
  XOR U34978 ( .A(b[27]), .B(a[219]), .Z(n34328) );
  NAND U34979 ( .A(n38343), .B(n34328), .Z(n34180) );
  AND U34980 ( .A(n34181), .B(n34180), .Z(n34391) );
  NAND U34981 ( .A(n183), .B(n34182), .Z(n34184) );
  XOR U34982 ( .A(a[241]), .B(b[5]), .Z(n34331) );
  NAND U34983 ( .A(n36296), .B(n34331), .Z(n34183) );
  AND U34984 ( .A(n34184), .B(n34183), .Z(n34389) );
  NAND U34985 ( .A(n190), .B(n34185), .Z(n34187) );
  XOR U34986 ( .A(b[19]), .B(a[227]), .Z(n34334) );
  NAND U34987 ( .A(n37821), .B(n34334), .Z(n34186) );
  NAND U34988 ( .A(n34187), .B(n34186), .Z(n34388) );
  XNOR U34989 ( .A(n34389), .B(n34388), .Z(n34390) );
  XNOR U34990 ( .A(n34391), .B(n34390), .Z(n34382) );
  NAND U34991 ( .A(n38470), .B(n34188), .Z(n34190) );
  XOR U34992 ( .A(b[31]), .B(a[215]), .Z(n34337) );
  NAND U34993 ( .A(n38453), .B(n34337), .Z(n34189) );
  AND U34994 ( .A(n34190), .B(n34189), .Z(n34349) );
  NAND U34995 ( .A(n181), .B(n34191), .Z(n34193) );
  XOR U34996 ( .A(a[243]), .B(b[3]), .Z(n34340) );
  NAND U34997 ( .A(n182), .B(n34340), .Z(n34192) );
  AND U34998 ( .A(n34193), .B(n34192), .Z(n34347) );
  NAND U34999 ( .A(n189), .B(n34194), .Z(n34196) );
  XOR U35000 ( .A(b[17]), .B(a[229]), .Z(n34343) );
  NAND U35001 ( .A(n37652), .B(n34343), .Z(n34195) );
  NAND U35002 ( .A(n34196), .B(n34195), .Z(n34346) );
  XNOR U35003 ( .A(n34347), .B(n34346), .Z(n34348) );
  XOR U35004 ( .A(n34349), .B(n34348), .Z(n34383) );
  XOR U35005 ( .A(n34382), .B(n34383), .Z(n34385) );
  XOR U35006 ( .A(n34384), .B(n34385), .Z(n34317) );
  NANDN U35007 ( .A(n34198), .B(n34197), .Z(n34202) );
  NANDN U35008 ( .A(n34200), .B(n34199), .Z(n34201) );
  AND U35009 ( .A(n34202), .B(n34201), .Z(n34370) );
  NANDN U35010 ( .A(n34204), .B(n34203), .Z(n34208) );
  NANDN U35011 ( .A(n34206), .B(n34205), .Z(n34207) );
  NAND U35012 ( .A(n34208), .B(n34207), .Z(n34371) );
  XNOR U35013 ( .A(n34370), .B(n34371), .Z(n34372) );
  NANDN U35014 ( .A(n34210), .B(n34209), .Z(n34214) );
  NANDN U35015 ( .A(n34212), .B(n34211), .Z(n34213) );
  NAND U35016 ( .A(n34214), .B(n34213), .Z(n34373) );
  XNOR U35017 ( .A(n34372), .B(n34373), .Z(n34316) );
  XNOR U35018 ( .A(n34317), .B(n34316), .Z(n34319) );
  NANDN U35019 ( .A(n34216), .B(n34215), .Z(n34220) );
  NANDN U35020 ( .A(n34218), .B(n34217), .Z(n34219) );
  AND U35021 ( .A(n34220), .B(n34219), .Z(n34318) );
  XOR U35022 ( .A(n34319), .B(n34318), .Z(n34433) );
  NANDN U35023 ( .A(n34222), .B(n34221), .Z(n34226) );
  NANDN U35024 ( .A(n34224), .B(n34223), .Z(n34225) );
  AND U35025 ( .A(n34226), .B(n34225), .Z(n34430) );
  NANDN U35026 ( .A(n34228), .B(n34227), .Z(n34232) );
  NANDN U35027 ( .A(n34230), .B(n34229), .Z(n34231) );
  AND U35028 ( .A(n34232), .B(n34231), .Z(n34313) );
  NANDN U35029 ( .A(n34234), .B(n34233), .Z(n34238) );
  OR U35030 ( .A(n34236), .B(n34235), .Z(n34237) );
  AND U35031 ( .A(n34238), .B(n34237), .Z(n34311) );
  NANDN U35032 ( .A(n34240), .B(n34239), .Z(n34244) );
  NANDN U35033 ( .A(n34242), .B(n34241), .Z(n34243) );
  AND U35034 ( .A(n34244), .B(n34243), .Z(n34377) );
  NANDN U35035 ( .A(n34246), .B(n34245), .Z(n34250) );
  NANDN U35036 ( .A(n34248), .B(n34247), .Z(n34249) );
  NAND U35037 ( .A(n34250), .B(n34249), .Z(n34376) );
  XNOR U35038 ( .A(n34377), .B(n34376), .Z(n34378) );
  NAND U35039 ( .A(b[0]), .B(a[245]), .Z(n34251) );
  XNOR U35040 ( .A(b[1]), .B(n34251), .Z(n34253) );
  NANDN U35041 ( .A(b[0]), .B(a[244]), .Z(n34252) );
  NAND U35042 ( .A(n34253), .B(n34252), .Z(n34325) );
  NAND U35043 ( .A(n194), .B(n34254), .Z(n34256) );
  XOR U35044 ( .A(b[29]), .B(a[217]), .Z(n34400) );
  NAND U35045 ( .A(n38456), .B(n34400), .Z(n34255) );
  AND U35046 ( .A(n34256), .B(n34255), .Z(n34323) );
  AND U35047 ( .A(b[31]), .B(a[213]), .Z(n34322) );
  XNOR U35048 ( .A(n34323), .B(n34322), .Z(n34324) );
  XNOR U35049 ( .A(n34325), .B(n34324), .Z(n34364) );
  NAND U35050 ( .A(n38185), .B(n34257), .Z(n34259) );
  XOR U35051 ( .A(b[23]), .B(a[223]), .Z(n34406) );
  NAND U35052 ( .A(n38132), .B(n34406), .Z(n34258) );
  AND U35053 ( .A(n34259), .B(n34258), .Z(n34397) );
  NAND U35054 ( .A(n184), .B(n34260), .Z(n34262) );
  XOR U35055 ( .A(a[239]), .B(b[7]), .Z(n34409) );
  NAND U35056 ( .A(n36592), .B(n34409), .Z(n34261) );
  AND U35057 ( .A(n34262), .B(n34261), .Z(n34395) );
  NAND U35058 ( .A(n38289), .B(n34263), .Z(n34265) );
  XOR U35059 ( .A(b[25]), .B(a[221]), .Z(n34412) );
  NAND U35060 ( .A(n38247), .B(n34412), .Z(n34264) );
  NAND U35061 ( .A(n34265), .B(n34264), .Z(n34394) );
  XNOR U35062 ( .A(n34395), .B(n34394), .Z(n34396) );
  XOR U35063 ( .A(n34397), .B(n34396), .Z(n34365) );
  XNOR U35064 ( .A(n34364), .B(n34365), .Z(n34366) );
  NAND U35065 ( .A(n187), .B(n34266), .Z(n34268) );
  XOR U35066 ( .A(b[13]), .B(a[233]), .Z(n34415) );
  NAND U35067 ( .A(n37295), .B(n34415), .Z(n34267) );
  AND U35068 ( .A(n34268), .B(n34267), .Z(n34359) );
  NAND U35069 ( .A(n186), .B(n34269), .Z(n34271) );
  XOR U35070 ( .A(b[11]), .B(a[235]), .Z(n34418) );
  NAND U35071 ( .A(n37097), .B(n34418), .Z(n34270) );
  NAND U35072 ( .A(n34271), .B(n34270), .Z(n34358) );
  XNOR U35073 ( .A(n34359), .B(n34358), .Z(n34360) );
  NAND U35074 ( .A(n188), .B(n34272), .Z(n34274) );
  XOR U35075 ( .A(b[15]), .B(a[231]), .Z(n34421) );
  NAND U35076 ( .A(n37382), .B(n34421), .Z(n34273) );
  AND U35077 ( .A(n34274), .B(n34273), .Z(n34355) );
  NAND U35078 ( .A(n38064), .B(n34275), .Z(n34277) );
  XOR U35079 ( .A(b[21]), .B(a[225]), .Z(n34424) );
  NAND U35080 ( .A(n37993), .B(n34424), .Z(n34276) );
  AND U35081 ( .A(n34277), .B(n34276), .Z(n34353) );
  NAND U35082 ( .A(n185), .B(n34278), .Z(n34280) );
  XOR U35083 ( .A(a[237]), .B(b[9]), .Z(n34427) );
  NAND U35084 ( .A(n36805), .B(n34427), .Z(n34279) );
  NAND U35085 ( .A(n34280), .B(n34279), .Z(n34352) );
  XNOR U35086 ( .A(n34353), .B(n34352), .Z(n34354) );
  XOR U35087 ( .A(n34355), .B(n34354), .Z(n34361) );
  XOR U35088 ( .A(n34360), .B(n34361), .Z(n34367) );
  XOR U35089 ( .A(n34366), .B(n34367), .Z(n34379) );
  XNOR U35090 ( .A(n34378), .B(n34379), .Z(n34310) );
  XNOR U35091 ( .A(n34311), .B(n34310), .Z(n34312) );
  XOR U35092 ( .A(n34313), .B(n34312), .Z(n34431) );
  XNOR U35093 ( .A(n34430), .B(n34431), .Z(n34432) );
  XNOR U35094 ( .A(n34433), .B(n34432), .Z(n34306) );
  XOR U35095 ( .A(n34307), .B(n34306), .Z(n34299) );
  NANDN U35096 ( .A(n34282), .B(n34281), .Z(n34286) );
  OR U35097 ( .A(n34284), .B(n34283), .Z(n34285) );
  AND U35098 ( .A(n34286), .B(n34285), .Z(n34298) );
  XNOR U35099 ( .A(n34299), .B(n34298), .Z(n34300) );
  XNOR U35100 ( .A(n34301), .B(n34300), .Z(n34292) );
  XNOR U35101 ( .A(n34293), .B(n34292), .Z(n34294) );
  XNOR U35102 ( .A(n34295), .B(n34294), .Z(n34436) );
  XNOR U35103 ( .A(sreg[469]), .B(n34436), .Z(n34438) );
  NANDN U35104 ( .A(sreg[468]), .B(n34287), .Z(n34291) );
  NAND U35105 ( .A(n34289), .B(n34288), .Z(n34290) );
  NAND U35106 ( .A(n34291), .B(n34290), .Z(n34437) );
  XNOR U35107 ( .A(n34438), .B(n34437), .Z(c[469]) );
  NANDN U35108 ( .A(n34293), .B(n34292), .Z(n34297) );
  NANDN U35109 ( .A(n34295), .B(n34294), .Z(n34296) );
  AND U35110 ( .A(n34297), .B(n34296), .Z(n34444) );
  NANDN U35111 ( .A(n34299), .B(n34298), .Z(n34303) );
  NANDN U35112 ( .A(n34301), .B(n34300), .Z(n34302) );
  AND U35113 ( .A(n34303), .B(n34302), .Z(n34442) );
  NANDN U35114 ( .A(n34305), .B(n34304), .Z(n34309) );
  NAND U35115 ( .A(n34307), .B(n34306), .Z(n34308) );
  AND U35116 ( .A(n34309), .B(n34308), .Z(n34449) );
  NANDN U35117 ( .A(n34311), .B(n34310), .Z(n34315) );
  NANDN U35118 ( .A(n34313), .B(n34312), .Z(n34314) );
  AND U35119 ( .A(n34315), .B(n34314), .Z(n34580) );
  NANDN U35120 ( .A(n34317), .B(n34316), .Z(n34321) );
  NAND U35121 ( .A(n34319), .B(n34318), .Z(n34320) );
  AND U35122 ( .A(n34321), .B(n34320), .Z(n34579) );
  XNOR U35123 ( .A(n34580), .B(n34579), .Z(n34582) );
  NANDN U35124 ( .A(n34323), .B(n34322), .Z(n34327) );
  NANDN U35125 ( .A(n34325), .B(n34324), .Z(n34326) );
  AND U35126 ( .A(n34327), .B(n34326), .Z(n34527) );
  NAND U35127 ( .A(n38385), .B(n34328), .Z(n34330) );
  XOR U35128 ( .A(b[27]), .B(a[220]), .Z(n34471) );
  NAND U35129 ( .A(n38343), .B(n34471), .Z(n34329) );
  AND U35130 ( .A(n34330), .B(n34329), .Z(n34534) );
  NAND U35131 ( .A(n183), .B(n34331), .Z(n34333) );
  XOR U35132 ( .A(a[242]), .B(b[5]), .Z(n34474) );
  NAND U35133 ( .A(n36296), .B(n34474), .Z(n34332) );
  AND U35134 ( .A(n34333), .B(n34332), .Z(n34532) );
  NAND U35135 ( .A(n190), .B(n34334), .Z(n34336) );
  XOR U35136 ( .A(b[19]), .B(a[228]), .Z(n34477) );
  NAND U35137 ( .A(n37821), .B(n34477), .Z(n34335) );
  NAND U35138 ( .A(n34336), .B(n34335), .Z(n34531) );
  XNOR U35139 ( .A(n34532), .B(n34531), .Z(n34533) );
  XNOR U35140 ( .A(n34534), .B(n34533), .Z(n34525) );
  NAND U35141 ( .A(n38470), .B(n34337), .Z(n34339) );
  XOR U35142 ( .A(b[31]), .B(a[216]), .Z(n34480) );
  NAND U35143 ( .A(n38453), .B(n34480), .Z(n34338) );
  AND U35144 ( .A(n34339), .B(n34338), .Z(n34492) );
  NAND U35145 ( .A(n181), .B(n34340), .Z(n34342) );
  XOR U35146 ( .A(a[244]), .B(b[3]), .Z(n34483) );
  NAND U35147 ( .A(n182), .B(n34483), .Z(n34341) );
  AND U35148 ( .A(n34342), .B(n34341), .Z(n34490) );
  NAND U35149 ( .A(n189), .B(n34343), .Z(n34345) );
  XOR U35150 ( .A(b[17]), .B(a[230]), .Z(n34486) );
  NAND U35151 ( .A(n37652), .B(n34486), .Z(n34344) );
  NAND U35152 ( .A(n34345), .B(n34344), .Z(n34489) );
  XNOR U35153 ( .A(n34490), .B(n34489), .Z(n34491) );
  XOR U35154 ( .A(n34492), .B(n34491), .Z(n34526) );
  XOR U35155 ( .A(n34525), .B(n34526), .Z(n34528) );
  XOR U35156 ( .A(n34527), .B(n34528), .Z(n34460) );
  NANDN U35157 ( .A(n34347), .B(n34346), .Z(n34351) );
  NANDN U35158 ( .A(n34349), .B(n34348), .Z(n34350) );
  AND U35159 ( .A(n34351), .B(n34350), .Z(n34513) );
  NANDN U35160 ( .A(n34353), .B(n34352), .Z(n34357) );
  NANDN U35161 ( .A(n34355), .B(n34354), .Z(n34356) );
  NAND U35162 ( .A(n34357), .B(n34356), .Z(n34514) );
  XNOR U35163 ( .A(n34513), .B(n34514), .Z(n34515) );
  NANDN U35164 ( .A(n34359), .B(n34358), .Z(n34363) );
  NANDN U35165 ( .A(n34361), .B(n34360), .Z(n34362) );
  NAND U35166 ( .A(n34363), .B(n34362), .Z(n34516) );
  XNOR U35167 ( .A(n34515), .B(n34516), .Z(n34459) );
  XNOR U35168 ( .A(n34460), .B(n34459), .Z(n34462) );
  NANDN U35169 ( .A(n34365), .B(n34364), .Z(n34369) );
  NANDN U35170 ( .A(n34367), .B(n34366), .Z(n34368) );
  AND U35171 ( .A(n34369), .B(n34368), .Z(n34461) );
  XOR U35172 ( .A(n34462), .B(n34461), .Z(n34576) );
  NANDN U35173 ( .A(n34371), .B(n34370), .Z(n34375) );
  NANDN U35174 ( .A(n34373), .B(n34372), .Z(n34374) );
  AND U35175 ( .A(n34375), .B(n34374), .Z(n34573) );
  NANDN U35176 ( .A(n34377), .B(n34376), .Z(n34381) );
  NANDN U35177 ( .A(n34379), .B(n34378), .Z(n34380) );
  AND U35178 ( .A(n34381), .B(n34380), .Z(n34456) );
  NANDN U35179 ( .A(n34383), .B(n34382), .Z(n34387) );
  OR U35180 ( .A(n34385), .B(n34384), .Z(n34386) );
  AND U35181 ( .A(n34387), .B(n34386), .Z(n34454) );
  NANDN U35182 ( .A(n34389), .B(n34388), .Z(n34393) );
  NANDN U35183 ( .A(n34391), .B(n34390), .Z(n34392) );
  AND U35184 ( .A(n34393), .B(n34392), .Z(n34520) );
  NANDN U35185 ( .A(n34395), .B(n34394), .Z(n34399) );
  NANDN U35186 ( .A(n34397), .B(n34396), .Z(n34398) );
  NAND U35187 ( .A(n34399), .B(n34398), .Z(n34519) );
  XNOR U35188 ( .A(n34520), .B(n34519), .Z(n34521) );
  NAND U35189 ( .A(n194), .B(n34400), .Z(n34402) );
  XOR U35190 ( .A(b[29]), .B(a[218]), .Z(n34543) );
  NAND U35191 ( .A(n38456), .B(n34543), .Z(n34401) );
  AND U35192 ( .A(n34402), .B(n34401), .Z(n34466) );
  AND U35193 ( .A(b[31]), .B(a[214]), .Z(n34465) );
  XNOR U35194 ( .A(n34466), .B(n34465), .Z(n34467) );
  NAND U35195 ( .A(b[0]), .B(a[246]), .Z(n34403) );
  XNOR U35196 ( .A(b[1]), .B(n34403), .Z(n34405) );
  NANDN U35197 ( .A(b[0]), .B(a[245]), .Z(n34404) );
  NAND U35198 ( .A(n34405), .B(n34404), .Z(n34468) );
  XNOR U35199 ( .A(n34467), .B(n34468), .Z(n34507) );
  NAND U35200 ( .A(n38185), .B(n34406), .Z(n34408) );
  XOR U35201 ( .A(b[23]), .B(a[224]), .Z(n34549) );
  NAND U35202 ( .A(n38132), .B(n34549), .Z(n34407) );
  AND U35203 ( .A(n34408), .B(n34407), .Z(n34540) );
  NAND U35204 ( .A(n184), .B(n34409), .Z(n34411) );
  XOR U35205 ( .A(a[240]), .B(b[7]), .Z(n34552) );
  NAND U35206 ( .A(n36592), .B(n34552), .Z(n34410) );
  AND U35207 ( .A(n34411), .B(n34410), .Z(n34538) );
  NAND U35208 ( .A(n38289), .B(n34412), .Z(n34414) );
  XOR U35209 ( .A(b[25]), .B(a[222]), .Z(n34555) );
  NAND U35210 ( .A(n38247), .B(n34555), .Z(n34413) );
  NAND U35211 ( .A(n34414), .B(n34413), .Z(n34537) );
  XNOR U35212 ( .A(n34538), .B(n34537), .Z(n34539) );
  XOR U35213 ( .A(n34540), .B(n34539), .Z(n34508) );
  XNOR U35214 ( .A(n34507), .B(n34508), .Z(n34509) );
  NAND U35215 ( .A(n187), .B(n34415), .Z(n34417) );
  XOR U35216 ( .A(b[13]), .B(a[234]), .Z(n34558) );
  NAND U35217 ( .A(n37295), .B(n34558), .Z(n34416) );
  AND U35218 ( .A(n34417), .B(n34416), .Z(n34502) );
  NAND U35219 ( .A(n186), .B(n34418), .Z(n34420) );
  XOR U35220 ( .A(b[11]), .B(a[236]), .Z(n34561) );
  NAND U35221 ( .A(n37097), .B(n34561), .Z(n34419) );
  NAND U35222 ( .A(n34420), .B(n34419), .Z(n34501) );
  XNOR U35223 ( .A(n34502), .B(n34501), .Z(n34503) );
  NAND U35224 ( .A(n188), .B(n34421), .Z(n34423) );
  XOR U35225 ( .A(b[15]), .B(a[232]), .Z(n34564) );
  NAND U35226 ( .A(n37382), .B(n34564), .Z(n34422) );
  AND U35227 ( .A(n34423), .B(n34422), .Z(n34498) );
  NAND U35228 ( .A(n38064), .B(n34424), .Z(n34426) );
  XOR U35229 ( .A(b[21]), .B(a[226]), .Z(n34567) );
  NAND U35230 ( .A(n37993), .B(n34567), .Z(n34425) );
  AND U35231 ( .A(n34426), .B(n34425), .Z(n34496) );
  NAND U35232 ( .A(n185), .B(n34427), .Z(n34429) );
  XOR U35233 ( .A(a[238]), .B(b[9]), .Z(n34570) );
  NAND U35234 ( .A(n36805), .B(n34570), .Z(n34428) );
  NAND U35235 ( .A(n34429), .B(n34428), .Z(n34495) );
  XNOR U35236 ( .A(n34496), .B(n34495), .Z(n34497) );
  XOR U35237 ( .A(n34498), .B(n34497), .Z(n34504) );
  XOR U35238 ( .A(n34503), .B(n34504), .Z(n34510) );
  XOR U35239 ( .A(n34509), .B(n34510), .Z(n34522) );
  XNOR U35240 ( .A(n34521), .B(n34522), .Z(n34453) );
  XNOR U35241 ( .A(n34454), .B(n34453), .Z(n34455) );
  XOR U35242 ( .A(n34456), .B(n34455), .Z(n34574) );
  XNOR U35243 ( .A(n34573), .B(n34574), .Z(n34575) );
  XNOR U35244 ( .A(n34576), .B(n34575), .Z(n34581) );
  XOR U35245 ( .A(n34582), .B(n34581), .Z(n34448) );
  NANDN U35246 ( .A(n34431), .B(n34430), .Z(n34435) );
  NANDN U35247 ( .A(n34433), .B(n34432), .Z(n34434) );
  AND U35248 ( .A(n34435), .B(n34434), .Z(n34447) );
  XOR U35249 ( .A(n34448), .B(n34447), .Z(n34450) );
  XNOR U35250 ( .A(n34449), .B(n34450), .Z(n34441) );
  XNOR U35251 ( .A(n34442), .B(n34441), .Z(n34443) );
  XNOR U35252 ( .A(n34444), .B(n34443), .Z(n34585) );
  XNOR U35253 ( .A(sreg[470]), .B(n34585), .Z(n34587) );
  NANDN U35254 ( .A(sreg[469]), .B(n34436), .Z(n34440) );
  NAND U35255 ( .A(n34438), .B(n34437), .Z(n34439) );
  NAND U35256 ( .A(n34440), .B(n34439), .Z(n34586) );
  XNOR U35257 ( .A(n34587), .B(n34586), .Z(c[470]) );
  NANDN U35258 ( .A(n34442), .B(n34441), .Z(n34446) );
  NANDN U35259 ( .A(n34444), .B(n34443), .Z(n34445) );
  AND U35260 ( .A(n34446), .B(n34445), .Z(n34593) );
  NANDN U35261 ( .A(n34448), .B(n34447), .Z(n34452) );
  NANDN U35262 ( .A(n34450), .B(n34449), .Z(n34451) );
  AND U35263 ( .A(n34452), .B(n34451), .Z(n34591) );
  NANDN U35264 ( .A(n34454), .B(n34453), .Z(n34458) );
  NANDN U35265 ( .A(n34456), .B(n34455), .Z(n34457) );
  AND U35266 ( .A(n34458), .B(n34457), .Z(n34729) );
  NANDN U35267 ( .A(n34460), .B(n34459), .Z(n34464) );
  NAND U35268 ( .A(n34462), .B(n34461), .Z(n34463) );
  AND U35269 ( .A(n34464), .B(n34463), .Z(n34728) );
  XNOR U35270 ( .A(n34729), .B(n34728), .Z(n34731) );
  NANDN U35271 ( .A(n34466), .B(n34465), .Z(n34470) );
  NANDN U35272 ( .A(n34468), .B(n34467), .Z(n34469) );
  AND U35273 ( .A(n34470), .B(n34469), .Z(n34676) );
  NAND U35274 ( .A(n38385), .B(n34471), .Z(n34473) );
  XOR U35275 ( .A(b[27]), .B(a[221]), .Z(n34620) );
  NAND U35276 ( .A(n38343), .B(n34620), .Z(n34472) );
  AND U35277 ( .A(n34473), .B(n34472), .Z(n34683) );
  NAND U35278 ( .A(n183), .B(n34474), .Z(n34476) );
  XOR U35279 ( .A(a[243]), .B(b[5]), .Z(n34623) );
  NAND U35280 ( .A(n36296), .B(n34623), .Z(n34475) );
  AND U35281 ( .A(n34476), .B(n34475), .Z(n34681) );
  NAND U35282 ( .A(n190), .B(n34477), .Z(n34479) );
  XOR U35283 ( .A(b[19]), .B(a[229]), .Z(n34626) );
  NAND U35284 ( .A(n37821), .B(n34626), .Z(n34478) );
  NAND U35285 ( .A(n34479), .B(n34478), .Z(n34680) );
  XNOR U35286 ( .A(n34681), .B(n34680), .Z(n34682) );
  XNOR U35287 ( .A(n34683), .B(n34682), .Z(n34674) );
  NAND U35288 ( .A(n38470), .B(n34480), .Z(n34482) );
  XOR U35289 ( .A(b[31]), .B(a[217]), .Z(n34629) );
  NAND U35290 ( .A(n38453), .B(n34629), .Z(n34481) );
  AND U35291 ( .A(n34482), .B(n34481), .Z(n34641) );
  NAND U35292 ( .A(n181), .B(n34483), .Z(n34485) );
  XOR U35293 ( .A(a[245]), .B(b[3]), .Z(n34632) );
  NAND U35294 ( .A(n182), .B(n34632), .Z(n34484) );
  AND U35295 ( .A(n34485), .B(n34484), .Z(n34639) );
  NAND U35296 ( .A(n189), .B(n34486), .Z(n34488) );
  XOR U35297 ( .A(b[17]), .B(a[231]), .Z(n34635) );
  NAND U35298 ( .A(n37652), .B(n34635), .Z(n34487) );
  NAND U35299 ( .A(n34488), .B(n34487), .Z(n34638) );
  XNOR U35300 ( .A(n34639), .B(n34638), .Z(n34640) );
  XOR U35301 ( .A(n34641), .B(n34640), .Z(n34675) );
  XOR U35302 ( .A(n34674), .B(n34675), .Z(n34677) );
  XOR U35303 ( .A(n34676), .B(n34677), .Z(n34609) );
  NANDN U35304 ( .A(n34490), .B(n34489), .Z(n34494) );
  NANDN U35305 ( .A(n34492), .B(n34491), .Z(n34493) );
  AND U35306 ( .A(n34494), .B(n34493), .Z(n34662) );
  NANDN U35307 ( .A(n34496), .B(n34495), .Z(n34500) );
  NANDN U35308 ( .A(n34498), .B(n34497), .Z(n34499) );
  NAND U35309 ( .A(n34500), .B(n34499), .Z(n34663) );
  XNOR U35310 ( .A(n34662), .B(n34663), .Z(n34664) );
  NANDN U35311 ( .A(n34502), .B(n34501), .Z(n34506) );
  NANDN U35312 ( .A(n34504), .B(n34503), .Z(n34505) );
  NAND U35313 ( .A(n34506), .B(n34505), .Z(n34665) );
  XNOR U35314 ( .A(n34664), .B(n34665), .Z(n34608) );
  XNOR U35315 ( .A(n34609), .B(n34608), .Z(n34611) );
  NANDN U35316 ( .A(n34508), .B(n34507), .Z(n34512) );
  NANDN U35317 ( .A(n34510), .B(n34509), .Z(n34511) );
  AND U35318 ( .A(n34512), .B(n34511), .Z(n34610) );
  XOR U35319 ( .A(n34611), .B(n34610), .Z(n34725) );
  NANDN U35320 ( .A(n34514), .B(n34513), .Z(n34518) );
  NANDN U35321 ( .A(n34516), .B(n34515), .Z(n34517) );
  AND U35322 ( .A(n34518), .B(n34517), .Z(n34722) );
  NANDN U35323 ( .A(n34520), .B(n34519), .Z(n34524) );
  NANDN U35324 ( .A(n34522), .B(n34521), .Z(n34523) );
  AND U35325 ( .A(n34524), .B(n34523), .Z(n34605) );
  NANDN U35326 ( .A(n34526), .B(n34525), .Z(n34530) );
  OR U35327 ( .A(n34528), .B(n34527), .Z(n34529) );
  AND U35328 ( .A(n34530), .B(n34529), .Z(n34603) );
  NANDN U35329 ( .A(n34532), .B(n34531), .Z(n34536) );
  NANDN U35330 ( .A(n34534), .B(n34533), .Z(n34535) );
  AND U35331 ( .A(n34536), .B(n34535), .Z(n34669) );
  NANDN U35332 ( .A(n34538), .B(n34537), .Z(n34542) );
  NANDN U35333 ( .A(n34540), .B(n34539), .Z(n34541) );
  NAND U35334 ( .A(n34542), .B(n34541), .Z(n34668) );
  XNOR U35335 ( .A(n34669), .B(n34668), .Z(n34670) );
  NAND U35336 ( .A(n194), .B(n34543), .Z(n34545) );
  XOR U35337 ( .A(b[29]), .B(a[219]), .Z(n34692) );
  NAND U35338 ( .A(n38456), .B(n34692), .Z(n34544) );
  AND U35339 ( .A(n34545), .B(n34544), .Z(n34615) );
  AND U35340 ( .A(b[31]), .B(a[215]), .Z(n34614) );
  XNOR U35341 ( .A(n34615), .B(n34614), .Z(n34616) );
  NAND U35342 ( .A(b[0]), .B(a[247]), .Z(n34546) );
  XNOR U35343 ( .A(b[1]), .B(n34546), .Z(n34548) );
  NANDN U35344 ( .A(b[0]), .B(a[246]), .Z(n34547) );
  NAND U35345 ( .A(n34548), .B(n34547), .Z(n34617) );
  XNOR U35346 ( .A(n34616), .B(n34617), .Z(n34656) );
  NAND U35347 ( .A(n38185), .B(n34549), .Z(n34551) );
  XOR U35348 ( .A(b[23]), .B(a[225]), .Z(n34698) );
  NAND U35349 ( .A(n38132), .B(n34698), .Z(n34550) );
  AND U35350 ( .A(n34551), .B(n34550), .Z(n34689) );
  NAND U35351 ( .A(n184), .B(n34552), .Z(n34554) );
  XOR U35352 ( .A(a[241]), .B(b[7]), .Z(n34701) );
  NAND U35353 ( .A(n36592), .B(n34701), .Z(n34553) );
  AND U35354 ( .A(n34554), .B(n34553), .Z(n34687) );
  NAND U35355 ( .A(n38289), .B(n34555), .Z(n34557) );
  XOR U35356 ( .A(b[25]), .B(a[223]), .Z(n34704) );
  NAND U35357 ( .A(n38247), .B(n34704), .Z(n34556) );
  NAND U35358 ( .A(n34557), .B(n34556), .Z(n34686) );
  XNOR U35359 ( .A(n34687), .B(n34686), .Z(n34688) );
  XOR U35360 ( .A(n34689), .B(n34688), .Z(n34657) );
  XNOR U35361 ( .A(n34656), .B(n34657), .Z(n34658) );
  NAND U35362 ( .A(n187), .B(n34558), .Z(n34560) );
  XOR U35363 ( .A(b[13]), .B(a[235]), .Z(n34707) );
  NAND U35364 ( .A(n37295), .B(n34707), .Z(n34559) );
  AND U35365 ( .A(n34560), .B(n34559), .Z(n34651) );
  NAND U35366 ( .A(n186), .B(n34561), .Z(n34563) );
  XOR U35367 ( .A(b[11]), .B(a[237]), .Z(n34710) );
  NAND U35368 ( .A(n37097), .B(n34710), .Z(n34562) );
  NAND U35369 ( .A(n34563), .B(n34562), .Z(n34650) );
  XNOR U35370 ( .A(n34651), .B(n34650), .Z(n34652) );
  NAND U35371 ( .A(n188), .B(n34564), .Z(n34566) );
  XOR U35372 ( .A(b[15]), .B(a[233]), .Z(n34713) );
  NAND U35373 ( .A(n37382), .B(n34713), .Z(n34565) );
  AND U35374 ( .A(n34566), .B(n34565), .Z(n34647) );
  NAND U35375 ( .A(n38064), .B(n34567), .Z(n34569) );
  XOR U35376 ( .A(b[21]), .B(a[227]), .Z(n34716) );
  NAND U35377 ( .A(n37993), .B(n34716), .Z(n34568) );
  AND U35378 ( .A(n34569), .B(n34568), .Z(n34645) );
  NAND U35379 ( .A(n185), .B(n34570), .Z(n34572) );
  XOR U35380 ( .A(a[239]), .B(b[9]), .Z(n34719) );
  NAND U35381 ( .A(n36805), .B(n34719), .Z(n34571) );
  NAND U35382 ( .A(n34572), .B(n34571), .Z(n34644) );
  XNOR U35383 ( .A(n34645), .B(n34644), .Z(n34646) );
  XOR U35384 ( .A(n34647), .B(n34646), .Z(n34653) );
  XOR U35385 ( .A(n34652), .B(n34653), .Z(n34659) );
  XOR U35386 ( .A(n34658), .B(n34659), .Z(n34671) );
  XNOR U35387 ( .A(n34670), .B(n34671), .Z(n34602) );
  XNOR U35388 ( .A(n34603), .B(n34602), .Z(n34604) );
  XOR U35389 ( .A(n34605), .B(n34604), .Z(n34723) );
  XNOR U35390 ( .A(n34722), .B(n34723), .Z(n34724) );
  XNOR U35391 ( .A(n34725), .B(n34724), .Z(n34730) );
  XOR U35392 ( .A(n34731), .B(n34730), .Z(n34597) );
  NANDN U35393 ( .A(n34574), .B(n34573), .Z(n34578) );
  NANDN U35394 ( .A(n34576), .B(n34575), .Z(n34577) );
  AND U35395 ( .A(n34578), .B(n34577), .Z(n34596) );
  XNOR U35396 ( .A(n34597), .B(n34596), .Z(n34598) );
  NANDN U35397 ( .A(n34580), .B(n34579), .Z(n34584) );
  NAND U35398 ( .A(n34582), .B(n34581), .Z(n34583) );
  NAND U35399 ( .A(n34584), .B(n34583), .Z(n34599) );
  XNOR U35400 ( .A(n34598), .B(n34599), .Z(n34590) );
  XNOR U35401 ( .A(n34591), .B(n34590), .Z(n34592) );
  XNOR U35402 ( .A(n34593), .B(n34592), .Z(n34734) );
  XNOR U35403 ( .A(sreg[471]), .B(n34734), .Z(n34736) );
  NANDN U35404 ( .A(sreg[470]), .B(n34585), .Z(n34589) );
  NAND U35405 ( .A(n34587), .B(n34586), .Z(n34588) );
  NAND U35406 ( .A(n34589), .B(n34588), .Z(n34735) );
  XNOR U35407 ( .A(n34736), .B(n34735), .Z(c[471]) );
  NANDN U35408 ( .A(n34591), .B(n34590), .Z(n34595) );
  NANDN U35409 ( .A(n34593), .B(n34592), .Z(n34594) );
  AND U35410 ( .A(n34595), .B(n34594), .Z(n34742) );
  NANDN U35411 ( .A(n34597), .B(n34596), .Z(n34601) );
  NANDN U35412 ( .A(n34599), .B(n34598), .Z(n34600) );
  AND U35413 ( .A(n34601), .B(n34600), .Z(n34740) );
  NANDN U35414 ( .A(n34603), .B(n34602), .Z(n34607) );
  NANDN U35415 ( .A(n34605), .B(n34604), .Z(n34606) );
  AND U35416 ( .A(n34607), .B(n34606), .Z(n34752) );
  NANDN U35417 ( .A(n34609), .B(n34608), .Z(n34613) );
  NAND U35418 ( .A(n34611), .B(n34610), .Z(n34612) );
  AND U35419 ( .A(n34613), .B(n34612), .Z(n34751) );
  XNOR U35420 ( .A(n34752), .B(n34751), .Z(n34754) );
  NANDN U35421 ( .A(n34615), .B(n34614), .Z(n34619) );
  NANDN U35422 ( .A(n34617), .B(n34616), .Z(n34618) );
  AND U35423 ( .A(n34619), .B(n34618), .Z(n34831) );
  NAND U35424 ( .A(n38385), .B(n34620), .Z(n34622) );
  XOR U35425 ( .A(b[27]), .B(a[222]), .Z(n34775) );
  NAND U35426 ( .A(n38343), .B(n34775), .Z(n34621) );
  AND U35427 ( .A(n34622), .B(n34621), .Z(n34838) );
  NAND U35428 ( .A(n183), .B(n34623), .Z(n34625) );
  XOR U35429 ( .A(a[244]), .B(b[5]), .Z(n34778) );
  NAND U35430 ( .A(n36296), .B(n34778), .Z(n34624) );
  AND U35431 ( .A(n34625), .B(n34624), .Z(n34836) );
  NAND U35432 ( .A(n190), .B(n34626), .Z(n34628) );
  XOR U35433 ( .A(b[19]), .B(a[230]), .Z(n34781) );
  NAND U35434 ( .A(n37821), .B(n34781), .Z(n34627) );
  NAND U35435 ( .A(n34628), .B(n34627), .Z(n34835) );
  XNOR U35436 ( .A(n34836), .B(n34835), .Z(n34837) );
  XNOR U35437 ( .A(n34838), .B(n34837), .Z(n34829) );
  NAND U35438 ( .A(n38470), .B(n34629), .Z(n34631) );
  XOR U35439 ( .A(b[31]), .B(a[218]), .Z(n34784) );
  NAND U35440 ( .A(n38453), .B(n34784), .Z(n34630) );
  AND U35441 ( .A(n34631), .B(n34630), .Z(n34796) );
  NAND U35442 ( .A(n181), .B(n34632), .Z(n34634) );
  XOR U35443 ( .A(a[246]), .B(b[3]), .Z(n34787) );
  NAND U35444 ( .A(n182), .B(n34787), .Z(n34633) );
  AND U35445 ( .A(n34634), .B(n34633), .Z(n34794) );
  NAND U35446 ( .A(n189), .B(n34635), .Z(n34637) );
  XOR U35447 ( .A(b[17]), .B(a[232]), .Z(n34790) );
  NAND U35448 ( .A(n37652), .B(n34790), .Z(n34636) );
  NAND U35449 ( .A(n34637), .B(n34636), .Z(n34793) );
  XNOR U35450 ( .A(n34794), .B(n34793), .Z(n34795) );
  XOR U35451 ( .A(n34796), .B(n34795), .Z(n34830) );
  XOR U35452 ( .A(n34829), .B(n34830), .Z(n34832) );
  XOR U35453 ( .A(n34831), .B(n34832), .Z(n34764) );
  NANDN U35454 ( .A(n34639), .B(n34638), .Z(n34643) );
  NANDN U35455 ( .A(n34641), .B(n34640), .Z(n34642) );
  AND U35456 ( .A(n34643), .B(n34642), .Z(n34817) );
  NANDN U35457 ( .A(n34645), .B(n34644), .Z(n34649) );
  NANDN U35458 ( .A(n34647), .B(n34646), .Z(n34648) );
  NAND U35459 ( .A(n34649), .B(n34648), .Z(n34818) );
  XNOR U35460 ( .A(n34817), .B(n34818), .Z(n34819) );
  NANDN U35461 ( .A(n34651), .B(n34650), .Z(n34655) );
  NANDN U35462 ( .A(n34653), .B(n34652), .Z(n34654) );
  NAND U35463 ( .A(n34655), .B(n34654), .Z(n34820) );
  XNOR U35464 ( .A(n34819), .B(n34820), .Z(n34763) );
  XNOR U35465 ( .A(n34764), .B(n34763), .Z(n34766) );
  NANDN U35466 ( .A(n34657), .B(n34656), .Z(n34661) );
  NANDN U35467 ( .A(n34659), .B(n34658), .Z(n34660) );
  AND U35468 ( .A(n34661), .B(n34660), .Z(n34765) );
  XOR U35469 ( .A(n34766), .B(n34765), .Z(n34880) );
  NANDN U35470 ( .A(n34663), .B(n34662), .Z(n34667) );
  NANDN U35471 ( .A(n34665), .B(n34664), .Z(n34666) );
  AND U35472 ( .A(n34667), .B(n34666), .Z(n34877) );
  NANDN U35473 ( .A(n34669), .B(n34668), .Z(n34673) );
  NANDN U35474 ( .A(n34671), .B(n34670), .Z(n34672) );
  AND U35475 ( .A(n34673), .B(n34672), .Z(n34760) );
  NANDN U35476 ( .A(n34675), .B(n34674), .Z(n34679) );
  OR U35477 ( .A(n34677), .B(n34676), .Z(n34678) );
  AND U35478 ( .A(n34679), .B(n34678), .Z(n34758) );
  NANDN U35479 ( .A(n34681), .B(n34680), .Z(n34685) );
  NANDN U35480 ( .A(n34683), .B(n34682), .Z(n34684) );
  AND U35481 ( .A(n34685), .B(n34684), .Z(n34824) );
  NANDN U35482 ( .A(n34687), .B(n34686), .Z(n34691) );
  NANDN U35483 ( .A(n34689), .B(n34688), .Z(n34690) );
  NAND U35484 ( .A(n34691), .B(n34690), .Z(n34823) );
  XNOR U35485 ( .A(n34824), .B(n34823), .Z(n34825) );
  NAND U35486 ( .A(n194), .B(n34692), .Z(n34694) );
  XOR U35487 ( .A(b[29]), .B(a[220]), .Z(n34850) );
  NAND U35488 ( .A(n38456), .B(n34850), .Z(n34693) );
  AND U35489 ( .A(n34694), .B(n34693), .Z(n34770) );
  AND U35490 ( .A(b[31]), .B(a[216]), .Z(n34769) );
  XNOR U35491 ( .A(n34770), .B(n34769), .Z(n34771) );
  NAND U35492 ( .A(b[0]), .B(a[248]), .Z(n34695) );
  XNOR U35493 ( .A(b[1]), .B(n34695), .Z(n34697) );
  NANDN U35494 ( .A(b[0]), .B(a[247]), .Z(n34696) );
  NAND U35495 ( .A(n34697), .B(n34696), .Z(n34772) );
  XNOR U35496 ( .A(n34771), .B(n34772), .Z(n34811) );
  NAND U35497 ( .A(n38185), .B(n34698), .Z(n34700) );
  XOR U35498 ( .A(b[23]), .B(a[226]), .Z(n34853) );
  NAND U35499 ( .A(n38132), .B(n34853), .Z(n34699) );
  AND U35500 ( .A(n34700), .B(n34699), .Z(n34844) );
  NAND U35501 ( .A(n184), .B(n34701), .Z(n34703) );
  XOR U35502 ( .A(a[242]), .B(b[7]), .Z(n34856) );
  NAND U35503 ( .A(n36592), .B(n34856), .Z(n34702) );
  AND U35504 ( .A(n34703), .B(n34702), .Z(n34842) );
  NAND U35505 ( .A(n38289), .B(n34704), .Z(n34706) );
  XOR U35506 ( .A(b[25]), .B(a[224]), .Z(n34859) );
  NAND U35507 ( .A(n38247), .B(n34859), .Z(n34705) );
  NAND U35508 ( .A(n34706), .B(n34705), .Z(n34841) );
  XNOR U35509 ( .A(n34842), .B(n34841), .Z(n34843) );
  XOR U35510 ( .A(n34844), .B(n34843), .Z(n34812) );
  XNOR U35511 ( .A(n34811), .B(n34812), .Z(n34813) );
  NAND U35512 ( .A(n187), .B(n34707), .Z(n34709) );
  XOR U35513 ( .A(b[13]), .B(a[236]), .Z(n34862) );
  NAND U35514 ( .A(n37295), .B(n34862), .Z(n34708) );
  AND U35515 ( .A(n34709), .B(n34708), .Z(n34806) );
  NAND U35516 ( .A(n186), .B(n34710), .Z(n34712) );
  XOR U35517 ( .A(a[238]), .B(b[11]), .Z(n34865) );
  NAND U35518 ( .A(n37097), .B(n34865), .Z(n34711) );
  NAND U35519 ( .A(n34712), .B(n34711), .Z(n34805) );
  XNOR U35520 ( .A(n34806), .B(n34805), .Z(n34807) );
  NAND U35521 ( .A(n188), .B(n34713), .Z(n34715) );
  XOR U35522 ( .A(b[15]), .B(a[234]), .Z(n34868) );
  NAND U35523 ( .A(n37382), .B(n34868), .Z(n34714) );
  AND U35524 ( .A(n34715), .B(n34714), .Z(n34802) );
  NAND U35525 ( .A(n38064), .B(n34716), .Z(n34718) );
  XOR U35526 ( .A(b[21]), .B(a[228]), .Z(n34871) );
  NAND U35527 ( .A(n37993), .B(n34871), .Z(n34717) );
  AND U35528 ( .A(n34718), .B(n34717), .Z(n34800) );
  NAND U35529 ( .A(n185), .B(n34719), .Z(n34721) );
  XOR U35530 ( .A(a[240]), .B(b[9]), .Z(n34874) );
  NAND U35531 ( .A(n36805), .B(n34874), .Z(n34720) );
  NAND U35532 ( .A(n34721), .B(n34720), .Z(n34799) );
  XNOR U35533 ( .A(n34800), .B(n34799), .Z(n34801) );
  XOR U35534 ( .A(n34802), .B(n34801), .Z(n34808) );
  XOR U35535 ( .A(n34807), .B(n34808), .Z(n34814) );
  XOR U35536 ( .A(n34813), .B(n34814), .Z(n34826) );
  XNOR U35537 ( .A(n34825), .B(n34826), .Z(n34757) );
  XNOR U35538 ( .A(n34758), .B(n34757), .Z(n34759) );
  XOR U35539 ( .A(n34760), .B(n34759), .Z(n34878) );
  XNOR U35540 ( .A(n34877), .B(n34878), .Z(n34879) );
  XNOR U35541 ( .A(n34880), .B(n34879), .Z(n34753) );
  XOR U35542 ( .A(n34754), .B(n34753), .Z(n34746) );
  NANDN U35543 ( .A(n34723), .B(n34722), .Z(n34727) );
  NANDN U35544 ( .A(n34725), .B(n34724), .Z(n34726) );
  AND U35545 ( .A(n34727), .B(n34726), .Z(n34745) );
  XNOR U35546 ( .A(n34746), .B(n34745), .Z(n34747) );
  NANDN U35547 ( .A(n34729), .B(n34728), .Z(n34733) );
  NAND U35548 ( .A(n34731), .B(n34730), .Z(n34732) );
  NAND U35549 ( .A(n34733), .B(n34732), .Z(n34748) );
  XNOR U35550 ( .A(n34747), .B(n34748), .Z(n34739) );
  XNOR U35551 ( .A(n34740), .B(n34739), .Z(n34741) );
  XNOR U35552 ( .A(n34742), .B(n34741), .Z(n34883) );
  XNOR U35553 ( .A(sreg[472]), .B(n34883), .Z(n34885) );
  NANDN U35554 ( .A(sreg[471]), .B(n34734), .Z(n34738) );
  NAND U35555 ( .A(n34736), .B(n34735), .Z(n34737) );
  NAND U35556 ( .A(n34738), .B(n34737), .Z(n34884) );
  XNOR U35557 ( .A(n34885), .B(n34884), .Z(c[472]) );
  NANDN U35558 ( .A(n34740), .B(n34739), .Z(n34744) );
  NANDN U35559 ( .A(n34742), .B(n34741), .Z(n34743) );
  AND U35560 ( .A(n34744), .B(n34743), .Z(n34891) );
  NANDN U35561 ( .A(n34746), .B(n34745), .Z(n34750) );
  NANDN U35562 ( .A(n34748), .B(n34747), .Z(n34749) );
  AND U35563 ( .A(n34750), .B(n34749), .Z(n34889) );
  NANDN U35564 ( .A(n34752), .B(n34751), .Z(n34756) );
  NAND U35565 ( .A(n34754), .B(n34753), .Z(n34755) );
  AND U35566 ( .A(n34756), .B(n34755), .Z(n34896) );
  NANDN U35567 ( .A(n34758), .B(n34757), .Z(n34762) );
  NANDN U35568 ( .A(n34760), .B(n34759), .Z(n34761) );
  AND U35569 ( .A(n34762), .B(n34761), .Z(n34901) );
  NANDN U35570 ( .A(n34764), .B(n34763), .Z(n34768) );
  NAND U35571 ( .A(n34766), .B(n34765), .Z(n34767) );
  AND U35572 ( .A(n34768), .B(n34767), .Z(n34900) );
  XNOR U35573 ( .A(n34901), .B(n34900), .Z(n34903) );
  NANDN U35574 ( .A(n34770), .B(n34769), .Z(n34774) );
  NANDN U35575 ( .A(n34772), .B(n34771), .Z(n34773) );
  AND U35576 ( .A(n34774), .B(n34773), .Z(n34980) );
  NAND U35577 ( .A(n38385), .B(n34775), .Z(n34777) );
  XOR U35578 ( .A(b[27]), .B(a[223]), .Z(n34924) );
  NAND U35579 ( .A(n38343), .B(n34924), .Z(n34776) );
  AND U35580 ( .A(n34777), .B(n34776), .Z(n34987) );
  NAND U35581 ( .A(n183), .B(n34778), .Z(n34780) );
  XOR U35582 ( .A(a[245]), .B(b[5]), .Z(n34927) );
  NAND U35583 ( .A(n36296), .B(n34927), .Z(n34779) );
  AND U35584 ( .A(n34780), .B(n34779), .Z(n34985) );
  NAND U35585 ( .A(n190), .B(n34781), .Z(n34783) );
  XOR U35586 ( .A(b[19]), .B(a[231]), .Z(n34930) );
  NAND U35587 ( .A(n37821), .B(n34930), .Z(n34782) );
  NAND U35588 ( .A(n34783), .B(n34782), .Z(n34984) );
  XNOR U35589 ( .A(n34985), .B(n34984), .Z(n34986) );
  XNOR U35590 ( .A(n34987), .B(n34986), .Z(n34978) );
  NAND U35591 ( .A(n38470), .B(n34784), .Z(n34786) );
  XOR U35592 ( .A(b[31]), .B(a[219]), .Z(n34933) );
  NAND U35593 ( .A(n38453), .B(n34933), .Z(n34785) );
  AND U35594 ( .A(n34786), .B(n34785), .Z(n34945) );
  NAND U35595 ( .A(n181), .B(n34787), .Z(n34789) );
  XOR U35596 ( .A(a[247]), .B(b[3]), .Z(n34936) );
  NAND U35597 ( .A(n182), .B(n34936), .Z(n34788) );
  AND U35598 ( .A(n34789), .B(n34788), .Z(n34943) );
  NAND U35599 ( .A(n189), .B(n34790), .Z(n34792) );
  XOR U35600 ( .A(b[17]), .B(a[233]), .Z(n34939) );
  NAND U35601 ( .A(n37652), .B(n34939), .Z(n34791) );
  NAND U35602 ( .A(n34792), .B(n34791), .Z(n34942) );
  XNOR U35603 ( .A(n34943), .B(n34942), .Z(n34944) );
  XOR U35604 ( .A(n34945), .B(n34944), .Z(n34979) );
  XOR U35605 ( .A(n34978), .B(n34979), .Z(n34981) );
  XOR U35606 ( .A(n34980), .B(n34981), .Z(n34913) );
  NANDN U35607 ( .A(n34794), .B(n34793), .Z(n34798) );
  NANDN U35608 ( .A(n34796), .B(n34795), .Z(n34797) );
  AND U35609 ( .A(n34798), .B(n34797), .Z(n34966) );
  NANDN U35610 ( .A(n34800), .B(n34799), .Z(n34804) );
  NANDN U35611 ( .A(n34802), .B(n34801), .Z(n34803) );
  NAND U35612 ( .A(n34804), .B(n34803), .Z(n34967) );
  XNOR U35613 ( .A(n34966), .B(n34967), .Z(n34968) );
  NANDN U35614 ( .A(n34806), .B(n34805), .Z(n34810) );
  NANDN U35615 ( .A(n34808), .B(n34807), .Z(n34809) );
  NAND U35616 ( .A(n34810), .B(n34809), .Z(n34969) );
  XNOR U35617 ( .A(n34968), .B(n34969), .Z(n34912) );
  XNOR U35618 ( .A(n34913), .B(n34912), .Z(n34915) );
  NANDN U35619 ( .A(n34812), .B(n34811), .Z(n34816) );
  NANDN U35620 ( .A(n34814), .B(n34813), .Z(n34815) );
  AND U35621 ( .A(n34816), .B(n34815), .Z(n34914) );
  XOR U35622 ( .A(n34915), .B(n34914), .Z(n35029) );
  NANDN U35623 ( .A(n34818), .B(n34817), .Z(n34822) );
  NANDN U35624 ( .A(n34820), .B(n34819), .Z(n34821) );
  AND U35625 ( .A(n34822), .B(n34821), .Z(n35026) );
  NANDN U35626 ( .A(n34824), .B(n34823), .Z(n34828) );
  NANDN U35627 ( .A(n34826), .B(n34825), .Z(n34827) );
  AND U35628 ( .A(n34828), .B(n34827), .Z(n34909) );
  NANDN U35629 ( .A(n34830), .B(n34829), .Z(n34834) );
  OR U35630 ( .A(n34832), .B(n34831), .Z(n34833) );
  AND U35631 ( .A(n34834), .B(n34833), .Z(n34907) );
  NANDN U35632 ( .A(n34836), .B(n34835), .Z(n34840) );
  NANDN U35633 ( .A(n34838), .B(n34837), .Z(n34839) );
  AND U35634 ( .A(n34840), .B(n34839), .Z(n34973) );
  NANDN U35635 ( .A(n34842), .B(n34841), .Z(n34846) );
  NANDN U35636 ( .A(n34844), .B(n34843), .Z(n34845) );
  NAND U35637 ( .A(n34846), .B(n34845), .Z(n34972) );
  XNOR U35638 ( .A(n34973), .B(n34972), .Z(n34974) );
  NAND U35639 ( .A(b[0]), .B(a[249]), .Z(n34847) );
  XNOR U35640 ( .A(b[1]), .B(n34847), .Z(n34849) );
  NANDN U35641 ( .A(b[0]), .B(a[248]), .Z(n34848) );
  NAND U35642 ( .A(n34849), .B(n34848), .Z(n34921) );
  NAND U35643 ( .A(n194), .B(n34850), .Z(n34852) );
  XOR U35644 ( .A(b[29]), .B(a[221]), .Z(n34996) );
  NAND U35645 ( .A(n38456), .B(n34996), .Z(n34851) );
  AND U35646 ( .A(n34852), .B(n34851), .Z(n34919) );
  AND U35647 ( .A(b[31]), .B(a[217]), .Z(n34918) );
  XNOR U35648 ( .A(n34919), .B(n34918), .Z(n34920) );
  XNOR U35649 ( .A(n34921), .B(n34920), .Z(n34960) );
  NAND U35650 ( .A(n38185), .B(n34853), .Z(n34855) );
  XOR U35651 ( .A(b[23]), .B(a[227]), .Z(n35002) );
  NAND U35652 ( .A(n38132), .B(n35002), .Z(n34854) );
  AND U35653 ( .A(n34855), .B(n34854), .Z(n34993) );
  NAND U35654 ( .A(n184), .B(n34856), .Z(n34858) );
  XOR U35655 ( .A(a[243]), .B(b[7]), .Z(n35005) );
  NAND U35656 ( .A(n36592), .B(n35005), .Z(n34857) );
  AND U35657 ( .A(n34858), .B(n34857), .Z(n34991) );
  NAND U35658 ( .A(n38289), .B(n34859), .Z(n34861) );
  XOR U35659 ( .A(b[25]), .B(a[225]), .Z(n35008) );
  NAND U35660 ( .A(n38247), .B(n35008), .Z(n34860) );
  NAND U35661 ( .A(n34861), .B(n34860), .Z(n34990) );
  XNOR U35662 ( .A(n34991), .B(n34990), .Z(n34992) );
  XOR U35663 ( .A(n34993), .B(n34992), .Z(n34961) );
  XNOR U35664 ( .A(n34960), .B(n34961), .Z(n34962) );
  NAND U35665 ( .A(n187), .B(n34862), .Z(n34864) );
  XOR U35666 ( .A(b[13]), .B(a[237]), .Z(n35011) );
  NAND U35667 ( .A(n37295), .B(n35011), .Z(n34863) );
  AND U35668 ( .A(n34864), .B(n34863), .Z(n34955) );
  NAND U35669 ( .A(n186), .B(n34865), .Z(n34867) );
  XOR U35670 ( .A(a[239]), .B(b[11]), .Z(n35014) );
  NAND U35671 ( .A(n37097), .B(n35014), .Z(n34866) );
  NAND U35672 ( .A(n34867), .B(n34866), .Z(n34954) );
  XNOR U35673 ( .A(n34955), .B(n34954), .Z(n34956) );
  NAND U35674 ( .A(n188), .B(n34868), .Z(n34870) );
  XOR U35675 ( .A(b[15]), .B(a[235]), .Z(n35017) );
  NAND U35676 ( .A(n37382), .B(n35017), .Z(n34869) );
  AND U35677 ( .A(n34870), .B(n34869), .Z(n34951) );
  NAND U35678 ( .A(n38064), .B(n34871), .Z(n34873) );
  XOR U35679 ( .A(b[21]), .B(a[229]), .Z(n35020) );
  NAND U35680 ( .A(n37993), .B(n35020), .Z(n34872) );
  AND U35681 ( .A(n34873), .B(n34872), .Z(n34949) );
  NAND U35682 ( .A(n185), .B(n34874), .Z(n34876) );
  XOR U35683 ( .A(a[241]), .B(b[9]), .Z(n35023) );
  NAND U35684 ( .A(n36805), .B(n35023), .Z(n34875) );
  NAND U35685 ( .A(n34876), .B(n34875), .Z(n34948) );
  XNOR U35686 ( .A(n34949), .B(n34948), .Z(n34950) );
  XOR U35687 ( .A(n34951), .B(n34950), .Z(n34957) );
  XOR U35688 ( .A(n34956), .B(n34957), .Z(n34963) );
  XOR U35689 ( .A(n34962), .B(n34963), .Z(n34975) );
  XNOR U35690 ( .A(n34974), .B(n34975), .Z(n34906) );
  XNOR U35691 ( .A(n34907), .B(n34906), .Z(n34908) );
  XOR U35692 ( .A(n34909), .B(n34908), .Z(n35027) );
  XNOR U35693 ( .A(n35026), .B(n35027), .Z(n35028) );
  XNOR U35694 ( .A(n35029), .B(n35028), .Z(n34902) );
  XOR U35695 ( .A(n34903), .B(n34902), .Z(n34895) );
  NANDN U35696 ( .A(n34878), .B(n34877), .Z(n34882) );
  NANDN U35697 ( .A(n34880), .B(n34879), .Z(n34881) );
  AND U35698 ( .A(n34882), .B(n34881), .Z(n34894) );
  XOR U35699 ( .A(n34895), .B(n34894), .Z(n34897) );
  XNOR U35700 ( .A(n34896), .B(n34897), .Z(n34888) );
  XNOR U35701 ( .A(n34889), .B(n34888), .Z(n34890) );
  XNOR U35702 ( .A(n34891), .B(n34890), .Z(n35032) );
  XNOR U35703 ( .A(sreg[473]), .B(n35032), .Z(n35034) );
  NANDN U35704 ( .A(sreg[472]), .B(n34883), .Z(n34887) );
  NAND U35705 ( .A(n34885), .B(n34884), .Z(n34886) );
  NAND U35706 ( .A(n34887), .B(n34886), .Z(n35033) );
  XNOR U35707 ( .A(n35034), .B(n35033), .Z(c[473]) );
  NANDN U35708 ( .A(n34889), .B(n34888), .Z(n34893) );
  NANDN U35709 ( .A(n34891), .B(n34890), .Z(n34892) );
  AND U35710 ( .A(n34893), .B(n34892), .Z(n35040) );
  NANDN U35711 ( .A(n34895), .B(n34894), .Z(n34899) );
  NANDN U35712 ( .A(n34897), .B(n34896), .Z(n34898) );
  AND U35713 ( .A(n34899), .B(n34898), .Z(n35038) );
  NANDN U35714 ( .A(n34901), .B(n34900), .Z(n34905) );
  NAND U35715 ( .A(n34903), .B(n34902), .Z(n34904) );
  AND U35716 ( .A(n34905), .B(n34904), .Z(n35045) );
  NANDN U35717 ( .A(n34907), .B(n34906), .Z(n34911) );
  NANDN U35718 ( .A(n34909), .B(n34908), .Z(n34910) );
  AND U35719 ( .A(n34911), .B(n34910), .Z(n35176) );
  NANDN U35720 ( .A(n34913), .B(n34912), .Z(n34917) );
  NAND U35721 ( .A(n34915), .B(n34914), .Z(n34916) );
  AND U35722 ( .A(n34917), .B(n34916), .Z(n35175) );
  XNOR U35723 ( .A(n35176), .B(n35175), .Z(n35178) );
  NANDN U35724 ( .A(n34919), .B(n34918), .Z(n34923) );
  NANDN U35725 ( .A(n34921), .B(n34920), .Z(n34922) );
  AND U35726 ( .A(n34923), .B(n34922), .Z(n35123) );
  NAND U35727 ( .A(n38385), .B(n34924), .Z(n34926) );
  XOR U35728 ( .A(b[27]), .B(a[224]), .Z(n35067) );
  NAND U35729 ( .A(n38343), .B(n35067), .Z(n34925) );
  AND U35730 ( .A(n34926), .B(n34925), .Z(n35130) );
  NAND U35731 ( .A(n183), .B(n34927), .Z(n34929) );
  XOR U35732 ( .A(a[246]), .B(b[5]), .Z(n35070) );
  NAND U35733 ( .A(n36296), .B(n35070), .Z(n34928) );
  AND U35734 ( .A(n34929), .B(n34928), .Z(n35128) );
  NAND U35735 ( .A(n190), .B(n34930), .Z(n34932) );
  XOR U35736 ( .A(b[19]), .B(a[232]), .Z(n35073) );
  NAND U35737 ( .A(n37821), .B(n35073), .Z(n34931) );
  NAND U35738 ( .A(n34932), .B(n34931), .Z(n35127) );
  XNOR U35739 ( .A(n35128), .B(n35127), .Z(n35129) );
  XNOR U35740 ( .A(n35130), .B(n35129), .Z(n35121) );
  NAND U35741 ( .A(n38470), .B(n34933), .Z(n34935) );
  XOR U35742 ( .A(b[31]), .B(a[220]), .Z(n35076) );
  NAND U35743 ( .A(n38453), .B(n35076), .Z(n34934) );
  AND U35744 ( .A(n34935), .B(n34934), .Z(n35088) );
  NAND U35745 ( .A(n181), .B(n34936), .Z(n34938) );
  XOR U35746 ( .A(a[248]), .B(b[3]), .Z(n35079) );
  NAND U35747 ( .A(n182), .B(n35079), .Z(n34937) );
  AND U35748 ( .A(n34938), .B(n34937), .Z(n35086) );
  NAND U35749 ( .A(n189), .B(n34939), .Z(n34941) );
  XOR U35750 ( .A(b[17]), .B(a[234]), .Z(n35082) );
  NAND U35751 ( .A(n37652), .B(n35082), .Z(n34940) );
  NAND U35752 ( .A(n34941), .B(n34940), .Z(n35085) );
  XNOR U35753 ( .A(n35086), .B(n35085), .Z(n35087) );
  XOR U35754 ( .A(n35088), .B(n35087), .Z(n35122) );
  XOR U35755 ( .A(n35121), .B(n35122), .Z(n35124) );
  XOR U35756 ( .A(n35123), .B(n35124), .Z(n35056) );
  NANDN U35757 ( .A(n34943), .B(n34942), .Z(n34947) );
  NANDN U35758 ( .A(n34945), .B(n34944), .Z(n34946) );
  AND U35759 ( .A(n34947), .B(n34946), .Z(n35109) );
  NANDN U35760 ( .A(n34949), .B(n34948), .Z(n34953) );
  NANDN U35761 ( .A(n34951), .B(n34950), .Z(n34952) );
  NAND U35762 ( .A(n34953), .B(n34952), .Z(n35110) );
  XNOR U35763 ( .A(n35109), .B(n35110), .Z(n35111) );
  NANDN U35764 ( .A(n34955), .B(n34954), .Z(n34959) );
  NANDN U35765 ( .A(n34957), .B(n34956), .Z(n34958) );
  NAND U35766 ( .A(n34959), .B(n34958), .Z(n35112) );
  XNOR U35767 ( .A(n35111), .B(n35112), .Z(n35055) );
  XNOR U35768 ( .A(n35056), .B(n35055), .Z(n35058) );
  NANDN U35769 ( .A(n34961), .B(n34960), .Z(n34965) );
  NANDN U35770 ( .A(n34963), .B(n34962), .Z(n34964) );
  AND U35771 ( .A(n34965), .B(n34964), .Z(n35057) );
  XOR U35772 ( .A(n35058), .B(n35057), .Z(n35172) );
  NANDN U35773 ( .A(n34967), .B(n34966), .Z(n34971) );
  NANDN U35774 ( .A(n34969), .B(n34968), .Z(n34970) );
  AND U35775 ( .A(n34971), .B(n34970), .Z(n35169) );
  NANDN U35776 ( .A(n34973), .B(n34972), .Z(n34977) );
  NANDN U35777 ( .A(n34975), .B(n34974), .Z(n34976) );
  AND U35778 ( .A(n34977), .B(n34976), .Z(n35052) );
  NANDN U35779 ( .A(n34979), .B(n34978), .Z(n34983) );
  OR U35780 ( .A(n34981), .B(n34980), .Z(n34982) );
  AND U35781 ( .A(n34983), .B(n34982), .Z(n35050) );
  NANDN U35782 ( .A(n34985), .B(n34984), .Z(n34989) );
  NANDN U35783 ( .A(n34987), .B(n34986), .Z(n34988) );
  AND U35784 ( .A(n34989), .B(n34988), .Z(n35116) );
  NANDN U35785 ( .A(n34991), .B(n34990), .Z(n34995) );
  NANDN U35786 ( .A(n34993), .B(n34992), .Z(n34994) );
  NAND U35787 ( .A(n34995), .B(n34994), .Z(n35115) );
  XNOR U35788 ( .A(n35116), .B(n35115), .Z(n35117) );
  NAND U35789 ( .A(n194), .B(n34996), .Z(n34998) );
  XOR U35790 ( .A(b[29]), .B(a[222]), .Z(n35142) );
  NAND U35791 ( .A(n38456), .B(n35142), .Z(n34997) );
  AND U35792 ( .A(n34998), .B(n34997), .Z(n35062) );
  AND U35793 ( .A(b[31]), .B(a[218]), .Z(n35061) );
  XNOR U35794 ( .A(n35062), .B(n35061), .Z(n35063) );
  NAND U35795 ( .A(b[0]), .B(a[250]), .Z(n34999) );
  XNOR U35796 ( .A(b[1]), .B(n34999), .Z(n35001) );
  NANDN U35797 ( .A(b[0]), .B(a[249]), .Z(n35000) );
  NAND U35798 ( .A(n35001), .B(n35000), .Z(n35064) );
  XNOR U35799 ( .A(n35063), .B(n35064), .Z(n35103) );
  NAND U35800 ( .A(n38185), .B(n35002), .Z(n35004) );
  XOR U35801 ( .A(b[23]), .B(a[228]), .Z(n35145) );
  NAND U35802 ( .A(n38132), .B(n35145), .Z(n35003) );
  AND U35803 ( .A(n35004), .B(n35003), .Z(n35136) );
  NAND U35804 ( .A(n184), .B(n35005), .Z(n35007) );
  XOR U35805 ( .A(a[244]), .B(b[7]), .Z(n35148) );
  NAND U35806 ( .A(n36592), .B(n35148), .Z(n35006) );
  AND U35807 ( .A(n35007), .B(n35006), .Z(n35134) );
  NAND U35808 ( .A(n38289), .B(n35008), .Z(n35010) );
  XOR U35809 ( .A(b[25]), .B(a[226]), .Z(n35151) );
  NAND U35810 ( .A(n38247), .B(n35151), .Z(n35009) );
  NAND U35811 ( .A(n35010), .B(n35009), .Z(n35133) );
  XNOR U35812 ( .A(n35134), .B(n35133), .Z(n35135) );
  XOR U35813 ( .A(n35136), .B(n35135), .Z(n35104) );
  XNOR U35814 ( .A(n35103), .B(n35104), .Z(n35105) );
  NAND U35815 ( .A(n187), .B(n35011), .Z(n35013) );
  XOR U35816 ( .A(b[13]), .B(a[238]), .Z(n35154) );
  NAND U35817 ( .A(n37295), .B(n35154), .Z(n35012) );
  AND U35818 ( .A(n35013), .B(n35012), .Z(n35098) );
  NAND U35819 ( .A(n186), .B(n35014), .Z(n35016) );
  XOR U35820 ( .A(a[240]), .B(b[11]), .Z(n35157) );
  NAND U35821 ( .A(n37097), .B(n35157), .Z(n35015) );
  NAND U35822 ( .A(n35016), .B(n35015), .Z(n35097) );
  XNOR U35823 ( .A(n35098), .B(n35097), .Z(n35099) );
  NAND U35824 ( .A(n188), .B(n35017), .Z(n35019) );
  XOR U35825 ( .A(b[15]), .B(a[236]), .Z(n35160) );
  NAND U35826 ( .A(n37382), .B(n35160), .Z(n35018) );
  AND U35827 ( .A(n35019), .B(n35018), .Z(n35094) );
  NAND U35828 ( .A(n38064), .B(n35020), .Z(n35022) );
  XOR U35829 ( .A(b[21]), .B(a[230]), .Z(n35163) );
  NAND U35830 ( .A(n37993), .B(n35163), .Z(n35021) );
  AND U35831 ( .A(n35022), .B(n35021), .Z(n35092) );
  NAND U35832 ( .A(n185), .B(n35023), .Z(n35025) );
  XOR U35833 ( .A(a[242]), .B(b[9]), .Z(n35166) );
  NAND U35834 ( .A(n36805), .B(n35166), .Z(n35024) );
  NAND U35835 ( .A(n35025), .B(n35024), .Z(n35091) );
  XNOR U35836 ( .A(n35092), .B(n35091), .Z(n35093) );
  XOR U35837 ( .A(n35094), .B(n35093), .Z(n35100) );
  XOR U35838 ( .A(n35099), .B(n35100), .Z(n35106) );
  XOR U35839 ( .A(n35105), .B(n35106), .Z(n35118) );
  XNOR U35840 ( .A(n35117), .B(n35118), .Z(n35049) );
  XNOR U35841 ( .A(n35050), .B(n35049), .Z(n35051) );
  XOR U35842 ( .A(n35052), .B(n35051), .Z(n35170) );
  XNOR U35843 ( .A(n35169), .B(n35170), .Z(n35171) );
  XNOR U35844 ( .A(n35172), .B(n35171), .Z(n35177) );
  XOR U35845 ( .A(n35178), .B(n35177), .Z(n35044) );
  NANDN U35846 ( .A(n35027), .B(n35026), .Z(n35031) );
  NANDN U35847 ( .A(n35029), .B(n35028), .Z(n35030) );
  AND U35848 ( .A(n35031), .B(n35030), .Z(n35043) );
  XOR U35849 ( .A(n35044), .B(n35043), .Z(n35046) );
  XNOR U35850 ( .A(n35045), .B(n35046), .Z(n35037) );
  XNOR U35851 ( .A(n35038), .B(n35037), .Z(n35039) );
  XNOR U35852 ( .A(n35040), .B(n35039), .Z(n35181) );
  XNOR U35853 ( .A(sreg[474]), .B(n35181), .Z(n35183) );
  NANDN U35854 ( .A(sreg[473]), .B(n35032), .Z(n35036) );
  NAND U35855 ( .A(n35034), .B(n35033), .Z(n35035) );
  NAND U35856 ( .A(n35036), .B(n35035), .Z(n35182) );
  XNOR U35857 ( .A(n35183), .B(n35182), .Z(c[474]) );
  NANDN U35858 ( .A(n35038), .B(n35037), .Z(n35042) );
  NANDN U35859 ( .A(n35040), .B(n35039), .Z(n35041) );
  AND U35860 ( .A(n35042), .B(n35041), .Z(n35189) );
  NANDN U35861 ( .A(n35044), .B(n35043), .Z(n35048) );
  NANDN U35862 ( .A(n35046), .B(n35045), .Z(n35047) );
  AND U35863 ( .A(n35048), .B(n35047), .Z(n35187) );
  NANDN U35864 ( .A(n35050), .B(n35049), .Z(n35054) );
  NANDN U35865 ( .A(n35052), .B(n35051), .Z(n35053) );
  AND U35866 ( .A(n35054), .B(n35053), .Z(n35325) );
  NANDN U35867 ( .A(n35056), .B(n35055), .Z(n35060) );
  NAND U35868 ( .A(n35058), .B(n35057), .Z(n35059) );
  AND U35869 ( .A(n35060), .B(n35059), .Z(n35324) );
  XNOR U35870 ( .A(n35325), .B(n35324), .Z(n35327) );
  NANDN U35871 ( .A(n35062), .B(n35061), .Z(n35066) );
  NANDN U35872 ( .A(n35064), .B(n35063), .Z(n35065) );
  AND U35873 ( .A(n35066), .B(n35065), .Z(n35272) );
  NAND U35874 ( .A(n38385), .B(n35067), .Z(n35069) );
  XOR U35875 ( .A(b[27]), .B(a[225]), .Z(n35216) );
  NAND U35876 ( .A(n38343), .B(n35216), .Z(n35068) );
  AND U35877 ( .A(n35069), .B(n35068), .Z(n35279) );
  NAND U35878 ( .A(n183), .B(n35070), .Z(n35072) );
  XOR U35879 ( .A(a[247]), .B(b[5]), .Z(n35219) );
  NAND U35880 ( .A(n36296), .B(n35219), .Z(n35071) );
  AND U35881 ( .A(n35072), .B(n35071), .Z(n35277) );
  NAND U35882 ( .A(n190), .B(n35073), .Z(n35075) );
  XOR U35883 ( .A(b[19]), .B(a[233]), .Z(n35222) );
  NAND U35884 ( .A(n37821), .B(n35222), .Z(n35074) );
  NAND U35885 ( .A(n35075), .B(n35074), .Z(n35276) );
  XNOR U35886 ( .A(n35277), .B(n35276), .Z(n35278) );
  XNOR U35887 ( .A(n35279), .B(n35278), .Z(n35270) );
  NAND U35888 ( .A(n38470), .B(n35076), .Z(n35078) );
  XOR U35889 ( .A(b[31]), .B(a[221]), .Z(n35225) );
  NAND U35890 ( .A(n38453), .B(n35225), .Z(n35077) );
  AND U35891 ( .A(n35078), .B(n35077), .Z(n35237) );
  NAND U35892 ( .A(n181), .B(n35079), .Z(n35081) );
  XOR U35893 ( .A(a[249]), .B(b[3]), .Z(n35228) );
  NAND U35894 ( .A(n182), .B(n35228), .Z(n35080) );
  AND U35895 ( .A(n35081), .B(n35080), .Z(n35235) );
  NAND U35896 ( .A(n189), .B(n35082), .Z(n35084) );
  XOR U35897 ( .A(b[17]), .B(a[235]), .Z(n35231) );
  NAND U35898 ( .A(n37652), .B(n35231), .Z(n35083) );
  NAND U35899 ( .A(n35084), .B(n35083), .Z(n35234) );
  XNOR U35900 ( .A(n35235), .B(n35234), .Z(n35236) );
  XOR U35901 ( .A(n35237), .B(n35236), .Z(n35271) );
  XOR U35902 ( .A(n35270), .B(n35271), .Z(n35273) );
  XOR U35903 ( .A(n35272), .B(n35273), .Z(n35205) );
  NANDN U35904 ( .A(n35086), .B(n35085), .Z(n35090) );
  NANDN U35905 ( .A(n35088), .B(n35087), .Z(n35089) );
  AND U35906 ( .A(n35090), .B(n35089), .Z(n35258) );
  NANDN U35907 ( .A(n35092), .B(n35091), .Z(n35096) );
  NANDN U35908 ( .A(n35094), .B(n35093), .Z(n35095) );
  NAND U35909 ( .A(n35096), .B(n35095), .Z(n35259) );
  XNOR U35910 ( .A(n35258), .B(n35259), .Z(n35260) );
  NANDN U35911 ( .A(n35098), .B(n35097), .Z(n35102) );
  NANDN U35912 ( .A(n35100), .B(n35099), .Z(n35101) );
  NAND U35913 ( .A(n35102), .B(n35101), .Z(n35261) );
  XNOR U35914 ( .A(n35260), .B(n35261), .Z(n35204) );
  XNOR U35915 ( .A(n35205), .B(n35204), .Z(n35207) );
  NANDN U35916 ( .A(n35104), .B(n35103), .Z(n35108) );
  NANDN U35917 ( .A(n35106), .B(n35105), .Z(n35107) );
  AND U35918 ( .A(n35108), .B(n35107), .Z(n35206) );
  XOR U35919 ( .A(n35207), .B(n35206), .Z(n35321) );
  NANDN U35920 ( .A(n35110), .B(n35109), .Z(n35114) );
  NANDN U35921 ( .A(n35112), .B(n35111), .Z(n35113) );
  AND U35922 ( .A(n35114), .B(n35113), .Z(n35318) );
  NANDN U35923 ( .A(n35116), .B(n35115), .Z(n35120) );
  NANDN U35924 ( .A(n35118), .B(n35117), .Z(n35119) );
  AND U35925 ( .A(n35120), .B(n35119), .Z(n35201) );
  NANDN U35926 ( .A(n35122), .B(n35121), .Z(n35126) );
  OR U35927 ( .A(n35124), .B(n35123), .Z(n35125) );
  AND U35928 ( .A(n35126), .B(n35125), .Z(n35199) );
  NANDN U35929 ( .A(n35128), .B(n35127), .Z(n35132) );
  NANDN U35930 ( .A(n35130), .B(n35129), .Z(n35131) );
  AND U35931 ( .A(n35132), .B(n35131), .Z(n35265) );
  NANDN U35932 ( .A(n35134), .B(n35133), .Z(n35138) );
  NANDN U35933 ( .A(n35136), .B(n35135), .Z(n35137) );
  NAND U35934 ( .A(n35138), .B(n35137), .Z(n35264) );
  XNOR U35935 ( .A(n35265), .B(n35264), .Z(n35266) );
  NAND U35936 ( .A(b[0]), .B(a[251]), .Z(n35139) );
  XNOR U35937 ( .A(b[1]), .B(n35139), .Z(n35141) );
  NANDN U35938 ( .A(b[0]), .B(a[250]), .Z(n35140) );
  NAND U35939 ( .A(n35141), .B(n35140), .Z(n35213) );
  NAND U35940 ( .A(n194), .B(n35142), .Z(n35144) );
  XOR U35941 ( .A(b[29]), .B(a[223]), .Z(n35291) );
  NAND U35942 ( .A(n38456), .B(n35291), .Z(n35143) );
  AND U35943 ( .A(n35144), .B(n35143), .Z(n35211) );
  AND U35944 ( .A(b[31]), .B(a[219]), .Z(n35210) );
  XNOR U35945 ( .A(n35211), .B(n35210), .Z(n35212) );
  XNOR U35946 ( .A(n35213), .B(n35212), .Z(n35252) );
  NAND U35947 ( .A(n38185), .B(n35145), .Z(n35147) );
  XOR U35948 ( .A(b[23]), .B(a[229]), .Z(n35294) );
  NAND U35949 ( .A(n38132), .B(n35294), .Z(n35146) );
  AND U35950 ( .A(n35147), .B(n35146), .Z(n35285) );
  NAND U35951 ( .A(n184), .B(n35148), .Z(n35150) );
  XOR U35952 ( .A(a[245]), .B(b[7]), .Z(n35297) );
  NAND U35953 ( .A(n36592), .B(n35297), .Z(n35149) );
  AND U35954 ( .A(n35150), .B(n35149), .Z(n35283) );
  NAND U35955 ( .A(n38289), .B(n35151), .Z(n35153) );
  XOR U35956 ( .A(b[25]), .B(a[227]), .Z(n35300) );
  NAND U35957 ( .A(n38247), .B(n35300), .Z(n35152) );
  NAND U35958 ( .A(n35153), .B(n35152), .Z(n35282) );
  XNOR U35959 ( .A(n35283), .B(n35282), .Z(n35284) );
  XOR U35960 ( .A(n35285), .B(n35284), .Z(n35253) );
  XNOR U35961 ( .A(n35252), .B(n35253), .Z(n35254) );
  NAND U35962 ( .A(n187), .B(n35154), .Z(n35156) );
  XOR U35963 ( .A(b[13]), .B(a[239]), .Z(n35303) );
  NAND U35964 ( .A(n37295), .B(n35303), .Z(n35155) );
  AND U35965 ( .A(n35156), .B(n35155), .Z(n35247) );
  NAND U35966 ( .A(n186), .B(n35157), .Z(n35159) );
  XOR U35967 ( .A(a[241]), .B(b[11]), .Z(n35306) );
  NAND U35968 ( .A(n37097), .B(n35306), .Z(n35158) );
  NAND U35969 ( .A(n35159), .B(n35158), .Z(n35246) );
  XNOR U35970 ( .A(n35247), .B(n35246), .Z(n35248) );
  NAND U35971 ( .A(n188), .B(n35160), .Z(n35162) );
  XOR U35972 ( .A(b[15]), .B(a[237]), .Z(n35309) );
  NAND U35973 ( .A(n37382), .B(n35309), .Z(n35161) );
  AND U35974 ( .A(n35162), .B(n35161), .Z(n35243) );
  NAND U35975 ( .A(n38064), .B(n35163), .Z(n35165) );
  XOR U35976 ( .A(b[21]), .B(a[231]), .Z(n35312) );
  NAND U35977 ( .A(n37993), .B(n35312), .Z(n35164) );
  AND U35978 ( .A(n35165), .B(n35164), .Z(n35241) );
  NAND U35979 ( .A(n185), .B(n35166), .Z(n35168) );
  XOR U35980 ( .A(a[243]), .B(b[9]), .Z(n35315) );
  NAND U35981 ( .A(n36805), .B(n35315), .Z(n35167) );
  NAND U35982 ( .A(n35168), .B(n35167), .Z(n35240) );
  XNOR U35983 ( .A(n35241), .B(n35240), .Z(n35242) );
  XOR U35984 ( .A(n35243), .B(n35242), .Z(n35249) );
  XOR U35985 ( .A(n35248), .B(n35249), .Z(n35255) );
  XOR U35986 ( .A(n35254), .B(n35255), .Z(n35267) );
  XNOR U35987 ( .A(n35266), .B(n35267), .Z(n35198) );
  XNOR U35988 ( .A(n35199), .B(n35198), .Z(n35200) );
  XOR U35989 ( .A(n35201), .B(n35200), .Z(n35319) );
  XNOR U35990 ( .A(n35318), .B(n35319), .Z(n35320) );
  XNOR U35991 ( .A(n35321), .B(n35320), .Z(n35326) );
  XOR U35992 ( .A(n35327), .B(n35326), .Z(n35193) );
  NANDN U35993 ( .A(n35170), .B(n35169), .Z(n35174) );
  NANDN U35994 ( .A(n35172), .B(n35171), .Z(n35173) );
  AND U35995 ( .A(n35174), .B(n35173), .Z(n35192) );
  XNOR U35996 ( .A(n35193), .B(n35192), .Z(n35194) );
  NANDN U35997 ( .A(n35176), .B(n35175), .Z(n35180) );
  NAND U35998 ( .A(n35178), .B(n35177), .Z(n35179) );
  NAND U35999 ( .A(n35180), .B(n35179), .Z(n35195) );
  XNOR U36000 ( .A(n35194), .B(n35195), .Z(n35186) );
  XNOR U36001 ( .A(n35187), .B(n35186), .Z(n35188) );
  XNOR U36002 ( .A(n35189), .B(n35188), .Z(n35330) );
  XNOR U36003 ( .A(sreg[475]), .B(n35330), .Z(n35332) );
  NANDN U36004 ( .A(sreg[474]), .B(n35181), .Z(n35185) );
  NAND U36005 ( .A(n35183), .B(n35182), .Z(n35184) );
  NAND U36006 ( .A(n35185), .B(n35184), .Z(n35331) );
  XNOR U36007 ( .A(n35332), .B(n35331), .Z(c[475]) );
  NANDN U36008 ( .A(n35187), .B(n35186), .Z(n35191) );
  NANDN U36009 ( .A(n35189), .B(n35188), .Z(n35190) );
  AND U36010 ( .A(n35191), .B(n35190), .Z(n35338) );
  NANDN U36011 ( .A(n35193), .B(n35192), .Z(n35197) );
  NANDN U36012 ( .A(n35195), .B(n35194), .Z(n35196) );
  AND U36013 ( .A(n35197), .B(n35196), .Z(n35336) );
  NANDN U36014 ( .A(n35199), .B(n35198), .Z(n35203) );
  NANDN U36015 ( .A(n35201), .B(n35200), .Z(n35202) );
  AND U36016 ( .A(n35203), .B(n35202), .Z(n35342) );
  NANDN U36017 ( .A(n35205), .B(n35204), .Z(n35209) );
  NAND U36018 ( .A(n35207), .B(n35206), .Z(n35208) );
  AND U36019 ( .A(n35209), .B(n35208), .Z(n35341) );
  XNOR U36020 ( .A(n35342), .B(n35341), .Z(n35344) );
  NANDN U36021 ( .A(n35211), .B(n35210), .Z(n35215) );
  NANDN U36022 ( .A(n35213), .B(n35212), .Z(n35214) );
  AND U36023 ( .A(n35215), .B(n35214), .Z(n35428) );
  NAND U36024 ( .A(n38385), .B(n35216), .Z(n35218) );
  XOR U36025 ( .A(b[27]), .B(a[226]), .Z(n35371) );
  NAND U36026 ( .A(n38343), .B(n35371), .Z(n35217) );
  NAND U36027 ( .A(n35218), .B(n35217), .Z(n35470) );
  NAND U36028 ( .A(n183), .B(n35219), .Z(n35221) );
  XOR U36029 ( .A(a[248]), .B(b[5]), .Z(n35374) );
  NAND U36030 ( .A(n36296), .B(n35374), .Z(n35220) );
  NAND U36031 ( .A(n35221), .B(n35220), .Z(n35468) );
  NAND U36032 ( .A(n190), .B(n35222), .Z(n35224) );
  XOR U36033 ( .A(b[19]), .B(a[234]), .Z(n35377) );
  NAND U36034 ( .A(n37821), .B(n35377), .Z(n35223) );
  NAND U36035 ( .A(n35224), .B(n35223), .Z(n35467) );
  NAND U36036 ( .A(n38470), .B(n35225), .Z(n35227) );
  XOR U36037 ( .A(b[31]), .B(a[222]), .Z(n35380) );
  NAND U36038 ( .A(n38453), .B(n35380), .Z(n35226) );
  NAND U36039 ( .A(n35227), .B(n35226), .Z(n35392) );
  NAND U36040 ( .A(n181), .B(n35228), .Z(n35230) );
  XOR U36041 ( .A(a[250]), .B(b[3]), .Z(n35383) );
  NAND U36042 ( .A(n182), .B(n35383), .Z(n35229) );
  NAND U36043 ( .A(n35230), .B(n35229), .Z(n35390) );
  NAND U36044 ( .A(n189), .B(n35231), .Z(n35233) );
  XOR U36045 ( .A(b[17]), .B(a[236]), .Z(n35386) );
  NAND U36046 ( .A(n37652), .B(n35386), .Z(n35232) );
  NAND U36047 ( .A(n35233), .B(n35232), .Z(n35389) );
  XOR U36048 ( .A(n35425), .B(n35426), .Z(n35427) );
  XOR U36049 ( .A(n35428), .B(n35427), .Z(n35360) );
  NANDN U36050 ( .A(n35235), .B(n35234), .Z(n35239) );
  NANDN U36051 ( .A(n35237), .B(n35236), .Z(n35238) );
  AND U36052 ( .A(n35239), .B(n35238), .Z(n35413) );
  NANDN U36053 ( .A(n35241), .B(n35240), .Z(n35245) );
  NANDN U36054 ( .A(n35243), .B(n35242), .Z(n35244) );
  NAND U36055 ( .A(n35245), .B(n35244), .Z(n35414) );
  XNOR U36056 ( .A(n35413), .B(n35414), .Z(n35415) );
  NANDN U36057 ( .A(n35247), .B(n35246), .Z(n35251) );
  NANDN U36058 ( .A(n35249), .B(n35248), .Z(n35250) );
  NAND U36059 ( .A(n35251), .B(n35250), .Z(n35416) );
  XNOR U36060 ( .A(n35415), .B(n35416), .Z(n35359) );
  XOR U36061 ( .A(n35360), .B(n35359), .Z(n35362) );
  NANDN U36062 ( .A(n35253), .B(n35252), .Z(n35257) );
  NANDN U36063 ( .A(n35255), .B(n35254), .Z(n35256) );
  AND U36064 ( .A(n35257), .B(n35256), .Z(n35361) );
  XOR U36065 ( .A(n35362), .B(n35361), .Z(n35350) );
  NANDN U36066 ( .A(n35259), .B(n35258), .Z(n35263) );
  NANDN U36067 ( .A(n35261), .B(n35260), .Z(n35262) );
  AND U36068 ( .A(n35263), .B(n35262), .Z(n35347) );
  NANDN U36069 ( .A(n35265), .B(n35264), .Z(n35269) );
  NANDN U36070 ( .A(n35267), .B(n35266), .Z(n35268) );
  AND U36071 ( .A(n35269), .B(n35268), .Z(n35356) );
  NANDN U36072 ( .A(n35271), .B(n35270), .Z(n35275) );
  OR U36073 ( .A(n35273), .B(n35272), .Z(n35274) );
  AND U36074 ( .A(n35275), .B(n35274), .Z(n35354) );
  NANDN U36075 ( .A(n35277), .B(n35276), .Z(n35281) );
  NANDN U36076 ( .A(n35279), .B(n35278), .Z(n35280) );
  AND U36077 ( .A(n35281), .B(n35280), .Z(n35420) );
  NANDN U36078 ( .A(n35283), .B(n35282), .Z(n35287) );
  NANDN U36079 ( .A(n35285), .B(n35284), .Z(n35286) );
  NAND U36080 ( .A(n35287), .B(n35286), .Z(n35419) );
  XNOR U36081 ( .A(n35420), .B(n35419), .Z(n35421) );
  NAND U36082 ( .A(b[0]), .B(a[252]), .Z(n35288) );
  XNOR U36083 ( .A(b[1]), .B(n35288), .Z(n35290) );
  NANDN U36084 ( .A(b[0]), .B(a[251]), .Z(n35289) );
  NAND U36085 ( .A(n35290), .B(n35289), .Z(n35368) );
  NAND U36086 ( .A(n194), .B(n35291), .Z(n35293) );
  XOR U36087 ( .A(b[29]), .B(a[224]), .Z(n35458) );
  NAND U36088 ( .A(n38456), .B(n35458), .Z(n35292) );
  NAND U36089 ( .A(n35293), .B(n35292), .Z(n35366) );
  AND U36090 ( .A(b[31]), .B(a[220]), .Z(n35365) );
  XNOR U36091 ( .A(n35368), .B(n35367), .Z(n35407) );
  NAND U36092 ( .A(n38185), .B(n35294), .Z(n35296) );
  XOR U36093 ( .A(b[23]), .B(a[230]), .Z(n35446) );
  NAND U36094 ( .A(n38132), .B(n35446), .Z(n35295) );
  NAND U36095 ( .A(n35296), .B(n35295), .Z(n35464) );
  NAND U36096 ( .A(n184), .B(n35297), .Z(n35299) );
  XOR U36097 ( .A(a[246]), .B(b[7]), .Z(n35449) );
  NAND U36098 ( .A(n36592), .B(n35449), .Z(n35298) );
  NAND U36099 ( .A(n35299), .B(n35298), .Z(n35462) );
  NAND U36100 ( .A(n38289), .B(n35300), .Z(n35302) );
  XOR U36101 ( .A(b[25]), .B(a[228]), .Z(n35452) );
  NAND U36102 ( .A(n38247), .B(n35452), .Z(n35301) );
  NAND U36103 ( .A(n35302), .B(n35301), .Z(n35461) );
  XNOR U36104 ( .A(n35407), .B(n35408), .Z(n35410) );
  NAND U36105 ( .A(n187), .B(n35303), .Z(n35305) );
  XOR U36106 ( .A(a[240]), .B(b[13]), .Z(n35431) );
  NAND U36107 ( .A(n37295), .B(n35431), .Z(n35304) );
  NAND U36108 ( .A(n35305), .B(n35304), .Z(n35402) );
  NAND U36109 ( .A(n186), .B(n35306), .Z(n35308) );
  XOR U36110 ( .A(a[242]), .B(b[11]), .Z(n35434) );
  NAND U36111 ( .A(n37097), .B(n35434), .Z(n35307) );
  NAND U36112 ( .A(n35308), .B(n35307), .Z(n35401) );
  NAND U36113 ( .A(n188), .B(n35309), .Z(n35311) );
  XOR U36114 ( .A(b[15]), .B(a[238]), .Z(n35437) );
  NAND U36115 ( .A(n37382), .B(n35437), .Z(n35310) );
  NAND U36116 ( .A(n35311), .B(n35310), .Z(n35398) );
  NAND U36117 ( .A(n38064), .B(n35312), .Z(n35314) );
  XOR U36118 ( .A(b[21]), .B(a[232]), .Z(n35440) );
  NAND U36119 ( .A(n37993), .B(n35440), .Z(n35313) );
  NAND U36120 ( .A(n35314), .B(n35313), .Z(n35396) );
  NAND U36121 ( .A(n185), .B(n35315), .Z(n35317) );
  XOR U36122 ( .A(a[244]), .B(b[9]), .Z(n35443) );
  NAND U36123 ( .A(n36805), .B(n35443), .Z(n35316) );
  NAND U36124 ( .A(n35317), .B(n35316), .Z(n35395) );
  XOR U36125 ( .A(n35404), .B(n35403), .Z(n35409) );
  XOR U36126 ( .A(n35410), .B(n35409), .Z(n35422) );
  XOR U36127 ( .A(n35421), .B(n35422), .Z(n35353) );
  XNOR U36128 ( .A(n35354), .B(n35353), .Z(n35355) );
  XOR U36129 ( .A(n35356), .B(n35355), .Z(n35348) );
  XNOR U36130 ( .A(n35347), .B(n35348), .Z(n35349) );
  XNOR U36131 ( .A(n35350), .B(n35349), .Z(n35343) );
  XOR U36132 ( .A(n35344), .B(n35343), .Z(n35474) );
  NANDN U36133 ( .A(n35319), .B(n35318), .Z(n35323) );
  NANDN U36134 ( .A(n35321), .B(n35320), .Z(n35322) );
  AND U36135 ( .A(n35323), .B(n35322), .Z(n35473) );
  XNOR U36136 ( .A(n35474), .B(n35473), .Z(n35475) );
  NANDN U36137 ( .A(n35325), .B(n35324), .Z(n35329) );
  NAND U36138 ( .A(n35327), .B(n35326), .Z(n35328) );
  NAND U36139 ( .A(n35329), .B(n35328), .Z(n35476) );
  XNOR U36140 ( .A(n35475), .B(n35476), .Z(n35335) );
  XNOR U36141 ( .A(n35336), .B(n35335), .Z(n35337) );
  XNOR U36142 ( .A(n35338), .B(n35337), .Z(n35479) );
  XNOR U36143 ( .A(sreg[476]), .B(n35479), .Z(n35481) );
  NANDN U36144 ( .A(sreg[475]), .B(n35330), .Z(n35334) );
  NAND U36145 ( .A(n35332), .B(n35331), .Z(n35333) );
  NAND U36146 ( .A(n35334), .B(n35333), .Z(n35480) );
  XNOR U36147 ( .A(n35481), .B(n35480), .Z(c[476]) );
  NANDN U36148 ( .A(n35336), .B(n35335), .Z(n35340) );
  NANDN U36149 ( .A(n35338), .B(n35337), .Z(n35339) );
  AND U36150 ( .A(n35340), .B(n35339), .Z(n35487) );
  NANDN U36151 ( .A(n35342), .B(n35341), .Z(n35346) );
  NAND U36152 ( .A(n35344), .B(n35343), .Z(n35345) );
  AND U36153 ( .A(n35346), .B(n35345), .Z(n35624) );
  NANDN U36154 ( .A(n35348), .B(n35347), .Z(n35352) );
  NANDN U36155 ( .A(n35350), .B(n35349), .Z(n35351) );
  AND U36156 ( .A(n35352), .B(n35351), .Z(n35623) );
  NANDN U36157 ( .A(n35354), .B(n35353), .Z(n35358) );
  NANDN U36158 ( .A(n35356), .B(n35355), .Z(n35357) );
  AND U36159 ( .A(n35358), .B(n35357), .Z(n35617) );
  NAND U36160 ( .A(n35360), .B(n35359), .Z(n35364) );
  NAND U36161 ( .A(n35362), .B(n35361), .Z(n35363) );
  AND U36162 ( .A(n35364), .B(n35363), .Z(n35616) );
  XNOR U36163 ( .A(n35617), .B(n35616), .Z(n35618) );
  NAND U36164 ( .A(n35366), .B(n35365), .Z(n35370) );
  NANDN U36165 ( .A(n35368), .B(n35367), .Z(n35369) );
  NAND U36166 ( .A(n35370), .B(n35369), .Z(n35553) );
  NAND U36167 ( .A(n38385), .B(n35371), .Z(n35373) );
  XOR U36168 ( .A(b[27]), .B(a[227]), .Z(n35508) );
  NAND U36169 ( .A(n38343), .B(n35508), .Z(n35372) );
  NAND U36170 ( .A(n35373), .B(n35372), .Z(n35589) );
  NAND U36171 ( .A(n183), .B(n35374), .Z(n35376) );
  XOR U36172 ( .A(a[249]), .B(b[5]), .Z(n35511) );
  NAND U36173 ( .A(n36296), .B(n35511), .Z(n35375) );
  NAND U36174 ( .A(n35376), .B(n35375), .Z(n35587) );
  NAND U36175 ( .A(n190), .B(n35377), .Z(n35379) );
  XOR U36176 ( .A(b[19]), .B(a[235]), .Z(n35514) );
  NAND U36177 ( .A(n37821), .B(n35514), .Z(n35378) );
  NAND U36178 ( .A(n35379), .B(n35378), .Z(n35586) );
  NAND U36179 ( .A(n38470), .B(n35380), .Z(n35382) );
  XOR U36180 ( .A(b[31]), .B(a[223]), .Z(n35517) );
  NAND U36181 ( .A(n38453), .B(n35517), .Z(n35381) );
  NAND U36182 ( .A(n35382), .B(n35381), .Z(n35535) );
  NAND U36183 ( .A(n181), .B(n35383), .Z(n35385) );
  XOR U36184 ( .A(a[251]), .B(b[3]), .Z(n35520) );
  NAND U36185 ( .A(n182), .B(n35520), .Z(n35384) );
  NAND U36186 ( .A(n35385), .B(n35384), .Z(n35533) );
  NAND U36187 ( .A(n189), .B(n35386), .Z(n35388) );
  XOR U36188 ( .A(b[17]), .B(a[237]), .Z(n35523) );
  NAND U36189 ( .A(n37652), .B(n35523), .Z(n35387) );
  NAND U36190 ( .A(n35388), .B(n35387), .Z(n35532) );
  XOR U36191 ( .A(n35551), .B(n35550), .Z(n35552) );
  NAND U36192 ( .A(n35390), .B(n35389), .Z(n35394) );
  NAND U36193 ( .A(n35392), .B(n35391), .Z(n35393) );
  AND U36194 ( .A(n35394), .B(n35393), .Z(n35598) );
  NAND U36195 ( .A(n35396), .B(n35395), .Z(n35400) );
  NAND U36196 ( .A(n35398), .B(n35397), .Z(n35399) );
  AND U36197 ( .A(n35400), .B(n35399), .Z(n35599) );
  NAND U36198 ( .A(n35402), .B(n35401), .Z(n35406) );
  NAND U36199 ( .A(n35404), .B(n35403), .Z(n35405) );
  AND U36200 ( .A(n35406), .B(n35405), .Z(n35601) );
  XOR U36201 ( .A(n35604), .B(n35605), .Z(n35607) );
  NANDN U36202 ( .A(n35408), .B(n35407), .Z(n35412) );
  NAND U36203 ( .A(n35410), .B(n35409), .Z(n35411) );
  AND U36204 ( .A(n35412), .B(n35411), .Z(n35606) );
  XOR U36205 ( .A(n35607), .B(n35606), .Z(n35493) );
  NANDN U36206 ( .A(n35414), .B(n35413), .Z(n35418) );
  NANDN U36207 ( .A(n35416), .B(n35415), .Z(n35417) );
  AND U36208 ( .A(n35418), .B(n35417), .Z(n35490) );
  NANDN U36209 ( .A(n35420), .B(n35419), .Z(n35424) );
  NAND U36210 ( .A(n35422), .B(n35421), .Z(n35423) );
  NAND U36211 ( .A(n35424), .B(n35423), .Z(n35613) );
  NAND U36212 ( .A(n35426), .B(n35425), .Z(n35430) );
  NANDN U36213 ( .A(n35428), .B(n35427), .Z(n35429) );
  NAND U36214 ( .A(n35430), .B(n35429), .Z(n35611) );
  NAND U36215 ( .A(n187), .B(n35431), .Z(n35433) );
  XOR U36216 ( .A(a[241]), .B(b[13]), .Z(n35556) );
  NAND U36217 ( .A(n37295), .B(n35556), .Z(n35432) );
  NAND U36218 ( .A(n35433), .B(n35432), .Z(n35541) );
  NAND U36219 ( .A(n186), .B(n35434), .Z(n35436) );
  XOR U36220 ( .A(a[243]), .B(b[11]), .Z(n35559) );
  NAND U36221 ( .A(n37097), .B(n35559), .Z(n35435) );
  NAND U36222 ( .A(n35436), .B(n35435), .Z(n35539) );
  NAND U36223 ( .A(n188), .B(n35437), .Z(n35439) );
  XOR U36224 ( .A(b[15]), .B(a[239]), .Z(n35562) );
  NAND U36225 ( .A(n37382), .B(n35562), .Z(n35438) );
  NAND U36226 ( .A(n35439), .B(n35438), .Z(n35529) );
  NAND U36227 ( .A(n38064), .B(n35440), .Z(n35442) );
  XOR U36228 ( .A(b[21]), .B(a[233]), .Z(n35565) );
  NAND U36229 ( .A(n37993), .B(n35565), .Z(n35441) );
  NAND U36230 ( .A(n35442), .B(n35441), .Z(n35527) );
  NAND U36231 ( .A(n185), .B(n35443), .Z(n35445) );
  XOR U36232 ( .A(a[245]), .B(b[9]), .Z(n35568) );
  NAND U36233 ( .A(n36805), .B(n35568), .Z(n35444) );
  NAND U36234 ( .A(n35445), .B(n35444), .Z(n35526) );
  NAND U36235 ( .A(n38185), .B(n35446), .Z(n35448) );
  XOR U36236 ( .A(b[23]), .B(a[231]), .Z(n35571) );
  NAND U36237 ( .A(n38132), .B(n35571), .Z(n35447) );
  NAND U36238 ( .A(n35448), .B(n35447), .Z(n35595) );
  NAND U36239 ( .A(n184), .B(n35449), .Z(n35451) );
  XOR U36240 ( .A(a[247]), .B(b[7]), .Z(n35574) );
  NAND U36241 ( .A(n36592), .B(n35574), .Z(n35450) );
  NAND U36242 ( .A(n35451), .B(n35450), .Z(n35593) );
  NAND U36243 ( .A(n38289), .B(n35452), .Z(n35454) );
  XOR U36244 ( .A(b[25]), .B(a[229]), .Z(n35577) );
  NAND U36245 ( .A(n38247), .B(n35577), .Z(n35453) );
  NAND U36246 ( .A(n35454), .B(n35453), .Z(n35592) );
  NAND U36247 ( .A(b[0]), .B(a[253]), .Z(n35455) );
  XNOR U36248 ( .A(b[1]), .B(n35455), .Z(n35457) );
  NANDN U36249 ( .A(b[0]), .B(a[252]), .Z(n35456) );
  NAND U36250 ( .A(n35457), .B(n35456), .Z(n35505) );
  NAND U36251 ( .A(n194), .B(n35458), .Z(n35460) );
  XOR U36252 ( .A(b[29]), .B(a[225]), .Z(n35583) );
  NAND U36253 ( .A(n38456), .B(n35583), .Z(n35459) );
  NAND U36254 ( .A(n35460), .B(n35459), .Z(n35503) );
  AND U36255 ( .A(b[31]), .B(a[221]), .Z(n35502) );
  XOR U36256 ( .A(n35505), .B(n35504), .Z(n35496) );
  XOR U36257 ( .A(n35497), .B(n35496), .Z(n35499) );
  XNOR U36258 ( .A(n35498), .B(n35499), .Z(n35546) );
  NAND U36259 ( .A(n35462), .B(n35461), .Z(n35466) );
  NAND U36260 ( .A(n35464), .B(n35463), .Z(n35465) );
  NAND U36261 ( .A(n35466), .B(n35465), .Z(n35545) );
  NAND U36262 ( .A(n35468), .B(n35467), .Z(n35472) );
  NAND U36263 ( .A(n35470), .B(n35469), .Z(n35471) );
  NAND U36264 ( .A(n35472), .B(n35471), .Z(n35544) );
  XOR U36265 ( .A(n35546), .B(n35547), .Z(n35610) );
  XOR U36266 ( .A(n35490), .B(n35491), .Z(n35492) );
  XOR U36267 ( .A(n35493), .B(n35492), .Z(n35619) );
  XNOR U36268 ( .A(n35618), .B(n35619), .Z(n35622) );
  XOR U36269 ( .A(n35623), .B(n35622), .Z(n35625) );
  XOR U36270 ( .A(n35624), .B(n35625), .Z(n35485) );
  NANDN U36271 ( .A(n35474), .B(n35473), .Z(n35478) );
  NANDN U36272 ( .A(n35476), .B(n35475), .Z(n35477) );
  NAND U36273 ( .A(n35478), .B(n35477), .Z(n35484) );
  XNOR U36274 ( .A(n35485), .B(n35484), .Z(n35486) );
  XNOR U36275 ( .A(n35487), .B(n35486), .Z(n35628) );
  XNOR U36276 ( .A(sreg[477]), .B(n35628), .Z(n35630) );
  NANDN U36277 ( .A(sreg[476]), .B(n35479), .Z(n35483) );
  NAND U36278 ( .A(n35481), .B(n35480), .Z(n35482) );
  NAND U36279 ( .A(n35483), .B(n35482), .Z(n35629) );
  XNOR U36280 ( .A(n35630), .B(n35629), .Z(c[477]) );
  NANDN U36281 ( .A(n35485), .B(n35484), .Z(n35489) );
  NANDN U36282 ( .A(n35487), .B(n35486), .Z(n35488) );
  AND U36283 ( .A(n35489), .B(n35488), .Z(n35636) );
  NAND U36284 ( .A(n35491), .B(n35490), .Z(n35495) );
  NANDN U36285 ( .A(n35493), .B(n35492), .Z(n35494) );
  AND U36286 ( .A(n35495), .B(n35494), .Z(n35772) );
  NAND U36287 ( .A(n35497), .B(n35496), .Z(n35501) );
  NAND U36288 ( .A(n35499), .B(n35498), .Z(n35500) );
  NAND U36289 ( .A(n35501), .B(n35500), .Z(n35768) );
  NAND U36290 ( .A(n35503), .B(n35502), .Z(n35507) );
  NANDN U36291 ( .A(n35505), .B(n35504), .Z(n35506) );
  NAND U36292 ( .A(n35507), .B(n35506), .Z(n35708) );
  NAND U36293 ( .A(n38385), .B(n35508), .Z(n35510) );
  XOR U36294 ( .A(b[27]), .B(a[228]), .Z(n35684) );
  NAND U36295 ( .A(n38343), .B(n35684), .Z(n35509) );
  NAND U36296 ( .A(n35510), .B(n35509), .Z(n35750) );
  NAND U36297 ( .A(n183), .B(n35511), .Z(n35513) );
  XOR U36298 ( .A(a[250]), .B(b[5]), .Z(n35687) );
  NAND U36299 ( .A(n36296), .B(n35687), .Z(n35512) );
  NAND U36300 ( .A(n35513), .B(n35512), .Z(n35748) );
  NAND U36301 ( .A(n190), .B(n35514), .Z(n35516) );
  XOR U36302 ( .A(b[19]), .B(a[236]), .Z(n35690) );
  NAND U36303 ( .A(n37821), .B(n35690), .Z(n35515) );
  NAND U36304 ( .A(n35516), .B(n35515), .Z(n35747) );
  NAND U36305 ( .A(n38470), .B(n35517), .Z(n35519) );
  XOR U36306 ( .A(b[31]), .B(a[224]), .Z(n35675) );
  NAND U36307 ( .A(n38453), .B(n35675), .Z(n35518) );
  NAND U36308 ( .A(n35519), .B(n35518), .Z(n35666) );
  NAND U36309 ( .A(n181), .B(n35520), .Z(n35522) );
  XOR U36310 ( .A(a[252]), .B(b[3]), .Z(n35678) );
  NAND U36311 ( .A(n182), .B(n35678), .Z(n35521) );
  NAND U36312 ( .A(n35522), .B(n35521), .Z(n35664) );
  NAND U36313 ( .A(n189), .B(n35523), .Z(n35525) );
  XOR U36314 ( .A(b[17]), .B(a[238]), .Z(n35681) );
  NAND U36315 ( .A(n37652), .B(n35681), .Z(n35524) );
  NAND U36316 ( .A(n35525), .B(n35524), .Z(n35663) );
  XOR U36317 ( .A(n35706), .B(n35705), .Z(n35707) );
  NAND U36318 ( .A(n35527), .B(n35526), .Z(n35531) );
  NAND U36319 ( .A(n35529), .B(n35528), .Z(n35530) );
  AND U36320 ( .A(n35531), .B(n35530), .Z(n35753) );
  NAND U36321 ( .A(n35533), .B(n35532), .Z(n35537) );
  NAND U36322 ( .A(n35535), .B(n35534), .Z(n35536) );
  AND U36323 ( .A(n35537), .B(n35536), .Z(n35754) );
  NAND U36324 ( .A(n35539), .B(n35538), .Z(n35543) );
  NAND U36325 ( .A(n35541), .B(n35540), .Z(n35542) );
  AND U36326 ( .A(n35543), .B(n35542), .Z(n35756) );
  XOR U36327 ( .A(n35765), .B(n35766), .Z(n35767) );
  NAND U36328 ( .A(n35545), .B(n35544), .Z(n35549) );
  NAND U36329 ( .A(n35547), .B(n35546), .Z(n35548) );
  NAND U36330 ( .A(n35549), .B(n35548), .Z(n35762) );
  NAND U36331 ( .A(n35551), .B(n35550), .Z(n35555) );
  NAND U36332 ( .A(n35553), .B(n35552), .Z(n35554) );
  NAND U36333 ( .A(n35555), .B(n35554), .Z(n35760) );
  NAND U36334 ( .A(n187), .B(n35556), .Z(n35558) );
  XOR U36335 ( .A(a[242]), .B(b[13]), .Z(n35711) );
  NAND U36336 ( .A(n37295), .B(n35711), .Z(n35557) );
  NAND U36337 ( .A(n35558), .B(n35557), .Z(n35672) );
  NAND U36338 ( .A(n186), .B(n35559), .Z(n35561) );
  XOR U36339 ( .A(a[244]), .B(b[11]), .Z(n35714) );
  NAND U36340 ( .A(n37097), .B(n35714), .Z(n35560) );
  NAND U36341 ( .A(n35561), .B(n35560), .Z(n35670) );
  NAND U36342 ( .A(n188), .B(n35562), .Z(n35564) );
  XOR U36343 ( .A(b[15]), .B(a[240]), .Z(n35717) );
  NAND U36344 ( .A(n37382), .B(n35717), .Z(n35563) );
  NAND U36345 ( .A(n35564), .B(n35563), .Z(n35660) );
  NAND U36346 ( .A(n38064), .B(n35565), .Z(n35567) );
  XOR U36347 ( .A(b[21]), .B(a[234]), .Z(n35720) );
  NAND U36348 ( .A(n37993), .B(n35720), .Z(n35566) );
  NAND U36349 ( .A(n35567), .B(n35566), .Z(n35658) );
  NAND U36350 ( .A(n185), .B(n35568), .Z(n35570) );
  XOR U36351 ( .A(a[246]), .B(b[9]), .Z(n35723) );
  NAND U36352 ( .A(n36805), .B(n35723), .Z(n35569) );
  NAND U36353 ( .A(n35570), .B(n35569), .Z(n35657) );
  XNOR U36354 ( .A(n35672), .B(n35671), .Z(n35653) );
  NAND U36355 ( .A(n38185), .B(n35571), .Z(n35573) );
  XOR U36356 ( .A(b[23]), .B(a[232]), .Z(n35726) );
  NAND U36357 ( .A(n38132), .B(n35726), .Z(n35572) );
  NAND U36358 ( .A(n35573), .B(n35572), .Z(n35744) );
  NAND U36359 ( .A(n184), .B(n35574), .Z(n35576) );
  XOR U36360 ( .A(a[248]), .B(b[7]), .Z(n35729) );
  NAND U36361 ( .A(n36592), .B(n35729), .Z(n35575) );
  NAND U36362 ( .A(n35576), .B(n35575), .Z(n35742) );
  NAND U36363 ( .A(n38289), .B(n35577), .Z(n35579) );
  XOR U36364 ( .A(b[25]), .B(a[230]), .Z(n35732) );
  NAND U36365 ( .A(n38247), .B(n35732), .Z(n35578) );
  NAND U36366 ( .A(n35579), .B(n35578), .Z(n35741) );
  NAND U36367 ( .A(b[0]), .B(a[254]), .Z(n35580) );
  XNOR U36368 ( .A(b[1]), .B(n35580), .Z(n35582) );
  NANDN U36369 ( .A(b[0]), .B(a[253]), .Z(n35581) );
  NAND U36370 ( .A(n35582), .B(n35581), .Z(n35696) );
  NAND U36371 ( .A(n194), .B(n35583), .Z(n35585) );
  XOR U36372 ( .A(b[29]), .B(a[226]), .Z(n35738) );
  NAND U36373 ( .A(n38456), .B(n35738), .Z(n35584) );
  NAND U36374 ( .A(n35585), .B(n35584), .Z(n35694) );
  AND U36375 ( .A(b[31]), .B(a[222]), .Z(n35693) );
  XOR U36376 ( .A(n35696), .B(n35695), .Z(n35651) );
  XOR U36377 ( .A(n35653), .B(n35654), .Z(n35701) );
  NAND U36378 ( .A(n35587), .B(n35586), .Z(n35591) );
  NAND U36379 ( .A(n35589), .B(n35588), .Z(n35590) );
  NAND U36380 ( .A(n35591), .B(n35590), .Z(n35700) );
  NAND U36381 ( .A(n35593), .B(n35592), .Z(n35597) );
  NAND U36382 ( .A(n35595), .B(n35594), .Z(n35596) );
  NAND U36383 ( .A(n35597), .B(n35596), .Z(n35699) );
  XOR U36384 ( .A(n35701), .B(n35702), .Z(n35759) );
  NAND U36385 ( .A(n35599), .B(n35598), .Z(n35603) );
  NAND U36386 ( .A(n35601), .B(n35600), .Z(n35602) );
  AND U36387 ( .A(n35603), .B(n35602), .Z(n35646) );
  XNOR U36388 ( .A(n35647), .B(n35648), .Z(n35641) );
  NAND U36389 ( .A(n35605), .B(n35604), .Z(n35609) );
  NAND U36390 ( .A(n35607), .B(n35606), .Z(n35608) );
  NAND U36391 ( .A(n35609), .B(n35608), .Z(n35640) );
  NAND U36392 ( .A(n35611), .B(n35610), .Z(n35615) );
  NAND U36393 ( .A(n35613), .B(n35612), .Z(n35614) );
  AND U36394 ( .A(n35615), .B(n35614), .Z(n35639) );
  XOR U36395 ( .A(n35641), .B(n35642), .Z(n35771) );
  XOR U36396 ( .A(n35772), .B(n35771), .Z(n35773) );
  NANDN U36397 ( .A(n35617), .B(n35616), .Z(n35621) );
  NANDN U36398 ( .A(n35619), .B(n35618), .Z(n35620) );
  AND U36399 ( .A(n35621), .B(n35620), .Z(n35774) );
  NANDN U36400 ( .A(n35623), .B(n35622), .Z(n35627) );
  OR U36401 ( .A(n35625), .B(n35624), .Z(n35626) );
  NAND U36402 ( .A(n35627), .B(n35626), .Z(n35634) );
  XNOR U36403 ( .A(n35633), .B(n35634), .Z(n35635) );
  XNOR U36404 ( .A(n35636), .B(n35635), .Z(n35777) );
  XNOR U36405 ( .A(sreg[478]), .B(n35777), .Z(n35779) );
  NANDN U36406 ( .A(sreg[477]), .B(n35628), .Z(n35632) );
  NAND U36407 ( .A(n35630), .B(n35629), .Z(n35631) );
  NAND U36408 ( .A(n35632), .B(n35631), .Z(n35778) );
  XNOR U36409 ( .A(n35779), .B(n35778), .Z(c[478]) );
  NANDN U36410 ( .A(n35634), .B(n35633), .Z(n35638) );
  NANDN U36411 ( .A(n35636), .B(n35635), .Z(n35637) );
  NAND U36412 ( .A(n35638), .B(n35637), .Z(n35790) );
  NAND U36413 ( .A(n35640), .B(n35639), .Z(n35644) );
  NAND U36414 ( .A(n35642), .B(n35641), .Z(n35643) );
  AND U36415 ( .A(n35644), .B(n35643), .Z(n35925) );
  NAND U36416 ( .A(n35646), .B(n35645), .Z(n35650) );
  NAND U36417 ( .A(n35648), .B(n35647), .Z(n35649) );
  NAND U36418 ( .A(n35650), .B(n35649), .Z(n35923) );
  NAND U36419 ( .A(n35652), .B(n35651), .Z(n35656) );
  NANDN U36420 ( .A(n35654), .B(n35653), .Z(n35655) );
  AND U36421 ( .A(n35656), .B(n35655), .Z(n35913) );
  NAND U36422 ( .A(n35658), .B(n35657), .Z(n35662) );
  NAND U36423 ( .A(n35660), .B(n35659), .Z(n35661) );
  AND U36424 ( .A(n35662), .B(n35661), .Z(n35799) );
  NAND U36425 ( .A(n35664), .B(n35663), .Z(n35668) );
  NAND U36426 ( .A(n35666), .B(n35665), .Z(n35667) );
  AND U36427 ( .A(n35668), .B(n35667), .Z(n35800) );
  NAND U36428 ( .A(n35670), .B(n35669), .Z(n35674) );
  NAND U36429 ( .A(n35672), .B(n35671), .Z(n35673) );
  AND U36430 ( .A(n35674), .B(n35673), .Z(n35801) );
  XNOR U36431 ( .A(n35802), .B(n35801), .Z(n35911) );
  NAND U36432 ( .A(n38470), .B(n35675), .Z(n35677) );
  XOR U36433 ( .A(b[31]), .B(a[225]), .Z(n35877) );
  NAND U36434 ( .A(n38453), .B(n35877), .Z(n35676) );
  NAND U36435 ( .A(n35677), .B(n35676), .Z(n35895) );
  NAND U36436 ( .A(n181), .B(n35678), .Z(n35680) );
  XOR U36437 ( .A(a[253]), .B(b[3]), .Z(n35880) );
  NAND U36438 ( .A(n182), .B(n35880), .Z(n35679) );
  NAND U36439 ( .A(n35680), .B(n35679), .Z(n35893) );
  NAND U36440 ( .A(n189), .B(n35681), .Z(n35683) );
  XOR U36441 ( .A(b[17]), .B(a[239]), .Z(n35883) );
  NAND U36442 ( .A(n37652), .B(n35883), .Z(n35682) );
  NAND U36443 ( .A(n35683), .B(n35682), .Z(n35892) );
  NAND U36444 ( .A(n38385), .B(n35684), .Z(n35686) );
  XOR U36445 ( .A(b[27]), .B(a[229]), .Z(n35868) );
  NAND U36446 ( .A(n38343), .B(n35868), .Z(n35685) );
  AND U36447 ( .A(n35686), .B(n35685), .Z(n35847) );
  NAND U36448 ( .A(n183), .B(n35687), .Z(n35689) );
  XOR U36449 ( .A(a[251]), .B(b[5]), .Z(n35871) );
  NAND U36450 ( .A(n36296), .B(n35871), .Z(n35688) );
  NAND U36451 ( .A(n35689), .B(n35688), .Z(n35845) );
  NAND U36452 ( .A(n190), .B(n35690), .Z(n35692) );
  XOR U36453 ( .A(b[19]), .B(a[237]), .Z(n35874) );
  NAND U36454 ( .A(n37821), .B(n35874), .Z(n35691) );
  NAND U36455 ( .A(n35692), .B(n35691), .Z(n35844) );
  XOR U36456 ( .A(n35847), .B(n35846), .Z(n35811) );
  XOR U36457 ( .A(n35812), .B(n35811), .Z(n35814) );
  NAND U36458 ( .A(n35694), .B(n35693), .Z(n35698) );
  NANDN U36459 ( .A(n35696), .B(n35695), .Z(n35697) );
  AND U36460 ( .A(n35698), .B(n35697), .Z(n35813) );
  XNOR U36461 ( .A(n35814), .B(n35813), .Z(n35910) );
  XNOR U36462 ( .A(n35913), .B(n35912), .Z(n35919) );
  NAND U36463 ( .A(n35700), .B(n35699), .Z(n35704) );
  NAND U36464 ( .A(n35702), .B(n35701), .Z(n35703) );
  NAND U36465 ( .A(n35704), .B(n35703), .Z(n35907) );
  NAND U36466 ( .A(n35706), .B(n35705), .Z(n35710) );
  NAND U36467 ( .A(n35708), .B(n35707), .Z(n35709) );
  NAND U36468 ( .A(n35710), .B(n35709), .Z(n35905) );
  NAND U36469 ( .A(n187), .B(n35711), .Z(n35713) );
  XOR U36470 ( .A(a[243]), .B(b[13]), .Z(n35832) );
  NAND U36471 ( .A(n37295), .B(n35832), .Z(n35712) );
  NAND U36472 ( .A(n35713), .B(n35712), .Z(n35901) );
  NAND U36473 ( .A(n186), .B(n35714), .Z(n35716) );
  XOR U36474 ( .A(a[245]), .B(b[11]), .Z(n35829) );
  NAND U36475 ( .A(n37097), .B(n35829), .Z(n35715) );
  NAND U36476 ( .A(n35716), .B(n35715), .Z(n35899) );
  NAND U36477 ( .A(n188), .B(n35717), .Z(n35719) );
  XOR U36478 ( .A(b[15]), .B(a[241]), .Z(n35835) );
  NAND U36479 ( .A(n37382), .B(n35835), .Z(n35718) );
  NAND U36480 ( .A(n35719), .B(n35718), .Z(n35889) );
  NAND U36481 ( .A(n38064), .B(n35720), .Z(n35722) );
  XOR U36482 ( .A(b[21]), .B(a[235]), .Z(n35838) );
  NAND U36483 ( .A(n37993), .B(n35838), .Z(n35721) );
  NAND U36484 ( .A(n35722), .B(n35721), .Z(n35887) );
  NAND U36485 ( .A(n185), .B(n35723), .Z(n35725) );
  XOR U36486 ( .A(a[247]), .B(b[9]), .Z(n35841) );
  NAND U36487 ( .A(n36805), .B(n35841), .Z(n35724) );
  NAND U36488 ( .A(n35725), .B(n35724), .Z(n35886) );
  NAND U36489 ( .A(n38185), .B(n35726), .Z(n35728) );
  XOR U36490 ( .A(b[23]), .B(a[233]), .Z(n35820) );
  NAND U36491 ( .A(n38132), .B(n35820), .Z(n35727) );
  NAND U36492 ( .A(n35728), .B(n35727), .Z(n35853) );
  NAND U36493 ( .A(n184), .B(n35729), .Z(n35731) );
  XOR U36494 ( .A(a[249]), .B(b[7]), .Z(n35823) );
  NAND U36495 ( .A(n36592), .B(n35823), .Z(n35730) );
  NAND U36496 ( .A(n35731), .B(n35730), .Z(n35851) );
  NAND U36497 ( .A(n38289), .B(n35732), .Z(n35734) );
  XOR U36498 ( .A(b[25]), .B(a[231]), .Z(n35826) );
  NAND U36499 ( .A(n38247), .B(n35826), .Z(n35733) );
  NAND U36500 ( .A(n35734), .B(n35733), .Z(n35850) );
  NAND U36501 ( .A(b[0]), .B(a[255]), .Z(n35735) );
  XNOR U36502 ( .A(b[1]), .B(n35735), .Z(n35737) );
  NANDN U36503 ( .A(b[0]), .B(a[254]), .Z(n35736) );
  NAND U36504 ( .A(n35737), .B(n35736), .Z(n35865) );
  NAND U36505 ( .A(n194), .B(n35738), .Z(n35740) );
  XOR U36506 ( .A(b[29]), .B(a[227]), .Z(n35817) );
  NAND U36507 ( .A(n38456), .B(n35817), .Z(n35739) );
  NAND U36508 ( .A(n35740), .B(n35739), .Z(n35863) );
  AND U36509 ( .A(b[31]), .B(a[223]), .Z(n35862) );
  XOR U36510 ( .A(n35865), .B(n35864), .Z(n35856) );
  XOR U36511 ( .A(n35857), .B(n35856), .Z(n35859) );
  XNOR U36512 ( .A(n35858), .B(n35859), .Z(n35807) );
  NAND U36513 ( .A(n35742), .B(n35741), .Z(n35746) );
  NAND U36514 ( .A(n35744), .B(n35743), .Z(n35745) );
  NAND U36515 ( .A(n35746), .B(n35745), .Z(n35806) );
  NAND U36516 ( .A(n35748), .B(n35747), .Z(n35752) );
  NAND U36517 ( .A(n35750), .B(n35749), .Z(n35751) );
  NAND U36518 ( .A(n35752), .B(n35751), .Z(n35805) );
  XOR U36519 ( .A(n35807), .B(n35808), .Z(n35904) );
  NAND U36520 ( .A(n35754), .B(n35753), .Z(n35758) );
  NAND U36521 ( .A(n35756), .B(n35755), .Z(n35757) );
  NAND U36522 ( .A(n35758), .B(n35757), .Z(n35916) );
  XOR U36523 ( .A(n35917), .B(n35916), .Z(n35918) );
  NAND U36524 ( .A(n35760), .B(n35759), .Z(n35764) );
  NAND U36525 ( .A(n35762), .B(n35761), .Z(n35763) );
  NAND U36526 ( .A(n35764), .B(n35763), .Z(n35794) );
  NAND U36527 ( .A(n35766), .B(n35765), .Z(n35770) );
  NAND U36528 ( .A(n35768), .B(n35767), .Z(n35769) );
  AND U36529 ( .A(n35770), .B(n35769), .Z(n35793) );
  XOR U36530 ( .A(n35795), .B(n35796), .Z(n35922) );
  XNOR U36531 ( .A(n35925), .B(n35924), .Z(n35788) );
  NAND U36532 ( .A(n35772), .B(n35771), .Z(n35776) );
  NAND U36533 ( .A(n35774), .B(n35773), .Z(n35775) );
  NAND U36534 ( .A(n35776), .B(n35775), .Z(n35787) );
  XNOR U36535 ( .A(sreg[479]), .B(n35782), .Z(n35784) );
  NANDN U36536 ( .A(sreg[478]), .B(n35777), .Z(n35781) );
  NAND U36537 ( .A(n35779), .B(n35778), .Z(n35780) );
  NAND U36538 ( .A(n35781), .B(n35780), .Z(n35783) );
  XNOR U36539 ( .A(n35784), .B(n35783), .Z(c[479]) );
  NANDN U36540 ( .A(sreg[479]), .B(n35782), .Z(n35786) );
  NAND U36541 ( .A(n35784), .B(n35783), .Z(n35785) );
  AND U36542 ( .A(n35786), .B(n35785), .Z(n35929) );
  NAND U36543 ( .A(n35788), .B(n35787), .Z(n35792) );
  NAND U36544 ( .A(n35790), .B(n35789), .Z(n35791) );
  AND U36545 ( .A(n35792), .B(n35791), .Z(n35933) );
  NAND U36546 ( .A(n35794), .B(n35793), .Z(n35798) );
  NAND U36547 ( .A(n35796), .B(n35795), .Z(n35797) );
  NAND U36548 ( .A(n35798), .B(n35797), .Z(n36068) );
  NAND U36549 ( .A(n35800), .B(n35799), .Z(n35804) );
  NAND U36550 ( .A(n35802), .B(n35801), .Z(n35803) );
  NAND U36551 ( .A(n35804), .B(n35803), .Z(n36060) );
  NAND U36552 ( .A(n35806), .B(n35805), .Z(n35810) );
  NAND U36553 ( .A(n35808), .B(n35807), .Z(n35809) );
  AND U36554 ( .A(n35810), .B(n35809), .Z(n35951) );
  NAND U36555 ( .A(n35812), .B(n35811), .Z(n35816) );
  NAND U36556 ( .A(n35814), .B(n35813), .Z(n35815) );
  NAND U36557 ( .A(n35816), .B(n35815), .Z(n35949) );
  NAND U36558 ( .A(n194), .B(n35817), .Z(n35819) );
  XOR U36559 ( .A(b[29]), .B(a[228]), .Z(n36032) );
  NAND U36560 ( .A(n38456), .B(n36032), .Z(n35818) );
  NAND U36561 ( .A(n35819), .B(n35818), .Z(n35979) );
  AND U36562 ( .A(b[31]), .B(a[224]), .Z(n35978) );
  NAND U36563 ( .A(n38185), .B(n35820), .Z(n35822) );
  XOR U36564 ( .A(b[23]), .B(a[234]), .Z(n36026) );
  NAND U36565 ( .A(n38132), .B(n36026), .Z(n35821) );
  AND U36566 ( .A(n35822), .B(n35821), .Z(n36038) );
  NAND U36567 ( .A(n184), .B(n35823), .Z(n35825) );
  XOR U36568 ( .A(a[250]), .B(b[7]), .Z(n36017) );
  NAND U36569 ( .A(n36592), .B(n36017), .Z(n35824) );
  NAND U36570 ( .A(n35825), .B(n35824), .Z(n36036) );
  NAND U36571 ( .A(n38289), .B(n35826), .Z(n35828) );
  XOR U36572 ( .A(b[25]), .B(a[232]), .Z(n35990) );
  NAND U36573 ( .A(n38247), .B(n35990), .Z(n35827) );
  NAND U36574 ( .A(n35828), .B(n35827), .Z(n36035) );
  XOR U36575 ( .A(n36038), .B(n36037), .Z(n35954) );
  XOR U36576 ( .A(n35955), .B(n35954), .Z(n35957) );
  NAND U36577 ( .A(n186), .B(n35829), .Z(n35831) );
  XOR U36578 ( .A(a[246]), .B(b[11]), .Z(n36008) );
  NAND U36579 ( .A(n37097), .B(n36008), .Z(n35830) );
  NAND U36580 ( .A(n35831), .B(n35830), .Z(n35975) );
  NAND U36581 ( .A(n187), .B(n35832), .Z(n35834) );
  XOR U36582 ( .A(a[244]), .B(b[13]), .Z(n36011) );
  NAND U36583 ( .A(n37295), .B(n36011), .Z(n35833) );
  NAND U36584 ( .A(n35834), .B(n35833), .Z(n35973) );
  NAND U36585 ( .A(n188), .B(n35835), .Z(n35837) );
  XOR U36586 ( .A(a[242]), .B(b[15]), .Z(n35987) );
  NAND U36587 ( .A(n37382), .B(n35987), .Z(n35836) );
  NAND U36588 ( .A(n35837), .B(n35836), .Z(n35963) );
  NAND U36589 ( .A(n38064), .B(n35838), .Z(n35840) );
  XOR U36590 ( .A(b[21]), .B(a[236]), .Z(n36020) );
  NAND U36591 ( .A(n37993), .B(n36020), .Z(n35839) );
  NAND U36592 ( .A(n35840), .B(n35839), .Z(n35961) );
  NAND U36593 ( .A(n185), .B(n35841), .Z(n35843) );
  XOR U36594 ( .A(a[248]), .B(b[9]), .Z(n36005) );
  NAND U36595 ( .A(n36805), .B(n36005), .Z(n35842) );
  NAND U36596 ( .A(n35843), .B(n35842), .Z(n35960) );
  XOR U36597 ( .A(n35957), .B(n35956), .Z(n36050) );
  NAND U36598 ( .A(n35845), .B(n35844), .Z(n35849) );
  NANDN U36599 ( .A(n35847), .B(n35846), .Z(n35848) );
  AND U36600 ( .A(n35849), .B(n35848), .Z(n36047) );
  NAND U36601 ( .A(n35851), .B(n35850), .Z(n35855) );
  NAND U36602 ( .A(n35853), .B(n35852), .Z(n35854) );
  AND U36603 ( .A(n35855), .B(n35854), .Z(n36048) );
  XOR U36604 ( .A(n36050), .B(n36049), .Z(n35948) );
  XOR U36605 ( .A(n35951), .B(n35950), .Z(n36059) );
  NAND U36606 ( .A(n35857), .B(n35856), .Z(n35861) );
  NAND U36607 ( .A(n35859), .B(n35858), .Z(n35860) );
  NAND U36608 ( .A(n35861), .B(n35860), .Z(n35945) );
  NAND U36609 ( .A(n35863), .B(n35862), .Z(n35867) );
  NANDN U36610 ( .A(n35865), .B(n35864), .Z(n35866) );
  NAND U36611 ( .A(n35867), .B(n35866), .Z(n36002) );
  NAND U36612 ( .A(n38385), .B(n35868), .Z(n35870) );
  XOR U36613 ( .A(b[27]), .B(a[230]), .Z(n35984) );
  NAND U36614 ( .A(n38343), .B(n35984), .Z(n35869) );
  NAND U36615 ( .A(n35870), .B(n35869), .Z(n36044) );
  NAND U36616 ( .A(n183), .B(n35871), .Z(n35873) );
  XOR U36617 ( .A(a[252]), .B(b[5]), .Z(n36023) );
  NAND U36618 ( .A(n36296), .B(n36023), .Z(n35872) );
  NAND U36619 ( .A(n35873), .B(n35872), .Z(n36042) );
  NAND U36620 ( .A(n190), .B(n35874), .Z(n35876) );
  XOR U36621 ( .A(b[19]), .B(a[238]), .Z(n36014) );
  NAND U36622 ( .A(n37821), .B(n36014), .Z(n35875) );
  NAND U36623 ( .A(n35876), .B(n35875), .Z(n36041) );
  NAND U36624 ( .A(n38470), .B(n35877), .Z(n35879) );
  XOR U36625 ( .A(b[31]), .B(a[226]), .Z(n36029) );
  NAND U36626 ( .A(n38453), .B(n36029), .Z(n35878) );
  NAND U36627 ( .A(n35879), .B(n35878), .Z(n35969) );
  NAND U36628 ( .A(n181), .B(n35880), .Z(n35882) );
  XOR U36629 ( .A(a[254]), .B(b[3]), .Z(n35993) );
  NAND U36630 ( .A(n182), .B(n35993), .Z(n35881) );
  NAND U36631 ( .A(n35882), .B(n35881), .Z(n35967) );
  NAND U36632 ( .A(n189), .B(n35883), .Z(n35885) );
  XOR U36633 ( .A(b[17]), .B(a[240]), .Z(n35996) );
  NAND U36634 ( .A(n37652), .B(n35996), .Z(n35884) );
  NAND U36635 ( .A(n35885), .B(n35884), .Z(n35966) );
  XOR U36636 ( .A(n36000), .B(n35999), .Z(n36001) );
  NAND U36637 ( .A(n35887), .B(n35886), .Z(n35891) );
  NAND U36638 ( .A(n35889), .B(n35888), .Z(n35890) );
  AND U36639 ( .A(n35891), .B(n35890), .Z(n36053) );
  NAND U36640 ( .A(n35893), .B(n35892), .Z(n35897) );
  NAND U36641 ( .A(n35895), .B(n35894), .Z(n35896) );
  AND U36642 ( .A(n35897), .B(n35896), .Z(n36054) );
  NAND U36643 ( .A(n35899), .B(n35898), .Z(n35903) );
  NAND U36644 ( .A(n35901), .B(n35900), .Z(n35902) );
  AND U36645 ( .A(n35903), .B(n35902), .Z(n36056) );
  XOR U36646 ( .A(n35942), .B(n35943), .Z(n35944) );
  XOR U36647 ( .A(n36062), .B(n36061), .Z(n35939) );
  NAND U36648 ( .A(n35905), .B(n35904), .Z(n35909) );
  NAND U36649 ( .A(n35907), .B(n35906), .Z(n35908) );
  AND U36650 ( .A(n35909), .B(n35908), .Z(n35936) );
  NAND U36651 ( .A(n35911), .B(n35910), .Z(n35915) );
  NAND U36652 ( .A(n35913), .B(n35912), .Z(n35914) );
  AND U36653 ( .A(n35915), .B(n35914), .Z(n35937) );
  XNOR U36654 ( .A(n35939), .B(n35938), .Z(n36066) );
  NAND U36655 ( .A(n35917), .B(n35916), .Z(n35921) );
  NAND U36656 ( .A(n35919), .B(n35918), .Z(n35920) );
  AND U36657 ( .A(n35921), .B(n35920), .Z(n36065) );
  NAND U36658 ( .A(n35923), .B(n35922), .Z(n35927) );
  NAND U36659 ( .A(n35925), .B(n35924), .Z(n35926) );
  AND U36660 ( .A(n35927), .B(n35926), .Z(n35931) );
  XOR U36661 ( .A(n35930), .B(n35931), .Z(n35932) );
  XOR U36662 ( .A(n35933), .B(n35932), .Z(n35928) );
  XOR U36663 ( .A(n35929), .B(n35928), .Z(c[480]) );
  AND U36664 ( .A(n35929), .B(n35928), .Z(n36072) );
  NAND U36665 ( .A(n35931), .B(n35930), .Z(n35935) );
  NANDN U36666 ( .A(n35933), .B(n35932), .Z(n35934) );
  AND U36667 ( .A(n35935), .B(n35934), .Z(n36076) );
  NAND U36668 ( .A(n35937), .B(n35936), .Z(n35941) );
  NAND U36669 ( .A(n35939), .B(n35938), .Z(n35940) );
  AND U36670 ( .A(n35941), .B(n35940), .Z(n36209) );
  NAND U36671 ( .A(n35943), .B(n35942), .Z(n35947) );
  NAND U36672 ( .A(n35945), .B(n35944), .Z(n35946) );
  AND U36673 ( .A(n35947), .B(n35946), .Z(n36079) );
  NAND U36674 ( .A(n35949), .B(n35948), .Z(n35953) );
  NAND U36675 ( .A(n35951), .B(n35950), .Z(n35952) );
  AND U36676 ( .A(n35953), .B(n35952), .Z(n36080) );
  NAND U36677 ( .A(n35955), .B(n35954), .Z(n35959) );
  NAND U36678 ( .A(n35957), .B(n35956), .Z(n35958) );
  NAND U36679 ( .A(n35959), .B(n35958), .Z(n36088) );
  NAND U36680 ( .A(n35961), .B(n35960), .Z(n35965) );
  NAND U36681 ( .A(n35963), .B(n35962), .Z(n35964) );
  AND U36682 ( .A(n35965), .B(n35964), .Z(n36188) );
  NAND U36683 ( .A(n35967), .B(n35966), .Z(n35971) );
  NAND U36684 ( .A(n35969), .B(n35968), .Z(n35970) );
  AND U36685 ( .A(n35971), .B(n35970), .Z(n36189) );
  NAND U36686 ( .A(n35973), .B(n35972), .Z(n35977) );
  NAND U36687 ( .A(n35975), .B(n35974), .Z(n35976) );
  AND U36688 ( .A(n35977), .B(n35976), .Z(n36191) );
  NAND U36689 ( .A(n35979), .B(n35978), .Z(n35983) );
  NAND U36690 ( .A(n35981), .B(n35980), .Z(n35982) );
  AND U36691 ( .A(n35983), .B(n35982), .Z(n36130) );
  NAND U36692 ( .A(n38385), .B(n35984), .Z(n35986) );
  XOR U36693 ( .A(b[27]), .B(a[231]), .Z(n36141) );
  NAND U36694 ( .A(n38343), .B(n36141), .Z(n35985) );
  NAND U36695 ( .A(n35986), .B(n35985), .Z(n36134) );
  NAND U36696 ( .A(n188), .B(n35987), .Z(n35989) );
  XOR U36697 ( .A(a[243]), .B(b[15]), .Z(n36168) );
  NAND U36698 ( .A(n37382), .B(n36168), .Z(n35988) );
  NAND U36699 ( .A(n35989), .B(n35988), .Z(n36133) );
  XNOR U36700 ( .A(b[1]), .B(n36133), .Z(n36135) );
  NAND U36701 ( .A(n38289), .B(n35990), .Z(n35992) );
  XOR U36702 ( .A(b[25]), .B(a[233]), .Z(n36112) );
  NAND U36703 ( .A(n38247), .B(n36112), .Z(n35991) );
  AND U36704 ( .A(n35992), .B(n35991), .Z(n36118) );
  NAND U36705 ( .A(n181), .B(n35993), .Z(n35995) );
  XOR U36706 ( .A(a[255]), .B(b[3]), .Z(n36147) );
  NAND U36707 ( .A(n182), .B(n36147), .Z(n35994) );
  NAND U36708 ( .A(n35995), .B(n35994), .Z(n36116) );
  NAND U36709 ( .A(n189), .B(n35996), .Z(n35998) );
  XOR U36710 ( .A(b[17]), .B(a[241]), .Z(n36144) );
  NAND U36711 ( .A(n37652), .B(n36144), .Z(n35997) );
  NAND U36712 ( .A(n35998), .B(n35997), .Z(n36115) );
  XOR U36713 ( .A(n36118), .B(n36117), .Z(n36127) );
  XOR U36714 ( .A(n36128), .B(n36127), .Z(n36129) );
  XOR U36715 ( .A(n36130), .B(n36129), .Z(n36085) );
  XOR U36716 ( .A(n36086), .B(n36085), .Z(n36087) );
  NAND U36717 ( .A(n36000), .B(n35999), .Z(n36004) );
  NAND U36718 ( .A(n36002), .B(n36001), .Z(n36003) );
  NAND U36719 ( .A(n36004), .B(n36003), .Z(n36195) );
  NAND U36720 ( .A(n185), .B(n36005), .Z(n36007) );
  XOR U36721 ( .A(a[249]), .B(b[9]), .Z(n36097) );
  NAND U36722 ( .A(n36805), .B(n36097), .Z(n36006) );
  NAND U36723 ( .A(n36007), .B(n36006), .Z(n36124) );
  NAND U36724 ( .A(n186), .B(n36008), .Z(n36010) );
  XOR U36725 ( .A(a[247]), .B(b[11]), .Z(n36109) );
  NAND U36726 ( .A(n37097), .B(n36109), .Z(n36009) );
  NAND U36727 ( .A(n36010), .B(n36009), .Z(n36122) );
  NAND U36728 ( .A(n187), .B(n36011), .Z(n36013) );
  XOR U36729 ( .A(a[245]), .B(b[13]), .Z(n36106) );
  NAND U36730 ( .A(n37295), .B(n36106), .Z(n36012) );
  NAND U36731 ( .A(n36013), .B(n36012), .Z(n36094) );
  NAND U36732 ( .A(n190), .B(n36014), .Z(n36016) );
  XOR U36733 ( .A(b[19]), .B(a[239]), .Z(n36153) );
  NAND U36734 ( .A(n37821), .B(n36153), .Z(n36015) );
  NAND U36735 ( .A(n36016), .B(n36015), .Z(n36092) );
  NAND U36736 ( .A(n184), .B(n36017), .Z(n36019) );
  XOR U36737 ( .A(a[251]), .B(b[7]), .Z(n36100) );
  NAND U36738 ( .A(n36592), .B(n36100), .Z(n36018) );
  NAND U36739 ( .A(n36019), .B(n36018), .Z(n36091) );
  XNOR U36740 ( .A(n36124), .B(n36123), .Z(n36158) );
  NAND U36741 ( .A(n38064), .B(n36020), .Z(n36022) );
  XOR U36742 ( .A(b[21]), .B(a[237]), .Z(n36103) );
  NAND U36743 ( .A(n37993), .B(n36103), .Z(n36021) );
  NAND U36744 ( .A(n36022), .B(n36021), .Z(n36185) );
  NAND U36745 ( .A(n183), .B(n36023), .Z(n36025) );
  XOR U36746 ( .A(a[253]), .B(b[5]), .Z(n36150) );
  NAND U36747 ( .A(n36296), .B(n36150), .Z(n36024) );
  NAND U36748 ( .A(n36025), .B(n36024), .Z(n36183) );
  NAND U36749 ( .A(n38185), .B(n36026), .Z(n36028) );
  XOR U36750 ( .A(b[23]), .B(a[235]), .Z(n36138) );
  NAND U36751 ( .A(n38132), .B(n36138), .Z(n36027) );
  NAND U36752 ( .A(n36028), .B(n36027), .Z(n36182) );
  NAND U36753 ( .A(n38470), .B(n36029), .Z(n36031) );
  XOR U36754 ( .A(b[31]), .B(a[227]), .Z(n36174) );
  NAND U36755 ( .A(n38453), .B(n36174), .Z(n36030) );
  NAND U36756 ( .A(n36031), .B(n36030), .Z(n36179) );
  AND U36757 ( .A(b[31]), .B(a[225]), .Z(n36410) );
  NAND U36758 ( .A(n194), .B(n36032), .Z(n36034) );
  XOR U36759 ( .A(b[29]), .B(a[229]), .Z(n36171) );
  NAND U36760 ( .A(n38456), .B(n36171), .Z(n36033) );
  NAND U36761 ( .A(n36034), .B(n36033), .Z(n36177) );
  XNOR U36762 ( .A(n36410), .B(n36177), .Z(n36178) );
  XNOR U36763 ( .A(n36179), .B(n36178), .Z(n36156) );
  XOR U36764 ( .A(n36158), .B(n36159), .Z(n36164) );
  NAND U36765 ( .A(n36036), .B(n36035), .Z(n36040) );
  NANDN U36766 ( .A(n36038), .B(n36037), .Z(n36039) );
  NAND U36767 ( .A(n36040), .B(n36039), .Z(n36163) );
  NAND U36768 ( .A(n36042), .B(n36041), .Z(n36046) );
  NAND U36769 ( .A(n36044), .B(n36043), .Z(n36045) );
  NAND U36770 ( .A(n36046), .B(n36045), .Z(n36162) );
  XOR U36771 ( .A(n36164), .B(n36165), .Z(n36194) );
  NAND U36772 ( .A(n36048), .B(n36047), .Z(n36052) );
  NAND U36773 ( .A(n36050), .B(n36049), .Z(n36051) );
  AND U36774 ( .A(n36052), .B(n36051), .Z(n36197) );
  NAND U36775 ( .A(n36054), .B(n36053), .Z(n36058) );
  NAND U36776 ( .A(n36056), .B(n36055), .Z(n36057) );
  AND U36777 ( .A(n36058), .B(n36057), .Z(n36201) );
  XOR U36778 ( .A(n36202), .B(n36203), .Z(n36081) );
  XOR U36779 ( .A(n36082), .B(n36081), .Z(n36206) );
  NAND U36780 ( .A(n36060), .B(n36059), .Z(n36064) );
  NAND U36781 ( .A(n36062), .B(n36061), .Z(n36063) );
  AND U36782 ( .A(n36064), .B(n36063), .Z(n36207) );
  XNOR U36783 ( .A(n36209), .B(n36208), .Z(n36074) );
  NAND U36784 ( .A(n36066), .B(n36065), .Z(n36070) );
  NAND U36785 ( .A(n36068), .B(n36067), .Z(n36069) );
  AND U36786 ( .A(n36070), .B(n36069), .Z(n36073) );
  XOR U36787 ( .A(n36076), .B(n36075), .Z(n36071) );
  XOR U36788 ( .A(n36072), .B(n36071), .Z(c[481]) );
  AND U36789 ( .A(n36072), .B(n36071), .Z(n36213) );
  NAND U36790 ( .A(n36074), .B(n36073), .Z(n36078) );
  NANDN U36791 ( .A(n36076), .B(n36075), .Z(n36077) );
  AND U36792 ( .A(n36078), .B(n36077), .Z(n36217) );
  NAND U36793 ( .A(n36080), .B(n36079), .Z(n36084) );
  NAND U36794 ( .A(n36082), .B(n36081), .Z(n36083) );
  AND U36795 ( .A(n36084), .B(n36083), .Z(n36223) );
  NAND U36796 ( .A(n36086), .B(n36085), .Z(n36090) );
  NAND U36797 ( .A(n36088), .B(n36087), .Z(n36089) );
  AND U36798 ( .A(n36090), .B(n36089), .Z(n36351) );
  NAND U36799 ( .A(n36092), .B(n36091), .Z(n36096) );
  NAND U36800 ( .A(n36094), .B(n36093), .Z(n36095) );
  AND U36801 ( .A(n36096), .B(n36095), .Z(n36280) );
  NAND U36802 ( .A(n185), .B(n36097), .Z(n36099) );
  XOR U36803 ( .A(a[250]), .B(b[9]), .Z(n36309) );
  NAND U36804 ( .A(n36805), .B(n36309), .Z(n36098) );
  NAND U36805 ( .A(n36099), .B(n36098), .Z(n36268) );
  NAND U36806 ( .A(n184), .B(n36100), .Z(n36102) );
  XOR U36807 ( .A(a[252]), .B(b[7]), .Z(n36321) );
  NAND U36808 ( .A(n36592), .B(n36321), .Z(n36101) );
  NAND U36809 ( .A(n36102), .B(n36101), .Z(n36266) );
  NAND U36810 ( .A(n38064), .B(n36103), .Z(n36105) );
  XOR U36811 ( .A(b[21]), .B(a[238]), .Z(n36327) );
  NAND U36812 ( .A(n37993), .B(n36327), .Z(n36104) );
  NAND U36813 ( .A(n36105), .B(n36104), .Z(n36265) );
  NAND U36814 ( .A(n187), .B(n36106), .Z(n36108) );
  XOR U36815 ( .A(a[246]), .B(b[13]), .Z(n36250) );
  NAND U36816 ( .A(n37295), .B(n36250), .Z(n36107) );
  AND U36817 ( .A(n36108), .B(n36107), .Z(n36292) );
  NAND U36818 ( .A(n186), .B(n36109), .Z(n36111) );
  XOR U36819 ( .A(a[248]), .B(b[11]), .Z(n36318) );
  NAND U36820 ( .A(n37097), .B(n36318), .Z(n36110) );
  NAND U36821 ( .A(n36111), .B(n36110), .Z(n36290) );
  NAND U36822 ( .A(n38289), .B(n36112), .Z(n36114) );
  XOR U36823 ( .A(b[25]), .B(a[234]), .Z(n36312) );
  NAND U36824 ( .A(n38247), .B(n36312), .Z(n36113) );
  NAND U36825 ( .A(n36114), .B(n36113), .Z(n36289) );
  XOR U36826 ( .A(n36292), .B(n36291), .Z(n36277) );
  XOR U36827 ( .A(n36278), .B(n36277), .Z(n36279) );
  XOR U36828 ( .A(n36280), .B(n36279), .Z(n36336) );
  NAND U36829 ( .A(n36116), .B(n36115), .Z(n36120) );
  NANDN U36830 ( .A(n36118), .B(n36117), .Z(n36119) );
  AND U36831 ( .A(n36120), .B(n36119), .Z(n36337) );
  NAND U36832 ( .A(n36122), .B(n36121), .Z(n36126) );
  NAND U36833 ( .A(n36124), .B(n36123), .Z(n36125) );
  AND U36834 ( .A(n36126), .B(n36125), .Z(n36338) );
  XNOR U36835 ( .A(n36339), .B(n36338), .Z(n36349) );
  NAND U36836 ( .A(n36128), .B(n36127), .Z(n36132) );
  NAND U36837 ( .A(n36130), .B(n36129), .Z(n36131) );
  AND U36838 ( .A(n36132), .B(n36131), .Z(n36235) );
  NANDN U36839 ( .A(b[1]), .B(n36133), .Z(n36137) );
  NAND U36840 ( .A(n36135), .B(n36134), .Z(n36136) );
  AND U36841 ( .A(n36137), .B(n36136), .Z(n36286) );
  NAND U36842 ( .A(n38185), .B(n36138), .Z(n36140) );
  XOR U36843 ( .A(b[23]), .B(a[236]), .Z(n36303) );
  NAND U36844 ( .A(n38132), .B(n36303), .Z(n36139) );
  NAND U36845 ( .A(n36140), .B(n36139), .Z(n36262) );
  NAND U36846 ( .A(n38385), .B(n36141), .Z(n36143) );
  XOR U36847 ( .A(b[27]), .B(a[232]), .Z(n36315) );
  NAND U36848 ( .A(n38343), .B(n36315), .Z(n36142) );
  NAND U36849 ( .A(n36143), .B(n36142), .Z(n36260) );
  NAND U36850 ( .A(n189), .B(n36144), .Z(n36146) );
  XOR U36851 ( .A(b[17]), .B(a[242]), .Z(n36247) );
  NAND U36852 ( .A(n37652), .B(n36247), .Z(n36145) );
  NAND U36853 ( .A(n36146), .B(n36145), .Z(n36259) );
  NAND U36854 ( .A(n182), .B(b[3]), .Z(n36149) );
  NANDN U36855 ( .A(n180), .B(n36147), .Z(n36148) );
  AND U36856 ( .A(n36149), .B(n36148), .Z(n36254) );
  NAND U36857 ( .A(b[31]), .B(a[226]), .Z(n36253) );
  XNOR U36858 ( .A(n36410), .B(n36255), .Z(n36274) );
  NAND U36859 ( .A(n183), .B(n36150), .Z(n36152) );
  XOR U36860 ( .A(a[254]), .B(b[5]), .Z(n36295) );
  NAND U36861 ( .A(n36296), .B(n36295), .Z(n36151) );
  NAND U36862 ( .A(n36152), .B(n36151), .Z(n36272) );
  NAND U36863 ( .A(n190), .B(n36153), .Z(n36155) );
  XOR U36864 ( .A(b[19]), .B(a[240]), .Z(n36299) );
  NAND U36865 ( .A(n37821), .B(n36299), .Z(n36154) );
  NAND U36866 ( .A(n36155), .B(n36154), .Z(n36271) );
  XNOR U36867 ( .A(n36274), .B(n36273), .Z(n36283) );
  XOR U36868 ( .A(n36284), .B(n36283), .Z(n36285) );
  XNOR U36869 ( .A(n36286), .B(n36285), .Z(n36233) );
  NAND U36870 ( .A(n36157), .B(n36156), .Z(n36161) );
  NANDN U36871 ( .A(n36159), .B(n36158), .Z(n36160) );
  AND U36872 ( .A(n36161), .B(n36160), .Z(n36232) );
  XOR U36873 ( .A(n36235), .B(n36234), .Z(n36348) );
  XNOR U36874 ( .A(n36351), .B(n36350), .Z(n36345) );
  NAND U36875 ( .A(n36163), .B(n36162), .Z(n36167) );
  NAND U36876 ( .A(n36165), .B(n36164), .Z(n36166) );
  NAND U36877 ( .A(n36167), .B(n36166), .Z(n36229) );
  NAND U36878 ( .A(n188), .B(n36168), .Z(n36170) );
  XOR U36879 ( .A(a[244]), .B(b[15]), .Z(n36244) );
  NAND U36880 ( .A(n37382), .B(n36244), .Z(n36169) );
  NAND U36881 ( .A(n36170), .B(n36169), .Z(n36333) );
  NAND U36882 ( .A(n194), .B(n36171), .Z(n36173) );
  XOR U36883 ( .A(b[29]), .B(a[230]), .Z(n36306) );
  NAND U36884 ( .A(n38456), .B(n36306), .Z(n36172) );
  NAND U36885 ( .A(n36173), .B(n36172), .Z(n36331) );
  NAND U36886 ( .A(n38470), .B(n36174), .Z(n36176) );
  XOR U36887 ( .A(b[31]), .B(a[228]), .Z(n36324) );
  NAND U36888 ( .A(n38453), .B(n36324), .Z(n36175) );
  NAND U36889 ( .A(n36176), .B(n36175), .Z(n36330) );
  IV U36890 ( .A(n36410), .Z(n36256) );
  NAND U36891 ( .A(n36256), .B(n36177), .Z(n36181) );
  NAND U36892 ( .A(n36179), .B(n36178), .Z(n36180) );
  AND U36893 ( .A(n36181), .B(n36180), .Z(n36239) );
  XOR U36894 ( .A(n36238), .B(n36239), .Z(n36241) );
  NAND U36895 ( .A(n36183), .B(n36182), .Z(n36187) );
  NAND U36896 ( .A(n36185), .B(n36184), .Z(n36186) );
  AND U36897 ( .A(n36187), .B(n36186), .Z(n36240) );
  XNOR U36898 ( .A(n36241), .B(n36240), .Z(n36227) );
  NAND U36899 ( .A(n36189), .B(n36188), .Z(n36193) );
  NAND U36900 ( .A(n36191), .B(n36190), .Z(n36192) );
  AND U36901 ( .A(n36193), .B(n36192), .Z(n36226) );
  NAND U36902 ( .A(n36195), .B(n36194), .Z(n36199) );
  NAND U36903 ( .A(n36197), .B(n36196), .Z(n36198) );
  AND U36904 ( .A(n36199), .B(n36198), .Z(n36343) );
  XOR U36905 ( .A(n36342), .B(n36343), .Z(n36344) );
  NAND U36906 ( .A(n36201), .B(n36200), .Z(n36205) );
  NAND U36907 ( .A(n36203), .B(n36202), .Z(n36204) );
  AND U36908 ( .A(n36205), .B(n36204), .Z(n36221) );
  XOR U36909 ( .A(n36223), .B(n36222), .Z(n36214) );
  NAND U36910 ( .A(n36207), .B(n36206), .Z(n36211) );
  NAND U36911 ( .A(n36209), .B(n36208), .Z(n36210) );
  AND U36912 ( .A(n36211), .B(n36210), .Z(n36215) );
  XOR U36913 ( .A(n36217), .B(n36216), .Z(n36212) );
  XOR U36914 ( .A(n36213), .B(n36212), .Z(c[482]) );
  AND U36915 ( .A(n36213), .B(n36212), .Z(n36355) );
  NAND U36916 ( .A(n36215), .B(n36214), .Z(n36219) );
  NANDN U36917 ( .A(n36217), .B(n36216), .Z(n36218) );
  AND U36918 ( .A(n36219), .B(n36218), .Z(n36359) );
  NAND U36919 ( .A(n36221), .B(n36220), .Z(n36225) );
  NAND U36920 ( .A(n36223), .B(n36222), .Z(n36224) );
  NAND U36921 ( .A(n36225), .B(n36224), .Z(n36357) );
  NAND U36922 ( .A(n36227), .B(n36226), .Z(n36231) );
  NAND U36923 ( .A(n36229), .B(n36228), .Z(n36230) );
  NAND U36924 ( .A(n36231), .B(n36230), .Z(n36369) );
  NAND U36925 ( .A(n36233), .B(n36232), .Z(n36237) );
  NAND U36926 ( .A(n36235), .B(n36234), .Z(n36236) );
  NAND U36927 ( .A(n36237), .B(n36236), .Z(n36368) );
  NAND U36928 ( .A(n36239), .B(n36238), .Z(n36243) );
  NAND U36929 ( .A(n36241), .B(n36240), .Z(n36242) );
  NAND U36930 ( .A(n36243), .B(n36242), .Z(n36474) );
  NAND U36931 ( .A(n188), .B(n36244), .Z(n36246) );
  XOR U36932 ( .A(a[245]), .B(b[15]), .Z(n36398) );
  NAND U36933 ( .A(n37382), .B(n36398), .Z(n36245) );
  NAND U36934 ( .A(n36246), .B(n36245), .Z(n36416) );
  NAND U36935 ( .A(n189), .B(n36247), .Z(n36249) );
  XOR U36936 ( .A(b[17]), .B(a[243]), .Z(n36401) );
  NAND U36937 ( .A(n37652), .B(n36401), .Z(n36248) );
  NAND U36938 ( .A(n36249), .B(n36248), .Z(n36414) );
  NAND U36939 ( .A(n187), .B(n36250), .Z(n36252) );
  XOR U36940 ( .A(a[247]), .B(b[13]), .Z(n36404) );
  NAND U36941 ( .A(n37295), .B(n36404), .Z(n36251) );
  NAND U36942 ( .A(n36252), .B(n36251), .Z(n36413) );
  OR U36943 ( .A(n36254), .B(n36253), .Z(n36258) );
  NAND U36944 ( .A(n36256), .B(n36255), .Z(n36257) );
  AND U36945 ( .A(n36258), .B(n36257), .Z(n36420) );
  XOR U36946 ( .A(n36419), .B(n36420), .Z(n36422) );
  NAND U36947 ( .A(n36260), .B(n36259), .Z(n36264) );
  NAND U36948 ( .A(n36262), .B(n36261), .Z(n36263) );
  AND U36949 ( .A(n36264), .B(n36263), .Z(n36421) );
  XNOR U36950 ( .A(n36422), .B(n36421), .Z(n36480) );
  NAND U36951 ( .A(n36266), .B(n36265), .Z(n36270) );
  NAND U36952 ( .A(n36268), .B(n36267), .Z(n36269) );
  NAND U36953 ( .A(n36270), .B(n36269), .Z(n36478) );
  NAND U36954 ( .A(n36272), .B(n36271), .Z(n36276) );
  NAND U36955 ( .A(n36274), .B(n36273), .Z(n36275) );
  NAND U36956 ( .A(n36276), .B(n36275), .Z(n36477) );
  NAND U36957 ( .A(n36278), .B(n36277), .Z(n36282) );
  NAND U36958 ( .A(n36280), .B(n36279), .Z(n36281) );
  NAND U36959 ( .A(n36282), .B(n36281), .Z(n36471) );
  XOR U36960 ( .A(n36472), .B(n36471), .Z(n36473) );
  NAND U36961 ( .A(n36284), .B(n36283), .Z(n36288) );
  NAND U36962 ( .A(n36286), .B(n36285), .Z(n36287) );
  NAND U36963 ( .A(n36288), .B(n36287), .Z(n36383) );
  NAND U36964 ( .A(n36290), .B(n36289), .Z(n36294) );
  NANDN U36965 ( .A(n36292), .B(n36291), .Z(n36293) );
  NAND U36966 ( .A(n36294), .B(n36293), .Z(n36492) );
  NAND U36967 ( .A(n183), .B(n36295), .Z(n36298) );
  XOR U36968 ( .A(a[255]), .B(b[5]), .Z(n36461) );
  NAND U36969 ( .A(n36296), .B(n36461), .Z(n36297) );
  NAND U36970 ( .A(n36298), .B(n36297), .Z(n36393) );
  NAND U36971 ( .A(n190), .B(n36299), .Z(n36301) );
  XOR U36972 ( .A(b[19]), .B(a[241]), .Z(n36440) );
  NAND U36973 ( .A(n37821), .B(n36440), .Z(n36300) );
  NAND U36974 ( .A(n36301), .B(n36300), .Z(n36392) );
  AND U36975 ( .A(b[31]), .B(a[227]), .Z(n36407) );
  XNOR U36976 ( .A(n36407), .B(n36302), .Z(n36409) );
  XOR U36977 ( .A(n36410), .B(n36409), .Z(n36394) );
  XOR U36978 ( .A(n36395), .B(n36394), .Z(n36490) );
  NAND U36979 ( .A(n38185), .B(n36303), .Z(n36305) );
  XOR U36980 ( .A(b[23]), .B(a[237]), .Z(n36425) );
  NAND U36981 ( .A(n38132), .B(n36425), .Z(n36304) );
  NAND U36982 ( .A(n36305), .B(n36304), .Z(n36468) );
  NAND U36983 ( .A(n194), .B(n36306), .Z(n36308) );
  XOR U36984 ( .A(b[29]), .B(a[231]), .Z(n36437) );
  NAND U36985 ( .A(n38456), .B(n36437), .Z(n36307) );
  NAND U36986 ( .A(n36308), .B(n36307), .Z(n36466) );
  NAND U36987 ( .A(n185), .B(n36309), .Z(n36311) );
  XOR U36988 ( .A(a[251]), .B(b[9]), .Z(n36452) );
  NAND U36989 ( .A(n36805), .B(n36452), .Z(n36310) );
  NAND U36990 ( .A(n36311), .B(n36310), .Z(n36465) );
  XOR U36991 ( .A(n36490), .B(n36489), .Z(n36491) );
  NAND U36992 ( .A(n38289), .B(n36312), .Z(n36314) );
  XOR U36993 ( .A(b[25]), .B(a[235]), .Z(n36428) );
  NAND U36994 ( .A(n38247), .B(n36428), .Z(n36313) );
  NAND U36995 ( .A(n36314), .B(n36313), .Z(n36446) );
  NAND U36996 ( .A(n38385), .B(n36315), .Z(n36317) );
  XOR U36997 ( .A(b[27]), .B(a[233]), .Z(n36449) );
  NAND U36998 ( .A(n38343), .B(n36449), .Z(n36316) );
  NAND U36999 ( .A(n36317), .B(n36316), .Z(n36444) );
  NAND U37000 ( .A(n186), .B(n36318), .Z(n36320) );
  XOR U37001 ( .A(a[249]), .B(b[11]), .Z(n36431) );
  NAND U37002 ( .A(n37097), .B(n36431), .Z(n36319) );
  NAND U37003 ( .A(n36320), .B(n36319), .Z(n36443) );
  NAND U37004 ( .A(n184), .B(n36321), .Z(n36323) );
  XOR U37005 ( .A(a[253]), .B(b[7]), .Z(n36434) );
  NAND U37006 ( .A(n36592), .B(n36434), .Z(n36322) );
  AND U37007 ( .A(n36323), .B(n36322), .Z(n36389) );
  NAND U37008 ( .A(n38470), .B(n36324), .Z(n36326) );
  XOR U37009 ( .A(b[31]), .B(a[229]), .Z(n36458) );
  NAND U37010 ( .A(n38453), .B(n36458), .Z(n36325) );
  NAND U37011 ( .A(n36326), .B(n36325), .Z(n36387) );
  NAND U37012 ( .A(n38064), .B(n36327), .Z(n36329) );
  XOR U37013 ( .A(b[21]), .B(a[239]), .Z(n36455) );
  NAND U37014 ( .A(n37993), .B(n36455), .Z(n36328) );
  NAND U37015 ( .A(n36329), .B(n36328), .Z(n36386) );
  XOR U37016 ( .A(n36389), .B(n36388), .Z(n36483) );
  XOR U37017 ( .A(n36484), .B(n36483), .Z(n36485) );
  NAND U37018 ( .A(n36331), .B(n36330), .Z(n36335) );
  NAND U37019 ( .A(n36333), .B(n36332), .Z(n36334) );
  AND U37020 ( .A(n36335), .B(n36334), .Z(n36486) );
  XOR U37021 ( .A(n36380), .B(n36381), .Z(n36382) );
  NAND U37022 ( .A(n36337), .B(n36336), .Z(n36341) );
  NAND U37023 ( .A(n36339), .B(n36338), .Z(n36340) );
  AND U37024 ( .A(n36341), .B(n36340), .Z(n36375) );
  XOR U37025 ( .A(n36374), .B(n36375), .Z(n36377) );
  XOR U37026 ( .A(n36376), .B(n36377), .Z(n36370) );
  XNOR U37027 ( .A(n36371), .B(n36370), .Z(n36365) );
  NAND U37028 ( .A(n36343), .B(n36342), .Z(n36347) );
  NAND U37029 ( .A(n36345), .B(n36344), .Z(n36346) );
  NAND U37030 ( .A(n36347), .B(n36346), .Z(n36363) );
  NAND U37031 ( .A(n36349), .B(n36348), .Z(n36353) );
  NAND U37032 ( .A(n36351), .B(n36350), .Z(n36352) );
  AND U37033 ( .A(n36353), .B(n36352), .Z(n36362) );
  XOR U37034 ( .A(n36359), .B(n36358), .Z(n36354) );
  XOR U37035 ( .A(n36355), .B(n36354), .Z(c[483]) );
  AND U37036 ( .A(n36355), .B(n36354), .Z(n36496) );
  NAND U37037 ( .A(n36357), .B(n36356), .Z(n36361) );
  NANDN U37038 ( .A(n36359), .B(n36358), .Z(n36360) );
  AND U37039 ( .A(n36361), .B(n36360), .Z(n36500) );
  NAND U37040 ( .A(n36363), .B(n36362), .Z(n36367) );
  NAND U37041 ( .A(n36365), .B(n36364), .Z(n36366) );
  NAND U37042 ( .A(n36367), .B(n36366), .Z(n36498) );
  NAND U37043 ( .A(n36369), .B(n36368), .Z(n36373) );
  NAND U37044 ( .A(n36371), .B(n36370), .Z(n36372) );
  AND U37045 ( .A(n36373), .B(n36372), .Z(n36506) );
  NAND U37046 ( .A(n36375), .B(n36374), .Z(n36379) );
  NAND U37047 ( .A(n36377), .B(n36376), .Z(n36378) );
  AND U37048 ( .A(n36379), .B(n36378), .Z(n36504) );
  NAND U37049 ( .A(n36381), .B(n36380), .Z(n36385) );
  NAND U37050 ( .A(n36383), .B(n36382), .Z(n36384) );
  NAND U37051 ( .A(n36385), .B(n36384), .Z(n36512) );
  NAND U37052 ( .A(n36387), .B(n36386), .Z(n36391) );
  NANDN U37053 ( .A(n36389), .B(n36388), .Z(n36390) );
  NAND U37054 ( .A(n36391), .B(n36390), .Z(n36516) );
  NAND U37055 ( .A(n36393), .B(n36392), .Z(n36397) );
  NAND U37056 ( .A(n36395), .B(n36394), .Z(n36396) );
  NAND U37057 ( .A(n36397), .B(n36396), .Z(n36515) );
  NAND U37058 ( .A(n188), .B(n36398), .Z(n36400) );
  XOR U37059 ( .A(a[246]), .B(b[15]), .Z(n36598) );
  NAND U37060 ( .A(n37382), .B(n36598), .Z(n36399) );
  NAND U37061 ( .A(n36400), .B(n36399), .Z(n36554) );
  NAND U37062 ( .A(n189), .B(n36401), .Z(n36403) );
  XOR U37063 ( .A(a[244]), .B(b[17]), .Z(n36604) );
  NAND U37064 ( .A(n37652), .B(n36604), .Z(n36402) );
  NAND U37065 ( .A(n36403), .B(n36402), .Z(n36552) );
  NAND U37066 ( .A(n187), .B(n36404), .Z(n36406) );
  XOR U37067 ( .A(a[248]), .B(b[13]), .Z(n36601) );
  NAND U37068 ( .A(n37295), .B(n36601), .Z(n36405) );
  NAND U37069 ( .A(n36406), .B(n36405), .Z(n36551) );
  NAND U37070 ( .A(n36408), .B(n36407), .Z(n36412) );
  NAND U37071 ( .A(n36410), .B(n36409), .Z(n36411) );
  NAND U37072 ( .A(n36412), .B(n36411), .Z(n36545) );
  XOR U37073 ( .A(n36546), .B(n36545), .Z(n36548) );
  NAND U37074 ( .A(n36414), .B(n36413), .Z(n36418) );
  NAND U37075 ( .A(n36416), .B(n36415), .Z(n36417) );
  NAND U37076 ( .A(n36418), .B(n36417), .Z(n36547) );
  XOR U37077 ( .A(n36548), .B(n36547), .Z(n36517) );
  XNOR U37078 ( .A(n36518), .B(n36517), .Z(n36510) );
  NAND U37079 ( .A(n36420), .B(n36419), .Z(n36424) );
  NAND U37080 ( .A(n36422), .B(n36421), .Z(n36423) );
  NAND U37081 ( .A(n36424), .B(n36423), .Z(n36542) );
  NAND U37082 ( .A(n38185), .B(n36425), .Z(n36427) );
  XOR U37083 ( .A(b[23]), .B(a[238]), .Z(n36573) );
  NAND U37084 ( .A(n38132), .B(n36573), .Z(n36426) );
  NAND U37085 ( .A(n36427), .B(n36426), .Z(n36616) );
  NAND U37086 ( .A(n38289), .B(n36428), .Z(n36430) );
  XOR U37087 ( .A(b[25]), .B(a[236]), .Z(n36607) );
  NAND U37088 ( .A(n38247), .B(n36607), .Z(n36429) );
  NAND U37089 ( .A(n36430), .B(n36429), .Z(n36614) );
  NAND U37090 ( .A(n186), .B(n36431), .Z(n36433) );
  XOR U37091 ( .A(a[250]), .B(b[11]), .Z(n36610) );
  NAND U37092 ( .A(n37097), .B(n36610), .Z(n36432) );
  NAND U37093 ( .A(n36433), .B(n36432), .Z(n36613) );
  NAND U37094 ( .A(n184), .B(n36434), .Z(n36436) );
  XOR U37095 ( .A(a[254]), .B(b[7]), .Z(n36591) );
  NAND U37096 ( .A(n36592), .B(n36591), .Z(n36435) );
  AND U37097 ( .A(n36436), .B(n36435), .Z(n36585) );
  NAND U37098 ( .A(n194), .B(n36437), .Z(n36439) );
  XOR U37099 ( .A(b[29]), .B(a[232]), .Z(n36588) );
  NAND U37100 ( .A(n38456), .B(n36588), .Z(n36438) );
  NAND U37101 ( .A(n36439), .B(n36438), .Z(n36583) );
  NAND U37102 ( .A(n190), .B(n36440), .Z(n36442) );
  XOR U37103 ( .A(b[19]), .B(a[242]), .Z(n36569) );
  NAND U37104 ( .A(n37821), .B(n36569), .Z(n36441) );
  NAND U37105 ( .A(n36442), .B(n36441), .Z(n36582) );
  XOR U37106 ( .A(n36585), .B(n36584), .Z(n36521) );
  XOR U37107 ( .A(n36522), .B(n36521), .Z(n36523) );
  NAND U37108 ( .A(n36444), .B(n36443), .Z(n36448) );
  NAND U37109 ( .A(n36446), .B(n36445), .Z(n36447) );
  AND U37110 ( .A(n36448), .B(n36447), .Z(n36524) );
  NAND U37111 ( .A(n38385), .B(n36449), .Z(n36451) );
  XOR U37112 ( .A(b[27]), .B(a[234]), .Z(n36579) );
  NAND U37113 ( .A(n38343), .B(n36579), .Z(n36450) );
  NAND U37114 ( .A(n36451), .B(n36450), .Z(n36560) );
  NAND U37115 ( .A(n185), .B(n36452), .Z(n36454) );
  XOR U37116 ( .A(a[252]), .B(b[9]), .Z(n36576) );
  NAND U37117 ( .A(n36805), .B(n36576), .Z(n36453) );
  NAND U37118 ( .A(n36454), .B(n36453), .Z(n36558) );
  NAND U37119 ( .A(n38064), .B(n36455), .Z(n36457) );
  XOR U37120 ( .A(b[21]), .B(a[240]), .Z(n36595) );
  NAND U37121 ( .A(n37993), .B(n36595), .Z(n36456) );
  NAND U37122 ( .A(n36457), .B(n36456), .Z(n36557) );
  NAND U37123 ( .A(n38470), .B(n36458), .Z(n36460) );
  XOR U37124 ( .A(b[31]), .B(a[230]), .Z(n36566) );
  NAND U37125 ( .A(n38453), .B(n36566), .Z(n36459) );
  AND U37126 ( .A(n36460), .B(n36459), .Z(n36565) );
  AND U37127 ( .A(b[31]), .B(a[228]), .Z(n36724) );
  AND U37128 ( .A(n36461), .B(n183), .Z(n36464) );
  XOR U37129 ( .A(b[4]), .B(b[3]), .Z(n36462) );
  NAND U37130 ( .A(b[5]), .B(n36462), .Z(n36463) );
  NANDN U37131 ( .A(n36464), .B(n36463), .Z(n36563) );
  XNOR U37132 ( .A(n36724), .B(n36563), .Z(n36564) );
  XOR U37133 ( .A(n36565), .B(n36564), .Z(n36527) );
  XOR U37134 ( .A(n36528), .B(n36527), .Z(n36529) );
  NAND U37135 ( .A(n36466), .B(n36465), .Z(n36470) );
  NAND U37136 ( .A(n36468), .B(n36467), .Z(n36469) );
  AND U37137 ( .A(n36470), .B(n36469), .Z(n36530) );
  XOR U37138 ( .A(n36540), .B(n36539), .Z(n36541) );
  NAND U37139 ( .A(n36472), .B(n36471), .Z(n36476) );
  NAND U37140 ( .A(n36474), .B(n36473), .Z(n36475) );
  NAND U37141 ( .A(n36476), .B(n36475), .Z(n36620) );
  NAND U37142 ( .A(n36478), .B(n36477), .Z(n36482) );
  NAND U37143 ( .A(n36480), .B(n36479), .Z(n36481) );
  AND U37144 ( .A(n36482), .B(n36481), .Z(n36536) );
  NAND U37145 ( .A(n36484), .B(n36483), .Z(n36488) );
  NAND U37146 ( .A(n36486), .B(n36485), .Z(n36487) );
  NAND U37147 ( .A(n36488), .B(n36487), .Z(n36534) );
  NAND U37148 ( .A(n36490), .B(n36489), .Z(n36494) );
  NAND U37149 ( .A(n36492), .B(n36491), .Z(n36493) );
  AND U37150 ( .A(n36494), .B(n36493), .Z(n36533) );
  XOR U37151 ( .A(n36536), .B(n36535), .Z(n36619) );
  XOR U37152 ( .A(n36622), .B(n36621), .Z(n36503) );
  XOR U37153 ( .A(n36504), .B(n36503), .Z(n36505) );
  XOR U37154 ( .A(n36506), .B(n36505), .Z(n36497) );
  XOR U37155 ( .A(n36500), .B(n36499), .Z(n36495) );
  XOR U37156 ( .A(n36496), .B(n36495), .Z(c[484]) );
  AND U37157 ( .A(n36496), .B(n36495), .Z(n36626) );
  NAND U37158 ( .A(n36498), .B(n36497), .Z(n36502) );
  NANDN U37159 ( .A(n36500), .B(n36499), .Z(n36501) );
  AND U37160 ( .A(n36502), .B(n36501), .Z(n36630) );
  NAND U37161 ( .A(n36504), .B(n36503), .Z(n36508) );
  NAND U37162 ( .A(n36506), .B(n36505), .Z(n36507) );
  NAND U37163 ( .A(n36508), .B(n36507), .Z(n36628) );
  NAND U37164 ( .A(n36510), .B(n36509), .Z(n36514) );
  NAND U37165 ( .A(n36512), .B(n36511), .Z(n36513) );
  AND U37166 ( .A(n36514), .B(n36513), .Z(n36636) );
  NAND U37167 ( .A(n36516), .B(n36515), .Z(n36520) );
  NAND U37168 ( .A(n36518), .B(n36517), .Z(n36519) );
  AND U37169 ( .A(n36520), .B(n36519), .Z(n36642) );
  NAND U37170 ( .A(n36522), .B(n36521), .Z(n36526) );
  NAND U37171 ( .A(n36524), .B(n36523), .Z(n36525) );
  NAND U37172 ( .A(n36526), .B(n36525), .Z(n36640) );
  NAND U37173 ( .A(n36528), .B(n36527), .Z(n36532) );
  NAND U37174 ( .A(n36530), .B(n36529), .Z(n36531) );
  NAND U37175 ( .A(n36532), .B(n36531), .Z(n36639) );
  XNOR U37176 ( .A(n36642), .B(n36641), .Z(n36634) );
  NAND U37177 ( .A(n36534), .B(n36533), .Z(n36538) );
  NAND U37178 ( .A(n36536), .B(n36535), .Z(n36537) );
  AND U37179 ( .A(n36538), .B(n36537), .Z(n36633) );
  XOR U37180 ( .A(n36636), .B(n36635), .Z(n36752) );
  NAND U37181 ( .A(n36540), .B(n36539), .Z(n36544) );
  NAND U37182 ( .A(n36542), .B(n36541), .Z(n36543) );
  AND U37183 ( .A(n36544), .B(n36543), .Z(n36748) );
  NAND U37184 ( .A(n36546), .B(n36545), .Z(n36550) );
  NAND U37185 ( .A(n36548), .B(n36547), .Z(n36549) );
  NAND U37186 ( .A(n36550), .B(n36549), .Z(n36746) );
  NAND U37187 ( .A(n36552), .B(n36551), .Z(n36556) );
  NAND U37188 ( .A(n36554), .B(n36553), .Z(n36555) );
  NAND U37189 ( .A(n36556), .B(n36555), .Z(n36707) );
  NAND U37190 ( .A(n36558), .B(n36557), .Z(n36562) );
  NAND U37191 ( .A(n36560), .B(n36559), .Z(n36561) );
  NAND U37192 ( .A(n36562), .B(n36561), .Z(n36706) );
  NAND U37193 ( .A(n38470), .B(n36566), .Z(n36568) );
  XOR U37194 ( .A(b[31]), .B(a[231]), .Z(n36687) );
  NAND U37195 ( .A(n38453), .B(n36687), .Z(n36567) );
  NAND U37196 ( .A(n36568), .B(n36567), .Z(n36695) );
  NAND U37197 ( .A(n190), .B(n36569), .Z(n36571) );
  XOR U37198 ( .A(b[19]), .B(a[243]), .Z(n36666) );
  NAND U37199 ( .A(n37821), .B(n36666), .Z(n36570) );
  NAND U37200 ( .A(n36571), .B(n36570), .Z(n36694) );
  AND U37201 ( .A(b[31]), .B(a[229]), .Z(n36726) );
  XNOR U37202 ( .A(n36572), .B(n36726), .Z(n36725) );
  XOR U37203 ( .A(n36724), .B(n36725), .Z(n36696) );
  XOR U37204 ( .A(n36697), .B(n36696), .Z(n36658) );
  NAND U37205 ( .A(n38185), .B(n36573), .Z(n36575) );
  XOR U37206 ( .A(b[23]), .B(a[239]), .Z(n36663) );
  NAND U37207 ( .A(n38132), .B(n36663), .Z(n36574) );
  NAND U37208 ( .A(n36575), .B(n36574), .Z(n36721) );
  NAND U37209 ( .A(n185), .B(n36576), .Z(n36578) );
  XOR U37210 ( .A(a[253]), .B(b[9]), .Z(n36681) );
  NAND U37211 ( .A(n36805), .B(n36681), .Z(n36577) );
  NAND U37212 ( .A(n36578), .B(n36577), .Z(n36719) );
  NAND U37213 ( .A(n38385), .B(n36579), .Z(n36581) );
  XOR U37214 ( .A(b[27]), .B(a[235]), .Z(n36669) );
  NAND U37215 ( .A(n38343), .B(n36669), .Z(n36580) );
  NAND U37216 ( .A(n36581), .B(n36580), .Z(n36718) );
  XOR U37217 ( .A(n36658), .B(n36657), .Z(n36659) );
  XOR U37218 ( .A(n36709), .B(n36708), .Z(n36648) );
  NAND U37219 ( .A(n36583), .B(n36582), .Z(n36587) );
  NANDN U37220 ( .A(n36585), .B(n36584), .Z(n36586) );
  NAND U37221 ( .A(n36587), .B(n36586), .Z(n36652) );
  NAND U37222 ( .A(n194), .B(n36588), .Z(n36590) );
  XOR U37223 ( .A(b[29]), .B(a[233]), .Z(n36672) );
  NAND U37224 ( .A(n38456), .B(n36672), .Z(n36589) );
  NAND U37225 ( .A(n36590), .B(n36589), .Z(n36742) );
  NAND U37226 ( .A(n184), .B(n36591), .Z(n36594) );
  XOR U37227 ( .A(a[255]), .B(b[7]), .Z(n36690) );
  NAND U37228 ( .A(n36592), .B(n36690), .Z(n36593) );
  NAND U37229 ( .A(n36594), .B(n36593), .Z(n36740) );
  NAND U37230 ( .A(n38064), .B(n36595), .Z(n36597) );
  XOR U37231 ( .A(b[21]), .B(a[241]), .Z(n36684) );
  NAND U37232 ( .A(n37993), .B(n36684), .Z(n36596) );
  NAND U37233 ( .A(n36597), .B(n36596), .Z(n36739) );
  NAND U37234 ( .A(n188), .B(n36598), .Z(n36600) );
  XOR U37235 ( .A(a[247]), .B(b[15]), .Z(n36730) );
  NAND U37236 ( .A(n37382), .B(n36730), .Z(n36599) );
  NAND U37237 ( .A(n36600), .B(n36599), .Z(n36715) );
  NAND U37238 ( .A(n187), .B(n36601), .Z(n36603) );
  XOR U37239 ( .A(a[249]), .B(b[13]), .Z(n36733) );
  NAND U37240 ( .A(n37295), .B(n36733), .Z(n36602) );
  NAND U37241 ( .A(n36603), .B(n36602), .Z(n36713) );
  NAND U37242 ( .A(n189), .B(n36604), .Z(n36606) );
  XOR U37243 ( .A(a[245]), .B(b[17]), .Z(n36675) );
  NAND U37244 ( .A(n37652), .B(n36675), .Z(n36605) );
  NAND U37245 ( .A(n36606), .B(n36605), .Z(n36703) );
  NAND U37246 ( .A(n38289), .B(n36607), .Z(n36609) );
  XOR U37247 ( .A(b[25]), .B(a[237]), .Z(n36736) );
  NAND U37248 ( .A(n38247), .B(n36736), .Z(n36608) );
  NAND U37249 ( .A(n36609), .B(n36608), .Z(n36701) );
  NAND U37250 ( .A(n186), .B(n36610), .Z(n36612) );
  XOR U37251 ( .A(a[251]), .B(b[11]), .Z(n36678) );
  NAND U37252 ( .A(n37097), .B(n36678), .Z(n36611) );
  NAND U37253 ( .A(n36612), .B(n36611), .Z(n36700) );
  XNOR U37254 ( .A(n36654), .B(n36653), .Z(n36646) );
  NAND U37255 ( .A(n36614), .B(n36613), .Z(n36618) );
  NAND U37256 ( .A(n36616), .B(n36615), .Z(n36617) );
  AND U37257 ( .A(n36618), .B(n36617), .Z(n36645) );
  XOR U37258 ( .A(n36648), .B(n36647), .Z(n36745) );
  XOR U37259 ( .A(n36748), .B(n36747), .Z(n36751) );
  XOR U37260 ( .A(n36752), .B(n36751), .Z(n36754) );
  NAND U37261 ( .A(n36620), .B(n36619), .Z(n36624) );
  NAND U37262 ( .A(n36622), .B(n36621), .Z(n36623) );
  AND U37263 ( .A(n36624), .B(n36623), .Z(n36753) );
  XNOR U37264 ( .A(n36754), .B(n36753), .Z(n36627) );
  XOR U37265 ( .A(n36630), .B(n36629), .Z(n36625) );
  XOR U37266 ( .A(n36626), .B(n36625), .Z(c[485]) );
  AND U37267 ( .A(n36626), .B(n36625), .Z(n36758) );
  NAND U37268 ( .A(n36628), .B(n36627), .Z(n36632) );
  NANDN U37269 ( .A(n36630), .B(n36629), .Z(n36631) );
  AND U37270 ( .A(n36632), .B(n36631), .Z(n36762) );
  NAND U37271 ( .A(n36634), .B(n36633), .Z(n36638) );
  NAND U37272 ( .A(n36636), .B(n36635), .Z(n36637) );
  NAND U37273 ( .A(n36638), .B(n36637), .Z(n36768) );
  NAND U37274 ( .A(n36640), .B(n36639), .Z(n36644) );
  NAND U37275 ( .A(n36642), .B(n36641), .Z(n36643) );
  NAND U37276 ( .A(n36644), .B(n36643), .Z(n36774) );
  NAND U37277 ( .A(n36646), .B(n36645), .Z(n36650) );
  NANDN U37278 ( .A(n36648), .B(n36647), .Z(n36649) );
  NAND U37279 ( .A(n36650), .B(n36649), .Z(n36772) );
  NAND U37280 ( .A(n36652), .B(n36651), .Z(n36656) );
  NAND U37281 ( .A(n36654), .B(n36653), .Z(n36655) );
  NAND U37282 ( .A(n36656), .B(n36655), .Z(n36874) );
  NAND U37283 ( .A(n36658), .B(n36657), .Z(n36662) );
  NAND U37284 ( .A(n36660), .B(n36659), .Z(n36661) );
  NAND U37285 ( .A(n36662), .B(n36661), .Z(n36872) );
  NAND U37286 ( .A(n38185), .B(n36663), .Z(n36665) );
  XOR U37287 ( .A(b[23]), .B(a[240]), .Z(n36817) );
  NAND U37288 ( .A(n38132), .B(n36817), .Z(n36664) );
  NAND U37289 ( .A(n36665), .B(n36664), .Z(n36850) );
  NAND U37290 ( .A(n190), .B(n36666), .Z(n36668) );
  XOR U37291 ( .A(a[244]), .B(b[19]), .Z(n36838) );
  NAND U37292 ( .A(n37821), .B(n36838), .Z(n36667) );
  NAND U37293 ( .A(n36668), .B(n36667), .Z(n36848) );
  NAND U37294 ( .A(n38385), .B(n36669), .Z(n36671) );
  XOR U37295 ( .A(b[27]), .B(a[236]), .Z(n36826) );
  NAND U37296 ( .A(n38343), .B(n36826), .Z(n36670) );
  NAND U37297 ( .A(n36671), .B(n36670), .Z(n36798) );
  NAND U37298 ( .A(n194), .B(n36672), .Z(n36674) );
  XOR U37299 ( .A(b[29]), .B(a[234]), .Z(n36811) );
  NAND U37300 ( .A(n38456), .B(n36811), .Z(n36673) );
  NAND U37301 ( .A(n36674), .B(n36673), .Z(n36796) );
  NAND U37302 ( .A(n189), .B(n36675), .Z(n36677) );
  XOR U37303 ( .A(a[246]), .B(b[17]), .Z(n36835) );
  NAND U37304 ( .A(n37652), .B(n36835), .Z(n36676) );
  NAND U37305 ( .A(n36677), .B(n36676), .Z(n36795) );
  NAND U37306 ( .A(n186), .B(n36678), .Z(n36680) );
  XOR U37307 ( .A(a[252]), .B(b[11]), .Z(n36829) );
  NAND U37308 ( .A(n37097), .B(n36829), .Z(n36679) );
  NAND U37309 ( .A(n36680), .B(n36679), .Z(n36792) );
  NAND U37310 ( .A(n185), .B(n36681), .Z(n36683) );
  XOR U37311 ( .A(a[254]), .B(b[9]), .Z(n36804) );
  NAND U37312 ( .A(n36805), .B(n36804), .Z(n36682) );
  NAND U37313 ( .A(n36683), .B(n36682), .Z(n36790) );
  NAND U37314 ( .A(n38064), .B(n36684), .Z(n36686) );
  XOR U37315 ( .A(b[21]), .B(a[242]), .Z(n36808) );
  NAND U37316 ( .A(n37993), .B(n36808), .Z(n36685) );
  NAND U37317 ( .A(n36686), .B(n36685), .Z(n36789) );
  NAND U37318 ( .A(n38470), .B(n36687), .Z(n36689) );
  XOR U37319 ( .A(b[31]), .B(a[232]), .Z(n36814) );
  NAND U37320 ( .A(n38453), .B(n36814), .Z(n36688) );
  AND U37321 ( .A(n36689), .B(n36688), .Z(n36803) );
  AND U37322 ( .A(b[31]), .B(a[230]), .Z(n36937) );
  AND U37323 ( .A(n36690), .B(n184), .Z(n36693) );
  XOR U37324 ( .A(b[6]), .B(b[5]), .Z(n36691) );
  NAND U37325 ( .A(b[7]), .B(n36691), .Z(n36692) );
  NANDN U37326 ( .A(n36693), .B(n36692), .Z(n36801) );
  XNOR U37327 ( .A(n36937), .B(n36801), .Z(n36802) );
  XOR U37328 ( .A(n36803), .B(n36802), .Z(n36865) );
  XOR U37329 ( .A(n36866), .B(n36865), .Z(n36868) );
  XNOR U37330 ( .A(n36867), .B(n36868), .Z(n36855) );
  NAND U37331 ( .A(n36695), .B(n36694), .Z(n36699) );
  NAND U37332 ( .A(n36697), .B(n36696), .Z(n36698) );
  NAND U37333 ( .A(n36699), .B(n36698), .Z(n36854) );
  NAND U37334 ( .A(n36701), .B(n36700), .Z(n36705) );
  NAND U37335 ( .A(n36703), .B(n36702), .Z(n36704) );
  NAND U37336 ( .A(n36705), .B(n36704), .Z(n36853) );
  XOR U37337 ( .A(n36855), .B(n36856), .Z(n36871) );
  NAND U37338 ( .A(n36707), .B(n36706), .Z(n36711) );
  NAND U37339 ( .A(n36709), .B(n36708), .Z(n36710) );
  AND U37340 ( .A(n36711), .B(n36710), .Z(n36778) );
  NAND U37341 ( .A(n36713), .B(n36712), .Z(n36717) );
  NAND U37342 ( .A(n36715), .B(n36714), .Z(n36716) );
  AND U37343 ( .A(n36717), .B(n36716), .Z(n36786) );
  NAND U37344 ( .A(n36719), .B(n36718), .Z(n36723) );
  NAND U37345 ( .A(n36721), .B(n36720), .Z(n36722) );
  NAND U37346 ( .A(n36723), .B(n36722), .Z(n36862) );
  AND U37347 ( .A(n36725), .B(n36724), .Z(n36729) );
  NAND U37348 ( .A(n36727), .B(n36726), .Z(n36728) );
  NANDN U37349 ( .A(n36729), .B(n36728), .Z(n36860) );
  NAND U37350 ( .A(n188), .B(n36730), .Z(n36732) );
  XOR U37351 ( .A(a[248]), .B(b[15]), .Z(n36844) );
  NAND U37352 ( .A(n37382), .B(n36844), .Z(n36731) );
  NAND U37353 ( .A(n36732), .B(n36731), .Z(n36823) );
  NAND U37354 ( .A(n187), .B(n36733), .Z(n36735) );
  XOR U37355 ( .A(a[250]), .B(b[13]), .Z(n36841) );
  NAND U37356 ( .A(n37295), .B(n36841), .Z(n36734) );
  NAND U37357 ( .A(n36735), .B(n36734), .Z(n36821) );
  NAND U37358 ( .A(n38289), .B(n36736), .Z(n36738) );
  XOR U37359 ( .A(b[25]), .B(a[238]), .Z(n36832) );
  NAND U37360 ( .A(n38247), .B(n36832), .Z(n36737) );
  NAND U37361 ( .A(n36738), .B(n36737), .Z(n36820) );
  NAND U37362 ( .A(n36740), .B(n36739), .Z(n36744) );
  NAND U37363 ( .A(n36742), .B(n36741), .Z(n36743) );
  AND U37364 ( .A(n36744), .B(n36743), .Z(n36784) );
  XOR U37365 ( .A(n36783), .B(n36784), .Z(n36785) );
  XOR U37366 ( .A(n36786), .B(n36785), .Z(n36777) );
  XOR U37367 ( .A(n36778), .B(n36777), .Z(n36780) );
  XOR U37368 ( .A(n36779), .B(n36780), .Z(n36771) );
  NAND U37369 ( .A(n36746), .B(n36745), .Z(n36750) );
  NAND U37370 ( .A(n36748), .B(n36747), .Z(n36749) );
  NAND U37371 ( .A(n36750), .B(n36749), .Z(n36765) );
  XOR U37372 ( .A(n36766), .B(n36765), .Z(n36767) );
  NAND U37373 ( .A(n36752), .B(n36751), .Z(n36756) );
  NAND U37374 ( .A(n36754), .B(n36753), .Z(n36755) );
  AND U37375 ( .A(n36756), .B(n36755), .Z(n36760) );
  XOR U37376 ( .A(n36759), .B(n36760), .Z(n36761) );
  XOR U37377 ( .A(n36762), .B(n36761), .Z(n36757) );
  XOR U37378 ( .A(n36758), .B(n36757), .Z(c[486]) );
  AND U37379 ( .A(n36758), .B(n36757), .Z(n36878) );
  NAND U37380 ( .A(n36760), .B(n36759), .Z(n36764) );
  NANDN U37381 ( .A(n36762), .B(n36761), .Z(n36763) );
  AND U37382 ( .A(n36764), .B(n36763), .Z(n36882) );
  NAND U37383 ( .A(n36766), .B(n36765), .Z(n36770) );
  NAND U37384 ( .A(n36768), .B(n36767), .Z(n36769) );
  AND U37385 ( .A(n36770), .B(n36769), .Z(n36880) );
  NAND U37386 ( .A(n36772), .B(n36771), .Z(n36776) );
  NAND U37387 ( .A(n36774), .B(n36773), .Z(n36775) );
  NAND U37388 ( .A(n36776), .B(n36775), .Z(n36888) );
  NAND U37389 ( .A(n36778), .B(n36777), .Z(n36782) );
  NAND U37390 ( .A(n36780), .B(n36779), .Z(n36781) );
  NAND U37391 ( .A(n36782), .B(n36781), .Z(n36886) );
  NAND U37392 ( .A(n36784), .B(n36783), .Z(n36788) );
  NAND U37393 ( .A(n36786), .B(n36785), .Z(n36787) );
  NAND U37394 ( .A(n36788), .B(n36787), .Z(n36998) );
  NAND U37395 ( .A(n36790), .B(n36789), .Z(n36794) );
  NAND U37396 ( .A(n36792), .B(n36791), .Z(n36793) );
  NAND U37397 ( .A(n36794), .B(n36793), .Z(n36972) );
  NAND U37398 ( .A(n36796), .B(n36795), .Z(n36800) );
  NAND U37399 ( .A(n36798), .B(n36797), .Z(n36799) );
  NAND U37400 ( .A(n36800), .B(n36799), .Z(n36971) );
  NAND U37401 ( .A(n185), .B(n36804), .Z(n36807) );
  XOR U37402 ( .A(a[255]), .B(b[9]), .Z(n36943) );
  NAND U37403 ( .A(n36805), .B(n36943), .Z(n36806) );
  NAND U37404 ( .A(n36807), .B(n36806), .Z(n36960) );
  NAND U37405 ( .A(n38064), .B(n36808), .Z(n36810) );
  XOR U37406 ( .A(b[21]), .B(a[243]), .Z(n36956) );
  NAND U37407 ( .A(n37993), .B(n36956), .Z(n36809) );
  NAND U37408 ( .A(n36810), .B(n36809), .Z(n36959) );
  AND U37409 ( .A(b[31]), .B(a[231]), .Z(n36940) );
  XOR U37410 ( .A(n36939), .B(n36940), .Z(n36938) );
  XOR U37411 ( .A(n36937), .B(n36938), .Z(n36961) );
  XOR U37412 ( .A(n36962), .B(n36961), .Z(n36984) );
  NAND U37413 ( .A(n194), .B(n36811), .Z(n36813) );
  XOR U37414 ( .A(b[29]), .B(a[235]), .Z(n36953) );
  NAND U37415 ( .A(n38456), .B(n36953), .Z(n36812) );
  NAND U37416 ( .A(n36813), .B(n36812), .Z(n36928) );
  NAND U37417 ( .A(n38470), .B(n36814), .Z(n36816) );
  XOR U37418 ( .A(b[31]), .B(a[233]), .Z(n36947) );
  NAND U37419 ( .A(n38453), .B(n36947), .Z(n36815) );
  NAND U37420 ( .A(n36816), .B(n36815), .Z(n36926) );
  NAND U37421 ( .A(n38185), .B(n36817), .Z(n36819) );
  XOR U37422 ( .A(b[23]), .B(a[241]), .Z(n36909) );
  NAND U37423 ( .A(n38132), .B(n36909), .Z(n36818) );
  NAND U37424 ( .A(n36819), .B(n36818), .Z(n36925) );
  XOR U37425 ( .A(n36984), .B(n36983), .Z(n36985) );
  XNOR U37426 ( .A(n36974), .B(n36973), .Z(n36996) );
  NAND U37427 ( .A(n36821), .B(n36820), .Z(n36825) );
  NAND U37428 ( .A(n36823), .B(n36822), .Z(n36824) );
  AND U37429 ( .A(n36825), .B(n36824), .Z(n36898) );
  NAND U37430 ( .A(n38385), .B(n36826), .Z(n36828) );
  XOR U37431 ( .A(b[27]), .B(a[237]), .Z(n36906) );
  NAND U37432 ( .A(n38343), .B(n36906), .Z(n36827) );
  NAND U37433 ( .A(n36828), .B(n36827), .Z(n36934) );
  NAND U37434 ( .A(n186), .B(n36829), .Z(n36831) );
  XOR U37435 ( .A(a[253]), .B(b[11]), .Z(n36950) );
  NAND U37436 ( .A(n37097), .B(n36950), .Z(n36830) );
  NAND U37437 ( .A(n36831), .B(n36830), .Z(n36932) );
  NAND U37438 ( .A(n38289), .B(n36832), .Z(n36834) );
  XOR U37439 ( .A(b[25]), .B(a[239]), .Z(n36903) );
  NAND U37440 ( .A(n38247), .B(n36903), .Z(n36833) );
  NAND U37441 ( .A(n36834), .B(n36833), .Z(n36931) );
  NAND U37442 ( .A(n189), .B(n36835), .Z(n36837) );
  XNOR U37443 ( .A(a[247]), .B(b[17]), .Z(n36921) );
  OR U37444 ( .A(n36921), .B(n36922), .Z(n36836) );
  NAND U37445 ( .A(n36837), .B(n36836), .Z(n36968) );
  NAND U37446 ( .A(n190), .B(n36838), .Z(n36840) );
  XOR U37447 ( .A(b[19]), .B(a[245]), .Z(n36915) );
  NAND U37448 ( .A(n37821), .B(n36915), .Z(n36839) );
  NAND U37449 ( .A(n36840), .B(n36839), .Z(n36966) );
  NAND U37450 ( .A(n187), .B(n36841), .Z(n36843) );
  XOR U37451 ( .A(a[251]), .B(b[13]), .Z(n36918) );
  NAND U37452 ( .A(n37295), .B(n36918), .Z(n36842) );
  NAND U37453 ( .A(n36843), .B(n36842), .Z(n36965) );
  NANDN U37454 ( .A(n178), .B(n36844), .Z(n36846) );
  XOR U37455 ( .A(a[249]), .B(b[15]), .Z(n36912) );
  NANDN U37456 ( .A(n37509), .B(n36912), .Z(n36845) );
  AND U37457 ( .A(n36846), .B(n36845), .Z(n36978) );
  XOR U37458 ( .A(n36977), .B(n36978), .Z(n36980) );
  XOR U37459 ( .A(n36979), .B(n36980), .Z(n36897) );
  XOR U37460 ( .A(n36898), .B(n36897), .Z(n36899) );
  NAND U37461 ( .A(n36848), .B(n36847), .Z(n36852) );
  NAND U37462 ( .A(n36850), .B(n36849), .Z(n36851) );
  AND U37463 ( .A(n36852), .B(n36851), .Z(n36900) );
  NAND U37464 ( .A(n36854), .B(n36853), .Z(n36858) );
  NAND U37465 ( .A(n36856), .B(n36855), .Z(n36857) );
  NAND U37466 ( .A(n36858), .B(n36857), .Z(n36992) );
  NAND U37467 ( .A(n36860), .B(n36859), .Z(n36864) );
  NAND U37468 ( .A(n36862), .B(n36861), .Z(n36863) );
  NAND U37469 ( .A(n36864), .B(n36863), .Z(n36990) );
  NAND U37470 ( .A(n36866), .B(n36865), .Z(n36870) );
  NAND U37471 ( .A(n36868), .B(n36867), .Z(n36869) );
  AND U37472 ( .A(n36870), .B(n36869), .Z(n36989) );
  NAND U37473 ( .A(n36872), .B(n36871), .Z(n36876) );
  NAND U37474 ( .A(n36874), .B(n36873), .Z(n36875) );
  AND U37475 ( .A(n36876), .B(n36875), .Z(n36892) );
  XOR U37476 ( .A(n36891), .B(n36892), .Z(n36893) );
  XOR U37477 ( .A(n36894), .B(n36893), .Z(n36885) );
  XOR U37478 ( .A(n36880), .B(n36879), .Z(n36881) );
  XOR U37479 ( .A(n36882), .B(n36881), .Z(n36877) );
  XOR U37480 ( .A(n36878), .B(n36877), .Z(c[487]) );
  AND U37481 ( .A(n36878), .B(n36877), .Z(n37002) );
  NAND U37482 ( .A(n36880), .B(n36879), .Z(n36884) );
  NANDN U37483 ( .A(n36882), .B(n36881), .Z(n36883) );
  AND U37484 ( .A(n36884), .B(n36883), .Z(n37006) );
  NAND U37485 ( .A(n36886), .B(n36885), .Z(n36890) );
  NAND U37486 ( .A(n36888), .B(n36887), .Z(n36889) );
  NAND U37487 ( .A(n36890), .B(n36889), .Z(n37004) );
  NAND U37488 ( .A(n36892), .B(n36891), .Z(n36896) );
  NAND U37489 ( .A(n36894), .B(n36893), .Z(n36895) );
  NAND U37490 ( .A(n36896), .B(n36895), .Z(n37012) );
  NAND U37491 ( .A(n36898), .B(n36897), .Z(n36902) );
  NAND U37492 ( .A(n36900), .B(n36899), .Z(n36901) );
  NAND U37493 ( .A(n36902), .B(n36901), .Z(n37024) );
  NAND U37494 ( .A(n38289), .B(n36903), .Z(n36905) );
  XOR U37495 ( .A(b[25]), .B(a[240]), .Z(n37075) );
  NAND U37496 ( .A(n38247), .B(n37075), .Z(n36904) );
  NAND U37497 ( .A(n36905), .B(n36904), .Z(n37054) );
  NAND U37498 ( .A(n38385), .B(n36906), .Z(n36908) );
  XOR U37499 ( .A(b[27]), .B(a[238]), .Z(n37078) );
  NAND U37500 ( .A(n38343), .B(n37078), .Z(n36907) );
  NAND U37501 ( .A(n36908), .B(n36907), .Z(n37052) );
  NAND U37502 ( .A(n38185), .B(n36909), .Z(n36911) );
  XOR U37503 ( .A(b[23]), .B(a[242]), .Z(n37100) );
  NAND U37504 ( .A(n38132), .B(n37100), .Z(n36910) );
  NAND U37505 ( .A(n36911), .B(n36910), .Z(n37051) );
  NAND U37506 ( .A(n188), .B(n36912), .Z(n36914) );
  XOR U37507 ( .A(a[250]), .B(b[15]), .Z(n37090) );
  NAND U37508 ( .A(n37382), .B(n37090), .Z(n36913) );
  NAND U37509 ( .A(n36914), .B(n36913), .Z(n37106) );
  NAND U37510 ( .A(n190), .B(n36915), .Z(n36917) );
  XOR U37511 ( .A(a[246]), .B(b[19]), .Z(n37081) );
  NAND U37512 ( .A(n37821), .B(n37081), .Z(n36916) );
  NAND U37513 ( .A(n36917), .B(n36916), .Z(n37104) );
  NAND U37514 ( .A(n187), .B(n36918), .Z(n36920) );
  XOR U37515 ( .A(a[252]), .B(b[13]), .Z(n37093) );
  NAND U37516 ( .A(n37295), .B(n37093), .Z(n36919) );
  NAND U37517 ( .A(n36920), .B(n36919), .Z(n37103) );
  OR U37518 ( .A(n36921), .B(n170), .Z(n36924) );
  XOR U37519 ( .A(a[248]), .B(b[17]), .Z(n37087) );
  NANDN U37520 ( .A(n36922), .B(n37087), .Z(n36923) );
  AND U37521 ( .A(n36924), .B(n36923), .Z(n37040) );
  XOR U37522 ( .A(n37039), .B(n37040), .Z(n37042) );
  XNOR U37523 ( .A(n37041), .B(n37042), .Z(n37029) );
  NAND U37524 ( .A(n36926), .B(n36925), .Z(n36930) );
  NAND U37525 ( .A(n36928), .B(n36927), .Z(n36929) );
  NAND U37526 ( .A(n36930), .B(n36929), .Z(n37028) );
  NAND U37527 ( .A(n36932), .B(n36931), .Z(n36936) );
  NAND U37528 ( .A(n36934), .B(n36933), .Z(n36935) );
  NAND U37529 ( .A(n36936), .B(n36935), .Z(n37048) );
  AND U37530 ( .A(n36938), .B(n36937), .Z(n36942) );
  NAND U37531 ( .A(n36940), .B(n36939), .Z(n36941) );
  NANDN U37532 ( .A(n36942), .B(n36941), .Z(n37046) );
  AND U37533 ( .A(n36943), .B(n185), .Z(n36946) );
  XOR U37534 ( .A(b[8]), .B(b[7]), .Z(n36944) );
  NAND U37535 ( .A(b[9]), .B(n36944), .Z(n36945) );
  NANDN U37536 ( .A(n36946), .B(n36945), .Z(n37059) );
  AND U37537 ( .A(b[31]), .B(a[232]), .Z(n37206) );
  NAND U37538 ( .A(n38470), .B(n36947), .Z(n36949) );
  XOR U37539 ( .A(b[31]), .B(a[234]), .Z(n37068) );
  NAND U37540 ( .A(n38453), .B(n37068), .Z(n36948) );
  NAND U37541 ( .A(n36949), .B(n36948), .Z(n37057) );
  XNOR U37542 ( .A(n37206), .B(n37057), .Z(n37058) );
  XNOR U37543 ( .A(n37029), .B(n37030), .Z(n37021) );
  NAND U37544 ( .A(n186), .B(n36950), .Z(n36952) );
  XOR U37545 ( .A(a[254]), .B(b[11]), .Z(n37096) );
  NAND U37546 ( .A(n37097), .B(n37096), .Z(n36951) );
  NAND U37547 ( .A(n36952), .B(n36951), .Z(n37065) );
  NAND U37548 ( .A(n194), .B(n36953), .Z(n36955) );
  XOR U37549 ( .A(b[29]), .B(a[236]), .Z(n37084) );
  NAND U37550 ( .A(n38456), .B(n37084), .Z(n36954) );
  NAND U37551 ( .A(n36955), .B(n36954), .Z(n37063) );
  NAND U37552 ( .A(n38064), .B(n36956), .Z(n36958) );
  XOR U37553 ( .A(b[21]), .B(a[244]), .Z(n37071) );
  NAND U37554 ( .A(n37993), .B(n37071), .Z(n36957) );
  NAND U37555 ( .A(n36958), .B(n36957), .Z(n37062) );
  NAND U37556 ( .A(n36960), .B(n36959), .Z(n36964) );
  NAND U37557 ( .A(n36962), .B(n36961), .Z(n36963) );
  AND U37558 ( .A(n36964), .B(n36963), .Z(n37034) );
  XOR U37559 ( .A(n37033), .B(n37034), .Z(n37035) );
  NAND U37560 ( .A(n36966), .B(n36965), .Z(n36970) );
  NAND U37561 ( .A(n36968), .B(n36967), .Z(n36969) );
  AND U37562 ( .A(n36970), .B(n36969), .Z(n37036) );
  XOR U37563 ( .A(n37021), .B(n37022), .Z(n37023) );
  NAND U37564 ( .A(n36972), .B(n36971), .Z(n36976) );
  NAND U37565 ( .A(n36974), .B(n36973), .Z(n36975) );
  AND U37566 ( .A(n36976), .B(n36975), .Z(n37112) );
  NAND U37567 ( .A(n36978), .B(n36977), .Z(n36982) );
  NAND U37568 ( .A(n36980), .B(n36979), .Z(n36981) );
  NAND U37569 ( .A(n36982), .B(n36981), .Z(n37110) );
  NAND U37570 ( .A(n36984), .B(n36983), .Z(n36988) );
  NAND U37571 ( .A(n36986), .B(n36985), .Z(n36987) );
  AND U37572 ( .A(n36988), .B(n36987), .Z(n37109) );
  XNOR U37573 ( .A(n37112), .B(n37111), .Z(n37016) );
  NAND U37574 ( .A(n36990), .B(n36989), .Z(n36994) );
  NAND U37575 ( .A(n36992), .B(n36991), .Z(n36993) );
  NAND U37576 ( .A(n36994), .B(n36993), .Z(n37015) );
  XNOR U37577 ( .A(n37017), .B(n37018), .Z(n37010) );
  NAND U37578 ( .A(n36996), .B(n36995), .Z(n37000) );
  NAND U37579 ( .A(n36998), .B(n36997), .Z(n36999) );
  NAND U37580 ( .A(n37000), .B(n36999), .Z(n37009) );
  XOR U37581 ( .A(n37010), .B(n37009), .Z(n37011) );
  XOR U37582 ( .A(n37006), .B(n37005), .Z(n37001) );
  XOR U37583 ( .A(n37002), .B(n37001), .Z(c[488]) );
  AND U37584 ( .A(n37002), .B(n37001), .Z(n37116) );
  NAND U37585 ( .A(n37004), .B(n37003), .Z(n37008) );
  NANDN U37586 ( .A(n37006), .B(n37005), .Z(n37007) );
  AND U37587 ( .A(n37008), .B(n37007), .Z(n37120) );
  NAND U37588 ( .A(n37010), .B(n37009), .Z(n37014) );
  NAND U37589 ( .A(n37012), .B(n37011), .Z(n37013) );
  NAND U37590 ( .A(n37014), .B(n37013), .Z(n37118) );
  NAND U37591 ( .A(n37016), .B(n37015), .Z(n37020) );
  NAND U37592 ( .A(n37018), .B(n37017), .Z(n37019) );
  AND U37593 ( .A(n37020), .B(n37019), .Z(n37126) );
  NAND U37594 ( .A(n37022), .B(n37021), .Z(n37026) );
  NAND U37595 ( .A(n37024), .B(n37023), .Z(n37025) );
  NAND U37596 ( .A(n37026), .B(n37025), .Z(n37124) );
  NAND U37597 ( .A(n37028), .B(n37027), .Z(n37032) );
  NAND U37598 ( .A(n37030), .B(n37029), .Z(n37031) );
  AND U37599 ( .A(n37032), .B(n37031), .Z(n37226) );
  NAND U37600 ( .A(n37034), .B(n37033), .Z(n37038) );
  NAND U37601 ( .A(n37036), .B(n37035), .Z(n37037) );
  NAND U37602 ( .A(n37038), .B(n37037), .Z(n37224) );
  NAND U37603 ( .A(n37040), .B(n37039), .Z(n37044) );
  NAND U37604 ( .A(n37042), .B(n37041), .Z(n37043) );
  NAND U37605 ( .A(n37044), .B(n37043), .Z(n37223) );
  XOR U37606 ( .A(n37226), .B(n37225), .Z(n37132) );
  NAND U37607 ( .A(n37046), .B(n37045), .Z(n37050) );
  NAND U37608 ( .A(n37048), .B(n37047), .Z(n37049) );
  AND U37609 ( .A(n37050), .B(n37049), .Z(n37138) );
  NAND U37610 ( .A(n37052), .B(n37051), .Z(n37056) );
  NAND U37611 ( .A(n37054), .B(n37053), .Z(n37055) );
  NAND U37612 ( .A(n37056), .B(n37055), .Z(n37218) );
  IV U37613 ( .A(n37206), .Z(n37074) );
  NAND U37614 ( .A(n37074), .B(n37057), .Z(n37061) );
  NAND U37615 ( .A(n37059), .B(n37058), .Z(n37060) );
  NAND U37616 ( .A(n37061), .B(n37060), .Z(n37217) );
  NAND U37617 ( .A(n37063), .B(n37062), .Z(n37067) );
  NAND U37618 ( .A(n37065), .B(n37064), .Z(n37066) );
  NAND U37619 ( .A(n37067), .B(n37066), .Z(n37190) );
  NAND U37620 ( .A(n38470), .B(n37068), .Z(n37070) );
  XOR U37621 ( .A(b[31]), .B(a[235]), .Z(n37147) );
  NAND U37622 ( .A(n38453), .B(n37147), .Z(n37069) );
  NAND U37623 ( .A(n37070), .B(n37069), .Z(n37142) );
  NAND U37624 ( .A(n38064), .B(n37071), .Z(n37073) );
  XOR U37625 ( .A(b[21]), .B(a[245]), .Z(n37157) );
  NAND U37626 ( .A(n37993), .B(n37157), .Z(n37072) );
  NAND U37627 ( .A(n37073), .B(n37072), .Z(n37141) );
  XNOR U37628 ( .A(n37074), .B(n37205), .Z(n37208) );
  AND U37629 ( .A(b[31]), .B(a[233]), .Z(n37207) );
  XOR U37630 ( .A(n37208), .B(n37207), .Z(n37143) );
  XOR U37631 ( .A(n37144), .B(n37143), .Z(n37188) );
  NAND U37632 ( .A(n38289), .B(n37075), .Z(n37077) );
  XOR U37633 ( .A(b[25]), .B(a[241]), .Z(n37154) );
  NAND U37634 ( .A(n38247), .B(n37154), .Z(n37076) );
  NAND U37635 ( .A(n37077), .B(n37076), .Z(n37184) );
  NAND U37636 ( .A(n38385), .B(n37078), .Z(n37080) );
  XOR U37637 ( .A(b[27]), .B(a[239]), .Z(n37169) );
  NAND U37638 ( .A(n38343), .B(n37169), .Z(n37079) );
  NAND U37639 ( .A(n37080), .B(n37079), .Z(n37182) );
  NAND U37640 ( .A(n190), .B(n37081), .Z(n37083) );
  XOR U37641 ( .A(a[247]), .B(b[19]), .Z(n37160) );
  NAND U37642 ( .A(n37821), .B(n37160), .Z(n37082) );
  NAND U37643 ( .A(n37083), .B(n37082), .Z(n37181) );
  XOR U37644 ( .A(n37188), .B(n37187), .Z(n37189) );
  XNOR U37645 ( .A(n37220), .B(n37219), .Z(n37136) );
  NAND U37646 ( .A(n194), .B(n37084), .Z(n37086) );
  XOR U37647 ( .A(b[29]), .B(a[237]), .Z(n37163) );
  NAND U37648 ( .A(n38456), .B(n37163), .Z(n37085) );
  NAND U37649 ( .A(n37086), .B(n37085), .Z(n37202) );
  NAND U37650 ( .A(n189), .B(n37087), .Z(n37089) );
  XOR U37651 ( .A(a[249]), .B(b[17]), .Z(n37166) );
  NAND U37652 ( .A(n37652), .B(n37166), .Z(n37088) );
  NAND U37653 ( .A(n37089), .B(n37088), .Z(n37200) );
  NAND U37654 ( .A(n188), .B(n37090), .Z(n37092) );
  XOR U37655 ( .A(a[251]), .B(b[15]), .Z(n37175) );
  NAND U37656 ( .A(n37382), .B(n37175), .Z(n37091) );
  NAND U37657 ( .A(n37092), .B(n37091), .Z(n37199) );
  NAND U37658 ( .A(n187), .B(n37093), .Z(n37095) );
  XOR U37659 ( .A(a[253]), .B(b[13]), .Z(n37178) );
  NAND U37660 ( .A(n37295), .B(n37178), .Z(n37094) );
  AND U37661 ( .A(n37095), .B(n37094), .Z(n37214) );
  NAND U37662 ( .A(n186), .B(n37096), .Z(n37099) );
  XOR U37663 ( .A(a[255]), .B(b[11]), .Z(n37150) );
  NAND U37664 ( .A(n37097), .B(n37150), .Z(n37098) );
  NAND U37665 ( .A(n37099), .B(n37098), .Z(n37212) );
  NAND U37666 ( .A(n38185), .B(n37100), .Z(n37102) );
  XOR U37667 ( .A(b[23]), .B(a[243]), .Z(n37172) );
  NAND U37668 ( .A(n38132), .B(n37172), .Z(n37101) );
  NAND U37669 ( .A(n37102), .B(n37101), .Z(n37211) );
  XOR U37670 ( .A(n37214), .B(n37213), .Z(n37193) );
  XOR U37671 ( .A(n37194), .B(n37193), .Z(n37195) );
  NAND U37672 ( .A(n37104), .B(n37103), .Z(n37108) );
  NAND U37673 ( .A(n37106), .B(n37105), .Z(n37107) );
  AND U37674 ( .A(n37108), .B(n37107), .Z(n37196) );
  XNOR U37675 ( .A(n37138), .B(n37137), .Z(n37130) );
  NAND U37676 ( .A(n37110), .B(n37109), .Z(n37114) );
  NAND U37677 ( .A(n37112), .B(n37111), .Z(n37113) );
  AND U37678 ( .A(n37114), .B(n37113), .Z(n37129) );
  XOR U37679 ( .A(n37132), .B(n37131), .Z(n37123) );
  XOR U37680 ( .A(n37126), .B(n37125), .Z(n37117) );
  XOR U37681 ( .A(n37120), .B(n37119), .Z(n37115) );
  XOR U37682 ( .A(n37116), .B(n37115), .Z(c[489]) );
  AND U37683 ( .A(n37116), .B(n37115), .Z(n37230) );
  NAND U37684 ( .A(n37118), .B(n37117), .Z(n37122) );
  NANDN U37685 ( .A(n37120), .B(n37119), .Z(n37121) );
  AND U37686 ( .A(n37122), .B(n37121), .Z(n37234) );
  NAND U37687 ( .A(n37124), .B(n37123), .Z(n37128) );
  NAND U37688 ( .A(n37126), .B(n37125), .Z(n37127) );
  NAND U37689 ( .A(n37128), .B(n37127), .Z(n37232) );
  NAND U37690 ( .A(n37130), .B(n37129), .Z(n37134) );
  NANDN U37691 ( .A(n37132), .B(n37131), .Z(n37133) );
  AND U37692 ( .A(n37134), .B(n37133), .Z(n37328) );
  NAND U37693 ( .A(n37136), .B(n37135), .Z(n37140) );
  NAND U37694 ( .A(n37138), .B(n37137), .Z(n37139) );
  NAND U37695 ( .A(n37140), .B(n37139), .Z(n37322) );
  NAND U37696 ( .A(n37142), .B(n37141), .Z(n37146) );
  NAND U37697 ( .A(n37144), .B(n37143), .Z(n37145) );
  NAND U37698 ( .A(n37146), .B(n37145), .Z(n37252) );
  NAND U37699 ( .A(n38470), .B(n37147), .Z(n37149) );
  XOR U37700 ( .A(b[31]), .B(a[236]), .Z(n37302) );
  NAND U37701 ( .A(n38453), .B(n37302), .Z(n37148) );
  NAND U37702 ( .A(n37149), .B(n37148), .Z(n37290) );
  AND U37703 ( .A(b[31]), .B(a[234]), .Z(n37389) );
  AND U37704 ( .A(n37150), .B(n186), .Z(n37153) );
  XOR U37705 ( .A(b[10]), .B(b[9]), .Z(n37151) );
  NAND U37706 ( .A(b[11]), .B(n37151), .Z(n37152) );
  NANDN U37707 ( .A(n37153), .B(n37152), .Z(n37288) );
  XNOR U37708 ( .A(n37389), .B(n37288), .Z(n37289) );
  NAND U37709 ( .A(n38289), .B(n37154), .Z(n37156) );
  XOR U37710 ( .A(b[25]), .B(a[242]), .Z(n37285) );
  NAND U37711 ( .A(n38247), .B(n37285), .Z(n37155) );
  NAND U37712 ( .A(n37156), .B(n37155), .Z(n37264) );
  NAND U37713 ( .A(n38064), .B(n37157), .Z(n37159) );
  XOR U37714 ( .A(b[21]), .B(a[246]), .Z(n37298) );
  NAND U37715 ( .A(n37993), .B(n37298), .Z(n37158) );
  NAND U37716 ( .A(n37159), .B(n37158), .Z(n37262) );
  NAND U37717 ( .A(n190), .B(n37160), .Z(n37162) );
  XOR U37718 ( .A(a[248]), .B(b[19]), .Z(n37279) );
  NAND U37719 ( .A(n37821), .B(n37279), .Z(n37161) );
  NAND U37720 ( .A(n37162), .B(n37161), .Z(n37261) );
  XOR U37721 ( .A(n37250), .B(n37249), .Z(n37251) );
  NAND U37722 ( .A(n194), .B(n37163), .Z(n37165) );
  XOR U37723 ( .A(b[29]), .B(a[238]), .Z(n37291) );
  NAND U37724 ( .A(n38456), .B(n37291), .Z(n37164) );
  NAND U37725 ( .A(n37165), .B(n37164), .Z(n37258) );
  NAND U37726 ( .A(n189), .B(n37166), .Z(n37168) );
  XOR U37727 ( .A(a[250]), .B(b[17]), .Z(n37273) );
  NAND U37728 ( .A(n37652), .B(n37273), .Z(n37167) );
  NAND U37729 ( .A(n37168), .B(n37167), .Z(n37256) );
  NAND U37730 ( .A(n38385), .B(n37169), .Z(n37171) );
  XOR U37731 ( .A(b[27]), .B(a[240]), .Z(n37282) );
  NAND U37732 ( .A(n38343), .B(n37282), .Z(n37170) );
  NAND U37733 ( .A(n37171), .B(n37170), .Z(n37255) );
  NAND U37734 ( .A(n38185), .B(n37172), .Z(n37174) );
  XOR U37735 ( .A(b[23]), .B(a[244]), .Z(n37305) );
  NAND U37736 ( .A(n38132), .B(n37305), .Z(n37173) );
  AND U37737 ( .A(n37174), .B(n37173), .Z(n37270) );
  NAND U37738 ( .A(n188), .B(n37175), .Z(n37177) );
  XOR U37739 ( .A(a[252]), .B(b[15]), .Z(n37276) );
  NAND U37740 ( .A(n37382), .B(n37276), .Z(n37176) );
  NAND U37741 ( .A(n37177), .B(n37176), .Z(n37268) );
  NAND U37742 ( .A(n187), .B(n37178), .Z(n37180) );
  XOR U37743 ( .A(a[254]), .B(b[13]), .Z(n37294) );
  NAND U37744 ( .A(n37295), .B(n37294), .Z(n37179) );
  NAND U37745 ( .A(n37180), .B(n37179), .Z(n37267) );
  XOR U37746 ( .A(n37270), .B(n37269), .Z(n37243) );
  XOR U37747 ( .A(n37244), .B(n37243), .Z(n37245) );
  NAND U37748 ( .A(n37182), .B(n37181), .Z(n37186) );
  NAND U37749 ( .A(n37184), .B(n37183), .Z(n37185) );
  AND U37750 ( .A(n37186), .B(n37185), .Z(n37246) );
  XOR U37751 ( .A(n37307), .B(n37308), .Z(n37309) );
  NAND U37752 ( .A(n37188), .B(n37187), .Z(n37192) );
  NAND U37753 ( .A(n37190), .B(n37189), .Z(n37191) );
  AND U37754 ( .A(n37192), .B(n37191), .Z(n37310) );
  NAND U37755 ( .A(n37194), .B(n37193), .Z(n37198) );
  NAND U37756 ( .A(n37196), .B(n37195), .Z(n37197) );
  NAND U37757 ( .A(n37198), .B(n37197), .Z(n37238) );
  NAND U37758 ( .A(n37200), .B(n37199), .Z(n37204) );
  NAND U37759 ( .A(n37202), .B(n37201), .Z(n37203) );
  AND U37760 ( .A(n37204), .B(n37203), .Z(n37316) );
  NAND U37761 ( .A(n37206), .B(n37205), .Z(n37210) );
  NAND U37762 ( .A(n37208), .B(n37207), .Z(n37209) );
  AND U37763 ( .A(n37210), .B(n37209), .Z(n37313) );
  NAND U37764 ( .A(n37212), .B(n37211), .Z(n37216) );
  NANDN U37765 ( .A(n37214), .B(n37213), .Z(n37215) );
  AND U37766 ( .A(n37216), .B(n37215), .Z(n37314) );
  XOR U37767 ( .A(n37316), .B(n37315), .Z(n37237) );
  XOR U37768 ( .A(n37240), .B(n37239), .Z(n37319) );
  NAND U37769 ( .A(n37218), .B(n37217), .Z(n37222) );
  NAND U37770 ( .A(n37220), .B(n37219), .Z(n37221) );
  AND U37771 ( .A(n37222), .B(n37221), .Z(n37320) );
  NAND U37772 ( .A(n37224), .B(n37223), .Z(n37228) );
  NAND U37773 ( .A(n37226), .B(n37225), .Z(n37227) );
  AND U37774 ( .A(n37228), .B(n37227), .Z(n37326) );
  XOR U37775 ( .A(n37325), .B(n37326), .Z(n37327) );
  XOR U37776 ( .A(n37328), .B(n37327), .Z(n37231) );
  XOR U37777 ( .A(n37234), .B(n37233), .Z(n37229) );
  XOR U37778 ( .A(n37230), .B(n37229), .Z(c[490]) );
  AND U37779 ( .A(n37230), .B(n37229), .Z(n37332) );
  NAND U37780 ( .A(n37232), .B(n37231), .Z(n37236) );
  NANDN U37781 ( .A(n37234), .B(n37233), .Z(n37235) );
  AND U37782 ( .A(n37236), .B(n37235), .Z(n37336) );
  NAND U37783 ( .A(n37238), .B(n37237), .Z(n37242) );
  NAND U37784 ( .A(n37240), .B(n37239), .Z(n37241) );
  AND U37785 ( .A(n37242), .B(n37241), .Z(n37340) );
  NAND U37786 ( .A(n37244), .B(n37243), .Z(n37248) );
  NAND U37787 ( .A(n37246), .B(n37245), .Z(n37247) );
  NAND U37788 ( .A(n37248), .B(n37247), .Z(n37352) );
  NAND U37789 ( .A(n37250), .B(n37249), .Z(n37254) );
  NAND U37790 ( .A(n37252), .B(n37251), .Z(n37253) );
  AND U37791 ( .A(n37254), .B(n37253), .Z(n37351) );
  NAND U37792 ( .A(n37256), .B(n37255), .Z(n37260) );
  NAND U37793 ( .A(n37258), .B(n37257), .Z(n37259) );
  AND U37794 ( .A(n37260), .B(n37259), .Z(n37428) );
  NAND U37795 ( .A(n37262), .B(n37261), .Z(n37266) );
  NAND U37796 ( .A(n37264), .B(n37263), .Z(n37265) );
  AND U37797 ( .A(n37266), .B(n37265), .Z(n37426) );
  NAND U37798 ( .A(n37268), .B(n37267), .Z(n37272) );
  NANDN U37799 ( .A(n37270), .B(n37269), .Z(n37271) );
  AND U37800 ( .A(n37272), .B(n37271), .Z(n37431) );
  NAND U37801 ( .A(n189), .B(n37273), .Z(n37275) );
  XOR U37802 ( .A(a[251]), .B(b[17]), .Z(n37378) );
  NAND U37803 ( .A(n37652), .B(n37378), .Z(n37274) );
  NAND U37804 ( .A(n37275), .B(n37274), .Z(n37360) );
  NAND U37805 ( .A(n188), .B(n37276), .Z(n37278) );
  XOR U37806 ( .A(a[253]), .B(b[15]), .Z(n37381) );
  NAND U37807 ( .A(n37382), .B(n37381), .Z(n37277) );
  NAND U37808 ( .A(n37278), .B(n37277), .Z(n37358) );
  NANDN U37809 ( .A(n174), .B(n37279), .Z(n37281) );
  XOR U37810 ( .A(a[249]), .B(b[19]), .Z(n37363) );
  NANDN U37811 ( .A(n37589), .B(n37363), .Z(n37280) );
  NAND U37812 ( .A(n37281), .B(n37280), .Z(n37420) );
  NAND U37813 ( .A(n38385), .B(n37282), .Z(n37284) );
  XOR U37814 ( .A(b[27]), .B(a[241]), .Z(n37369) );
  NAND U37815 ( .A(n38343), .B(n37369), .Z(n37283) );
  NAND U37816 ( .A(n37284), .B(n37283), .Z(n37419) );
  XOR U37817 ( .A(n37420), .B(n37419), .Z(n37422) );
  NANDN U37818 ( .A(n191), .B(n37285), .Z(n37287) );
  XOR U37819 ( .A(b[25]), .B(a[243]), .Z(n37385) );
  NANDN U37820 ( .A(n37513), .B(n37385), .Z(n37286) );
  NAND U37821 ( .A(n37287), .B(n37286), .Z(n37421) );
  XOR U37822 ( .A(n37422), .B(n37421), .Z(n37357) );
  NAND U37823 ( .A(n194), .B(n37291), .Z(n37293) );
  XOR U37824 ( .A(b[29]), .B(a[239]), .Z(n37372) );
  NAND U37825 ( .A(n38456), .B(n37372), .Z(n37292) );
  NAND U37826 ( .A(n37293), .B(n37292), .Z(n37397) );
  NAND U37827 ( .A(n187), .B(n37294), .Z(n37297) );
  XOR U37828 ( .A(a[255]), .B(b[13]), .Z(n37412) );
  NAND U37829 ( .A(n37295), .B(n37412), .Z(n37296) );
  NAND U37830 ( .A(n37297), .B(n37296), .Z(n37395) );
  NAND U37831 ( .A(n38064), .B(n37298), .Z(n37300) );
  XOR U37832 ( .A(b[21]), .B(a[247]), .Z(n37366) );
  NAND U37833 ( .A(n37993), .B(n37366), .Z(n37299) );
  NAND U37834 ( .A(n37300), .B(n37299), .Z(n37394) );
  AND U37835 ( .A(b[31]), .B(a[235]), .Z(n37391) );
  XNOR U37836 ( .A(n37301), .B(n37391), .Z(n37388) );
  XNOR U37837 ( .A(n37389), .B(n37388), .Z(n37406) );
  NANDN U37838 ( .A(n195), .B(n37302), .Z(n37304) );
  XOR U37839 ( .A(b[31]), .B(a[237]), .Z(n37416) );
  NANDN U37840 ( .A(n38493), .B(n37416), .Z(n37303) );
  AND U37841 ( .A(n37304), .B(n37303), .Z(n37407) );
  XOR U37842 ( .A(n37406), .B(n37407), .Z(n37408) );
  XOR U37843 ( .A(b[23]), .B(a[245]), .Z(n37375) );
  XOR U37844 ( .A(n37400), .B(n37401), .Z(n37402) );
  XOR U37845 ( .A(n37403), .B(n37402), .Z(n37433) );
  XOR U37846 ( .A(n37434), .B(n37433), .Z(n37425) );
  XOR U37847 ( .A(n37426), .B(n37425), .Z(n37427) );
  XOR U37848 ( .A(n37428), .B(n37427), .Z(n37353) );
  XNOR U37849 ( .A(n37354), .B(n37353), .Z(n37348) );
  NAND U37850 ( .A(n37308), .B(n37307), .Z(n37312) );
  NAND U37851 ( .A(n37310), .B(n37309), .Z(n37311) );
  AND U37852 ( .A(n37312), .B(n37311), .Z(n37345) );
  NAND U37853 ( .A(n37314), .B(n37313), .Z(n37318) );
  NAND U37854 ( .A(n37316), .B(n37315), .Z(n37317) );
  AND U37855 ( .A(n37318), .B(n37317), .Z(n37346) );
  XOR U37856 ( .A(n37340), .B(n37339), .Z(n37342) );
  NAND U37857 ( .A(n37320), .B(n37319), .Z(n37324) );
  NAND U37858 ( .A(n37322), .B(n37321), .Z(n37323) );
  AND U37859 ( .A(n37324), .B(n37323), .Z(n37341) );
  XNOR U37860 ( .A(n37342), .B(n37341), .Z(n37334) );
  NAND U37861 ( .A(n37326), .B(n37325), .Z(n37330) );
  NANDN U37862 ( .A(n37328), .B(n37327), .Z(n37329) );
  AND U37863 ( .A(n37330), .B(n37329), .Z(n37333) );
  XOR U37864 ( .A(n37336), .B(n37335), .Z(n37331) );
  XOR U37865 ( .A(n37332), .B(n37331), .Z(c[491]) );
  AND U37866 ( .A(n37332), .B(n37331), .Z(n37438) );
  NAND U37867 ( .A(n37334), .B(n37333), .Z(n37338) );
  NANDN U37868 ( .A(n37336), .B(n37335), .Z(n37337) );
  AND U37869 ( .A(n37338), .B(n37337), .Z(n37442) );
  NAND U37870 ( .A(n37340), .B(n37339), .Z(n37344) );
  NAND U37871 ( .A(n37342), .B(n37341), .Z(n37343) );
  AND U37872 ( .A(n37344), .B(n37343), .Z(n37440) );
  NAND U37873 ( .A(n37346), .B(n37345), .Z(n37350) );
  NAND U37874 ( .A(n37348), .B(n37347), .Z(n37349) );
  AND U37875 ( .A(n37350), .B(n37349), .Z(n37448) );
  NAND U37876 ( .A(n37352), .B(n37351), .Z(n37356) );
  NAND U37877 ( .A(n37354), .B(n37353), .Z(n37355) );
  NAND U37878 ( .A(n37356), .B(n37355), .Z(n37446) );
  NAND U37879 ( .A(n37358), .B(n37357), .Z(n37362) );
  NAND U37880 ( .A(n37360), .B(n37359), .Z(n37361) );
  AND U37881 ( .A(n37362), .B(n37361), .Z(n37460) );
  NAND U37882 ( .A(n190), .B(n37363), .Z(n37365) );
  XOR U37883 ( .A(a[250]), .B(b[19]), .Z(n37484) );
  NAND U37884 ( .A(n37821), .B(n37484), .Z(n37364) );
  NAND U37885 ( .A(n37365), .B(n37364), .Z(n37498) );
  NAND U37886 ( .A(n38064), .B(n37366), .Z(n37368) );
  XOR U37887 ( .A(a[248]), .B(b[21]), .Z(n37487) );
  NAND U37888 ( .A(n37993), .B(n37487), .Z(n37367) );
  NAND U37889 ( .A(n37368), .B(n37367), .Z(n37496) );
  NAND U37890 ( .A(n38385), .B(n37369), .Z(n37371) );
  XOR U37891 ( .A(b[27]), .B(a[242]), .Z(n37478) );
  NAND U37892 ( .A(n38343), .B(n37478), .Z(n37370) );
  NAND U37893 ( .A(n37371), .B(n37370), .Z(n37504) );
  NAND U37894 ( .A(n194), .B(n37372), .Z(n37374) );
  XOR U37895 ( .A(b[29]), .B(a[240]), .Z(n37481) );
  NAND U37896 ( .A(n38456), .B(n37481), .Z(n37373) );
  NAND U37897 ( .A(n37374), .B(n37373), .Z(n37502) );
  NAND U37898 ( .A(n38185), .B(n37375), .Z(n37377) );
  XOR U37899 ( .A(b[23]), .B(a[246]), .Z(n37475) );
  NAND U37900 ( .A(n38132), .B(n37475), .Z(n37376) );
  NAND U37901 ( .A(n37377), .B(n37376), .Z(n37501) );
  NAND U37902 ( .A(n189), .B(n37378), .Z(n37380) );
  XOR U37903 ( .A(a[252]), .B(b[17]), .Z(n37469) );
  NAND U37904 ( .A(n37652), .B(n37469), .Z(n37379) );
  NAND U37905 ( .A(n37380), .B(n37379), .Z(n37492) );
  NAND U37906 ( .A(n188), .B(n37381), .Z(n37384) );
  XOR U37907 ( .A(a[254]), .B(b[15]), .Z(n37508) );
  NAND U37908 ( .A(n37382), .B(n37508), .Z(n37383) );
  NAND U37909 ( .A(n37384), .B(n37383), .Z(n37490) );
  NAND U37910 ( .A(n38289), .B(n37385), .Z(n37387) );
  XOR U37911 ( .A(b[25]), .B(a[244]), .Z(n37512) );
  NAND U37912 ( .A(n38247), .B(n37512), .Z(n37386) );
  NAND U37913 ( .A(n37387), .B(n37386), .Z(n37489) );
  NAND U37914 ( .A(n37389), .B(n37388), .Z(n37393) );
  AND U37915 ( .A(n37391), .B(n37390), .Z(n37392) );
  ANDN U37916 ( .B(n37393), .A(n37392), .Z(n37520) );
  XOR U37917 ( .A(n37519), .B(n37520), .Z(n37522) );
  XOR U37918 ( .A(n37521), .B(n37522), .Z(n37457) );
  NAND U37919 ( .A(n37395), .B(n37394), .Z(n37399) );
  NAND U37920 ( .A(n37397), .B(n37396), .Z(n37398) );
  AND U37921 ( .A(n37399), .B(n37398), .Z(n37458) );
  XOR U37922 ( .A(n37460), .B(n37459), .Z(n37454) );
  NAND U37923 ( .A(n37401), .B(n37400), .Z(n37405) );
  NAND U37924 ( .A(n37403), .B(n37402), .Z(n37404) );
  NAND U37925 ( .A(n37405), .B(n37404), .Z(n37452) );
  NAND U37926 ( .A(n37407), .B(n37406), .Z(n37411) );
  NAND U37927 ( .A(n37409), .B(n37408), .Z(n37410) );
  NAND U37928 ( .A(n37411), .B(n37410), .Z(n37466) );
  AND U37929 ( .A(n37412), .B(n187), .Z(n37415) );
  XOR U37930 ( .A(b[12]), .B(b[11]), .Z(n37413) );
  NAND U37931 ( .A(b[13]), .B(n37413), .Z(n37414) );
  NANDN U37932 ( .A(n37415), .B(n37414), .Z(n37518) );
  AND U37933 ( .A(b[31]), .B(a[236]), .Z(n37551) );
  NAND U37934 ( .A(n38470), .B(n37416), .Z(n37418) );
  XOR U37935 ( .A(b[31]), .B(a[238]), .Z(n37472) );
  NAND U37936 ( .A(n38453), .B(n37472), .Z(n37417) );
  NAND U37937 ( .A(n37418), .B(n37417), .Z(n37516) );
  XNOR U37938 ( .A(n37551), .B(n37516), .Z(n37517) );
  NAND U37939 ( .A(n37420), .B(n37419), .Z(n37424) );
  NAND U37940 ( .A(n37422), .B(n37421), .Z(n37423) );
  AND U37941 ( .A(n37424), .B(n37423), .Z(n37464) );
  XOR U37942 ( .A(n37463), .B(n37464), .Z(n37465) );
  XOR U37943 ( .A(n37454), .B(n37453), .Z(n37528) );
  NAND U37944 ( .A(n37426), .B(n37425), .Z(n37430) );
  NAND U37945 ( .A(n37428), .B(n37427), .Z(n37429) );
  NAND U37946 ( .A(n37430), .B(n37429), .Z(n37526) );
  NAND U37947 ( .A(n37432), .B(n37431), .Z(n37436) );
  NAND U37948 ( .A(n37434), .B(n37433), .Z(n37435) );
  NAND U37949 ( .A(n37436), .B(n37435), .Z(n37525) );
  XOR U37950 ( .A(n37528), .B(n37527), .Z(n37445) );
  XOR U37951 ( .A(n37448), .B(n37447), .Z(n37439) );
  XOR U37952 ( .A(n37440), .B(n37439), .Z(n37441) );
  XOR U37953 ( .A(n37442), .B(n37441), .Z(n37437) );
  XOR U37954 ( .A(n37438), .B(n37437), .Z(c[492]) );
  AND U37955 ( .A(n37438), .B(n37437), .Z(n37532) );
  NAND U37956 ( .A(n37440), .B(n37439), .Z(n37444) );
  NANDN U37957 ( .A(n37442), .B(n37441), .Z(n37443) );
  AND U37958 ( .A(n37444), .B(n37443), .Z(n37536) );
  NAND U37959 ( .A(n37446), .B(n37445), .Z(n37450) );
  NAND U37960 ( .A(n37448), .B(n37447), .Z(n37449) );
  NAND U37961 ( .A(n37450), .B(n37449), .Z(n37534) );
  NAND U37962 ( .A(n37452), .B(n37451), .Z(n37456) );
  NAND U37963 ( .A(n37454), .B(n37453), .Z(n37455) );
  AND U37964 ( .A(n37456), .B(n37455), .Z(n37623) );
  NAND U37965 ( .A(n37458), .B(n37457), .Z(n37462) );
  NAND U37966 ( .A(n37460), .B(n37459), .Z(n37461) );
  AND U37967 ( .A(n37462), .B(n37461), .Z(n37539) );
  NAND U37968 ( .A(n37464), .B(n37463), .Z(n37468) );
  NAND U37969 ( .A(n37466), .B(n37465), .Z(n37467) );
  AND U37970 ( .A(n37468), .B(n37467), .Z(n37540) );
  NAND U37971 ( .A(n189), .B(n37469), .Z(n37471) );
  XOR U37972 ( .A(a[253]), .B(b[17]), .Z(n37585) );
  NAND U37973 ( .A(n37652), .B(n37585), .Z(n37470) );
  NAND U37974 ( .A(n37471), .B(n37470), .Z(n37601) );
  NAND U37975 ( .A(n38470), .B(n37472), .Z(n37474) );
  XOR U37976 ( .A(b[31]), .B(a[239]), .Z(n37561) );
  NAND U37977 ( .A(n38453), .B(n37561), .Z(n37473) );
  NAND U37978 ( .A(n37474), .B(n37473), .Z(n37599) );
  NAND U37979 ( .A(n38185), .B(n37475), .Z(n37477) );
  XOR U37980 ( .A(b[23]), .B(a[247]), .Z(n37582) );
  NAND U37981 ( .A(n38132), .B(n37582), .Z(n37476) );
  NAND U37982 ( .A(n37477), .B(n37476), .Z(n37598) );
  NAND U37983 ( .A(n38385), .B(n37478), .Z(n37480) );
  XOR U37984 ( .A(b[27]), .B(a[243]), .Z(n37570) );
  NAND U37985 ( .A(n38343), .B(n37570), .Z(n37479) );
  NAND U37986 ( .A(n37480), .B(n37479), .Z(n37595) );
  NAND U37987 ( .A(n194), .B(n37481), .Z(n37483) );
  XOR U37988 ( .A(b[29]), .B(a[241]), .Z(n37573) );
  NAND U37989 ( .A(n38456), .B(n37573), .Z(n37482) );
  NAND U37990 ( .A(n37483), .B(n37482), .Z(n37593) );
  NAND U37991 ( .A(n190), .B(n37484), .Z(n37486) );
  XOR U37992 ( .A(a[251]), .B(b[19]), .Z(n37588) );
  NAND U37993 ( .A(n37821), .B(n37588), .Z(n37485) );
  NAND U37994 ( .A(n37486), .B(n37485), .Z(n37592) );
  XOR U37995 ( .A(a[249]), .B(b[21]), .Z(n37579) );
  XOR U37996 ( .A(n37545), .B(n37546), .Z(n37548) );
  XOR U37997 ( .A(n37547), .B(n37548), .Z(n37610) );
  NAND U37998 ( .A(n37490), .B(n37489), .Z(n37494) );
  NAND U37999 ( .A(n37492), .B(n37491), .Z(n37493) );
  AND U38000 ( .A(n37494), .B(n37493), .Z(n37611) );
  NAND U38001 ( .A(n37496), .B(n37495), .Z(n37500) );
  NAND U38002 ( .A(n37498), .B(n37497), .Z(n37499) );
  AND U38003 ( .A(n37500), .B(n37499), .Z(n37612) );
  XNOR U38004 ( .A(n37613), .B(n37612), .Z(n37619) );
  NAND U38005 ( .A(n37502), .B(n37501), .Z(n37506) );
  NAND U38006 ( .A(n37504), .B(n37503), .Z(n37505) );
  AND U38007 ( .A(n37506), .B(n37505), .Z(n37605) );
  AND U38008 ( .A(b[31]), .B(a[237]), .Z(n37553) );
  XNOR U38009 ( .A(n37507), .B(n37553), .Z(n37552) );
  XNOR U38010 ( .A(n37551), .B(n37552), .Z(n37564) );
  NANDN U38011 ( .A(n178), .B(n37508), .Z(n37511) );
  XOR U38012 ( .A(a[255]), .B(b[15]), .Z(n37557) );
  NANDN U38013 ( .A(n37509), .B(n37557), .Z(n37510) );
  AND U38014 ( .A(n37511), .B(n37510), .Z(n37565) );
  XOR U38015 ( .A(n37564), .B(n37565), .Z(n37566) );
  NANDN U38016 ( .A(n191), .B(n37512), .Z(n37515) );
  XOR U38017 ( .A(b[25]), .B(a[245]), .Z(n37576) );
  NANDN U38018 ( .A(n37513), .B(n37576), .Z(n37514) );
  AND U38019 ( .A(n37515), .B(n37514), .Z(n37567) );
  XOR U38020 ( .A(n37605), .B(n37604), .Z(n37607) );
  XNOR U38021 ( .A(n37607), .B(n37606), .Z(n37617) );
  NAND U38022 ( .A(n37520), .B(n37519), .Z(n37524) );
  NAND U38023 ( .A(n37522), .B(n37521), .Z(n37523) );
  AND U38024 ( .A(n37524), .B(n37523), .Z(n37616) );
  XOR U38025 ( .A(n37542), .B(n37541), .Z(n37622) );
  XOR U38026 ( .A(n37623), .B(n37622), .Z(n37625) );
  NAND U38027 ( .A(n37526), .B(n37525), .Z(n37530) );
  NAND U38028 ( .A(n37528), .B(n37527), .Z(n37529) );
  AND U38029 ( .A(n37530), .B(n37529), .Z(n37624) );
  XNOR U38030 ( .A(n37625), .B(n37624), .Z(n37533) );
  XOR U38031 ( .A(n37536), .B(n37535), .Z(n37531) );
  XOR U38032 ( .A(n37532), .B(n37531), .Z(c[493]) );
  AND U38033 ( .A(n37532), .B(n37531), .Z(n37629) );
  NAND U38034 ( .A(n37534), .B(n37533), .Z(n37538) );
  NANDN U38035 ( .A(n37536), .B(n37535), .Z(n37537) );
  AND U38036 ( .A(n37538), .B(n37537), .Z(n37633) );
  NAND U38037 ( .A(n37540), .B(n37539), .Z(n37544) );
  NAND U38038 ( .A(n37542), .B(n37541), .Z(n37543) );
  NAND U38039 ( .A(n37544), .B(n37543), .Z(n37639) );
  NAND U38040 ( .A(n37546), .B(n37545), .Z(n37550) );
  NAND U38041 ( .A(n37548), .B(n37547), .Z(n37549) );
  AND U38042 ( .A(n37550), .B(n37549), .Z(n37708) );
  AND U38043 ( .A(n37552), .B(n37551), .Z(n37556) );
  NAND U38044 ( .A(n37554), .B(n37553), .Z(n37555) );
  NANDN U38045 ( .A(n37556), .B(n37555), .Z(n37696) );
  AND U38046 ( .A(n37557), .B(n188), .Z(n37560) );
  XOR U38047 ( .A(b[14]), .B(b[13]), .Z(n37558) );
  NAND U38048 ( .A(b[15]), .B(n37558), .Z(n37559) );
  NANDN U38049 ( .A(n37560), .B(n37559), .Z(n37678) );
  AND U38050 ( .A(b[31]), .B(a[238]), .Z(n37767) );
  NAND U38051 ( .A(n38470), .B(n37561), .Z(n37563) );
  XOR U38052 ( .A(b[31]), .B(a[240]), .Z(n37679) );
  NAND U38053 ( .A(n38453), .B(n37679), .Z(n37562) );
  NAND U38054 ( .A(n37563), .B(n37562), .Z(n37676) );
  XNOR U38055 ( .A(n37767), .B(n37676), .Z(n37677) );
  NAND U38056 ( .A(n37565), .B(n37564), .Z(n37569) );
  NAND U38057 ( .A(n37567), .B(n37566), .Z(n37568) );
  AND U38058 ( .A(n37569), .B(n37568), .Z(n37698) );
  XOR U38059 ( .A(n37708), .B(n37707), .Z(n37710) );
  NAND U38060 ( .A(n38385), .B(n37570), .Z(n37572) );
  XOR U38061 ( .A(b[27]), .B(a[244]), .Z(n37686) );
  NAND U38062 ( .A(n38343), .B(n37686), .Z(n37571) );
  NAND U38063 ( .A(n37572), .B(n37571), .Z(n37661) );
  NAND U38064 ( .A(n194), .B(n37573), .Z(n37575) );
  XOR U38065 ( .A(b[29]), .B(a[242]), .Z(n37689) );
  NAND U38066 ( .A(n38456), .B(n37689), .Z(n37574) );
  NAND U38067 ( .A(n37575), .B(n37574), .Z(n37659) );
  NAND U38068 ( .A(n38289), .B(n37576), .Z(n37578) );
  XOR U38069 ( .A(b[25]), .B(a[246]), .Z(n37682) );
  NAND U38070 ( .A(n38247), .B(n37682), .Z(n37577) );
  NAND U38071 ( .A(n37578), .B(n37577), .Z(n37658) );
  NAND U38072 ( .A(n38064), .B(n37579), .Z(n37581) );
  XOR U38073 ( .A(a[250]), .B(b[21]), .Z(n37692) );
  NAND U38074 ( .A(n37993), .B(n37692), .Z(n37580) );
  NAND U38075 ( .A(n37581), .B(n37580), .Z(n37667) );
  NAND U38076 ( .A(n38185), .B(n37582), .Z(n37584) );
  XOR U38077 ( .A(b[23]), .B(a[248]), .Z(n37655) );
  NAND U38078 ( .A(n38132), .B(n37655), .Z(n37583) );
  NAND U38079 ( .A(n37584), .B(n37583), .Z(n37665) );
  NAND U38080 ( .A(n189), .B(n37585), .Z(n37587) );
  XOR U38081 ( .A(a[254]), .B(b[17]), .Z(n37651) );
  NAND U38082 ( .A(n37652), .B(n37651), .Z(n37586) );
  NAND U38083 ( .A(n37587), .B(n37586), .Z(n37664) );
  NANDN U38084 ( .A(n174), .B(n37588), .Z(n37591) );
  XOR U38085 ( .A(a[252]), .B(b[19]), .Z(n37648) );
  NANDN U38086 ( .A(n37589), .B(n37648), .Z(n37590) );
  AND U38087 ( .A(n37591), .B(n37590), .Z(n37671) );
  XOR U38088 ( .A(n37670), .B(n37671), .Z(n37673) );
  XNOR U38089 ( .A(n37672), .B(n37673), .Z(n37703) );
  NAND U38090 ( .A(n37593), .B(n37592), .Z(n37597) );
  NAND U38091 ( .A(n37595), .B(n37594), .Z(n37596) );
  NAND U38092 ( .A(n37597), .B(n37596), .Z(n37702) );
  NAND U38093 ( .A(n37599), .B(n37598), .Z(n37603) );
  NAND U38094 ( .A(n37601), .B(n37600), .Z(n37602) );
  NAND U38095 ( .A(n37603), .B(n37602), .Z(n37701) );
  XOR U38096 ( .A(n37703), .B(n37704), .Z(n37709) );
  XNOR U38097 ( .A(n37710), .B(n37709), .Z(n37645) );
  NAND U38098 ( .A(n37605), .B(n37604), .Z(n37609) );
  NAND U38099 ( .A(n37607), .B(n37606), .Z(n37608) );
  NAND U38100 ( .A(n37609), .B(n37608), .Z(n37643) );
  NAND U38101 ( .A(n37611), .B(n37610), .Z(n37615) );
  NAND U38102 ( .A(n37613), .B(n37612), .Z(n37614) );
  NAND U38103 ( .A(n37615), .B(n37614), .Z(n37642) );
  NAND U38104 ( .A(n37617), .B(n37616), .Z(n37621) );
  NAND U38105 ( .A(n37619), .B(n37618), .Z(n37620) );
  NAND U38106 ( .A(n37621), .B(n37620), .Z(n37636) );
  XOR U38107 ( .A(n37637), .B(n37636), .Z(n37638) );
  NAND U38108 ( .A(n37623), .B(n37622), .Z(n37627) );
  NAND U38109 ( .A(n37625), .B(n37624), .Z(n37626) );
  AND U38110 ( .A(n37627), .B(n37626), .Z(n37631) );
  XOR U38111 ( .A(n37630), .B(n37631), .Z(n37632) );
  XOR U38112 ( .A(n37633), .B(n37632), .Z(n37628) );
  XOR U38113 ( .A(n37629), .B(n37628), .Z(c[494]) );
  AND U38114 ( .A(n37629), .B(n37628), .Z(n37714) );
  NAND U38115 ( .A(n37631), .B(n37630), .Z(n37635) );
  NANDN U38116 ( .A(n37633), .B(n37632), .Z(n37634) );
  AND U38117 ( .A(n37635), .B(n37634), .Z(n37718) );
  NAND U38118 ( .A(n37637), .B(n37636), .Z(n37641) );
  NAND U38119 ( .A(n37639), .B(n37638), .Z(n37640) );
  AND U38120 ( .A(n37641), .B(n37640), .Z(n37716) );
  NAND U38121 ( .A(n37643), .B(n37642), .Z(n37647) );
  NAND U38122 ( .A(n37645), .B(n37644), .Z(n37646) );
  NAND U38123 ( .A(n37647), .B(n37646), .Z(n37724) );
  NAND U38124 ( .A(n190), .B(n37648), .Z(n37650) );
  XOR U38125 ( .A(a[253]), .B(b[19]), .Z(n37742) );
  NAND U38126 ( .A(n37821), .B(n37742), .Z(n37649) );
  NAND U38127 ( .A(n37650), .B(n37649), .Z(n37758) );
  NAND U38128 ( .A(n189), .B(n37651), .Z(n37654) );
  XOR U38129 ( .A(a[255]), .B(b[17]), .Z(n37751) );
  NAND U38130 ( .A(n37652), .B(n37751), .Z(n37653) );
  NAND U38131 ( .A(n37654), .B(n37653), .Z(n37756) );
  NAND U38132 ( .A(n38185), .B(n37655), .Z(n37657) );
  XOR U38133 ( .A(b[23]), .B(a[249]), .Z(n37779) );
  NAND U38134 ( .A(n38132), .B(n37779), .Z(n37656) );
  NAND U38135 ( .A(n37657), .B(n37656), .Z(n37755) );
  NAND U38136 ( .A(n37659), .B(n37658), .Z(n37663) );
  NAND U38137 ( .A(n37661), .B(n37660), .Z(n37662) );
  AND U38138 ( .A(n37663), .B(n37662), .Z(n37783) );
  XOR U38139 ( .A(n37782), .B(n37783), .Z(n37785) );
  NAND U38140 ( .A(n37665), .B(n37664), .Z(n37669) );
  NAND U38141 ( .A(n37667), .B(n37666), .Z(n37668) );
  AND U38142 ( .A(n37669), .B(n37668), .Z(n37784) );
  XNOR U38143 ( .A(n37785), .B(n37784), .Z(n37797) );
  NAND U38144 ( .A(n37671), .B(n37670), .Z(n37675) );
  NAND U38145 ( .A(n37673), .B(n37672), .Z(n37674) );
  AND U38146 ( .A(n37675), .B(n37674), .Z(n37795) );
  NAND U38147 ( .A(n38470), .B(n37679), .Z(n37681) );
  XOR U38148 ( .A(b[31]), .B(a[241]), .Z(n37748) );
  NAND U38149 ( .A(n38453), .B(n37748), .Z(n37680) );
  NAND U38150 ( .A(n37681), .B(n37680), .Z(n37734) );
  NAND U38151 ( .A(n38289), .B(n37682), .Z(n37684) );
  XOR U38152 ( .A(b[25]), .B(a[247]), .Z(n37773) );
  NAND U38153 ( .A(n38247), .B(n37773), .Z(n37683) );
  NAND U38154 ( .A(n37684), .B(n37683), .Z(n37733) );
  AND U38155 ( .A(b[31]), .B(a[239]), .Z(n37769) );
  XNOR U38156 ( .A(n37685), .B(n37769), .Z(n37768) );
  XOR U38157 ( .A(n37767), .B(n37768), .Z(n37735) );
  XOR U38158 ( .A(n37736), .B(n37735), .Z(n37789) );
  NAND U38159 ( .A(n38385), .B(n37686), .Z(n37688) );
  XOR U38160 ( .A(b[27]), .B(a[245]), .Z(n37745) );
  NAND U38161 ( .A(n38343), .B(n37745), .Z(n37687) );
  NAND U38162 ( .A(n37688), .B(n37687), .Z(n37764) );
  NAND U38163 ( .A(n194), .B(n37689), .Z(n37691) );
  XOR U38164 ( .A(b[29]), .B(a[243]), .Z(n37776) );
  NAND U38165 ( .A(n38456), .B(n37776), .Z(n37690) );
  NAND U38166 ( .A(n37691), .B(n37690), .Z(n37762) );
  NAND U38167 ( .A(n38064), .B(n37692), .Z(n37694) );
  XOR U38168 ( .A(a[251]), .B(b[21]), .Z(n37739) );
  NAND U38169 ( .A(n37993), .B(n37739), .Z(n37693) );
  NAND U38170 ( .A(n37694), .B(n37693), .Z(n37761) );
  XOR U38171 ( .A(n37789), .B(n37788), .Z(n37790) );
  XOR U38172 ( .A(n37795), .B(n37794), .Z(n37796) );
  NAND U38173 ( .A(n37696), .B(n37695), .Z(n37700) );
  NAND U38174 ( .A(n37698), .B(n37697), .Z(n37699) );
  AND U38175 ( .A(n37700), .B(n37699), .Z(n37727) );
  NAND U38176 ( .A(n37702), .B(n37701), .Z(n37706) );
  NAND U38177 ( .A(n37704), .B(n37703), .Z(n37705) );
  AND U38178 ( .A(n37706), .B(n37705), .Z(n37728) );
  XOR U38179 ( .A(n37729), .B(n37730), .Z(n37721) );
  NAND U38180 ( .A(n37708), .B(n37707), .Z(n37712) );
  NAND U38181 ( .A(n37710), .B(n37709), .Z(n37711) );
  AND U38182 ( .A(n37712), .B(n37711), .Z(n37722) );
  XOR U38183 ( .A(n37716), .B(n37715), .Z(n37717) );
  XOR U38184 ( .A(n37718), .B(n37717), .Z(n37713) );
  XOR U38185 ( .A(n37714), .B(n37713), .Z(c[495]) );
  AND U38186 ( .A(n37714), .B(n37713), .Z(n37801) );
  NAND U38187 ( .A(n37716), .B(n37715), .Z(n37720) );
  NANDN U38188 ( .A(n37718), .B(n37717), .Z(n37719) );
  AND U38189 ( .A(n37720), .B(n37719), .Z(n37805) );
  NAND U38190 ( .A(n37722), .B(n37721), .Z(n37726) );
  NAND U38191 ( .A(n37724), .B(n37723), .Z(n37725) );
  NAND U38192 ( .A(n37726), .B(n37725), .Z(n37803) );
  NAND U38193 ( .A(n37728), .B(n37727), .Z(n37732) );
  NAND U38194 ( .A(n37730), .B(n37729), .Z(n37731) );
  NAND U38195 ( .A(n37732), .B(n37731), .Z(n37811) );
  NAND U38196 ( .A(n37734), .B(n37733), .Z(n37738) );
  NAND U38197 ( .A(n37736), .B(n37735), .Z(n37737) );
  NAND U38198 ( .A(n37738), .B(n37737), .Z(n37873) );
  NAND U38199 ( .A(n38064), .B(n37739), .Z(n37741) );
  XOR U38200 ( .A(a[252]), .B(b[21]), .Z(n37833) );
  NAND U38201 ( .A(n37993), .B(n37833), .Z(n37740) );
  NAND U38202 ( .A(n37741), .B(n37740), .Z(n37863) );
  NAND U38203 ( .A(n190), .B(n37742), .Z(n37744) );
  XOR U38204 ( .A(a[254]), .B(b[19]), .Z(n37820) );
  NAND U38205 ( .A(n37821), .B(n37820), .Z(n37743) );
  NAND U38206 ( .A(n37744), .B(n37743), .Z(n37861) );
  NAND U38207 ( .A(n38385), .B(n37745), .Z(n37747) );
  XOR U38208 ( .A(b[27]), .B(a[246]), .Z(n37824) );
  NAND U38209 ( .A(n38343), .B(n37824), .Z(n37746) );
  NAND U38210 ( .A(n37747), .B(n37746), .Z(n37860) );
  NAND U38211 ( .A(n38470), .B(n37748), .Z(n37750) );
  XOR U38212 ( .A(b[31]), .B(a[242]), .Z(n37836) );
  NAND U38213 ( .A(n38453), .B(n37836), .Z(n37749) );
  AND U38214 ( .A(n37750), .B(n37749), .Z(n37869) );
  AND U38215 ( .A(b[31]), .B(a[240]), .Z(n37938) );
  AND U38216 ( .A(n37751), .B(n189), .Z(n37754) );
  XOR U38217 ( .A(b[16]), .B(b[15]), .Z(n37752) );
  NAND U38218 ( .A(b[17]), .B(n37752), .Z(n37753) );
  NANDN U38219 ( .A(n37754), .B(n37753), .Z(n37866) );
  XNOR U38220 ( .A(n37938), .B(n37866), .Z(n37868) );
  XOR U38221 ( .A(n37869), .B(n37868), .Z(n37848) );
  XOR U38222 ( .A(n37849), .B(n37848), .Z(n37851) );
  NAND U38223 ( .A(n37756), .B(n37755), .Z(n37760) );
  NAND U38224 ( .A(n37758), .B(n37757), .Z(n37759) );
  AND U38225 ( .A(n37760), .B(n37759), .Z(n37850) );
  XNOR U38226 ( .A(n37851), .B(n37850), .Z(n37872) );
  NAND U38227 ( .A(n37762), .B(n37761), .Z(n37766) );
  NAND U38228 ( .A(n37764), .B(n37763), .Z(n37765) );
  NAND U38229 ( .A(n37766), .B(n37765), .Z(n37857) );
  AND U38230 ( .A(n37768), .B(n37767), .Z(n37772) );
  NAND U38231 ( .A(n37770), .B(n37769), .Z(n37771) );
  NANDN U38232 ( .A(n37772), .B(n37771), .Z(n37855) );
  NAND U38233 ( .A(n38289), .B(n37773), .Z(n37775) );
  XOR U38234 ( .A(b[25]), .B(a[248]), .Z(n37839) );
  NAND U38235 ( .A(n38247), .B(n37839), .Z(n37774) );
  NAND U38236 ( .A(n37775), .B(n37774), .Z(n37845) );
  NAND U38237 ( .A(n194), .B(n37776), .Z(n37778) );
  XOR U38238 ( .A(b[29]), .B(a[244]), .Z(n37827) );
  NAND U38239 ( .A(n38456), .B(n37827), .Z(n37777) );
  NAND U38240 ( .A(n37778), .B(n37777), .Z(n37843) );
  NAND U38241 ( .A(n38185), .B(n37779), .Z(n37781) );
  XOR U38242 ( .A(a[250]), .B(b[23]), .Z(n37830) );
  NAND U38243 ( .A(n38132), .B(n37830), .Z(n37780) );
  NAND U38244 ( .A(n37781), .B(n37780), .Z(n37842) );
  XNOR U38245 ( .A(n37875), .B(n37874), .Z(n37817) );
  NAND U38246 ( .A(n37783), .B(n37782), .Z(n37787) );
  NAND U38247 ( .A(n37785), .B(n37784), .Z(n37786) );
  NAND U38248 ( .A(n37787), .B(n37786), .Z(n37815) );
  NAND U38249 ( .A(n37789), .B(n37788), .Z(n37793) );
  NAND U38250 ( .A(n37791), .B(n37790), .Z(n37792) );
  AND U38251 ( .A(n37793), .B(n37792), .Z(n37814) );
  NAND U38252 ( .A(n37795), .B(n37794), .Z(n37799) );
  NAND U38253 ( .A(n37797), .B(n37796), .Z(n37798) );
  AND U38254 ( .A(n37799), .B(n37798), .Z(n37809) );
  XOR U38255 ( .A(n37805), .B(n37804), .Z(n37800) );
  XOR U38256 ( .A(n37801), .B(n37800), .Z(c[496]) );
  AND U38257 ( .A(n37801), .B(n37800), .Z(n37879) );
  NAND U38258 ( .A(n37803), .B(n37802), .Z(n37807) );
  NANDN U38259 ( .A(n37805), .B(n37804), .Z(n37806) );
  AND U38260 ( .A(n37807), .B(n37806), .Z(n37883) );
  NAND U38261 ( .A(n37809), .B(n37808), .Z(n37813) );
  NAND U38262 ( .A(n37811), .B(n37810), .Z(n37812) );
  NAND U38263 ( .A(n37813), .B(n37812), .Z(n37881) );
  NAND U38264 ( .A(n37815), .B(n37814), .Z(n37819) );
  NAND U38265 ( .A(n37817), .B(n37816), .Z(n37818) );
  NAND U38266 ( .A(n37819), .B(n37818), .Z(n37889) );
  NAND U38267 ( .A(n190), .B(n37820), .Z(n37823) );
  XOR U38268 ( .A(a[255]), .B(b[19]), .Z(n37947) );
  NAND U38269 ( .A(n37821), .B(n37947), .Z(n37822) );
  NAND U38270 ( .A(n37823), .B(n37822), .Z(n37933) );
  NAND U38271 ( .A(n38385), .B(n37824), .Z(n37826) );
  XOR U38272 ( .A(b[27]), .B(a[247]), .Z(n37928) );
  NAND U38273 ( .A(n38343), .B(n37928), .Z(n37825) );
  NAND U38274 ( .A(n37826), .B(n37825), .Z(n37932) );
  IV U38275 ( .A(n37938), .Z(n37867) );
  AND U38276 ( .A(b[31]), .B(a[241]), .Z(n37941) );
  XOR U38277 ( .A(n37940), .B(n37941), .Z(n37939) );
  XNOR U38278 ( .A(n37867), .B(n37939), .Z(n37934) );
  XNOR U38279 ( .A(n37935), .B(n37934), .Z(n37905) );
  NAND U38280 ( .A(n194), .B(n37827), .Z(n37829) );
  XOR U38281 ( .A(b[29]), .B(a[245]), .Z(n37925) );
  NAND U38282 ( .A(n38456), .B(n37925), .Z(n37828) );
  AND U38283 ( .A(n37829), .B(n37828), .Z(n37954) );
  NAND U38284 ( .A(n38185), .B(n37830), .Z(n37832) );
  XOR U38285 ( .A(a[251]), .B(b[23]), .Z(n37916) );
  NAND U38286 ( .A(n38132), .B(n37916), .Z(n37831) );
  NAND U38287 ( .A(n37832), .B(n37831), .Z(n37952) );
  NAND U38288 ( .A(n38064), .B(n37833), .Z(n37835) );
  XOR U38289 ( .A(a[253]), .B(b[21]), .Z(n37919) );
  NAND U38290 ( .A(n37993), .B(n37919), .Z(n37834) );
  NAND U38291 ( .A(n37835), .B(n37834), .Z(n37913) );
  NAND U38292 ( .A(n38470), .B(n37836), .Z(n37838) );
  XOR U38293 ( .A(b[31]), .B(a[243]), .Z(n37944) );
  NAND U38294 ( .A(n38453), .B(n37944), .Z(n37837) );
  NAND U38295 ( .A(n37838), .B(n37837), .Z(n37911) );
  NAND U38296 ( .A(n38289), .B(n37839), .Z(n37841) );
  XOR U38297 ( .A(b[25]), .B(a[249]), .Z(n37922) );
  NAND U38298 ( .A(n38247), .B(n37922), .Z(n37840) );
  NAND U38299 ( .A(n37841), .B(n37840), .Z(n37910) );
  XOR U38300 ( .A(n37954), .B(n37953), .Z(n37904) );
  NAND U38301 ( .A(n37843), .B(n37842), .Z(n37847) );
  NAND U38302 ( .A(n37845), .B(n37844), .Z(n37846) );
  AND U38303 ( .A(n37847), .B(n37846), .Z(n37906) );
  XNOR U38304 ( .A(n37907), .B(n37906), .Z(n37893) );
  NAND U38305 ( .A(n37849), .B(n37848), .Z(n37853) );
  NAND U38306 ( .A(n37851), .B(n37850), .Z(n37852) );
  AND U38307 ( .A(n37853), .B(n37852), .Z(n37892) );
  NAND U38308 ( .A(n37855), .B(n37854), .Z(n37859) );
  NAND U38309 ( .A(n37857), .B(n37856), .Z(n37858) );
  NAND U38310 ( .A(n37859), .B(n37858), .Z(n37901) );
  NAND U38311 ( .A(n37861), .B(n37860), .Z(n37865) );
  NAND U38312 ( .A(n37863), .B(n37862), .Z(n37864) );
  NAND U38313 ( .A(n37865), .B(n37864), .Z(n37899) );
  NAND U38314 ( .A(n37867), .B(n37866), .Z(n37871) );
  NANDN U38315 ( .A(n37869), .B(n37868), .Z(n37870) );
  NAND U38316 ( .A(n37871), .B(n37870), .Z(n37898) );
  XNOR U38317 ( .A(n37895), .B(n37894), .Z(n37887) );
  NAND U38318 ( .A(n37873), .B(n37872), .Z(n37877) );
  NAND U38319 ( .A(n37875), .B(n37874), .Z(n37876) );
  AND U38320 ( .A(n37877), .B(n37876), .Z(n37886) );
  XOR U38321 ( .A(n37883), .B(n37882), .Z(n37878) );
  XOR U38322 ( .A(n37879), .B(n37878), .Z(c[497]) );
  AND U38323 ( .A(n37879), .B(n37878), .Z(n37958) );
  NAND U38324 ( .A(n37881), .B(n37880), .Z(n37885) );
  NANDN U38325 ( .A(n37883), .B(n37882), .Z(n37884) );
  AND U38326 ( .A(n37885), .B(n37884), .Z(n37962) );
  NAND U38327 ( .A(n37887), .B(n37886), .Z(n37891) );
  NAND U38328 ( .A(n37889), .B(n37888), .Z(n37890) );
  NAND U38329 ( .A(n37891), .B(n37890), .Z(n37960) );
  NAND U38330 ( .A(n37893), .B(n37892), .Z(n37897) );
  NAND U38331 ( .A(n37895), .B(n37894), .Z(n37896) );
  AND U38332 ( .A(n37897), .B(n37896), .Z(n37968) );
  NAND U38333 ( .A(n37899), .B(n37898), .Z(n37903) );
  NAND U38334 ( .A(n37901), .B(n37900), .Z(n37902) );
  AND U38335 ( .A(n37903), .B(n37902), .Z(n37966) );
  NAND U38336 ( .A(n37905), .B(n37904), .Z(n37909) );
  NAND U38337 ( .A(n37907), .B(n37906), .Z(n37908) );
  NAND U38338 ( .A(n37909), .B(n37908), .Z(n38020) );
  NAND U38339 ( .A(n37911), .B(n37910), .Z(n37915) );
  NAND U38340 ( .A(n37913), .B(n37912), .Z(n37914) );
  NAND U38341 ( .A(n37915), .B(n37914), .Z(n38012) );
  NAND U38342 ( .A(n38185), .B(n37916), .Z(n37918) );
  XOR U38343 ( .A(a[252]), .B(b[23]), .Z(n37986) );
  NAND U38344 ( .A(n38132), .B(n37986), .Z(n37917) );
  NAND U38345 ( .A(n37918), .B(n37917), .Z(n38002) );
  NAND U38346 ( .A(n38064), .B(n37919), .Z(n37921) );
  XOR U38347 ( .A(a[254]), .B(b[21]), .Z(n37992) );
  NAND U38348 ( .A(n37993), .B(n37992), .Z(n37920) );
  NAND U38349 ( .A(n37921), .B(n37920), .Z(n38000) );
  NAND U38350 ( .A(n38289), .B(n37922), .Z(n37924) );
  XOR U38351 ( .A(b[25]), .B(a[250]), .Z(n37983) );
  NAND U38352 ( .A(n38247), .B(n37983), .Z(n37923) );
  NAND U38353 ( .A(n37924), .B(n37923), .Z(n37974) );
  IV U38354 ( .A(n37974), .Z(n37931) );
  NAND U38355 ( .A(n194), .B(n37925), .Z(n37927) );
  XOR U38356 ( .A(b[29]), .B(a[246]), .Z(n37980) );
  NAND U38357 ( .A(n38456), .B(n37980), .Z(n37926) );
  NAND U38358 ( .A(n37927), .B(n37926), .Z(n37972) );
  NAND U38359 ( .A(n38385), .B(n37928), .Z(n37930) );
  XOR U38360 ( .A(b[27]), .B(a[248]), .Z(n37996) );
  NAND U38361 ( .A(n38343), .B(n37996), .Z(n37929) );
  NAND U38362 ( .A(n37930), .B(n37929), .Z(n37971) );
  XNOR U38363 ( .A(n37931), .B(n37973), .Z(n37999) );
  NAND U38364 ( .A(n37933), .B(n37932), .Z(n37937) );
  NAND U38365 ( .A(n37935), .B(n37934), .Z(n37936) );
  NAND U38366 ( .A(n37937), .B(n37936), .Z(n38008) );
  AND U38367 ( .A(n37939), .B(n37938), .Z(n37943) );
  NAND U38368 ( .A(n37941), .B(n37940), .Z(n37942) );
  NANDN U38369 ( .A(n37943), .B(n37942), .Z(n38006) );
  NAND U38370 ( .A(n38470), .B(n37944), .Z(n37946) );
  XOR U38371 ( .A(b[31]), .B(a[244]), .Z(n37989) );
  NAND U38372 ( .A(n38453), .B(n37989), .Z(n37945) );
  NAND U38373 ( .A(n37946), .B(n37945), .Z(n37979) );
  AND U38374 ( .A(b[31]), .B(a[242]), .Z(n38044) );
  AND U38375 ( .A(n37947), .B(n190), .Z(n37950) );
  XOR U38376 ( .A(b[18]), .B(b[17]), .Z(n37948) );
  NAND U38377 ( .A(b[19]), .B(n37948), .Z(n37949) );
  NANDN U38378 ( .A(n37950), .B(n37949), .Z(n37977) );
  XNOR U38379 ( .A(n38044), .B(n37977), .Z(n37978) );
  XNOR U38380 ( .A(n38014), .B(n38013), .Z(n38018) );
  NAND U38381 ( .A(n37952), .B(n37951), .Z(n37956) );
  NANDN U38382 ( .A(n37954), .B(n37953), .Z(n37955) );
  AND U38383 ( .A(n37956), .B(n37955), .Z(n38017) );
  XOR U38384 ( .A(n37966), .B(n37965), .Z(n37967) );
  XOR U38385 ( .A(n37968), .B(n37967), .Z(n37959) );
  XOR U38386 ( .A(n37962), .B(n37961), .Z(n37957) );
  XOR U38387 ( .A(n37958), .B(n37957), .Z(c[498]) );
  AND U38388 ( .A(n37958), .B(n37957), .Z(n38024) );
  NAND U38389 ( .A(n37960), .B(n37959), .Z(n37964) );
  NANDN U38390 ( .A(n37962), .B(n37961), .Z(n37963) );
  AND U38391 ( .A(n37964), .B(n37963), .Z(n38028) );
  NAND U38392 ( .A(n37966), .B(n37965), .Z(n37970) );
  NAND U38393 ( .A(n37968), .B(n37967), .Z(n37969) );
  NAND U38394 ( .A(n37970), .B(n37969), .Z(n38026) );
  NAND U38395 ( .A(n37972), .B(n37971), .Z(n37976) );
  NAND U38396 ( .A(n37974), .B(n37973), .Z(n37975) );
  NAND U38397 ( .A(n37976), .B(n37975), .Z(n38088) );
  NAND U38398 ( .A(n194), .B(n37980), .Z(n37982) );
  XOR U38399 ( .A(b[29]), .B(a[247]), .Z(n38078) );
  NAND U38400 ( .A(n38456), .B(n38078), .Z(n37981) );
  NAND U38401 ( .A(n37982), .B(n37981), .Z(n38082) );
  NAND U38402 ( .A(n38289), .B(n37983), .Z(n37985) );
  XOR U38403 ( .A(b[25]), .B(a[251]), .Z(n38069) );
  NAND U38404 ( .A(n38247), .B(n38069), .Z(n37984) );
  NAND U38405 ( .A(n37985), .B(n37984), .Z(n38058) );
  NAND U38406 ( .A(n38185), .B(n37986), .Z(n37988) );
  XOR U38407 ( .A(a[253]), .B(b[23]), .Z(n38072) );
  NAND U38408 ( .A(n38132), .B(n38072), .Z(n37987) );
  NAND U38409 ( .A(n37988), .B(n37987), .Z(n38056) );
  NAND U38410 ( .A(n38470), .B(n37989), .Z(n37991) );
  XOR U38411 ( .A(b[31]), .B(a[245]), .Z(n38061) );
  NAND U38412 ( .A(n38453), .B(n38061), .Z(n37990) );
  NAND U38413 ( .A(n37991), .B(n37990), .Z(n38055) );
  NAND U38414 ( .A(n38064), .B(n37992), .Z(n37995) );
  XOR U38415 ( .A(a[255]), .B(b[21]), .Z(n38065) );
  NAND U38416 ( .A(n37993), .B(n38065), .Z(n37994) );
  NAND U38417 ( .A(n37995), .B(n37994), .Z(n38050) );
  NAND U38418 ( .A(n38385), .B(n37996), .Z(n37998) );
  XOR U38419 ( .A(b[27]), .B(a[249]), .Z(n38075) );
  NAND U38420 ( .A(n38343), .B(n38075), .Z(n37997) );
  NAND U38421 ( .A(n37998), .B(n37997), .Z(n38049) );
  AND U38422 ( .A(b[31]), .B(a[243]), .Z(n38046) );
  XOR U38423 ( .A(n38045), .B(n38046), .Z(n38043) );
  XOR U38424 ( .A(n38044), .B(n38043), .Z(n38051) );
  XOR U38425 ( .A(n38052), .B(n38051), .Z(n38083) );
  XOR U38426 ( .A(n38084), .B(n38083), .Z(n38089) );
  XNOR U38427 ( .A(n38090), .B(n38089), .Z(n38040) );
  NAND U38428 ( .A(n38000), .B(n37999), .Z(n38004) );
  NAND U38429 ( .A(n38002), .B(n38001), .Z(n38003) );
  AND U38430 ( .A(n38004), .B(n38003), .Z(n38037) );
  NAND U38431 ( .A(n38006), .B(n38005), .Z(n38010) );
  NAND U38432 ( .A(n38008), .B(n38007), .Z(n38009) );
  AND U38433 ( .A(n38010), .B(n38009), .Z(n38038) );
  NAND U38434 ( .A(n38012), .B(n38011), .Z(n38016) );
  NAND U38435 ( .A(n38014), .B(n38013), .Z(n38015) );
  NAND U38436 ( .A(n38016), .B(n38015), .Z(n38031) );
  XOR U38437 ( .A(n38032), .B(n38031), .Z(n38034) );
  NAND U38438 ( .A(n38018), .B(n38017), .Z(n38022) );
  NAND U38439 ( .A(n38020), .B(n38019), .Z(n38021) );
  AND U38440 ( .A(n38022), .B(n38021), .Z(n38033) );
  XNOR U38441 ( .A(n38034), .B(n38033), .Z(n38025) );
  XOR U38442 ( .A(n38028), .B(n38027), .Z(n38023) );
  XOR U38443 ( .A(n38024), .B(n38023), .Z(c[499]) );
  AND U38444 ( .A(n38024), .B(n38023), .Z(n38094) );
  NAND U38445 ( .A(n38026), .B(n38025), .Z(n38030) );
  NANDN U38446 ( .A(n38028), .B(n38027), .Z(n38029) );
  AND U38447 ( .A(n38030), .B(n38029), .Z(n38098) );
  NAND U38448 ( .A(n38032), .B(n38031), .Z(n38036) );
  NAND U38449 ( .A(n38034), .B(n38033), .Z(n38035) );
  AND U38450 ( .A(n38036), .B(n38035), .Z(n38096) );
  NAND U38451 ( .A(n38038), .B(n38037), .Z(n38042) );
  NAND U38452 ( .A(n38040), .B(n38039), .Z(n38041) );
  NAND U38453 ( .A(n38042), .B(n38041), .Z(n38104) );
  NAND U38454 ( .A(n38044), .B(n38043), .Z(n38048) );
  AND U38455 ( .A(n38046), .B(n38045), .Z(n38047) );
  ANDN U38456 ( .B(n38048), .A(n38047), .Z(n38113) );
  NAND U38457 ( .A(n38050), .B(n38049), .Z(n38054) );
  NAND U38458 ( .A(n38052), .B(n38051), .Z(n38053) );
  AND U38459 ( .A(n38054), .B(n38053), .Z(n38114) );
  NAND U38460 ( .A(n38056), .B(n38055), .Z(n38060) );
  NAND U38461 ( .A(n38058), .B(n38057), .Z(n38059) );
  AND U38462 ( .A(n38060), .B(n38059), .Z(n38115) );
  XNOR U38463 ( .A(n38116), .B(n38115), .Z(n38110) );
  NAND U38464 ( .A(n38470), .B(n38061), .Z(n38063) );
  XOR U38465 ( .A(b[31]), .B(a[246]), .Z(n38144) );
  NAND U38466 ( .A(n38453), .B(n38144), .Z(n38062) );
  NAND U38467 ( .A(n38063), .B(n38062), .Z(n38150) );
  AND U38468 ( .A(b[31]), .B(a[244]), .Z(n38203) );
  AND U38469 ( .A(n38065), .B(n38064), .Z(n38068) );
  XOR U38470 ( .A(b[20]), .B(b[19]), .Z(n38066) );
  NAND U38471 ( .A(b[21]), .B(n38066), .Z(n38067) );
  NANDN U38472 ( .A(n38068), .B(n38067), .Z(n38147) );
  XNOR U38473 ( .A(n38203), .B(n38147), .Z(n38149) );
  NAND U38474 ( .A(n38289), .B(n38069), .Z(n38071) );
  XOR U38475 ( .A(a[252]), .B(b[25]), .Z(n38138) );
  NAND U38476 ( .A(n38247), .B(n38138), .Z(n38070) );
  NAND U38477 ( .A(n38071), .B(n38070), .Z(n38128) );
  NAND U38478 ( .A(n38185), .B(n38072), .Z(n38074) );
  XOR U38479 ( .A(a[254]), .B(b[23]), .Z(n38131) );
  NAND U38480 ( .A(n38132), .B(n38131), .Z(n38073) );
  NAND U38481 ( .A(n38074), .B(n38073), .Z(n38126) );
  NAND U38482 ( .A(n38385), .B(n38075), .Z(n38077) );
  XOR U38483 ( .A(b[27]), .B(a[250]), .Z(n38135) );
  NAND U38484 ( .A(n38343), .B(n38135), .Z(n38076) );
  NAND U38485 ( .A(n38077), .B(n38076), .Z(n38125) );
  NANDN U38486 ( .A(n177), .B(n38078), .Z(n38080) );
  XOR U38487 ( .A(b[29]), .B(a[248]), .Z(n38141) );
  NANDN U38488 ( .A(n193), .B(n38141), .Z(n38079) );
  AND U38489 ( .A(n38080), .B(n38079), .Z(n38120) );
  XOR U38490 ( .A(n38119), .B(n38120), .Z(n38122) );
  XNOR U38491 ( .A(n38121), .B(n38122), .Z(n38108) );
  NAND U38492 ( .A(n38082), .B(n38081), .Z(n38086) );
  NAND U38493 ( .A(n38084), .B(n38083), .Z(n38085) );
  NAND U38494 ( .A(n38086), .B(n38085), .Z(n38107) );
  XOR U38495 ( .A(n38108), .B(n38107), .Z(n38109) );
  NAND U38496 ( .A(n38088), .B(n38087), .Z(n38092) );
  NAND U38497 ( .A(n38090), .B(n38089), .Z(n38091) );
  AND U38498 ( .A(n38092), .B(n38091), .Z(n38102) );
  XOR U38499 ( .A(n38101), .B(n38102), .Z(n38103) );
  XOR U38500 ( .A(n38096), .B(n38095), .Z(n38097) );
  XOR U38501 ( .A(n38098), .B(n38097), .Z(n38093) );
  XOR U38502 ( .A(n38094), .B(n38093), .Z(c[500]) );
  AND U38503 ( .A(n38094), .B(n38093), .Z(n38154) );
  NAND U38504 ( .A(n38096), .B(n38095), .Z(n38100) );
  NANDN U38505 ( .A(n38098), .B(n38097), .Z(n38099) );
  AND U38506 ( .A(n38100), .B(n38099), .Z(n38158) );
  NAND U38507 ( .A(n38102), .B(n38101), .Z(n38106) );
  NAND U38508 ( .A(n38104), .B(n38103), .Z(n38105) );
  NAND U38509 ( .A(n38106), .B(n38105), .Z(n38156) );
  NAND U38510 ( .A(n38108), .B(n38107), .Z(n38112) );
  NAND U38511 ( .A(n38110), .B(n38109), .Z(n38111) );
  AND U38512 ( .A(n38112), .B(n38111), .Z(n38164) );
  NAND U38513 ( .A(n38114), .B(n38113), .Z(n38118) );
  NAND U38514 ( .A(n38116), .B(n38115), .Z(n38117) );
  NAND U38515 ( .A(n38118), .B(n38117), .Z(n38162) );
  NAND U38516 ( .A(n38120), .B(n38119), .Z(n38124) );
  NAND U38517 ( .A(n38122), .B(n38121), .Z(n38123) );
  NAND U38518 ( .A(n38124), .B(n38123), .Z(n38170) );
  NAND U38519 ( .A(n38126), .B(n38125), .Z(n38130) );
  NAND U38520 ( .A(n38128), .B(n38127), .Z(n38129) );
  NAND U38521 ( .A(n38130), .B(n38129), .Z(n38211) );
  NAND U38522 ( .A(n38185), .B(n38131), .Z(n38134) );
  XOR U38523 ( .A(a[255]), .B(b[23]), .Z(n38186) );
  NAND U38524 ( .A(n38132), .B(n38186), .Z(n38133) );
  NAND U38525 ( .A(n38134), .B(n38133), .Z(n38197) );
  NAND U38526 ( .A(n38385), .B(n38135), .Z(n38137) );
  XOR U38527 ( .A(b[27]), .B(a[251]), .Z(n38173) );
  NAND U38528 ( .A(n38343), .B(n38173), .Z(n38136) );
  NAND U38529 ( .A(n38137), .B(n38136), .Z(n38196) );
  IV U38530 ( .A(n38203), .Z(n38148) );
  XNOR U38531 ( .A(n38148), .B(n38202), .Z(n38205) );
  AND U38532 ( .A(b[31]), .B(a[245]), .Z(n38204) );
  XOR U38533 ( .A(n38205), .B(n38204), .Z(n38198) );
  XOR U38534 ( .A(n38199), .B(n38198), .Z(n38209) );
  NAND U38535 ( .A(n38289), .B(n38138), .Z(n38140) );
  XOR U38536 ( .A(a[253]), .B(b[25]), .Z(n38176) );
  NAND U38537 ( .A(n38247), .B(n38176), .Z(n38139) );
  NAND U38538 ( .A(n38140), .B(n38139), .Z(n38193) );
  NAND U38539 ( .A(n194), .B(n38141), .Z(n38143) );
  XOR U38540 ( .A(b[29]), .B(a[249]), .Z(n38179) );
  NAND U38541 ( .A(n38456), .B(n38179), .Z(n38142) );
  NAND U38542 ( .A(n38143), .B(n38142), .Z(n38191) );
  NAND U38543 ( .A(n38470), .B(n38144), .Z(n38146) );
  XOR U38544 ( .A(b[31]), .B(a[247]), .Z(n38182) );
  NAND U38545 ( .A(n38453), .B(n38182), .Z(n38145) );
  NAND U38546 ( .A(n38146), .B(n38145), .Z(n38190) );
  XOR U38547 ( .A(n38209), .B(n38208), .Z(n38210) );
  NAND U38548 ( .A(n38148), .B(n38147), .Z(n38152) );
  NAND U38549 ( .A(n38150), .B(n38149), .Z(n38151) );
  AND U38550 ( .A(n38152), .B(n38151), .Z(n38168) );
  XOR U38551 ( .A(n38167), .B(n38168), .Z(n38169) );
  XOR U38552 ( .A(n38164), .B(n38163), .Z(n38155) );
  XOR U38553 ( .A(n38158), .B(n38157), .Z(n38153) );
  XOR U38554 ( .A(n38154), .B(n38153), .Z(c[501]) );
  AND U38555 ( .A(n38154), .B(n38153), .Z(n38215) );
  NAND U38556 ( .A(n38156), .B(n38155), .Z(n38160) );
  NANDN U38557 ( .A(n38158), .B(n38157), .Z(n38159) );
  AND U38558 ( .A(n38160), .B(n38159), .Z(n38219) );
  NAND U38559 ( .A(n38162), .B(n38161), .Z(n38166) );
  NAND U38560 ( .A(n38164), .B(n38163), .Z(n38165) );
  NAND U38561 ( .A(n38166), .B(n38165), .Z(n38217) );
  NAND U38562 ( .A(n38168), .B(n38167), .Z(n38172) );
  NAND U38563 ( .A(n38170), .B(n38169), .Z(n38171) );
  NAND U38564 ( .A(n38172), .B(n38171), .Z(n38225) );
  NAND U38565 ( .A(n38385), .B(n38173), .Z(n38175) );
  XOR U38566 ( .A(b[27]), .B(a[252]), .Z(n38243) );
  NAND U38567 ( .A(n38343), .B(n38243), .Z(n38174) );
  NAND U38568 ( .A(n38175), .B(n38174), .Z(n38234) );
  NAND U38569 ( .A(n38289), .B(n38176), .Z(n38178) );
  XOR U38570 ( .A(a[254]), .B(b[25]), .Z(n38246) );
  NAND U38571 ( .A(n38247), .B(n38246), .Z(n38177) );
  NAND U38572 ( .A(n38178), .B(n38177), .Z(n38232) );
  NAND U38573 ( .A(n194), .B(n38179), .Z(n38181) );
  XOR U38574 ( .A(b[29]), .B(a[250]), .Z(n38250) );
  NAND U38575 ( .A(n38456), .B(n38250), .Z(n38180) );
  NAND U38576 ( .A(n38181), .B(n38180), .Z(n38231) );
  NAND U38577 ( .A(n38470), .B(n38182), .Z(n38184) );
  XOR U38578 ( .A(b[31]), .B(a[248]), .Z(n38240) );
  NAND U38579 ( .A(n38453), .B(n38240), .Z(n38183) );
  AND U38580 ( .A(n38184), .B(n38183), .Z(n38239) );
  AND U38581 ( .A(b[31]), .B(a[246]), .Z(n38295) );
  AND U38582 ( .A(n38186), .B(n38185), .Z(n38189) );
  XOR U38583 ( .A(b[22]), .B(b[21]), .Z(n38187) );
  NAND U38584 ( .A(b[23]), .B(n38187), .Z(n38188) );
  NANDN U38585 ( .A(n38189), .B(n38188), .Z(n38237) );
  XNOR U38586 ( .A(n38295), .B(n38237), .Z(n38238) );
  XOR U38587 ( .A(n38239), .B(n38238), .Z(n38254) );
  XOR U38588 ( .A(n38255), .B(n38254), .Z(n38257) );
  NAND U38589 ( .A(n38191), .B(n38190), .Z(n38195) );
  NAND U38590 ( .A(n38193), .B(n38192), .Z(n38194) );
  AND U38591 ( .A(n38195), .B(n38194), .Z(n38256) );
  XNOR U38592 ( .A(n38257), .B(n38256), .Z(n38230) );
  NAND U38593 ( .A(n38197), .B(n38196), .Z(n38201) );
  NAND U38594 ( .A(n38199), .B(n38198), .Z(n38200) );
  NAND U38595 ( .A(n38201), .B(n38200), .Z(n38229) );
  NAND U38596 ( .A(n38203), .B(n38202), .Z(n38207) );
  NAND U38597 ( .A(n38205), .B(n38204), .Z(n38206) );
  AND U38598 ( .A(n38207), .B(n38206), .Z(n38228) );
  NAND U38599 ( .A(n38209), .B(n38208), .Z(n38213) );
  NAND U38600 ( .A(n38211), .B(n38210), .Z(n38212) );
  AND U38601 ( .A(n38213), .B(n38212), .Z(n38223) );
  XOR U38602 ( .A(n38219), .B(n38218), .Z(n38214) );
  XOR U38603 ( .A(n38215), .B(n38214), .Z(c[502]) );
  AND U38604 ( .A(n38215), .B(n38214), .Z(n38261) );
  NAND U38605 ( .A(n38217), .B(n38216), .Z(n38221) );
  NANDN U38606 ( .A(n38219), .B(n38218), .Z(n38220) );
  AND U38607 ( .A(n38221), .B(n38220), .Z(n38265) );
  NAND U38608 ( .A(n38223), .B(n38222), .Z(n38227) );
  NAND U38609 ( .A(n38225), .B(n38224), .Z(n38226) );
  NAND U38610 ( .A(n38227), .B(n38226), .Z(n38263) );
  NAND U38611 ( .A(n38232), .B(n38231), .Z(n38236) );
  NAND U38612 ( .A(n38234), .B(n38233), .Z(n38235) );
  NAND U38613 ( .A(n38236), .B(n38235), .Z(n38277) );
  NAND U38614 ( .A(n38470), .B(n38240), .Z(n38242) );
  XOR U38615 ( .A(b[31]), .B(a[249]), .Z(n38286) );
  NAND U38616 ( .A(n38453), .B(n38286), .Z(n38241) );
  NAND U38617 ( .A(n38242), .B(n38241), .Z(n38310) );
  NAND U38618 ( .A(n38385), .B(n38243), .Z(n38245) );
  XOR U38619 ( .A(b[27]), .B(a[253]), .Z(n38304) );
  NAND U38620 ( .A(n38343), .B(n38304), .Z(n38244) );
  NAND U38621 ( .A(n38245), .B(n38244), .Z(n38308) );
  NAND U38622 ( .A(n38289), .B(n38246), .Z(n38249) );
  XOR U38623 ( .A(a[255]), .B(b[25]), .Z(n38290) );
  NAND U38624 ( .A(n38247), .B(n38290), .Z(n38248) );
  NAND U38625 ( .A(n38249), .B(n38248), .Z(n38281) );
  NAND U38626 ( .A(n194), .B(n38250), .Z(n38252) );
  XOR U38627 ( .A(b[29]), .B(a[251]), .Z(n38301) );
  NAND U38628 ( .A(n38456), .B(n38301), .Z(n38251) );
  NAND U38629 ( .A(n38252), .B(n38251), .Z(n38280) );
  AND U38630 ( .A(b[31]), .B(a[247]), .Z(n38297) );
  XNOR U38631 ( .A(n38253), .B(n38297), .Z(n38296) );
  XOR U38632 ( .A(n38295), .B(n38296), .Z(n38282) );
  XOR U38633 ( .A(n38283), .B(n38282), .Z(n38307) );
  NAND U38634 ( .A(n38255), .B(n38254), .Z(n38259) );
  NAND U38635 ( .A(n38257), .B(n38256), .Z(n38258) );
  NAND U38636 ( .A(n38259), .B(n38258), .Z(n38268) );
  XOR U38637 ( .A(n38269), .B(n38268), .Z(n38270) );
  XNOR U38638 ( .A(n38271), .B(n38270), .Z(n38262) );
  XOR U38639 ( .A(n38265), .B(n38264), .Z(n38260) );
  XOR U38640 ( .A(n38261), .B(n38260), .Z(c[503]) );
  AND U38641 ( .A(n38261), .B(n38260), .Z(n38314) );
  NAND U38642 ( .A(n38263), .B(n38262), .Z(n38267) );
  NANDN U38643 ( .A(n38265), .B(n38264), .Z(n38266) );
  AND U38644 ( .A(n38267), .B(n38266), .Z(n38318) );
  NAND U38645 ( .A(n38269), .B(n38268), .Z(n38273) );
  NANDN U38646 ( .A(n38271), .B(n38270), .Z(n38272) );
  NAND U38647 ( .A(n38273), .B(n38272), .Z(n38316) );
  NAND U38648 ( .A(n38275), .B(n38274), .Z(n38279) );
  NAND U38649 ( .A(n38277), .B(n38276), .Z(n38278) );
  AND U38650 ( .A(n38279), .B(n38278), .Z(n38324) );
  NAND U38651 ( .A(n38281), .B(n38280), .Z(n38285) );
  NAND U38652 ( .A(n38283), .B(n38282), .Z(n38284) );
  NAND U38653 ( .A(n38285), .B(n38284), .Z(n38328) );
  NAND U38654 ( .A(n38470), .B(n38286), .Z(n38288) );
  XOR U38655 ( .A(b[31]), .B(a[250]), .Z(n38349) );
  NAND U38656 ( .A(n38453), .B(n38349), .Z(n38287) );
  NAND U38657 ( .A(n38288), .B(n38287), .Z(n38341) );
  IV U38658 ( .A(n38341), .Z(n38294) );
  AND U38659 ( .A(b[31]), .B(a[248]), .Z(n38376) );
  AND U38660 ( .A(n38290), .B(n38289), .Z(n38293) );
  XOR U38661 ( .A(b[24]), .B(b[23]), .Z(n38291) );
  NAND U38662 ( .A(b[25]), .B(n38291), .Z(n38292) );
  NANDN U38663 ( .A(n38293), .B(n38292), .Z(n38339) );
  XNOR U38664 ( .A(n38376), .B(n38339), .Z(n38340) );
  XNOR U38665 ( .A(n38294), .B(n38340), .Z(n38327) );
  AND U38666 ( .A(n38296), .B(n38295), .Z(n38300) );
  NAND U38667 ( .A(n38298), .B(n38297), .Z(n38299) );
  NANDN U38668 ( .A(n38300), .B(n38299), .Z(n38336) );
  NAND U38669 ( .A(n194), .B(n38301), .Z(n38303) );
  XOR U38670 ( .A(b[29]), .B(a[252]), .Z(n38346) );
  NAND U38671 ( .A(n38456), .B(n38346), .Z(n38302) );
  NAND U38672 ( .A(n38303), .B(n38302), .Z(n38334) );
  NAND U38673 ( .A(n38385), .B(n38304), .Z(n38306) );
  XOR U38674 ( .A(b[27]), .B(a[254]), .Z(n38342) );
  NAND U38675 ( .A(n38343), .B(n38342), .Z(n38305) );
  NAND U38676 ( .A(n38306), .B(n38305), .Z(n38333) );
  XNOR U38677 ( .A(n38330), .B(n38329), .Z(n38322) );
  NAND U38678 ( .A(n38308), .B(n38307), .Z(n38312) );
  NAND U38679 ( .A(n38310), .B(n38309), .Z(n38311) );
  AND U38680 ( .A(n38312), .B(n38311), .Z(n38321) );
  XOR U38681 ( .A(n38324), .B(n38323), .Z(n38315) );
  XOR U38682 ( .A(n38318), .B(n38317), .Z(n38313) );
  XOR U38683 ( .A(n38314), .B(n38313), .Z(c[504]) );
  AND U38684 ( .A(n38314), .B(n38313), .Z(n38354) );
  NAND U38685 ( .A(n38316), .B(n38315), .Z(n38320) );
  NANDN U38686 ( .A(n38318), .B(n38317), .Z(n38319) );
  AND U38687 ( .A(n38320), .B(n38319), .Z(n38358) );
  NAND U38688 ( .A(n38322), .B(n38321), .Z(n38326) );
  NAND U38689 ( .A(n38324), .B(n38323), .Z(n38325) );
  NAND U38690 ( .A(n38326), .B(n38325), .Z(n38356) );
  NAND U38691 ( .A(n38328), .B(n38327), .Z(n38332) );
  NAND U38692 ( .A(n38330), .B(n38329), .Z(n38331) );
  AND U38693 ( .A(n38332), .B(n38331), .Z(n38393) );
  NAND U38694 ( .A(n38334), .B(n38333), .Z(n38338) );
  NAND U38695 ( .A(n38336), .B(n38335), .Z(n38337) );
  NAND U38696 ( .A(n38338), .B(n38337), .Z(n38391) );
  NAND U38697 ( .A(n38385), .B(n38342), .Z(n38345) );
  XOR U38698 ( .A(b[27]), .B(a[255]), .Z(n38386) );
  NAND U38699 ( .A(n38343), .B(n38386), .Z(n38344) );
  NAND U38700 ( .A(n38345), .B(n38344), .Z(n38362) );
  NAND U38701 ( .A(n194), .B(n38346), .Z(n38348) );
  XOR U38702 ( .A(b[29]), .B(a[253]), .Z(n38373) );
  NAND U38703 ( .A(n38456), .B(n38373), .Z(n38347) );
  NAND U38704 ( .A(n38348), .B(n38347), .Z(n38368) );
  NAND U38705 ( .A(n38470), .B(n38349), .Z(n38351) );
  XOR U38706 ( .A(b[31]), .B(a[251]), .Z(n38382) );
  NAND U38707 ( .A(n38453), .B(n38382), .Z(n38350) );
  NAND U38708 ( .A(n38351), .B(n38350), .Z(n38367) );
  AND U38709 ( .A(b[31]), .B(a[249]), .Z(n38378) );
  XNOR U38710 ( .A(n38352), .B(n38378), .Z(n38377) );
  XOR U38711 ( .A(n38376), .B(n38377), .Z(n38369) );
  XOR U38712 ( .A(n38370), .B(n38369), .Z(n38361) );
  XOR U38713 ( .A(n38393), .B(n38392), .Z(n38355) );
  XOR U38714 ( .A(n38358), .B(n38357), .Z(n38353) );
  XOR U38715 ( .A(n38354), .B(n38353), .Z(c[505]) );
  AND U38716 ( .A(n38354), .B(n38353), .Z(n38397) );
  NAND U38717 ( .A(n38356), .B(n38355), .Z(n38360) );
  NANDN U38718 ( .A(n38358), .B(n38357), .Z(n38359) );
  AND U38719 ( .A(n38360), .B(n38359), .Z(n38401) );
  NAND U38720 ( .A(n38362), .B(n38361), .Z(n38366) );
  NAND U38721 ( .A(n38364), .B(n38363), .Z(n38365) );
  NAND U38722 ( .A(n38366), .B(n38365), .Z(n38407) );
  NAND U38723 ( .A(n38368), .B(n38367), .Z(n38372) );
  NAND U38724 ( .A(n38370), .B(n38369), .Z(n38371) );
  NAND U38725 ( .A(n38372), .B(n38371), .Z(n38405) );
  NAND U38726 ( .A(n194), .B(n38373), .Z(n38375) );
  XOR U38727 ( .A(b[29]), .B(a[254]), .Z(n38419) );
  NAND U38728 ( .A(n38456), .B(n38419), .Z(n38374) );
  NAND U38729 ( .A(n38375), .B(n38374), .Z(n38411) );
  AND U38730 ( .A(n38377), .B(n38376), .Z(n38381) );
  NAND U38731 ( .A(n38379), .B(n38378), .Z(n38380) );
  NANDN U38732 ( .A(n38381), .B(n38380), .Z(n38410) );
  NAND U38733 ( .A(n38470), .B(n38382), .Z(n38384) );
  XOR U38734 ( .A(b[31]), .B(a[252]), .Z(n38416) );
  NAND U38735 ( .A(n38453), .B(n38416), .Z(n38383) );
  NAND U38736 ( .A(n38384), .B(n38383), .Z(n38423) );
  AND U38737 ( .A(b[31]), .B(a[250]), .Z(n38446) );
  AND U38738 ( .A(n38386), .B(n38385), .Z(n38389) );
  XOR U38739 ( .A(b[26]), .B(b[25]), .Z(n38387) );
  NAND U38740 ( .A(b[27]), .B(n38387), .Z(n38388) );
  NANDN U38741 ( .A(n38389), .B(n38388), .Z(n38420) );
  XNOR U38742 ( .A(n38446), .B(n38420), .Z(n38422) );
  XOR U38743 ( .A(n38413), .B(n38412), .Z(n38404) );
  NAND U38744 ( .A(n38391), .B(n38390), .Z(n38395) );
  NANDN U38745 ( .A(n38393), .B(n38392), .Z(n38394) );
  AND U38746 ( .A(n38395), .B(n38394), .Z(n38399) );
  XOR U38747 ( .A(n38398), .B(n38399), .Z(n38400) );
  XOR U38748 ( .A(n38401), .B(n38400), .Z(n38396) );
  XOR U38749 ( .A(n38397), .B(n38396), .Z(c[506]) );
  AND U38750 ( .A(n38397), .B(n38396), .Z(n38427) );
  NAND U38751 ( .A(n38399), .B(n38398), .Z(n38403) );
  NANDN U38752 ( .A(n38401), .B(n38400), .Z(n38402) );
  AND U38753 ( .A(n38403), .B(n38402), .Z(n38431) );
  NAND U38754 ( .A(n38405), .B(n38404), .Z(n38409) );
  NAND U38755 ( .A(n38407), .B(n38406), .Z(n38408) );
  AND U38756 ( .A(n38409), .B(n38408), .Z(n38429) );
  NAND U38757 ( .A(n38411), .B(n38410), .Z(n38415) );
  NAND U38758 ( .A(n38413), .B(n38412), .Z(n38414) );
  AND U38759 ( .A(n38415), .B(n38414), .Z(n38437) );
  NAND U38760 ( .A(n38470), .B(n38416), .Z(n38418) );
  XOR U38761 ( .A(b[31]), .B(a[253]), .Z(n38452) );
  NAND U38762 ( .A(n38453), .B(n38452), .Z(n38417) );
  NAND U38763 ( .A(n38418), .B(n38417), .Z(n38441) );
  XNOR U38764 ( .A(b[29]), .B(a[255]), .Z(n38457) );
  IV U38765 ( .A(n38446), .Z(n38421) );
  AND U38766 ( .A(b[31]), .B(a[251]), .Z(n38449) );
  XOR U38767 ( .A(n38448), .B(n38449), .Z(n38447) );
  XNOR U38768 ( .A(n38421), .B(n38447), .Z(n38442) );
  XNOR U38769 ( .A(n38443), .B(n38442), .Z(n38435) );
  NAND U38770 ( .A(n38421), .B(n38420), .Z(n38425) );
  NAND U38771 ( .A(n38423), .B(n38422), .Z(n38424) );
  AND U38772 ( .A(n38425), .B(n38424), .Z(n38434) );
  XOR U38773 ( .A(n38437), .B(n38436), .Z(n38428) );
  XOR U38774 ( .A(n38429), .B(n38428), .Z(n38430) );
  XOR U38775 ( .A(n38431), .B(n38430), .Z(n38426) );
  XOR U38776 ( .A(n38427), .B(n38426), .Z(c[507]) );
  AND U38777 ( .A(n38427), .B(n38426), .Z(n38461) );
  NAND U38778 ( .A(n38429), .B(n38428), .Z(n38433) );
  NANDN U38779 ( .A(n38431), .B(n38430), .Z(n38432) );
  AND U38780 ( .A(n38433), .B(n38432), .Z(n38465) );
  NAND U38781 ( .A(n38435), .B(n38434), .Z(n38439) );
  NAND U38782 ( .A(n38437), .B(n38436), .Z(n38438) );
  NAND U38783 ( .A(n38439), .B(n38438), .Z(n38463) );
  NAND U38784 ( .A(n38441), .B(n38440), .Z(n38445) );
  NAND U38785 ( .A(n38443), .B(n38442), .Z(n38444) );
  AND U38786 ( .A(n38445), .B(n38444), .Z(n38481) );
  AND U38787 ( .A(n38447), .B(n38446), .Z(n38451) );
  NAND U38788 ( .A(n38449), .B(n38448), .Z(n38450) );
  NANDN U38789 ( .A(n38451), .B(n38450), .Z(n38479) );
  NAND U38790 ( .A(n38470), .B(n38452), .Z(n38455) );
  XOR U38791 ( .A(b[31]), .B(a[254]), .Z(n38469) );
  NAND U38792 ( .A(n38453), .B(n38469), .Z(n38454) );
  NAND U38793 ( .A(n38455), .B(n38454), .Z(n38475) );
  NAND U38794 ( .A(n38456), .B(b[29]), .Z(n38459) );
  NANDN U38795 ( .A(n38457), .B(n194), .Z(n38458) );
  AND U38796 ( .A(n38459), .B(n38458), .Z(n38473) );
  AND U38797 ( .A(b[31]), .B(a[252]), .Z(n38468) );
  IV U38798 ( .A(n38468), .Z(n38488) );
  XNOR U38799 ( .A(n38473), .B(n38488), .Z(n38474) );
  XOR U38800 ( .A(n38481), .B(n38480), .Z(n38462) );
  XOR U38801 ( .A(n38465), .B(n38464), .Z(n38460) );
  XOR U38802 ( .A(n38461), .B(n38460), .Z(c[508]) );
  AND U38803 ( .A(n38461), .B(n38460), .Z(n38485) );
  NAND U38804 ( .A(n38463), .B(n38462), .Z(n38467) );
  NANDN U38805 ( .A(n38465), .B(n38464), .Z(n38466) );
  AND U38806 ( .A(n38467), .B(n38466), .Z(n38499) );
  AND U38807 ( .A(b[31]), .B(a[253]), .Z(n38487) );
  XNOR U38808 ( .A(n38486), .B(n38487), .Z(n38489) );
  XNOR U38809 ( .A(n38468), .B(n38489), .Z(n38502) );
  NAND U38810 ( .A(n38470), .B(n38469), .Z(n38472) );
  XNOR U38811 ( .A(b[31]), .B(a[255]), .Z(n38492) );
  OR U38812 ( .A(n38492), .B(n38493), .Z(n38471) );
  NAND U38813 ( .A(n38472), .B(n38471), .Z(n38503) );
  NANDN U38814 ( .A(n38473), .B(n38488), .Z(n38477) );
  NAND U38815 ( .A(n38475), .B(n38474), .Z(n38476) );
  NAND U38816 ( .A(n38477), .B(n38476), .Z(n38504) );
  XNOR U38817 ( .A(n38505), .B(n38504), .Z(n38497) );
  NAND U38818 ( .A(n38479), .B(n38478), .Z(n38483) );
  NANDN U38819 ( .A(n38481), .B(n38480), .Z(n38482) );
  AND U38820 ( .A(n38483), .B(n38482), .Z(n38496) );
  XOR U38821 ( .A(n38499), .B(n38498), .Z(n38484) );
  XOR U38822 ( .A(n38485), .B(n38484), .Z(c[509]) );
  AND U38823 ( .A(n38485), .B(n38484), .Z(n38509) );
  AND U38824 ( .A(n38487), .B(n38486), .Z(n38491) );
  OR U38825 ( .A(n38489), .B(n38488), .Z(n38490) );
  NANDN U38826 ( .A(n38491), .B(n38490), .Z(n38524) );
  NAND U38827 ( .A(b[31]), .B(a[254]), .Z(n38522) );
  OR U38828 ( .A(n38492), .B(n195), .Z(n38495) );
  NANDN U38829 ( .A(n38493), .B(b[31]), .Z(n38494) );
  NAND U38830 ( .A(n38495), .B(n38494), .Z(n38521) );
  XOR U38831 ( .A(n38522), .B(n38521), .Z(n38523) );
  NAND U38832 ( .A(n38497), .B(n38496), .Z(n38501) );
  NANDN U38833 ( .A(n38499), .B(n38498), .Z(n38500) );
  NAND U38834 ( .A(n38501), .B(n38500), .Z(n38510) );
  NAND U38835 ( .A(n38503), .B(n38502), .Z(n38507) );
  NAND U38836 ( .A(n38505), .B(n38504), .Z(n38506) );
  AND U38837 ( .A(n38507), .B(n38506), .Z(n38511) );
  XNOR U38838 ( .A(n38512), .B(n38513), .Z(n38508) );
  XOR U38839 ( .A(n38509), .B(n38508), .Z(c[510]) );
  NAND U38840 ( .A(n38509), .B(n38508), .Z(n38517) );
  AND U38841 ( .A(n38511), .B(n38510), .Z(n38515) );
  AND U38842 ( .A(n38513), .B(n38512), .Z(n38514) );
  OR U38843 ( .A(n38515), .B(n38514), .Z(n38516) );
  AND U38844 ( .A(n38517), .B(n38516), .Z(n38530) );
  XNOR U38845 ( .A(a[254]), .B(a[255]), .Z(n38518) );
  XNOR U38846 ( .A(n38519), .B(n38518), .Z(n38520) );
  ANDN U38847 ( .B(b[31]), .A(n38520), .Z(n38528) );
  AND U38848 ( .A(n38522), .B(n38521), .Z(n38526) );
  AND U38849 ( .A(n38524), .B(n38523), .Z(n38525) );
  OR U38850 ( .A(n38526), .B(n38525), .Z(n38527) );
  XNOR U38851 ( .A(n38528), .B(n38527), .Z(n38529) );
  XNOR U38852 ( .A(n38530), .B(n38529), .Z(c[511]) );
endmodule

