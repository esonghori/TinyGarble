
module mult_N256_CC128 ( clk, rst, a, b, c );
  input [255:0] a;
  input [1:0] b;
  output [511:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063;
  wire   [511:0] sreg;

  DFF \sreg_reg[509]  ( .D(c[511]), .CLK(clk), .RST(rst), .Q(sreg[509]) );
  DFF \sreg_reg[508]  ( .D(c[510]), .CLK(clk), .RST(rst), .Q(sreg[508]) );
  DFF \sreg_reg[507]  ( .D(c[509]), .CLK(clk), .RST(rst), .Q(sreg[507]) );
  DFF \sreg_reg[506]  ( .D(c[508]), .CLK(clk), .RST(rst), .Q(sreg[506]) );
  DFF \sreg_reg[505]  ( .D(c[507]), .CLK(clk), .RST(rst), .Q(sreg[505]) );
  DFF \sreg_reg[504]  ( .D(c[506]), .CLK(clk), .RST(rst), .Q(sreg[504]) );
  DFF \sreg_reg[503]  ( .D(c[505]), .CLK(clk), .RST(rst), .Q(sreg[503]) );
  DFF \sreg_reg[502]  ( .D(c[504]), .CLK(clk), .RST(rst), .Q(sreg[502]) );
  DFF \sreg_reg[501]  ( .D(c[503]), .CLK(clk), .RST(rst), .Q(sreg[501]) );
  DFF \sreg_reg[500]  ( .D(c[502]), .CLK(clk), .RST(rst), .Q(sreg[500]) );
  DFF \sreg_reg[499]  ( .D(c[501]), .CLK(clk), .RST(rst), .Q(sreg[499]) );
  DFF \sreg_reg[498]  ( .D(c[500]), .CLK(clk), .RST(rst), .Q(sreg[498]) );
  DFF \sreg_reg[497]  ( .D(c[499]), .CLK(clk), .RST(rst), .Q(sreg[497]) );
  DFF \sreg_reg[496]  ( .D(c[498]), .CLK(clk), .RST(rst), .Q(sreg[496]) );
  DFF \sreg_reg[495]  ( .D(c[497]), .CLK(clk), .RST(rst), .Q(sreg[495]) );
  DFF \sreg_reg[494]  ( .D(c[496]), .CLK(clk), .RST(rst), .Q(sreg[494]) );
  DFF \sreg_reg[493]  ( .D(c[495]), .CLK(clk), .RST(rst), .Q(sreg[493]) );
  DFF \sreg_reg[492]  ( .D(c[494]), .CLK(clk), .RST(rst), .Q(sreg[492]) );
  DFF \sreg_reg[491]  ( .D(c[493]), .CLK(clk), .RST(rst), .Q(sreg[491]) );
  DFF \sreg_reg[490]  ( .D(c[492]), .CLK(clk), .RST(rst), .Q(sreg[490]) );
  DFF \sreg_reg[489]  ( .D(c[491]), .CLK(clk), .RST(rst), .Q(sreg[489]) );
  DFF \sreg_reg[488]  ( .D(c[490]), .CLK(clk), .RST(rst), .Q(sreg[488]) );
  DFF \sreg_reg[487]  ( .D(c[489]), .CLK(clk), .RST(rst), .Q(sreg[487]) );
  DFF \sreg_reg[486]  ( .D(c[488]), .CLK(clk), .RST(rst), .Q(sreg[486]) );
  DFF \sreg_reg[485]  ( .D(c[487]), .CLK(clk), .RST(rst), .Q(sreg[485]) );
  DFF \sreg_reg[484]  ( .D(c[486]), .CLK(clk), .RST(rst), .Q(sreg[484]) );
  DFF \sreg_reg[483]  ( .D(c[485]), .CLK(clk), .RST(rst), .Q(sreg[483]) );
  DFF \sreg_reg[482]  ( .D(c[484]), .CLK(clk), .RST(rst), .Q(sreg[482]) );
  DFF \sreg_reg[481]  ( .D(c[483]), .CLK(clk), .RST(rst), .Q(sreg[481]) );
  DFF \sreg_reg[480]  ( .D(c[482]), .CLK(clk), .RST(rst), .Q(sreg[480]) );
  DFF \sreg_reg[479]  ( .D(c[481]), .CLK(clk), .RST(rst), .Q(sreg[479]) );
  DFF \sreg_reg[478]  ( .D(c[480]), .CLK(clk), .RST(rst), .Q(sreg[478]) );
  DFF \sreg_reg[477]  ( .D(c[479]), .CLK(clk), .RST(rst), .Q(sreg[477]) );
  DFF \sreg_reg[476]  ( .D(c[478]), .CLK(clk), .RST(rst), .Q(sreg[476]) );
  DFF \sreg_reg[475]  ( .D(c[477]), .CLK(clk), .RST(rst), .Q(sreg[475]) );
  DFF \sreg_reg[474]  ( .D(c[476]), .CLK(clk), .RST(rst), .Q(sreg[474]) );
  DFF \sreg_reg[473]  ( .D(c[475]), .CLK(clk), .RST(rst), .Q(sreg[473]) );
  DFF \sreg_reg[472]  ( .D(c[474]), .CLK(clk), .RST(rst), .Q(sreg[472]) );
  DFF \sreg_reg[471]  ( .D(c[473]), .CLK(clk), .RST(rst), .Q(sreg[471]) );
  DFF \sreg_reg[470]  ( .D(c[472]), .CLK(clk), .RST(rst), .Q(sreg[470]) );
  DFF \sreg_reg[469]  ( .D(c[471]), .CLK(clk), .RST(rst), .Q(sreg[469]) );
  DFF \sreg_reg[468]  ( .D(c[470]), .CLK(clk), .RST(rst), .Q(sreg[468]) );
  DFF \sreg_reg[467]  ( .D(c[469]), .CLK(clk), .RST(rst), .Q(sreg[467]) );
  DFF \sreg_reg[466]  ( .D(c[468]), .CLK(clk), .RST(rst), .Q(sreg[466]) );
  DFF \sreg_reg[465]  ( .D(c[467]), .CLK(clk), .RST(rst), .Q(sreg[465]) );
  DFF \sreg_reg[464]  ( .D(c[466]), .CLK(clk), .RST(rst), .Q(sreg[464]) );
  DFF \sreg_reg[463]  ( .D(c[465]), .CLK(clk), .RST(rst), .Q(sreg[463]) );
  DFF \sreg_reg[462]  ( .D(c[464]), .CLK(clk), .RST(rst), .Q(sreg[462]) );
  DFF \sreg_reg[461]  ( .D(c[463]), .CLK(clk), .RST(rst), .Q(sreg[461]) );
  DFF \sreg_reg[460]  ( .D(c[462]), .CLK(clk), .RST(rst), .Q(sreg[460]) );
  DFF \sreg_reg[459]  ( .D(c[461]), .CLK(clk), .RST(rst), .Q(sreg[459]) );
  DFF \sreg_reg[458]  ( .D(c[460]), .CLK(clk), .RST(rst), .Q(sreg[458]) );
  DFF \sreg_reg[457]  ( .D(c[459]), .CLK(clk), .RST(rst), .Q(sreg[457]) );
  DFF \sreg_reg[456]  ( .D(c[458]), .CLK(clk), .RST(rst), .Q(sreg[456]) );
  DFF \sreg_reg[455]  ( .D(c[457]), .CLK(clk), .RST(rst), .Q(sreg[455]) );
  DFF \sreg_reg[454]  ( .D(c[456]), .CLK(clk), .RST(rst), .Q(sreg[454]) );
  DFF \sreg_reg[453]  ( .D(c[455]), .CLK(clk), .RST(rst), .Q(sreg[453]) );
  DFF \sreg_reg[452]  ( .D(c[454]), .CLK(clk), .RST(rst), .Q(sreg[452]) );
  DFF \sreg_reg[451]  ( .D(c[453]), .CLK(clk), .RST(rst), .Q(sreg[451]) );
  DFF \sreg_reg[450]  ( .D(c[452]), .CLK(clk), .RST(rst), .Q(sreg[450]) );
  DFF \sreg_reg[449]  ( .D(c[451]), .CLK(clk), .RST(rst), .Q(sreg[449]) );
  DFF \sreg_reg[448]  ( .D(c[450]), .CLK(clk), .RST(rst), .Q(sreg[448]) );
  DFF \sreg_reg[447]  ( .D(c[449]), .CLK(clk), .RST(rst), .Q(sreg[447]) );
  DFF \sreg_reg[446]  ( .D(c[448]), .CLK(clk), .RST(rst), .Q(sreg[446]) );
  DFF \sreg_reg[445]  ( .D(c[447]), .CLK(clk), .RST(rst), .Q(sreg[445]) );
  DFF \sreg_reg[444]  ( .D(c[446]), .CLK(clk), .RST(rst), .Q(sreg[444]) );
  DFF \sreg_reg[443]  ( .D(c[445]), .CLK(clk), .RST(rst), .Q(sreg[443]) );
  DFF \sreg_reg[442]  ( .D(c[444]), .CLK(clk), .RST(rst), .Q(sreg[442]) );
  DFF \sreg_reg[441]  ( .D(c[443]), .CLK(clk), .RST(rst), .Q(sreg[441]) );
  DFF \sreg_reg[440]  ( .D(c[442]), .CLK(clk), .RST(rst), .Q(sreg[440]) );
  DFF \sreg_reg[439]  ( .D(c[441]), .CLK(clk), .RST(rst), .Q(sreg[439]) );
  DFF \sreg_reg[438]  ( .D(c[440]), .CLK(clk), .RST(rst), .Q(sreg[438]) );
  DFF \sreg_reg[437]  ( .D(c[439]), .CLK(clk), .RST(rst), .Q(sreg[437]) );
  DFF \sreg_reg[436]  ( .D(c[438]), .CLK(clk), .RST(rst), .Q(sreg[436]) );
  DFF \sreg_reg[435]  ( .D(c[437]), .CLK(clk), .RST(rst), .Q(sreg[435]) );
  DFF \sreg_reg[434]  ( .D(c[436]), .CLK(clk), .RST(rst), .Q(sreg[434]) );
  DFF \sreg_reg[433]  ( .D(c[435]), .CLK(clk), .RST(rst), .Q(sreg[433]) );
  DFF \sreg_reg[432]  ( .D(c[434]), .CLK(clk), .RST(rst), .Q(sreg[432]) );
  DFF \sreg_reg[431]  ( .D(c[433]), .CLK(clk), .RST(rst), .Q(sreg[431]) );
  DFF \sreg_reg[430]  ( .D(c[432]), .CLK(clk), .RST(rst), .Q(sreg[430]) );
  DFF \sreg_reg[429]  ( .D(c[431]), .CLK(clk), .RST(rst), .Q(sreg[429]) );
  DFF \sreg_reg[428]  ( .D(c[430]), .CLK(clk), .RST(rst), .Q(sreg[428]) );
  DFF \sreg_reg[427]  ( .D(c[429]), .CLK(clk), .RST(rst), .Q(sreg[427]) );
  DFF \sreg_reg[426]  ( .D(c[428]), .CLK(clk), .RST(rst), .Q(sreg[426]) );
  DFF \sreg_reg[425]  ( .D(c[427]), .CLK(clk), .RST(rst), .Q(sreg[425]) );
  DFF \sreg_reg[424]  ( .D(c[426]), .CLK(clk), .RST(rst), .Q(sreg[424]) );
  DFF \sreg_reg[423]  ( .D(c[425]), .CLK(clk), .RST(rst), .Q(sreg[423]) );
  DFF \sreg_reg[422]  ( .D(c[424]), .CLK(clk), .RST(rst), .Q(sreg[422]) );
  DFF \sreg_reg[421]  ( .D(c[423]), .CLK(clk), .RST(rst), .Q(sreg[421]) );
  DFF \sreg_reg[420]  ( .D(c[422]), .CLK(clk), .RST(rst), .Q(sreg[420]) );
  DFF \sreg_reg[419]  ( .D(c[421]), .CLK(clk), .RST(rst), .Q(sreg[419]) );
  DFF \sreg_reg[418]  ( .D(c[420]), .CLK(clk), .RST(rst), .Q(sreg[418]) );
  DFF \sreg_reg[417]  ( .D(c[419]), .CLK(clk), .RST(rst), .Q(sreg[417]) );
  DFF \sreg_reg[416]  ( .D(c[418]), .CLK(clk), .RST(rst), .Q(sreg[416]) );
  DFF \sreg_reg[415]  ( .D(c[417]), .CLK(clk), .RST(rst), .Q(sreg[415]) );
  DFF \sreg_reg[414]  ( .D(c[416]), .CLK(clk), .RST(rst), .Q(sreg[414]) );
  DFF \sreg_reg[413]  ( .D(c[415]), .CLK(clk), .RST(rst), .Q(sreg[413]) );
  DFF \sreg_reg[412]  ( .D(c[414]), .CLK(clk), .RST(rst), .Q(sreg[412]) );
  DFF \sreg_reg[411]  ( .D(c[413]), .CLK(clk), .RST(rst), .Q(sreg[411]) );
  DFF \sreg_reg[410]  ( .D(c[412]), .CLK(clk), .RST(rst), .Q(sreg[410]) );
  DFF \sreg_reg[409]  ( .D(c[411]), .CLK(clk), .RST(rst), .Q(sreg[409]) );
  DFF \sreg_reg[408]  ( .D(c[410]), .CLK(clk), .RST(rst), .Q(sreg[408]) );
  DFF \sreg_reg[407]  ( .D(c[409]), .CLK(clk), .RST(rst), .Q(sreg[407]) );
  DFF \sreg_reg[406]  ( .D(c[408]), .CLK(clk), .RST(rst), .Q(sreg[406]) );
  DFF \sreg_reg[405]  ( .D(c[407]), .CLK(clk), .RST(rst), .Q(sreg[405]) );
  DFF \sreg_reg[404]  ( .D(c[406]), .CLK(clk), .RST(rst), .Q(sreg[404]) );
  DFF \sreg_reg[403]  ( .D(c[405]), .CLK(clk), .RST(rst), .Q(sreg[403]) );
  DFF \sreg_reg[402]  ( .D(c[404]), .CLK(clk), .RST(rst), .Q(sreg[402]) );
  DFF \sreg_reg[401]  ( .D(c[403]), .CLK(clk), .RST(rst), .Q(sreg[401]) );
  DFF \sreg_reg[400]  ( .D(c[402]), .CLK(clk), .RST(rst), .Q(sreg[400]) );
  DFF \sreg_reg[399]  ( .D(c[401]), .CLK(clk), .RST(rst), .Q(sreg[399]) );
  DFF \sreg_reg[398]  ( .D(c[400]), .CLK(clk), .RST(rst), .Q(sreg[398]) );
  DFF \sreg_reg[397]  ( .D(c[399]), .CLK(clk), .RST(rst), .Q(sreg[397]) );
  DFF \sreg_reg[396]  ( .D(c[398]), .CLK(clk), .RST(rst), .Q(sreg[396]) );
  DFF \sreg_reg[395]  ( .D(c[397]), .CLK(clk), .RST(rst), .Q(sreg[395]) );
  DFF \sreg_reg[394]  ( .D(c[396]), .CLK(clk), .RST(rst), .Q(sreg[394]) );
  DFF \sreg_reg[393]  ( .D(c[395]), .CLK(clk), .RST(rst), .Q(sreg[393]) );
  DFF \sreg_reg[392]  ( .D(c[394]), .CLK(clk), .RST(rst), .Q(sreg[392]) );
  DFF \sreg_reg[391]  ( .D(c[393]), .CLK(clk), .RST(rst), .Q(sreg[391]) );
  DFF \sreg_reg[390]  ( .D(c[392]), .CLK(clk), .RST(rst), .Q(sreg[390]) );
  DFF \sreg_reg[389]  ( .D(c[391]), .CLK(clk), .RST(rst), .Q(sreg[389]) );
  DFF \sreg_reg[388]  ( .D(c[390]), .CLK(clk), .RST(rst), .Q(sreg[388]) );
  DFF \sreg_reg[387]  ( .D(c[389]), .CLK(clk), .RST(rst), .Q(sreg[387]) );
  DFF \sreg_reg[386]  ( .D(c[388]), .CLK(clk), .RST(rst), .Q(sreg[386]) );
  DFF \sreg_reg[385]  ( .D(c[387]), .CLK(clk), .RST(rst), .Q(sreg[385]) );
  DFF \sreg_reg[384]  ( .D(c[386]), .CLK(clk), .RST(rst), .Q(sreg[384]) );
  DFF \sreg_reg[383]  ( .D(c[385]), .CLK(clk), .RST(rst), .Q(sreg[383]) );
  DFF \sreg_reg[382]  ( .D(c[384]), .CLK(clk), .RST(rst), .Q(sreg[382]) );
  DFF \sreg_reg[381]  ( .D(c[383]), .CLK(clk), .RST(rst), .Q(sreg[381]) );
  DFF \sreg_reg[380]  ( .D(c[382]), .CLK(clk), .RST(rst), .Q(sreg[380]) );
  DFF \sreg_reg[379]  ( .D(c[381]), .CLK(clk), .RST(rst), .Q(sreg[379]) );
  DFF \sreg_reg[378]  ( .D(c[380]), .CLK(clk), .RST(rst), .Q(sreg[378]) );
  DFF \sreg_reg[377]  ( .D(c[379]), .CLK(clk), .RST(rst), .Q(sreg[377]) );
  DFF \sreg_reg[376]  ( .D(c[378]), .CLK(clk), .RST(rst), .Q(sreg[376]) );
  DFF \sreg_reg[375]  ( .D(c[377]), .CLK(clk), .RST(rst), .Q(sreg[375]) );
  DFF \sreg_reg[374]  ( .D(c[376]), .CLK(clk), .RST(rst), .Q(sreg[374]) );
  DFF \sreg_reg[373]  ( .D(c[375]), .CLK(clk), .RST(rst), .Q(sreg[373]) );
  DFF \sreg_reg[372]  ( .D(c[374]), .CLK(clk), .RST(rst), .Q(sreg[372]) );
  DFF \sreg_reg[371]  ( .D(c[373]), .CLK(clk), .RST(rst), .Q(sreg[371]) );
  DFF \sreg_reg[370]  ( .D(c[372]), .CLK(clk), .RST(rst), .Q(sreg[370]) );
  DFF \sreg_reg[369]  ( .D(c[371]), .CLK(clk), .RST(rst), .Q(sreg[369]) );
  DFF \sreg_reg[368]  ( .D(c[370]), .CLK(clk), .RST(rst), .Q(sreg[368]) );
  DFF \sreg_reg[367]  ( .D(c[369]), .CLK(clk), .RST(rst), .Q(sreg[367]) );
  DFF \sreg_reg[366]  ( .D(c[368]), .CLK(clk), .RST(rst), .Q(sreg[366]) );
  DFF \sreg_reg[365]  ( .D(c[367]), .CLK(clk), .RST(rst), .Q(sreg[365]) );
  DFF \sreg_reg[364]  ( .D(c[366]), .CLK(clk), .RST(rst), .Q(sreg[364]) );
  DFF \sreg_reg[363]  ( .D(c[365]), .CLK(clk), .RST(rst), .Q(sreg[363]) );
  DFF \sreg_reg[362]  ( .D(c[364]), .CLK(clk), .RST(rst), .Q(sreg[362]) );
  DFF \sreg_reg[361]  ( .D(c[363]), .CLK(clk), .RST(rst), .Q(sreg[361]) );
  DFF \sreg_reg[360]  ( .D(c[362]), .CLK(clk), .RST(rst), .Q(sreg[360]) );
  DFF \sreg_reg[359]  ( .D(c[361]), .CLK(clk), .RST(rst), .Q(sreg[359]) );
  DFF \sreg_reg[358]  ( .D(c[360]), .CLK(clk), .RST(rst), .Q(sreg[358]) );
  DFF \sreg_reg[357]  ( .D(c[359]), .CLK(clk), .RST(rst), .Q(sreg[357]) );
  DFF \sreg_reg[356]  ( .D(c[358]), .CLK(clk), .RST(rst), .Q(sreg[356]) );
  DFF \sreg_reg[355]  ( .D(c[357]), .CLK(clk), .RST(rst), .Q(sreg[355]) );
  DFF \sreg_reg[354]  ( .D(c[356]), .CLK(clk), .RST(rst), .Q(sreg[354]) );
  DFF \sreg_reg[353]  ( .D(c[355]), .CLK(clk), .RST(rst), .Q(sreg[353]) );
  DFF \sreg_reg[352]  ( .D(c[354]), .CLK(clk), .RST(rst), .Q(sreg[352]) );
  DFF \sreg_reg[351]  ( .D(c[353]), .CLK(clk), .RST(rst), .Q(sreg[351]) );
  DFF \sreg_reg[350]  ( .D(c[352]), .CLK(clk), .RST(rst), .Q(sreg[350]) );
  DFF \sreg_reg[349]  ( .D(c[351]), .CLK(clk), .RST(rst), .Q(sreg[349]) );
  DFF \sreg_reg[348]  ( .D(c[350]), .CLK(clk), .RST(rst), .Q(sreg[348]) );
  DFF \sreg_reg[347]  ( .D(c[349]), .CLK(clk), .RST(rst), .Q(sreg[347]) );
  DFF \sreg_reg[346]  ( .D(c[348]), .CLK(clk), .RST(rst), .Q(sreg[346]) );
  DFF \sreg_reg[345]  ( .D(c[347]), .CLK(clk), .RST(rst), .Q(sreg[345]) );
  DFF \sreg_reg[344]  ( .D(c[346]), .CLK(clk), .RST(rst), .Q(sreg[344]) );
  DFF \sreg_reg[343]  ( .D(c[345]), .CLK(clk), .RST(rst), .Q(sreg[343]) );
  DFF \sreg_reg[342]  ( .D(c[344]), .CLK(clk), .RST(rst), .Q(sreg[342]) );
  DFF \sreg_reg[341]  ( .D(c[343]), .CLK(clk), .RST(rst), .Q(sreg[341]) );
  DFF \sreg_reg[340]  ( .D(c[342]), .CLK(clk), .RST(rst), .Q(sreg[340]) );
  DFF \sreg_reg[339]  ( .D(c[341]), .CLK(clk), .RST(rst), .Q(sreg[339]) );
  DFF \sreg_reg[338]  ( .D(c[340]), .CLK(clk), .RST(rst), .Q(sreg[338]) );
  DFF \sreg_reg[337]  ( .D(c[339]), .CLK(clk), .RST(rst), .Q(sreg[337]) );
  DFF \sreg_reg[336]  ( .D(c[338]), .CLK(clk), .RST(rst), .Q(sreg[336]) );
  DFF \sreg_reg[335]  ( .D(c[337]), .CLK(clk), .RST(rst), .Q(sreg[335]) );
  DFF \sreg_reg[334]  ( .D(c[336]), .CLK(clk), .RST(rst), .Q(sreg[334]) );
  DFF \sreg_reg[333]  ( .D(c[335]), .CLK(clk), .RST(rst), .Q(sreg[333]) );
  DFF \sreg_reg[332]  ( .D(c[334]), .CLK(clk), .RST(rst), .Q(sreg[332]) );
  DFF \sreg_reg[331]  ( .D(c[333]), .CLK(clk), .RST(rst), .Q(sreg[331]) );
  DFF \sreg_reg[330]  ( .D(c[332]), .CLK(clk), .RST(rst), .Q(sreg[330]) );
  DFF \sreg_reg[329]  ( .D(c[331]), .CLK(clk), .RST(rst), .Q(sreg[329]) );
  DFF \sreg_reg[328]  ( .D(c[330]), .CLK(clk), .RST(rst), .Q(sreg[328]) );
  DFF \sreg_reg[327]  ( .D(c[329]), .CLK(clk), .RST(rst), .Q(sreg[327]) );
  DFF \sreg_reg[326]  ( .D(c[328]), .CLK(clk), .RST(rst), .Q(sreg[326]) );
  DFF \sreg_reg[325]  ( .D(c[327]), .CLK(clk), .RST(rst), .Q(sreg[325]) );
  DFF \sreg_reg[324]  ( .D(c[326]), .CLK(clk), .RST(rst), .Q(sreg[324]) );
  DFF \sreg_reg[323]  ( .D(c[325]), .CLK(clk), .RST(rst), .Q(sreg[323]) );
  DFF \sreg_reg[322]  ( .D(c[324]), .CLK(clk), .RST(rst), .Q(sreg[322]) );
  DFF \sreg_reg[321]  ( .D(c[323]), .CLK(clk), .RST(rst), .Q(sreg[321]) );
  DFF \sreg_reg[320]  ( .D(c[322]), .CLK(clk), .RST(rst), .Q(sreg[320]) );
  DFF \sreg_reg[319]  ( .D(c[321]), .CLK(clk), .RST(rst), .Q(sreg[319]) );
  DFF \sreg_reg[318]  ( .D(c[320]), .CLK(clk), .RST(rst), .Q(sreg[318]) );
  DFF \sreg_reg[317]  ( .D(c[319]), .CLK(clk), .RST(rst), .Q(sreg[317]) );
  DFF \sreg_reg[316]  ( .D(c[318]), .CLK(clk), .RST(rst), .Q(sreg[316]) );
  DFF \sreg_reg[315]  ( .D(c[317]), .CLK(clk), .RST(rst), .Q(sreg[315]) );
  DFF \sreg_reg[314]  ( .D(c[316]), .CLK(clk), .RST(rst), .Q(sreg[314]) );
  DFF \sreg_reg[313]  ( .D(c[315]), .CLK(clk), .RST(rst), .Q(sreg[313]) );
  DFF \sreg_reg[312]  ( .D(c[314]), .CLK(clk), .RST(rst), .Q(sreg[312]) );
  DFF \sreg_reg[311]  ( .D(c[313]), .CLK(clk), .RST(rst), .Q(sreg[311]) );
  DFF \sreg_reg[310]  ( .D(c[312]), .CLK(clk), .RST(rst), .Q(sreg[310]) );
  DFF \sreg_reg[309]  ( .D(c[311]), .CLK(clk), .RST(rst), .Q(sreg[309]) );
  DFF \sreg_reg[308]  ( .D(c[310]), .CLK(clk), .RST(rst), .Q(sreg[308]) );
  DFF \sreg_reg[307]  ( .D(c[309]), .CLK(clk), .RST(rst), .Q(sreg[307]) );
  DFF \sreg_reg[306]  ( .D(c[308]), .CLK(clk), .RST(rst), .Q(sreg[306]) );
  DFF \sreg_reg[305]  ( .D(c[307]), .CLK(clk), .RST(rst), .Q(sreg[305]) );
  DFF \sreg_reg[304]  ( .D(c[306]), .CLK(clk), .RST(rst), .Q(sreg[304]) );
  DFF \sreg_reg[303]  ( .D(c[305]), .CLK(clk), .RST(rst), .Q(sreg[303]) );
  DFF \sreg_reg[302]  ( .D(c[304]), .CLK(clk), .RST(rst), .Q(sreg[302]) );
  DFF \sreg_reg[301]  ( .D(c[303]), .CLK(clk), .RST(rst), .Q(sreg[301]) );
  DFF \sreg_reg[300]  ( .D(c[302]), .CLK(clk), .RST(rst), .Q(sreg[300]) );
  DFF \sreg_reg[299]  ( .D(c[301]), .CLK(clk), .RST(rst), .Q(sreg[299]) );
  DFF \sreg_reg[298]  ( .D(c[300]), .CLK(clk), .RST(rst), .Q(sreg[298]) );
  DFF \sreg_reg[297]  ( .D(c[299]), .CLK(clk), .RST(rst), .Q(sreg[297]) );
  DFF \sreg_reg[296]  ( .D(c[298]), .CLK(clk), .RST(rst), .Q(sreg[296]) );
  DFF \sreg_reg[295]  ( .D(c[297]), .CLK(clk), .RST(rst), .Q(sreg[295]) );
  DFF \sreg_reg[294]  ( .D(c[296]), .CLK(clk), .RST(rst), .Q(sreg[294]) );
  DFF \sreg_reg[293]  ( .D(c[295]), .CLK(clk), .RST(rst), .Q(sreg[293]) );
  DFF \sreg_reg[292]  ( .D(c[294]), .CLK(clk), .RST(rst), .Q(sreg[292]) );
  DFF \sreg_reg[291]  ( .D(c[293]), .CLK(clk), .RST(rst), .Q(sreg[291]) );
  DFF \sreg_reg[290]  ( .D(c[292]), .CLK(clk), .RST(rst), .Q(sreg[290]) );
  DFF \sreg_reg[289]  ( .D(c[291]), .CLK(clk), .RST(rst), .Q(sreg[289]) );
  DFF \sreg_reg[288]  ( .D(c[290]), .CLK(clk), .RST(rst), .Q(sreg[288]) );
  DFF \sreg_reg[287]  ( .D(c[289]), .CLK(clk), .RST(rst), .Q(sreg[287]) );
  DFF \sreg_reg[286]  ( .D(c[288]), .CLK(clk), .RST(rst), .Q(sreg[286]) );
  DFF \sreg_reg[285]  ( .D(c[287]), .CLK(clk), .RST(rst), .Q(sreg[285]) );
  DFF \sreg_reg[284]  ( .D(c[286]), .CLK(clk), .RST(rst), .Q(sreg[284]) );
  DFF \sreg_reg[283]  ( .D(c[285]), .CLK(clk), .RST(rst), .Q(sreg[283]) );
  DFF \sreg_reg[282]  ( .D(c[284]), .CLK(clk), .RST(rst), .Q(sreg[282]) );
  DFF \sreg_reg[281]  ( .D(c[283]), .CLK(clk), .RST(rst), .Q(sreg[281]) );
  DFF \sreg_reg[280]  ( .D(c[282]), .CLK(clk), .RST(rst), .Q(sreg[280]) );
  DFF \sreg_reg[279]  ( .D(c[281]), .CLK(clk), .RST(rst), .Q(sreg[279]) );
  DFF \sreg_reg[278]  ( .D(c[280]), .CLK(clk), .RST(rst), .Q(sreg[278]) );
  DFF \sreg_reg[277]  ( .D(c[279]), .CLK(clk), .RST(rst), .Q(sreg[277]) );
  DFF \sreg_reg[276]  ( .D(c[278]), .CLK(clk), .RST(rst), .Q(sreg[276]) );
  DFF \sreg_reg[275]  ( .D(c[277]), .CLK(clk), .RST(rst), .Q(sreg[275]) );
  DFF \sreg_reg[274]  ( .D(c[276]), .CLK(clk), .RST(rst), .Q(sreg[274]) );
  DFF \sreg_reg[273]  ( .D(c[275]), .CLK(clk), .RST(rst), .Q(sreg[273]) );
  DFF \sreg_reg[272]  ( .D(c[274]), .CLK(clk), .RST(rst), .Q(sreg[272]) );
  DFF \sreg_reg[271]  ( .D(c[273]), .CLK(clk), .RST(rst), .Q(sreg[271]) );
  DFF \sreg_reg[270]  ( .D(c[272]), .CLK(clk), .RST(rst), .Q(sreg[270]) );
  DFF \sreg_reg[269]  ( .D(c[271]), .CLK(clk), .RST(rst), .Q(sreg[269]) );
  DFF \sreg_reg[268]  ( .D(c[270]), .CLK(clk), .RST(rst), .Q(sreg[268]) );
  DFF \sreg_reg[267]  ( .D(c[269]), .CLK(clk), .RST(rst), .Q(sreg[267]) );
  DFF \sreg_reg[266]  ( .D(c[268]), .CLK(clk), .RST(rst), .Q(sreg[266]) );
  DFF \sreg_reg[265]  ( .D(c[267]), .CLK(clk), .RST(rst), .Q(sreg[265]) );
  DFF \sreg_reg[264]  ( .D(c[266]), .CLK(clk), .RST(rst), .Q(sreg[264]) );
  DFF \sreg_reg[263]  ( .D(c[265]), .CLK(clk), .RST(rst), .Q(sreg[263]) );
  DFF \sreg_reg[262]  ( .D(c[264]), .CLK(clk), .RST(rst), .Q(sreg[262]) );
  DFF \sreg_reg[261]  ( .D(c[263]), .CLK(clk), .RST(rst), .Q(sreg[261]) );
  DFF \sreg_reg[260]  ( .D(c[262]), .CLK(clk), .RST(rst), .Q(sreg[260]) );
  DFF \sreg_reg[259]  ( .D(c[261]), .CLK(clk), .RST(rst), .Q(sreg[259]) );
  DFF \sreg_reg[258]  ( .D(c[260]), .CLK(clk), .RST(rst), .Q(sreg[258]) );
  DFF \sreg_reg[257]  ( .D(c[259]), .CLK(clk), .RST(rst), .Q(sreg[257]) );
  DFF \sreg_reg[256]  ( .D(c[258]), .CLK(clk), .RST(rst), .Q(sreg[256]) );
  DFF \sreg_reg[255]  ( .D(c[257]), .CLK(clk), .RST(rst), .Q(sreg[255]) );
  DFF \sreg_reg[254]  ( .D(c[256]), .CLK(clk), .RST(rst), .Q(sreg[254]) );
  DFF \sreg_reg[253]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(c[253]) );
  DFF \sreg_reg[252]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(c[252]) );
  DFF \sreg_reg[251]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(c[251]) );
  DFF \sreg_reg[250]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(c[250]) );
  DFF \sreg_reg[249]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(c[249]) );
  DFF \sreg_reg[248]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(c[248]) );
  DFF \sreg_reg[247]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(c[247]) );
  DFF \sreg_reg[246]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(c[246]) );
  DFF \sreg_reg[245]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(c[245]) );
  DFF \sreg_reg[244]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(c[244]) );
  DFF \sreg_reg[243]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(c[243]) );
  DFF \sreg_reg[242]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(c[242]) );
  DFF \sreg_reg[241]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(c[241]) );
  DFF \sreg_reg[240]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(c[240]) );
  DFF \sreg_reg[239]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(c[239]) );
  DFF \sreg_reg[238]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(c[238]) );
  DFF \sreg_reg[237]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(c[237]) );
  DFF \sreg_reg[236]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(c[236]) );
  DFF \sreg_reg[235]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(c[235]) );
  DFF \sreg_reg[234]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(c[234]) );
  DFF \sreg_reg[233]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(c[233]) );
  DFF \sreg_reg[232]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(c[232]) );
  DFF \sreg_reg[231]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(c[231]) );
  DFF \sreg_reg[230]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(c[230]) );
  DFF \sreg_reg[229]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(c[229]) );
  DFF \sreg_reg[228]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(c[228]) );
  DFF \sreg_reg[227]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(c[227]) );
  DFF \sreg_reg[226]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(c[226]) );
  DFF \sreg_reg[225]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(c[225]) );
  DFF \sreg_reg[224]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(c[224]) );
  DFF \sreg_reg[223]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(c[223]) );
  DFF \sreg_reg[222]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(c[222]) );
  DFF \sreg_reg[221]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(c[221]) );
  DFF \sreg_reg[220]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(c[220]) );
  DFF \sreg_reg[219]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(c[219]) );
  DFF \sreg_reg[218]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(c[218]) );
  DFF \sreg_reg[217]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(c[217]) );
  DFF \sreg_reg[216]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(c[216]) );
  DFF \sreg_reg[215]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(c[215]) );
  DFF \sreg_reg[214]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(c[214]) );
  DFF \sreg_reg[213]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(c[213]) );
  DFF \sreg_reg[212]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(c[212]) );
  DFF \sreg_reg[211]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(c[211]) );
  DFF \sreg_reg[210]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(c[210]) );
  DFF \sreg_reg[209]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(c[209]) );
  DFF \sreg_reg[208]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(c[208]) );
  DFF \sreg_reg[207]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(c[207]) );
  DFF \sreg_reg[206]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(c[206]) );
  DFF \sreg_reg[205]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(c[205]) );
  DFF \sreg_reg[204]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(c[204]) );
  DFF \sreg_reg[203]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(c[203]) );
  DFF \sreg_reg[202]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(c[202]) );
  DFF \sreg_reg[201]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(c[201]) );
  DFF \sreg_reg[200]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(c[200]) );
  DFF \sreg_reg[199]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(c[199]) );
  DFF \sreg_reg[198]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(c[198]) );
  DFF \sreg_reg[197]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(c[197]) );
  DFF \sreg_reg[196]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(c[196]) );
  DFF \sreg_reg[195]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(c[195]) );
  DFF \sreg_reg[194]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(c[194]) );
  DFF \sreg_reg[193]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(c[193]) );
  DFF \sreg_reg[192]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(c[192]) );
  DFF \sreg_reg[191]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(c[191]) );
  DFF \sreg_reg[190]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(c[190]) );
  DFF \sreg_reg[189]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(c[189]) );
  DFF \sreg_reg[188]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(c[188]) );
  DFF \sreg_reg[187]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(c[187]) );
  DFF \sreg_reg[186]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(c[186]) );
  DFF \sreg_reg[185]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(c[185]) );
  DFF \sreg_reg[184]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(c[184]) );
  DFF \sreg_reg[183]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(c[183]) );
  DFF \sreg_reg[182]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(c[182]) );
  DFF \sreg_reg[181]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(c[181]) );
  DFF \sreg_reg[180]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(c[180]) );
  DFF \sreg_reg[179]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(c[179]) );
  DFF \sreg_reg[178]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(c[178]) );
  DFF \sreg_reg[177]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(c[177]) );
  DFF \sreg_reg[176]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(c[176]) );
  DFF \sreg_reg[175]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(c[175]) );
  DFF \sreg_reg[174]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(c[174]) );
  DFF \sreg_reg[173]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(c[173]) );
  DFF \sreg_reg[172]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(c[172]) );
  DFF \sreg_reg[171]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(c[171]) );
  DFF \sreg_reg[170]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(c[170]) );
  DFF \sreg_reg[169]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(c[169]) );
  DFF \sreg_reg[168]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(c[168]) );
  DFF \sreg_reg[167]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(c[167]) );
  DFF \sreg_reg[166]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(c[166]) );
  DFF \sreg_reg[165]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(c[165]) );
  DFF \sreg_reg[164]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(c[164]) );
  DFF \sreg_reg[163]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(c[163]) );
  DFF \sreg_reg[162]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(c[162]) );
  DFF \sreg_reg[161]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(c[161]) );
  DFF \sreg_reg[160]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(c[160]) );
  DFF \sreg_reg[159]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(c[159]) );
  DFF \sreg_reg[158]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(c[158]) );
  DFF \sreg_reg[157]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(c[157]) );
  DFF \sreg_reg[156]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(c[156]) );
  DFF \sreg_reg[155]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(c[155]) );
  DFF \sreg_reg[154]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(c[154]) );
  DFF \sreg_reg[153]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(c[153]) );
  DFF \sreg_reg[152]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(c[152]) );
  DFF \sreg_reg[151]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(c[151]) );
  DFF \sreg_reg[150]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(c[150]) );
  DFF \sreg_reg[149]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(c[149]) );
  DFF \sreg_reg[148]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(c[148]) );
  DFF \sreg_reg[147]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(c[147]) );
  DFF \sreg_reg[146]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(c[146]) );
  DFF \sreg_reg[145]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(c[145]) );
  DFF \sreg_reg[144]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(c[144]) );
  DFF \sreg_reg[143]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(c[143]) );
  DFF \sreg_reg[142]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(c[142]) );
  DFF \sreg_reg[141]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(c[141]) );
  DFF \sreg_reg[140]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(c[140]) );
  DFF \sreg_reg[139]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(c[139]) );
  DFF \sreg_reg[138]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(c[138]) );
  DFF \sreg_reg[137]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(c[137]) );
  DFF \sreg_reg[136]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(c[136]) );
  DFF \sreg_reg[135]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(c[135]) );
  DFF \sreg_reg[134]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(c[134]) );
  DFF \sreg_reg[133]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(c[133]) );
  DFF \sreg_reg[132]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(c[132]) );
  DFF \sreg_reg[131]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(c[131]) );
  DFF \sreg_reg[130]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(c[130]) );
  DFF \sreg_reg[129]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(c[129]) );
  DFF \sreg_reg[128]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(c[128]) );
  DFF \sreg_reg[127]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(c[127]) );
  DFF \sreg_reg[126]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(c[126]) );
  DFF \sreg_reg[125]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[125]) );
  DFF \sreg_reg[124]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[124]) );
  DFF \sreg_reg[123]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[123]) );
  DFF \sreg_reg[122]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[122]) );
  DFF \sreg_reg[121]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[121]) );
  DFF \sreg_reg[120]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[120]) );
  DFF \sreg_reg[119]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[118]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[117]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[116]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[115]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[114]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[113]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[112]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[111]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[110]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[109]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[108]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[107]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[106]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[105]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[104]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[103]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[102]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[101]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[100]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[99]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[98]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[97]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[96]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[95]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[94]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[93]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[92]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[91]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[90]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[89]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[88]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[87]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[86]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[85]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[84]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[83]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[82]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[81]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[80]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[79]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[78]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[77]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[76]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[75]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[74]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[73]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[72]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[71]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[70]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[69]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[68]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[67]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[66]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[65]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[64]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[63]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[62]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[3]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[2]), .CLK(clk), .RST(rst), .Q(c[0]) );
  NANDN U5 ( .A(n1321), .B(n1322), .Z(n1) );
  NANDN U6 ( .A(n1324), .B(n1323), .Z(n2) );
  NAND U7 ( .A(n1), .B(n2), .Z(n1330) );
  NANDN U8 ( .A(n1342), .B(n1343), .Z(n3) );
  NANDN U9 ( .A(n1345), .B(n1344), .Z(n4) );
  NAND U10 ( .A(n3), .B(n4), .Z(n1351) );
  NANDN U11 ( .A(n1363), .B(n1364), .Z(n5) );
  NANDN U12 ( .A(n1366), .B(n1365), .Z(n6) );
  AND U13 ( .A(n5), .B(n6), .Z(n1372) );
  NANDN U14 ( .A(n1386), .B(n1387), .Z(n7) );
  NANDN U15 ( .A(n1384), .B(n1385), .Z(n8) );
  NAND U16 ( .A(n7), .B(n8), .Z(n1393) );
  NANDN U17 ( .A(n1407), .B(n1408), .Z(n9) );
  NANDN U18 ( .A(n1405), .B(n1406), .Z(n10) );
  NAND U19 ( .A(n9), .B(n10), .Z(n1414) );
  NANDN U20 ( .A(n1426), .B(n1427), .Z(n11) );
  NANDN U21 ( .A(n1429), .B(n1428), .Z(n12) );
  AND U22 ( .A(n11), .B(n12), .Z(n1435) );
  NANDN U23 ( .A(n1447), .B(n1448), .Z(n13) );
  NANDN U24 ( .A(n1450), .B(n1449), .Z(n14) );
  NAND U25 ( .A(n13), .B(n14), .Z(n1456) );
  NANDN U26 ( .A(n1470), .B(n1471), .Z(n15) );
  NANDN U27 ( .A(n1468), .B(n1469), .Z(n16) );
  NAND U28 ( .A(n15), .B(n16), .Z(n1477) );
  NANDN U29 ( .A(n1489), .B(n1490), .Z(n17) );
  NANDN U30 ( .A(n1492), .B(n1491), .Z(n18) );
  AND U31 ( .A(n17), .B(n18), .Z(n1498) );
  NANDN U32 ( .A(n1510), .B(n1511), .Z(n19) );
  NANDN U33 ( .A(n1512), .B(n1513), .Z(n20) );
  AND U34 ( .A(n19), .B(n20), .Z(n1519) );
  NANDN U35 ( .A(n1531), .B(n1532), .Z(n21) );
  NANDN U36 ( .A(n1534), .B(n1533), .Z(n22) );
  NAND U37 ( .A(n21), .B(n22), .Z(n1540) );
  NANDN U38 ( .A(n1554), .B(n1555), .Z(n23) );
  NANDN U39 ( .A(n1552), .B(n1553), .Z(n24) );
  NAND U40 ( .A(n23), .B(n24), .Z(n1561) );
  NANDN U41 ( .A(n1573), .B(n1574), .Z(n25) );
  NANDN U42 ( .A(n1576), .B(n1575), .Z(n26) );
  AND U43 ( .A(n25), .B(n26), .Z(n1582) );
  NANDN U44 ( .A(n1596), .B(n1597), .Z(n27) );
  NANDN U45 ( .A(n1594), .B(n1595), .Z(n28) );
  NAND U46 ( .A(n27), .B(n28), .Z(n1603) );
  NANDN U47 ( .A(n1615), .B(n1616), .Z(n29) );
  NANDN U48 ( .A(n1618), .B(n1617), .Z(n30) );
  NAND U49 ( .A(n29), .B(n30), .Z(n1624) );
  NANDN U50 ( .A(n1636), .B(n1637), .Z(n31) );
  NANDN U51 ( .A(n1639), .B(n1638), .Z(n32) );
  AND U52 ( .A(n31), .B(n32), .Z(n1645) );
  NANDN U53 ( .A(n1657), .B(n1658), .Z(n33) );
  NANDN U54 ( .A(n1659), .B(n1660), .Z(n34) );
  AND U55 ( .A(n33), .B(n34), .Z(n1666) );
  NANDN U56 ( .A(n1678), .B(n1679), .Z(n35) );
  NANDN U57 ( .A(n1681), .B(n1680), .Z(n36) );
  NAND U58 ( .A(n35), .B(n36), .Z(n1687) );
  NANDN U59 ( .A(n1699), .B(n1700), .Z(n37) );
  NANDN U60 ( .A(n1702), .B(n1701), .Z(n38) );
  AND U61 ( .A(n37), .B(n38), .Z(n1708) );
  NANDN U62 ( .A(n1722), .B(n1723), .Z(n39) );
  NANDN U63 ( .A(n1720), .B(n1721), .Z(n40) );
  NAND U64 ( .A(n39), .B(n40), .Z(n1729) );
  NANDN U65 ( .A(n1741), .B(n1742), .Z(n41) );
  NANDN U66 ( .A(n1744), .B(n1743), .Z(n42) );
  NAND U67 ( .A(n41), .B(n42), .Z(n1750) );
  NANDN U68 ( .A(n1764), .B(n1765), .Z(n43) );
  NANDN U69 ( .A(n1762), .B(n1763), .Z(n44) );
  NAND U70 ( .A(n43), .B(n44), .Z(n1771) );
  NANDN U71 ( .A(n1783), .B(n1784), .Z(n45) );
  NANDN U72 ( .A(n1786), .B(n1785), .Z(n46) );
  NAND U73 ( .A(n45), .B(n46), .Z(n1792) );
  NANDN U74 ( .A(n1804), .B(n1805), .Z(n47) );
  NANDN U75 ( .A(n1807), .B(n1806), .Z(n48) );
  NAND U76 ( .A(n47), .B(n48), .Z(n1813) );
  NANDN U77 ( .A(n1825), .B(n1826), .Z(n49) );
  NANDN U78 ( .A(n1828), .B(n1827), .Z(n50) );
  NAND U79 ( .A(n49), .B(n50), .Z(n1834) );
  NANDN U80 ( .A(n1846), .B(n1847), .Z(n51) );
  NANDN U81 ( .A(n1849), .B(n1848), .Z(n52) );
  AND U82 ( .A(n51), .B(n52), .Z(n1855) );
  NANDN U83 ( .A(n1869), .B(n1870), .Z(n53) );
  NANDN U84 ( .A(n1867), .B(n1868), .Z(n54) );
  NAND U85 ( .A(n53), .B(n54), .Z(n1876) );
  NANDN U86 ( .A(n1888), .B(n1889), .Z(n55) );
  NANDN U87 ( .A(n1891), .B(n1890), .Z(n56) );
  NAND U88 ( .A(n55), .B(n56), .Z(n1897) );
  NANDN U89 ( .A(n1909), .B(n1910), .Z(n57) );
  NANDN U90 ( .A(n1912), .B(n1911), .Z(n58) );
  AND U91 ( .A(n57), .B(n58), .Z(n1918) );
  NANDN U92 ( .A(n1932), .B(n1933), .Z(n59) );
  NANDN U93 ( .A(n1930), .B(n1931), .Z(n60) );
  NAND U94 ( .A(n59), .B(n60), .Z(n1939) );
  NANDN U95 ( .A(n1951), .B(n1952), .Z(n61) );
  NANDN U96 ( .A(n1954), .B(n1953), .Z(n62) );
  AND U97 ( .A(n61), .B(n62), .Z(n1960) );
  NANDN U98 ( .A(n1972), .B(n1973), .Z(n63) );
  NANDN U99 ( .A(n1975), .B(n1974), .Z(n64) );
  NAND U100 ( .A(n63), .B(n64), .Z(n1981) );
  NANDN U101 ( .A(n1993), .B(n1994), .Z(n65) );
  NANDN U102 ( .A(n1995), .B(n1996), .Z(n66) );
  AND U103 ( .A(n65), .B(n66), .Z(n2002) );
  NANDN U104 ( .A(n2014), .B(n2015), .Z(n67) );
  NANDN U105 ( .A(n2017), .B(n2016), .Z(n68) );
  NAND U106 ( .A(n67), .B(n68), .Z(n2023) );
  NANDN U107 ( .A(n2035), .B(n2036), .Z(n69) );
  NANDN U108 ( .A(n2038), .B(n2037), .Z(n70) );
  AND U109 ( .A(n69), .B(n70), .Z(n2044) );
  NANDN U110 ( .A(n2056), .B(n2057), .Z(n71) );
  NANDN U111 ( .A(n2059), .B(n2058), .Z(n72) );
  NAND U112 ( .A(n71), .B(n72), .Z(n2065) );
  NANDN U113 ( .A(n2079), .B(n2080), .Z(n73) );
  NANDN U114 ( .A(n2077), .B(n2078), .Z(n74) );
  NAND U115 ( .A(n73), .B(n74), .Z(n2086) );
  NANDN U116 ( .A(n2098), .B(n2099), .Z(n75) );
  NANDN U117 ( .A(n2101), .B(n2100), .Z(n76) );
  AND U118 ( .A(n75), .B(n76), .Z(n2107) );
  NANDN U119 ( .A(n2119), .B(n2120), .Z(n77) );
  NANDN U120 ( .A(n2122), .B(n2121), .Z(n78) );
  NAND U121 ( .A(n77), .B(n78), .Z(n2128) );
  NANDN U122 ( .A(n2142), .B(n2143), .Z(n79) );
  NANDN U123 ( .A(n2140), .B(n2141), .Z(n80) );
  NAND U124 ( .A(n79), .B(n80), .Z(n2149) );
  NANDN U125 ( .A(n2161), .B(n2162), .Z(n81) );
  NANDN U126 ( .A(n2164), .B(n2163), .Z(n82) );
  AND U127 ( .A(n81), .B(n82), .Z(n2170) );
  NANDN U128 ( .A(n2184), .B(n2185), .Z(n83) );
  NANDN U129 ( .A(n2182), .B(n2183), .Z(n84) );
  NAND U130 ( .A(n83), .B(n84), .Z(n2191) );
  NANDN U131 ( .A(n2203), .B(n2204), .Z(n85) );
  NANDN U132 ( .A(n2206), .B(n2205), .Z(n86) );
  NAND U133 ( .A(n85), .B(n86), .Z(n2212) );
  NANDN U134 ( .A(n2226), .B(n2227), .Z(n87) );
  NANDN U135 ( .A(n2224), .B(n2225), .Z(n88) );
  NAND U136 ( .A(n87), .B(n88), .Z(n2233) );
  NANDN U137 ( .A(n2245), .B(n2246), .Z(n89) );
  NANDN U138 ( .A(n2248), .B(n2247), .Z(n90) );
  AND U139 ( .A(n89), .B(n90), .Z(n2254) );
  NANDN U140 ( .A(n2268), .B(n2269), .Z(n91) );
  NANDN U141 ( .A(n2266), .B(n2267), .Z(n92) );
  NAND U142 ( .A(n91), .B(n92), .Z(n2275) );
  NANDN U143 ( .A(n2287), .B(n2288), .Z(n93) );
  NANDN U144 ( .A(n2290), .B(n2289), .Z(n94) );
  NAND U145 ( .A(n93), .B(n94), .Z(n2296) );
  NANDN U146 ( .A(n2308), .B(n2309), .Z(n95) );
  NANDN U147 ( .A(n2311), .B(n2310), .Z(n96) );
  AND U148 ( .A(n95), .B(n96), .Z(n2317) );
  NANDN U149 ( .A(n2331), .B(n2332), .Z(n97) );
  NANDN U150 ( .A(n2329), .B(n2330), .Z(n98) );
  NAND U151 ( .A(n97), .B(n98), .Z(n2338) );
  NANDN U152 ( .A(n2350), .B(n2351), .Z(n99) );
  NANDN U153 ( .A(n2353), .B(n2352), .Z(n100) );
  NAND U154 ( .A(n99), .B(n100), .Z(n2359) );
  NANDN U155 ( .A(n2371), .B(n2372), .Z(n101) );
  NANDN U156 ( .A(n2374), .B(n2373), .Z(n102) );
  AND U157 ( .A(n101), .B(n102), .Z(n2380) );
  NANDN U158 ( .A(n2394), .B(n2395), .Z(n103) );
  NANDN U159 ( .A(n2392), .B(n2393), .Z(n104) );
  NAND U160 ( .A(n103), .B(n104), .Z(n2401) );
  NANDN U161 ( .A(n2413), .B(n2414), .Z(n105) );
  NANDN U162 ( .A(n2416), .B(n2415), .Z(n106) );
  AND U163 ( .A(n105), .B(n106), .Z(n2422) );
  NANDN U164 ( .A(n2434), .B(n2435), .Z(n107) );
  NANDN U165 ( .A(n2437), .B(n2436), .Z(n108) );
  NAND U166 ( .A(n107), .B(n108), .Z(n2443) );
  NANDN U167 ( .A(n2455), .B(n2456), .Z(n109) );
  NANDN U168 ( .A(n2458), .B(n2457), .Z(n110) );
  NAND U169 ( .A(n109), .B(n110), .Z(n2464) );
  NANDN U170 ( .A(n2476), .B(n2477), .Z(n111) );
  NANDN U171 ( .A(n2478), .B(n2479), .Z(n112) );
  AND U172 ( .A(n111), .B(n112), .Z(n2485) );
  NANDN U173 ( .A(n2497), .B(n2498), .Z(n113) );
  NANDN U174 ( .A(n2500), .B(n2499), .Z(n114) );
  NAND U175 ( .A(n113), .B(n114), .Z(n2506) );
  NANDN U176 ( .A(n2518), .B(n2519), .Z(n115) );
  NANDN U177 ( .A(n2521), .B(n2520), .Z(n116) );
  AND U178 ( .A(n115), .B(n116), .Z(n2527) );
  NANDN U179 ( .A(n2541), .B(n2542), .Z(n117) );
  NANDN U180 ( .A(n2539), .B(n2540), .Z(n118) );
  NAND U181 ( .A(n117), .B(n118), .Z(n2548) );
  NANDN U182 ( .A(n2560), .B(n2561), .Z(n119) );
  NANDN U183 ( .A(n2563), .B(n2562), .Z(n120) );
  AND U184 ( .A(n119), .B(n120), .Z(n2569) );
  NANDN U185 ( .A(n2581), .B(n2582), .Z(n121) );
  NANDN U186 ( .A(n2584), .B(n2583), .Z(n122) );
  AND U187 ( .A(n121), .B(n122), .Z(n2590) );
  NANDN U188 ( .A(n2604), .B(n2605), .Z(n123) );
  NANDN U189 ( .A(n2602), .B(n2603), .Z(n124) );
  NAND U190 ( .A(n123), .B(n124), .Z(n2611) );
  NANDN U191 ( .A(n2623), .B(n2624), .Z(n125) );
  NANDN U192 ( .A(n2626), .B(n2625), .Z(n126) );
  AND U193 ( .A(n125), .B(n126), .Z(n2632) );
  NANDN U194 ( .A(n2644), .B(n2645), .Z(n127) );
  NANDN U195 ( .A(n2647), .B(n2646), .Z(n128) );
  NAND U196 ( .A(n127), .B(n128), .Z(n2653) );
  NANDN U197 ( .A(n2665), .B(n2666), .Z(n129) );
  NANDN U198 ( .A(n2668), .B(n2667), .Z(n130) );
  AND U199 ( .A(n129), .B(n130), .Z(n2674) );
  NANDN U200 ( .A(n2686), .B(n2687), .Z(n131) );
  NANDN U201 ( .A(n2689), .B(n2688), .Z(n132) );
  NAND U202 ( .A(n131), .B(n132), .Z(n2695) );
  NANDN U203 ( .A(n2707), .B(n2708), .Z(n133) );
  NANDN U204 ( .A(n2710), .B(n2709), .Z(n134) );
  AND U205 ( .A(n133), .B(n134), .Z(n2716) );
  NANDN U206 ( .A(n2728), .B(n2729), .Z(n135) );
  NANDN U207 ( .A(n2731), .B(n2730), .Z(n136) );
  NAND U208 ( .A(n135), .B(n136), .Z(n2737) );
  NANDN U209 ( .A(n2751), .B(n2752), .Z(n137) );
  NANDN U210 ( .A(n2749), .B(n2750), .Z(n138) );
  NAND U211 ( .A(n137), .B(n138), .Z(n2758) );
  NANDN U212 ( .A(n2770), .B(n2771), .Z(n139) );
  NANDN U213 ( .A(n2773), .B(n2772), .Z(n140) );
  NAND U214 ( .A(n139), .B(n140), .Z(n2779) );
  NANDN U215 ( .A(n2791), .B(n2792), .Z(n141) );
  NANDN U216 ( .A(n2794), .B(n2793), .Z(n142) );
  NAND U217 ( .A(n141), .B(n142), .Z(n2800) );
  NANDN U218 ( .A(n2812), .B(n2813), .Z(n143) );
  NANDN U219 ( .A(n2814), .B(n2815), .Z(n144) );
  AND U220 ( .A(n143), .B(n144), .Z(n2821) );
  NANDN U221 ( .A(n2833), .B(n2834), .Z(n145) );
  NANDN U222 ( .A(n2836), .B(n2835), .Z(n146) );
  AND U223 ( .A(n145), .B(n146), .Z(n2842) );
  NANDN U224 ( .A(n2854), .B(n2855), .Z(n147) );
  NANDN U225 ( .A(n2857), .B(n2856), .Z(n148) );
  AND U226 ( .A(n147), .B(n148), .Z(n2863) );
  NANDN U227 ( .A(n2875), .B(n2876), .Z(n149) );
  NANDN U228 ( .A(n2878), .B(n2877), .Z(n150) );
  AND U229 ( .A(n149), .B(n150), .Z(n2884) );
  NANDN U230 ( .A(n2898), .B(n2899), .Z(n151) );
  NANDN U231 ( .A(n2896), .B(n2897), .Z(n152) );
  NAND U232 ( .A(n151), .B(n152), .Z(n2905) );
  NANDN U233 ( .A(n2917), .B(n2918), .Z(n153) );
  NANDN U234 ( .A(n2920), .B(n2919), .Z(n154) );
  NAND U235 ( .A(n153), .B(n154), .Z(n2926) );
  NANDN U236 ( .A(n2940), .B(n2941), .Z(n155) );
  NANDN U237 ( .A(n2938), .B(n2939), .Z(n156) );
  NAND U238 ( .A(n155), .B(n156), .Z(n2947) );
  NANDN U239 ( .A(n2959), .B(n2960), .Z(n157) );
  NANDN U240 ( .A(n2962), .B(n2961), .Z(n158) );
  NAND U241 ( .A(n157), .B(n158), .Z(n2968) );
  NANDN U242 ( .A(n2980), .B(n2981), .Z(n159) );
  NANDN U243 ( .A(n2983), .B(n2982), .Z(n160) );
  AND U244 ( .A(n159), .B(n160), .Z(n2989) );
  NANDN U245 ( .A(n3003), .B(n3004), .Z(n161) );
  NANDN U246 ( .A(n3001), .B(n3002), .Z(n162) );
  NAND U247 ( .A(n161), .B(n162), .Z(n3010) );
  NANDN U248 ( .A(n3022), .B(n3023), .Z(n163) );
  NANDN U249 ( .A(n3025), .B(n3024), .Z(n164) );
  NAND U250 ( .A(n163), .B(n164), .Z(n3031) );
  NANDN U251 ( .A(n1328), .B(n1329), .Z(n165) );
  NANDN U252 ( .A(n1331), .B(n1330), .Z(n166) );
  AND U253 ( .A(n165), .B(n166), .Z(n1337) );
  NANDN U254 ( .A(n1349), .B(n1350), .Z(n167) );
  NANDN U255 ( .A(n1352), .B(n1351), .Z(n168) );
  AND U256 ( .A(n167), .B(n168), .Z(n1358) );
  NANDN U257 ( .A(n1370), .B(n1371), .Z(n169) );
  NANDN U258 ( .A(n1372), .B(n1373), .Z(n170) );
  AND U259 ( .A(n169), .B(n170), .Z(n1379) );
  NANDN U260 ( .A(n1391), .B(n1392), .Z(n171) );
  NANDN U261 ( .A(n1394), .B(n1393), .Z(n172) );
  NAND U262 ( .A(n171), .B(n172), .Z(n1400) );
  NANDN U263 ( .A(n1412), .B(n1413), .Z(n173) );
  NANDN U264 ( .A(n1415), .B(n1414), .Z(n174) );
  AND U265 ( .A(n173), .B(n174), .Z(n1421) );
  NANDN U266 ( .A(n1435), .B(n1436), .Z(n175) );
  NANDN U267 ( .A(n1433), .B(n1434), .Z(n176) );
  NAND U268 ( .A(n175), .B(n176), .Z(n1442) );
  NANDN U269 ( .A(n1454), .B(n1455), .Z(n177) );
  NANDN U270 ( .A(n1457), .B(n1456), .Z(n178) );
  NAND U271 ( .A(n177), .B(n178), .Z(n1463) );
  NANDN U272 ( .A(n1475), .B(n1476), .Z(n179) );
  NANDN U273 ( .A(n1478), .B(n1477), .Z(n180) );
  AND U274 ( .A(n179), .B(n180), .Z(n1484) );
  NANDN U275 ( .A(n1498), .B(n1499), .Z(n181) );
  NANDN U276 ( .A(n1496), .B(n1497), .Z(n182) );
  NAND U277 ( .A(n181), .B(n182), .Z(n1505) );
  NANDN U278 ( .A(n1519), .B(n1520), .Z(n183) );
  NANDN U279 ( .A(n1517), .B(n1518), .Z(n184) );
  NAND U280 ( .A(n183), .B(n184), .Z(n1526) );
  NANDN U281 ( .A(n1538), .B(n1539), .Z(n185) );
  NANDN U282 ( .A(n1541), .B(n1540), .Z(n186) );
  NAND U283 ( .A(n185), .B(n186), .Z(n1547) );
  NANDN U284 ( .A(n1559), .B(n1560), .Z(n187) );
  NANDN U285 ( .A(n1562), .B(n1561), .Z(n188) );
  NAND U286 ( .A(n187), .B(n188), .Z(n1568) );
  NANDN U287 ( .A(n1582), .B(n1583), .Z(n189) );
  NANDN U288 ( .A(n1580), .B(n1581), .Z(n190) );
  NAND U289 ( .A(n189), .B(n190), .Z(n1589) );
  NANDN U290 ( .A(n1601), .B(n1602), .Z(n191) );
  NANDN U291 ( .A(n1604), .B(n1603), .Z(n192) );
  NAND U292 ( .A(n191), .B(n192), .Z(n1610) );
  NANDN U293 ( .A(n1622), .B(n1623), .Z(n193) );
  NANDN U294 ( .A(n1625), .B(n1624), .Z(n194) );
  AND U295 ( .A(n193), .B(n194), .Z(n1631) );
  NANDN U296 ( .A(n1645), .B(n1646), .Z(n195) );
  NANDN U297 ( .A(n1643), .B(n1644), .Z(n196) );
  NAND U298 ( .A(n195), .B(n196), .Z(n1652) );
  NANDN U299 ( .A(n1664), .B(n1665), .Z(n197) );
  NANDN U300 ( .A(n1666), .B(n1667), .Z(n198) );
  AND U301 ( .A(n197), .B(n198), .Z(n1673) );
  NANDN U302 ( .A(n1685), .B(n1686), .Z(n199) );
  NANDN U303 ( .A(n1688), .B(n1687), .Z(n200) );
  NAND U304 ( .A(n199), .B(n200), .Z(n1694) );
  NANDN U305 ( .A(n1708), .B(n1709), .Z(n201) );
  NANDN U306 ( .A(n1706), .B(n1707), .Z(n202) );
  NAND U307 ( .A(n201), .B(n202), .Z(n1715) );
  NANDN U308 ( .A(n1727), .B(n1728), .Z(n203) );
  NANDN U309 ( .A(n1730), .B(n1729), .Z(n204) );
  AND U310 ( .A(n203), .B(n204), .Z(n1736) );
  NANDN U311 ( .A(n1748), .B(n1749), .Z(n205) );
  NANDN U312 ( .A(n1751), .B(n1750), .Z(n206) );
  NAND U313 ( .A(n205), .B(n206), .Z(n1757) );
  NANDN U314 ( .A(n1769), .B(n1770), .Z(n207) );
  NANDN U315 ( .A(n1772), .B(n1771), .Z(n208) );
  NAND U316 ( .A(n207), .B(n208), .Z(n1778) );
  NANDN U317 ( .A(n1790), .B(n1791), .Z(n209) );
  NANDN U318 ( .A(n1793), .B(n1792), .Z(n210) );
  NAND U319 ( .A(n209), .B(n210), .Z(n1799) );
  NANDN U320 ( .A(n1811), .B(n1812), .Z(n211) );
  NANDN U321 ( .A(n1814), .B(n1813), .Z(n212) );
  AND U322 ( .A(n211), .B(n212), .Z(n1820) );
  NANDN U323 ( .A(n1832), .B(n1833), .Z(n213) );
  NANDN U324 ( .A(n1835), .B(n1834), .Z(n214) );
  NAND U325 ( .A(n213), .B(n214), .Z(n1841) );
  NANDN U326 ( .A(n1855), .B(n1856), .Z(n215) );
  NANDN U327 ( .A(n1853), .B(n1854), .Z(n216) );
  NAND U328 ( .A(n215), .B(n216), .Z(n1862) );
  NANDN U329 ( .A(n1874), .B(n1875), .Z(n217) );
  NANDN U330 ( .A(n1877), .B(n1876), .Z(n218) );
  AND U331 ( .A(n217), .B(n218), .Z(n1883) );
  NANDN U332 ( .A(n1895), .B(n1896), .Z(n219) );
  NANDN U333 ( .A(n1898), .B(n1897), .Z(n220) );
  NAND U334 ( .A(n219), .B(n220), .Z(n1904) );
  NANDN U335 ( .A(n1918), .B(n1919), .Z(n221) );
  NANDN U336 ( .A(n1916), .B(n1917), .Z(n222) );
  NAND U337 ( .A(n221), .B(n222), .Z(n1925) );
  NANDN U338 ( .A(n1937), .B(n1938), .Z(n223) );
  NANDN U339 ( .A(n1940), .B(n1939), .Z(n224) );
  AND U340 ( .A(n223), .B(n224), .Z(n1946) );
  NANDN U341 ( .A(n1960), .B(n1961), .Z(n225) );
  NANDN U342 ( .A(n1958), .B(n1959), .Z(n226) );
  NAND U343 ( .A(n225), .B(n226), .Z(n1967) );
  NANDN U344 ( .A(n1979), .B(n1980), .Z(n227) );
  NANDN U345 ( .A(n1982), .B(n1981), .Z(n228) );
  NAND U346 ( .A(n227), .B(n228), .Z(n1988) );
  NANDN U347 ( .A(n2002), .B(n2003), .Z(n229) );
  NANDN U348 ( .A(n2000), .B(n2001), .Z(n230) );
  NAND U349 ( .A(n229), .B(n230), .Z(n2009) );
  NANDN U350 ( .A(n2021), .B(n2022), .Z(n231) );
  NANDN U351 ( .A(n2024), .B(n2023), .Z(n232) );
  AND U352 ( .A(n231), .B(n232), .Z(n2030) );
  NANDN U353 ( .A(n2042), .B(n2043), .Z(n233) );
  NANDN U354 ( .A(n2044), .B(n2045), .Z(n234) );
  AND U355 ( .A(n233), .B(n234), .Z(n2051) );
  NANDN U356 ( .A(n2063), .B(n2064), .Z(n235) );
  NANDN U357 ( .A(n2066), .B(n2065), .Z(n236) );
  NAND U358 ( .A(n235), .B(n236), .Z(n2072) );
  NANDN U359 ( .A(n2084), .B(n2085), .Z(n237) );
  NANDN U360 ( .A(n2087), .B(n2086), .Z(n238) );
  NAND U361 ( .A(n237), .B(n238), .Z(n2093) );
  NANDN U362 ( .A(n2107), .B(n2108), .Z(n239) );
  NANDN U363 ( .A(n2105), .B(n2106), .Z(n240) );
  NAND U364 ( .A(n239), .B(n240), .Z(n2114) );
  NANDN U365 ( .A(n2126), .B(n2127), .Z(n241) );
  NANDN U366 ( .A(n2129), .B(n2128), .Z(n242) );
  NAND U367 ( .A(n241), .B(n242), .Z(n2135) );
  NANDN U368 ( .A(n2147), .B(n2148), .Z(n243) );
  NANDN U369 ( .A(n2150), .B(n2149), .Z(n244) );
  AND U370 ( .A(n243), .B(n244), .Z(n2156) );
  NANDN U371 ( .A(n2170), .B(n2171), .Z(n245) );
  NANDN U372 ( .A(n2168), .B(n2169), .Z(n246) );
  NAND U373 ( .A(n245), .B(n246), .Z(n2177) );
  NANDN U374 ( .A(n2189), .B(n2190), .Z(n247) );
  NANDN U375 ( .A(n2192), .B(n2191), .Z(n248) );
  AND U376 ( .A(n247), .B(n248), .Z(n2198) );
  NANDN U377 ( .A(n2210), .B(n2211), .Z(n249) );
  NANDN U378 ( .A(n2213), .B(n2212), .Z(n250) );
  NAND U379 ( .A(n249), .B(n250), .Z(n2219) );
  NANDN U380 ( .A(n2231), .B(n2232), .Z(n251) );
  NANDN U381 ( .A(n2234), .B(n2233), .Z(n252) );
  NAND U382 ( .A(n251), .B(n252), .Z(n2240) );
  NANDN U383 ( .A(n2254), .B(n2255), .Z(n253) );
  NANDN U384 ( .A(n2252), .B(n2253), .Z(n254) );
  NAND U385 ( .A(n253), .B(n254), .Z(n2261) );
  NANDN U386 ( .A(n2273), .B(n2274), .Z(n255) );
  NANDN U387 ( .A(n2276), .B(n2275), .Z(n256) );
  AND U388 ( .A(n255), .B(n256), .Z(n2282) );
  NANDN U389 ( .A(n2294), .B(n2295), .Z(n257) );
  NANDN U390 ( .A(n2297), .B(n2296), .Z(n258) );
  AND U391 ( .A(n257), .B(n258), .Z(n2303) );
  NANDN U392 ( .A(n2315), .B(n2316), .Z(n259) );
  NANDN U393 ( .A(n2317), .B(n2318), .Z(n260) );
  AND U394 ( .A(n259), .B(n260), .Z(n2324) );
  NANDN U395 ( .A(n2336), .B(n2337), .Z(n261) );
  NANDN U396 ( .A(n2339), .B(n2338), .Z(n262) );
  NAND U397 ( .A(n261), .B(n262), .Z(n2345) );
  NANDN U398 ( .A(n2357), .B(n2358), .Z(n263) );
  NANDN U399 ( .A(n2360), .B(n2359), .Z(n264) );
  NAND U400 ( .A(n263), .B(n264), .Z(n2366) );
  NANDN U401 ( .A(n2380), .B(n2381), .Z(n265) );
  NANDN U402 ( .A(n2378), .B(n2379), .Z(n266) );
  NAND U403 ( .A(n265), .B(n266), .Z(n2387) );
  NANDN U404 ( .A(n2399), .B(n2400), .Z(n267) );
  NANDN U405 ( .A(n2402), .B(n2401), .Z(n268) );
  AND U406 ( .A(n267), .B(n268), .Z(n2408) );
  NANDN U407 ( .A(n2422), .B(n2423), .Z(n269) );
  NANDN U408 ( .A(n2420), .B(n2421), .Z(n270) );
  NAND U409 ( .A(n269), .B(n270), .Z(n2429) );
  NANDN U410 ( .A(n2441), .B(n2442), .Z(n271) );
  NANDN U411 ( .A(n2444), .B(n2443), .Z(n272) );
  NAND U412 ( .A(n271), .B(n272), .Z(n2450) );
  NANDN U413 ( .A(n2462), .B(n2463), .Z(n273) );
  NANDN U414 ( .A(n2465), .B(n2464), .Z(n274) );
  NAND U415 ( .A(n273), .B(n274), .Z(n2471) );
  NANDN U416 ( .A(n2483), .B(n2484), .Z(n275) );
  NANDN U417 ( .A(n2485), .B(n2486), .Z(n276) );
  AND U418 ( .A(n275), .B(n276), .Z(n2492) );
  NANDN U419 ( .A(n2504), .B(n2505), .Z(n277) );
  NANDN U420 ( .A(n2507), .B(n2506), .Z(n278) );
  NAND U421 ( .A(n277), .B(n278), .Z(n2513) );
  NANDN U422 ( .A(n2525), .B(n2526), .Z(n279) );
  NANDN U423 ( .A(n2527), .B(n2528), .Z(n280) );
  AND U424 ( .A(n279), .B(n280), .Z(n2534) );
  NANDN U425 ( .A(n2546), .B(n2547), .Z(n281) );
  NANDN U426 ( .A(n2549), .B(n2548), .Z(n282) );
  AND U427 ( .A(n281), .B(n282), .Z(n2555) );
  NANDN U428 ( .A(n2569), .B(n2570), .Z(n283) );
  NANDN U429 ( .A(n2567), .B(n2568), .Z(n284) );
  NAND U430 ( .A(n283), .B(n284), .Z(n2576) );
  NANDN U431 ( .A(n2590), .B(n2591), .Z(n285) );
  NANDN U432 ( .A(n2588), .B(n2589), .Z(n286) );
  NAND U433 ( .A(n285), .B(n286), .Z(n2597) );
  NANDN U434 ( .A(n2609), .B(n2610), .Z(n287) );
  NANDN U435 ( .A(n2612), .B(n2611), .Z(n288) );
  AND U436 ( .A(n287), .B(n288), .Z(n2618) );
  NANDN U437 ( .A(n2632), .B(n2633), .Z(n289) );
  NANDN U438 ( .A(n2630), .B(n2631), .Z(n290) );
  NAND U439 ( .A(n289), .B(n290), .Z(n2639) );
  NANDN U440 ( .A(n2651), .B(n2652), .Z(n291) );
  NANDN U441 ( .A(n2654), .B(n2653), .Z(n292) );
  AND U442 ( .A(n291), .B(n292), .Z(n2660) );
  NANDN U443 ( .A(n2674), .B(n2675), .Z(n293) );
  NANDN U444 ( .A(n2672), .B(n2673), .Z(n294) );
  NAND U445 ( .A(n293), .B(n294), .Z(n2681) );
  NANDN U446 ( .A(n2693), .B(n2694), .Z(n295) );
  NANDN U447 ( .A(n2696), .B(n2695), .Z(n296) );
  AND U448 ( .A(n295), .B(n296), .Z(n2702) );
  NANDN U449 ( .A(n2716), .B(n2717), .Z(n297) );
  NANDN U450 ( .A(n2714), .B(n2715), .Z(n298) );
  NAND U451 ( .A(n297), .B(n298), .Z(n2723) );
  NANDN U452 ( .A(n2735), .B(n2736), .Z(n299) );
  NANDN U453 ( .A(n2738), .B(n2737), .Z(n300) );
  NAND U454 ( .A(n299), .B(n300), .Z(n2744) );
  NANDN U455 ( .A(n2756), .B(n2757), .Z(n301) );
  NANDN U456 ( .A(n2759), .B(n2758), .Z(n302) );
  AND U457 ( .A(n301), .B(n302), .Z(n2765) );
  NANDN U458 ( .A(n2777), .B(n2778), .Z(n303) );
  NANDN U459 ( .A(n2780), .B(n2779), .Z(n304) );
  NAND U460 ( .A(n303), .B(n304), .Z(n2786) );
  NANDN U461 ( .A(n2798), .B(n2799), .Z(n305) );
  NANDN U462 ( .A(n2801), .B(n2800), .Z(n306) );
  NAND U463 ( .A(n305), .B(n306), .Z(n2807) );
  NANDN U464 ( .A(n2819), .B(n2820), .Z(n307) );
  NANDN U465 ( .A(n2821), .B(n2822), .Z(n308) );
  AND U466 ( .A(n307), .B(n308), .Z(n2828) );
  NANDN U467 ( .A(n2842), .B(n2843), .Z(n309) );
  NANDN U468 ( .A(n2840), .B(n2841), .Z(n310) );
  NAND U469 ( .A(n309), .B(n310), .Z(n2849) );
  NANDN U470 ( .A(n2863), .B(n2864), .Z(n311) );
  NANDN U471 ( .A(n2861), .B(n2862), .Z(n312) );
  NAND U472 ( .A(n311), .B(n312), .Z(n2870) );
  NANDN U473 ( .A(n2882), .B(n2883), .Z(n313) );
  NANDN U474 ( .A(n2884), .B(n2885), .Z(n314) );
  AND U475 ( .A(n313), .B(n314), .Z(n2891) );
  NANDN U476 ( .A(n2903), .B(n2904), .Z(n315) );
  NANDN U477 ( .A(n2906), .B(n2905), .Z(n316) );
  NAND U478 ( .A(n315), .B(n316), .Z(n2912) );
  NANDN U479 ( .A(n2924), .B(n2925), .Z(n317) );
  NANDN U480 ( .A(n2927), .B(n2926), .Z(n318) );
  NAND U481 ( .A(n317), .B(n318), .Z(n2933) );
  NANDN U482 ( .A(n2945), .B(n2946), .Z(n319) );
  NANDN U483 ( .A(n2948), .B(n2947), .Z(n320) );
  NAND U484 ( .A(n319), .B(n320), .Z(n2954) );
  NANDN U485 ( .A(n2966), .B(n2967), .Z(n321) );
  NANDN U486 ( .A(n2969), .B(n2968), .Z(n322) );
  AND U487 ( .A(n321), .B(n322), .Z(n2975) );
  NANDN U488 ( .A(n2989), .B(n2990), .Z(n323) );
  NANDN U489 ( .A(n2987), .B(n2988), .Z(n324) );
  NAND U490 ( .A(n323), .B(n324), .Z(n2996) );
  NANDN U491 ( .A(n3008), .B(n3009), .Z(n325) );
  NANDN U492 ( .A(n3011), .B(n3010), .Z(n326) );
  NAND U493 ( .A(n325), .B(n326), .Z(n3017) );
  NANDN U494 ( .A(n3029), .B(n3030), .Z(n327) );
  NANDN U495 ( .A(n3032), .B(n3031), .Z(n328) );
  AND U496 ( .A(n327), .B(n328), .Z(n3038) );
  NANDN U497 ( .A(n1316), .B(n1317), .Z(n329) );
  NANDN U498 ( .A(n1314), .B(n1315), .Z(n330) );
  NAND U499 ( .A(n329), .B(n330), .Z(n1323) );
  NANDN U500 ( .A(n1337), .B(n1338), .Z(n331) );
  NANDN U501 ( .A(n1335), .B(n1336), .Z(n332) );
  NAND U502 ( .A(n331), .B(n332), .Z(n1344) );
  NANDN U503 ( .A(n1358), .B(n1359), .Z(n333) );
  NANDN U504 ( .A(n1356), .B(n1357), .Z(n334) );
  NAND U505 ( .A(n333), .B(n334), .Z(n1365) );
  NANDN U506 ( .A(n1377), .B(n1378), .Z(n335) );
  NANDN U507 ( .A(n1379), .B(n1380), .Z(n336) );
  AND U508 ( .A(n335), .B(n336), .Z(n1386) );
  NANDN U509 ( .A(n1398), .B(n1399), .Z(n337) );
  NANDN U510 ( .A(n1401), .B(n1400), .Z(n338) );
  AND U511 ( .A(n337), .B(n338), .Z(n1407) );
  NANDN U512 ( .A(n1421), .B(n1422), .Z(n339) );
  NANDN U513 ( .A(n1419), .B(n1420), .Z(n340) );
  NAND U514 ( .A(n339), .B(n340), .Z(n1428) );
  NANDN U515 ( .A(n1440), .B(n1441), .Z(n341) );
  NANDN U516 ( .A(n1443), .B(n1442), .Z(n342) );
  NAND U517 ( .A(n341), .B(n342), .Z(n1449) );
  NANDN U518 ( .A(n1461), .B(n1462), .Z(n343) );
  NANDN U519 ( .A(n1464), .B(n1463), .Z(n344) );
  AND U520 ( .A(n343), .B(n344), .Z(n1470) );
  NANDN U521 ( .A(n1484), .B(n1485), .Z(n345) );
  NANDN U522 ( .A(n1482), .B(n1483), .Z(n346) );
  NAND U523 ( .A(n345), .B(n346), .Z(n1491) );
  NANDN U524 ( .A(n1503), .B(n1504), .Z(n347) );
  NANDN U525 ( .A(n1506), .B(n1505), .Z(n348) );
  AND U526 ( .A(n347), .B(n348), .Z(n1512) );
  NANDN U527 ( .A(n1524), .B(n1525), .Z(n349) );
  NANDN U528 ( .A(n1527), .B(n1526), .Z(n350) );
  NAND U529 ( .A(n349), .B(n350), .Z(n1533) );
  NANDN U530 ( .A(n1545), .B(n1546), .Z(n351) );
  NANDN U531 ( .A(n1548), .B(n1547), .Z(n352) );
  AND U532 ( .A(n351), .B(n352), .Z(n1554) );
  NANDN U533 ( .A(n1566), .B(n1567), .Z(n353) );
  NANDN U534 ( .A(n1569), .B(n1568), .Z(n354) );
  NAND U535 ( .A(n353), .B(n354), .Z(n1575) );
  NANDN U536 ( .A(n1587), .B(n1588), .Z(n355) );
  NANDN U537 ( .A(n1590), .B(n1589), .Z(n356) );
  AND U538 ( .A(n355), .B(n356), .Z(n1596) );
  NANDN U539 ( .A(n1608), .B(n1609), .Z(n357) );
  NANDN U540 ( .A(n1611), .B(n1610), .Z(n358) );
  NAND U541 ( .A(n357), .B(n358), .Z(n1617) );
  NANDN U542 ( .A(n1631), .B(n1632), .Z(n359) );
  NANDN U543 ( .A(n1629), .B(n1630), .Z(n360) );
  NAND U544 ( .A(n359), .B(n360), .Z(n1638) );
  NANDN U545 ( .A(n1650), .B(n1651), .Z(n361) );
  NANDN U546 ( .A(n1653), .B(n1652), .Z(n362) );
  AND U547 ( .A(n361), .B(n362), .Z(n1659) );
  NANDN U548 ( .A(n1673), .B(n1674), .Z(n363) );
  NANDN U549 ( .A(n1671), .B(n1672), .Z(n364) );
  NAND U550 ( .A(n363), .B(n364), .Z(n1680) );
  NANDN U551 ( .A(n1692), .B(n1693), .Z(n365) );
  NANDN U552 ( .A(n1695), .B(n1694), .Z(n366) );
  NAND U553 ( .A(n365), .B(n366), .Z(n1701) );
  NANDN U554 ( .A(n1713), .B(n1714), .Z(n367) );
  NANDN U555 ( .A(n1716), .B(n1715), .Z(n368) );
  AND U556 ( .A(n367), .B(n368), .Z(n1722) );
  NANDN U557 ( .A(n1736), .B(n1737), .Z(n369) );
  NANDN U558 ( .A(n1734), .B(n1735), .Z(n370) );
  NAND U559 ( .A(n369), .B(n370), .Z(n1743) );
  NANDN U560 ( .A(n1755), .B(n1756), .Z(n371) );
  NANDN U561 ( .A(n1758), .B(n1757), .Z(n372) );
  AND U562 ( .A(n371), .B(n372), .Z(n1764) );
  NANDN U563 ( .A(n1776), .B(n1777), .Z(n373) );
  NANDN U564 ( .A(n1779), .B(n1778), .Z(n374) );
  NAND U565 ( .A(n373), .B(n374), .Z(n1785) );
  NANDN U566 ( .A(n1797), .B(n1798), .Z(n375) );
  NANDN U567 ( .A(n1800), .B(n1799), .Z(n376) );
  NAND U568 ( .A(n375), .B(n376), .Z(n1806) );
  NANDN U569 ( .A(n1820), .B(n1821), .Z(n377) );
  NANDN U570 ( .A(n1818), .B(n1819), .Z(n378) );
  NAND U571 ( .A(n377), .B(n378), .Z(n1827) );
  NANDN U572 ( .A(n1839), .B(n1840), .Z(n379) );
  NANDN U573 ( .A(n1842), .B(n1841), .Z(n380) );
  NAND U574 ( .A(n379), .B(n380), .Z(n1848) );
  NANDN U575 ( .A(n1860), .B(n1861), .Z(n381) );
  NANDN U576 ( .A(n1863), .B(n1862), .Z(n382) );
  AND U577 ( .A(n381), .B(n382), .Z(n1869) );
  NANDN U578 ( .A(n1883), .B(n1884), .Z(n383) );
  NANDN U579 ( .A(n1881), .B(n1882), .Z(n384) );
  NAND U580 ( .A(n383), .B(n384), .Z(n1890) );
  NANDN U581 ( .A(n1902), .B(n1903), .Z(n385) );
  NANDN U582 ( .A(n1905), .B(n1904), .Z(n386) );
  NAND U583 ( .A(n385), .B(n386), .Z(n1911) );
  NANDN U584 ( .A(n1923), .B(n1924), .Z(n387) );
  NANDN U585 ( .A(n1926), .B(n1925), .Z(n388) );
  AND U586 ( .A(n387), .B(n388), .Z(n1932) );
  NANDN U587 ( .A(n1946), .B(n1947), .Z(n389) );
  NANDN U588 ( .A(n1944), .B(n1945), .Z(n390) );
  NAND U589 ( .A(n389), .B(n390), .Z(n1953) );
  NANDN U590 ( .A(n1965), .B(n1966), .Z(n391) );
  NANDN U591 ( .A(n1968), .B(n1967), .Z(n392) );
  NAND U592 ( .A(n391), .B(n392), .Z(n1974) );
  NANDN U593 ( .A(n1986), .B(n1987), .Z(n393) );
  NANDN U594 ( .A(n1989), .B(n1988), .Z(n394) );
  AND U595 ( .A(n393), .B(n394), .Z(n1995) );
  NANDN U596 ( .A(n2007), .B(n2008), .Z(n395) );
  NANDN U597 ( .A(n2010), .B(n2009), .Z(n396) );
  NAND U598 ( .A(n395), .B(n396), .Z(n2016) );
  NANDN U599 ( .A(n2030), .B(n2031), .Z(n397) );
  NANDN U600 ( .A(n2028), .B(n2029), .Z(n398) );
  NAND U601 ( .A(n397), .B(n398), .Z(n2037) );
  NANDN U602 ( .A(n2051), .B(n2052), .Z(n399) );
  NANDN U603 ( .A(n2049), .B(n2050), .Z(n400) );
  NAND U604 ( .A(n399), .B(n400), .Z(n2058) );
  NANDN U605 ( .A(n2070), .B(n2071), .Z(n401) );
  NANDN U606 ( .A(n2073), .B(n2072), .Z(n402) );
  AND U607 ( .A(n401), .B(n402), .Z(n2079) );
  NANDN U608 ( .A(n2091), .B(n2092), .Z(n403) );
  NANDN U609 ( .A(n2094), .B(n2093), .Z(n404) );
  NAND U610 ( .A(n403), .B(n404), .Z(n2100) );
  NANDN U611 ( .A(n2112), .B(n2113), .Z(n405) );
  NANDN U612 ( .A(n2115), .B(n2114), .Z(n406) );
  NAND U613 ( .A(n405), .B(n406), .Z(n2121) );
  NANDN U614 ( .A(n2133), .B(n2134), .Z(n407) );
  NANDN U615 ( .A(n2136), .B(n2135), .Z(n408) );
  AND U616 ( .A(n407), .B(n408), .Z(n2142) );
  NANDN U617 ( .A(n2156), .B(n2157), .Z(n409) );
  NANDN U618 ( .A(n2154), .B(n2155), .Z(n410) );
  NAND U619 ( .A(n409), .B(n410), .Z(n2163) );
  NANDN U620 ( .A(n2175), .B(n2176), .Z(n411) );
  NANDN U621 ( .A(n2178), .B(n2177), .Z(n412) );
  AND U622 ( .A(n411), .B(n412), .Z(n2184) );
  NANDN U623 ( .A(n2198), .B(n2199), .Z(n413) );
  NANDN U624 ( .A(n2196), .B(n2197), .Z(n414) );
  NAND U625 ( .A(n413), .B(n414), .Z(n2205) );
  NANDN U626 ( .A(n2217), .B(n2218), .Z(n415) );
  NANDN U627 ( .A(n2220), .B(n2219), .Z(n416) );
  AND U628 ( .A(n415), .B(n416), .Z(n2226) );
  NANDN U629 ( .A(n2238), .B(n2239), .Z(n417) );
  NANDN U630 ( .A(n2241), .B(n2240), .Z(n418) );
  NAND U631 ( .A(n417), .B(n418), .Z(n2247) );
  NANDN U632 ( .A(n2259), .B(n2260), .Z(n419) );
  NANDN U633 ( .A(n2262), .B(n2261), .Z(n420) );
  AND U634 ( .A(n419), .B(n420), .Z(n2268) );
  NANDN U635 ( .A(n2282), .B(n2283), .Z(n421) );
  NANDN U636 ( .A(n2280), .B(n2281), .Z(n422) );
  NAND U637 ( .A(n421), .B(n422), .Z(n2289) );
  NANDN U638 ( .A(n2303), .B(n2304), .Z(n423) );
  NANDN U639 ( .A(n2301), .B(n2302), .Z(n424) );
  NAND U640 ( .A(n423), .B(n424), .Z(n2310) );
  NANDN U641 ( .A(n2322), .B(n2323), .Z(n425) );
  NANDN U642 ( .A(n2324), .B(n2325), .Z(n426) );
  AND U643 ( .A(n425), .B(n426), .Z(n2331) );
  NANDN U644 ( .A(n2343), .B(n2344), .Z(n427) );
  NANDN U645 ( .A(n2346), .B(n2345), .Z(n428) );
  NAND U646 ( .A(n427), .B(n428), .Z(n2352) );
  NANDN U647 ( .A(n2364), .B(n2365), .Z(n429) );
  NANDN U648 ( .A(n2367), .B(n2366), .Z(n430) );
  NAND U649 ( .A(n429), .B(n430), .Z(n2373) );
  NANDN U650 ( .A(n2385), .B(n2386), .Z(n431) );
  NANDN U651 ( .A(n2388), .B(n2387), .Z(n432) );
  AND U652 ( .A(n431), .B(n432), .Z(n2394) );
  NANDN U653 ( .A(n2408), .B(n2409), .Z(n433) );
  NANDN U654 ( .A(n2406), .B(n2407), .Z(n434) );
  NAND U655 ( .A(n433), .B(n434), .Z(n2415) );
  NANDN U656 ( .A(n2427), .B(n2428), .Z(n435) );
  NANDN U657 ( .A(n2430), .B(n2429), .Z(n436) );
  NAND U658 ( .A(n435), .B(n436), .Z(n2436) );
  NANDN U659 ( .A(n2448), .B(n2449), .Z(n437) );
  NANDN U660 ( .A(n2451), .B(n2450), .Z(n438) );
  NAND U661 ( .A(n437), .B(n438), .Z(n2457) );
  NANDN U662 ( .A(n2469), .B(n2470), .Z(n439) );
  NANDN U663 ( .A(n2472), .B(n2471), .Z(n440) );
  AND U664 ( .A(n439), .B(n440), .Z(n2478) );
  NANDN U665 ( .A(n2492), .B(n2493), .Z(n441) );
  NANDN U666 ( .A(n2490), .B(n2491), .Z(n442) );
  NAND U667 ( .A(n441), .B(n442), .Z(n2499) );
  NANDN U668 ( .A(n2511), .B(n2512), .Z(n443) );
  NANDN U669 ( .A(n2514), .B(n2513), .Z(n444) );
  NAND U670 ( .A(n443), .B(n444), .Z(n2520) );
  NANDN U671 ( .A(n2532), .B(n2533), .Z(n445) );
  NANDN U672 ( .A(n2534), .B(n2535), .Z(n446) );
  AND U673 ( .A(n445), .B(n446), .Z(n2541) );
  NANDN U674 ( .A(n2555), .B(n2556), .Z(n447) );
  NANDN U675 ( .A(n2553), .B(n2554), .Z(n448) );
  NAND U676 ( .A(n447), .B(n448), .Z(n2562) );
  NANDN U677 ( .A(n2574), .B(n2575), .Z(n449) );
  NANDN U678 ( .A(n2577), .B(n2576), .Z(n450) );
  NAND U679 ( .A(n449), .B(n450), .Z(n2583) );
  NANDN U680 ( .A(n2595), .B(n2596), .Z(n451) );
  NANDN U681 ( .A(n2598), .B(n2597), .Z(n452) );
  AND U682 ( .A(n451), .B(n452), .Z(n2604) );
  NANDN U683 ( .A(n2618), .B(n2619), .Z(n453) );
  NANDN U684 ( .A(n2616), .B(n2617), .Z(n454) );
  NAND U685 ( .A(n453), .B(n454), .Z(n2625) );
  NANDN U686 ( .A(n2637), .B(n2638), .Z(n455) );
  NANDN U687 ( .A(n2640), .B(n2639), .Z(n456) );
  NAND U688 ( .A(n455), .B(n456), .Z(n2646) );
  NANDN U689 ( .A(n2660), .B(n2661), .Z(n457) );
  NANDN U690 ( .A(n2658), .B(n2659), .Z(n458) );
  NAND U691 ( .A(n457), .B(n458), .Z(n2667) );
  NANDN U692 ( .A(n2679), .B(n2680), .Z(n459) );
  NANDN U693 ( .A(n2682), .B(n2681), .Z(n460) );
  NAND U694 ( .A(n459), .B(n460), .Z(n2688) );
  NANDN U695 ( .A(n2702), .B(n2703), .Z(n461) );
  NANDN U696 ( .A(n2700), .B(n2701), .Z(n462) );
  NAND U697 ( .A(n461), .B(n462), .Z(n2709) );
  NANDN U698 ( .A(n2721), .B(n2722), .Z(n463) );
  NANDN U699 ( .A(n2724), .B(n2723), .Z(n464) );
  NAND U700 ( .A(n463), .B(n464), .Z(n2730) );
  NANDN U701 ( .A(n2742), .B(n2743), .Z(n465) );
  NANDN U702 ( .A(n2745), .B(n2744), .Z(n466) );
  AND U703 ( .A(n465), .B(n466), .Z(n2751) );
  NANDN U704 ( .A(n2765), .B(n2766), .Z(n467) );
  NANDN U705 ( .A(n2763), .B(n2764), .Z(n468) );
  NAND U706 ( .A(n467), .B(n468), .Z(n2772) );
  NANDN U707 ( .A(n2784), .B(n2785), .Z(n469) );
  NANDN U708 ( .A(n2787), .B(n2786), .Z(n470) );
  NAND U709 ( .A(n469), .B(n470), .Z(n2793) );
  NANDN U710 ( .A(n2805), .B(n2806), .Z(n471) );
  NANDN U711 ( .A(n2808), .B(n2807), .Z(n472) );
  AND U712 ( .A(n471), .B(n472), .Z(n2814) );
  NANDN U713 ( .A(n2828), .B(n2829), .Z(n473) );
  NANDN U714 ( .A(n2826), .B(n2827), .Z(n474) );
  NAND U715 ( .A(n473), .B(n474), .Z(n2835) );
  NANDN U716 ( .A(n2847), .B(n2848), .Z(n475) );
  NANDN U717 ( .A(n2850), .B(n2849), .Z(n476) );
  NAND U718 ( .A(n475), .B(n476), .Z(n2856) );
  NANDN U719 ( .A(n2868), .B(n2869), .Z(n477) );
  NANDN U720 ( .A(n2871), .B(n2870), .Z(n478) );
  NAND U721 ( .A(n477), .B(n478), .Z(n2877) );
  NANDN U722 ( .A(n2889), .B(n2890), .Z(n479) );
  NANDN U723 ( .A(n2891), .B(n2892), .Z(n480) );
  AND U724 ( .A(n479), .B(n480), .Z(n2898) );
  NANDN U725 ( .A(n2910), .B(n2911), .Z(n481) );
  NANDN U726 ( .A(n2913), .B(n2912), .Z(n482) );
  NAND U727 ( .A(n481), .B(n482), .Z(n2919) );
  NANDN U728 ( .A(n2931), .B(n2932), .Z(n483) );
  NANDN U729 ( .A(n2934), .B(n2933), .Z(n484) );
  AND U730 ( .A(n483), .B(n484), .Z(n2940) );
  NANDN U731 ( .A(n2952), .B(n2953), .Z(n485) );
  NANDN U732 ( .A(n2955), .B(n2954), .Z(n486) );
  NAND U733 ( .A(n485), .B(n486), .Z(n2961) );
  NANDN U734 ( .A(n2975), .B(n2976), .Z(n487) );
  NANDN U735 ( .A(n2973), .B(n2974), .Z(n488) );
  NAND U736 ( .A(n487), .B(n488), .Z(n2982) );
  NANDN U737 ( .A(n2994), .B(n2995), .Z(n489) );
  NANDN U738 ( .A(n2997), .B(n2996), .Z(n490) );
  AND U739 ( .A(n489), .B(n490), .Z(n3003) );
  NANDN U740 ( .A(n3015), .B(n3016), .Z(n491) );
  NANDN U741 ( .A(n3018), .B(n3017), .Z(n492) );
  NAND U742 ( .A(n491), .B(n492), .Z(n3024) );
  NANDN U743 ( .A(n3038), .B(n3039), .Z(n493) );
  NANDN U744 ( .A(n3036), .B(n3037), .Z(n494) );
  NAND U745 ( .A(n493), .B(n494), .Z(n3044) );
  NANDN U746 ( .A(n3053), .B(n3043), .Z(n495) );
  NANDN U747 ( .A(n3045), .B(n3044), .Z(n496) );
  AND U748 ( .A(n495), .B(n496), .Z(n3055) );
  NAND U749 ( .A(n1283), .B(n1284), .Z(n497) );
  XOR U750 ( .A(n1283), .B(n1284), .Z(n498) );
  NAND U751 ( .A(n498), .B(sreg[257]), .Z(n499) );
  NAND U752 ( .A(n497), .B(n499), .Z(n1294) );
  NAND U753 ( .A(n1319), .B(n1318), .Z(n500) );
  XOR U754 ( .A(n1319), .B(n1318), .Z(n501) );
  NANDN U755 ( .A(sreg[261]), .B(n501), .Z(n502) );
  NAND U756 ( .A(n500), .B(n502), .Z(n1325) );
  XOR U757 ( .A(sreg[264]), .B(n1339), .Z(n503) );
  NANDN U758 ( .A(n1340), .B(n503), .Z(n504) );
  NAND U759 ( .A(sreg[264]), .B(n1339), .Z(n505) );
  AND U760 ( .A(n504), .B(n505), .Z(n1346) );
  XOR U761 ( .A(sreg[267]), .B(n1360), .Z(n506) );
  NANDN U762 ( .A(n1361), .B(n506), .Z(n507) );
  NAND U763 ( .A(sreg[267]), .B(n1360), .Z(n508) );
  AND U764 ( .A(n507), .B(n508), .Z(n1367) );
  NAND U765 ( .A(n1381), .B(n1382), .Z(n509) );
  XOR U766 ( .A(n1381), .B(n1382), .Z(n510) );
  NANDN U767 ( .A(sreg[270]), .B(n510), .Z(n511) );
  NAND U768 ( .A(n509), .B(n511), .Z(n1388) );
  NAND U769 ( .A(n1402), .B(n1403), .Z(n512) );
  XOR U770 ( .A(n1402), .B(n1403), .Z(n513) );
  NAND U771 ( .A(n513), .B(sreg[273]), .Z(n514) );
  NAND U772 ( .A(n512), .B(n514), .Z(n1409) );
  XOR U773 ( .A(sreg[276]), .B(n1423), .Z(n515) );
  NANDN U774 ( .A(n1424), .B(n515), .Z(n516) );
  NAND U775 ( .A(sreg[276]), .B(n1423), .Z(n517) );
  AND U776 ( .A(n516), .B(n517), .Z(n1430) );
  NAND U777 ( .A(sreg[279]), .B(n1445), .Z(n518) );
  XOR U778 ( .A(sreg[279]), .B(n1445), .Z(n519) );
  NANDN U779 ( .A(n1444), .B(n519), .Z(n520) );
  NAND U780 ( .A(n518), .B(n520), .Z(n1451) );
  NAND U781 ( .A(sreg[282]), .B(n1466), .Z(n521) );
  XOR U782 ( .A(sreg[282]), .B(n1466), .Z(n522) );
  NAND U783 ( .A(n522), .B(n1465), .Z(n523) );
  NAND U784 ( .A(n521), .B(n523), .Z(n1472) );
  XOR U785 ( .A(sreg[285]), .B(n1486), .Z(n524) );
  NANDN U786 ( .A(n1487), .B(n524), .Z(n525) );
  NAND U787 ( .A(sreg[285]), .B(n1486), .Z(n526) );
  AND U788 ( .A(n525), .B(n526), .Z(n1493) );
  NAND U789 ( .A(sreg[288]), .B(n1508), .Z(n527) );
  XOR U790 ( .A(sreg[288]), .B(n1508), .Z(n528) );
  NANDN U791 ( .A(n1507), .B(n528), .Z(n529) );
  NAND U792 ( .A(n527), .B(n529), .Z(n1514) );
  NAND U793 ( .A(sreg[291]), .B(n1529), .Z(n530) );
  XOR U794 ( .A(sreg[291]), .B(n1529), .Z(n531) );
  NANDN U795 ( .A(n1528), .B(n531), .Z(n532) );
  NAND U796 ( .A(n530), .B(n532), .Z(n1535) );
  NAND U797 ( .A(n1549), .B(n1550), .Z(n533) );
  XOR U798 ( .A(n1549), .B(n1550), .Z(n534) );
  NAND U799 ( .A(n534), .B(sreg[294]), .Z(n535) );
  NAND U800 ( .A(n533), .B(n535), .Z(n1556) );
  NAND U801 ( .A(n1570), .B(n1571), .Z(n536) );
  XOR U802 ( .A(n1570), .B(n1571), .Z(n537) );
  NAND U803 ( .A(n537), .B(sreg[297]), .Z(n538) );
  NAND U804 ( .A(n536), .B(n538), .Z(n1577) );
  NAND U805 ( .A(sreg[300]), .B(n1592), .Z(n539) );
  XOR U806 ( .A(sreg[300]), .B(n1592), .Z(n540) );
  NANDN U807 ( .A(n1591), .B(n540), .Z(n541) );
  NAND U808 ( .A(n539), .B(n541), .Z(n1598) );
  NAND U809 ( .A(n1612), .B(n1613), .Z(n542) );
  XOR U810 ( .A(n1612), .B(n1613), .Z(n543) );
  NAND U811 ( .A(n543), .B(sreg[303]), .Z(n544) );
  NAND U812 ( .A(n542), .B(n544), .Z(n1619) );
  XOR U813 ( .A(sreg[306]), .B(n1633), .Z(n545) );
  NANDN U814 ( .A(n1634), .B(n545), .Z(n546) );
  NAND U815 ( .A(sreg[306]), .B(n1633), .Z(n547) );
  AND U816 ( .A(n546), .B(n547), .Z(n1640) );
  NAND U817 ( .A(sreg[309]), .B(n1655), .Z(n548) );
  XOR U818 ( .A(sreg[309]), .B(n1655), .Z(n549) );
  NANDN U819 ( .A(n1654), .B(n549), .Z(n550) );
  NAND U820 ( .A(n548), .B(n550), .Z(n1661) );
  NAND U821 ( .A(n1675), .B(n1676), .Z(n551) );
  XOR U822 ( .A(n1675), .B(n1676), .Z(n552) );
  NANDN U823 ( .A(sreg[312]), .B(n552), .Z(n553) );
  NAND U824 ( .A(n551), .B(n553), .Z(n1682) );
  NAND U825 ( .A(n1696), .B(n1697), .Z(n554) );
  XOR U826 ( .A(n1696), .B(n1697), .Z(n555) );
  NAND U827 ( .A(n555), .B(sreg[315]), .Z(n556) );
  NAND U828 ( .A(n554), .B(n556), .Z(n1703) );
  NAND U829 ( .A(sreg[318]), .B(n1718), .Z(n557) );
  XOR U830 ( .A(sreg[318]), .B(n1718), .Z(n558) );
  NANDN U831 ( .A(n1717), .B(n558), .Z(n559) );
  NAND U832 ( .A(n557), .B(n559), .Z(n1724) );
  XOR U833 ( .A(sreg[321]), .B(n1738), .Z(n560) );
  NANDN U834 ( .A(n1739), .B(n560), .Z(n561) );
  NAND U835 ( .A(sreg[321]), .B(n1738), .Z(n562) );
  AND U836 ( .A(n561), .B(n562), .Z(n1745) );
  NAND U837 ( .A(n1759), .B(n1760), .Z(n563) );
  XOR U838 ( .A(n1759), .B(n1760), .Z(n564) );
  NAND U839 ( .A(n564), .B(sreg[324]), .Z(n565) );
  NAND U840 ( .A(n563), .B(n565), .Z(n1766) );
  NAND U841 ( .A(n1780), .B(n1781), .Z(n566) );
  XOR U842 ( .A(n1780), .B(n1781), .Z(n567) );
  NAND U843 ( .A(n567), .B(sreg[327]), .Z(n568) );
  NAND U844 ( .A(n566), .B(n568), .Z(n1787) );
  NAND U845 ( .A(n1801), .B(n1802), .Z(n569) );
  XOR U846 ( .A(n1801), .B(n1802), .Z(n570) );
  NAND U847 ( .A(n570), .B(sreg[330]), .Z(n571) );
  NAND U848 ( .A(n569), .B(n571), .Z(n1808) );
  XOR U849 ( .A(sreg[333]), .B(n1822), .Z(n572) );
  NANDN U850 ( .A(n1823), .B(n572), .Z(n573) );
  NAND U851 ( .A(sreg[333]), .B(n1822), .Z(n574) );
  AND U852 ( .A(n573), .B(n574), .Z(n1829) );
  NAND U853 ( .A(n1843), .B(n1844), .Z(n575) );
  XOR U854 ( .A(n1843), .B(n1844), .Z(n576) );
  NAND U855 ( .A(n576), .B(sreg[336]), .Z(n577) );
  NAND U856 ( .A(n575), .B(n577), .Z(n1850) );
  NAND U857 ( .A(sreg[339]), .B(n1865), .Z(n578) );
  XOR U858 ( .A(sreg[339]), .B(n1865), .Z(n579) );
  NANDN U859 ( .A(n1864), .B(n579), .Z(n580) );
  NAND U860 ( .A(n578), .B(n580), .Z(n1871) );
  XOR U861 ( .A(sreg[342]), .B(n1885), .Z(n581) );
  NANDN U862 ( .A(n1886), .B(n581), .Z(n582) );
  NAND U863 ( .A(sreg[342]), .B(n1885), .Z(n583) );
  AND U864 ( .A(n582), .B(n583), .Z(n1892) );
  NAND U865 ( .A(n1906), .B(n1907), .Z(n584) );
  XOR U866 ( .A(n1906), .B(n1907), .Z(n585) );
  NAND U867 ( .A(n585), .B(sreg[345]), .Z(n586) );
  NAND U868 ( .A(n584), .B(n586), .Z(n1913) );
  NAND U869 ( .A(sreg[348]), .B(n1928), .Z(n587) );
  XOR U870 ( .A(sreg[348]), .B(n1928), .Z(n588) );
  NANDN U871 ( .A(n1927), .B(n588), .Z(n589) );
  NAND U872 ( .A(n587), .B(n589), .Z(n1934) );
  XOR U873 ( .A(sreg[351]), .B(n1948), .Z(n590) );
  NANDN U874 ( .A(n1949), .B(n590), .Z(n591) );
  NAND U875 ( .A(sreg[351]), .B(n1948), .Z(n592) );
  AND U876 ( .A(n591), .B(n592), .Z(n1955) );
  NAND U877 ( .A(sreg[354]), .B(n1970), .Z(n593) );
  XOR U878 ( .A(sreg[354]), .B(n1970), .Z(n594) );
  NANDN U879 ( .A(n1969), .B(n594), .Z(n595) );
  NAND U880 ( .A(n593), .B(n595), .Z(n1976) );
  NAND U881 ( .A(n1990), .B(n1991), .Z(n596) );
  XOR U882 ( .A(n1990), .B(n1991), .Z(n597) );
  NAND U883 ( .A(n597), .B(sreg[357]), .Z(n598) );
  NAND U884 ( .A(n596), .B(n598), .Z(n1997) );
  NAND U885 ( .A(sreg[360]), .B(n2012), .Z(n599) );
  XOR U886 ( .A(sreg[360]), .B(n2012), .Z(n600) );
  NANDN U887 ( .A(n2011), .B(n600), .Z(n601) );
  NAND U888 ( .A(n599), .B(n601), .Z(n2018) );
  XOR U889 ( .A(sreg[363]), .B(n2032), .Z(n602) );
  NANDN U890 ( .A(n2033), .B(n602), .Z(n603) );
  NAND U891 ( .A(sreg[363]), .B(n2032), .Z(n604) );
  AND U892 ( .A(n603), .B(n604), .Z(n2039) );
  NAND U893 ( .A(n2053), .B(n2054), .Z(n605) );
  XOR U894 ( .A(n2053), .B(n2054), .Z(n606) );
  NANDN U895 ( .A(sreg[366]), .B(n606), .Z(n607) );
  NAND U896 ( .A(n605), .B(n607), .Z(n2060) );
  NAND U897 ( .A(n2074), .B(n2075), .Z(n608) );
  XOR U898 ( .A(n2074), .B(n2075), .Z(n609) );
  NAND U899 ( .A(n609), .B(sreg[369]), .Z(n610) );
  NAND U900 ( .A(n608), .B(n610), .Z(n2081) );
  NAND U901 ( .A(n2095), .B(n2096), .Z(n611) );
  XOR U902 ( .A(n2095), .B(n2096), .Z(n612) );
  NAND U903 ( .A(n612), .B(sreg[372]), .Z(n613) );
  NAND U904 ( .A(n611), .B(n613), .Z(n2102) );
  NAND U905 ( .A(sreg[375]), .B(n2117), .Z(n614) );
  XOR U906 ( .A(sreg[375]), .B(n2117), .Z(n615) );
  NANDN U907 ( .A(n2116), .B(n615), .Z(n616) );
  NAND U908 ( .A(n614), .B(n616), .Z(n2123) );
  NAND U909 ( .A(n2137), .B(n2138), .Z(n617) );
  XOR U910 ( .A(n2137), .B(n2138), .Z(n618) );
  NAND U911 ( .A(n618), .B(sreg[378]), .Z(n619) );
  NAND U912 ( .A(n617), .B(n619), .Z(n2144) );
  XOR U913 ( .A(sreg[381]), .B(n2158), .Z(n620) );
  NANDN U914 ( .A(n2159), .B(n620), .Z(n621) );
  NAND U915 ( .A(sreg[381]), .B(n2158), .Z(n622) );
  AND U916 ( .A(n621), .B(n622), .Z(n2165) );
  NAND U917 ( .A(sreg[384]), .B(n2180), .Z(n623) );
  XOR U918 ( .A(sreg[384]), .B(n2180), .Z(n624) );
  NANDN U919 ( .A(n2179), .B(n624), .Z(n625) );
  NAND U920 ( .A(n623), .B(n625), .Z(n2186) );
  XOR U921 ( .A(sreg[387]), .B(n2200), .Z(n626) );
  NANDN U922 ( .A(n2201), .B(n626), .Z(n627) );
  NAND U923 ( .A(sreg[387]), .B(n2200), .Z(n628) );
  AND U924 ( .A(n627), .B(n628), .Z(n2207) );
  NAND U925 ( .A(n2221), .B(n2222), .Z(n629) );
  XOR U926 ( .A(n2221), .B(n2222), .Z(n630) );
  NAND U927 ( .A(n630), .B(sreg[390]), .Z(n631) );
  NAND U928 ( .A(n629), .B(n631), .Z(n2228) );
  NAND U929 ( .A(n2242), .B(n2243), .Z(n632) );
  XOR U930 ( .A(n2242), .B(n2243), .Z(n633) );
  NAND U931 ( .A(n633), .B(sreg[393]), .Z(n634) );
  NAND U932 ( .A(n632), .B(n634), .Z(n2249) );
  NAND U933 ( .A(sreg[396]), .B(n2264), .Z(n635) );
  XOR U934 ( .A(sreg[396]), .B(n2264), .Z(n636) );
  NANDN U935 ( .A(n2263), .B(n636), .Z(n637) );
  NAND U936 ( .A(n635), .B(n637), .Z(n2270) );
  XOR U937 ( .A(sreg[399]), .B(n2284), .Z(n638) );
  NANDN U938 ( .A(n2285), .B(n638), .Z(n639) );
  NAND U939 ( .A(sreg[399]), .B(n2284), .Z(n640) );
  AND U940 ( .A(n639), .B(n640), .Z(n2291) );
  XOR U941 ( .A(sreg[402]), .B(n2305), .Z(n641) );
  NANDN U942 ( .A(n2306), .B(n641), .Z(n642) );
  NAND U943 ( .A(sreg[402]), .B(n2305), .Z(n643) );
  AND U944 ( .A(n642), .B(n643), .Z(n2312) );
  NAND U945 ( .A(n2326), .B(n2327), .Z(n644) );
  XOR U946 ( .A(n2326), .B(n2327), .Z(n645) );
  NANDN U947 ( .A(sreg[405]), .B(n645), .Z(n646) );
  NAND U948 ( .A(n644), .B(n646), .Z(n2333) );
  NAND U949 ( .A(n2347), .B(n2348), .Z(n647) );
  XOR U950 ( .A(n2347), .B(n2348), .Z(n648) );
  NAND U951 ( .A(n648), .B(sreg[408]), .Z(n649) );
  NAND U952 ( .A(n647), .B(n649), .Z(n2354) );
  NAND U953 ( .A(n2368), .B(n2369), .Z(n650) );
  XOR U954 ( .A(n2368), .B(n2369), .Z(n651) );
  NAND U955 ( .A(n651), .B(sreg[411]), .Z(n652) );
  NAND U956 ( .A(n650), .B(n652), .Z(n2375) );
  NAND U957 ( .A(sreg[414]), .B(n2390), .Z(n653) );
  XOR U958 ( .A(sreg[414]), .B(n2390), .Z(n654) );
  NANDN U959 ( .A(n2389), .B(n654), .Z(n655) );
  NAND U960 ( .A(n653), .B(n655), .Z(n2396) );
  XOR U961 ( .A(sreg[417]), .B(n2410), .Z(n656) );
  NANDN U962 ( .A(n2411), .B(n656), .Z(n657) );
  NAND U963 ( .A(sreg[417]), .B(n2410), .Z(n658) );
  AND U964 ( .A(n657), .B(n658), .Z(n2417) );
  NAND U965 ( .A(sreg[420]), .B(n2432), .Z(n659) );
  XOR U966 ( .A(sreg[420]), .B(n2432), .Z(n660) );
  NANDN U967 ( .A(n2431), .B(n660), .Z(n661) );
  NAND U968 ( .A(n659), .B(n661), .Z(n2438) );
  NAND U969 ( .A(n2452), .B(n2453), .Z(n662) );
  XOR U970 ( .A(n2452), .B(n2453), .Z(n663) );
  NAND U971 ( .A(n663), .B(sreg[423]), .Z(n664) );
  NAND U972 ( .A(n662), .B(n664), .Z(n2459) );
  NAND U973 ( .A(n2473), .B(n2474), .Z(n665) );
  XOR U974 ( .A(n2473), .B(n2474), .Z(n666) );
  NAND U975 ( .A(n666), .B(sreg[426]), .Z(n667) );
  NAND U976 ( .A(n665), .B(n667), .Z(n2480) );
  NAND U977 ( .A(n2494), .B(n2495), .Z(n668) );
  XOR U978 ( .A(n2494), .B(n2495), .Z(n669) );
  NANDN U979 ( .A(sreg[429]), .B(n669), .Z(n670) );
  NAND U980 ( .A(n668), .B(n670), .Z(n2501) );
  NAND U981 ( .A(n2515), .B(n2516), .Z(n671) );
  XOR U982 ( .A(n2515), .B(n2516), .Z(n672) );
  NAND U983 ( .A(n672), .B(sreg[432]), .Z(n673) );
  NAND U984 ( .A(n671), .B(n673), .Z(n2522) );
  NAND U985 ( .A(n2536), .B(n2537), .Z(n674) );
  XOR U986 ( .A(n2536), .B(n2537), .Z(n675) );
  NANDN U987 ( .A(sreg[435]), .B(n675), .Z(n676) );
  NAND U988 ( .A(n674), .B(n676), .Z(n2543) );
  XOR U989 ( .A(sreg[438]), .B(n2557), .Z(n677) );
  NANDN U990 ( .A(n2558), .B(n677), .Z(n678) );
  NAND U991 ( .A(sreg[438]), .B(n2557), .Z(n679) );
  AND U992 ( .A(n678), .B(n679), .Z(n2564) );
  NAND U993 ( .A(sreg[441]), .B(n2579), .Z(n680) );
  XOR U994 ( .A(sreg[441]), .B(n2579), .Z(n681) );
  NANDN U995 ( .A(n2578), .B(n681), .Z(n682) );
  NAND U996 ( .A(n680), .B(n682), .Z(n2585) );
  NAND U997 ( .A(sreg[444]), .B(n2600), .Z(n683) );
  XOR U998 ( .A(sreg[444]), .B(n2600), .Z(n684) );
  NANDN U999 ( .A(n2599), .B(n684), .Z(n685) );
  NAND U1000 ( .A(n683), .B(n685), .Z(n2606) );
  XOR U1001 ( .A(sreg[447]), .B(n2620), .Z(n686) );
  NANDN U1002 ( .A(n2621), .B(n686), .Z(n687) );
  NAND U1003 ( .A(sreg[447]), .B(n2620), .Z(n688) );
  AND U1004 ( .A(n687), .B(n688), .Z(n2627) );
  NAND U1005 ( .A(sreg[450]), .B(n2642), .Z(n689) );
  XOR U1006 ( .A(sreg[450]), .B(n2642), .Z(n690) );
  NANDN U1007 ( .A(n2641), .B(n690), .Z(n691) );
  NAND U1008 ( .A(n689), .B(n691), .Z(n2648) );
  XOR U1009 ( .A(sreg[453]), .B(n2662), .Z(n692) );
  NANDN U1010 ( .A(n2663), .B(n692), .Z(n693) );
  NAND U1011 ( .A(sreg[453]), .B(n2662), .Z(n694) );
  AND U1012 ( .A(n693), .B(n694), .Z(n2669) );
  NAND U1013 ( .A(sreg[456]), .B(n2684), .Z(n695) );
  XOR U1014 ( .A(sreg[456]), .B(n2684), .Z(n696) );
  NANDN U1015 ( .A(n2683), .B(n696), .Z(n697) );
  NAND U1016 ( .A(n695), .B(n697), .Z(n2690) );
  XOR U1017 ( .A(sreg[459]), .B(n2704), .Z(n698) );
  NANDN U1018 ( .A(n2705), .B(n698), .Z(n699) );
  NAND U1019 ( .A(sreg[459]), .B(n2704), .Z(n700) );
  AND U1020 ( .A(n699), .B(n700), .Z(n2711) );
  NAND U1021 ( .A(sreg[462]), .B(n2726), .Z(n701) );
  XOR U1022 ( .A(sreg[462]), .B(n2726), .Z(n702) );
  NANDN U1023 ( .A(n2725), .B(n702), .Z(n703) );
  NAND U1024 ( .A(n701), .B(n703), .Z(n2732) );
  NAND U1025 ( .A(n2746), .B(n2747), .Z(n704) );
  XOR U1026 ( .A(n2746), .B(n2747), .Z(n705) );
  NAND U1027 ( .A(n705), .B(sreg[465]), .Z(n706) );
  NAND U1028 ( .A(n704), .B(n706), .Z(n2753) );
  XOR U1029 ( .A(sreg[468]), .B(n2767), .Z(n707) );
  NANDN U1030 ( .A(n2768), .B(n707), .Z(n708) );
  NAND U1031 ( .A(sreg[468]), .B(n2767), .Z(n709) );
  AND U1032 ( .A(n708), .B(n709), .Z(n2774) );
  NAND U1033 ( .A(n2788), .B(n2789), .Z(n710) );
  XOR U1034 ( .A(n2788), .B(n2789), .Z(n711) );
  NAND U1035 ( .A(n711), .B(sreg[471]), .Z(n712) );
  NAND U1036 ( .A(n710), .B(n712), .Z(n2795) );
  NAND U1037 ( .A(n2809), .B(n2810), .Z(n713) );
  XOR U1038 ( .A(n2809), .B(n2810), .Z(n714) );
  NAND U1039 ( .A(n714), .B(sreg[474]), .Z(n715) );
  NAND U1040 ( .A(n713), .B(n715), .Z(n2816) );
  NAND U1041 ( .A(n2830), .B(n2831), .Z(n716) );
  XOR U1042 ( .A(n2830), .B(n2831), .Z(n717) );
  NANDN U1043 ( .A(sreg[477]), .B(n717), .Z(n718) );
  NAND U1044 ( .A(n716), .B(n718), .Z(n2837) );
  NAND U1045 ( .A(sreg[480]), .B(n2852), .Z(n719) );
  XOR U1046 ( .A(sreg[480]), .B(n2852), .Z(n720) );
  NANDN U1047 ( .A(n2851), .B(n720), .Z(n721) );
  NAND U1048 ( .A(n719), .B(n721), .Z(n2858) );
  NAND U1049 ( .A(sreg[483]), .B(n2873), .Z(n722) );
  XOR U1050 ( .A(sreg[483]), .B(n2873), .Z(n723) );
  NANDN U1051 ( .A(n2872), .B(n723), .Z(n724) );
  NAND U1052 ( .A(n722), .B(n724), .Z(n2879) );
  NAND U1053 ( .A(n2893), .B(n2894), .Z(n725) );
  XOR U1054 ( .A(n2893), .B(n2894), .Z(n726) );
  NANDN U1055 ( .A(sreg[486]), .B(n726), .Z(n727) );
  NAND U1056 ( .A(n725), .B(n727), .Z(n2900) );
  NAND U1057 ( .A(n2914), .B(n2915), .Z(n728) );
  XOR U1058 ( .A(n2914), .B(n2915), .Z(n729) );
  NAND U1059 ( .A(n729), .B(sreg[489]), .Z(n730) );
  NAND U1060 ( .A(n728), .B(n730), .Z(n2921) );
  NAND U1061 ( .A(n2935), .B(n2936), .Z(n731) );
  XOR U1062 ( .A(n2935), .B(n2936), .Z(n732) );
  NAND U1063 ( .A(n732), .B(sreg[492]), .Z(n733) );
  NAND U1064 ( .A(n731), .B(n733), .Z(n2942) );
  NAND U1065 ( .A(n2956), .B(n2957), .Z(n734) );
  XOR U1066 ( .A(n2956), .B(n2957), .Z(n735) );
  NAND U1067 ( .A(n735), .B(sreg[495]), .Z(n736) );
  NAND U1068 ( .A(n734), .B(n736), .Z(n2963) );
  XOR U1069 ( .A(sreg[498]), .B(n2977), .Z(n737) );
  NANDN U1070 ( .A(n2978), .B(n737), .Z(n738) );
  NAND U1071 ( .A(sreg[498]), .B(n2977), .Z(n739) );
  AND U1072 ( .A(n738), .B(n739), .Z(n2984) );
  NAND U1073 ( .A(sreg[501]), .B(n2999), .Z(n740) );
  XOR U1074 ( .A(sreg[501]), .B(n2999), .Z(n741) );
  NANDN U1075 ( .A(n2998), .B(n741), .Z(n742) );
  NAND U1076 ( .A(n740), .B(n742), .Z(n3005) );
  NAND U1077 ( .A(n3019), .B(n3020), .Z(n743) );
  XOR U1078 ( .A(n3019), .B(n3020), .Z(n744) );
  NAND U1079 ( .A(n744), .B(sreg[504]), .Z(n745) );
  NAND U1080 ( .A(n743), .B(n745), .Z(n3026) );
  XOR U1081 ( .A(sreg[507]), .B(n3040), .Z(n746) );
  NANDN U1082 ( .A(n3041), .B(n746), .Z(n747) );
  NAND U1083 ( .A(sreg[507]), .B(n3040), .Z(n748) );
  AND U1084 ( .A(n747), .B(n748), .Z(n3048) );
  NAND U1085 ( .A(n1264), .B(n1263), .Z(n749) );
  XOR U1086 ( .A(n1264), .B(n1263), .Z(n750) );
  NANDN U1087 ( .A(sreg[255]), .B(n750), .Z(n751) );
  NAND U1088 ( .A(n749), .B(n751), .Z(n1268) );
  XOR U1089 ( .A(sreg[258]), .B(n1294), .Z(n752) );
  NANDN U1090 ( .A(n1295), .B(n752), .Z(n753) );
  NAND U1091 ( .A(sreg[258]), .B(n1294), .Z(n754) );
  AND U1092 ( .A(n753), .B(n754), .Z(n1297) );
  NAND U1093 ( .A(sreg[262]), .B(n1326), .Z(n755) );
  XOR U1094 ( .A(sreg[262]), .B(n1326), .Z(n756) );
  NANDN U1095 ( .A(n1325), .B(n756), .Z(n757) );
  NAND U1096 ( .A(n755), .B(n757), .Z(n1332) );
  NAND U1097 ( .A(sreg[265]), .B(n1347), .Z(n758) );
  XOR U1098 ( .A(sreg[265]), .B(n1347), .Z(n759) );
  NANDN U1099 ( .A(n1346), .B(n759), .Z(n760) );
  NAND U1100 ( .A(n758), .B(n760), .Z(n1353) );
  NAND U1101 ( .A(sreg[268]), .B(n1368), .Z(n761) );
  XOR U1102 ( .A(sreg[268]), .B(n1368), .Z(n762) );
  NANDN U1103 ( .A(n1367), .B(n762), .Z(n763) );
  NAND U1104 ( .A(n761), .B(n763), .Z(n1374) );
  NAND U1105 ( .A(n1388), .B(n1389), .Z(n764) );
  XOR U1106 ( .A(n1388), .B(n1389), .Z(n765) );
  NANDN U1107 ( .A(sreg[271]), .B(n765), .Z(n766) );
  NAND U1108 ( .A(n764), .B(n766), .Z(n1395) );
  XOR U1109 ( .A(sreg[274]), .B(n1409), .Z(n767) );
  NANDN U1110 ( .A(n1410), .B(n767), .Z(n768) );
  NAND U1111 ( .A(sreg[274]), .B(n1409), .Z(n769) );
  AND U1112 ( .A(n768), .B(n769), .Z(n1416) );
  NAND U1113 ( .A(sreg[277]), .B(n1431), .Z(n770) );
  XOR U1114 ( .A(sreg[277]), .B(n1431), .Z(n771) );
  NANDN U1115 ( .A(n1430), .B(n771), .Z(n772) );
  NAND U1116 ( .A(n770), .B(n772), .Z(n1437) );
  NAND U1117 ( .A(n1451), .B(n1452), .Z(n773) );
  XOR U1118 ( .A(n1451), .B(n1452), .Z(n774) );
  NAND U1119 ( .A(n774), .B(sreg[280]), .Z(n775) );
  NAND U1120 ( .A(n773), .B(n775), .Z(n1458) );
  XOR U1121 ( .A(sreg[283]), .B(n1472), .Z(n776) );
  NANDN U1122 ( .A(n1473), .B(n776), .Z(n777) );
  NAND U1123 ( .A(sreg[283]), .B(n1472), .Z(n778) );
  AND U1124 ( .A(n777), .B(n778), .Z(n1479) );
  NAND U1125 ( .A(sreg[286]), .B(n1494), .Z(n779) );
  XOR U1126 ( .A(sreg[286]), .B(n1494), .Z(n780) );
  NANDN U1127 ( .A(n1493), .B(n780), .Z(n781) );
  NAND U1128 ( .A(n779), .B(n781), .Z(n1500) );
  XOR U1129 ( .A(sreg[289]), .B(n1514), .Z(n782) );
  NANDN U1130 ( .A(n1515), .B(n782), .Z(n783) );
  NAND U1131 ( .A(sreg[289]), .B(n1514), .Z(n784) );
  AND U1132 ( .A(n783), .B(n784), .Z(n1521) );
  NAND U1133 ( .A(n1535), .B(n1536), .Z(n785) );
  XOR U1134 ( .A(n1535), .B(n1536), .Z(n786) );
  NAND U1135 ( .A(n786), .B(sreg[292]), .Z(n787) );
  NAND U1136 ( .A(n785), .B(n787), .Z(n1542) );
  XOR U1137 ( .A(sreg[295]), .B(n1556), .Z(n788) );
  NANDN U1138 ( .A(n1557), .B(n788), .Z(n789) );
  NAND U1139 ( .A(sreg[295]), .B(n1556), .Z(n790) );
  AND U1140 ( .A(n789), .B(n790), .Z(n1563) );
  NAND U1141 ( .A(n1577), .B(n1578), .Z(n791) );
  XOR U1142 ( .A(n1577), .B(n1578), .Z(n792) );
  NAND U1143 ( .A(n792), .B(sreg[298]), .Z(n793) );
  NAND U1144 ( .A(n791), .B(n793), .Z(n1584) );
  XOR U1145 ( .A(sreg[301]), .B(n1598), .Z(n794) );
  NANDN U1146 ( .A(n1599), .B(n794), .Z(n795) );
  NAND U1147 ( .A(sreg[301]), .B(n1598), .Z(n796) );
  AND U1148 ( .A(n795), .B(n796), .Z(n1605) );
  NAND U1149 ( .A(n1619), .B(n1620), .Z(n797) );
  XOR U1150 ( .A(n1619), .B(n1620), .Z(n798) );
  NAND U1151 ( .A(n798), .B(sreg[304]), .Z(n799) );
  NAND U1152 ( .A(n797), .B(n799), .Z(n1626) );
  NAND U1153 ( .A(sreg[307]), .B(n1641), .Z(n800) );
  XOR U1154 ( .A(sreg[307]), .B(n1641), .Z(n801) );
  NANDN U1155 ( .A(n1640), .B(n801), .Z(n802) );
  NAND U1156 ( .A(n800), .B(n802), .Z(n1647) );
  XOR U1157 ( .A(sreg[310]), .B(n1661), .Z(n803) );
  NANDN U1158 ( .A(n1662), .B(n803), .Z(n804) );
  NAND U1159 ( .A(sreg[310]), .B(n1661), .Z(n805) );
  AND U1160 ( .A(n804), .B(n805), .Z(n1668) );
  NAND U1161 ( .A(sreg[313]), .B(n1683), .Z(n806) );
  XOR U1162 ( .A(sreg[313]), .B(n1683), .Z(n807) );
  NANDN U1163 ( .A(n1682), .B(n807), .Z(n808) );
  NAND U1164 ( .A(n806), .B(n808), .Z(n1689) );
  NAND U1165 ( .A(n1703), .B(n1704), .Z(n809) );
  XOR U1166 ( .A(n1703), .B(n1704), .Z(n810) );
  NAND U1167 ( .A(n810), .B(sreg[316]), .Z(n811) );
  NAND U1168 ( .A(n809), .B(n811), .Z(n1710) );
  XOR U1169 ( .A(sreg[319]), .B(n1724), .Z(n812) );
  NANDN U1170 ( .A(n1725), .B(n812), .Z(n813) );
  NAND U1171 ( .A(sreg[319]), .B(n1724), .Z(n814) );
  AND U1172 ( .A(n813), .B(n814), .Z(n1731) );
  NAND U1173 ( .A(sreg[322]), .B(n1746), .Z(n815) );
  XOR U1174 ( .A(sreg[322]), .B(n1746), .Z(n816) );
  NANDN U1175 ( .A(n1745), .B(n816), .Z(n817) );
  NAND U1176 ( .A(n815), .B(n817), .Z(n1752) );
  XOR U1177 ( .A(sreg[325]), .B(n1766), .Z(n818) );
  NANDN U1178 ( .A(n1767), .B(n818), .Z(n819) );
  NAND U1179 ( .A(sreg[325]), .B(n1766), .Z(n820) );
  AND U1180 ( .A(n819), .B(n820), .Z(n1773) );
  NAND U1181 ( .A(n1787), .B(n1788), .Z(n821) );
  XOR U1182 ( .A(n1787), .B(n1788), .Z(n822) );
  NAND U1183 ( .A(n822), .B(sreg[328]), .Z(n823) );
  NAND U1184 ( .A(n821), .B(n823), .Z(n1794) );
  NAND U1185 ( .A(n1808), .B(n1809), .Z(n824) );
  XOR U1186 ( .A(n1808), .B(n1809), .Z(n825) );
  NAND U1187 ( .A(n825), .B(sreg[331]), .Z(n826) );
  NAND U1188 ( .A(n824), .B(n826), .Z(n1815) );
  NAND U1189 ( .A(sreg[334]), .B(n1830), .Z(n827) );
  XOR U1190 ( .A(sreg[334]), .B(n1830), .Z(n828) );
  NANDN U1191 ( .A(n1829), .B(n828), .Z(n829) );
  NAND U1192 ( .A(n827), .B(n829), .Z(n1836) );
  NAND U1193 ( .A(n1850), .B(n1851), .Z(n830) );
  XOR U1194 ( .A(n1850), .B(n1851), .Z(n831) );
  NAND U1195 ( .A(n831), .B(sreg[337]), .Z(n832) );
  NAND U1196 ( .A(n830), .B(n832), .Z(n1857) );
  XOR U1197 ( .A(sreg[340]), .B(n1871), .Z(n833) );
  NANDN U1198 ( .A(n1872), .B(n833), .Z(n834) );
  NAND U1199 ( .A(sreg[340]), .B(n1871), .Z(n835) );
  AND U1200 ( .A(n834), .B(n835), .Z(n1878) );
  NAND U1201 ( .A(sreg[343]), .B(n1893), .Z(n836) );
  XOR U1202 ( .A(sreg[343]), .B(n1893), .Z(n837) );
  NANDN U1203 ( .A(n1892), .B(n837), .Z(n838) );
  NAND U1204 ( .A(n836), .B(n838), .Z(n1899) );
  NAND U1205 ( .A(n1913), .B(n1914), .Z(n839) );
  XOR U1206 ( .A(n1913), .B(n1914), .Z(n840) );
  NAND U1207 ( .A(n840), .B(sreg[346]), .Z(n841) );
  NAND U1208 ( .A(n839), .B(n841), .Z(n1920) );
  XOR U1209 ( .A(sreg[349]), .B(n1934), .Z(n842) );
  NANDN U1210 ( .A(n1935), .B(n842), .Z(n843) );
  NAND U1211 ( .A(sreg[349]), .B(n1934), .Z(n844) );
  AND U1212 ( .A(n843), .B(n844), .Z(n1941) );
  NAND U1213 ( .A(sreg[352]), .B(n1956), .Z(n845) );
  XOR U1214 ( .A(sreg[352]), .B(n1956), .Z(n846) );
  NANDN U1215 ( .A(n1955), .B(n846), .Z(n847) );
  NAND U1216 ( .A(n845), .B(n847), .Z(n1962) );
  NAND U1217 ( .A(n1976), .B(n1977), .Z(n848) );
  XOR U1218 ( .A(n1976), .B(n1977), .Z(n849) );
  NAND U1219 ( .A(n849), .B(sreg[355]), .Z(n850) );
  NAND U1220 ( .A(n848), .B(n850), .Z(n1983) );
  XOR U1221 ( .A(sreg[358]), .B(n1997), .Z(n851) );
  NANDN U1222 ( .A(n1998), .B(n851), .Z(n852) );
  NAND U1223 ( .A(sreg[358]), .B(n1997), .Z(n853) );
  AND U1224 ( .A(n852), .B(n853), .Z(n2004) );
  NAND U1225 ( .A(n2018), .B(n2019), .Z(n854) );
  XOR U1226 ( .A(n2018), .B(n2019), .Z(n855) );
  NAND U1227 ( .A(n855), .B(sreg[361]), .Z(n856) );
  NAND U1228 ( .A(n854), .B(n856), .Z(n2025) );
  NAND U1229 ( .A(sreg[364]), .B(n2040), .Z(n857) );
  XOR U1230 ( .A(sreg[364]), .B(n2040), .Z(n858) );
  NANDN U1231 ( .A(n2039), .B(n858), .Z(n859) );
  NAND U1232 ( .A(n857), .B(n859), .Z(n2046) );
  NAND U1233 ( .A(sreg[367]), .B(n2061), .Z(n860) );
  XOR U1234 ( .A(sreg[367]), .B(n2061), .Z(n861) );
  NANDN U1235 ( .A(n2060), .B(n861), .Z(n862) );
  NAND U1236 ( .A(n860), .B(n862), .Z(n2067) );
  XOR U1237 ( .A(sreg[370]), .B(n2081), .Z(n863) );
  NANDN U1238 ( .A(n2082), .B(n863), .Z(n864) );
  NAND U1239 ( .A(sreg[370]), .B(n2081), .Z(n865) );
  AND U1240 ( .A(n864), .B(n865), .Z(n2088) );
  NAND U1241 ( .A(n2102), .B(n2103), .Z(n866) );
  XOR U1242 ( .A(n2102), .B(n2103), .Z(n867) );
  NAND U1243 ( .A(n867), .B(sreg[373]), .Z(n868) );
  NAND U1244 ( .A(n866), .B(n868), .Z(n2109) );
  NAND U1245 ( .A(n2123), .B(n2124), .Z(n869) );
  XOR U1246 ( .A(n2123), .B(n2124), .Z(n870) );
  NAND U1247 ( .A(n870), .B(sreg[376]), .Z(n871) );
  NAND U1248 ( .A(n869), .B(n871), .Z(n2130) );
  XOR U1249 ( .A(sreg[379]), .B(n2144), .Z(n872) );
  NANDN U1250 ( .A(n2145), .B(n872), .Z(n873) );
  NAND U1251 ( .A(sreg[379]), .B(n2144), .Z(n874) );
  AND U1252 ( .A(n873), .B(n874), .Z(n2151) );
  NAND U1253 ( .A(sreg[382]), .B(n2166), .Z(n875) );
  XOR U1254 ( .A(sreg[382]), .B(n2166), .Z(n876) );
  NANDN U1255 ( .A(n2165), .B(n876), .Z(n877) );
  NAND U1256 ( .A(n875), .B(n877), .Z(n2172) );
  XOR U1257 ( .A(sreg[385]), .B(n2186), .Z(n878) );
  NANDN U1258 ( .A(n2187), .B(n878), .Z(n879) );
  NAND U1259 ( .A(sreg[385]), .B(n2186), .Z(n880) );
  AND U1260 ( .A(n879), .B(n880), .Z(n2193) );
  NAND U1261 ( .A(sreg[388]), .B(n2208), .Z(n881) );
  XOR U1262 ( .A(sreg[388]), .B(n2208), .Z(n882) );
  NANDN U1263 ( .A(n2207), .B(n882), .Z(n883) );
  NAND U1264 ( .A(n881), .B(n883), .Z(n2214) );
  XOR U1265 ( .A(sreg[391]), .B(n2228), .Z(n884) );
  NANDN U1266 ( .A(n2229), .B(n884), .Z(n885) );
  NAND U1267 ( .A(sreg[391]), .B(n2228), .Z(n886) );
  AND U1268 ( .A(n885), .B(n886), .Z(n2235) );
  NAND U1269 ( .A(n2249), .B(n2250), .Z(n887) );
  XOR U1270 ( .A(n2249), .B(n2250), .Z(n888) );
  NAND U1271 ( .A(n888), .B(sreg[394]), .Z(n889) );
  NAND U1272 ( .A(n887), .B(n889), .Z(n2256) );
  XOR U1273 ( .A(sreg[397]), .B(n2270), .Z(n890) );
  NANDN U1274 ( .A(n2271), .B(n890), .Z(n891) );
  NAND U1275 ( .A(sreg[397]), .B(n2270), .Z(n892) );
  AND U1276 ( .A(n891), .B(n892), .Z(n2277) );
  NAND U1277 ( .A(sreg[400]), .B(n2292), .Z(n893) );
  XOR U1278 ( .A(sreg[400]), .B(n2292), .Z(n894) );
  NANDN U1279 ( .A(n2291), .B(n894), .Z(n895) );
  NAND U1280 ( .A(n893), .B(n895), .Z(n2298) );
  NAND U1281 ( .A(sreg[403]), .B(n2313), .Z(n896) );
  XOR U1282 ( .A(sreg[403]), .B(n2313), .Z(n897) );
  NANDN U1283 ( .A(n2312), .B(n897), .Z(n898) );
  NAND U1284 ( .A(n896), .B(n898), .Z(n2319) );
  NAND U1285 ( .A(n2333), .B(n2334), .Z(n899) );
  XOR U1286 ( .A(n2333), .B(n2334), .Z(n900) );
  NANDN U1287 ( .A(sreg[406]), .B(n900), .Z(n901) );
  NAND U1288 ( .A(n899), .B(n901), .Z(n2340) );
  NAND U1289 ( .A(n2354), .B(n2355), .Z(n902) );
  XOR U1290 ( .A(n2354), .B(n2355), .Z(n903) );
  NAND U1291 ( .A(n903), .B(sreg[409]), .Z(n904) );
  NAND U1292 ( .A(n902), .B(n904), .Z(n2361) );
  NAND U1293 ( .A(n2375), .B(n2376), .Z(n905) );
  XOR U1294 ( .A(n2375), .B(n2376), .Z(n906) );
  NAND U1295 ( .A(n906), .B(sreg[412]), .Z(n907) );
  NAND U1296 ( .A(n905), .B(n907), .Z(n2382) );
  XOR U1297 ( .A(sreg[415]), .B(n2396), .Z(n908) );
  NANDN U1298 ( .A(n2397), .B(n908), .Z(n909) );
  NAND U1299 ( .A(sreg[415]), .B(n2396), .Z(n910) );
  AND U1300 ( .A(n909), .B(n910), .Z(n2403) );
  NAND U1301 ( .A(sreg[418]), .B(n2418), .Z(n911) );
  XOR U1302 ( .A(sreg[418]), .B(n2418), .Z(n912) );
  NANDN U1303 ( .A(n2417), .B(n912), .Z(n913) );
  NAND U1304 ( .A(n911), .B(n913), .Z(n2424) );
  NAND U1305 ( .A(n2438), .B(n2439), .Z(n914) );
  XOR U1306 ( .A(n2438), .B(n2439), .Z(n915) );
  NAND U1307 ( .A(n915), .B(sreg[421]), .Z(n916) );
  NAND U1308 ( .A(n914), .B(n916), .Z(n2445) );
  NAND U1309 ( .A(n2459), .B(n2460), .Z(n917) );
  XOR U1310 ( .A(n2459), .B(n2460), .Z(n918) );
  NAND U1311 ( .A(n918), .B(sreg[424]), .Z(n919) );
  NAND U1312 ( .A(n917), .B(n919), .Z(n2466) );
  XOR U1313 ( .A(sreg[427]), .B(n2480), .Z(n920) );
  NANDN U1314 ( .A(n2481), .B(n920), .Z(n921) );
  NAND U1315 ( .A(sreg[427]), .B(n2480), .Z(n922) );
  AND U1316 ( .A(n921), .B(n922), .Z(n2487) );
  NAND U1317 ( .A(sreg[430]), .B(n2502), .Z(n923) );
  XOR U1318 ( .A(sreg[430]), .B(n2502), .Z(n924) );
  NANDN U1319 ( .A(n2501), .B(n924), .Z(n925) );
  NAND U1320 ( .A(n923), .B(n925), .Z(n2508) );
  NAND U1321 ( .A(n2522), .B(n2523), .Z(n926) );
  XOR U1322 ( .A(n2522), .B(n2523), .Z(n927) );
  NAND U1323 ( .A(n927), .B(sreg[433]), .Z(n928) );
  NAND U1324 ( .A(n926), .B(n928), .Z(n2529) );
  NAND U1325 ( .A(n2543), .B(n2544), .Z(n929) );
  XOR U1326 ( .A(n2543), .B(n2544), .Z(n930) );
  NANDN U1327 ( .A(sreg[436]), .B(n930), .Z(n931) );
  NAND U1328 ( .A(n929), .B(n931), .Z(n2550) );
  NAND U1329 ( .A(sreg[439]), .B(n2565), .Z(n932) );
  XOR U1330 ( .A(sreg[439]), .B(n2565), .Z(n933) );
  NANDN U1331 ( .A(n2564), .B(n933), .Z(n934) );
  NAND U1332 ( .A(n932), .B(n934), .Z(n2571) );
  NAND U1333 ( .A(n2585), .B(n2586), .Z(n935) );
  XOR U1334 ( .A(n2585), .B(n2586), .Z(n936) );
  NAND U1335 ( .A(n936), .B(sreg[442]), .Z(n937) );
  NAND U1336 ( .A(n935), .B(n937), .Z(n2592) );
  XOR U1337 ( .A(sreg[445]), .B(n2606), .Z(n938) );
  NANDN U1338 ( .A(n2607), .B(n938), .Z(n939) );
  NAND U1339 ( .A(sreg[445]), .B(n2606), .Z(n940) );
  AND U1340 ( .A(n939), .B(n940), .Z(n2613) );
  NAND U1341 ( .A(sreg[448]), .B(n2628), .Z(n941) );
  XOR U1342 ( .A(sreg[448]), .B(n2628), .Z(n942) );
  NANDN U1343 ( .A(n2627), .B(n942), .Z(n943) );
  NAND U1344 ( .A(n941), .B(n943), .Z(n2634) );
  NAND U1345 ( .A(n2648), .B(n2649), .Z(n944) );
  XOR U1346 ( .A(n2648), .B(n2649), .Z(n945) );
  NAND U1347 ( .A(n945), .B(sreg[451]), .Z(n946) );
  NAND U1348 ( .A(n944), .B(n946), .Z(n2655) );
  NAND U1349 ( .A(sreg[454]), .B(n2670), .Z(n947) );
  XOR U1350 ( .A(sreg[454]), .B(n2670), .Z(n948) );
  NANDN U1351 ( .A(n2669), .B(n948), .Z(n949) );
  NAND U1352 ( .A(n947), .B(n949), .Z(n2676) );
  NAND U1353 ( .A(n2690), .B(n2691), .Z(n950) );
  XOR U1354 ( .A(n2690), .B(n2691), .Z(n951) );
  NAND U1355 ( .A(n951), .B(sreg[457]), .Z(n952) );
  NAND U1356 ( .A(n950), .B(n952), .Z(n2697) );
  NAND U1357 ( .A(sreg[460]), .B(n2712), .Z(n953) );
  XOR U1358 ( .A(sreg[460]), .B(n2712), .Z(n954) );
  NANDN U1359 ( .A(n2711), .B(n954), .Z(n955) );
  NAND U1360 ( .A(n953), .B(n955), .Z(n2718) );
  NAND U1361 ( .A(n2732), .B(n2733), .Z(n956) );
  XOR U1362 ( .A(n2732), .B(n2733), .Z(n957) );
  NAND U1363 ( .A(n957), .B(sreg[463]), .Z(n958) );
  NAND U1364 ( .A(n956), .B(n958), .Z(n2739) );
  XOR U1365 ( .A(sreg[466]), .B(n2753), .Z(n959) );
  NANDN U1366 ( .A(n2754), .B(n959), .Z(n960) );
  NAND U1367 ( .A(sreg[466]), .B(n2753), .Z(n961) );
  AND U1368 ( .A(n960), .B(n961), .Z(n2760) );
  NAND U1369 ( .A(sreg[469]), .B(n2775), .Z(n962) );
  XOR U1370 ( .A(sreg[469]), .B(n2775), .Z(n963) );
  NANDN U1371 ( .A(n2774), .B(n963), .Z(n964) );
  NAND U1372 ( .A(n962), .B(n964), .Z(n2781) );
  NAND U1373 ( .A(n2795), .B(n2796), .Z(n965) );
  XOR U1374 ( .A(n2795), .B(n2796), .Z(n966) );
  NAND U1375 ( .A(n966), .B(sreg[472]), .Z(n967) );
  NAND U1376 ( .A(n965), .B(n967), .Z(n2802) );
  XOR U1377 ( .A(sreg[475]), .B(n2816), .Z(n968) );
  NANDN U1378 ( .A(n2817), .B(n968), .Z(n969) );
  NAND U1379 ( .A(sreg[475]), .B(n2816), .Z(n970) );
  AND U1380 ( .A(n969), .B(n970), .Z(n2823) );
  NAND U1381 ( .A(sreg[478]), .B(n2838), .Z(n971) );
  XOR U1382 ( .A(sreg[478]), .B(n2838), .Z(n972) );
  NANDN U1383 ( .A(n2837), .B(n972), .Z(n973) );
  NAND U1384 ( .A(n971), .B(n973), .Z(n2844) );
  NAND U1385 ( .A(n2858), .B(n2859), .Z(n974) );
  XOR U1386 ( .A(n2858), .B(n2859), .Z(n975) );
  NAND U1387 ( .A(n975), .B(sreg[481]), .Z(n976) );
  NAND U1388 ( .A(n974), .B(n976), .Z(n2865) );
  NAND U1389 ( .A(n2879), .B(n2880), .Z(n977) );
  XOR U1390 ( .A(n2879), .B(n2880), .Z(n978) );
  NAND U1391 ( .A(n978), .B(sreg[484]), .Z(n979) );
  NAND U1392 ( .A(n977), .B(n979), .Z(n2886) );
  NAND U1393 ( .A(n2900), .B(n2901), .Z(n980) );
  XOR U1394 ( .A(n2900), .B(n2901), .Z(n981) );
  NANDN U1395 ( .A(sreg[487]), .B(n981), .Z(n982) );
  NAND U1396 ( .A(n980), .B(n982), .Z(n2907) );
  NAND U1397 ( .A(n2921), .B(n2922), .Z(n983) );
  XOR U1398 ( .A(n2921), .B(n2922), .Z(n984) );
  NAND U1399 ( .A(n984), .B(sreg[490]), .Z(n985) );
  NAND U1400 ( .A(n983), .B(n985), .Z(n2928) );
  XOR U1401 ( .A(sreg[493]), .B(n2942), .Z(n986) );
  NANDN U1402 ( .A(n2943), .B(n986), .Z(n987) );
  NAND U1403 ( .A(sreg[493]), .B(n2942), .Z(n988) );
  AND U1404 ( .A(n987), .B(n988), .Z(n2949) );
  NAND U1405 ( .A(n2963), .B(n2964), .Z(n989) );
  XOR U1406 ( .A(n2963), .B(n2964), .Z(n990) );
  NAND U1407 ( .A(n990), .B(sreg[496]), .Z(n991) );
  NAND U1408 ( .A(n989), .B(n991), .Z(n2970) );
  NAND U1409 ( .A(sreg[499]), .B(n2985), .Z(n992) );
  XOR U1410 ( .A(sreg[499]), .B(n2985), .Z(n993) );
  NANDN U1411 ( .A(n2984), .B(n993), .Z(n994) );
  NAND U1412 ( .A(n992), .B(n994), .Z(n2991) );
  XOR U1413 ( .A(sreg[502]), .B(n3005), .Z(n995) );
  NANDN U1414 ( .A(n3006), .B(n995), .Z(n996) );
  NAND U1415 ( .A(sreg[502]), .B(n3005), .Z(n997) );
  AND U1416 ( .A(n996), .B(n997), .Z(n3012) );
  NAND U1417 ( .A(n3026), .B(n3027), .Z(n998) );
  XOR U1418 ( .A(n3026), .B(n3027), .Z(n999) );
  NAND U1419 ( .A(n999), .B(sreg[505]), .Z(n1000) );
  NAND U1420 ( .A(n998), .B(n1000), .Z(n3033) );
  NAND U1421 ( .A(sreg[508]), .B(n3049), .Z(n1001) );
  XOR U1422 ( .A(sreg[508]), .B(n3049), .Z(n1002) );
  NANDN U1423 ( .A(n3048), .B(n1002), .Z(n1003) );
  NAND U1424 ( .A(n1001), .B(n1003), .Z(n3051) );
  NAND U1425 ( .A(n1307), .B(n1306), .Z(n1004) );
  NANDN U1426 ( .A(n1304), .B(n1305), .Z(n1005) );
  AND U1427 ( .A(n1004), .B(n1005), .Z(n1316) );
  NANDN U1428 ( .A(n1266), .B(sreg[256]), .Z(n1006) );
  NANDN U1429 ( .A(n1268), .B(n1267), .Z(n1007) );
  NAND U1430 ( .A(n1006), .B(n1007), .Z(n1283) );
  NAND U1431 ( .A(n1297), .B(n1298), .Z(n1008) );
  XOR U1432 ( .A(n1297), .B(n1298), .Z(n1009) );
  NANDN U1433 ( .A(sreg[259]), .B(n1009), .Z(n1010) );
  NAND U1434 ( .A(n1008), .B(n1010), .Z(n1309) );
  NAND U1435 ( .A(n1332), .B(n1333), .Z(n1011) );
  XOR U1436 ( .A(n1332), .B(n1333), .Z(n1012) );
  NAND U1437 ( .A(n1012), .B(sreg[263]), .Z(n1013) );
  NAND U1438 ( .A(n1011), .B(n1013), .Z(n1339) );
  NAND U1439 ( .A(n1353), .B(n1354), .Z(n1014) );
  XOR U1440 ( .A(n1353), .B(n1354), .Z(n1015) );
  NAND U1441 ( .A(n1015), .B(sreg[266]), .Z(n1016) );
  NAND U1442 ( .A(n1014), .B(n1016), .Z(n1360) );
  XOR U1443 ( .A(sreg[269]), .B(n1374), .Z(n1017) );
  NANDN U1444 ( .A(n1375), .B(n1017), .Z(n1018) );
  NAND U1445 ( .A(sreg[269]), .B(n1374), .Z(n1019) );
  AND U1446 ( .A(n1018), .B(n1019), .Z(n1381) );
  NAND U1447 ( .A(sreg[272]), .B(n1396), .Z(n1020) );
  XOR U1448 ( .A(sreg[272]), .B(n1396), .Z(n1021) );
  NANDN U1449 ( .A(n1395), .B(n1021), .Z(n1022) );
  NAND U1450 ( .A(n1020), .B(n1022), .Z(n1402) );
  NAND U1451 ( .A(sreg[275]), .B(n1417), .Z(n1023) );
  XOR U1452 ( .A(sreg[275]), .B(n1417), .Z(n1024) );
  NANDN U1453 ( .A(n1416), .B(n1024), .Z(n1025) );
  NAND U1454 ( .A(n1023), .B(n1025), .Z(n1423) );
  XOR U1455 ( .A(sreg[278]), .B(n1437), .Z(n1026) );
  NANDN U1456 ( .A(n1438), .B(n1026), .Z(n1027) );
  NAND U1457 ( .A(sreg[278]), .B(n1437), .Z(n1028) );
  AND U1458 ( .A(n1027), .B(n1028), .Z(n1444) );
  NAND U1459 ( .A(n1458), .B(n1459), .Z(n1029) );
  XOR U1460 ( .A(n1458), .B(n1459), .Z(n1030) );
  NAND U1461 ( .A(n1030), .B(sreg[281]), .Z(n1031) );
  NAND U1462 ( .A(n1029), .B(n1031), .Z(n1466) );
  NAND U1463 ( .A(sreg[284]), .B(n1480), .Z(n1032) );
  XOR U1464 ( .A(sreg[284]), .B(n1480), .Z(n1033) );
  NANDN U1465 ( .A(n1479), .B(n1033), .Z(n1034) );
  NAND U1466 ( .A(n1032), .B(n1034), .Z(n1486) );
  XOR U1467 ( .A(sreg[287]), .B(n1500), .Z(n1035) );
  NANDN U1468 ( .A(n1501), .B(n1035), .Z(n1036) );
  NAND U1469 ( .A(sreg[287]), .B(n1500), .Z(n1037) );
  AND U1470 ( .A(n1036), .B(n1037), .Z(n1507) );
  NAND U1471 ( .A(n1521), .B(n1522), .Z(n1038) );
  XOR U1472 ( .A(n1521), .B(n1522), .Z(n1039) );
  NANDN U1473 ( .A(sreg[290]), .B(n1039), .Z(n1040) );
  NAND U1474 ( .A(n1038), .B(n1040), .Z(n1528) );
  NAND U1475 ( .A(n1542), .B(n1543), .Z(n1041) );
  XOR U1476 ( .A(n1542), .B(n1543), .Z(n1042) );
  NAND U1477 ( .A(n1042), .B(sreg[293]), .Z(n1043) );
  NAND U1478 ( .A(n1041), .B(n1043), .Z(n1549) );
  NAND U1479 ( .A(sreg[296]), .B(n1564), .Z(n1044) );
  XOR U1480 ( .A(sreg[296]), .B(n1564), .Z(n1045) );
  NANDN U1481 ( .A(n1563), .B(n1045), .Z(n1046) );
  NAND U1482 ( .A(n1044), .B(n1046), .Z(n1570) );
  XOR U1483 ( .A(sreg[299]), .B(n1584), .Z(n1047) );
  NANDN U1484 ( .A(n1585), .B(n1047), .Z(n1048) );
  NAND U1485 ( .A(sreg[299]), .B(n1584), .Z(n1049) );
  AND U1486 ( .A(n1048), .B(n1049), .Z(n1591) );
  NAND U1487 ( .A(sreg[302]), .B(n1606), .Z(n1050) );
  XOR U1488 ( .A(sreg[302]), .B(n1606), .Z(n1051) );
  NANDN U1489 ( .A(n1605), .B(n1051), .Z(n1052) );
  NAND U1490 ( .A(n1050), .B(n1052), .Z(n1612) );
  NAND U1491 ( .A(n1626), .B(n1627), .Z(n1053) );
  XOR U1492 ( .A(n1626), .B(n1627), .Z(n1054) );
  NAND U1493 ( .A(n1054), .B(sreg[305]), .Z(n1055) );
  NAND U1494 ( .A(n1053), .B(n1055), .Z(n1633) );
  XOR U1495 ( .A(sreg[308]), .B(n1647), .Z(n1056) );
  NANDN U1496 ( .A(n1648), .B(n1056), .Z(n1057) );
  NAND U1497 ( .A(sreg[308]), .B(n1647), .Z(n1058) );
  AND U1498 ( .A(n1057), .B(n1058), .Z(n1654) );
  NAND U1499 ( .A(n1668), .B(n1669), .Z(n1059) );
  XOR U1500 ( .A(n1668), .B(n1669), .Z(n1060) );
  NANDN U1501 ( .A(sreg[311]), .B(n1060), .Z(n1061) );
  NAND U1502 ( .A(n1059), .B(n1061), .Z(n1675) );
  NAND U1503 ( .A(n1689), .B(n1690), .Z(n1062) );
  XOR U1504 ( .A(n1689), .B(n1690), .Z(n1063) );
  NAND U1505 ( .A(n1063), .B(sreg[314]), .Z(n1064) );
  NAND U1506 ( .A(n1062), .B(n1064), .Z(n1696) );
  XOR U1507 ( .A(sreg[317]), .B(n1710), .Z(n1065) );
  NANDN U1508 ( .A(n1711), .B(n1065), .Z(n1066) );
  NAND U1509 ( .A(sreg[317]), .B(n1710), .Z(n1067) );
  AND U1510 ( .A(n1066), .B(n1067), .Z(n1717) );
  NAND U1511 ( .A(sreg[320]), .B(n1732), .Z(n1068) );
  XOR U1512 ( .A(sreg[320]), .B(n1732), .Z(n1069) );
  NANDN U1513 ( .A(n1731), .B(n1069), .Z(n1070) );
  NAND U1514 ( .A(n1068), .B(n1070), .Z(n1738) );
  NAND U1515 ( .A(n1752), .B(n1753), .Z(n1071) );
  XOR U1516 ( .A(n1752), .B(n1753), .Z(n1072) );
  NAND U1517 ( .A(n1072), .B(sreg[323]), .Z(n1073) );
  NAND U1518 ( .A(n1071), .B(n1073), .Z(n1759) );
  NAND U1519 ( .A(sreg[326]), .B(n1774), .Z(n1074) );
  XOR U1520 ( .A(sreg[326]), .B(n1774), .Z(n1075) );
  NANDN U1521 ( .A(n1773), .B(n1075), .Z(n1076) );
  NAND U1522 ( .A(n1074), .B(n1076), .Z(n1780) );
  NAND U1523 ( .A(n1794), .B(n1795), .Z(n1077) );
  XOR U1524 ( .A(n1794), .B(n1795), .Z(n1078) );
  NAND U1525 ( .A(n1078), .B(sreg[329]), .Z(n1079) );
  NAND U1526 ( .A(n1077), .B(n1079), .Z(n1801) );
  NAND U1527 ( .A(n1815), .B(n1816), .Z(n1080) );
  XOR U1528 ( .A(n1815), .B(n1816), .Z(n1081) );
  NAND U1529 ( .A(n1081), .B(sreg[332]), .Z(n1082) );
  NAND U1530 ( .A(n1080), .B(n1082), .Z(n1822) );
  NAND U1531 ( .A(n1836), .B(n1837), .Z(n1083) );
  XOR U1532 ( .A(n1836), .B(n1837), .Z(n1084) );
  NAND U1533 ( .A(n1084), .B(sreg[335]), .Z(n1085) );
  NAND U1534 ( .A(n1083), .B(n1085), .Z(n1843) );
  XOR U1535 ( .A(sreg[338]), .B(n1857), .Z(n1086) );
  NANDN U1536 ( .A(n1858), .B(n1086), .Z(n1087) );
  NAND U1537 ( .A(sreg[338]), .B(n1857), .Z(n1088) );
  AND U1538 ( .A(n1087), .B(n1088), .Z(n1864) );
  NAND U1539 ( .A(sreg[341]), .B(n1879), .Z(n1089) );
  XOR U1540 ( .A(sreg[341]), .B(n1879), .Z(n1090) );
  NANDN U1541 ( .A(n1878), .B(n1090), .Z(n1091) );
  NAND U1542 ( .A(n1089), .B(n1091), .Z(n1885) );
  NAND U1543 ( .A(n1899), .B(n1900), .Z(n1092) );
  XOR U1544 ( .A(n1899), .B(n1900), .Z(n1093) );
  NAND U1545 ( .A(n1093), .B(sreg[344]), .Z(n1094) );
  NAND U1546 ( .A(n1092), .B(n1094), .Z(n1906) );
  XOR U1547 ( .A(sreg[347]), .B(n1920), .Z(n1095) );
  NANDN U1548 ( .A(n1921), .B(n1095), .Z(n1096) );
  NAND U1549 ( .A(sreg[347]), .B(n1920), .Z(n1097) );
  AND U1550 ( .A(n1096), .B(n1097), .Z(n1927) );
  NAND U1551 ( .A(sreg[350]), .B(n1942), .Z(n1098) );
  XOR U1552 ( .A(sreg[350]), .B(n1942), .Z(n1099) );
  NANDN U1553 ( .A(n1941), .B(n1099), .Z(n1100) );
  NAND U1554 ( .A(n1098), .B(n1100), .Z(n1948) );
  XOR U1555 ( .A(sreg[353]), .B(n1962), .Z(n1101) );
  NANDN U1556 ( .A(n1963), .B(n1101), .Z(n1102) );
  NAND U1557 ( .A(sreg[353]), .B(n1962), .Z(n1103) );
  AND U1558 ( .A(n1102), .B(n1103), .Z(n1969) );
  NAND U1559 ( .A(n1983), .B(n1984), .Z(n1104) );
  XOR U1560 ( .A(n1983), .B(n1984), .Z(n1105) );
  NAND U1561 ( .A(n1105), .B(sreg[356]), .Z(n1106) );
  NAND U1562 ( .A(n1104), .B(n1106), .Z(n1990) );
  NAND U1563 ( .A(n2004), .B(n2005), .Z(n1107) );
  XOR U1564 ( .A(n2004), .B(n2005), .Z(n1108) );
  NANDN U1565 ( .A(sreg[359]), .B(n1108), .Z(n1109) );
  NAND U1566 ( .A(n1107), .B(n1109), .Z(n2011) );
  NAND U1567 ( .A(n2025), .B(n2026), .Z(n1110) );
  XOR U1568 ( .A(n2025), .B(n2026), .Z(n1111) );
  NAND U1569 ( .A(n1111), .B(sreg[362]), .Z(n1112) );
  NAND U1570 ( .A(n1110), .B(n1112), .Z(n2032) );
  XOR U1571 ( .A(sreg[365]), .B(n2046), .Z(n1113) );
  NANDN U1572 ( .A(n2047), .B(n1113), .Z(n1114) );
  NAND U1573 ( .A(sreg[365]), .B(n2046), .Z(n1115) );
  AND U1574 ( .A(n1114), .B(n1115), .Z(n2053) );
  NAND U1575 ( .A(n2067), .B(n2068), .Z(n1116) );
  XOR U1576 ( .A(n2067), .B(n2068), .Z(n1117) );
  NAND U1577 ( .A(n1117), .B(sreg[368]), .Z(n1118) );
  NAND U1578 ( .A(n1116), .B(n1118), .Z(n2074) );
  NAND U1579 ( .A(sreg[371]), .B(n2089), .Z(n1119) );
  XOR U1580 ( .A(sreg[371]), .B(n2089), .Z(n1120) );
  NANDN U1581 ( .A(n2088), .B(n1120), .Z(n1121) );
  NAND U1582 ( .A(n1119), .B(n1121), .Z(n2095) );
  XOR U1583 ( .A(sreg[374]), .B(n2109), .Z(n1122) );
  NANDN U1584 ( .A(n2110), .B(n1122), .Z(n1123) );
  NAND U1585 ( .A(sreg[374]), .B(n2109), .Z(n1124) );
  AND U1586 ( .A(n1123), .B(n1124), .Z(n2116) );
  NAND U1587 ( .A(n2130), .B(n2131), .Z(n1125) );
  XOR U1588 ( .A(n2130), .B(n2131), .Z(n1126) );
  NAND U1589 ( .A(n1126), .B(sreg[377]), .Z(n1127) );
  NAND U1590 ( .A(n1125), .B(n1127), .Z(n2137) );
  NAND U1591 ( .A(sreg[380]), .B(n2152), .Z(n1128) );
  XOR U1592 ( .A(sreg[380]), .B(n2152), .Z(n1129) );
  NANDN U1593 ( .A(n2151), .B(n1129), .Z(n1130) );
  NAND U1594 ( .A(n1128), .B(n1130), .Z(n2158) );
  XOR U1595 ( .A(sreg[383]), .B(n2172), .Z(n1131) );
  NANDN U1596 ( .A(n2173), .B(n1131), .Z(n1132) );
  NAND U1597 ( .A(sreg[383]), .B(n2172), .Z(n1133) );
  AND U1598 ( .A(n1132), .B(n1133), .Z(n2179) );
  NAND U1599 ( .A(sreg[386]), .B(n2194), .Z(n1134) );
  XOR U1600 ( .A(sreg[386]), .B(n2194), .Z(n1135) );
  NANDN U1601 ( .A(n2193), .B(n1135), .Z(n1136) );
  NAND U1602 ( .A(n1134), .B(n1136), .Z(n2200) );
  NAND U1603 ( .A(n2214), .B(n2215), .Z(n1137) );
  XOR U1604 ( .A(n2214), .B(n2215), .Z(n1138) );
  NAND U1605 ( .A(n1138), .B(sreg[389]), .Z(n1139) );
  NAND U1606 ( .A(n1137), .B(n1139), .Z(n2221) );
  NAND U1607 ( .A(sreg[392]), .B(n2236), .Z(n1140) );
  XOR U1608 ( .A(sreg[392]), .B(n2236), .Z(n1141) );
  NANDN U1609 ( .A(n2235), .B(n1141), .Z(n1142) );
  NAND U1610 ( .A(n1140), .B(n1142), .Z(n2242) );
  XOR U1611 ( .A(sreg[395]), .B(n2256), .Z(n1143) );
  NANDN U1612 ( .A(n2257), .B(n1143), .Z(n1144) );
  NAND U1613 ( .A(sreg[395]), .B(n2256), .Z(n1145) );
  AND U1614 ( .A(n1144), .B(n1145), .Z(n2263) );
  NAND U1615 ( .A(sreg[398]), .B(n2278), .Z(n1146) );
  XOR U1616 ( .A(sreg[398]), .B(n2278), .Z(n1147) );
  NANDN U1617 ( .A(n2277), .B(n1147), .Z(n1148) );
  NAND U1618 ( .A(n1146), .B(n1148), .Z(n2284) );
  NAND U1619 ( .A(n2298), .B(n2299), .Z(n1149) );
  XOR U1620 ( .A(n2298), .B(n2299), .Z(n1150) );
  NAND U1621 ( .A(n1150), .B(sreg[401]), .Z(n1151) );
  NAND U1622 ( .A(n1149), .B(n1151), .Z(n2305) );
  XOR U1623 ( .A(sreg[404]), .B(n2319), .Z(n1152) );
  NANDN U1624 ( .A(n2320), .B(n1152), .Z(n1153) );
  NAND U1625 ( .A(sreg[404]), .B(n2319), .Z(n1154) );
  AND U1626 ( .A(n1153), .B(n1154), .Z(n2326) );
  NAND U1627 ( .A(sreg[407]), .B(n2341), .Z(n1155) );
  XOR U1628 ( .A(sreg[407]), .B(n2341), .Z(n1156) );
  NANDN U1629 ( .A(n2340), .B(n1156), .Z(n1157) );
  NAND U1630 ( .A(n1155), .B(n1157), .Z(n2347) );
  NAND U1631 ( .A(n2361), .B(n2362), .Z(n1158) );
  XOR U1632 ( .A(n2361), .B(n2362), .Z(n1159) );
  NAND U1633 ( .A(n1159), .B(sreg[410]), .Z(n1160) );
  NAND U1634 ( .A(n1158), .B(n1160), .Z(n2368) );
  XOR U1635 ( .A(sreg[413]), .B(n2382), .Z(n1161) );
  NANDN U1636 ( .A(n2383), .B(n1161), .Z(n1162) );
  NAND U1637 ( .A(sreg[413]), .B(n2382), .Z(n1163) );
  AND U1638 ( .A(n1162), .B(n1163), .Z(n2389) );
  NAND U1639 ( .A(sreg[416]), .B(n2404), .Z(n1164) );
  XOR U1640 ( .A(sreg[416]), .B(n2404), .Z(n1165) );
  NANDN U1641 ( .A(n2403), .B(n1165), .Z(n1166) );
  NAND U1642 ( .A(n1164), .B(n1166), .Z(n2410) );
  XOR U1643 ( .A(sreg[419]), .B(n2424), .Z(n1167) );
  NANDN U1644 ( .A(n2425), .B(n1167), .Z(n1168) );
  NAND U1645 ( .A(sreg[419]), .B(n2424), .Z(n1169) );
  AND U1646 ( .A(n1168), .B(n1169), .Z(n2431) );
  NAND U1647 ( .A(n2445), .B(n2446), .Z(n1170) );
  XOR U1648 ( .A(n2445), .B(n2446), .Z(n1171) );
  NAND U1649 ( .A(n1171), .B(sreg[422]), .Z(n1172) );
  NAND U1650 ( .A(n1170), .B(n1172), .Z(n2452) );
  NAND U1651 ( .A(n2466), .B(n2467), .Z(n1173) );
  XOR U1652 ( .A(n2466), .B(n2467), .Z(n1174) );
  NAND U1653 ( .A(n1174), .B(sreg[425]), .Z(n1175) );
  NAND U1654 ( .A(n1173), .B(n1175), .Z(n2473) );
  NAND U1655 ( .A(n2487), .B(n2488), .Z(n1176) );
  XOR U1656 ( .A(n2487), .B(n2488), .Z(n1177) );
  NANDN U1657 ( .A(sreg[428]), .B(n1177), .Z(n1178) );
  NAND U1658 ( .A(n1176), .B(n1178), .Z(n2494) );
  NAND U1659 ( .A(n2508), .B(n2509), .Z(n1179) );
  XOR U1660 ( .A(n2508), .B(n2509), .Z(n1180) );
  NAND U1661 ( .A(n1180), .B(sreg[431]), .Z(n1181) );
  NAND U1662 ( .A(n1179), .B(n1181), .Z(n2515) );
  XOR U1663 ( .A(sreg[434]), .B(n2529), .Z(n1182) );
  NANDN U1664 ( .A(n2530), .B(n1182), .Z(n1183) );
  NAND U1665 ( .A(sreg[434]), .B(n2529), .Z(n1184) );
  AND U1666 ( .A(n1183), .B(n1184), .Z(n2536) );
  NAND U1667 ( .A(sreg[437]), .B(n2551), .Z(n1185) );
  XOR U1668 ( .A(sreg[437]), .B(n2551), .Z(n1186) );
  NANDN U1669 ( .A(n2550), .B(n1186), .Z(n1187) );
  NAND U1670 ( .A(n1185), .B(n1187), .Z(n2557) );
  XOR U1671 ( .A(sreg[440]), .B(n2571), .Z(n1188) );
  NANDN U1672 ( .A(n2572), .B(n1188), .Z(n1189) );
  NAND U1673 ( .A(sreg[440]), .B(n2571), .Z(n1190) );
  AND U1674 ( .A(n1189), .B(n1190), .Z(n2578) );
  XOR U1675 ( .A(sreg[443]), .B(n2592), .Z(n1191) );
  NANDN U1676 ( .A(n2593), .B(n1191), .Z(n1192) );
  NAND U1677 ( .A(sreg[443]), .B(n2592), .Z(n1193) );
  AND U1678 ( .A(n1192), .B(n1193), .Z(n2599) );
  NAND U1679 ( .A(sreg[446]), .B(n2614), .Z(n1194) );
  XOR U1680 ( .A(sreg[446]), .B(n2614), .Z(n1195) );
  NANDN U1681 ( .A(n2613), .B(n1195), .Z(n1196) );
  NAND U1682 ( .A(n1194), .B(n1196), .Z(n2620) );
  XOR U1683 ( .A(sreg[449]), .B(n2634), .Z(n1197) );
  NANDN U1684 ( .A(n2635), .B(n1197), .Z(n1198) );
  NAND U1685 ( .A(sreg[449]), .B(n2634), .Z(n1199) );
  AND U1686 ( .A(n1198), .B(n1199), .Z(n2641) );
  NAND U1687 ( .A(n2655), .B(n2656), .Z(n1200) );
  XOR U1688 ( .A(n2655), .B(n2656), .Z(n1201) );
  NAND U1689 ( .A(n1201), .B(sreg[452]), .Z(n1202) );
  NAND U1690 ( .A(n1200), .B(n1202), .Z(n2662) );
  XOR U1691 ( .A(sreg[455]), .B(n2676), .Z(n1203) );
  NANDN U1692 ( .A(n2677), .B(n1203), .Z(n1204) );
  NAND U1693 ( .A(sreg[455]), .B(n2676), .Z(n1205) );
  AND U1694 ( .A(n1204), .B(n1205), .Z(n2683) );
  NAND U1695 ( .A(n2697), .B(n2698), .Z(n1206) );
  XOR U1696 ( .A(n2697), .B(n2698), .Z(n1207) );
  NAND U1697 ( .A(n1207), .B(sreg[458]), .Z(n1208) );
  NAND U1698 ( .A(n1206), .B(n1208), .Z(n2704) );
  XOR U1699 ( .A(sreg[461]), .B(n2718), .Z(n1209) );
  NANDN U1700 ( .A(n2719), .B(n1209), .Z(n1210) );
  NAND U1701 ( .A(sreg[461]), .B(n2718), .Z(n1211) );
  AND U1702 ( .A(n1210), .B(n1211), .Z(n2725) );
  NAND U1703 ( .A(n2739), .B(n2740), .Z(n1212) );
  XOR U1704 ( .A(n2739), .B(n2740), .Z(n1213) );
  NAND U1705 ( .A(n1213), .B(sreg[464]), .Z(n1214) );
  NAND U1706 ( .A(n1212), .B(n1214), .Z(n2746) );
  NAND U1707 ( .A(sreg[467]), .B(n2761), .Z(n1215) );
  XOR U1708 ( .A(sreg[467]), .B(n2761), .Z(n1216) );
  NANDN U1709 ( .A(n2760), .B(n1216), .Z(n1217) );
  NAND U1710 ( .A(n1215), .B(n1217), .Z(n2767) );
  NAND U1711 ( .A(n2781), .B(n2782), .Z(n1218) );
  XOR U1712 ( .A(n2781), .B(n2782), .Z(n1219) );
  NAND U1713 ( .A(n1219), .B(sreg[470]), .Z(n1220) );
  NAND U1714 ( .A(n1218), .B(n1220), .Z(n2788) );
  NAND U1715 ( .A(n2802), .B(n2803), .Z(n1221) );
  XOR U1716 ( .A(n2802), .B(n2803), .Z(n1222) );
  NAND U1717 ( .A(n1222), .B(sreg[473]), .Z(n1223) );
  NAND U1718 ( .A(n1221), .B(n1223), .Z(n2809) );
  NAND U1719 ( .A(n2823), .B(n2824), .Z(n1224) );
  XOR U1720 ( .A(n2823), .B(n2824), .Z(n1225) );
  NANDN U1721 ( .A(sreg[476]), .B(n1225), .Z(n1226) );
  NAND U1722 ( .A(n1224), .B(n1226), .Z(n2830) );
  XOR U1723 ( .A(sreg[479]), .B(n2844), .Z(n1227) );
  NANDN U1724 ( .A(n2845), .B(n1227), .Z(n1228) );
  NAND U1725 ( .A(sreg[479]), .B(n2844), .Z(n1229) );
  AND U1726 ( .A(n1228), .B(n1229), .Z(n2851) );
  XOR U1727 ( .A(sreg[482]), .B(n2865), .Z(n1230) );
  NANDN U1728 ( .A(n2866), .B(n1230), .Z(n1231) );
  NAND U1729 ( .A(sreg[482]), .B(n2865), .Z(n1232) );
  AND U1730 ( .A(n1231), .B(n1232), .Z(n2872) );
  XOR U1731 ( .A(sreg[485]), .B(n2886), .Z(n1233) );
  NANDN U1732 ( .A(n2887), .B(n1233), .Z(n1234) );
  NAND U1733 ( .A(sreg[485]), .B(n2886), .Z(n1235) );
  AND U1734 ( .A(n1234), .B(n1235), .Z(n2893) );
  NAND U1735 ( .A(sreg[488]), .B(n2908), .Z(n1236) );
  XOR U1736 ( .A(sreg[488]), .B(n2908), .Z(n1237) );
  NANDN U1737 ( .A(n2907), .B(n1237), .Z(n1238) );
  NAND U1738 ( .A(n1236), .B(n1238), .Z(n2914) );
  NAND U1739 ( .A(n2928), .B(n2929), .Z(n1239) );
  XOR U1740 ( .A(n2928), .B(n2929), .Z(n1240) );
  NAND U1741 ( .A(n1240), .B(sreg[491]), .Z(n1241) );
  NAND U1742 ( .A(n1239), .B(n1241), .Z(n2935) );
  NAND U1743 ( .A(sreg[494]), .B(n2950), .Z(n1242) );
  XOR U1744 ( .A(sreg[494]), .B(n2950), .Z(n1243) );
  NANDN U1745 ( .A(n2949), .B(n1243), .Z(n1244) );
  NAND U1746 ( .A(n1242), .B(n1244), .Z(n2956) );
  NAND U1747 ( .A(n2970), .B(n2971), .Z(n1245) );
  XOR U1748 ( .A(n2970), .B(n2971), .Z(n1246) );
  NAND U1749 ( .A(n1246), .B(sreg[497]), .Z(n1247) );
  NAND U1750 ( .A(n1245), .B(n1247), .Z(n2977) );
  XOR U1751 ( .A(sreg[500]), .B(n2991), .Z(n1248) );
  NANDN U1752 ( .A(n2992), .B(n1248), .Z(n1249) );
  NAND U1753 ( .A(sreg[500]), .B(n2991), .Z(n1250) );
  AND U1754 ( .A(n1249), .B(n1250), .Z(n2998) );
  NAND U1755 ( .A(sreg[503]), .B(n3013), .Z(n1251) );
  XOR U1756 ( .A(sreg[503]), .B(n3013), .Z(n1252) );
  NANDN U1757 ( .A(n3012), .B(n1252), .Z(n1253) );
  NAND U1758 ( .A(n1251), .B(n1253), .Z(n3019) );
  NAND U1759 ( .A(n3033), .B(n3034), .Z(n1254) );
  XOR U1760 ( .A(n3033), .B(n3034), .Z(n1255) );
  NAND U1761 ( .A(n1255), .B(sreg[506]), .Z(n1256) );
  NAND U1762 ( .A(n1254), .B(n1256), .Z(n3040) );
  XOR U1763 ( .A(sreg[509]), .B(n3051), .Z(n1257) );
  NANDN U1764 ( .A(n3052), .B(n1257), .Z(n1258) );
  NAND U1765 ( .A(sreg[509]), .B(n3051), .Z(n1259) );
  AND U1766 ( .A(n1258), .B(n1259), .Z(n3060) );
  AND U1767 ( .A(b[0]), .B(a[0]), .Z(n1270) );
  IV U1768 ( .A(n1270), .Z(n1265) );
  XNOR U1769 ( .A(sreg[254]), .B(n1265), .Z(c[254]) );
  NAND U1770 ( .A(n1270), .B(sreg[254]), .Z(n1264) );
  AND U1771 ( .A(b[0]), .B(a[1]), .Z(n1261) );
  AND U1772 ( .A(a[0]), .B(b[1]), .Z(n1260) );
  XNOR U1773 ( .A(n1261), .B(n1260), .Z(n1263) );
  XNOR U1774 ( .A(sreg[255]), .B(n1263), .Z(n1262) );
  XNOR U1775 ( .A(n1264), .B(n1262), .Z(c[255]) );
  AND U1776 ( .A(b[0]), .B(a[2]), .Z(n1277) );
  AND U1777 ( .A(b[1]), .B(a[1]), .Z(n1269) );
  AND U1778 ( .A(n1269), .B(n1265), .Z(n1271) );
  XNOR U1779 ( .A(n1277), .B(n1271), .Z(n1266) );
  XNOR U1780 ( .A(sreg[256]), .B(n1266), .Z(n1267) );
  XNOR U1781 ( .A(n1268), .B(n1267), .Z(c[256]) );
  NAND U1782 ( .A(n1270), .B(n1269), .Z(n1273) );
  NAND U1783 ( .A(n1271), .B(n1277), .Z(n1272) );
  AND U1784 ( .A(n1273), .B(n1272), .Z(n1279) );
  AND U1785 ( .A(a[3]), .B(b[0]), .Z(n1287) );
  NAND U1786 ( .A(a[2]), .B(b[1]), .Z(n1274) );
  XNOR U1787 ( .A(n1287), .B(n1274), .Z(n1278) );
  XNOR U1788 ( .A(n1279), .B(n1278), .Z(n1284) );
  XNOR U1789 ( .A(sreg[257]), .B(n1284), .Z(n1275) );
  XNOR U1790 ( .A(n1283), .B(n1275), .Z(c[257]) );
  AND U1791 ( .A(b[1]), .B(a[3]), .Z(n1276) );
  NAND U1792 ( .A(n1277), .B(n1276), .Z(n1281) );
  NANDN U1793 ( .A(n1279), .B(n1278), .Z(n1280) );
  AND U1794 ( .A(n1281), .B(n1280), .Z(n1288) );
  AND U1795 ( .A(a[4]), .B(b[0]), .Z(n1299) );
  NAND U1796 ( .A(a[3]), .B(b[1]), .Z(n1282) );
  XOR U1797 ( .A(n1299), .B(n1282), .Z(n1289) );
  XNOR U1798 ( .A(n1288), .B(n1289), .Z(n1295) );
  XOR U1799 ( .A(n1294), .B(sreg[258]), .Z(n1285) );
  XNOR U1800 ( .A(n1295), .B(n1285), .Z(c[258]) );
  AND U1801 ( .A(b[1]), .B(a[4]), .Z(n1286) );
  NAND U1802 ( .A(n1287), .B(n1286), .Z(n1291) );
  OR U1803 ( .A(n1289), .B(n1288), .Z(n1290) );
  AND U1804 ( .A(n1291), .B(n1290), .Z(n1300) );
  AND U1805 ( .A(b[0]), .B(a[5]), .Z(n1293) );
  NAND U1806 ( .A(a[4]), .B(b[1]), .Z(n1292) );
  XOR U1807 ( .A(n1293), .B(n1292), .Z(n1301) );
  XNOR U1808 ( .A(n1300), .B(n1301), .Z(n1298) );
  XNOR U1809 ( .A(n1297), .B(sreg[259]), .Z(n1296) );
  XNOR U1810 ( .A(n1298), .B(n1296), .Z(c[259]) );
  AND U1811 ( .A(b[1]), .B(a[5]), .Z(n1304) );
  NAND U1812 ( .A(n1304), .B(n1299), .Z(n1303) );
  OR U1813 ( .A(n1301), .B(n1300), .Z(n1302) );
  AND U1814 ( .A(n1303), .B(n1302), .Z(n1307) );
  NAND U1815 ( .A(b[0]), .B(a[6]), .Z(n1305) );
  XNOR U1816 ( .A(n1304), .B(n1305), .Z(n1306) );
  XNOR U1817 ( .A(n1307), .B(n1306), .Z(n1308) );
  XNOR U1818 ( .A(sreg[260]), .B(n1308), .Z(n1310) );
  XOR U1819 ( .A(n1309), .B(n1310), .Z(c[260]) );
  AND U1820 ( .A(b[0]), .B(a[7]), .Z(n1314) );
  NAND U1821 ( .A(b[1]), .B(a[6]), .Z(n1315) );
  XNOR U1822 ( .A(n1314), .B(n1315), .Z(n1317) );
  XNOR U1823 ( .A(n1316), .B(n1317), .Z(n1319) );
  NAND U1824 ( .A(sreg[260]), .B(n1308), .Z(n1312) );
  OR U1825 ( .A(n1310), .B(n1309), .Z(n1311) );
  AND U1826 ( .A(n1312), .B(n1311), .Z(n1318) );
  XNOR U1827 ( .A(n1318), .B(sreg[261]), .Z(n1313) );
  XNOR U1828 ( .A(n1319), .B(n1313), .Z(c[261]) );
  AND U1829 ( .A(b[0]), .B(a[8]), .Z(n1321) );
  NAND U1830 ( .A(b[1]), .B(a[7]), .Z(n1322) );
  XOR U1831 ( .A(n1321), .B(n1322), .Z(n1324) );
  XOR U1832 ( .A(n1323), .B(n1324), .Z(n1326) );
  XOR U1833 ( .A(sreg[262]), .B(n1325), .Z(n1320) );
  XNOR U1834 ( .A(n1326), .B(n1320), .Z(c[262]) );
  AND U1835 ( .A(b[0]), .B(a[9]), .Z(n1328) );
  NAND U1836 ( .A(b[1]), .B(a[8]), .Z(n1329) );
  XOR U1837 ( .A(n1328), .B(n1329), .Z(n1331) );
  XOR U1838 ( .A(n1330), .B(n1331), .Z(n1333) );
  XNOR U1839 ( .A(sreg[263]), .B(n1332), .Z(n1327) );
  XNOR U1840 ( .A(n1333), .B(n1327), .Z(c[263]) );
  AND U1841 ( .A(b[0]), .B(a[10]), .Z(n1335) );
  NAND U1842 ( .A(b[1]), .B(a[9]), .Z(n1336) );
  XNOR U1843 ( .A(n1335), .B(n1336), .Z(n1338) );
  XNOR U1844 ( .A(n1337), .B(n1338), .Z(n1340) );
  XOR U1845 ( .A(n1339), .B(sreg[264]), .Z(n1334) );
  XNOR U1846 ( .A(n1340), .B(n1334), .Z(c[264]) );
  AND U1847 ( .A(b[0]), .B(a[11]), .Z(n1342) );
  NAND U1848 ( .A(b[1]), .B(a[10]), .Z(n1343) );
  XOR U1849 ( .A(n1342), .B(n1343), .Z(n1345) );
  XOR U1850 ( .A(n1344), .B(n1345), .Z(n1347) );
  XOR U1851 ( .A(sreg[265]), .B(n1346), .Z(n1341) );
  XNOR U1852 ( .A(n1347), .B(n1341), .Z(c[265]) );
  AND U1853 ( .A(b[0]), .B(a[12]), .Z(n1349) );
  NAND U1854 ( .A(b[1]), .B(a[11]), .Z(n1350) );
  XOR U1855 ( .A(n1349), .B(n1350), .Z(n1352) );
  XOR U1856 ( .A(n1351), .B(n1352), .Z(n1354) );
  XNOR U1857 ( .A(sreg[266]), .B(n1353), .Z(n1348) );
  XNOR U1858 ( .A(n1354), .B(n1348), .Z(c[266]) );
  AND U1859 ( .A(b[0]), .B(a[13]), .Z(n1356) );
  NAND U1860 ( .A(b[1]), .B(a[12]), .Z(n1357) );
  XNOR U1861 ( .A(n1356), .B(n1357), .Z(n1359) );
  XNOR U1862 ( .A(n1358), .B(n1359), .Z(n1361) );
  XOR U1863 ( .A(n1360), .B(sreg[267]), .Z(n1355) );
  XNOR U1864 ( .A(n1361), .B(n1355), .Z(c[267]) );
  AND U1865 ( .A(b[0]), .B(a[14]), .Z(n1363) );
  NAND U1866 ( .A(b[1]), .B(a[13]), .Z(n1364) );
  XOR U1867 ( .A(n1363), .B(n1364), .Z(n1366) );
  XOR U1868 ( .A(n1365), .B(n1366), .Z(n1368) );
  XOR U1869 ( .A(sreg[268]), .B(n1367), .Z(n1362) );
  XNOR U1870 ( .A(n1368), .B(n1362), .Z(c[268]) );
  AND U1871 ( .A(b[0]), .B(a[15]), .Z(n1370) );
  NAND U1872 ( .A(b[1]), .B(a[14]), .Z(n1371) );
  XNOR U1873 ( .A(n1370), .B(n1371), .Z(n1373) );
  XNOR U1874 ( .A(n1372), .B(n1373), .Z(n1375) );
  XOR U1875 ( .A(n1374), .B(sreg[269]), .Z(n1369) );
  XNOR U1876 ( .A(n1375), .B(n1369), .Z(c[269]) );
  AND U1877 ( .A(b[0]), .B(a[16]), .Z(n1377) );
  NAND U1878 ( .A(b[1]), .B(a[15]), .Z(n1378) );
  XNOR U1879 ( .A(n1377), .B(n1378), .Z(n1380) );
  XNOR U1880 ( .A(n1379), .B(n1380), .Z(n1382) );
  XNOR U1881 ( .A(n1381), .B(sreg[270]), .Z(n1376) );
  XNOR U1882 ( .A(n1382), .B(n1376), .Z(c[270]) );
  AND U1883 ( .A(b[0]), .B(a[17]), .Z(n1384) );
  NAND U1884 ( .A(b[1]), .B(a[16]), .Z(n1385) );
  XNOR U1885 ( .A(n1384), .B(n1385), .Z(n1387) );
  XNOR U1886 ( .A(n1386), .B(n1387), .Z(n1389) );
  XNOR U1887 ( .A(n1388), .B(sreg[271]), .Z(n1383) );
  XNOR U1888 ( .A(n1389), .B(n1383), .Z(c[271]) );
  AND U1889 ( .A(b[0]), .B(a[18]), .Z(n1391) );
  NAND U1890 ( .A(b[1]), .B(a[17]), .Z(n1392) );
  XOR U1891 ( .A(n1391), .B(n1392), .Z(n1394) );
  XOR U1892 ( .A(n1393), .B(n1394), .Z(n1396) );
  XOR U1893 ( .A(sreg[272]), .B(n1395), .Z(n1390) );
  XNOR U1894 ( .A(n1396), .B(n1390), .Z(c[272]) );
  AND U1895 ( .A(b[0]), .B(a[19]), .Z(n1398) );
  NAND U1896 ( .A(b[1]), .B(a[18]), .Z(n1399) );
  XOR U1897 ( .A(n1398), .B(n1399), .Z(n1401) );
  XOR U1898 ( .A(n1400), .B(n1401), .Z(n1403) );
  XNOR U1899 ( .A(sreg[273]), .B(n1402), .Z(n1397) );
  XNOR U1900 ( .A(n1403), .B(n1397), .Z(c[273]) );
  AND U1901 ( .A(b[0]), .B(a[20]), .Z(n1405) );
  NAND U1902 ( .A(b[1]), .B(a[19]), .Z(n1406) );
  XNOR U1903 ( .A(n1405), .B(n1406), .Z(n1408) );
  XNOR U1904 ( .A(n1407), .B(n1408), .Z(n1410) );
  XOR U1905 ( .A(n1409), .B(sreg[274]), .Z(n1404) );
  XNOR U1906 ( .A(n1410), .B(n1404), .Z(c[274]) );
  AND U1907 ( .A(b[0]), .B(a[21]), .Z(n1412) );
  NAND U1908 ( .A(b[1]), .B(a[20]), .Z(n1413) );
  XOR U1909 ( .A(n1412), .B(n1413), .Z(n1415) );
  XOR U1910 ( .A(n1414), .B(n1415), .Z(n1417) );
  XOR U1911 ( .A(sreg[275]), .B(n1416), .Z(n1411) );
  XNOR U1912 ( .A(n1417), .B(n1411), .Z(c[275]) );
  AND U1913 ( .A(b[0]), .B(a[22]), .Z(n1419) );
  NAND U1914 ( .A(b[1]), .B(a[21]), .Z(n1420) );
  XNOR U1915 ( .A(n1419), .B(n1420), .Z(n1422) );
  XNOR U1916 ( .A(n1421), .B(n1422), .Z(n1424) );
  XOR U1917 ( .A(n1423), .B(sreg[276]), .Z(n1418) );
  XNOR U1918 ( .A(n1424), .B(n1418), .Z(c[276]) );
  AND U1919 ( .A(b[0]), .B(a[23]), .Z(n1426) );
  NAND U1920 ( .A(b[1]), .B(a[22]), .Z(n1427) );
  XOR U1921 ( .A(n1426), .B(n1427), .Z(n1429) );
  XOR U1922 ( .A(n1428), .B(n1429), .Z(n1431) );
  XOR U1923 ( .A(sreg[277]), .B(n1430), .Z(n1425) );
  XNOR U1924 ( .A(n1431), .B(n1425), .Z(c[277]) );
  AND U1925 ( .A(b[0]), .B(a[24]), .Z(n1433) );
  NAND U1926 ( .A(b[1]), .B(a[23]), .Z(n1434) );
  XNOR U1927 ( .A(n1433), .B(n1434), .Z(n1436) );
  XNOR U1928 ( .A(n1435), .B(n1436), .Z(n1438) );
  XOR U1929 ( .A(n1437), .B(sreg[278]), .Z(n1432) );
  XNOR U1930 ( .A(n1438), .B(n1432), .Z(c[278]) );
  AND U1931 ( .A(b[0]), .B(a[25]), .Z(n1440) );
  NAND U1932 ( .A(b[1]), .B(a[24]), .Z(n1441) );
  XOR U1933 ( .A(n1440), .B(n1441), .Z(n1443) );
  XOR U1934 ( .A(n1442), .B(n1443), .Z(n1445) );
  XOR U1935 ( .A(sreg[279]), .B(n1444), .Z(n1439) );
  XNOR U1936 ( .A(n1445), .B(n1439), .Z(c[279]) );
  AND U1937 ( .A(b[0]), .B(a[26]), .Z(n1447) );
  NAND U1938 ( .A(b[1]), .B(a[25]), .Z(n1448) );
  XOR U1939 ( .A(n1447), .B(n1448), .Z(n1450) );
  XOR U1940 ( .A(n1449), .B(n1450), .Z(n1452) );
  XNOR U1941 ( .A(sreg[280]), .B(n1451), .Z(n1446) );
  XNOR U1942 ( .A(n1452), .B(n1446), .Z(c[280]) );
  AND U1943 ( .A(b[0]), .B(a[27]), .Z(n1454) );
  NAND U1944 ( .A(b[1]), .B(a[26]), .Z(n1455) );
  XOR U1945 ( .A(n1454), .B(n1455), .Z(n1457) );
  XOR U1946 ( .A(n1456), .B(n1457), .Z(n1459) );
  XNOR U1947 ( .A(sreg[281]), .B(n1458), .Z(n1453) );
  XNOR U1948 ( .A(n1459), .B(n1453), .Z(c[281]) );
  AND U1949 ( .A(b[0]), .B(a[28]), .Z(n1461) );
  NAND U1950 ( .A(b[1]), .B(a[27]), .Z(n1462) );
  XOR U1951 ( .A(n1461), .B(n1462), .Z(n1464) );
  XOR U1952 ( .A(n1463), .B(n1464), .Z(n1465) );
  XNOR U1953 ( .A(sreg[282]), .B(n1466), .Z(n1460) );
  XNOR U1954 ( .A(n1465), .B(n1460), .Z(c[282]) );
  AND U1955 ( .A(b[0]), .B(a[29]), .Z(n1468) );
  NAND U1956 ( .A(b[1]), .B(a[28]), .Z(n1469) );
  XNOR U1957 ( .A(n1468), .B(n1469), .Z(n1471) );
  XNOR U1958 ( .A(n1470), .B(n1471), .Z(n1473) );
  XOR U1959 ( .A(n1472), .B(sreg[283]), .Z(n1467) );
  XNOR U1960 ( .A(n1473), .B(n1467), .Z(c[283]) );
  AND U1961 ( .A(b[0]), .B(a[30]), .Z(n1475) );
  NAND U1962 ( .A(b[1]), .B(a[29]), .Z(n1476) );
  XOR U1963 ( .A(n1475), .B(n1476), .Z(n1478) );
  XOR U1964 ( .A(n1477), .B(n1478), .Z(n1480) );
  XOR U1965 ( .A(sreg[284]), .B(n1479), .Z(n1474) );
  XNOR U1966 ( .A(n1480), .B(n1474), .Z(c[284]) );
  AND U1967 ( .A(b[0]), .B(a[31]), .Z(n1482) );
  NAND U1968 ( .A(b[1]), .B(a[30]), .Z(n1483) );
  XNOR U1969 ( .A(n1482), .B(n1483), .Z(n1485) );
  XNOR U1970 ( .A(n1484), .B(n1485), .Z(n1487) );
  XOR U1971 ( .A(n1486), .B(sreg[285]), .Z(n1481) );
  XNOR U1972 ( .A(n1487), .B(n1481), .Z(c[285]) );
  AND U1973 ( .A(b[0]), .B(a[32]), .Z(n1489) );
  NAND U1974 ( .A(b[1]), .B(a[31]), .Z(n1490) );
  XOR U1975 ( .A(n1489), .B(n1490), .Z(n1492) );
  XOR U1976 ( .A(n1491), .B(n1492), .Z(n1494) );
  XOR U1977 ( .A(sreg[286]), .B(n1493), .Z(n1488) );
  XNOR U1978 ( .A(n1494), .B(n1488), .Z(c[286]) );
  AND U1979 ( .A(b[0]), .B(a[33]), .Z(n1496) );
  NAND U1980 ( .A(b[1]), .B(a[32]), .Z(n1497) );
  XNOR U1981 ( .A(n1496), .B(n1497), .Z(n1499) );
  XNOR U1982 ( .A(n1498), .B(n1499), .Z(n1501) );
  XOR U1983 ( .A(n1500), .B(sreg[287]), .Z(n1495) );
  XNOR U1984 ( .A(n1501), .B(n1495), .Z(c[287]) );
  AND U1985 ( .A(b[0]), .B(a[34]), .Z(n1503) );
  NAND U1986 ( .A(b[1]), .B(a[33]), .Z(n1504) );
  XOR U1987 ( .A(n1503), .B(n1504), .Z(n1506) );
  XOR U1988 ( .A(n1505), .B(n1506), .Z(n1508) );
  XOR U1989 ( .A(sreg[288]), .B(n1507), .Z(n1502) );
  XNOR U1990 ( .A(n1508), .B(n1502), .Z(c[288]) );
  AND U1991 ( .A(b[0]), .B(a[35]), .Z(n1510) );
  NAND U1992 ( .A(b[1]), .B(a[34]), .Z(n1511) );
  XNOR U1993 ( .A(n1510), .B(n1511), .Z(n1513) );
  XNOR U1994 ( .A(n1512), .B(n1513), .Z(n1515) );
  XOR U1995 ( .A(n1514), .B(sreg[289]), .Z(n1509) );
  XNOR U1996 ( .A(n1515), .B(n1509), .Z(c[289]) );
  AND U1997 ( .A(b[0]), .B(a[36]), .Z(n1517) );
  NAND U1998 ( .A(b[1]), .B(a[35]), .Z(n1518) );
  XNOR U1999 ( .A(n1517), .B(n1518), .Z(n1520) );
  XNOR U2000 ( .A(n1519), .B(n1520), .Z(n1522) );
  XNOR U2001 ( .A(n1521), .B(sreg[290]), .Z(n1516) );
  XNOR U2002 ( .A(n1522), .B(n1516), .Z(c[290]) );
  AND U2003 ( .A(b[0]), .B(a[37]), .Z(n1524) );
  NAND U2004 ( .A(b[1]), .B(a[36]), .Z(n1525) );
  XOR U2005 ( .A(n1524), .B(n1525), .Z(n1527) );
  XOR U2006 ( .A(n1526), .B(n1527), .Z(n1529) );
  XOR U2007 ( .A(sreg[291]), .B(n1528), .Z(n1523) );
  XNOR U2008 ( .A(n1529), .B(n1523), .Z(c[291]) );
  AND U2009 ( .A(b[0]), .B(a[38]), .Z(n1531) );
  NAND U2010 ( .A(b[1]), .B(a[37]), .Z(n1532) );
  XOR U2011 ( .A(n1531), .B(n1532), .Z(n1534) );
  XOR U2012 ( .A(n1533), .B(n1534), .Z(n1536) );
  XNOR U2013 ( .A(sreg[292]), .B(n1535), .Z(n1530) );
  XNOR U2014 ( .A(n1536), .B(n1530), .Z(c[292]) );
  AND U2015 ( .A(b[0]), .B(a[39]), .Z(n1538) );
  NAND U2016 ( .A(b[1]), .B(a[38]), .Z(n1539) );
  XOR U2017 ( .A(n1538), .B(n1539), .Z(n1541) );
  XOR U2018 ( .A(n1540), .B(n1541), .Z(n1543) );
  XNOR U2019 ( .A(sreg[293]), .B(n1542), .Z(n1537) );
  XNOR U2020 ( .A(n1543), .B(n1537), .Z(c[293]) );
  AND U2021 ( .A(b[0]), .B(a[40]), .Z(n1545) );
  NAND U2022 ( .A(b[1]), .B(a[39]), .Z(n1546) );
  XOR U2023 ( .A(n1545), .B(n1546), .Z(n1548) );
  XOR U2024 ( .A(n1547), .B(n1548), .Z(n1550) );
  XNOR U2025 ( .A(sreg[294]), .B(n1549), .Z(n1544) );
  XNOR U2026 ( .A(n1550), .B(n1544), .Z(c[294]) );
  AND U2027 ( .A(b[0]), .B(a[41]), .Z(n1552) );
  NAND U2028 ( .A(b[1]), .B(a[40]), .Z(n1553) );
  XNOR U2029 ( .A(n1552), .B(n1553), .Z(n1555) );
  XNOR U2030 ( .A(n1554), .B(n1555), .Z(n1557) );
  XOR U2031 ( .A(n1556), .B(sreg[295]), .Z(n1551) );
  XNOR U2032 ( .A(n1557), .B(n1551), .Z(c[295]) );
  AND U2033 ( .A(b[0]), .B(a[42]), .Z(n1559) );
  NAND U2034 ( .A(b[1]), .B(a[41]), .Z(n1560) );
  XOR U2035 ( .A(n1559), .B(n1560), .Z(n1562) );
  XOR U2036 ( .A(n1561), .B(n1562), .Z(n1564) );
  XOR U2037 ( .A(sreg[296]), .B(n1563), .Z(n1558) );
  XNOR U2038 ( .A(n1564), .B(n1558), .Z(c[296]) );
  AND U2039 ( .A(b[0]), .B(a[43]), .Z(n1566) );
  NAND U2040 ( .A(b[1]), .B(a[42]), .Z(n1567) );
  XOR U2041 ( .A(n1566), .B(n1567), .Z(n1569) );
  XOR U2042 ( .A(n1568), .B(n1569), .Z(n1571) );
  XNOR U2043 ( .A(sreg[297]), .B(n1570), .Z(n1565) );
  XNOR U2044 ( .A(n1571), .B(n1565), .Z(c[297]) );
  AND U2045 ( .A(b[0]), .B(a[44]), .Z(n1573) );
  NAND U2046 ( .A(b[1]), .B(a[43]), .Z(n1574) );
  XOR U2047 ( .A(n1573), .B(n1574), .Z(n1576) );
  XOR U2048 ( .A(n1575), .B(n1576), .Z(n1578) );
  XNOR U2049 ( .A(sreg[298]), .B(n1577), .Z(n1572) );
  XNOR U2050 ( .A(n1578), .B(n1572), .Z(c[298]) );
  AND U2051 ( .A(b[0]), .B(a[45]), .Z(n1580) );
  NAND U2052 ( .A(b[1]), .B(a[44]), .Z(n1581) );
  XNOR U2053 ( .A(n1580), .B(n1581), .Z(n1583) );
  XNOR U2054 ( .A(n1582), .B(n1583), .Z(n1585) );
  XOR U2055 ( .A(n1584), .B(sreg[299]), .Z(n1579) );
  XNOR U2056 ( .A(n1585), .B(n1579), .Z(c[299]) );
  AND U2057 ( .A(b[0]), .B(a[46]), .Z(n1587) );
  NAND U2058 ( .A(b[1]), .B(a[45]), .Z(n1588) );
  XOR U2059 ( .A(n1587), .B(n1588), .Z(n1590) );
  XOR U2060 ( .A(n1589), .B(n1590), .Z(n1592) );
  XOR U2061 ( .A(sreg[300]), .B(n1591), .Z(n1586) );
  XNOR U2062 ( .A(n1592), .B(n1586), .Z(c[300]) );
  AND U2063 ( .A(b[0]), .B(a[47]), .Z(n1594) );
  NAND U2064 ( .A(b[1]), .B(a[46]), .Z(n1595) );
  XNOR U2065 ( .A(n1594), .B(n1595), .Z(n1597) );
  XNOR U2066 ( .A(n1596), .B(n1597), .Z(n1599) );
  XOR U2067 ( .A(n1598), .B(sreg[301]), .Z(n1593) );
  XNOR U2068 ( .A(n1599), .B(n1593), .Z(c[301]) );
  AND U2069 ( .A(b[0]), .B(a[48]), .Z(n1601) );
  NAND U2070 ( .A(b[1]), .B(a[47]), .Z(n1602) );
  XOR U2071 ( .A(n1601), .B(n1602), .Z(n1604) );
  XOR U2072 ( .A(n1603), .B(n1604), .Z(n1606) );
  XOR U2073 ( .A(sreg[302]), .B(n1605), .Z(n1600) );
  XNOR U2074 ( .A(n1606), .B(n1600), .Z(c[302]) );
  AND U2075 ( .A(b[0]), .B(a[49]), .Z(n1608) );
  NAND U2076 ( .A(b[1]), .B(a[48]), .Z(n1609) );
  XOR U2077 ( .A(n1608), .B(n1609), .Z(n1611) );
  XOR U2078 ( .A(n1610), .B(n1611), .Z(n1613) );
  XNOR U2079 ( .A(sreg[303]), .B(n1612), .Z(n1607) );
  XNOR U2080 ( .A(n1613), .B(n1607), .Z(c[303]) );
  AND U2081 ( .A(b[0]), .B(a[50]), .Z(n1615) );
  NAND U2082 ( .A(b[1]), .B(a[49]), .Z(n1616) );
  XOR U2083 ( .A(n1615), .B(n1616), .Z(n1618) );
  XOR U2084 ( .A(n1617), .B(n1618), .Z(n1620) );
  XNOR U2085 ( .A(sreg[304]), .B(n1619), .Z(n1614) );
  XNOR U2086 ( .A(n1620), .B(n1614), .Z(c[304]) );
  AND U2087 ( .A(b[0]), .B(a[51]), .Z(n1622) );
  NAND U2088 ( .A(b[1]), .B(a[50]), .Z(n1623) );
  XOR U2089 ( .A(n1622), .B(n1623), .Z(n1625) );
  XOR U2090 ( .A(n1624), .B(n1625), .Z(n1627) );
  XNOR U2091 ( .A(sreg[305]), .B(n1626), .Z(n1621) );
  XNOR U2092 ( .A(n1627), .B(n1621), .Z(c[305]) );
  AND U2093 ( .A(b[0]), .B(a[52]), .Z(n1629) );
  NAND U2094 ( .A(b[1]), .B(a[51]), .Z(n1630) );
  XNOR U2095 ( .A(n1629), .B(n1630), .Z(n1632) );
  XNOR U2096 ( .A(n1631), .B(n1632), .Z(n1634) );
  XOR U2097 ( .A(n1633), .B(sreg[306]), .Z(n1628) );
  XNOR U2098 ( .A(n1634), .B(n1628), .Z(c[306]) );
  AND U2099 ( .A(b[0]), .B(a[53]), .Z(n1636) );
  NAND U2100 ( .A(b[1]), .B(a[52]), .Z(n1637) );
  XOR U2101 ( .A(n1636), .B(n1637), .Z(n1639) );
  XOR U2102 ( .A(n1638), .B(n1639), .Z(n1641) );
  XOR U2103 ( .A(sreg[307]), .B(n1640), .Z(n1635) );
  XNOR U2104 ( .A(n1641), .B(n1635), .Z(c[307]) );
  AND U2105 ( .A(b[0]), .B(a[54]), .Z(n1643) );
  NAND U2106 ( .A(b[1]), .B(a[53]), .Z(n1644) );
  XNOR U2107 ( .A(n1643), .B(n1644), .Z(n1646) );
  XNOR U2108 ( .A(n1645), .B(n1646), .Z(n1648) );
  XOR U2109 ( .A(n1647), .B(sreg[308]), .Z(n1642) );
  XNOR U2110 ( .A(n1648), .B(n1642), .Z(c[308]) );
  AND U2111 ( .A(b[0]), .B(a[55]), .Z(n1650) );
  NAND U2112 ( .A(b[1]), .B(a[54]), .Z(n1651) );
  XOR U2113 ( .A(n1650), .B(n1651), .Z(n1653) );
  XOR U2114 ( .A(n1652), .B(n1653), .Z(n1655) );
  XOR U2115 ( .A(sreg[309]), .B(n1654), .Z(n1649) );
  XNOR U2116 ( .A(n1655), .B(n1649), .Z(c[309]) );
  AND U2117 ( .A(b[0]), .B(a[56]), .Z(n1657) );
  NAND U2118 ( .A(b[1]), .B(a[55]), .Z(n1658) );
  XNOR U2119 ( .A(n1657), .B(n1658), .Z(n1660) );
  XNOR U2120 ( .A(n1659), .B(n1660), .Z(n1662) );
  XOR U2121 ( .A(n1661), .B(sreg[310]), .Z(n1656) );
  XNOR U2122 ( .A(n1662), .B(n1656), .Z(c[310]) );
  AND U2123 ( .A(b[0]), .B(a[57]), .Z(n1664) );
  NAND U2124 ( .A(b[1]), .B(a[56]), .Z(n1665) );
  XNOR U2125 ( .A(n1664), .B(n1665), .Z(n1667) );
  XNOR U2126 ( .A(n1666), .B(n1667), .Z(n1669) );
  XNOR U2127 ( .A(n1668), .B(sreg[311]), .Z(n1663) );
  XNOR U2128 ( .A(n1669), .B(n1663), .Z(c[311]) );
  AND U2129 ( .A(b[0]), .B(a[58]), .Z(n1671) );
  NAND U2130 ( .A(b[1]), .B(a[57]), .Z(n1672) );
  XNOR U2131 ( .A(n1671), .B(n1672), .Z(n1674) );
  XNOR U2132 ( .A(n1673), .B(n1674), .Z(n1676) );
  XNOR U2133 ( .A(n1675), .B(sreg[312]), .Z(n1670) );
  XNOR U2134 ( .A(n1676), .B(n1670), .Z(c[312]) );
  AND U2135 ( .A(b[0]), .B(a[59]), .Z(n1678) );
  NAND U2136 ( .A(b[1]), .B(a[58]), .Z(n1679) );
  XOR U2137 ( .A(n1678), .B(n1679), .Z(n1681) );
  XOR U2138 ( .A(n1680), .B(n1681), .Z(n1683) );
  XOR U2139 ( .A(sreg[313]), .B(n1682), .Z(n1677) );
  XNOR U2140 ( .A(n1683), .B(n1677), .Z(c[313]) );
  AND U2141 ( .A(b[0]), .B(a[60]), .Z(n1685) );
  NAND U2142 ( .A(b[1]), .B(a[59]), .Z(n1686) );
  XOR U2143 ( .A(n1685), .B(n1686), .Z(n1688) );
  XOR U2144 ( .A(n1687), .B(n1688), .Z(n1690) );
  XNOR U2145 ( .A(sreg[314]), .B(n1689), .Z(n1684) );
  XNOR U2146 ( .A(n1690), .B(n1684), .Z(c[314]) );
  AND U2147 ( .A(b[0]), .B(a[61]), .Z(n1692) );
  NAND U2148 ( .A(b[1]), .B(a[60]), .Z(n1693) );
  XOR U2149 ( .A(n1692), .B(n1693), .Z(n1695) );
  XOR U2150 ( .A(n1694), .B(n1695), .Z(n1697) );
  XNOR U2151 ( .A(sreg[315]), .B(n1696), .Z(n1691) );
  XNOR U2152 ( .A(n1697), .B(n1691), .Z(c[315]) );
  AND U2153 ( .A(b[0]), .B(a[62]), .Z(n1699) );
  NAND U2154 ( .A(b[1]), .B(a[61]), .Z(n1700) );
  XOR U2155 ( .A(n1699), .B(n1700), .Z(n1702) );
  XOR U2156 ( .A(n1701), .B(n1702), .Z(n1704) );
  XNOR U2157 ( .A(sreg[316]), .B(n1703), .Z(n1698) );
  XNOR U2158 ( .A(n1704), .B(n1698), .Z(c[316]) );
  AND U2159 ( .A(b[0]), .B(a[63]), .Z(n1706) );
  NAND U2160 ( .A(b[1]), .B(a[62]), .Z(n1707) );
  XNOR U2161 ( .A(n1706), .B(n1707), .Z(n1709) );
  XNOR U2162 ( .A(n1708), .B(n1709), .Z(n1711) );
  XOR U2163 ( .A(n1710), .B(sreg[317]), .Z(n1705) );
  XNOR U2164 ( .A(n1711), .B(n1705), .Z(c[317]) );
  AND U2165 ( .A(b[0]), .B(a[64]), .Z(n1713) );
  NAND U2166 ( .A(b[1]), .B(a[63]), .Z(n1714) );
  XOR U2167 ( .A(n1713), .B(n1714), .Z(n1716) );
  XOR U2168 ( .A(n1715), .B(n1716), .Z(n1718) );
  XOR U2169 ( .A(sreg[318]), .B(n1717), .Z(n1712) );
  XNOR U2170 ( .A(n1718), .B(n1712), .Z(c[318]) );
  AND U2171 ( .A(b[0]), .B(a[65]), .Z(n1720) );
  NAND U2172 ( .A(b[1]), .B(a[64]), .Z(n1721) );
  XNOR U2173 ( .A(n1720), .B(n1721), .Z(n1723) );
  XNOR U2174 ( .A(n1722), .B(n1723), .Z(n1725) );
  XOR U2175 ( .A(n1724), .B(sreg[319]), .Z(n1719) );
  XNOR U2176 ( .A(n1725), .B(n1719), .Z(c[319]) );
  AND U2177 ( .A(b[0]), .B(a[66]), .Z(n1727) );
  NAND U2178 ( .A(b[1]), .B(a[65]), .Z(n1728) );
  XOR U2179 ( .A(n1727), .B(n1728), .Z(n1730) );
  XOR U2180 ( .A(n1729), .B(n1730), .Z(n1732) );
  XOR U2181 ( .A(sreg[320]), .B(n1731), .Z(n1726) );
  XNOR U2182 ( .A(n1732), .B(n1726), .Z(c[320]) );
  AND U2183 ( .A(b[0]), .B(a[67]), .Z(n1734) );
  NAND U2184 ( .A(b[1]), .B(a[66]), .Z(n1735) );
  XNOR U2185 ( .A(n1734), .B(n1735), .Z(n1737) );
  XNOR U2186 ( .A(n1736), .B(n1737), .Z(n1739) );
  XOR U2187 ( .A(n1738), .B(sreg[321]), .Z(n1733) );
  XNOR U2188 ( .A(n1739), .B(n1733), .Z(c[321]) );
  AND U2189 ( .A(b[0]), .B(a[68]), .Z(n1741) );
  NAND U2190 ( .A(b[1]), .B(a[67]), .Z(n1742) );
  XOR U2191 ( .A(n1741), .B(n1742), .Z(n1744) );
  XOR U2192 ( .A(n1743), .B(n1744), .Z(n1746) );
  XOR U2193 ( .A(sreg[322]), .B(n1745), .Z(n1740) );
  XNOR U2194 ( .A(n1746), .B(n1740), .Z(c[322]) );
  AND U2195 ( .A(b[0]), .B(a[69]), .Z(n1748) );
  NAND U2196 ( .A(b[1]), .B(a[68]), .Z(n1749) );
  XOR U2197 ( .A(n1748), .B(n1749), .Z(n1751) );
  XOR U2198 ( .A(n1750), .B(n1751), .Z(n1753) );
  XNOR U2199 ( .A(sreg[323]), .B(n1752), .Z(n1747) );
  XNOR U2200 ( .A(n1753), .B(n1747), .Z(c[323]) );
  AND U2201 ( .A(b[0]), .B(a[70]), .Z(n1755) );
  NAND U2202 ( .A(b[1]), .B(a[69]), .Z(n1756) );
  XOR U2203 ( .A(n1755), .B(n1756), .Z(n1758) );
  XOR U2204 ( .A(n1757), .B(n1758), .Z(n1760) );
  XNOR U2205 ( .A(sreg[324]), .B(n1759), .Z(n1754) );
  XNOR U2206 ( .A(n1760), .B(n1754), .Z(c[324]) );
  AND U2207 ( .A(b[0]), .B(a[71]), .Z(n1762) );
  NAND U2208 ( .A(b[1]), .B(a[70]), .Z(n1763) );
  XNOR U2209 ( .A(n1762), .B(n1763), .Z(n1765) );
  XNOR U2210 ( .A(n1764), .B(n1765), .Z(n1767) );
  XOR U2211 ( .A(n1766), .B(sreg[325]), .Z(n1761) );
  XNOR U2212 ( .A(n1767), .B(n1761), .Z(c[325]) );
  AND U2213 ( .A(b[0]), .B(a[72]), .Z(n1769) );
  NAND U2214 ( .A(b[1]), .B(a[71]), .Z(n1770) );
  XOR U2215 ( .A(n1769), .B(n1770), .Z(n1772) );
  XOR U2216 ( .A(n1771), .B(n1772), .Z(n1774) );
  XOR U2217 ( .A(sreg[326]), .B(n1773), .Z(n1768) );
  XNOR U2218 ( .A(n1774), .B(n1768), .Z(c[326]) );
  AND U2219 ( .A(b[0]), .B(a[73]), .Z(n1776) );
  NAND U2220 ( .A(b[1]), .B(a[72]), .Z(n1777) );
  XOR U2221 ( .A(n1776), .B(n1777), .Z(n1779) );
  XOR U2222 ( .A(n1778), .B(n1779), .Z(n1781) );
  XNOR U2223 ( .A(sreg[327]), .B(n1780), .Z(n1775) );
  XNOR U2224 ( .A(n1781), .B(n1775), .Z(c[327]) );
  AND U2225 ( .A(b[0]), .B(a[74]), .Z(n1783) );
  NAND U2226 ( .A(b[1]), .B(a[73]), .Z(n1784) );
  XOR U2227 ( .A(n1783), .B(n1784), .Z(n1786) );
  XOR U2228 ( .A(n1785), .B(n1786), .Z(n1788) );
  XNOR U2229 ( .A(sreg[328]), .B(n1787), .Z(n1782) );
  XNOR U2230 ( .A(n1788), .B(n1782), .Z(c[328]) );
  AND U2231 ( .A(b[0]), .B(a[75]), .Z(n1790) );
  NAND U2232 ( .A(b[1]), .B(a[74]), .Z(n1791) );
  XOR U2233 ( .A(n1790), .B(n1791), .Z(n1793) );
  XOR U2234 ( .A(n1792), .B(n1793), .Z(n1795) );
  XNOR U2235 ( .A(sreg[329]), .B(n1794), .Z(n1789) );
  XNOR U2236 ( .A(n1795), .B(n1789), .Z(c[329]) );
  AND U2237 ( .A(b[0]), .B(a[76]), .Z(n1797) );
  NAND U2238 ( .A(b[1]), .B(a[75]), .Z(n1798) );
  XOR U2239 ( .A(n1797), .B(n1798), .Z(n1800) );
  XOR U2240 ( .A(n1799), .B(n1800), .Z(n1802) );
  XNOR U2241 ( .A(sreg[330]), .B(n1801), .Z(n1796) );
  XNOR U2242 ( .A(n1802), .B(n1796), .Z(c[330]) );
  AND U2243 ( .A(b[0]), .B(a[77]), .Z(n1804) );
  NAND U2244 ( .A(b[1]), .B(a[76]), .Z(n1805) );
  XOR U2245 ( .A(n1804), .B(n1805), .Z(n1807) );
  XOR U2246 ( .A(n1806), .B(n1807), .Z(n1809) );
  XNOR U2247 ( .A(sreg[331]), .B(n1808), .Z(n1803) );
  XNOR U2248 ( .A(n1809), .B(n1803), .Z(c[331]) );
  AND U2249 ( .A(b[0]), .B(a[78]), .Z(n1811) );
  NAND U2250 ( .A(b[1]), .B(a[77]), .Z(n1812) );
  XOR U2251 ( .A(n1811), .B(n1812), .Z(n1814) );
  XOR U2252 ( .A(n1813), .B(n1814), .Z(n1816) );
  XNOR U2253 ( .A(sreg[332]), .B(n1815), .Z(n1810) );
  XNOR U2254 ( .A(n1816), .B(n1810), .Z(c[332]) );
  AND U2255 ( .A(b[0]), .B(a[79]), .Z(n1818) );
  NAND U2256 ( .A(b[1]), .B(a[78]), .Z(n1819) );
  XNOR U2257 ( .A(n1818), .B(n1819), .Z(n1821) );
  XNOR U2258 ( .A(n1820), .B(n1821), .Z(n1823) );
  XOR U2259 ( .A(n1822), .B(sreg[333]), .Z(n1817) );
  XNOR U2260 ( .A(n1823), .B(n1817), .Z(c[333]) );
  AND U2261 ( .A(b[0]), .B(a[80]), .Z(n1825) );
  NAND U2262 ( .A(b[1]), .B(a[79]), .Z(n1826) );
  XOR U2263 ( .A(n1825), .B(n1826), .Z(n1828) );
  XOR U2264 ( .A(n1827), .B(n1828), .Z(n1830) );
  XOR U2265 ( .A(sreg[334]), .B(n1829), .Z(n1824) );
  XNOR U2266 ( .A(n1830), .B(n1824), .Z(c[334]) );
  AND U2267 ( .A(b[0]), .B(a[81]), .Z(n1832) );
  NAND U2268 ( .A(b[1]), .B(a[80]), .Z(n1833) );
  XOR U2269 ( .A(n1832), .B(n1833), .Z(n1835) );
  XOR U2270 ( .A(n1834), .B(n1835), .Z(n1837) );
  XNOR U2271 ( .A(sreg[335]), .B(n1836), .Z(n1831) );
  XNOR U2272 ( .A(n1837), .B(n1831), .Z(c[335]) );
  AND U2273 ( .A(b[0]), .B(a[82]), .Z(n1839) );
  NAND U2274 ( .A(b[1]), .B(a[81]), .Z(n1840) );
  XOR U2275 ( .A(n1839), .B(n1840), .Z(n1842) );
  XOR U2276 ( .A(n1841), .B(n1842), .Z(n1844) );
  XNOR U2277 ( .A(sreg[336]), .B(n1843), .Z(n1838) );
  XNOR U2278 ( .A(n1844), .B(n1838), .Z(c[336]) );
  AND U2279 ( .A(b[0]), .B(a[83]), .Z(n1846) );
  NAND U2280 ( .A(b[1]), .B(a[82]), .Z(n1847) );
  XOR U2281 ( .A(n1846), .B(n1847), .Z(n1849) );
  XOR U2282 ( .A(n1848), .B(n1849), .Z(n1851) );
  XNOR U2283 ( .A(sreg[337]), .B(n1850), .Z(n1845) );
  XNOR U2284 ( .A(n1851), .B(n1845), .Z(c[337]) );
  AND U2285 ( .A(b[0]), .B(a[84]), .Z(n1853) );
  NAND U2286 ( .A(b[1]), .B(a[83]), .Z(n1854) );
  XNOR U2287 ( .A(n1853), .B(n1854), .Z(n1856) );
  XNOR U2288 ( .A(n1855), .B(n1856), .Z(n1858) );
  XOR U2289 ( .A(n1857), .B(sreg[338]), .Z(n1852) );
  XNOR U2290 ( .A(n1858), .B(n1852), .Z(c[338]) );
  AND U2291 ( .A(b[0]), .B(a[85]), .Z(n1860) );
  NAND U2292 ( .A(b[1]), .B(a[84]), .Z(n1861) );
  XOR U2293 ( .A(n1860), .B(n1861), .Z(n1863) );
  XOR U2294 ( .A(n1862), .B(n1863), .Z(n1865) );
  XOR U2295 ( .A(sreg[339]), .B(n1864), .Z(n1859) );
  XNOR U2296 ( .A(n1865), .B(n1859), .Z(c[339]) );
  AND U2297 ( .A(b[0]), .B(a[86]), .Z(n1867) );
  NAND U2298 ( .A(b[1]), .B(a[85]), .Z(n1868) );
  XNOR U2299 ( .A(n1867), .B(n1868), .Z(n1870) );
  XNOR U2300 ( .A(n1869), .B(n1870), .Z(n1872) );
  XOR U2301 ( .A(n1871), .B(sreg[340]), .Z(n1866) );
  XNOR U2302 ( .A(n1872), .B(n1866), .Z(c[340]) );
  AND U2303 ( .A(b[0]), .B(a[87]), .Z(n1874) );
  NAND U2304 ( .A(b[1]), .B(a[86]), .Z(n1875) );
  XOR U2305 ( .A(n1874), .B(n1875), .Z(n1877) );
  XOR U2306 ( .A(n1876), .B(n1877), .Z(n1879) );
  XOR U2307 ( .A(sreg[341]), .B(n1878), .Z(n1873) );
  XNOR U2308 ( .A(n1879), .B(n1873), .Z(c[341]) );
  AND U2309 ( .A(b[0]), .B(a[88]), .Z(n1881) );
  NAND U2310 ( .A(b[1]), .B(a[87]), .Z(n1882) );
  XNOR U2311 ( .A(n1881), .B(n1882), .Z(n1884) );
  XNOR U2312 ( .A(n1883), .B(n1884), .Z(n1886) );
  XOR U2313 ( .A(n1885), .B(sreg[342]), .Z(n1880) );
  XNOR U2314 ( .A(n1886), .B(n1880), .Z(c[342]) );
  AND U2315 ( .A(b[0]), .B(a[89]), .Z(n1888) );
  NAND U2316 ( .A(b[1]), .B(a[88]), .Z(n1889) );
  XOR U2317 ( .A(n1888), .B(n1889), .Z(n1891) );
  XOR U2318 ( .A(n1890), .B(n1891), .Z(n1893) );
  XOR U2319 ( .A(sreg[343]), .B(n1892), .Z(n1887) );
  XNOR U2320 ( .A(n1893), .B(n1887), .Z(c[343]) );
  AND U2321 ( .A(b[0]), .B(a[90]), .Z(n1895) );
  NAND U2322 ( .A(b[1]), .B(a[89]), .Z(n1896) );
  XOR U2323 ( .A(n1895), .B(n1896), .Z(n1898) );
  XOR U2324 ( .A(n1897), .B(n1898), .Z(n1900) );
  XNOR U2325 ( .A(sreg[344]), .B(n1899), .Z(n1894) );
  XNOR U2326 ( .A(n1900), .B(n1894), .Z(c[344]) );
  AND U2327 ( .A(b[0]), .B(a[91]), .Z(n1902) );
  NAND U2328 ( .A(b[1]), .B(a[90]), .Z(n1903) );
  XOR U2329 ( .A(n1902), .B(n1903), .Z(n1905) );
  XOR U2330 ( .A(n1904), .B(n1905), .Z(n1907) );
  XNOR U2331 ( .A(sreg[345]), .B(n1906), .Z(n1901) );
  XNOR U2332 ( .A(n1907), .B(n1901), .Z(c[345]) );
  AND U2333 ( .A(b[0]), .B(a[92]), .Z(n1909) );
  NAND U2334 ( .A(b[1]), .B(a[91]), .Z(n1910) );
  XOR U2335 ( .A(n1909), .B(n1910), .Z(n1912) );
  XOR U2336 ( .A(n1911), .B(n1912), .Z(n1914) );
  XNOR U2337 ( .A(sreg[346]), .B(n1913), .Z(n1908) );
  XNOR U2338 ( .A(n1914), .B(n1908), .Z(c[346]) );
  AND U2339 ( .A(b[0]), .B(a[93]), .Z(n1916) );
  NAND U2340 ( .A(b[1]), .B(a[92]), .Z(n1917) );
  XNOR U2341 ( .A(n1916), .B(n1917), .Z(n1919) );
  XNOR U2342 ( .A(n1918), .B(n1919), .Z(n1921) );
  XOR U2343 ( .A(n1920), .B(sreg[347]), .Z(n1915) );
  XNOR U2344 ( .A(n1921), .B(n1915), .Z(c[347]) );
  AND U2345 ( .A(b[0]), .B(a[94]), .Z(n1923) );
  NAND U2346 ( .A(b[1]), .B(a[93]), .Z(n1924) );
  XOR U2347 ( .A(n1923), .B(n1924), .Z(n1926) );
  XOR U2348 ( .A(n1925), .B(n1926), .Z(n1928) );
  XOR U2349 ( .A(sreg[348]), .B(n1927), .Z(n1922) );
  XNOR U2350 ( .A(n1928), .B(n1922), .Z(c[348]) );
  AND U2351 ( .A(b[0]), .B(a[95]), .Z(n1930) );
  NAND U2352 ( .A(b[1]), .B(a[94]), .Z(n1931) );
  XNOR U2353 ( .A(n1930), .B(n1931), .Z(n1933) );
  XNOR U2354 ( .A(n1932), .B(n1933), .Z(n1935) );
  XOR U2355 ( .A(n1934), .B(sreg[349]), .Z(n1929) );
  XNOR U2356 ( .A(n1935), .B(n1929), .Z(c[349]) );
  AND U2357 ( .A(b[0]), .B(a[96]), .Z(n1937) );
  NAND U2358 ( .A(b[1]), .B(a[95]), .Z(n1938) );
  XOR U2359 ( .A(n1937), .B(n1938), .Z(n1940) );
  XOR U2360 ( .A(n1939), .B(n1940), .Z(n1942) );
  XOR U2361 ( .A(sreg[350]), .B(n1941), .Z(n1936) );
  XNOR U2362 ( .A(n1942), .B(n1936), .Z(c[350]) );
  AND U2363 ( .A(b[0]), .B(a[97]), .Z(n1944) );
  NAND U2364 ( .A(b[1]), .B(a[96]), .Z(n1945) );
  XNOR U2365 ( .A(n1944), .B(n1945), .Z(n1947) );
  XNOR U2366 ( .A(n1946), .B(n1947), .Z(n1949) );
  XOR U2367 ( .A(n1948), .B(sreg[351]), .Z(n1943) );
  XNOR U2368 ( .A(n1949), .B(n1943), .Z(c[351]) );
  AND U2369 ( .A(b[0]), .B(a[98]), .Z(n1951) );
  NAND U2370 ( .A(b[1]), .B(a[97]), .Z(n1952) );
  XOR U2371 ( .A(n1951), .B(n1952), .Z(n1954) );
  XOR U2372 ( .A(n1953), .B(n1954), .Z(n1956) );
  XOR U2373 ( .A(sreg[352]), .B(n1955), .Z(n1950) );
  XNOR U2374 ( .A(n1956), .B(n1950), .Z(c[352]) );
  AND U2375 ( .A(b[0]), .B(a[99]), .Z(n1958) );
  NAND U2376 ( .A(b[1]), .B(a[98]), .Z(n1959) );
  XNOR U2377 ( .A(n1958), .B(n1959), .Z(n1961) );
  XNOR U2378 ( .A(n1960), .B(n1961), .Z(n1963) );
  XOR U2379 ( .A(n1962), .B(sreg[353]), .Z(n1957) );
  XNOR U2380 ( .A(n1963), .B(n1957), .Z(c[353]) );
  AND U2381 ( .A(b[0]), .B(a[100]), .Z(n1965) );
  NAND U2382 ( .A(b[1]), .B(a[99]), .Z(n1966) );
  XOR U2383 ( .A(n1965), .B(n1966), .Z(n1968) );
  XOR U2384 ( .A(n1967), .B(n1968), .Z(n1970) );
  XOR U2385 ( .A(sreg[354]), .B(n1969), .Z(n1964) );
  XNOR U2386 ( .A(n1970), .B(n1964), .Z(c[354]) );
  AND U2387 ( .A(b[0]), .B(a[101]), .Z(n1972) );
  NAND U2388 ( .A(b[1]), .B(a[100]), .Z(n1973) );
  XOR U2389 ( .A(n1972), .B(n1973), .Z(n1975) );
  XOR U2390 ( .A(n1974), .B(n1975), .Z(n1977) );
  XNOR U2391 ( .A(sreg[355]), .B(n1976), .Z(n1971) );
  XNOR U2392 ( .A(n1977), .B(n1971), .Z(c[355]) );
  AND U2393 ( .A(b[0]), .B(a[102]), .Z(n1979) );
  NAND U2394 ( .A(b[1]), .B(a[101]), .Z(n1980) );
  XOR U2395 ( .A(n1979), .B(n1980), .Z(n1982) );
  XOR U2396 ( .A(n1981), .B(n1982), .Z(n1984) );
  XNOR U2397 ( .A(sreg[356]), .B(n1983), .Z(n1978) );
  XNOR U2398 ( .A(n1984), .B(n1978), .Z(c[356]) );
  AND U2399 ( .A(b[0]), .B(a[103]), .Z(n1986) );
  NAND U2400 ( .A(b[1]), .B(a[102]), .Z(n1987) );
  XOR U2401 ( .A(n1986), .B(n1987), .Z(n1989) );
  XOR U2402 ( .A(n1988), .B(n1989), .Z(n1991) );
  XNOR U2403 ( .A(sreg[357]), .B(n1990), .Z(n1985) );
  XNOR U2404 ( .A(n1991), .B(n1985), .Z(c[357]) );
  AND U2405 ( .A(b[0]), .B(a[104]), .Z(n1993) );
  NAND U2406 ( .A(b[1]), .B(a[103]), .Z(n1994) );
  XNOR U2407 ( .A(n1993), .B(n1994), .Z(n1996) );
  XNOR U2408 ( .A(n1995), .B(n1996), .Z(n1998) );
  XOR U2409 ( .A(n1997), .B(sreg[358]), .Z(n1992) );
  XNOR U2410 ( .A(n1998), .B(n1992), .Z(c[358]) );
  AND U2411 ( .A(b[0]), .B(a[105]), .Z(n2000) );
  NAND U2412 ( .A(b[1]), .B(a[104]), .Z(n2001) );
  XNOR U2413 ( .A(n2000), .B(n2001), .Z(n2003) );
  XNOR U2414 ( .A(n2002), .B(n2003), .Z(n2005) );
  XNOR U2415 ( .A(n2004), .B(sreg[359]), .Z(n1999) );
  XNOR U2416 ( .A(n2005), .B(n1999), .Z(c[359]) );
  AND U2417 ( .A(b[0]), .B(a[106]), .Z(n2007) );
  NAND U2418 ( .A(b[1]), .B(a[105]), .Z(n2008) );
  XOR U2419 ( .A(n2007), .B(n2008), .Z(n2010) );
  XOR U2420 ( .A(n2009), .B(n2010), .Z(n2012) );
  XOR U2421 ( .A(sreg[360]), .B(n2011), .Z(n2006) );
  XNOR U2422 ( .A(n2012), .B(n2006), .Z(c[360]) );
  AND U2423 ( .A(b[0]), .B(a[107]), .Z(n2014) );
  NAND U2424 ( .A(b[1]), .B(a[106]), .Z(n2015) );
  XOR U2425 ( .A(n2014), .B(n2015), .Z(n2017) );
  XOR U2426 ( .A(n2016), .B(n2017), .Z(n2019) );
  XNOR U2427 ( .A(sreg[361]), .B(n2018), .Z(n2013) );
  XNOR U2428 ( .A(n2019), .B(n2013), .Z(c[361]) );
  AND U2429 ( .A(b[0]), .B(a[108]), .Z(n2021) );
  NAND U2430 ( .A(b[1]), .B(a[107]), .Z(n2022) );
  XOR U2431 ( .A(n2021), .B(n2022), .Z(n2024) );
  XOR U2432 ( .A(n2023), .B(n2024), .Z(n2026) );
  XNOR U2433 ( .A(sreg[362]), .B(n2025), .Z(n2020) );
  XNOR U2434 ( .A(n2026), .B(n2020), .Z(c[362]) );
  AND U2435 ( .A(b[0]), .B(a[109]), .Z(n2028) );
  NAND U2436 ( .A(b[1]), .B(a[108]), .Z(n2029) );
  XNOR U2437 ( .A(n2028), .B(n2029), .Z(n2031) );
  XNOR U2438 ( .A(n2030), .B(n2031), .Z(n2033) );
  XOR U2439 ( .A(n2032), .B(sreg[363]), .Z(n2027) );
  XNOR U2440 ( .A(n2033), .B(n2027), .Z(c[363]) );
  AND U2441 ( .A(b[0]), .B(a[110]), .Z(n2035) );
  NAND U2442 ( .A(b[1]), .B(a[109]), .Z(n2036) );
  XOR U2443 ( .A(n2035), .B(n2036), .Z(n2038) );
  XOR U2444 ( .A(n2037), .B(n2038), .Z(n2040) );
  XOR U2445 ( .A(sreg[364]), .B(n2039), .Z(n2034) );
  XNOR U2446 ( .A(n2040), .B(n2034), .Z(c[364]) );
  AND U2447 ( .A(b[0]), .B(a[111]), .Z(n2042) );
  NAND U2448 ( .A(b[1]), .B(a[110]), .Z(n2043) );
  XNOR U2449 ( .A(n2042), .B(n2043), .Z(n2045) );
  XNOR U2450 ( .A(n2044), .B(n2045), .Z(n2047) );
  XOR U2451 ( .A(n2046), .B(sreg[365]), .Z(n2041) );
  XNOR U2452 ( .A(n2047), .B(n2041), .Z(c[365]) );
  AND U2453 ( .A(b[0]), .B(a[112]), .Z(n2049) );
  NAND U2454 ( .A(b[1]), .B(a[111]), .Z(n2050) );
  XNOR U2455 ( .A(n2049), .B(n2050), .Z(n2052) );
  XNOR U2456 ( .A(n2051), .B(n2052), .Z(n2054) );
  XNOR U2457 ( .A(n2053), .B(sreg[366]), .Z(n2048) );
  XNOR U2458 ( .A(n2054), .B(n2048), .Z(c[366]) );
  AND U2459 ( .A(b[0]), .B(a[113]), .Z(n2056) );
  NAND U2460 ( .A(b[1]), .B(a[112]), .Z(n2057) );
  XOR U2461 ( .A(n2056), .B(n2057), .Z(n2059) );
  XOR U2462 ( .A(n2058), .B(n2059), .Z(n2061) );
  XOR U2463 ( .A(sreg[367]), .B(n2060), .Z(n2055) );
  XNOR U2464 ( .A(n2061), .B(n2055), .Z(c[367]) );
  AND U2465 ( .A(b[0]), .B(a[114]), .Z(n2063) );
  NAND U2466 ( .A(b[1]), .B(a[113]), .Z(n2064) );
  XOR U2467 ( .A(n2063), .B(n2064), .Z(n2066) );
  XOR U2468 ( .A(n2065), .B(n2066), .Z(n2068) );
  XNOR U2469 ( .A(sreg[368]), .B(n2067), .Z(n2062) );
  XNOR U2470 ( .A(n2068), .B(n2062), .Z(c[368]) );
  AND U2471 ( .A(b[0]), .B(a[115]), .Z(n2070) );
  NAND U2472 ( .A(b[1]), .B(a[114]), .Z(n2071) );
  XOR U2473 ( .A(n2070), .B(n2071), .Z(n2073) );
  XOR U2474 ( .A(n2072), .B(n2073), .Z(n2075) );
  XNOR U2475 ( .A(sreg[369]), .B(n2074), .Z(n2069) );
  XNOR U2476 ( .A(n2075), .B(n2069), .Z(c[369]) );
  AND U2477 ( .A(b[0]), .B(a[116]), .Z(n2077) );
  NAND U2478 ( .A(b[1]), .B(a[115]), .Z(n2078) );
  XNOR U2479 ( .A(n2077), .B(n2078), .Z(n2080) );
  XNOR U2480 ( .A(n2079), .B(n2080), .Z(n2082) );
  XOR U2481 ( .A(n2081), .B(sreg[370]), .Z(n2076) );
  XNOR U2482 ( .A(n2082), .B(n2076), .Z(c[370]) );
  AND U2483 ( .A(b[0]), .B(a[117]), .Z(n2084) );
  NAND U2484 ( .A(b[1]), .B(a[116]), .Z(n2085) );
  XOR U2485 ( .A(n2084), .B(n2085), .Z(n2087) );
  XOR U2486 ( .A(n2086), .B(n2087), .Z(n2089) );
  XOR U2487 ( .A(sreg[371]), .B(n2088), .Z(n2083) );
  XNOR U2488 ( .A(n2089), .B(n2083), .Z(c[371]) );
  AND U2489 ( .A(b[0]), .B(a[118]), .Z(n2091) );
  NAND U2490 ( .A(b[1]), .B(a[117]), .Z(n2092) );
  XOR U2491 ( .A(n2091), .B(n2092), .Z(n2094) );
  XOR U2492 ( .A(n2093), .B(n2094), .Z(n2096) );
  XNOR U2493 ( .A(sreg[372]), .B(n2095), .Z(n2090) );
  XNOR U2494 ( .A(n2096), .B(n2090), .Z(c[372]) );
  AND U2495 ( .A(b[0]), .B(a[119]), .Z(n2098) );
  NAND U2496 ( .A(b[1]), .B(a[118]), .Z(n2099) );
  XOR U2497 ( .A(n2098), .B(n2099), .Z(n2101) );
  XOR U2498 ( .A(n2100), .B(n2101), .Z(n2103) );
  XNOR U2499 ( .A(sreg[373]), .B(n2102), .Z(n2097) );
  XNOR U2500 ( .A(n2103), .B(n2097), .Z(c[373]) );
  AND U2501 ( .A(b[0]), .B(a[120]), .Z(n2105) );
  NAND U2502 ( .A(b[1]), .B(a[119]), .Z(n2106) );
  XNOR U2503 ( .A(n2105), .B(n2106), .Z(n2108) );
  XNOR U2504 ( .A(n2107), .B(n2108), .Z(n2110) );
  XOR U2505 ( .A(n2109), .B(sreg[374]), .Z(n2104) );
  XNOR U2506 ( .A(n2110), .B(n2104), .Z(c[374]) );
  AND U2507 ( .A(b[0]), .B(a[121]), .Z(n2112) );
  NAND U2508 ( .A(b[1]), .B(a[120]), .Z(n2113) );
  XOR U2509 ( .A(n2112), .B(n2113), .Z(n2115) );
  XOR U2510 ( .A(n2114), .B(n2115), .Z(n2117) );
  XOR U2511 ( .A(sreg[375]), .B(n2116), .Z(n2111) );
  XNOR U2512 ( .A(n2117), .B(n2111), .Z(c[375]) );
  AND U2513 ( .A(b[0]), .B(a[122]), .Z(n2119) );
  NAND U2514 ( .A(b[1]), .B(a[121]), .Z(n2120) );
  XOR U2515 ( .A(n2119), .B(n2120), .Z(n2122) );
  XOR U2516 ( .A(n2121), .B(n2122), .Z(n2124) );
  XNOR U2517 ( .A(sreg[376]), .B(n2123), .Z(n2118) );
  XNOR U2518 ( .A(n2124), .B(n2118), .Z(c[376]) );
  AND U2519 ( .A(b[0]), .B(a[123]), .Z(n2126) );
  NAND U2520 ( .A(b[1]), .B(a[122]), .Z(n2127) );
  XOR U2521 ( .A(n2126), .B(n2127), .Z(n2129) );
  XOR U2522 ( .A(n2128), .B(n2129), .Z(n2131) );
  XNOR U2523 ( .A(sreg[377]), .B(n2130), .Z(n2125) );
  XNOR U2524 ( .A(n2131), .B(n2125), .Z(c[377]) );
  AND U2525 ( .A(b[0]), .B(a[124]), .Z(n2133) );
  NAND U2526 ( .A(b[1]), .B(a[123]), .Z(n2134) );
  XOR U2527 ( .A(n2133), .B(n2134), .Z(n2136) );
  XOR U2528 ( .A(n2135), .B(n2136), .Z(n2138) );
  XNOR U2529 ( .A(sreg[378]), .B(n2137), .Z(n2132) );
  XNOR U2530 ( .A(n2138), .B(n2132), .Z(c[378]) );
  AND U2531 ( .A(b[0]), .B(a[125]), .Z(n2140) );
  NAND U2532 ( .A(b[1]), .B(a[124]), .Z(n2141) );
  XNOR U2533 ( .A(n2140), .B(n2141), .Z(n2143) );
  XNOR U2534 ( .A(n2142), .B(n2143), .Z(n2145) );
  XOR U2535 ( .A(n2144), .B(sreg[379]), .Z(n2139) );
  XNOR U2536 ( .A(n2145), .B(n2139), .Z(c[379]) );
  AND U2537 ( .A(b[0]), .B(a[126]), .Z(n2147) );
  NAND U2538 ( .A(b[1]), .B(a[125]), .Z(n2148) );
  XOR U2539 ( .A(n2147), .B(n2148), .Z(n2150) );
  XOR U2540 ( .A(n2149), .B(n2150), .Z(n2152) );
  XOR U2541 ( .A(sreg[380]), .B(n2151), .Z(n2146) );
  XNOR U2542 ( .A(n2152), .B(n2146), .Z(c[380]) );
  AND U2543 ( .A(b[0]), .B(a[127]), .Z(n2154) );
  NAND U2544 ( .A(b[1]), .B(a[126]), .Z(n2155) );
  XNOR U2545 ( .A(n2154), .B(n2155), .Z(n2157) );
  XNOR U2546 ( .A(n2156), .B(n2157), .Z(n2159) );
  XOR U2547 ( .A(n2158), .B(sreg[381]), .Z(n2153) );
  XNOR U2548 ( .A(n2159), .B(n2153), .Z(c[381]) );
  AND U2549 ( .A(b[0]), .B(a[128]), .Z(n2161) );
  NAND U2550 ( .A(b[1]), .B(a[127]), .Z(n2162) );
  XOR U2551 ( .A(n2161), .B(n2162), .Z(n2164) );
  XOR U2552 ( .A(n2163), .B(n2164), .Z(n2166) );
  XOR U2553 ( .A(sreg[382]), .B(n2165), .Z(n2160) );
  XNOR U2554 ( .A(n2166), .B(n2160), .Z(c[382]) );
  AND U2555 ( .A(b[0]), .B(a[129]), .Z(n2168) );
  NAND U2556 ( .A(b[1]), .B(a[128]), .Z(n2169) );
  XNOR U2557 ( .A(n2168), .B(n2169), .Z(n2171) );
  XNOR U2558 ( .A(n2170), .B(n2171), .Z(n2173) );
  XOR U2559 ( .A(n2172), .B(sreg[383]), .Z(n2167) );
  XNOR U2560 ( .A(n2173), .B(n2167), .Z(c[383]) );
  AND U2561 ( .A(b[0]), .B(a[130]), .Z(n2175) );
  NAND U2562 ( .A(b[1]), .B(a[129]), .Z(n2176) );
  XOR U2563 ( .A(n2175), .B(n2176), .Z(n2178) );
  XOR U2564 ( .A(n2177), .B(n2178), .Z(n2180) );
  XOR U2565 ( .A(sreg[384]), .B(n2179), .Z(n2174) );
  XNOR U2566 ( .A(n2180), .B(n2174), .Z(c[384]) );
  AND U2567 ( .A(b[0]), .B(a[131]), .Z(n2182) );
  NAND U2568 ( .A(b[1]), .B(a[130]), .Z(n2183) );
  XNOR U2569 ( .A(n2182), .B(n2183), .Z(n2185) );
  XNOR U2570 ( .A(n2184), .B(n2185), .Z(n2187) );
  XOR U2571 ( .A(n2186), .B(sreg[385]), .Z(n2181) );
  XNOR U2572 ( .A(n2187), .B(n2181), .Z(c[385]) );
  AND U2573 ( .A(b[0]), .B(a[132]), .Z(n2189) );
  NAND U2574 ( .A(b[1]), .B(a[131]), .Z(n2190) );
  XOR U2575 ( .A(n2189), .B(n2190), .Z(n2192) );
  XOR U2576 ( .A(n2191), .B(n2192), .Z(n2194) );
  XOR U2577 ( .A(sreg[386]), .B(n2193), .Z(n2188) );
  XNOR U2578 ( .A(n2194), .B(n2188), .Z(c[386]) );
  AND U2579 ( .A(b[0]), .B(a[133]), .Z(n2196) );
  NAND U2580 ( .A(b[1]), .B(a[132]), .Z(n2197) );
  XNOR U2581 ( .A(n2196), .B(n2197), .Z(n2199) );
  XNOR U2582 ( .A(n2198), .B(n2199), .Z(n2201) );
  XOR U2583 ( .A(n2200), .B(sreg[387]), .Z(n2195) );
  XNOR U2584 ( .A(n2201), .B(n2195), .Z(c[387]) );
  AND U2585 ( .A(b[0]), .B(a[134]), .Z(n2203) );
  NAND U2586 ( .A(b[1]), .B(a[133]), .Z(n2204) );
  XOR U2587 ( .A(n2203), .B(n2204), .Z(n2206) );
  XOR U2588 ( .A(n2205), .B(n2206), .Z(n2208) );
  XOR U2589 ( .A(sreg[388]), .B(n2207), .Z(n2202) );
  XNOR U2590 ( .A(n2208), .B(n2202), .Z(c[388]) );
  AND U2591 ( .A(b[0]), .B(a[135]), .Z(n2210) );
  NAND U2592 ( .A(b[1]), .B(a[134]), .Z(n2211) );
  XOR U2593 ( .A(n2210), .B(n2211), .Z(n2213) );
  XOR U2594 ( .A(n2212), .B(n2213), .Z(n2215) );
  XNOR U2595 ( .A(sreg[389]), .B(n2214), .Z(n2209) );
  XNOR U2596 ( .A(n2215), .B(n2209), .Z(c[389]) );
  AND U2597 ( .A(b[0]), .B(a[136]), .Z(n2217) );
  NAND U2598 ( .A(b[1]), .B(a[135]), .Z(n2218) );
  XOR U2599 ( .A(n2217), .B(n2218), .Z(n2220) );
  XOR U2600 ( .A(n2219), .B(n2220), .Z(n2222) );
  XNOR U2601 ( .A(sreg[390]), .B(n2221), .Z(n2216) );
  XNOR U2602 ( .A(n2222), .B(n2216), .Z(c[390]) );
  AND U2603 ( .A(b[0]), .B(a[137]), .Z(n2224) );
  NAND U2604 ( .A(b[1]), .B(a[136]), .Z(n2225) );
  XNOR U2605 ( .A(n2224), .B(n2225), .Z(n2227) );
  XNOR U2606 ( .A(n2226), .B(n2227), .Z(n2229) );
  XOR U2607 ( .A(n2228), .B(sreg[391]), .Z(n2223) );
  XNOR U2608 ( .A(n2229), .B(n2223), .Z(c[391]) );
  AND U2609 ( .A(b[0]), .B(a[138]), .Z(n2231) );
  NAND U2610 ( .A(b[1]), .B(a[137]), .Z(n2232) );
  XOR U2611 ( .A(n2231), .B(n2232), .Z(n2234) );
  XOR U2612 ( .A(n2233), .B(n2234), .Z(n2236) );
  XOR U2613 ( .A(sreg[392]), .B(n2235), .Z(n2230) );
  XNOR U2614 ( .A(n2236), .B(n2230), .Z(c[392]) );
  AND U2615 ( .A(b[0]), .B(a[139]), .Z(n2238) );
  NAND U2616 ( .A(b[1]), .B(a[138]), .Z(n2239) );
  XOR U2617 ( .A(n2238), .B(n2239), .Z(n2241) );
  XOR U2618 ( .A(n2240), .B(n2241), .Z(n2243) );
  XNOR U2619 ( .A(sreg[393]), .B(n2242), .Z(n2237) );
  XNOR U2620 ( .A(n2243), .B(n2237), .Z(c[393]) );
  AND U2621 ( .A(b[0]), .B(a[140]), .Z(n2245) );
  NAND U2622 ( .A(b[1]), .B(a[139]), .Z(n2246) );
  XOR U2623 ( .A(n2245), .B(n2246), .Z(n2248) );
  XOR U2624 ( .A(n2247), .B(n2248), .Z(n2250) );
  XNOR U2625 ( .A(sreg[394]), .B(n2249), .Z(n2244) );
  XNOR U2626 ( .A(n2250), .B(n2244), .Z(c[394]) );
  AND U2627 ( .A(b[0]), .B(a[141]), .Z(n2252) );
  NAND U2628 ( .A(b[1]), .B(a[140]), .Z(n2253) );
  XNOR U2629 ( .A(n2252), .B(n2253), .Z(n2255) );
  XNOR U2630 ( .A(n2254), .B(n2255), .Z(n2257) );
  XOR U2631 ( .A(n2256), .B(sreg[395]), .Z(n2251) );
  XNOR U2632 ( .A(n2257), .B(n2251), .Z(c[395]) );
  AND U2633 ( .A(b[0]), .B(a[142]), .Z(n2259) );
  NAND U2634 ( .A(b[1]), .B(a[141]), .Z(n2260) );
  XOR U2635 ( .A(n2259), .B(n2260), .Z(n2262) );
  XOR U2636 ( .A(n2261), .B(n2262), .Z(n2264) );
  XOR U2637 ( .A(sreg[396]), .B(n2263), .Z(n2258) );
  XNOR U2638 ( .A(n2264), .B(n2258), .Z(c[396]) );
  AND U2639 ( .A(b[0]), .B(a[143]), .Z(n2266) );
  NAND U2640 ( .A(b[1]), .B(a[142]), .Z(n2267) );
  XNOR U2641 ( .A(n2266), .B(n2267), .Z(n2269) );
  XNOR U2642 ( .A(n2268), .B(n2269), .Z(n2271) );
  XOR U2643 ( .A(n2270), .B(sreg[397]), .Z(n2265) );
  XNOR U2644 ( .A(n2271), .B(n2265), .Z(c[397]) );
  AND U2645 ( .A(b[0]), .B(a[144]), .Z(n2273) );
  NAND U2646 ( .A(b[1]), .B(a[143]), .Z(n2274) );
  XOR U2647 ( .A(n2273), .B(n2274), .Z(n2276) );
  XOR U2648 ( .A(n2275), .B(n2276), .Z(n2278) );
  XOR U2649 ( .A(sreg[398]), .B(n2277), .Z(n2272) );
  XNOR U2650 ( .A(n2278), .B(n2272), .Z(c[398]) );
  AND U2651 ( .A(b[0]), .B(a[145]), .Z(n2280) );
  NAND U2652 ( .A(b[1]), .B(a[144]), .Z(n2281) );
  XNOR U2653 ( .A(n2280), .B(n2281), .Z(n2283) );
  XNOR U2654 ( .A(n2282), .B(n2283), .Z(n2285) );
  XOR U2655 ( .A(n2284), .B(sreg[399]), .Z(n2279) );
  XNOR U2656 ( .A(n2285), .B(n2279), .Z(c[399]) );
  AND U2657 ( .A(b[0]), .B(a[146]), .Z(n2287) );
  NAND U2658 ( .A(b[1]), .B(a[145]), .Z(n2288) );
  XOR U2659 ( .A(n2287), .B(n2288), .Z(n2290) );
  XOR U2660 ( .A(n2289), .B(n2290), .Z(n2292) );
  XOR U2661 ( .A(sreg[400]), .B(n2291), .Z(n2286) );
  XNOR U2662 ( .A(n2292), .B(n2286), .Z(c[400]) );
  AND U2663 ( .A(b[0]), .B(a[147]), .Z(n2294) );
  NAND U2664 ( .A(b[1]), .B(a[146]), .Z(n2295) );
  XOR U2665 ( .A(n2294), .B(n2295), .Z(n2297) );
  XOR U2666 ( .A(n2296), .B(n2297), .Z(n2299) );
  XNOR U2667 ( .A(sreg[401]), .B(n2298), .Z(n2293) );
  XNOR U2668 ( .A(n2299), .B(n2293), .Z(c[401]) );
  AND U2669 ( .A(b[0]), .B(a[148]), .Z(n2301) );
  NAND U2670 ( .A(b[1]), .B(a[147]), .Z(n2302) );
  XNOR U2671 ( .A(n2301), .B(n2302), .Z(n2304) );
  XNOR U2672 ( .A(n2303), .B(n2304), .Z(n2306) );
  XOR U2673 ( .A(n2305), .B(sreg[402]), .Z(n2300) );
  XNOR U2674 ( .A(n2306), .B(n2300), .Z(c[402]) );
  AND U2675 ( .A(b[0]), .B(a[149]), .Z(n2308) );
  NAND U2676 ( .A(b[1]), .B(a[148]), .Z(n2309) );
  XOR U2677 ( .A(n2308), .B(n2309), .Z(n2311) );
  XOR U2678 ( .A(n2310), .B(n2311), .Z(n2313) );
  XOR U2679 ( .A(sreg[403]), .B(n2312), .Z(n2307) );
  XNOR U2680 ( .A(n2313), .B(n2307), .Z(c[403]) );
  AND U2681 ( .A(b[0]), .B(a[150]), .Z(n2315) );
  NAND U2682 ( .A(b[1]), .B(a[149]), .Z(n2316) );
  XNOR U2683 ( .A(n2315), .B(n2316), .Z(n2318) );
  XNOR U2684 ( .A(n2317), .B(n2318), .Z(n2320) );
  XOR U2685 ( .A(n2319), .B(sreg[404]), .Z(n2314) );
  XNOR U2686 ( .A(n2320), .B(n2314), .Z(c[404]) );
  AND U2687 ( .A(b[0]), .B(a[151]), .Z(n2322) );
  NAND U2688 ( .A(b[1]), .B(a[150]), .Z(n2323) );
  XNOR U2689 ( .A(n2322), .B(n2323), .Z(n2325) );
  XNOR U2690 ( .A(n2324), .B(n2325), .Z(n2327) );
  XNOR U2691 ( .A(n2326), .B(sreg[405]), .Z(n2321) );
  XNOR U2692 ( .A(n2327), .B(n2321), .Z(c[405]) );
  AND U2693 ( .A(b[0]), .B(a[152]), .Z(n2329) );
  NAND U2694 ( .A(b[1]), .B(a[151]), .Z(n2330) );
  XNOR U2695 ( .A(n2329), .B(n2330), .Z(n2332) );
  XNOR U2696 ( .A(n2331), .B(n2332), .Z(n2334) );
  XNOR U2697 ( .A(n2333), .B(sreg[406]), .Z(n2328) );
  XNOR U2698 ( .A(n2334), .B(n2328), .Z(c[406]) );
  AND U2699 ( .A(b[0]), .B(a[153]), .Z(n2336) );
  NAND U2700 ( .A(b[1]), .B(a[152]), .Z(n2337) );
  XOR U2701 ( .A(n2336), .B(n2337), .Z(n2339) );
  XOR U2702 ( .A(n2338), .B(n2339), .Z(n2341) );
  XOR U2703 ( .A(sreg[407]), .B(n2340), .Z(n2335) );
  XNOR U2704 ( .A(n2341), .B(n2335), .Z(c[407]) );
  AND U2705 ( .A(b[0]), .B(a[154]), .Z(n2343) );
  NAND U2706 ( .A(b[1]), .B(a[153]), .Z(n2344) );
  XOR U2707 ( .A(n2343), .B(n2344), .Z(n2346) );
  XOR U2708 ( .A(n2345), .B(n2346), .Z(n2348) );
  XNOR U2709 ( .A(sreg[408]), .B(n2347), .Z(n2342) );
  XNOR U2710 ( .A(n2348), .B(n2342), .Z(c[408]) );
  AND U2711 ( .A(b[0]), .B(a[155]), .Z(n2350) );
  NAND U2712 ( .A(b[1]), .B(a[154]), .Z(n2351) );
  XOR U2713 ( .A(n2350), .B(n2351), .Z(n2353) );
  XOR U2714 ( .A(n2352), .B(n2353), .Z(n2355) );
  XNOR U2715 ( .A(sreg[409]), .B(n2354), .Z(n2349) );
  XNOR U2716 ( .A(n2355), .B(n2349), .Z(c[409]) );
  AND U2717 ( .A(b[0]), .B(a[156]), .Z(n2357) );
  NAND U2718 ( .A(b[1]), .B(a[155]), .Z(n2358) );
  XOR U2719 ( .A(n2357), .B(n2358), .Z(n2360) );
  XOR U2720 ( .A(n2359), .B(n2360), .Z(n2362) );
  XNOR U2721 ( .A(sreg[410]), .B(n2361), .Z(n2356) );
  XNOR U2722 ( .A(n2362), .B(n2356), .Z(c[410]) );
  AND U2723 ( .A(b[0]), .B(a[157]), .Z(n2364) );
  NAND U2724 ( .A(b[1]), .B(a[156]), .Z(n2365) );
  XOR U2725 ( .A(n2364), .B(n2365), .Z(n2367) );
  XOR U2726 ( .A(n2366), .B(n2367), .Z(n2369) );
  XNOR U2727 ( .A(sreg[411]), .B(n2368), .Z(n2363) );
  XNOR U2728 ( .A(n2369), .B(n2363), .Z(c[411]) );
  AND U2729 ( .A(b[0]), .B(a[158]), .Z(n2371) );
  NAND U2730 ( .A(b[1]), .B(a[157]), .Z(n2372) );
  XOR U2731 ( .A(n2371), .B(n2372), .Z(n2374) );
  XOR U2732 ( .A(n2373), .B(n2374), .Z(n2376) );
  XNOR U2733 ( .A(sreg[412]), .B(n2375), .Z(n2370) );
  XNOR U2734 ( .A(n2376), .B(n2370), .Z(c[412]) );
  AND U2735 ( .A(b[0]), .B(a[159]), .Z(n2378) );
  NAND U2736 ( .A(b[1]), .B(a[158]), .Z(n2379) );
  XNOR U2737 ( .A(n2378), .B(n2379), .Z(n2381) );
  XNOR U2738 ( .A(n2380), .B(n2381), .Z(n2383) );
  XOR U2739 ( .A(n2382), .B(sreg[413]), .Z(n2377) );
  XNOR U2740 ( .A(n2383), .B(n2377), .Z(c[413]) );
  AND U2741 ( .A(b[0]), .B(a[160]), .Z(n2385) );
  NAND U2742 ( .A(b[1]), .B(a[159]), .Z(n2386) );
  XOR U2743 ( .A(n2385), .B(n2386), .Z(n2388) );
  XOR U2744 ( .A(n2387), .B(n2388), .Z(n2390) );
  XOR U2745 ( .A(sreg[414]), .B(n2389), .Z(n2384) );
  XNOR U2746 ( .A(n2390), .B(n2384), .Z(c[414]) );
  AND U2747 ( .A(b[0]), .B(a[161]), .Z(n2392) );
  NAND U2748 ( .A(b[1]), .B(a[160]), .Z(n2393) );
  XNOR U2749 ( .A(n2392), .B(n2393), .Z(n2395) );
  XNOR U2750 ( .A(n2394), .B(n2395), .Z(n2397) );
  XOR U2751 ( .A(n2396), .B(sreg[415]), .Z(n2391) );
  XNOR U2752 ( .A(n2397), .B(n2391), .Z(c[415]) );
  AND U2753 ( .A(b[0]), .B(a[162]), .Z(n2399) );
  NAND U2754 ( .A(b[1]), .B(a[161]), .Z(n2400) );
  XOR U2755 ( .A(n2399), .B(n2400), .Z(n2402) );
  XOR U2756 ( .A(n2401), .B(n2402), .Z(n2404) );
  XOR U2757 ( .A(sreg[416]), .B(n2403), .Z(n2398) );
  XNOR U2758 ( .A(n2404), .B(n2398), .Z(c[416]) );
  AND U2759 ( .A(b[0]), .B(a[163]), .Z(n2406) );
  NAND U2760 ( .A(b[1]), .B(a[162]), .Z(n2407) );
  XNOR U2761 ( .A(n2406), .B(n2407), .Z(n2409) );
  XNOR U2762 ( .A(n2408), .B(n2409), .Z(n2411) );
  XOR U2763 ( .A(n2410), .B(sreg[417]), .Z(n2405) );
  XNOR U2764 ( .A(n2411), .B(n2405), .Z(c[417]) );
  AND U2765 ( .A(b[0]), .B(a[164]), .Z(n2413) );
  NAND U2766 ( .A(b[1]), .B(a[163]), .Z(n2414) );
  XOR U2767 ( .A(n2413), .B(n2414), .Z(n2416) );
  XOR U2768 ( .A(n2415), .B(n2416), .Z(n2418) );
  XOR U2769 ( .A(sreg[418]), .B(n2417), .Z(n2412) );
  XNOR U2770 ( .A(n2418), .B(n2412), .Z(c[418]) );
  AND U2771 ( .A(b[0]), .B(a[165]), .Z(n2420) );
  NAND U2772 ( .A(b[1]), .B(a[164]), .Z(n2421) );
  XNOR U2773 ( .A(n2420), .B(n2421), .Z(n2423) );
  XNOR U2774 ( .A(n2422), .B(n2423), .Z(n2425) );
  XOR U2775 ( .A(n2424), .B(sreg[419]), .Z(n2419) );
  XNOR U2776 ( .A(n2425), .B(n2419), .Z(c[419]) );
  AND U2777 ( .A(b[0]), .B(a[166]), .Z(n2427) );
  NAND U2778 ( .A(b[1]), .B(a[165]), .Z(n2428) );
  XOR U2779 ( .A(n2427), .B(n2428), .Z(n2430) );
  XOR U2780 ( .A(n2429), .B(n2430), .Z(n2432) );
  XOR U2781 ( .A(sreg[420]), .B(n2431), .Z(n2426) );
  XNOR U2782 ( .A(n2432), .B(n2426), .Z(c[420]) );
  AND U2783 ( .A(b[0]), .B(a[167]), .Z(n2434) );
  NAND U2784 ( .A(b[1]), .B(a[166]), .Z(n2435) );
  XOR U2785 ( .A(n2434), .B(n2435), .Z(n2437) );
  XOR U2786 ( .A(n2436), .B(n2437), .Z(n2439) );
  XNOR U2787 ( .A(sreg[421]), .B(n2438), .Z(n2433) );
  XNOR U2788 ( .A(n2439), .B(n2433), .Z(c[421]) );
  AND U2789 ( .A(b[0]), .B(a[168]), .Z(n2441) );
  NAND U2790 ( .A(b[1]), .B(a[167]), .Z(n2442) );
  XOR U2791 ( .A(n2441), .B(n2442), .Z(n2444) );
  XOR U2792 ( .A(n2443), .B(n2444), .Z(n2446) );
  XNOR U2793 ( .A(sreg[422]), .B(n2445), .Z(n2440) );
  XNOR U2794 ( .A(n2446), .B(n2440), .Z(c[422]) );
  AND U2795 ( .A(b[0]), .B(a[169]), .Z(n2448) );
  NAND U2796 ( .A(b[1]), .B(a[168]), .Z(n2449) );
  XOR U2797 ( .A(n2448), .B(n2449), .Z(n2451) );
  XOR U2798 ( .A(n2450), .B(n2451), .Z(n2453) );
  XNOR U2799 ( .A(sreg[423]), .B(n2452), .Z(n2447) );
  XNOR U2800 ( .A(n2453), .B(n2447), .Z(c[423]) );
  AND U2801 ( .A(b[0]), .B(a[170]), .Z(n2455) );
  NAND U2802 ( .A(b[1]), .B(a[169]), .Z(n2456) );
  XOR U2803 ( .A(n2455), .B(n2456), .Z(n2458) );
  XOR U2804 ( .A(n2457), .B(n2458), .Z(n2460) );
  XNOR U2805 ( .A(sreg[424]), .B(n2459), .Z(n2454) );
  XNOR U2806 ( .A(n2460), .B(n2454), .Z(c[424]) );
  AND U2807 ( .A(b[0]), .B(a[171]), .Z(n2462) );
  NAND U2808 ( .A(b[1]), .B(a[170]), .Z(n2463) );
  XOR U2809 ( .A(n2462), .B(n2463), .Z(n2465) );
  XOR U2810 ( .A(n2464), .B(n2465), .Z(n2467) );
  XNOR U2811 ( .A(sreg[425]), .B(n2466), .Z(n2461) );
  XNOR U2812 ( .A(n2467), .B(n2461), .Z(c[425]) );
  AND U2813 ( .A(b[0]), .B(a[172]), .Z(n2469) );
  NAND U2814 ( .A(b[1]), .B(a[171]), .Z(n2470) );
  XOR U2815 ( .A(n2469), .B(n2470), .Z(n2472) );
  XOR U2816 ( .A(n2471), .B(n2472), .Z(n2474) );
  XNOR U2817 ( .A(sreg[426]), .B(n2473), .Z(n2468) );
  XNOR U2818 ( .A(n2474), .B(n2468), .Z(c[426]) );
  AND U2819 ( .A(b[0]), .B(a[173]), .Z(n2476) );
  NAND U2820 ( .A(b[1]), .B(a[172]), .Z(n2477) );
  XNOR U2821 ( .A(n2476), .B(n2477), .Z(n2479) );
  XNOR U2822 ( .A(n2478), .B(n2479), .Z(n2481) );
  XOR U2823 ( .A(n2480), .B(sreg[427]), .Z(n2475) );
  XNOR U2824 ( .A(n2481), .B(n2475), .Z(c[427]) );
  AND U2825 ( .A(b[0]), .B(a[174]), .Z(n2483) );
  NAND U2826 ( .A(b[1]), .B(a[173]), .Z(n2484) );
  XNOR U2827 ( .A(n2483), .B(n2484), .Z(n2486) );
  XNOR U2828 ( .A(n2485), .B(n2486), .Z(n2488) );
  XNOR U2829 ( .A(n2487), .B(sreg[428]), .Z(n2482) );
  XNOR U2830 ( .A(n2488), .B(n2482), .Z(c[428]) );
  AND U2831 ( .A(b[0]), .B(a[175]), .Z(n2490) );
  NAND U2832 ( .A(b[1]), .B(a[174]), .Z(n2491) );
  XNOR U2833 ( .A(n2490), .B(n2491), .Z(n2493) );
  XNOR U2834 ( .A(n2492), .B(n2493), .Z(n2495) );
  XNOR U2835 ( .A(n2494), .B(sreg[429]), .Z(n2489) );
  XNOR U2836 ( .A(n2495), .B(n2489), .Z(c[429]) );
  AND U2837 ( .A(b[0]), .B(a[176]), .Z(n2497) );
  NAND U2838 ( .A(b[1]), .B(a[175]), .Z(n2498) );
  XOR U2839 ( .A(n2497), .B(n2498), .Z(n2500) );
  XOR U2840 ( .A(n2499), .B(n2500), .Z(n2502) );
  XOR U2841 ( .A(sreg[430]), .B(n2501), .Z(n2496) );
  XNOR U2842 ( .A(n2502), .B(n2496), .Z(c[430]) );
  AND U2843 ( .A(b[0]), .B(a[177]), .Z(n2504) );
  NAND U2844 ( .A(b[1]), .B(a[176]), .Z(n2505) );
  XOR U2845 ( .A(n2504), .B(n2505), .Z(n2507) );
  XOR U2846 ( .A(n2506), .B(n2507), .Z(n2509) );
  XNOR U2847 ( .A(sreg[431]), .B(n2508), .Z(n2503) );
  XNOR U2848 ( .A(n2509), .B(n2503), .Z(c[431]) );
  AND U2849 ( .A(b[0]), .B(a[178]), .Z(n2511) );
  NAND U2850 ( .A(b[1]), .B(a[177]), .Z(n2512) );
  XOR U2851 ( .A(n2511), .B(n2512), .Z(n2514) );
  XOR U2852 ( .A(n2513), .B(n2514), .Z(n2516) );
  XNOR U2853 ( .A(sreg[432]), .B(n2515), .Z(n2510) );
  XNOR U2854 ( .A(n2516), .B(n2510), .Z(c[432]) );
  AND U2855 ( .A(b[0]), .B(a[179]), .Z(n2518) );
  NAND U2856 ( .A(b[1]), .B(a[178]), .Z(n2519) );
  XOR U2857 ( .A(n2518), .B(n2519), .Z(n2521) );
  XOR U2858 ( .A(n2520), .B(n2521), .Z(n2523) );
  XNOR U2859 ( .A(sreg[433]), .B(n2522), .Z(n2517) );
  XNOR U2860 ( .A(n2523), .B(n2517), .Z(c[433]) );
  AND U2861 ( .A(b[0]), .B(a[180]), .Z(n2525) );
  NAND U2862 ( .A(b[1]), .B(a[179]), .Z(n2526) );
  XNOR U2863 ( .A(n2525), .B(n2526), .Z(n2528) );
  XNOR U2864 ( .A(n2527), .B(n2528), .Z(n2530) );
  XOR U2865 ( .A(n2529), .B(sreg[434]), .Z(n2524) );
  XNOR U2866 ( .A(n2530), .B(n2524), .Z(c[434]) );
  AND U2867 ( .A(b[0]), .B(a[181]), .Z(n2532) );
  NAND U2868 ( .A(b[1]), .B(a[180]), .Z(n2533) );
  XNOR U2869 ( .A(n2532), .B(n2533), .Z(n2535) );
  XNOR U2870 ( .A(n2534), .B(n2535), .Z(n2537) );
  XNOR U2871 ( .A(n2536), .B(sreg[435]), .Z(n2531) );
  XNOR U2872 ( .A(n2537), .B(n2531), .Z(c[435]) );
  AND U2873 ( .A(b[0]), .B(a[182]), .Z(n2539) );
  NAND U2874 ( .A(b[1]), .B(a[181]), .Z(n2540) );
  XNOR U2875 ( .A(n2539), .B(n2540), .Z(n2542) );
  XNOR U2876 ( .A(n2541), .B(n2542), .Z(n2544) );
  XNOR U2877 ( .A(n2543), .B(sreg[436]), .Z(n2538) );
  XNOR U2878 ( .A(n2544), .B(n2538), .Z(c[436]) );
  AND U2879 ( .A(b[0]), .B(a[183]), .Z(n2546) );
  NAND U2880 ( .A(b[1]), .B(a[182]), .Z(n2547) );
  XOR U2881 ( .A(n2546), .B(n2547), .Z(n2549) );
  XOR U2882 ( .A(n2548), .B(n2549), .Z(n2551) );
  XOR U2883 ( .A(sreg[437]), .B(n2550), .Z(n2545) );
  XNOR U2884 ( .A(n2551), .B(n2545), .Z(c[437]) );
  AND U2885 ( .A(b[0]), .B(a[184]), .Z(n2553) );
  NAND U2886 ( .A(b[1]), .B(a[183]), .Z(n2554) );
  XNOR U2887 ( .A(n2553), .B(n2554), .Z(n2556) );
  XNOR U2888 ( .A(n2555), .B(n2556), .Z(n2558) );
  XOR U2889 ( .A(n2557), .B(sreg[438]), .Z(n2552) );
  XNOR U2890 ( .A(n2558), .B(n2552), .Z(c[438]) );
  AND U2891 ( .A(b[0]), .B(a[185]), .Z(n2560) );
  NAND U2892 ( .A(b[1]), .B(a[184]), .Z(n2561) );
  XOR U2893 ( .A(n2560), .B(n2561), .Z(n2563) );
  XOR U2894 ( .A(n2562), .B(n2563), .Z(n2565) );
  XOR U2895 ( .A(sreg[439]), .B(n2564), .Z(n2559) );
  XNOR U2896 ( .A(n2565), .B(n2559), .Z(c[439]) );
  AND U2897 ( .A(b[0]), .B(a[186]), .Z(n2567) );
  NAND U2898 ( .A(b[1]), .B(a[185]), .Z(n2568) );
  XNOR U2899 ( .A(n2567), .B(n2568), .Z(n2570) );
  XNOR U2900 ( .A(n2569), .B(n2570), .Z(n2572) );
  XOR U2901 ( .A(n2571), .B(sreg[440]), .Z(n2566) );
  XNOR U2902 ( .A(n2572), .B(n2566), .Z(c[440]) );
  AND U2903 ( .A(b[0]), .B(a[187]), .Z(n2574) );
  NAND U2904 ( .A(b[1]), .B(a[186]), .Z(n2575) );
  XOR U2905 ( .A(n2574), .B(n2575), .Z(n2577) );
  XOR U2906 ( .A(n2576), .B(n2577), .Z(n2579) );
  XOR U2907 ( .A(sreg[441]), .B(n2578), .Z(n2573) );
  XNOR U2908 ( .A(n2579), .B(n2573), .Z(c[441]) );
  AND U2909 ( .A(b[0]), .B(a[188]), .Z(n2581) );
  NAND U2910 ( .A(b[1]), .B(a[187]), .Z(n2582) );
  XOR U2911 ( .A(n2581), .B(n2582), .Z(n2584) );
  XOR U2912 ( .A(n2583), .B(n2584), .Z(n2586) );
  XNOR U2913 ( .A(sreg[442]), .B(n2585), .Z(n2580) );
  XNOR U2914 ( .A(n2586), .B(n2580), .Z(c[442]) );
  AND U2915 ( .A(b[0]), .B(a[189]), .Z(n2588) );
  NAND U2916 ( .A(b[1]), .B(a[188]), .Z(n2589) );
  XNOR U2917 ( .A(n2588), .B(n2589), .Z(n2591) );
  XNOR U2918 ( .A(n2590), .B(n2591), .Z(n2593) );
  XOR U2919 ( .A(n2592), .B(sreg[443]), .Z(n2587) );
  XNOR U2920 ( .A(n2593), .B(n2587), .Z(c[443]) );
  AND U2921 ( .A(b[0]), .B(a[190]), .Z(n2595) );
  NAND U2922 ( .A(b[1]), .B(a[189]), .Z(n2596) );
  XOR U2923 ( .A(n2595), .B(n2596), .Z(n2598) );
  XOR U2924 ( .A(n2597), .B(n2598), .Z(n2600) );
  XOR U2925 ( .A(sreg[444]), .B(n2599), .Z(n2594) );
  XNOR U2926 ( .A(n2600), .B(n2594), .Z(c[444]) );
  AND U2927 ( .A(b[0]), .B(a[191]), .Z(n2602) );
  NAND U2928 ( .A(b[1]), .B(a[190]), .Z(n2603) );
  XNOR U2929 ( .A(n2602), .B(n2603), .Z(n2605) );
  XNOR U2930 ( .A(n2604), .B(n2605), .Z(n2607) );
  XOR U2931 ( .A(n2606), .B(sreg[445]), .Z(n2601) );
  XNOR U2932 ( .A(n2607), .B(n2601), .Z(c[445]) );
  AND U2933 ( .A(b[0]), .B(a[192]), .Z(n2609) );
  NAND U2934 ( .A(b[1]), .B(a[191]), .Z(n2610) );
  XOR U2935 ( .A(n2609), .B(n2610), .Z(n2612) );
  XOR U2936 ( .A(n2611), .B(n2612), .Z(n2614) );
  XOR U2937 ( .A(sreg[446]), .B(n2613), .Z(n2608) );
  XNOR U2938 ( .A(n2614), .B(n2608), .Z(c[446]) );
  AND U2939 ( .A(b[0]), .B(a[193]), .Z(n2616) );
  NAND U2940 ( .A(b[1]), .B(a[192]), .Z(n2617) );
  XNOR U2941 ( .A(n2616), .B(n2617), .Z(n2619) );
  XNOR U2942 ( .A(n2618), .B(n2619), .Z(n2621) );
  XOR U2943 ( .A(n2620), .B(sreg[447]), .Z(n2615) );
  XNOR U2944 ( .A(n2621), .B(n2615), .Z(c[447]) );
  AND U2945 ( .A(b[0]), .B(a[194]), .Z(n2623) );
  NAND U2946 ( .A(b[1]), .B(a[193]), .Z(n2624) );
  XOR U2947 ( .A(n2623), .B(n2624), .Z(n2626) );
  XOR U2948 ( .A(n2625), .B(n2626), .Z(n2628) );
  XOR U2949 ( .A(sreg[448]), .B(n2627), .Z(n2622) );
  XNOR U2950 ( .A(n2628), .B(n2622), .Z(c[448]) );
  AND U2951 ( .A(b[0]), .B(a[195]), .Z(n2630) );
  NAND U2952 ( .A(b[1]), .B(a[194]), .Z(n2631) );
  XNOR U2953 ( .A(n2630), .B(n2631), .Z(n2633) );
  XNOR U2954 ( .A(n2632), .B(n2633), .Z(n2635) );
  XOR U2955 ( .A(n2634), .B(sreg[449]), .Z(n2629) );
  XNOR U2956 ( .A(n2635), .B(n2629), .Z(c[449]) );
  AND U2957 ( .A(b[0]), .B(a[196]), .Z(n2637) );
  NAND U2958 ( .A(b[1]), .B(a[195]), .Z(n2638) );
  XOR U2959 ( .A(n2637), .B(n2638), .Z(n2640) );
  XOR U2960 ( .A(n2639), .B(n2640), .Z(n2642) );
  XOR U2961 ( .A(sreg[450]), .B(n2641), .Z(n2636) );
  XNOR U2962 ( .A(n2642), .B(n2636), .Z(c[450]) );
  AND U2963 ( .A(b[0]), .B(a[197]), .Z(n2644) );
  NAND U2964 ( .A(b[1]), .B(a[196]), .Z(n2645) );
  XOR U2965 ( .A(n2644), .B(n2645), .Z(n2647) );
  XOR U2966 ( .A(n2646), .B(n2647), .Z(n2649) );
  XNOR U2967 ( .A(sreg[451]), .B(n2648), .Z(n2643) );
  XNOR U2968 ( .A(n2649), .B(n2643), .Z(c[451]) );
  AND U2969 ( .A(b[0]), .B(a[198]), .Z(n2651) );
  NAND U2970 ( .A(b[1]), .B(a[197]), .Z(n2652) );
  XOR U2971 ( .A(n2651), .B(n2652), .Z(n2654) );
  XOR U2972 ( .A(n2653), .B(n2654), .Z(n2656) );
  XNOR U2973 ( .A(sreg[452]), .B(n2655), .Z(n2650) );
  XNOR U2974 ( .A(n2656), .B(n2650), .Z(c[452]) );
  AND U2975 ( .A(b[0]), .B(a[199]), .Z(n2658) );
  NAND U2976 ( .A(b[1]), .B(a[198]), .Z(n2659) );
  XNOR U2977 ( .A(n2658), .B(n2659), .Z(n2661) );
  XNOR U2978 ( .A(n2660), .B(n2661), .Z(n2663) );
  XOR U2979 ( .A(n2662), .B(sreg[453]), .Z(n2657) );
  XNOR U2980 ( .A(n2663), .B(n2657), .Z(c[453]) );
  AND U2981 ( .A(b[0]), .B(a[200]), .Z(n2665) );
  NAND U2982 ( .A(b[1]), .B(a[199]), .Z(n2666) );
  XOR U2983 ( .A(n2665), .B(n2666), .Z(n2668) );
  XOR U2984 ( .A(n2667), .B(n2668), .Z(n2670) );
  XOR U2985 ( .A(sreg[454]), .B(n2669), .Z(n2664) );
  XNOR U2986 ( .A(n2670), .B(n2664), .Z(c[454]) );
  AND U2987 ( .A(b[0]), .B(a[201]), .Z(n2672) );
  NAND U2988 ( .A(b[1]), .B(a[200]), .Z(n2673) );
  XNOR U2989 ( .A(n2672), .B(n2673), .Z(n2675) );
  XNOR U2990 ( .A(n2674), .B(n2675), .Z(n2677) );
  XOR U2991 ( .A(n2676), .B(sreg[455]), .Z(n2671) );
  XNOR U2992 ( .A(n2677), .B(n2671), .Z(c[455]) );
  AND U2993 ( .A(b[0]), .B(a[202]), .Z(n2679) );
  NAND U2994 ( .A(b[1]), .B(a[201]), .Z(n2680) );
  XOR U2995 ( .A(n2679), .B(n2680), .Z(n2682) );
  XOR U2996 ( .A(n2681), .B(n2682), .Z(n2684) );
  XOR U2997 ( .A(sreg[456]), .B(n2683), .Z(n2678) );
  XNOR U2998 ( .A(n2684), .B(n2678), .Z(c[456]) );
  AND U2999 ( .A(b[0]), .B(a[203]), .Z(n2686) );
  NAND U3000 ( .A(b[1]), .B(a[202]), .Z(n2687) );
  XOR U3001 ( .A(n2686), .B(n2687), .Z(n2689) );
  XOR U3002 ( .A(n2688), .B(n2689), .Z(n2691) );
  XNOR U3003 ( .A(sreg[457]), .B(n2690), .Z(n2685) );
  XNOR U3004 ( .A(n2691), .B(n2685), .Z(c[457]) );
  AND U3005 ( .A(b[0]), .B(a[204]), .Z(n2693) );
  NAND U3006 ( .A(b[1]), .B(a[203]), .Z(n2694) );
  XOR U3007 ( .A(n2693), .B(n2694), .Z(n2696) );
  XOR U3008 ( .A(n2695), .B(n2696), .Z(n2698) );
  XNOR U3009 ( .A(sreg[458]), .B(n2697), .Z(n2692) );
  XNOR U3010 ( .A(n2698), .B(n2692), .Z(c[458]) );
  AND U3011 ( .A(b[0]), .B(a[205]), .Z(n2700) );
  NAND U3012 ( .A(b[1]), .B(a[204]), .Z(n2701) );
  XNOR U3013 ( .A(n2700), .B(n2701), .Z(n2703) );
  XNOR U3014 ( .A(n2702), .B(n2703), .Z(n2705) );
  XOR U3015 ( .A(n2704), .B(sreg[459]), .Z(n2699) );
  XNOR U3016 ( .A(n2705), .B(n2699), .Z(c[459]) );
  AND U3017 ( .A(b[0]), .B(a[206]), .Z(n2707) );
  NAND U3018 ( .A(b[1]), .B(a[205]), .Z(n2708) );
  XOR U3019 ( .A(n2707), .B(n2708), .Z(n2710) );
  XOR U3020 ( .A(n2709), .B(n2710), .Z(n2712) );
  XOR U3021 ( .A(sreg[460]), .B(n2711), .Z(n2706) );
  XNOR U3022 ( .A(n2712), .B(n2706), .Z(c[460]) );
  AND U3023 ( .A(b[0]), .B(a[207]), .Z(n2714) );
  NAND U3024 ( .A(b[1]), .B(a[206]), .Z(n2715) );
  XNOR U3025 ( .A(n2714), .B(n2715), .Z(n2717) );
  XNOR U3026 ( .A(n2716), .B(n2717), .Z(n2719) );
  XOR U3027 ( .A(n2718), .B(sreg[461]), .Z(n2713) );
  XNOR U3028 ( .A(n2719), .B(n2713), .Z(c[461]) );
  AND U3029 ( .A(b[0]), .B(a[208]), .Z(n2721) );
  NAND U3030 ( .A(b[1]), .B(a[207]), .Z(n2722) );
  XOR U3031 ( .A(n2721), .B(n2722), .Z(n2724) );
  XOR U3032 ( .A(n2723), .B(n2724), .Z(n2726) );
  XOR U3033 ( .A(sreg[462]), .B(n2725), .Z(n2720) );
  XNOR U3034 ( .A(n2726), .B(n2720), .Z(c[462]) );
  AND U3035 ( .A(b[0]), .B(a[209]), .Z(n2728) );
  NAND U3036 ( .A(b[1]), .B(a[208]), .Z(n2729) );
  XOR U3037 ( .A(n2728), .B(n2729), .Z(n2731) );
  XOR U3038 ( .A(n2730), .B(n2731), .Z(n2733) );
  XNOR U3039 ( .A(sreg[463]), .B(n2732), .Z(n2727) );
  XNOR U3040 ( .A(n2733), .B(n2727), .Z(c[463]) );
  AND U3041 ( .A(b[0]), .B(a[210]), .Z(n2735) );
  NAND U3042 ( .A(b[1]), .B(a[209]), .Z(n2736) );
  XOR U3043 ( .A(n2735), .B(n2736), .Z(n2738) );
  XOR U3044 ( .A(n2737), .B(n2738), .Z(n2740) );
  XNOR U3045 ( .A(sreg[464]), .B(n2739), .Z(n2734) );
  XNOR U3046 ( .A(n2740), .B(n2734), .Z(c[464]) );
  AND U3047 ( .A(b[0]), .B(a[211]), .Z(n2742) );
  NAND U3048 ( .A(b[1]), .B(a[210]), .Z(n2743) );
  XOR U3049 ( .A(n2742), .B(n2743), .Z(n2745) );
  XOR U3050 ( .A(n2744), .B(n2745), .Z(n2747) );
  XNOR U3051 ( .A(sreg[465]), .B(n2746), .Z(n2741) );
  XNOR U3052 ( .A(n2747), .B(n2741), .Z(c[465]) );
  AND U3053 ( .A(b[0]), .B(a[212]), .Z(n2749) );
  NAND U3054 ( .A(b[1]), .B(a[211]), .Z(n2750) );
  XNOR U3055 ( .A(n2749), .B(n2750), .Z(n2752) );
  XNOR U3056 ( .A(n2751), .B(n2752), .Z(n2754) );
  XOR U3057 ( .A(n2753), .B(sreg[466]), .Z(n2748) );
  XNOR U3058 ( .A(n2754), .B(n2748), .Z(c[466]) );
  AND U3059 ( .A(b[0]), .B(a[213]), .Z(n2756) );
  NAND U3060 ( .A(b[1]), .B(a[212]), .Z(n2757) );
  XOR U3061 ( .A(n2756), .B(n2757), .Z(n2759) );
  XOR U3062 ( .A(n2758), .B(n2759), .Z(n2761) );
  XOR U3063 ( .A(sreg[467]), .B(n2760), .Z(n2755) );
  XNOR U3064 ( .A(n2761), .B(n2755), .Z(c[467]) );
  AND U3065 ( .A(b[0]), .B(a[214]), .Z(n2763) );
  NAND U3066 ( .A(b[1]), .B(a[213]), .Z(n2764) );
  XNOR U3067 ( .A(n2763), .B(n2764), .Z(n2766) );
  XNOR U3068 ( .A(n2765), .B(n2766), .Z(n2768) );
  XOR U3069 ( .A(n2767), .B(sreg[468]), .Z(n2762) );
  XNOR U3070 ( .A(n2768), .B(n2762), .Z(c[468]) );
  AND U3071 ( .A(b[0]), .B(a[215]), .Z(n2770) );
  NAND U3072 ( .A(b[1]), .B(a[214]), .Z(n2771) );
  XOR U3073 ( .A(n2770), .B(n2771), .Z(n2773) );
  XOR U3074 ( .A(n2772), .B(n2773), .Z(n2775) );
  XOR U3075 ( .A(sreg[469]), .B(n2774), .Z(n2769) );
  XNOR U3076 ( .A(n2775), .B(n2769), .Z(c[469]) );
  AND U3077 ( .A(b[0]), .B(a[216]), .Z(n2777) );
  NAND U3078 ( .A(b[1]), .B(a[215]), .Z(n2778) );
  XOR U3079 ( .A(n2777), .B(n2778), .Z(n2780) );
  XOR U3080 ( .A(n2779), .B(n2780), .Z(n2782) );
  XNOR U3081 ( .A(sreg[470]), .B(n2781), .Z(n2776) );
  XNOR U3082 ( .A(n2782), .B(n2776), .Z(c[470]) );
  AND U3083 ( .A(b[0]), .B(a[217]), .Z(n2784) );
  NAND U3084 ( .A(b[1]), .B(a[216]), .Z(n2785) );
  XOR U3085 ( .A(n2784), .B(n2785), .Z(n2787) );
  XOR U3086 ( .A(n2786), .B(n2787), .Z(n2789) );
  XNOR U3087 ( .A(sreg[471]), .B(n2788), .Z(n2783) );
  XNOR U3088 ( .A(n2789), .B(n2783), .Z(c[471]) );
  AND U3089 ( .A(b[0]), .B(a[218]), .Z(n2791) );
  NAND U3090 ( .A(b[1]), .B(a[217]), .Z(n2792) );
  XOR U3091 ( .A(n2791), .B(n2792), .Z(n2794) );
  XOR U3092 ( .A(n2793), .B(n2794), .Z(n2796) );
  XNOR U3093 ( .A(sreg[472]), .B(n2795), .Z(n2790) );
  XNOR U3094 ( .A(n2796), .B(n2790), .Z(c[472]) );
  AND U3095 ( .A(b[0]), .B(a[219]), .Z(n2798) );
  NAND U3096 ( .A(b[1]), .B(a[218]), .Z(n2799) );
  XOR U3097 ( .A(n2798), .B(n2799), .Z(n2801) );
  XOR U3098 ( .A(n2800), .B(n2801), .Z(n2803) );
  XNOR U3099 ( .A(sreg[473]), .B(n2802), .Z(n2797) );
  XNOR U3100 ( .A(n2803), .B(n2797), .Z(c[473]) );
  AND U3101 ( .A(b[0]), .B(a[220]), .Z(n2805) );
  NAND U3102 ( .A(b[1]), .B(a[219]), .Z(n2806) );
  XOR U3103 ( .A(n2805), .B(n2806), .Z(n2808) );
  XOR U3104 ( .A(n2807), .B(n2808), .Z(n2810) );
  XNOR U3105 ( .A(sreg[474]), .B(n2809), .Z(n2804) );
  XNOR U3106 ( .A(n2810), .B(n2804), .Z(c[474]) );
  AND U3107 ( .A(b[0]), .B(a[221]), .Z(n2812) );
  NAND U3108 ( .A(b[1]), .B(a[220]), .Z(n2813) );
  XNOR U3109 ( .A(n2812), .B(n2813), .Z(n2815) );
  XNOR U3110 ( .A(n2814), .B(n2815), .Z(n2817) );
  XOR U3111 ( .A(n2816), .B(sreg[475]), .Z(n2811) );
  XNOR U3112 ( .A(n2817), .B(n2811), .Z(c[475]) );
  AND U3113 ( .A(b[0]), .B(a[222]), .Z(n2819) );
  NAND U3114 ( .A(b[1]), .B(a[221]), .Z(n2820) );
  XNOR U3115 ( .A(n2819), .B(n2820), .Z(n2822) );
  XNOR U3116 ( .A(n2821), .B(n2822), .Z(n2824) );
  XNOR U3117 ( .A(n2823), .B(sreg[476]), .Z(n2818) );
  XNOR U3118 ( .A(n2824), .B(n2818), .Z(c[476]) );
  AND U3119 ( .A(b[0]), .B(a[223]), .Z(n2826) );
  NAND U3120 ( .A(b[1]), .B(a[222]), .Z(n2827) );
  XNOR U3121 ( .A(n2826), .B(n2827), .Z(n2829) );
  XNOR U3122 ( .A(n2828), .B(n2829), .Z(n2831) );
  XNOR U3123 ( .A(n2830), .B(sreg[477]), .Z(n2825) );
  XNOR U3124 ( .A(n2831), .B(n2825), .Z(c[477]) );
  AND U3125 ( .A(b[0]), .B(a[224]), .Z(n2833) );
  NAND U3126 ( .A(b[1]), .B(a[223]), .Z(n2834) );
  XOR U3127 ( .A(n2833), .B(n2834), .Z(n2836) );
  XOR U3128 ( .A(n2835), .B(n2836), .Z(n2838) );
  XOR U3129 ( .A(sreg[478]), .B(n2837), .Z(n2832) );
  XNOR U3130 ( .A(n2838), .B(n2832), .Z(c[478]) );
  AND U3131 ( .A(b[0]), .B(a[225]), .Z(n2840) );
  NAND U3132 ( .A(b[1]), .B(a[224]), .Z(n2841) );
  XNOR U3133 ( .A(n2840), .B(n2841), .Z(n2843) );
  XNOR U3134 ( .A(n2842), .B(n2843), .Z(n2845) );
  XOR U3135 ( .A(n2844), .B(sreg[479]), .Z(n2839) );
  XNOR U3136 ( .A(n2845), .B(n2839), .Z(c[479]) );
  AND U3137 ( .A(b[0]), .B(a[226]), .Z(n2847) );
  NAND U3138 ( .A(b[1]), .B(a[225]), .Z(n2848) );
  XOR U3139 ( .A(n2847), .B(n2848), .Z(n2850) );
  XOR U3140 ( .A(n2849), .B(n2850), .Z(n2852) );
  XOR U3141 ( .A(sreg[480]), .B(n2851), .Z(n2846) );
  XNOR U3142 ( .A(n2852), .B(n2846), .Z(c[480]) );
  AND U3143 ( .A(b[0]), .B(a[227]), .Z(n2854) );
  NAND U3144 ( .A(b[1]), .B(a[226]), .Z(n2855) );
  XOR U3145 ( .A(n2854), .B(n2855), .Z(n2857) );
  XOR U3146 ( .A(n2856), .B(n2857), .Z(n2859) );
  XNOR U3147 ( .A(sreg[481]), .B(n2858), .Z(n2853) );
  XNOR U3148 ( .A(n2859), .B(n2853), .Z(c[481]) );
  AND U3149 ( .A(b[0]), .B(a[228]), .Z(n2861) );
  NAND U3150 ( .A(b[1]), .B(a[227]), .Z(n2862) );
  XNOR U3151 ( .A(n2861), .B(n2862), .Z(n2864) );
  XNOR U3152 ( .A(n2863), .B(n2864), .Z(n2866) );
  XOR U3153 ( .A(n2865), .B(sreg[482]), .Z(n2860) );
  XNOR U3154 ( .A(n2866), .B(n2860), .Z(c[482]) );
  AND U3155 ( .A(b[0]), .B(a[229]), .Z(n2868) );
  NAND U3156 ( .A(b[1]), .B(a[228]), .Z(n2869) );
  XOR U3157 ( .A(n2868), .B(n2869), .Z(n2871) );
  XOR U3158 ( .A(n2870), .B(n2871), .Z(n2873) );
  XOR U3159 ( .A(sreg[483]), .B(n2872), .Z(n2867) );
  XNOR U3160 ( .A(n2873), .B(n2867), .Z(c[483]) );
  AND U3161 ( .A(b[0]), .B(a[230]), .Z(n2875) );
  NAND U3162 ( .A(b[1]), .B(a[229]), .Z(n2876) );
  XOR U3163 ( .A(n2875), .B(n2876), .Z(n2878) );
  XOR U3164 ( .A(n2877), .B(n2878), .Z(n2880) );
  XNOR U3165 ( .A(sreg[484]), .B(n2879), .Z(n2874) );
  XNOR U3166 ( .A(n2880), .B(n2874), .Z(c[484]) );
  AND U3167 ( .A(b[0]), .B(a[231]), .Z(n2882) );
  NAND U3168 ( .A(b[1]), .B(a[230]), .Z(n2883) );
  XNOR U3169 ( .A(n2882), .B(n2883), .Z(n2885) );
  XNOR U3170 ( .A(n2884), .B(n2885), .Z(n2887) );
  XOR U3171 ( .A(n2886), .B(sreg[485]), .Z(n2881) );
  XNOR U3172 ( .A(n2887), .B(n2881), .Z(c[485]) );
  AND U3173 ( .A(b[0]), .B(a[232]), .Z(n2889) );
  NAND U3174 ( .A(b[1]), .B(a[231]), .Z(n2890) );
  XNOR U3175 ( .A(n2889), .B(n2890), .Z(n2892) );
  XNOR U3176 ( .A(n2891), .B(n2892), .Z(n2894) );
  XNOR U3177 ( .A(n2893), .B(sreg[486]), .Z(n2888) );
  XNOR U3178 ( .A(n2894), .B(n2888), .Z(c[486]) );
  AND U3179 ( .A(b[0]), .B(a[233]), .Z(n2896) );
  NAND U3180 ( .A(b[1]), .B(a[232]), .Z(n2897) );
  XNOR U3181 ( .A(n2896), .B(n2897), .Z(n2899) );
  XNOR U3182 ( .A(n2898), .B(n2899), .Z(n2901) );
  XNOR U3183 ( .A(n2900), .B(sreg[487]), .Z(n2895) );
  XNOR U3184 ( .A(n2901), .B(n2895), .Z(c[487]) );
  AND U3185 ( .A(b[0]), .B(a[234]), .Z(n2903) );
  NAND U3186 ( .A(b[1]), .B(a[233]), .Z(n2904) );
  XOR U3187 ( .A(n2903), .B(n2904), .Z(n2906) );
  XOR U3188 ( .A(n2905), .B(n2906), .Z(n2908) );
  XOR U3189 ( .A(sreg[488]), .B(n2907), .Z(n2902) );
  XNOR U3190 ( .A(n2908), .B(n2902), .Z(c[488]) );
  AND U3191 ( .A(b[0]), .B(a[235]), .Z(n2910) );
  NAND U3192 ( .A(b[1]), .B(a[234]), .Z(n2911) );
  XOR U3193 ( .A(n2910), .B(n2911), .Z(n2913) );
  XOR U3194 ( .A(n2912), .B(n2913), .Z(n2915) );
  XNOR U3195 ( .A(sreg[489]), .B(n2914), .Z(n2909) );
  XNOR U3196 ( .A(n2915), .B(n2909), .Z(c[489]) );
  AND U3197 ( .A(b[0]), .B(a[236]), .Z(n2917) );
  NAND U3198 ( .A(b[1]), .B(a[235]), .Z(n2918) );
  XOR U3199 ( .A(n2917), .B(n2918), .Z(n2920) );
  XOR U3200 ( .A(n2919), .B(n2920), .Z(n2922) );
  XNOR U3201 ( .A(sreg[490]), .B(n2921), .Z(n2916) );
  XNOR U3202 ( .A(n2922), .B(n2916), .Z(c[490]) );
  AND U3203 ( .A(b[0]), .B(a[237]), .Z(n2924) );
  NAND U3204 ( .A(b[1]), .B(a[236]), .Z(n2925) );
  XOR U3205 ( .A(n2924), .B(n2925), .Z(n2927) );
  XOR U3206 ( .A(n2926), .B(n2927), .Z(n2929) );
  XNOR U3207 ( .A(sreg[491]), .B(n2928), .Z(n2923) );
  XNOR U3208 ( .A(n2929), .B(n2923), .Z(c[491]) );
  AND U3209 ( .A(b[0]), .B(a[238]), .Z(n2931) );
  NAND U3210 ( .A(b[1]), .B(a[237]), .Z(n2932) );
  XOR U3211 ( .A(n2931), .B(n2932), .Z(n2934) );
  XOR U3212 ( .A(n2933), .B(n2934), .Z(n2936) );
  XNOR U3213 ( .A(sreg[492]), .B(n2935), .Z(n2930) );
  XNOR U3214 ( .A(n2936), .B(n2930), .Z(c[492]) );
  AND U3215 ( .A(b[0]), .B(a[239]), .Z(n2938) );
  NAND U3216 ( .A(b[1]), .B(a[238]), .Z(n2939) );
  XNOR U3217 ( .A(n2938), .B(n2939), .Z(n2941) );
  XNOR U3218 ( .A(n2940), .B(n2941), .Z(n2943) );
  XOR U3219 ( .A(n2942), .B(sreg[493]), .Z(n2937) );
  XNOR U3220 ( .A(n2943), .B(n2937), .Z(c[493]) );
  AND U3221 ( .A(b[0]), .B(a[240]), .Z(n2945) );
  NAND U3222 ( .A(b[1]), .B(a[239]), .Z(n2946) );
  XOR U3223 ( .A(n2945), .B(n2946), .Z(n2948) );
  XOR U3224 ( .A(n2947), .B(n2948), .Z(n2950) );
  XOR U3225 ( .A(sreg[494]), .B(n2949), .Z(n2944) );
  XNOR U3226 ( .A(n2950), .B(n2944), .Z(c[494]) );
  AND U3227 ( .A(b[0]), .B(a[241]), .Z(n2952) );
  NAND U3228 ( .A(b[1]), .B(a[240]), .Z(n2953) );
  XOR U3229 ( .A(n2952), .B(n2953), .Z(n2955) );
  XOR U3230 ( .A(n2954), .B(n2955), .Z(n2957) );
  XNOR U3231 ( .A(sreg[495]), .B(n2956), .Z(n2951) );
  XNOR U3232 ( .A(n2957), .B(n2951), .Z(c[495]) );
  AND U3233 ( .A(b[0]), .B(a[242]), .Z(n2959) );
  NAND U3234 ( .A(b[1]), .B(a[241]), .Z(n2960) );
  XOR U3235 ( .A(n2959), .B(n2960), .Z(n2962) );
  XOR U3236 ( .A(n2961), .B(n2962), .Z(n2964) );
  XNOR U3237 ( .A(sreg[496]), .B(n2963), .Z(n2958) );
  XNOR U3238 ( .A(n2964), .B(n2958), .Z(c[496]) );
  AND U3239 ( .A(b[0]), .B(a[243]), .Z(n2966) );
  NAND U3240 ( .A(b[1]), .B(a[242]), .Z(n2967) );
  XOR U3241 ( .A(n2966), .B(n2967), .Z(n2969) );
  XOR U3242 ( .A(n2968), .B(n2969), .Z(n2971) );
  XNOR U3243 ( .A(sreg[497]), .B(n2970), .Z(n2965) );
  XNOR U3244 ( .A(n2971), .B(n2965), .Z(c[497]) );
  AND U3245 ( .A(b[0]), .B(a[244]), .Z(n2973) );
  NAND U3246 ( .A(b[1]), .B(a[243]), .Z(n2974) );
  XNOR U3247 ( .A(n2973), .B(n2974), .Z(n2976) );
  XNOR U3248 ( .A(n2975), .B(n2976), .Z(n2978) );
  XOR U3249 ( .A(n2977), .B(sreg[498]), .Z(n2972) );
  XNOR U3250 ( .A(n2978), .B(n2972), .Z(c[498]) );
  AND U3251 ( .A(b[0]), .B(a[245]), .Z(n2980) );
  NAND U3252 ( .A(b[1]), .B(a[244]), .Z(n2981) );
  XOR U3253 ( .A(n2980), .B(n2981), .Z(n2983) );
  XOR U3254 ( .A(n2982), .B(n2983), .Z(n2985) );
  XOR U3255 ( .A(sreg[499]), .B(n2984), .Z(n2979) );
  XNOR U3256 ( .A(n2985), .B(n2979), .Z(c[499]) );
  AND U3257 ( .A(b[0]), .B(a[246]), .Z(n2987) );
  NAND U3258 ( .A(b[1]), .B(a[245]), .Z(n2988) );
  XNOR U3259 ( .A(n2987), .B(n2988), .Z(n2990) );
  XNOR U3260 ( .A(n2989), .B(n2990), .Z(n2992) );
  XOR U3261 ( .A(n2991), .B(sreg[500]), .Z(n2986) );
  XNOR U3262 ( .A(n2992), .B(n2986), .Z(c[500]) );
  AND U3263 ( .A(b[0]), .B(a[247]), .Z(n2994) );
  NAND U3264 ( .A(b[1]), .B(a[246]), .Z(n2995) );
  XOR U3265 ( .A(n2994), .B(n2995), .Z(n2997) );
  XOR U3266 ( .A(n2996), .B(n2997), .Z(n2999) );
  XOR U3267 ( .A(sreg[501]), .B(n2998), .Z(n2993) );
  XNOR U3268 ( .A(n2999), .B(n2993), .Z(c[501]) );
  AND U3269 ( .A(b[0]), .B(a[248]), .Z(n3001) );
  NAND U3270 ( .A(b[1]), .B(a[247]), .Z(n3002) );
  XNOR U3271 ( .A(n3001), .B(n3002), .Z(n3004) );
  XNOR U3272 ( .A(n3003), .B(n3004), .Z(n3006) );
  XOR U3273 ( .A(n3005), .B(sreg[502]), .Z(n3000) );
  XNOR U3274 ( .A(n3006), .B(n3000), .Z(c[502]) );
  AND U3275 ( .A(b[0]), .B(a[249]), .Z(n3008) );
  NAND U3276 ( .A(b[1]), .B(a[248]), .Z(n3009) );
  XOR U3277 ( .A(n3008), .B(n3009), .Z(n3011) );
  XOR U3278 ( .A(n3010), .B(n3011), .Z(n3013) );
  XOR U3279 ( .A(sreg[503]), .B(n3012), .Z(n3007) );
  XNOR U3280 ( .A(n3013), .B(n3007), .Z(c[503]) );
  AND U3281 ( .A(b[0]), .B(a[250]), .Z(n3015) );
  NAND U3282 ( .A(b[1]), .B(a[249]), .Z(n3016) );
  XOR U3283 ( .A(n3015), .B(n3016), .Z(n3018) );
  XOR U3284 ( .A(n3017), .B(n3018), .Z(n3020) );
  XNOR U3285 ( .A(sreg[504]), .B(n3019), .Z(n3014) );
  XNOR U3286 ( .A(n3020), .B(n3014), .Z(c[504]) );
  AND U3287 ( .A(b[0]), .B(a[251]), .Z(n3022) );
  NAND U3288 ( .A(b[1]), .B(a[250]), .Z(n3023) );
  XOR U3289 ( .A(n3022), .B(n3023), .Z(n3025) );
  XOR U3290 ( .A(n3024), .B(n3025), .Z(n3027) );
  XNOR U3291 ( .A(sreg[505]), .B(n3026), .Z(n3021) );
  XNOR U3292 ( .A(n3027), .B(n3021), .Z(c[505]) );
  AND U3293 ( .A(b[0]), .B(a[252]), .Z(n3029) );
  NAND U3294 ( .A(b[1]), .B(a[251]), .Z(n3030) );
  XOR U3295 ( .A(n3029), .B(n3030), .Z(n3032) );
  XOR U3296 ( .A(n3031), .B(n3032), .Z(n3034) );
  XNOR U3297 ( .A(sreg[506]), .B(n3033), .Z(n3028) );
  XNOR U3298 ( .A(n3034), .B(n3028), .Z(c[506]) );
  AND U3299 ( .A(b[0]), .B(a[253]), .Z(n3036) );
  NAND U3300 ( .A(b[1]), .B(a[252]), .Z(n3037) );
  XNOR U3301 ( .A(n3036), .B(n3037), .Z(n3039) );
  XNOR U3302 ( .A(n3038), .B(n3039), .Z(n3041) );
  XOR U3303 ( .A(n3040), .B(sreg[507]), .Z(n3035) );
  XNOR U3304 ( .A(n3041), .B(n3035), .Z(c[507]) );
  AND U3305 ( .A(b[0]), .B(a[254]), .Z(n3053) );
  NAND U3306 ( .A(b[1]), .B(a[253]), .Z(n3043) );
  XOR U3307 ( .A(n3053), .B(n3043), .Z(n3045) );
  XOR U3308 ( .A(n3044), .B(n3045), .Z(n3049) );
  XOR U3309 ( .A(sreg[508]), .B(n3048), .Z(n3042) );
  XNOR U3310 ( .A(n3049), .B(n3042), .Z(c[508]) );
  AND U3311 ( .A(b[0]), .B(a[255]), .Z(n3047) );
  NAND U3312 ( .A(a[254]), .B(b[1]), .Z(n3046) );
  XNOR U3313 ( .A(n3047), .B(n3046), .Z(n3054) );
  XNOR U3314 ( .A(n3055), .B(n3054), .Z(n3052) );
  XOR U3315 ( .A(n3051), .B(sreg[509]), .Z(n3050) );
  XNOR U3316 ( .A(n3052), .B(n3050), .Z(c[509]) );
  AND U3317 ( .A(b[1]), .B(a[255]), .Z(n3061) );
  XNOR U3318 ( .A(n3061), .B(n3060), .Z(n3058) );
  NAND U3319 ( .A(n3053), .B(n3061), .Z(n3057) );
  NAND U3320 ( .A(n3055), .B(n3054), .Z(n3056) );
  AND U3321 ( .A(n3057), .B(n3056), .Z(n3059) );
  XNOR U3322 ( .A(n3058), .B(n3059), .Z(c[510]) );
  NAND U3323 ( .A(n3059), .B(n3058), .Z(n3063) );
  NANDN U3324 ( .A(n3061), .B(n3060), .Z(n3062) );
  AND U3325 ( .A(n3063), .B(n3062), .Z(c[511]) );
endmodule

