
module hamming_N16000_CC4_DW01_add_0 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57;

  XOR U1 ( .A(n1), .B(n2), .Z(SUM[9]) );
  XNOR U2 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[8]) );
  XNOR U4 ( .A(B[8]), .B(A[8]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[7]) );
  XNOR U6 ( .A(B[7]), .B(A[7]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[6]) );
  XNOR U8 ( .A(B[6]), .B(A[6]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[5]) );
  XNOR U10 ( .A(B[5]), .B(A[5]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[3]) );
  XNOR U14 ( .A(B[3]), .B(A[3]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U16 ( .A(B[2]), .B(A[2]), .Z(n16) );
  XOR U17 ( .A(n17), .B(n18), .Z(SUM[1]) );
  XOR U18 ( .A(B[1]), .B(A[1]), .Z(n18) );
  XOR U19 ( .A(A[13]), .B(n19), .Z(SUM[13]) );
  ANDN U20 ( .B(A[12]), .A(n20), .Z(n19) );
  XNOR U21 ( .A(A[12]), .B(n20), .Z(SUM[12]) );
  AND U22 ( .A(n21), .B(n22), .Z(n20) );
  NAND U23 ( .A(n23), .B(B[11]), .Z(n22) );
  NANDN U24 ( .A(A[11]), .B(n24), .Z(n23) );
  NANDN U25 ( .A(n24), .B(A[11]), .Z(n21) );
  XOR U26 ( .A(n24), .B(n25), .Z(SUM[11]) );
  XNOR U27 ( .A(B[11]), .B(A[11]), .Z(n25) );
  AND U28 ( .A(n26), .B(n27), .Z(n24) );
  NAND U29 ( .A(n28), .B(B[10]), .Z(n27) );
  NANDN U30 ( .A(A[10]), .B(n29), .Z(n28) );
  NANDN U31 ( .A(n29), .B(A[10]), .Z(n26) );
  XOR U32 ( .A(n29), .B(n30), .Z(SUM[10]) );
  XNOR U33 ( .A(B[10]), .B(A[10]), .Z(n30) );
  AND U34 ( .A(n31), .B(n32), .Z(n29) );
  NAND U35 ( .A(n33), .B(B[9]), .Z(n32) );
  NANDN U36 ( .A(A[9]), .B(n1), .Z(n33) );
  NANDN U37 ( .A(n1), .B(A[9]), .Z(n31) );
  AND U38 ( .A(n34), .B(n35), .Z(n1) );
  NAND U39 ( .A(n36), .B(B[8]), .Z(n35) );
  NANDN U40 ( .A(A[8]), .B(n3), .Z(n36) );
  NANDN U41 ( .A(n3), .B(A[8]), .Z(n34) );
  AND U42 ( .A(n37), .B(n38), .Z(n3) );
  NAND U43 ( .A(n39), .B(B[7]), .Z(n38) );
  NANDN U44 ( .A(A[7]), .B(n5), .Z(n39) );
  NANDN U45 ( .A(n5), .B(A[7]), .Z(n37) );
  AND U46 ( .A(n40), .B(n41), .Z(n5) );
  NAND U47 ( .A(n42), .B(B[6]), .Z(n41) );
  NANDN U48 ( .A(A[6]), .B(n7), .Z(n42) );
  NANDN U49 ( .A(n7), .B(A[6]), .Z(n40) );
  AND U50 ( .A(n43), .B(n44), .Z(n7) );
  NAND U51 ( .A(n45), .B(B[5]), .Z(n44) );
  NANDN U52 ( .A(A[5]), .B(n9), .Z(n45) );
  NANDN U53 ( .A(n9), .B(A[5]), .Z(n43) );
  AND U54 ( .A(n46), .B(n47), .Z(n9) );
  NAND U55 ( .A(n48), .B(B[4]), .Z(n47) );
  NANDN U56 ( .A(A[4]), .B(n11), .Z(n48) );
  NANDN U57 ( .A(n11), .B(A[4]), .Z(n46) );
  AND U58 ( .A(n49), .B(n50), .Z(n11) );
  NAND U59 ( .A(n51), .B(B[3]), .Z(n50) );
  NANDN U60 ( .A(A[3]), .B(n13), .Z(n51) );
  NANDN U61 ( .A(n13), .B(A[3]), .Z(n49) );
  AND U62 ( .A(n52), .B(n53), .Z(n13) );
  NAND U63 ( .A(n54), .B(B[2]), .Z(n53) );
  NANDN U64 ( .A(A[2]), .B(n15), .Z(n54) );
  NANDN U65 ( .A(n15), .B(A[2]), .Z(n52) );
  AND U66 ( .A(n55), .B(n56), .Z(n15) );
  NAND U67 ( .A(n57), .B(B[1]), .Z(n56) );
  OR U68 ( .A(n17), .B(A[1]), .Z(n57) );
  NAND U69 ( .A(n17), .B(A[1]), .Z(n55) );
  AND U70 ( .A(B[0]), .B(A[0]), .Z(n17) );
  XOR U71 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_1 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52;

  IV U1 ( .A(B[11]), .Z(n1) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[9]) );
  XNOR U3 ( .A(B[9]), .B(A[9]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[8]) );
  XNOR U5 ( .A(B[8]), .B(A[8]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[7]) );
  XNOR U7 ( .A(B[7]), .B(A[7]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[6]) );
  XNOR U9 ( .A(B[6]), .B(A[6]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XNOR U11 ( .A(B[5]), .B(A[5]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[4]) );
  XNOR U13 ( .A(B[4]), .B(A[4]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[3]) );
  XNOR U15 ( .A(B[3]), .B(A[3]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[2]) );
  XNOR U17 ( .A(B[2]), .B(A[2]), .Z(n17) );
  XOR U18 ( .A(n18), .B(n19), .Z(SUM[1]) );
  XOR U19 ( .A(B[1]), .B(A[1]), .Z(n19) );
  XOR U20 ( .A(n20), .B(n1), .Z(SUM[11]) );
  AND U21 ( .A(n21), .B(n22), .Z(n20) );
  NAND U22 ( .A(n23), .B(B[10]), .Z(n22) );
  NANDN U23 ( .A(A[10]), .B(n24), .Z(n23) );
  NANDN U24 ( .A(n24), .B(A[10]), .Z(n21) );
  XOR U25 ( .A(n24), .B(n25), .Z(SUM[10]) );
  XNOR U26 ( .A(B[10]), .B(A[10]), .Z(n25) );
  AND U27 ( .A(n26), .B(n27), .Z(n24) );
  NAND U28 ( .A(n28), .B(B[9]), .Z(n27) );
  NANDN U29 ( .A(A[9]), .B(n2), .Z(n28) );
  NANDN U30 ( .A(n2), .B(A[9]), .Z(n26) );
  AND U31 ( .A(n29), .B(n30), .Z(n2) );
  NAND U32 ( .A(n31), .B(B[8]), .Z(n30) );
  NANDN U33 ( .A(A[8]), .B(n4), .Z(n31) );
  NANDN U34 ( .A(n4), .B(A[8]), .Z(n29) );
  AND U35 ( .A(n32), .B(n33), .Z(n4) );
  NAND U36 ( .A(n34), .B(B[7]), .Z(n33) );
  NANDN U37 ( .A(A[7]), .B(n6), .Z(n34) );
  NANDN U38 ( .A(n6), .B(A[7]), .Z(n32) );
  AND U39 ( .A(n35), .B(n36), .Z(n6) );
  NAND U40 ( .A(n37), .B(B[6]), .Z(n36) );
  NANDN U41 ( .A(A[6]), .B(n8), .Z(n37) );
  NANDN U42 ( .A(n8), .B(A[6]), .Z(n35) );
  AND U43 ( .A(n38), .B(n39), .Z(n8) );
  NAND U44 ( .A(n40), .B(B[5]), .Z(n39) );
  NANDN U45 ( .A(A[5]), .B(n10), .Z(n40) );
  NANDN U46 ( .A(n10), .B(A[5]), .Z(n38) );
  AND U47 ( .A(n41), .B(n42), .Z(n10) );
  NAND U48 ( .A(n43), .B(B[4]), .Z(n42) );
  NANDN U49 ( .A(A[4]), .B(n12), .Z(n43) );
  NANDN U50 ( .A(n12), .B(A[4]), .Z(n41) );
  AND U51 ( .A(n44), .B(n45), .Z(n12) );
  NAND U52 ( .A(n46), .B(B[3]), .Z(n45) );
  NANDN U53 ( .A(A[3]), .B(n14), .Z(n46) );
  NANDN U54 ( .A(n14), .B(A[3]), .Z(n44) );
  AND U55 ( .A(n47), .B(n48), .Z(n14) );
  NAND U56 ( .A(n49), .B(B[2]), .Z(n48) );
  NANDN U57 ( .A(A[2]), .B(n16), .Z(n49) );
  NANDN U58 ( .A(n16), .B(A[2]), .Z(n47) );
  AND U59 ( .A(n50), .B(n51), .Z(n16) );
  NAND U60 ( .A(n52), .B(B[1]), .Z(n51) );
  OR U61 ( .A(n18), .B(A[1]), .Z(n52) );
  NAND U62 ( .A(n18), .B(A[1]), .Z(n50) );
  AND U63 ( .A(B[0]), .B(A[0]), .Z(n18) );
  XOR U64 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_2 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51;

  NAND U1 ( .A(n20), .B(n21), .Z(SUM[11]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[9]) );
  XNOR U3 ( .A(B[9]), .B(A[9]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[8]) );
  XNOR U5 ( .A(B[8]), .B(A[8]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[7]) );
  XNOR U7 ( .A(B[7]), .B(A[7]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[6]) );
  XNOR U9 ( .A(B[6]), .B(A[6]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XNOR U11 ( .A(B[5]), .B(A[5]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[4]) );
  XNOR U13 ( .A(B[4]), .B(A[4]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[3]) );
  XNOR U15 ( .A(B[3]), .B(A[3]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[2]) );
  XNOR U17 ( .A(B[2]), .B(A[2]), .Z(n17) );
  XOR U18 ( .A(n18), .B(n19), .Z(SUM[1]) );
  XOR U19 ( .A(B[1]), .B(A[1]), .Z(n19) );
  NAND U20 ( .A(n22), .B(B[10]), .Z(n21) );
  NANDN U21 ( .A(A[10]), .B(n23), .Z(n22) );
  NANDN U22 ( .A(n23), .B(A[10]), .Z(n20) );
  XOR U23 ( .A(n23), .B(n24), .Z(SUM[10]) );
  XNOR U24 ( .A(B[10]), .B(A[10]), .Z(n24) );
  AND U25 ( .A(n25), .B(n26), .Z(n23) );
  NAND U26 ( .A(n27), .B(B[9]), .Z(n26) );
  NANDN U27 ( .A(A[9]), .B(n2), .Z(n27) );
  NANDN U28 ( .A(n2), .B(A[9]), .Z(n25) );
  AND U29 ( .A(n28), .B(n29), .Z(n2) );
  NAND U30 ( .A(n30), .B(B[8]), .Z(n29) );
  NANDN U31 ( .A(A[8]), .B(n4), .Z(n30) );
  NANDN U32 ( .A(n4), .B(A[8]), .Z(n28) );
  AND U33 ( .A(n31), .B(n32), .Z(n4) );
  NAND U34 ( .A(n33), .B(B[7]), .Z(n32) );
  NANDN U35 ( .A(A[7]), .B(n6), .Z(n33) );
  NANDN U36 ( .A(n6), .B(A[7]), .Z(n31) );
  AND U37 ( .A(n34), .B(n35), .Z(n6) );
  NAND U38 ( .A(n36), .B(B[6]), .Z(n35) );
  NANDN U39 ( .A(A[6]), .B(n8), .Z(n36) );
  NANDN U40 ( .A(n8), .B(A[6]), .Z(n34) );
  AND U41 ( .A(n37), .B(n38), .Z(n8) );
  NAND U42 ( .A(n39), .B(B[5]), .Z(n38) );
  NANDN U43 ( .A(A[5]), .B(n10), .Z(n39) );
  NANDN U44 ( .A(n10), .B(A[5]), .Z(n37) );
  AND U45 ( .A(n40), .B(n41), .Z(n10) );
  NAND U46 ( .A(n42), .B(B[4]), .Z(n41) );
  NANDN U47 ( .A(A[4]), .B(n12), .Z(n42) );
  NANDN U48 ( .A(n12), .B(A[4]), .Z(n40) );
  AND U49 ( .A(n43), .B(n44), .Z(n12) );
  NAND U50 ( .A(n45), .B(B[3]), .Z(n44) );
  NANDN U51 ( .A(A[3]), .B(n14), .Z(n45) );
  NANDN U52 ( .A(n14), .B(A[3]), .Z(n43) );
  AND U53 ( .A(n46), .B(n47), .Z(n14) );
  NAND U54 ( .A(n48), .B(B[2]), .Z(n47) );
  NANDN U55 ( .A(A[2]), .B(n16), .Z(n48) );
  NANDN U56 ( .A(n16), .B(A[2]), .Z(n46) );
  AND U57 ( .A(n49), .B(n50), .Z(n16) );
  NAND U58 ( .A(n51), .B(B[1]), .Z(n50) );
  OR U59 ( .A(n18), .B(A[1]), .Z(n51) );
  NAND U60 ( .A(n18), .B(A[1]), .Z(n49) );
  AND U61 ( .A(B[0]), .B(A[0]), .Z(n18) );
  XOR U62 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_3 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46;

  NAND U1 ( .A(n20), .B(n21), .Z(SUM[10]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[9]) );
  XNOR U3 ( .A(B[9]), .B(A[9]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[8]) );
  XNOR U5 ( .A(B[8]), .B(A[8]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[7]) );
  XNOR U7 ( .A(B[7]), .B(A[7]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[6]) );
  XNOR U9 ( .A(B[6]), .B(A[6]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XNOR U11 ( .A(B[5]), .B(A[5]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[4]) );
  XNOR U13 ( .A(B[4]), .B(A[4]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[3]) );
  XNOR U15 ( .A(B[3]), .B(A[3]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[2]) );
  XNOR U17 ( .A(B[2]), .B(A[2]), .Z(n17) );
  XOR U18 ( .A(n18), .B(n19), .Z(SUM[1]) );
  XOR U19 ( .A(B[1]), .B(A[1]), .Z(n19) );
  NAND U20 ( .A(n22), .B(B[9]), .Z(n21) );
  NANDN U21 ( .A(A[9]), .B(n2), .Z(n22) );
  NANDN U22 ( .A(n2), .B(A[9]), .Z(n20) );
  AND U23 ( .A(n23), .B(n24), .Z(n2) );
  NAND U24 ( .A(n25), .B(B[8]), .Z(n24) );
  NANDN U25 ( .A(A[8]), .B(n4), .Z(n25) );
  NANDN U26 ( .A(n4), .B(A[8]), .Z(n23) );
  AND U27 ( .A(n26), .B(n27), .Z(n4) );
  NAND U28 ( .A(n28), .B(B[7]), .Z(n27) );
  NANDN U29 ( .A(A[7]), .B(n6), .Z(n28) );
  NANDN U30 ( .A(n6), .B(A[7]), .Z(n26) );
  AND U31 ( .A(n29), .B(n30), .Z(n6) );
  NAND U32 ( .A(n31), .B(B[6]), .Z(n30) );
  NANDN U33 ( .A(A[6]), .B(n8), .Z(n31) );
  NANDN U34 ( .A(n8), .B(A[6]), .Z(n29) );
  AND U35 ( .A(n32), .B(n33), .Z(n8) );
  NAND U36 ( .A(n34), .B(B[5]), .Z(n33) );
  NANDN U37 ( .A(A[5]), .B(n10), .Z(n34) );
  NANDN U38 ( .A(n10), .B(A[5]), .Z(n32) );
  AND U39 ( .A(n35), .B(n36), .Z(n10) );
  NAND U40 ( .A(n37), .B(B[4]), .Z(n36) );
  NANDN U41 ( .A(A[4]), .B(n12), .Z(n37) );
  NANDN U42 ( .A(n12), .B(A[4]), .Z(n35) );
  AND U43 ( .A(n38), .B(n39), .Z(n12) );
  NAND U44 ( .A(n40), .B(B[3]), .Z(n39) );
  NANDN U45 ( .A(A[3]), .B(n14), .Z(n40) );
  NANDN U46 ( .A(n14), .B(A[3]), .Z(n38) );
  AND U47 ( .A(n41), .B(n42), .Z(n14) );
  NAND U48 ( .A(n43), .B(B[2]), .Z(n42) );
  NANDN U49 ( .A(A[2]), .B(n16), .Z(n43) );
  NANDN U50 ( .A(n16), .B(A[2]), .Z(n41) );
  AND U51 ( .A(n44), .B(n45), .Z(n16) );
  NAND U52 ( .A(n46), .B(B[1]), .Z(n45) );
  OR U53 ( .A(n18), .B(A[1]), .Z(n46) );
  NAND U54 ( .A(n18), .B(A[1]), .Z(n44) );
  AND U55 ( .A(B[0]), .B(A[0]), .Z(n18) );
  XOR U56 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_4 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46;

  NAND U1 ( .A(n20), .B(n21), .Z(SUM[10]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[9]) );
  XNOR U3 ( .A(B[9]), .B(A[9]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[8]) );
  XNOR U5 ( .A(B[8]), .B(A[8]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[7]) );
  XNOR U7 ( .A(B[7]), .B(A[7]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[6]) );
  XNOR U9 ( .A(B[6]), .B(A[6]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XNOR U11 ( .A(B[5]), .B(A[5]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[4]) );
  XNOR U13 ( .A(B[4]), .B(A[4]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[3]) );
  XNOR U15 ( .A(B[3]), .B(A[3]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[2]) );
  XNOR U17 ( .A(B[2]), .B(A[2]), .Z(n17) );
  XOR U18 ( .A(n18), .B(n19), .Z(SUM[1]) );
  XOR U19 ( .A(B[1]), .B(A[1]), .Z(n19) );
  NAND U20 ( .A(n22), .B(B[9]), .Z(n21) );
  NANDN U21 ( .A(A[9]), .B(n2), .Z(n22) );
  NANDN U22 ( .A(n2), .B(A[9]), .Z(n20) );
  AND U23 ( .A(n23), .B(n24), .Z(n2) );
  NAND U24 ( .A(n25), .B(B[8]), .Z(n24) );
  NANDN U25 ( .A(A[8]), .B(n4), .Z(n25) );
  NANDN U26 ( .A(n4), .B(A[8]), .Z(n23) );
  AND U27 ( .A(n26), .B(n27), .Z(n4) );
  NAND U28 ( .A(n28), .B(B[7]), .Z(n27) );
  NANDN U29 ( .A(A[7]), .B(n6), .Z(n28) );
  NANDN U30 ( .A(n6), .B(A[7]), .Z(n26) );
  AND U31 ( .A(n29), .B(n30), .Z(n6) );
  NAND U32 ( .A(n31), .B(B[6]), .Z(n30) );
  NANDN U33 ( .A(A[6]), .B(n8), .Z(n31) );
  NANDN U34 ( .A(n8), .B(A[6]), .Z(n29) );
  AND U35 ( .A(n32), .B(n33), .Z(n8) );
  NAND U36 ( .A(n34), .B(B[5]), .Z(n33) );
  NANDN U37 ( .A(A[5]), .B(n10), .Z(n34) );
  NANDN U38 ( .A(n10), .B(A[5]), .Z(n32) );
  AND U39 ( .A(n35), .B(n36), .Z(n10) );
  NAND U40 ( .A(n37), .B(B[4]), .Z(n36) );
  NANDN U41 ( .A(A[4]), .B(n12), .Z(n37) );
  NANDN U42 ( .A(n12), .B(A[4]), .Z(n35) );
  AND U43 ( .A(n38), .B(n39), .Z(n12) );
  NAND U44 ( .A(n40), .B(B[3]), .Z(n39) );
  NANDN U45 ( .A(A[3]), .B(n14), .Z(n40) );
  NANDN U46 ( .A(n14), .B(A[3]), .Z(n38) );
  AND U47 ( .A(n41), .B(n42), .Z(n14) );
  NAND U48 ( .A(n43), .B(B[2]), .Z(n42) );
  NANDN U49 ( .A(A[2]), .B(n16), .Z(n43) );
  NANDN U50 ( .A(n16), .B(A[2]), .Z(n41) );
  AND U51 ( .A(n44), .B(n45), .Z(n16) );
  NAND U52 ( .A(n46), .B(B[1]), .Z(n45) );
  OR U53 ( .A(n18), .B(A[1]), .Z(n46) );
  NAND U54 ( .A(n18), .B(A[1]), .Z(n44) );
  AND U55 ( .A(B[0]), .B(A[0]), .Z(n18) );
  XOR U56 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_5 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44;

  AND U1 ( .A(n2), .B(B[9]), .Z(SUM[10]) );
  IV U2 ( .A(n4), .Z(n2) );
  IV U3 ( .A(B[9]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n3), .Z(SUM[9]) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[8]) );
  XNOR U6 ( .A(B[8]), .B(A[8]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[7]) );
  XNOR U8 ( .A(B[7]), .B(A[7]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[6]) );
  XNOR U10 ( .A(B[6]), .B(A[6]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[5]) );
  XNOR U12 ( .A(B[5]), .B(A[5]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[4]) );
  XNOR U14 ( .A(B[4]), .B(A[4]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[3]) );
  XNOR U16 ( .A(B[3]), .B(A[3]), .Z(n16) );
  XOR U17 ( .A(n17), .B(n18), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n18) );
  XOR U19 ( .A(n19), .B(n20), .Z(SUM[1]) );
  XOR U20 ( .A(B[1]), .B(A[1]), .Z(n20) );
  AND U21 ( .A(n21), .B(n22), .Z(n4) );
  NAND U22 ( .A(n23), .B(B[8]), .Z(n22) );
  NANDN U23 ( .A(A[8]), .B(n5), .Z(n23) );
  NANDN U24 ( .A(n5), .B(A[8]), .Z(n21) );
  AND U25 ( .A(n24), .B(n25), .Z(n5) );
  NAND U26 ( .A(n26), .B(B[7]), .Z(n25) );
  NANDN U27 ( .A(A[7]), .B(n7), .Z(n26) );
  NANDN U28 ( .A(n7), .B(A[7]), .Z(n24) );
  AND U29 ( .A(n27), .B(n28), .Z(n7) );
  NAND U30 ( .A(n29), .B(B[6]), .Z(n28) );
  NANDN U31 ( .A(A[6]), .B(n9), .Z(n29) );
  NANDN U32 ( .A(n9), .B(A[6]), .Z(n27) );
  AND U33 ( .A(n30), .B(n31), .Z(n9) );
  NAND U34 ( .A(n32), .B(B[5]), .Z(n31) );
  NANDN U35 ( .A(A[5]), .B(n11), .Z(n32) );
  NANDN U36 ( .A(n11), .B(A[5]), .Z(n30) );
  AND U37 ( .A(n33), .B(n34), .Z(n11) );
  NAND U38 ( .A(n35), .B(B[4]), .Z(n34) );
  NANDN U39 ( .A(A[4]), .B(n13), .Z(n35) );
  NANDN U40 ( .A(n13), .B(A[4]), .Z(n33) );
  AND U41 ( .A(n36), .B(n37), .Z(n13) );
  NAND U42 ( .A(n38), .B(B[3]), .Z(n37) );
  NANDN U43 ( .A(A[3]), .B(n15), .Z(n38) );
  NANDN U44 ( .A(n15), .B(A[3]), .Z(n36) );
  AND U45 ( .A(n39), .B(n40), .Z(n15) );
  NAND U46 ( .A(n41), .B(B[2]), .Z(n40) );
  NANDN U47 ( .A(A[2]), .B(n17), .Z(n41) );
  NANDN U48 ( .A(n17), .B(A[2]), .Z(n39) );
  AND U49 ( .A(n42), .B(n43), .Z(n17) );
  NAND U50 ( .A(n44), .B(B[1]), .Z(n43) );
  OR U51 ( .A(n19), .B(A[1]), .Z(n44) );
  NAND U52 ( .A(n19), .B(A[1]), .Z(n42) );
  AND U53 ( .A(B[0]), .B(A[0]), .Z(n19) );
  XOR U54 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_6 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41;

  NAND U1 ( .A(n18), .B(n19), .Z(SUM[9]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[8]) );
  XNOR U3 ( .A(B[8]), .B(A[8]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[7]) );
  XNOR U5 ( .A(B[7]), .B(A[7]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[6]) );
  XNOR U7 ( .A(B[6]), .B(A[6]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[5]) );
  XNOR U9 ( .A(B[5]), .B(A[5]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[4]) );
  XNOR U11 ( .A(B[4]), .B(A[4]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[3]) );
  XNOR U13 ( .A(B[3]), .B(A[3]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[2]) );
  XNOR U15 ( .A(B[2]), .B(A[2]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[1]) );
  XOR U17 ( .A(B[1]), .B(A[1]), .Z(n17) );
  NAND U18 ( .A(n20), .B(B[8]), .Z(n19) );
  NANDN U19 ( .A(A[8]), .B(n2), .Z(n20) );
  NANDN U20 ( .A(n2), .B(A[8]), .Z(n18) );
  AND U21 ( .A(n21), .B(n22), .Z(n2) );
  NAND U22 ( .A(n23), .B(B[7]), .Z(n22) );
  NANDN U23 ( .A(A[7]), .B(n4), .Z(n23) );
  NANDN U24 ( .A(n4), .B(A[7]), .Z(n21) );
  AND U25 ( .A(n24), .B(n25), .Z(n4) );
  NAND U26 ( .A(n26), .B(B[6]), .Z(n25) );
  NANDN U27 ( .A(A[6]), .B(n6), .Z(n26) );
  NANDN U28 ( .A(n6), .B(A[6]), .Z(n24) );
  AND U29 ( .A(n27), .B(n28), .Z(n6) );
  NAND U30 ( .A(n29), .B(B[5]), .Z(n28) );
  NANDN U31 ( .A(A[5]), .B(n8), .Z(n29) );
  NANDN U32 ( .A(n8), .B(A[5]), .Z(n27) );
  AND U33 ( .A(n30), .B(n31), .Z(n8) );
  NAND U34 ( .A(n32), .B(B[4]), .Z(n31) );
  NANDN U35 ( .A(A[4]), .B(n10), .Z(n32) );
  NANDN U36 ( .A(n10), .B(A[4]), .Z(n30) );
  AND U37 ( .A(n33), .B(n34), .Z(n10) );
  NAND U38 ( .A(n35), .B(B[3]), .Z(n34) );
  NANDN U39 ( .A(A[3]), .B(n12), .Z(n35) );
  NANDN U40 ( .A(n12), .B(A[3]), .Z(n33) );
  AND U41 ( .A(n36), .B(n37), .Z(n12) );
  NAND U42 ( .A(n38), .B(B[2]), .Z(n37) );
  NANDN U43 ( .A(A[2]), .B(n14), .Z(n38) );
  NANDN U44 ( .A(n14), .B(A[2]), .Z(n36) );
  AND U45 ( .A(n39), .B(n40), .Z(n14) );
  NAND U46 ( .A(n41), .B(B[1]), .Z(n40) );
  OR U47 ( .A(n16), .B(A[1]), .Z(n41) );
  NAND U48 ( .A(n16), .B(A[1]), .Z(n39) );
  AND U49 ( .A(B[0]), .B(A[0]), .Z(n16) );
  XOR U50 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_7 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41;

  NAND U1 ( .A(n18), .B(n19), .Z(SUM[9]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[8]) );
  XNOR U3 ( .A(B[8]), .B(A[8]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[7]) );
  XNOR U5 ( .A(B[7]), .B(A[7]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[6]) );
  XNOR U7 ( .A(B[6]), .B(A[6]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[5]) );
  XNOR U9 ( .A(B[5]), .B(A[5]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[4]) );
  XNOR U11 ( .A(B[4]), .B(A[4]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[3]) );
  XNOR U13 ( .A(B[3]), .B(A[3]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[2]) );
  XNOR U15 ( .A(B[2]), .B(A[2]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[1]) );
  XOR U17 ( .A(B[1]), .B(A[1]), .Z(n17) );
  NAND U18 ( .A(n20), .B(B[8]), .Z(n19) );
  NANDN U19 ( .A(A[8]), .B(n2), .Z(n20) );
  NANDN U20 ( .A(n2), .B(A[8]), .Z(n18) );
  AND U21 ( .A(n21), .B(n22), .Z(n2) );
  NAND U22 ( .A(n23), .B(B[7]), .Z(n22) );
  NANDN U23 ( .A(A[7]), .B(n4), .Z(n23) );
  NANDN U24 ( .A(n4), .B(A[7]), .Z(n21) );
  AND U25 ( .A(n24), .B(n25), .Z(n4) );
  NAND U26 ( .A(n26), .B(B[6]), .Z(n25) );
  NANDN U27 ( .A(A[6]), .B(n6), .Z(n26) );
  NANDN U28 ( .A(n6), .B(A[6]), .Z(n24) );
  AND U29 ( .A(n27), .B(n28), .Z(n6) );
  NAND U30 ( .A(n29), .B(B[5]), .Z(n28) );
  NANDN U31 ( .A(A[5]), .B(n8), .Z(n29) );
  NANDN U32 ( .A(n8), .B(A[5]), .Z(n27) );
  AND U33 ( .A(n30), .B(n31), .Z(n8) );
  NAND U34 ( .A(n32), .B(B[4]), .Z(n31) );
  NANDN U35 ( .A(A[4]), .B(n10), .Z(n32) );
  NANDN U36 ( .A(n10), .B(A[4]), .Z(n30) );
  AND U37 ( .A(n33), .B(n34), .Z(n10) );
  NAND U38 ( .A(n35), .B(B[3]), .Z(n34) );
  NANDN U39 ( .A(A[3]), .B(n12), .Z(n35) );
  NANDN U40 ( .A(n12), .B(A[3]), .Z(n33) );
  AND U41 ( .A(n36), .B(n37), .Z(n12) );
  NAND U42 ( .A(n38), .B(B[2]), .Z(n37) );
  NANDN U43 ( .A(A[2]), .B(n14), .Z(n38) );
  NANDN U44 ( .A(n14), .B(A[2]), .Z(n36) );
  AND U45 ( .A(n39), .B(n40), .Z(n14) );
  NAND U46 ( .A(n41), .B(B[1]), .Z(n40) );
  OR U47 ( .A(n16), .B(A[1]), .Z(n41) );
  NAND U48 ( .A(n16), .B(A[1]), .Z(n39) );
  AND U49 ( .A(B[0]), .B(A[0]), .Z(n16) );
  XOR U50 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_8 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41;

  NAND U1 ( .A(n18), .B(n19), .Z(SUM[9]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[8]) );
  XNOR U3 ( .A(B[8]), .B(A[8]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[7]) );
  XNOR U5 ( .A(B[7]), .B(A[7]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[6]) );
  XNOR U7 ( .A(B[6]), .B(A[6]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[5]) );
  XNOR U9 ( .A(B[5]), .B(A[5]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[4]) );
  XNOR U11 ( .A(B[4]), .B(A[4]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[3]) );
  XNOR U13 ( .A(B[3]), .B(A[3]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[2]) );
  XNOR U15 ( .A(B[2]), .B(A[2]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[1]) );
  XOR U17 ( .A(B[1]), .B(A[1]), .Z(n17) );
  NAND U18 ( .A(n20), .B(B[8]), .Z(n19) );
  NANDN U19 ( .A(A[8]), .B(n2), .Z(n20) );
  NANDN U20 ( .A(n2), .B(A[8]), .Z(n18) );
  AND U21 ( .A(n21), .B(n22), .Z(n2) );
  NAND U22 ( .A(n23), .B(B[7]), .Z(n22) );
  NANDN U23 ( .A(A[7]), .B(n4), .Z(n23) );
  NANDN U24 ( .A(n4), .B(A[7]), .Z(n21) );
  AND U25 ( .A(n24), .B(n25), .Z(n4) );
  NAND U26 ( .A(n26), .B(B[6]), .Z(n25) );
  NANDN U27 ( .A(A[6]), .B(n6), .Z(n26) );
  NANDN U28 ( .A(n6), .B(A[6]), .Z(n24) );
  AND U29 ( .A(n27), .B(n28), .Z(n6) );
  NAND U30 ( .A(n29), .B(B[5]), .Z(n28) );
  NANDN U31 ( .A(A[5]), .B(n8), .Z(n29) );
  NANDN U32 ( .A(n8), .B(A[5]), .Z(n27) );
  AND U33 ( .A(n30), .B(n31), .Z(n8) );
  NAND U34 ( .A(n32), .B(B[4]), .Z(n31) );
  NANDN U35 ( .A(A[4]), .B(n10), .Z(n32) );
  NANDN U36 ( .A(n10), .B(A[4]), .Z(n30) );
  AND U37 ( .A(n33), .B(n34), .Z(n10) );
  NAND U38 ( .A(n35), .B(B[3]), .Z(n34) );
  NANDN U39 ( .A(A[3]), .B(n12), .Z(n35) );
  NANDN U40 ( .A(n12), .B(A[3]), .Z(n33) );
  AND U41 ( .A(n36), .B(n37), .Z(n12) );
  NAND U42 ( .A(n38), .B(B[2]), .Z(n37) );
  NANDN U43 ( .A(A[2]), .B(n14), .Z(n38) );
  NANDN U44 ( .A(n14), .B(A[2]), .Z(n36) );
  AND U45 ( .A(n39), .B(n40), .Z(n14) );
  NAND U46 ( .A(n41), .B(B[1]), .Z(n40) );
  OR U47 ( .A(n16), .B(A[1]), .Z(n41) );
  NAND U48 ( .A(n16), .B(A[1]), .Z(n39) );
  AND U49 ( .A(B[0]), .B(A[0]), .Z(n16) );
  XOR U50 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_9 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41;

  NAND U1 ( .A(n18), .B(n19), .Z(SUM[9]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[8]) );
  XNOR U3 ( .A(B[8]), .B(A[8]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[7]) );
  XNOR U5 ( .A(B[7]), .B(A[7]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[6]) );
  XNOR U7 ( .A(B[6]), .B(A[6]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[5]) );
  XNOR U9 ( .A(B[5]), .B(A[5]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[4]) );
  XNOR U11 ( .A(B[4]), .B(A[4]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[3]) );
  XNOR U13 ( .A(B[3]), .B(A[3]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[2]) );
  XNOR U15 ( .A(B[2]), .B(A[2]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[1]) );
  XOR U17 ( .A(B[1]), .B(A[1]), .Z(n17) );
  NAND U18 ( .A(n20), .B(B[8]), .Z(n19) );
  NANDN U19 ( .A(A[8]), .B(n2), .Z(n20) );
  NANDN U20 ( .A(n2), .B(A[8]), .Z(n18) );
  AND U21 ( .A(n21), .B(n22), .Z(n2) );
  NAND U22 ( .A(n23), .B(B[7]), .Z(n22) );
  NANDN U23 ( .A(A[7]), .B(n4), .Z(n23) );
  NANDN U24 ( .A(n4), .B(A[7]), .Z(n21) );
  AND U25 ( .A(n24), .B(n25), .Z(n4) );
  NAND U26 ( .A(n26), .B(B[6]), .Z(n25) );
  NANDN U27 ( .A(A[6]), .B(n6), .Z(n26) );
  NANDN U28 ( .A(n6), .B(A[6]), .Z(n24) );
  AND U29 ( .A(n27), .B(n28), .Z(n6) );
  NAND U30 ( .A(n29), .B(B[5]), .Z(n28) );
  NANDN U31 ( .A(A[5]), .B(n8), .Z(n29) );
  NANDN U32 ( .A(n8), .B(A[5]), .Z(n27) );
  AND U33 ( .A(n30), .B(n31), .Z(n8) );
  NAND U34 ( .A(n32), .B(B[4]), .Z(n31) );
  NANDN U35 ( .A(A[4]), .B(n10), .Z(n32) );
  NANDN U36 ( .A(n10), .B(A[4]), .Z(n30) );
  AND U37 ( .A(n33), .B(n34), .Z(n10) );
  NAND U38 ( .A(n35), .B(B[3]), .Z(n34) );
  NANDN U39 ( .A(A[3]), .B(n12), .Z(n35) );
  NANDN U40 ( .A(n12), .B(A[3]), .Z(n33) );
  AND U41 ( .A(n36), .B(n37), .Z(n12) );
  NAND U42 ( .A(n38), .B(B[2]), .Z(n37) );
  NANDN U43 ( .A(A[2]), .B(n14), .Z(n38) );
  NANDN U44 ( .A(n14), .B(A[2]), .Z(n36) );
  AND U45 ( .A(n39), .B(n40), .Z(n14) );
  NAND U46 ( .A(n41), .B(B[1]), .Z(n40) );
  OR U47 ( .A(n16), .B(A[1]), .Z(n41) );
  NAND U48 ( .A(n16), .B(A[1]), .Z(n39) );
  AND U49 ( .A(B[0]), .B(A[0]), .Z(n16) );
  XOR U50 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_10 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39;

  AND U1 ( .A(n2), .B(B[8]), .Z(SUM[9]) );
  IV U2 ( .A(n4), .Z(n2) );
  IV U3 ( .A(B[8]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n3), .Z(SUM[8]) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[7]) );
  XNOR U6 ( .A(B[7]), .B(A[7]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[6]) );
  XNOR U8 ( .A(B[6]), .B(A[6]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[5]) );
  XNOR U10 ( .A(B[5]), .B(A[5]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[3]) );
  XNOR U14 ( .A(B[3]), .B(A[3]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U16 ( .A(B[2]), .B(A[2]), .Z(n16) );
  XOR U17 ( .A(n17), .B(n18), .Z(SUM[1]) );
  XOR U18 ( .A(B[1]), .B(A[1]), .Z(n18) );
  AND U19 ( .A(n19), .B(n20), .Z(n4) );
  NAND U20 ( .A(n21), .B(B[7]), .Z(n20) );
  NANDN U21 ( .A(A[7]), .B(n5), .Z(n21) );
  NANDN U22 ( .A(n5), .B(A[7]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n5) );
  NAND U24 ( .A(n24), .B(B[6]), .Z(n23) );
  NANDN U25 ( .A(A[6]), .B(n7), .Z(n24) );
  NANDN U26 ( .A(n7), .B(A[6]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n7) );
  NAND U28 ( .A(n27), .B(B[5]), .Z(n26) );
  NANDN U29 ( .A(A[5]), .B(n9), .Z(n27) );
  NANDN U30 ( .A(n9), .B(A[5]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n9) );
  NAND U32 ( .A(n30), .B(B[4]), .Z(n29) );
  NANDN U33 ( .A(A[4]), .B(n11), .Z(n30) );
  NANDN U34 ( .A(n11), .B(A[4]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n11) );
  NAND U36 ( .A(n33), .B(B[3]), .Z(n32) );
  NANDN U37 ( .A(A[3]), .B(n13), .Z(n33) );
  NANDN U38 ( .A(n13), .B(A[3]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n13) );
  NAND U40 ( .A(n36), .B(B[2]), .Z(n35) );
  NANDN U41 ( .A(A[2]), .B(n15), .Z(n36) );
  NANDN U42 ( .A(n15), .B(A[2]), .Z(n34) );
  AND U43 ( .A(n37), .B(n38), .Z(n15) );
  NAND U44 ( .A(n39), .B(B[1]), .Z(n38) );
  OR U45 ( .A(n17), .B(A[1]), .Z(n39) );
  NAND U46 ( .A(n17), .B(A[1]), .Z(n37) );
  AND U47 ( .A(B[0]), .B(A[0]), .Z(n17) );
  XOR U48 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_11 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_12 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_13 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_14 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_15 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_16 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_17 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_18 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_19 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_20 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_21 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_22 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_23 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_24 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_25 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_26 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_27 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_28 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_29 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_30 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_31 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_32 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_33 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_34 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_35 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_36 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_37 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_38 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_39 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_40 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_41 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_42 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_43 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_44 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_45 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_46 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_47 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_48 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_49 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_50 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_51 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_52 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_53 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_54 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_55 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_56 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_57 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_58 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_59 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_60 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_61 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_62 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_63 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_64 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_65 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_66 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_67 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_68 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_69 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_70 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_71 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_72 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_73 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_74 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_75 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_76 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_77 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_78 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_79 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_80 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_81 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_82 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_83 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24;

  AND U1 ( .A(n2), .B(B[5]), .Z(SUM[6]) );
  IV U2 ( .A(n4), .Z(n2) );
  IV U3 ( .A(B[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n3), .Z(SUM[5]) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[3]) );
  XNOR U8 ( .A(B[3]), .B(A[3]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[2]) );
  XNOR U10 ( .A(B[2]), .B(A[2]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[1]) );
  XOR U12 ( .A(B[1]), .B(A[1]), .Z(n12) );
  AND U13 ( .A(n13), .B(n14), .Z(n4) );
  NAND U14 ( .A(n15), .B(B[4]), .Z(n14) );
  NANDN U15 ( .A(A[4]), .B(n5), .Z(n15) );
  NANDN U16 ( .A(n5), .B(A[4]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n5) );
  NAND U18 ( .A(n18), .B(B[3]), .Z(n17) );
  NANDN U19 ( .A(A[3]), .B(n7), .Z(n18) );
  NANDN U20 ( .A(n7), .B(A[3]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n7) );
  NAND U22 ( .A(n21), .B(B[2]), .Z(n20) );
  NANDN U23 ( .A(A[2]), .B(n9), .Z(n21) );
  NANDN U24 ( .A(n9), .B(A[2]), .Z(n19) );
  AND U25 ( .A(n22), .B(n23), .Z(n9) );
  NAND U26 ( .A(n24), .B(B[1]), .Z(n23) );
  OR U27 ( .A(n11), .B(A[1]), .Z(n24) );
  NAND U28 ( .A(n11), .B(A[1]), .Z(n22) );
  AND U29 ( .A(B[0]), .B(A[0]), .Z(n11) );
  XOR U30 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_84 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_85 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_86 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_87 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_88 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_89 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_90 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_91 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_92 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_93 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_94 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_95 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_96 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_97 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_98 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_99 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_100 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_101 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_102 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_103 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_104 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_105 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_106 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_107 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_108 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_109 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_110 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_111 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_112 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_113 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_114 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_115 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_116 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_117 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_118 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_119 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_120 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_121 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_122 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_123 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_124 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_125 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_126 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_127 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_128 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_129 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_130 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_131 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_132 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_133 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_134 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_135 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_136 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_137 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_138 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_139 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_140 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_141 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_142 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_143 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_144 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_145 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_146 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_147 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_148 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_149 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_150 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_151 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_152 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_153 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_154 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_155 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_156 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_157 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_158 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_159 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_160 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_161 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_162 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_163 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_164 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_165 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_166 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4 ( clk, rst, x, y, o );
  input [3999:0] x;
  input [3999:0] y;
  output [13:0] o;
  input clk, rst;
  wire   N27929, N27930, N27931, N27932, N27933, N27941, N27942, N27943,
         N27944, N27945, N27953, N27954, N27955, N27956, N27957, N27965,
         N27966, N27967, N27968, N27969, N27977, N27978, N27979, N27980,
         N27981, N27989, N27990, N27991, N27992, N27993, N28001, N28002,
         N28003, N28004, N28005, N28013, N28014, N28015, N28016, N28017,
         N28025, N28026, N28027, N28028, N28029, N28037, N28038, N28039,
         N28040, N28041, N28049, N28050, N28051, N28052, N28053, N28061,
         N28062, N28063, N28064, N28065, N28073, N28074, N28075, N28076,
         N28077, N28085, N28086, N28087, N28088, N28089, N28097, N28098,
         N28099, N28100, N28101, N28109, N28110, N28111, N28112, N28113,
         N28121, N28122, N28123, N28124, N28125, N28133, N28134, N28135,
         N28136, N28137, N28145, N28146, N28147, N28148, N28149, N28157,
         N28158, N28159, N28160, N28161, N28169, N28170, N28171, N28172,
         N28173, N28181, N28182, N28183, N28184, N28185, N28193, N28194,
         N28195, N28196, N28197, N28205, N28206, N28207, N28208, N28209,
         N28217, N28218, N28219, N28220, N28221, N28229, N28230, N28231,
         N28232, N28233, N28241, N28242, N28243, N28244, N28245, N28253,
         N28254, N28255, N28256, N28257, N28265, N28266, N28267, N28268,
         N28269, N28277, N28278, N28279, N28280, N28281, N28289, N28290,
         N28291, N28292, N28293, N28301, N28302, N28303, N28304, N28305,
         N28313, N28314, N28315, N28316, N28317, N28325, N28326, N28327,
         N28328, N28329, N28337, N28338, N28339, N28340, N28341, N28349,
         N28350, N28351, N28352, N28353, N28361, N28362, N28363, N28364,
         N28365, N28373, N28374, N28375, N28376, N28377, N28385, N28386,
         N28387, N28388, N28389, N28397, N28398, N28399, N28400, N28401,
         N28409, N28410, N28411, N28412, N28413, N28421, N28422, N28423,
         N28424, N28425, N28433, N28434, N28435, N28436, N28437, N28445,
         N28446, N28447, N28448, N28449, N28457, N28458, N28459, N28460,
         N28461, N28469, N28470, N28471, N28472, N28473, N28481, N28482,
         N28483, N28484, N28485, N28493, N28494, N28495, N28496, N28497,
         N28505, N28506, N28507, N28508, N28509, N28517, N28518, N28519,
         N28520, N28521, N28529, N28530, N28531, N28532, N28533, N28541,
         N28542, N28543, N28544, N28545, N28553, N28554, N28555, N28556,
         N28557, N28565, N28566, N28567, N28568, N28569, N28577, N28578,
         N28579, N28580, N28581, N28589, N28590, N28591, N28592, N28593,
         N28601, N28602, N28603, N28604, N28605, N28613, N28614, N28615,
         N28616, N28617, N28625, N28626, N28627, N28628, N28629, N28637,
         N28638, N28639, N28640, N28641, N28649, N28650, N28651, N28652,
         N28653, N28661, N28662, N28663, N28664, N28665, N28673, N28674,
         N28675, N28676, N28677, N28685, N28686, N28687, N28688, N28689,
         N28697, N28698, N28699, N28700, N28701, N28709, N28710, N28711,
         N28712, N28713, N28721, N28722, N28723, N28724, N28725, N28733,
         N28734, N28735, N28736, N28737, N28745, N28746, N28747, N28748,
         N28749, N28757, N28758, N28759, N28760, N28761, N28769, N28770,
         N28771, N28772, N28773, N28781, N28782, N28783, N28784, N28785,
         N28793, N28794, N28795, N28796, N28797, N28805, N28806, N28807,
         N28808, N28809, N28817, N28818, N28819, N28820, N28821, N28829,
         N28830, N28831, N28832, N28833, N28841, N28842, N28843, N28844,
         N28845, N28853, N28854, N28855, N28856, N28857, N28865, N28866,
         N28867, N28868, N28869, N28877, N28878, N28879, N28880, N28881,
         N28889, N28890, N28891, N28892, N28893, N28901, N28902, N28903,
         N28904, N28905, N28913, N28914, N28915, N28916, N28917, N28925,
         N28926, N28927, N28928, N28929, N28937, N28938, N28939, N28940,
         N28941, N28949, N28950, N28951, N28952, N28953, N28961, N28962,
         N28963, N28964, N28965, N28973, N28974, N28975, N28976, N28977,
         N28985, N28986, N28987, N28988, N28989, N28997, N28998, N28999,
         N29000, N29001, N29009, N29010, N29011, N29012, N29013, N29021,
         N29022, N29023, N29024, N29025, N29033, N29034, N29035, N29036,
         N29037, N29045, N29046, N29047, N29048, N29049, N29057, N29058,
         N29059, N29060, N29061, N29069, N29070, N29071, N29072, N29073,
         N29081, N29082, N29083, N29084, N29085, N29093, N29094, N29095,
         N29096, N29097, N29105, N29106, N29107, N29108, N29109, N29117,
         N29118, N29119, N29120, N29121, N29129, N29130, N29131, N29132,
         N29133, N29141, N29142, N29143, N29144, N29145, N29153, N29154,
         N29155, N29156, N29157, N29165, N29166, N29167, N29168, N29169,
         N29177, N29178, N29179, N29180, N29181, N29189, N29190, N29191,
         N29192, N29193, N29201, N29202, N29203, N29204, N29205, N29213,
         N29214, N29215, N29216, N29217, N29225, N29226, N29227, N29228,
         N29229, N29237, N29238, N29239, N29240, N29241, N29249, N29250,
         N29251, N29252, N29253, N29261, N29262, N29263, N29264, N29265,
         N29273, N29274, N29275, N29276, N29277, N29285, N29286, N29287,
         N29288, N29289, N29297, N29298, N29299, N29300, N29301, N29309,
         N29310, N29311, N29312, N29313, N29321, N29322, N29323, N29324,
         N29325, N29333, N29334, N29335, N29336, N29337, N29345, N29346,
         N29347, N29348, N29349, N29357, N29358, N29359, N29360, N29361,
         N29369, N29370, N29371, N29372, N29373, N29381, N29382, N29383,
         N29384, N29385, N29393, N29394, N29395, N29396, N29397, N29405,
         N29406, N29407, N29408, N29409, N29417, N29418, N29419, N29420,
         N29421, N29429, N29430, N29431, N29432, N29433, N29441, N29442,
         N29443, N29444, N29445, N29453, N29454, N29455, N29456, N29457,
         N29465, N29466, N29467, N29468, N29469, N29477, N29478, N29479,
         N29480, N29481, N29489, N29490, N29491, N29492, N29493, N29501,
         N29502, N29503, N29504, N29505, N29513, N29514, N29515, N29516,
         N29517, N29525, N29526, N29527, N29528, N29529, N29537, N29538,
         N29539, N29540, N29541, N29549, N29550, N29551, N29552, N29553,
         N29561, N29562, N29563, N29564, N29565, N29573, N29574, N29575,
         N29576, N29577, N29585, N29586, N29587, N29588, N29589, N29597,
         N29598, N29599, N29600, N29601, N29609, N29610, N29611, N29612,
         N29613, N29621, N29622, N29623, N29624, N29625, N29633, N29634,
         N29635, N29636, N29637, N29645, N29646, N29647, N29648, N29649,
         N29657, N29658, N29659, N29660, N29661, N29669, N29670, N29671,
         N29672, N29673, N29681, N29682, N29683, N29684, N29685, N29693,
         N29694, N29695, N29696, N29697, N29705, N29706, N29707, N29708,
         N29709, N29717, N29718, N29719, N29720, N29721, N29729, N29730,
         N29731, N29732, N29733, N29741, N29742, N29743, N29744, N29745,
         N29753, N29754, N29755, N29756, N29757, N29765, N29766, N29767,
         N29768, N29769, N29777, N29778, N29779, N29780, N29781, N29789,
         N29790, N29791, N29792, N29793, N29801, N29802, N29803, N29804,
         N29805, N29813, N29814, N29815, N29816, N29817, N29825, N29826,
         N29827, N29828, N29829, N29837, N29838, N29839, N29840, N29841,
         N29849, N29850, N29851, N29852, N29853, N29861, N29862, N29863,
         N29864, N29865, N29873, N29874, N29875, N29876, N29877, N29885,
         N29886, N29887, N29888, N29889, N29897, N29898, N29899, N29900,
         N29901, N29909, N29910, N29911, N29912, N29913, N29921, N29922,
         N29923, N29924, N29925, N29933, N29934, N29935, N29936, N29937,
         N29938, N29945, N29946, N29947, N29948, N29949, N29950, N29957,
         N29958, N29959, N29960, N29961, N29962, N29969, N29970, N29971,
         N29972, N29973, N29974, N29981, N29982, N29983, N29984, N29985,
         N29986, N29993, N29994, N29995, N29996, N29997, N29998, N30005,
         N30006, N30007, N30008, N30009, N30010, N30017, N30018, N30019,
         N30020, N30021, N30022, N30029, N30030, N30031, N30032, N30033,
         N30034, N30041, N30042, N30043, N30044, N30045, N30046, N30053,
         N30054, N30055, N30056, N30057, N30058, N30065, N30066, N30067,
         N30068, N30069, N30070, N30077, N30078, N30079, N30080, N30081,
         N30082, N30089, N30090, N30091, N30092, N30093, N30094, N30101,
         N30102, N30103, N30104, N30105, N30106, N30113, N30114, N30115,
         N30116, N30117, N30118, N30125, N30126, N30127, N30128, N30129,
         N30130, N30137, N30138, N30139, N30140, N30141, N30142, N30149,
         N30150, N30151, N30152, N30153, N30154, N30161, N30162, N30163,
         N30164, N30165, N30166, N30173, N30174, N30175, N30176, N30177,
         N30178, N30185, N30186, N30187, N30188, N30189, N30190, N30197,
         N30198, N30199, N30200, N30201, N30202, N30209, N30210, N30211,
         N30212, N30213, N30214, N30221, N30222, N30223, N30224, N30225,
         N30226, N30233, N30234, N30235, N30236, N30237, N30238, N30245,
         N30246, N30247, N30248, N30249, N30250, N30257, N30258, N30259,
         N30260, N30261, N30262, N30269, N30270, N30271, N30272, N30273,
         N30274, N30281, N30282, N30283, N30284, N30285, N30286, N30293,
         N30294, N30295, N30296, N30297, N30298, N30305, N30306, N30307,
         N30308, N30309, N30310, N30317, N30318, N30319, N30320, N30321,
         N30322, N30329, N30330, N30331, N30332, N30333, N30334, N30341,
         N30342, N30343, N30344, N30345, N30346, N30353, N30354, N30355,
         N30356, N30357, N30358, N30365, N30366, N30367, N30368, N30369,
         N30370, N30377, N30378, N30379, N30380, N30381, N30382, N30389,
         N30390, N30391, N30392, N30393, N30394, N30401, N30402, N30403,
         N30404, N30405, N30406, N30413, N30414, N30415, N30416, N30417,
         N30418, N30425, N30426, N30427, N30428, N30429, N30430, N30437,
         N30438, N30439, N30440, N30441, N30442, N30449, N30450, N30451,
         N30452, N30453, N30454, N30461, N30462, N30463, N30464, N30465,
         N30466, N30473, N30474, N30475, N30476, N30477, N30478, N30485,
         N30486, N30487, N30488, N30489, N30490, N30497, N30498, N30499,
         N30500, N30501, N30502, N30509, N30510, N30511, N30512, N30513,
         N30514, N30521, N30522, N30523, N30524, N30525, N30526, N30533,
         N30534, N30535, N30536, N30537, N30538, N30545, N30546, N30547,
         N30548, N30549, N30550, N30557, N30558, N30559, N30560, N30561,
         N30562, N30569, N30570, N30571, N30572, N30573, N30574, N30581,
         N30582, N30583, N30584, N30585, N30586, N30593, N30594, N30595,
         N30596, N30597, N30598, N30605, N30606, N30607, N30608, N30609,
         N30610, N30617, N30618, N30619, N30620, N30621, N30622, N30629,
         N30630, N30631, N30632, N30633, N30634, N30641, N30642, N30643,
         N30644, N30645, N30646, N30653, N30654, N30655, N30656, N30657,
         N30658, N30665, N30666, N30667, N30668, N30669, N30670, N30677,
         N30678, N30679, N30680, N30681, N30682, N30689, N30690, N30691,
         N30692, N30693, N30694, N30701, N30702, N30703, N30704, N30705,
         N30706, N30713, N30714, N30715, N30716, N30717, N30718, N30725,
         N30726, N30727, N30728, N30729, N30730, N30737, N30738, N30739,
         N30740, N30741, N30742, N30749, N30750, N30751, N30752, N30753,
         N30754, N30761, N30762, N30763, N30764, N30765, N30766, N30773,
         N30774, N30775, N30776, N30777, N30778, N30785, N30786, N30787,
         N30788, N30789, N30790, N30797, N30798, N30799, N30800, N30801,
         N30802, N30809, N30810, N30811, N30812, N30813, N30814, N30821,
         N30822, N30823, N30824, N30825, N30826, N30833, N30834, N30835,
         N30836, N30837, N30838, N30845, N30846, N30847, N30848, N30849,
         N30850, N30857, N30858, N30859, N30860, N30861, N30862, N30869,
         N30870, N30871, N30872, N30873, N30874, N30881, N30882, N30883,
         N30884, N30885, N30886, N30893, N30894, N30895, N30896, N30897,
         N30898, N30905, N30906, N30907, N30908, N30909, N30910, N30917,
         N30918, N30919, N30920, N30921, N30922, N30929, N30930, N30931,
         N30932, N30933, N30934, N30935, N30941, N30942, N30943, N30944,
         N30945, N30946, N30947, N30953, N30954, N30955, N30956, N30957,
         N30958, N30959, N30965, N30966, N30967, N30968, N30969, N30970,
         N30971, N30977, N30978, N30979, N30980, N30981, N30982, N30983,
         N30989, N30990, N30991, N30992, N30993, N30994, N30995, N31001,
         N31002, N31003, N31004, N31005, N31006, N31007, N31013, N31014,
         N31015, N31016, N31017, N31018, N31019, N31025, N31026, N31027,
         N31028, N31029, N31030, N31031, N31037, N31038, N31039, N31040,
         N31041, N31042, N31043, N31049, N31050, N31051, N31052, N31053,
         N31054, N31055, N31061, N31062, N31063, N31064, N31065, N31066,
         N31067, N31073, N31074, N31075, N31076, N31077, N31078, N31079,
         N31085, N31086, N31087, N31088, N31089, N31090, N31091, N31097,
         N31098, N31099, N31100, N31101, N31102, N31103, N31109, N31110,
         N31111, N31112, N31113, N31114, N31115, N31121, N31122, N31123,
         N31124, N31125, N31126, N31127, N31133, N31134, N31135, N31136,
         N31137, N31138, N31139, N31145, N31146, N31147, N31148, N31149,
         N31150, N31151, N31157, N31158, N31159, N31160, N31161, N31162,
         N31163, N31169, N31170, N31171, N31172, N31173, N31174, N31175,
         N31181, N31182, N31183, N31184, N31185, N31186, N31187, N31193,
         N31194, N31195, N31196, N31197, N31198, N31199, N31205, N31206,
         N31207, N31208, N31209, N31210, N31211, N31217, N31218, N31219,
         N31220, N31221, N31222, N31223, N31229, N31230, N31231, N31232,
         N31233, N31234, N31235, N31241, N31242, N31243, N31244, N31245,
         N31246, N31247, N31253, N31254, N31255, N31256, N31257, N31258,
         N31259, N31265, N31266, N31267, N31268, N31269, N31270, N31271,
         N31277, N31278, N31279, N31280, N31281, N31282, N31283, N31289,
         N31290, N31291, N31292, N31293, N31294, N31295, N31301, N31302,
         N31303, N31304, N31305, N31306, N31307, N31313, N31314, N31315,
         N31316, N31317, N31318, N31319, N31325, N31326, N31327, N31328,
         N31329, N31330, N31331, N31337, N31338, N31339, N31340, N31341,
         N31342, N31343, N31349, N31350, N31351, N31352, N31353, N31354,
         N31355, N31361, N31362, N31363, N31364, N31365, N31366, N31367,
         N31373, N31374, N31375, N31376, N31377, N31378, N31379, N31385,
         N31386, N31387, N31388, N31389, N31390, N31391, N31397, N31398,
         N31399, N31400, N31401, N31402, N31403, N31409, N31410, N31411,
         N31412, N31413, N31414, N31415, N31421, N31422, N31423, N31424,
         N31425, N31426, N31427, N31433, N31434, N31435, N31436, N31437,
         N31438, N31439, N31440, N31445, N31446, N31447, N31448, N31449,
         N31450, N31451, N31452, N31457, N31458, N31459, N31460, N31461,
         N31462, N31463, N31464, N31469, N31470, N31471, N31472, N31473,
         N31474, N31475, N31476, N31481, N31482, N31483, N31484, N31485,
         N31486, N31487, N31488, N31493, N31494, N31495, N31496, N31497,
         N31498, N31499, N31500, N31505, N31506, N31507, N31508, N31509,
         N31510, N31511, N31512, N31517, N31518, N31519, N31520, N31521,
         N31522, N31523, N31524, N31529, N31530, N31531, N31532, N31533,
         N31534, N31535, N31536, N31541, N31542, N31543, N31544, N31545,
         N31546, N31547, N31548, N31553, N31554, N31555, N31556, N31557,
         N31558, N31559, N31560, N31565, N31566, N31567, N31568, N31569,
         N31570, N31571, N31572, N31577, N31578, N31579, N31580, N31581,
         N31582, N31583, N31584, N31589, N31590, N31591, N31592, N31593,
         N31594, N31595, N31596, N31601, N31602, N31603, N31604, N31605,
         N31606, N31607, N31608, N31613, N31614, N31615, N31616, N31617,
         N31618, N31619, N31620, N31625, N31626, N31627, N31628, N31629,
         N31630, N31631, N31632, N31637, N31638, N31639, N31640, N31641,
         N31642, N31643, N31644, N31649, N31650, N31651, N31652, N31653,
         N31654, N31655, N31656, N31661, N31662, N31663, N31664, N31665,
         N31666, N31667, N31668, N31673, N31674, N31675, N31676, N31677,
         N31678, N31679, N31680, N31685, N31686, N31687, N31688, N31689,
         N31690, N31691, N31692, N31693, N31697, N31698, N31699, N31700,
         N31701, N31702, N31703, N31704, N31705, N31709, N31710, N31711,
         N31712, N31713, N31714, N31715, N31716, N31717, N31721, N31722,
         N31723, N31724, N31725, N31726, N31727, N31728, N31729, N31733,
         N31734, N31735, N31736, N31737, N31738, N31739, N31740, N31741,
         N31745, N31746, N31747, N31748, N31749, N31750, N31751, N31752,
         N31753, N31757, N31758, N31759, N31760, N31761, N31762, N31763,
         N31764, N31765, N31769, N31770, N31771, N31772, N31773, N31774,
         N31775, N31776, N31777, N31781, N31782, N31783, N31784, N31785,
         N31786, N31787, N31788, N31789, N31793, N31794, N31795, N31796,
         N31797, N31798, N31799, N31800, N31801, N31805, N31806, N31807,
         N31808, N31809, N31810, N31811, N31812, N31813, N31814, N31817,
         N31818, N31819, N31820, N31821, N31822, N31823, N31824, N31825,
         N31826, N31829, N31830, N31831, N31832, N31833, N31834, N31835,
         N31836, N31837, N31838, N31841, N31842, N31843, N31844, N31845,
         N31846, N31847, N31848, N31849, N31850, N31853, N31854, N31855,
         N31856, N31857, N31858, N31859, N31860, N31861, N31862, N31865,
         N31866, N31867, N31868, N31869, N31870, N31871, N31872, N31873,
         N31874, N31875, N31877, N31878, N31879, N31880, N31881, N31882,
         N31883, N31884, N31885, N31886, N31887, N31889, N31890, N31891,
         N31892, N31893, N31894, N31895, N31896, N31897, N31898, N31899,
         N31901, N31902, N31903, N31904, N31905, N31906, N31907, N31908,
         N31909, N31910, N31911, N31912, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,
         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,
         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,
         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
         n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,
         n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
         n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
         n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
         n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,
         n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
         n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,
         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
         n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,
         n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,
         n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,
         n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
         n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
         n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
         n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,
         n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,
         n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
         n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
         n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,
         n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
         n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
         n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,
         n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
         n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432,
         n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440,
         n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,
         n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
         n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
         n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
         n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,
         n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,
         n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
         n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504,
         n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,
         n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,
         n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528,
         n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536,
         n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544,
         n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,
         n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,
         n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568,
         n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576,
         n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,
         n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,
         n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600,
         n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608,
         n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616,
         n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624,
         n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632,
         n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640,
         n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648,
         n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656,
         n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664,
         n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672,
         n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680,
         n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688,
         n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,
         n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704,
         n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,
         n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720,
         n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,
         n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
         n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
         n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
         n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,
         n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
         n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,
         n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,
         n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,
         n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,
         n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,
         n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
         n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,
         n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,
         n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
         n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,
         n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
         n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,
         n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,
         n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,
         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
         n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,
         n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
         n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
         n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,
         n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
         n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,
         n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,
         n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,
         n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
         n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968,
         n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,
         n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
         n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992,
         n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
         n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
         n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016,
         n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024,
         n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,
         n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040,
         n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048,
         n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056,
         n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064,
         n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072,
         n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080,
         n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088,
         n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096,
         n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104,
         n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112,
         n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120,
         n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128,
         n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136,
         n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144,
         n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152,
         n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160,
         n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168,
         n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176,
         n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184,
         n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192,
         n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200,
         n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208,
         n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216,
         n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224,
         n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232,
         n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240,
         n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248,
         n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256,
         n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264,
         n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272,
         n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280,
         n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288,
         n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296,
         n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304,
         n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312,
         n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320,
         n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328,
         n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336,
         n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344,
         n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352,
         n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360,
         n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368,
         n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376,
         n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384,
         n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392,
         n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400,
         n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408,
         n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416,
         n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424,
         n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432,
         n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440,
         n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448,
         n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456,
         n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464,
         n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472,
         n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480,
         n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488,
         n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496,
         n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504,
         n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512,
         n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520,
         n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528,
         n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536,
         n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544,
         n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552,
         n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560,
         n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568,
         n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576,
         n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584,
         n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592,
         n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600,
         n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608,
         n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616,
         n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624,
         n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632,
         n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640,
         n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648,
         n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656,
         n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664,
         n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672,
         n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680,
         n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688,
         n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696,
         n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704,
         n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712,
         n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720,
         n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728,
         n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736,
         n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744,
         n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752,
         n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760,
         n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768,
         n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776,
         n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784,
         n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792,
         n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800,
         n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808,
         n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816,
         n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824,
         n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832,
         n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840,
         n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848,
         n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856,
         n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864,
         n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872,
         n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880,
         n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888,
         n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896,
         n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904,
         n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912,
         n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920,
         n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928,
         n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936,
         n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944,
         n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952,
         n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960,
         n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968,
         n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976,
         n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984,
         n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992,
         n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000,
         n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008,
         n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016,
         n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024,
         n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032,
         n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040,
         n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048,
         n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056,
         n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064,
         n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072,
         n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080,
         n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088,
         n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096,
         n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104,
         n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112,
         n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120,
         n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128,
         n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136,
         n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144,
         n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152,
         n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160,
         n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168,
         n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176,
         n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184,
         n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192,
         n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200,
         n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208,
         n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216,
         n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224,
         n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232,
         n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240,
         n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248,
         n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256,
         n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264,
         n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272,
         n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280,
         n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288,
         n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296,
         n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304,
         n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312,
         n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320,
         n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328,
         n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336,
         n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344,
         n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352,
         n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360,
         n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368,
         n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376,
         n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384,
         n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392,
         n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,
         n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408,
         n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416,
         n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,
         n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432,
         n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440,
         n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448,
         n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456,
         n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464,
         n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472,
         n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480,
         n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488,
         n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496,
         n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504,
         n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512,
         n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520,
         n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528,
         n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536,
         n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544,
         n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552,
         n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560,
         n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568,
         n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576,
         n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584,
         n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592,
         n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600,
         n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608,
         n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616,
         n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624,
         n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632,
         n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640,
         n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648,
         n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656,
         n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664,
         n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672,
         n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680,
         n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688,
         n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696,
         n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704,
         n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712,
         n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720,
         n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728,
         n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736,
         n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744,
         n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752,
         n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760,
         n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768,
         n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776,
         n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784,
         n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792,
         n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800,
         n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808,
         n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816,
         n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824,
         n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832,
         n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840,
         n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848,
         n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856,
         n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864,
         n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872,
         n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880,
         n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888,
         n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896,
         n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904,
         n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912,
         n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920,
         n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928,
         n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936,
         n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944,
         n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952,
         n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960,
         n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968,
         n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976,
         n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984,
         n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992,
         n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000,
         n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008,
         n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016,
         n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024,
         n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032,
         n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040,
         n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048,
         n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056,
         n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064,
         n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072,
         n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080,
         n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088,
         n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096,
         n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104,
         n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112,
         n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120,
         n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128,
         n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136,
         n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144,
         n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152,
         n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160,
         n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168,
         n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176,
         n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184,
         n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192,
         n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200,
         n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208,
         n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216,
         n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224,
         n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232,
         n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240,
         n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248,
         n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256,
         n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264,
         n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272,
         n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280,
         n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288,
         n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296,
         n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304,
         n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312,
         n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320,
         n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328,
         n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336,
         n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344,
         n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352,
         n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360,
         n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368,
         n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376,
         n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384,
         n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392,
         n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400,
         n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408,
         n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416,
         n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424,
         n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432,
         n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440,
         n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448,
         n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456,
         n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464,
         n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472,
         n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480,
         n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488,
         n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496,
         n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504,
         n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512,
         n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520,
         n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528,
         n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536,
         n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544,
         n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552,
         n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560,
         n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568,
         n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576,
         n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584,
         n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592,
         n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600,
         n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608,
         n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616,
         n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624,
         n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632,
         n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640,
         n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648,
         n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656,
         n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664,
         n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672,
         n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680,
         n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688,
         n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696,
         n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704,
         n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712,
         n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720,
         n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728,
         n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736,
         n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744,
         n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752,
         n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760,
         n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768,
         n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776,
         n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784,
         n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792,
         n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800,
         n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808,
         n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816,
         n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824,
         n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832,
         n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840,
         n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848,
         n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856,
         n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864,
         n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872,
         n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880,
         n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888,
         n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896,
         n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904,
         n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912,
         n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920,
         n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928,
         n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936,
         n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944,
         n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952,
         n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960,
         n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968,
         n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976,
         n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984,
         n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992,
         n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000,
         n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008,
         n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016,
         n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024,
         n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032,
         n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040,
         n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048,
         n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056,
         n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064,
         n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072,
         n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080,
         n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088,
         n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096,
         n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104,
         n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112,
         n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120,
         n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128,
         n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136,
         n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144,
         n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152,
         n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160,
         n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168,
         n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176,
         n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184,
         n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192,
         n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200,
         n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208,
         n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216,
         n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224,
         n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232,
         n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240,
         n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248,
         n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256,
         n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264,
         n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272,
         n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280,
         n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288,
         n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296,
         n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304,
         n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312,
         n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320,
         n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328,
         n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336,
         n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344,
         n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352,
         n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360,
         n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368,
         n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376,
         n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384,
         n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392,
         n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400,
         n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408,
         n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416,
         n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424,
         n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432,
         n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440,
         n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448,
         n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456,
         n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464,
         n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472,
         n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480,
         n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488,
         n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496,
         n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504,
         n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512,
         n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520,
         n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528,
         n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536,
         n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544,
         n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552,
         n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560,
         n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568,
         n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576,
         n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584,
         n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592,
         n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600,
         n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608,
         n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616,
         n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624,
         n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632,
         n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640,
         n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648,
         n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656,
         n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664,
         n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672,
         n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680,
         n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688,
         n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696,
         n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704,
         n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712,
         n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720,
         n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728,
         n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736,
         n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744,
         n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752,
         n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760,
         n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768,
         n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776,
         n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784,
         n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792,
         n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800,
         n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808,
         n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816,
         n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824,
         n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832,
         n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840,
         n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848,
         n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856,
         n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864,
         n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872,
         n20873, n20874, n20875, n20876, n20877, n20878, n20879, n20880,
         n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888,
         n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896,
         n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904,
         n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912,
         n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920,
         n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928,
         n20929, n20930, n20931, n20932, n20933, n20934, n20935, n20936,
         n20937, n20938, n20939, n20940, n20941, n20942, n20943, n20944,
         n20945, n20946, n20947, n20948, n20949, n20950, n20951, n20952,
         n20953, n20954, n20955, n20956, n20957, n20958, n20959, n20960,
         n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968,
         n20969, n20970, n20971, n20972, n20973, n20974, n20975, n20976,
         n20977, n20978, n20979, n20980, n20981, n20982, n20983, n20984,
         n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992,
         n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000,
         n21001, n21002, n21003, n21004, n21005, n21006, n21007, n21008,
         n21009, n21010, n21011, n21012, n21013, n21014, n21015, n21016,
         n21017, n21018, n21019, n21020, n21021, n21022, n21023, n21024,
         n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032,
         n21033, n21034, n21035, n21036, n21037, n21038, n21039, n21040,
         n21041, n21042, n21043, n21044, n21045, n21046, n21047, n21048,
         n21049, n21050, n21051, n21052, n21053, n21054, n21055, n21056,
         n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21064,
         n21065, n21066, n21067, n21068, n21069, n21070, n21071, n21072,
         n21073, n21074, n21075, n21076, n21077, n21078, n21079, n21080,
         n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088,
         n21089, n21090, n21091, n21092, n21093, n21094, n21095, n21096,
         n21097, n21098, n21099, n21100, n21101, n21102, n21103, n21104,
         n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21112,
         n21113, n21114, n21115, n21116, n21117, n21118, n21119, n21120,
         n21121, n21122, n21123, n21124, n21125, n21126, n21127, n21128,
         n21129, n21130, n21131, n21132, n21133, n21134, n21135, n21136,
         n21137, n21138, n21139, n21140, n21141, n21142, n21143, n21144,
         n21145, n21146, n21147, n21148, n21149, n21150, n21151, n21152,
         n21153, n21154, n21155, n21156, n21157, n21158, n21159, n21160,
         n21161, n21162, n21163, n21164, n21165, n21166, n21167, n21168,
         n21169, n21170, n21171, n21172, n21173, n21174, n21175, n21176,
         n21177, n21178, n21179, n21180, n21181, n21182, n21183, n21184,
         n21185, n21186, n21187, n21188, n21189, n21190, n21191, n21192,
         n21193, n21194, n21195, n21196, n21197, n21198, n21199, n21200,
         n21201, n21202, n21203, n21204, n21205, n21206, n21207, n21208,
         n21209, n21210, n21211, n21212, n21213, n21214, n21215, n21216,
         n21217, n21218, n21219, n21220, n21221, n21222, n21223, n21224,
         n21225, n21226, n21227, n21228, n21229, n21230, n21231, n21232,
         n21233, n21234, n21235, n21236, n21237, n21238, n21239, n21240,
         n21241, n21242, n21243, n21244, n21245, n21246, n21247, n21248,
         n21249, n21250, n21251, n21252, n21253, n21254, n21255, n21256,
         n21257, n21258, n21259, n21260, n21261, n21262, n21263, n21264,
         n21265, n21266, n21267, n21268, n21269, n21270, n21271, n21272,
         n21273, n21274, n21275, n21276, n21277, n21278, n21279, n21280,
         n21281, n21282, n21283, n21284, n21285, n21286, n21287, n21288,
         n21289, n21290, n21291, n21292, n21293, n21294, n21295, n21296,
         n21297, n21298, n21299, n21300, n21301, n21302, n21303, n21304,
         n21305, n21306, n21307, n21308, n21309, n21310, n21311, n21312,
         n21313, n21314, n21315, n21316, n21317, n21318, n21319, n21320,
         n21321, n21322, n21323, n21324, n21325, n21326, n21327, n21328,
         n21329, n21330, n21331, n21332, n21333, n21334, n21335, n21336,
         n21337, n21338, n21339, n21340, n21341, n21342, n21343, n21344,
         n21345, n21346, n21347, n21348, n21349, n21350, n21351, n21352,
         n21353, n21354, n21355, n21356, n21357, n21358, n21359, n21360,
         n21361, n21362, n21363, n21364, n21365, n21366, n21367, n21368,
         n21369, n21370, n21371, n21372, n21373, n21374, n21375, n21376,
         n21377, n21378, n21379, n21380, n21381, n21382, n21383, n21384,
         n21385, n21386, n21387, n21388, n21389, n21390, n21391, n21392,
         n21393, n21394, n21395, n21396, n21397, n21398, n21399, n21400,
         n21401, n21402, n21403, n21404, n21405, n21406, n21407, n21408,
         n21409, n21410, n21411, n21412, n21413, n21414, n21415, n21416,
         n21417, n21418, n21419, n21420, n21421, n21422, n21423, n21424,
         n21425, n21426, n21427, n21428, n21429, n21430, n21431, n21432,
         n21433, n21434, n21435, n21436, n21437, n21438, n21439, n21440,
         n21441, n21442, n21443, n21444, n21445, n21446, n21447, n21448,
         n21449, n21450, n21451, n21452, n21453, n21454, n21455, n21456,
         n21457, n21458, n21459, n21460, n21461, n21462, n21463, n21464,
         n21465, n21466, n21467, n21468, n21469, n21470, n21471, n21472,
         n21473, n21474, n21475, n21476, n21477, n21478, n21479, n21480,
         n21481, n21482, n21483, n21484, n21485, n21486, n21487, n21488,
         n21489, n21490, n21491, n21492, n21493, n21494, n21495, n21496,
         n21497, n21498, n21499, n21500, n21501, n21502, n21503, n21504,
         n21505, n21506, n21507, n21508, n21509, n21510, n21511, n21512,
         n21513, n21514, n21515, n21516, n21517, n21518, n21519, n21520,
         n21521, n21522, n21523, n21524, n21525, n21526, n21527, n21528,
         n21529, n21530, n21531, n21532, n21533, n21534, n21535, n21536,
         n21537, n21538, n21539, n21540, n21541, n21542, n21543, n21544,
         n21545, n21546, n21547, n21548, n21549, n21550, n21551, n21552,
         n21553, n21554, n21555, n21556, n21557, n21558, n21559, n21560,
         n21561, n21562, n21563, n21564, n21565, n21566, n21567, n21568,
         n21569, n21570, n21571, n21572, n21573, n21574, n21575, n21576,
         n21577, n21578, n21579, n21580, n21581, n21582, n21583, n21584,
         n21585, n21586, n21587, n21588, n21589, n21590, n21591, n21592,
         n21593, n21594, n21595, n21596, n21597, n21598, n21599, n21600,
         n21601, n21602, n21603, n21604, n21605, n21606, n21607, n21608,
         n21609, n21610, n21611, n21612, n21613, n21614, n21615, n21616,
         n21617, n21618, n21619, n21620, n21621, n21622, n21623, n21624,
         n21625, n21626, n21627, n21628, n21629, n21630, n21631, n21632,
         n21633, n21634, n21635, n21636, n21637, n21638, n21639, n21640,
         n21641, n21642, n21643, n21644, n21645, n21646, n21647, n21648,
         n21649, n21650, n21651, n21652, n21653, n21654, n21655, n21656,
         n21657, n21658, n21659, n21660, n21661, n21662, n21663, n21664,
         n21665, n21666, n21667, n21668, n21669, n21670, n21671, n21672,
         n21673, n21674, n21675, n21676, n21677, n21678, n21679, n21680,
         n21681, n21682, n21683, n21684, n21685, n21686, n21687, n21688,
         n21689, n21690, n21691, n21692, n21693, n21694, n21695, n21696,
         n21697, n21698, n21699, n21700, n21701, n21702, n21703, n21704,
         n21705, n21706, n21707, n21708, n21709, n21710, n21711, n21712,
         n21713, n21714, n21715, n21716, n21717, n21718, n21719, n21720,
         n21721, n21722, n21723, n21724, n21725, n21726, n21727, n21728,
         n21729, n21730, n21731, n21732, n21733, n21734, n21735, n21736,
         n21737, n21738, n21739, n21740, n21741, n21742, n21743, n21744,
         n21745, n21746, n21747, n21748, n21749, n21750, n21751, n21752,
         n21753, n21754, n21755, n21756, n21757, n21758, n21759, n21760,
         n21761, n21762, n21763, n21764, n21765, n21766, n21767, n21768,
         n21769, n21770, n21771, n21772, n21773, n21774, n21775, n21776,
         n21777, n21778, n21779, n21780, n21781, n21782, n21783, n21784,
         n21785, n21786, n21787, n21788, n21789, n21790, n21791, n21792,
         n21793, n21794, n21795, n21796, n21797, n21798, n21799, n21800,
         n21801, n21802, n21803, n21804, n21805, n21806, n21807, n21808,
         n21809, n21810, n21811, n21812, n21813, n21814, n21815, n21816,
         n21817, n21818, n21819, n21820, n21821, n21822, n21823, n21824,
         n21825, n21826, n21827, n21828, n21829, n21830, n21831, n21832,
         n21833, n21834, n21835, n21836, n21837, n21838, n21839, n21840,
         n21841, n21842, n21843, n21844, n21845, n21846, n21847, n21848,
         n21849, n21850, n21851, n21852, n21853, n21854, n21855, n21856,
         n21857, n21858, n21859, n21860, n21861, n21862, n21863, n21864,
         n21865, n21866, n21867, n21868, n21869, n21870, n21871, n21872,
         n21873, n21874, n21875, n21876, n21877, n21878, n21879, n21880,
         n21881, n21882, n21883, n21884, n21885, n21886, n21887, n21888,
         n21889, n21890, n21891, n21892, n21893, n21894, n21895, n21896,
         n21897, n21898, n21899, n21900, n21901, n21902, n21903, n21904,
         n21905, n21906, n21907, n21908, n21909, n21910, n21911, n21912,
         n21913, n21914, n21915, n21916, n21917, n21918, n21919, n21920,
         n21921, n21922, n21923, n21924, n21925, n21926, n21927, n21928,
         n21929, n21930, n21931, n21932, n21933, n21934, n21935, n21936,
         n21937, n21938, n21939, n21940, n21941, n21942, n21943, n21944,
         n21945, n21946, n21947, n21948, n21949, n21950, n21951, n21952,
         n21953, n21954, n21955, n21956, n21957, n21958, n21959, n21960,
         n21961, n21962, n21963, n21964, n21965, n21966, n21967, n21968,
         n21969, n21970, n21971, n21972, n21973, n21974, n21975, n21976,
         n21977, n21978, n21979, n21980, n21981, n21982, n21983, n21984,
         n21985, n21986, n21987, n21988, n21989, n21990, n21991, n21992,
         n21993, n21994, n21995, n21996, n21997, n21998, n21999, n22000,
         n22001, n22002, n22003, n22004, n22005, n22006, n22007, n22008,
         n22009, n22010, n22011, n22012, n22013, n22014, n22015, n22016,
         n22017, n22018, n22019, n22020, n22021, n22022, n22023, n22024,
         n22025, n22026, n22027, n22028, n22029, n22030, n22031, n22032,
         n22033, n22034, n22035, n22036, n22037, n22038, n22039, n22040,
         n22041, n22042, n22043, n22044, n22045, n22046, n22047, n22048,
         n22049, n22050, n22051, n22052, n22053, n22054, n22055, n22056,
         n22057, n22058, n22059, n22060, n22061, n22062, n22063, n22064,
         n22065, n22066, n22067, n22068, n22069, n22070, n22071, n22072,
         n22073, n22074, n22075, n22076, n22077, n22078, n22079, n22080,
         n22081, n22082, n22083, n22084, n22085, n22086, n22087, n22088,
         n22089, n22090, n22091, n22092, n22093, n22094, n22095, n22096,
         n22097, n22098, n22099, n22100, n22101, n22102, n22103, n22104,
         n22105, n22106, n22107, n22108, n22109, n22110, n22111, n22112,
         n22113, n22114, n22115, n22116, n22117, n22118, n22119, n22120,
         n22121, n22122, n22123, n22124, n22125, n22126, n22127, n22128,
         n22129, n22130, n22131, n22132, n22133, n22134, n22135, n22136,
         n22137, n22138, n22139, n22140, n22141, n22142, n22143, n22144,
         n22145, n22146, n22147, n22148, n22149, n22150, n22151, n22152,
         n22153, n22154, n22155, n22156, n22157, n22158, n22159, n22160,
         n22161, n22162, n22163, n22164, n22165, n22166, n22167, n22168,
         n22169, n22170, n22171, n22172, n22173, n22174, n22175, n22176,
         n22177, n22178, n22179, n22180, n22181, n22182, n22183, n22184,
         n22185, n22186, n22187, n22188, n22189, n22190, n22191, n22192,
         n22193, n22194, n22195, n22196, n22197, n22198, n22199, n22200,
         n22201, n22202, n22203, n22204, n22205, n22206, n22207, n22208,
         n22209, n22210, n22211, n22212, n22213, n22214, n22215, n22216,
         n22217, n22218, n22219, n22220, n22221, n22222, n22223, n22224,
         n22225, n22226, n22227, n22228, n22229, n22230, n22231, n22232,
         n22233, n22234, n22235, n22236, n22237, n22238, n22239, n22240,
         n22241, n22242, n22243, n22244, n22245, n22246, n22247, n22248,
         n22249, n22250, n22251, n22252, n22253, n22254, n22255, n22256,
         n22257, n22258, n22259, n22260, n22261, n22262, n22263, n22264,
         n22265, n22266, n22267, n22268, n22269, n22270, n22271, n22272,
         n22273, n22274, n22275, n22276, n22277, n22278, n22279, n22280,
         n22281, n22282, n22283, n22284, n22285, n22286, n22287, n22288,
         n22289, n22290, n22291, n22292, n22293, n22294, n22295, n22296,
         n22297, n22298, n22299, n22300, n22301, n22302, n22303, n22304,
         n22305, n22306, n22307, n22308, n22309, n22310, n22311, n22312,
         n22313, n22314, n22315, n22316, n22317, n22318, n22319, n22320,
         n22321, n22322, n22323, n22324, n22325, n22326, n22327, n22328,
         n22329, n22330, n22331, n22332, n22333, n22334, n22335, n22336,
         n22337, n22338, n22339, n22340, n22341, n22342, n22343, n22344,
         n22345, n22346, n22347, n22348, n22349, n22350, n22351, n22352,
         n22353, n22354, n22355, n22356, n22357, n22358, n22359, n22360,
         n22361, n22362, n22363, n22364, n22365, n22366, n22367, n22368,
         n22369, n22370, n22371, n22372, n22373, n22374, n22375, n22376,
         n22377, n22378, n22379, n22380, n22381, n22382, n22383, n22384,
         n22385, n22386, n22387, n22388, n22389, n22390, n22391, n22392,
         n22393, n22394, n22395, n22396, n22397, n22398, n22399, n22400,
         n22401, n22402, n22403, n22404, n22405, n22406, n22407, n22408,
         n22409, n22410, n22411, n22412, n22413, n22414, n22415, n22416,
         n22417, n22418, n22419, n22420, n22421, n22422, n22423, n22424,
         n22425, n22426, n22427, n22428, n22429, n22430, n22431, n22432,
         n22433, n22434, n22435, n22436, n22437, n22438, n22439, n22440,
         n22441, n22442, n22443, n22444, n22445, n22446, n22447, n22448,
         n22449, n22450, n22451, n22452, n22453, n22454, n22455, n22456,
         n22457, n22458, n22459, n22460, n22461, n22462, n22463, n22464,
         n22465, n22466, n22467, n22468, n22469, n22470, n22471, n22472,
         n22473, n22474, n22475, n22476, n22477, n22478, n22479, n22480,
         n22481, n22482, n22483, n22484, n22485, n22486, n22487, n22488,
         n22489, n22490, n22491, n22492, n22493, n22494, n22495, n22496,
         n22497, n22498, n22499, n22500, n22501, n22502, n22503, n22504,
         n22505, n22506, n22507, n22508, n22509, n22510, n22511, n22512,
         n22513, n22514, n22515, n22516, n22517, n22518, n22519, n22520,
         n22521, n22522, n22523, n22524, n22525, n22526, n22527, n22528,
         n22529, n22530, n22531, n22532, n22533, n22534, n22535, n22536,
         n22537, n22538, n22539, n22540, n22541, n22542, n22543, n22544,
         n22545, n22546, n22547, n22548, n22549, n22550, n22551, n22552,
         n22553, n22554, n22555, n22556, n22557, n22558, n22559, n22560,
         n22561, n22562, n22563, n22564, n22565, n22566, n22567, n22568,
         n22569, n22570, n22571, n22572, n22573, n22574, n22575, n22576,
         n22577, n22578, n22579, n22580, n22581, n22582, n22583, n22584,
         n22585, n22586, n22587, n22588, n22589, n22590, n22591, n22592,
         n22593, n22594, n22595, n22596, n22597, n22598, n22599, n22600,
         n22601, n22602, n22603, n22604, n22605, n22606, n22607, n22608,
         n22609, n22610, n22611, n22612, n22613, n22614, n22615, n22616,
         n22617, n22618, n22619, n22620, n22621, n22622, n22623, n22624,
         n22625, n22626, n22627, n22628, n22629, n22630, n22631, n22632,
         n22633, n22634, n22635, n22636, n22637, n22638, n22639, n22640,
         n22641, n22642, n22643, n22644, n22645, n22646, n22647, n22648,
         n22649, n22650, n22651, n22652, n22653, n22654, n22655, n22656,
         n22657, n22658, n22659, n22660, n22661, n22662, n22663, n22664,
         n22665, n22666, n22667, n22668, n22669, n22670, n22671, n22672,
         n22673, n22674, n22675, n22676, n22677, n22678, n22679, n22680,
         n22681, n22682, n22683, n22684, n22685, n22686, n22687, n22688,
         n22689, n22690, n22691, n22692, n22693, n22694, n22695, n22696,
         n22697, n22698, n22699, n22700, n22701, n22702, n22703, n22704,
         n22705, n22706, n22707, n22708, n22709, n22710, n22711, n22712,
         n22713, n22714, n22715, n22716, n22717, n22718, n22719, n22720,
         n22721, n22722, n22723, n22724, n22725, n22726, n22727, n22728,
         n22729, n22730, n22731, n22732, n22733, n22734, n22735, n22736,
         n22737, n22738, n22739, n22740, n22741, n22742, n22743, n22744,
         n22745, n22746, n22747, n22748, n22749, n22750, n22751, n22752,
         n22753, n22754, n22755, n22756, n22757, n22758, n22759, n22760,
         n22761, n22762, n22763, n22764, n22765, n22766, n22767, n22768,
         n22769, n22770, n22771, n22772, n22773, n22774, n22775, n22776,
         n22777, n22778, n22779, n22780, n22781, n22782, n22783, n22784,
         n22785, n22786, n22787, n22788, n22789, n22790, n22791, n22792,
         n22793, n22794, n22795, n22796, n22797, n22798, n22799, n22800,
         n22801, n22802, n22803, n22804, n22805, n22806, n22807, n22808,
         n22809, n22810, n22811, n22812, n22813, n22814, n22815, n22816,
         n22817, n22818, n22819, n22820, n22821, n22822, n22823, n22824,
         n22825, n22826, n22827, n22828, n22829, n22830, n22831, n22832,
         n22833, n22834, n22835, n22836, n22837, n22838, n22839, n22840,
         n22841, n22842, n22843, n22844, n22845, n22846, n22847, n22848,
         n22849, n22850, n22851, n22852, n22853, n22854, n22855, n22856,
         n22857, n22858, n22859, n22860, n22861, n22862, n22863, n22864,
         n22865, n22866, n22867, n22868, n22869, n22870, n22871, n22872,
         n22873, n22874, n22875, n22876, n22877, n22878, n22879, n22880,
         n22881, n22882, n22883, n22884, n22885, n22886, n22887, n22888,
         n22889, n22890, n22891, n22892, n22893, n22894, n22895, n22896,
         n22897, n22898, n22899, n22900, n22901, n22902, n22903, n22904,
         n22905, n22906, n22907, n22908, n22909, n22910, n22911, n22912,
         n22913, n22914, n22915, n22916, n22917, n22918, n22919, n22920,
         n22921, n22922, n22923, n22924, n22925, n22926, n22927, n22928,
         n22929, n22930, n22931, n22932, n22933, n22934, n22935, n22936,
         n22937, n22938, n22939, n22940, n22941, n22942, n22943, n22944,
         n22945, n22946, n22947, n22948, n22949, n22950, n22951, n22952,
         n22953, n22954, n22955, n22956, n22957, n22958, n22959, n22960,
         n22961, n22962, n22963, n22964, n22965, n22966, n22967, n22968,
         n22969, n22970, n22971, n22972, n22973, n22974, n22975, n22976,
         n22977, n22978, n22979, n22980, n22981, n22982, n22983, n22984,
         n22985, n22986, n22987, n22988, n22989, n22990, n22991, n22992,
         n22993, n22994, n22995, n22996, n22997, n22998, n22999, n23000,
         n23001, n23002, n23003, n23004, n23005, n23006, n23007, n23008,
         n23009, n23010, n23011, n23012, n23013, n23014, n23015, n23016,
         n23017, n23018, n23019, n23020, n23021, n23022, n23023, n23024,
         n23025, n23026, n23027, n23028, n23029, n23030, n23031, n23032,
         n23033, n23034, n23035, n23036, n23037, n23038, n23039, n23040,
         n23041, n23042, n23043, n23044, n23045, n23046, n23047, n23048,
         n23049, n23050, n23051, n23052, n23053, n23054, n23055, n23056,
         n23057, n23058, n23059, n23060, n23061, n23062, n23063, n23064,
         n23065, n23066, n23067, n23068, n23069, n23070, n23071, n23072,
         n23073, n23074, n23075, n23076, n23077, n23078, n23079, n23080,
         n23081, n23082, n23083, n23084, n23085, n23086, n23087, n23088,
         n23089, n23090, n23091, n23092, n23093, n23094, n23095, n23096,
         n23097, n23098, n23099, n23100, n23101, n23102, n23103, n23104,
         n23105, n23106, n23107, n23108, n23109, n23110, n23111, n23112,
         n23113, n23114, n23115, n23116, n23117, n23118, n23119, n23120,
         n23121, n23122, n23123, n23124, n23125, n23126, n23127, n23128,
         n23129, n23130, n23131, n23132, n23133, n23134, n23135, n23136,
         n23137, n23138, n23139, n23140, n23141, n23142, n23143, n23144,
         n23145, n23146, n23147, n23148, n23149, n23150, n23151, n23152,
         n23153, n23154, n23155, n23156, n23157, n23158, n23159, n23160,
         n23161, n23162, n23163, n23164, n23165, n23166, n23167, n23168,
         n23169, n23170, n23171, n23172, n23173, n23174, n23175, n23176,
         n23177, n23178, n23179, n23180, n23181, n23182, n23183, n23184,
         n23185, n23186, n23187, n23188, n23189, n23190, n23191, n23192,
         n23193, n23194, n23195, n23196, n23197, n23198, n23199, n23200,
         n23201, n23202, n23203, n23204, n23205, n23206, n23207, n23208,
         n23209, n23210, n23211, n23212, n23213, n23214, n23215, n23216,
         n23217, n23218, n23219, n23220, n23221, n23222, n23223, n23224,
         n23225, n23226, n23227, n23228, n23229, n23230, n23231, n23232,
         n23233, n23234, n23235, n23236, n23237, n23238, n23239, n23240,
         n23241, n23242, n23243, n23244, n23245, n23246, n23247, n23248,
         n23249, n23250, n23251, n23252, n23253, n23254, n23255, n23256,
         n23257, n23258, n23259, n23260, n23261, n23262, n23263, n23264,
         n23265, n23266, n23267, n23268, n23269, n23270, n23271, n23272,
         n23273, n23274, n23275, n23276, n23277, n23278, n23279, n23280,
         n23281, n23282, n23283, n23284, n23285, n23286, n23287, n23288,
         n23289, n23290, n23291, n23292, n23293, n23294, n23295, n23296,
         n23297, n23298, n23299, n23300, n23301, n23302, n23303, n23304,
         n23305, n23306, n23307, n23308, n23309, n23310, n23311, n23312,
         n23313, n23314, n23315, n23316, n23317, n23318, n23319, n23320,
         n23321, n23322, n23323, n23324, n23325, n23326, n23327, n23328,
         n23329, n23330, n23331, n23332, n23333, n23334, n23335, n23336,
         n23337, n23338, n23339, n23340, n23341, n23342, n23343, n23344,
         n23345, n23346, n23347, n23348, n23349, n23350, n23351, n23352,
         n23353, n23354, n23355, n23356, n23357, n23358, n23359, n23360,
         n23361, n23362, n23363, n23364, n23365, n23366, n23367, n23368,
         n23369, n23370, n23371, n23372, n23373, n23374, n23375, n23376,
         n23377, n23378, n23379, n23380, n23381, n23382, n23383, n23384,
         n23385, n23386, n23387, n23388, n23389, n23390, n23391, n23392,
         n23393, n23394, n23395, n23396, n23397, n23398, n23399, n23400,
         n23401, n23402, n23403, n23404, n23405, n23406, n23407, n23408,
         n23409, n23410, n23411, n23412, n23413, n23414, n23415, n23416,
         n23417, n23418, n23419, n23420, n23421, n23422, n23423, n23424,
         n23425, n23426, n23427, n23428, n23429, n23430, n23431, n23432,
         n23433, n23434, n23435, n23436, n23437, n23438, n23439, n23440,
         n23441, n23442, n23443, n23444, n23445, n23446, n23447, n23448,
         n23449, n23450, n23451, n23452, n23453, n23454, n23455, n23456,
         n23457, n23458, n23459, n23460, n23461, n23462, n23463, n23464,
         n23465, n23466, n23467, n23468, n23469, n23470, n23471, n23472,
         n23473, n23474, n23475, n23476, n23477, n23478, n23479, n23480,
         n23481, n23482, n23483, n23484, n23485, n23486, n23487, n23488,
         n23489, n23490, n23491, n23492, n23493, n23494, n23495, n23496,
         n23497, n23498, n23499, n23500, n23501, n23502, n23503, n23504,
         n23505, n23506, n23507, n23508, n23509, n23510, n23511, n23512,
         n23513, n23514, n23515, n23516, n23517, n23518, n23519, n23520,
         n23521, n23522, n23523, n23524, n23525, n23526, n23527, n23528,
         n23529, n23530, n23531, n23532, n23533, n23534, n23535, n23536,
         n23537, n23538, n23539, n23540, n23541, n23542, n23543, n23544,
         n23545, n23546, n23547, n23548, n23549, n23550, n23551, n23552,
         n23553, n23554, n23555, n23556, n23557, n23558, n23559, n23560,
         n23561, n23562, n23563, n23564, n23565, n23566, n23567, n23568,
         n23569, n23570, n23571, n23572, n23573, n23574, n23575, n23576,
         n23577, n23578, n23579, n23580, n23581, n23582, n23583, n23584,
         n23585, n23586, n23587, n23588, n23589, n23590, n23591, n23592,
         n23593, n23594, n23595, n23596, n23597, n23598, n23599, n23600,
         n23601, n23602, n23603, n23604, n23605, n23606, n23607, n23608,
         n23609, n23610, n23611, n23612, n23613, n23614, n23615, n23616,
         n23617, n23618, n23619, n23620, n23621, n23622, n23623, n23624,
         n23625, n23626, n23627, n23628, n23629, n23630, n23631, n23632,
         n23633, n23634, n23635, n23636, n23637, n23638, n23639, n23640,
         n23641, n23642, n23643, n23644, n23645, n23646, n23647, n23648,
         n23649, n23650, n23651, n23652, n23653, n23654, n23655, n23656,
         n23657, n23658, n23659, n23660, n23661, n23662, n23663, n23664,
         n23665, n23666, n23667, n23668, n23669, n23670, n23671, n23672,
         n23673, n23674, n23675, n23676, n23677, n23678, n23679, n23680,
         n23681, n23682, n23683, n23684, n23685, n23686, n23687, n23688,
         n23689, n23690, n23691, n23692, n23693, n23694, n23695, n23696,
         n23697, n23698, n23699, n23700, n23701, n23702, n23703, n23704,
         n23705, n23706, n23707, n23708, n23709, n23710, n23711, n23712,
         n23713, n23714, n23715, n23716, n23717, n23718, n23719, n23720,
         n23721, n23722, n23723, n23724, n23725, n23726, n23727, n23728,
         n23729, n23730, n23731, n23732, n23733, n23734, n23735, n23736,
         n23737, n23738, n23739, n23740, n23741, n23742, n23743, n23744,
         n23745, n23746, n23747, n23748, n23749, n23750, n23751, n23752,
         n23753, n23754, n23755, n23756, n23757, n23758, n23759, n23760,
         n23761, n23762, n23763, n23764, n23765, n23766, n23767, n23768,
         n23769, n23770, n23771, n23772, n23773, n23774, n23775, n23776,
         n23777, n23778, n23779, n23780, n23781, n23782, n23783, n23784,
         n23785, n23786, n23787, n23788, n23789, n23790, n23791, n23792,
         n23793, n23794, n23795, n23796, n23797, n23798, n23799, n23800,
         n23801, n23802, n23803, n23804, n23805, n23806, n23807, n23808,
         n23809, n23810, n23811, n23812, n23813, n23814, n23815, n23816,
         n23817, n23818, n23819, n23820, n23821, n23822, n23823, n23824,
         n23825, n23826, n23827, n23828, n23829, n23830, n23831, n23832,
         n23833, n23834, n23835, n23836, n23837, n23838, n23839, n23840,
         n23841, n23842, n23843, n23844, n23845, n23846, n23847, n23848,
         n23849, n23850, n23851, n23852, n23853, n23854, n23855, n23856,
         n23857, n23858, n23859, n23860, n23861, n23862, n23863, n23864,
         n23865, n23866, n23867, n23868, n23869, n23870, n23871, n23872,
         n23873, n23874, n23875, n23876, n23877, n23878, n23879, n23880,
         n23881, n23882, n23883, n23884, n23885, n23886, n23887, n23888,
         n23889, n23890, n23891, n23892, n23893, n23894, n23895, n23896,
         n23897, n23898, n23899, n23900, n23901, n23902, n23903, n23904,
         n23905, n23906, n23907, n23908, n23909, n23910, n23911, n23912,
         n23913, n23914, n23915, n23916, n23917, n23918, n23919, n23920,
         n23921, n23922, n23923, n23924, n23925, n23926, n23927, n23928,
         n23929, n23930, n23931, n23932, n23933, n23934, n23935, n23936,
         n23937, n23938, n23939, n23940, n23941, n23942, n23943, n23944,
         n23945, n23946, n23947, n23948, n23949, n23950, n23951, n23952,
         n23953, n23954, n23955, n23956, n23957, n23958, n23959, n23960,
         n23961, n23962, n23963, n23964, n23965, n23966, n23967, n23968,
         n23969, n23970, n23971, n23972, n23973, n23974, n23975, n23976,
         n23977, n23978, n23979, n23980, n23981, n23982, n23983, n23984,
         n23985, n23986, n23987, n23988, n23989, n23990, n23991, n23992,
         n23993, n23994, n23995, n23996, n23997, n23998, n23999, n24000,
         n24001, n24002, n24003, n24004, n24005, n24006, n24007, n24008,
         n24009, n24010, n24011, n24012, n24013, n24014, n24015, n24016,
         n24017, n24018, n24019, n24020, n24021, n24022, n24023, n24024,
         n24025, n24026, n24027, n24028, n24029, n24030, n24031, n24032,
         n24033, n24034, n24035, n24036, n24037, n24038, n24039, n24040,
         n24041, n24042, n24043, n24044, n24045, n24046, n24047, n24048,
         n24049, n24050, n24051, n24052, n24053, n24054, n24055, n24056,
         n24057, n24058, n24059, n24060, n24061, n24062, n24063, n24064,
         n24065, n24066, n24067, n24068, n24069, n24070, n24071, n24072,
         n24073, n24074, n24075, n24076, n24077, n24078, n24079, n24080,
         n24081, n24082, n24083, n24084, n24085, n24086, n24087, n24088,
         n24089, n24090, n24091, n24092, n24093, n24094, n24095, n24096,
         n24097, n24098, n24099, n24100, n24101, n24102, n24103, n24104,
         n24105, n24106, n24107, n24108, n24109, n24110, n24111, n24112,
         n24113, n24114, n24115, n24116, n24117, n24118, n24119, n24120,
         n24121, n24122, n24123, n24124, n24125, n24126, n24127, n24128,
         n24129, n24130, n24131, n24132, n24133, n24134, n24135, n24136,
         n24137, n24138, n24139, n24140, n24141, n24142, n24143, n24144,
         n24145, n24146, n24147, n24148, n24149, n24150, n24151, n24152,
         n24153, n24154, n24155, n24156, n24157, n24158, n24159, n24160,
         n24161, n24162, n24163, n24164, n24165, n24166, n24167, n24168,
         n24169, n24170, n24171, n24172, n24173, n24174, n24175, n24176,
         n24177, n24178, n24179, n24180, n24181, n24182, n24183, n24184,
         n24185, n24186, n24187, n24188, n24189, n24190, n24191, n24192,
         n24193, n24194, n24195, n24196, n24197, n24198, n24199, n24200,
         n24201, n24202, n24203, n24204, n24205, n24206, n24207, n24208,
         n24209, n24210, n24211, n24212, n24213, n24214, n24215, n24216,
         n24217, n24218, n24219, n24220, n24221, n24222, n24223, n24224,
         n24225, n24226, n24227, n24228, n24229, n24230, n24231, n24232,
         n24233, n24234, n24235, n24236, n24237, n24238, n24239, n24240,
         n24241, n24242, n24243, n24244, n24245, n24246, n24247, n24248,
         n24249, n24250, n24251, n24252, n24253, n24254, n24255, n24256,
         n24257, n24258, n24259, n24260, n24261, n24262, n24263, n24264,
         n24265, n24266, n24267, n24268, n24269, n24270, n24271, n24272,
         n24273, n24274, n24275, n24276, n24277, n24278, n24279, n24280,
         n24281, n24282, n24283, n24284, n24285, n24286, n24287, n24288,
         n24289, n24290, n24291, n24292, n24293, n24294, n24295, n24296,
         n24297, n24298, n24299, n24300, n24301, n24302, n24303, n24304,
         n24305, n24306, n24307, n24308, n24309, n24310, n24311, n24312,
         n24313, n24314, n24315, n24316, n24317, n24318, n24319, n24320,
         n24321, n24322, n24323, n24324, n24325, n24326, n24327, n24328,
         n24329, n24330, n24331, n24332, n24333, n24334, n24335, n24336,
         n24337, n24338, n24339, n24340, n24341, n24342, n24343, n24344,
         n24345, n24346, n24347, n24348, n24349, n24350, n24351, n24352,
         n24353, n24354, n24355, n24356, n24357, n24358, n24359, n24360,
         n24361, n24362, n24363, n24364, n24365, n24366, n24367, n24368,
         n24369, n24370, n24371, n24372, n24373, n24374, n24375, n24376,
         n24377, n24378, n24379, n24380, n24381, n24382, n24383, n24384,
         n24385, n24386, n24387, n24388, n24389, n24390, n24391, n24392,
         n24393, n24394, n24395, n24396, n24397, n24398, n24399, n24400,
         n24401, n24402, n24403, n24404, n24405, n24406, n24407, n24408,
         n24409, n24410, n24411, n24412, n24413, n24414, n24415, n24416,
         n24417, n24418, n24419, n24420, n24421, n24422, n24423, n24424,
         n24425, n24426, n24427, n24428, n24429, n24430, n24431, n24432,
         n24433, n24434, n24435, n24436, n24437, n24438, n24439, n24440,
         n24441, n24442, n24443, n24444, n24445, n24446, n24447, n24448,
         n24449, n24450, n24451, n24452, n24453, n24454, n24455, n24456,
         n24457, n24458, n24459, n24460, n24461, n24462, n24463, n24464,
         n24465, n24466, n24467, n24468, n24469, n24470, n24471, n24472,
         n24473, n24474, n24475, n24476, n24477, n24478, n24479, n24480,
         n24481, n24482, n24483, n24484, n24485, n24486, n24487, n24488,
         n24489, n24490, n24491, n24492, n24493, n24494, n24495, n24496,
         n24497, n24498, n24499, n24500, n24501, n24502, n24503, n24504,
         n24505, n24506, n24507, n24508, n24509, n24510, n24511, n24512,
         n24513, n24514, n24515, n24516, n24517, n24518, n24519, n24520,
         n24521, n24522, n24523, n24524, n24525, n24526, n24527, n24528,
         n24529, n24530, n24531, n24532, n24533, n24534, n24535, n24536,
         n24537, n24538, n24539, n24540, n24541, n24542, n24543, n24544,
         n24545, n24546, n24547, n24548, n24549, n24550, n24551, n24552,
         n24553, n24554, n24555, n24556, n24557, n24558, n24559, n24560,
         n24561, n24562, n24563, n24564, n24565, n24566, n24567, n24568,
         n24569, n24570, n24571, n24572, n24573, n24574, n24575, n24576,
         n24577, n24578, n24579, n24580, n24581, n24582, n24583, n24584,
         n24585, n24586, n24587, n24588, n24589, n24590, n24591, n24592,
         n24593, n24594, n24595, n24596, n24597, n24598, n24599, n24600,
         n24601, n24602, n24603, n24604, n24605, n24606, n24607, n24608,
         n24609, n24610, n24611, n24612, n24613, n24614, n24615, n24616,
         n24617, n24618, n24619, n24620, n24621, n24622, n24623, n24624,
         n24625, n24626, n24627, n24628, n24629, n24630, n24631, n24632,
         n24633, n24634, n24635, n24636, n24637, n24638, n24639, n24640,
         n24641, n24642, n24643, n24644, n24645, n24646, n24647, n24648,
         n24649, n24650, n24651, n24652, n24653, n24654, n24655, n24656,
         n24657, n24658, n24659, n24660, n24661, n24662, n24663, n24664,
         n24665, n24666, n24667, n24668, n24669, n24670, n24671, n24672,
         n24673, n24674, n24675, n24676, n24677, n24678, n24679, n24680,
         n24681, n24682, n24683, n24684, n24685, n24686, n24687, n24688,
         n24689, n24690, n24691, n24692, n24693, n24694, n24695, n24696,
         n24697, n24698, n24699, n24700, n24701, n24702, n24703, n24704,
         n24705, n24706, n24707, n24708, n24709, n24710, n24711, n24712,
         n24713, n24714, n24715, n24716, n24717, n24718, n24719, n24720,
         n24721, n24722, n24723, n24724, n24725, n24726, n24727, n24728,
         n24729, n24730, n24731, n24732, n24733, n24734, n24735, n24736,
         n24737, n24738, n24739, n24740, n24741, n24742, n24743, n24744,
         n24745, n24746, n24747, n24748, n24749, n24750, n24751, n24752,
         n24753, n24754, n24755, n24756, n24757, n24758, n24759, n24760,
         n24761, n24762, n24763, n24764, n24765, n24766, n24767, n24768,
         n24769, n24770, n24771, n24772, n24773, n24774, n24775, n24776,
         n24777, n24778, n24779, n24780, n24781, n24782, n24783, n24784,
         n24785, n24786, n24787, n24788, n24789, n24790, n24791, n24792,
         n24793, n24794, n24795, n24796, n24797, n24798, n24799, n24800,
         n24801, n24802, n24803, n24804, n24805, n24806, n24807, n24808,
         n24809, n24810, n24811, n24812, n24813, n24814, n24815, n24816,
         n24817, n24818, n24819, n24820, n24821, n24822, n24823, n24824,
         n24825, n24826, n24827, n24828, n24829, n24830, n24831, n24832,
         n24833, n24834, n24835, n24836, n24837, n24838, n24839, n24840,
         n24841, n24842, n24843, n24844, n24845, n24846, n24847, n24848,
         n24849, n24850, n24851, n24852, n24853, n24854, n24855, n24856,
         n24857, n24858, n24859, n24860, n24861, n24862, n24863, n24864,
         n24865, n24866, n24867, n24868, n24869, n24870, n24871, n24872,
         n24873, n24874, n24875, n24876, n24877, n24878, n24879, n24880,
         n24881, n24882, n24883, n24884, n24885, n24886, n24887, n24888,
         n24889, n24890, n24891, n24892, n24893, n24894, n24895, n24896,
         n24897, n24898, n24899, n24900, n24901, n24902, n24903, n24904,
         n24905, n24906, n24907, n24908, n24909, n24910, n24911, n24912,
         n24913, n24914, n24915, n24916, n24917, n24918, n24919, n24920,
         n24921, n24922, n24923, n24924, n24925, n24926, n24927, n24928,
         n24929, n24930, n24931, n24932, n24933, n24934, n24935, n24936,
         n24937, n24938, n24939, n24940, n24941, n24942, n24943, n24944,
         n24945, n24946, n24947, n24948, n24949, n24950, n24951, n24952,
         n24953, n24954, n24955, n24956, n24957, n24958, n24959, n24960,
         n24961, n24962, n24963, n24964, n24965, n24966, n24967, n24968,
         n24969, n24970, n24971, n24972, n24973, n24974, n24975, n24976,
         n24977, n24978, n24979, n24980, n24981, n24982, n24983, n24984,
         n24985, n24986, n24987, n24988, n24989, n24990, n24991, n24992,
         n24993, n24994, n24995, n24996, n24997, n24998, n24999, n25000,
         n25001, n25002, n25003, n25004, n25005, n25006, n25007, n25008,
         n25009, n25010, n25011, n25012, n25013, n25014, n25015, n25016,
         n25017, n25018, n25019, n25020, n25021, n25022, n25023, n25024,
         n25025, n25026, n25027, n25028, n25029, n25030, n25031, n25032,
         n25033, n25034, n25035, n25036, n25037, n25038, n25039, n25040,
         n25041, n25042, n25043, n25044, n25045, n25046, n25047, n25048,
         n25049, n25050, n25051, n25052, n25053, n25054, n25055, n25056,
         n25057, n25058, n25059, n25060, n25061, n25062, n25063, n25064,
         n25065, n25066, n25067, n25068, n25069, n25070, n25071, n25072,
         n25073, n25074, n25075, n25076, n25077, n25078, n25079, n25080,
         n25081, n25082, n25083, n25084, n25085, n25086, n25087, n25088,
         n25089, n25090, n25091, n25092, n25093, n25094, n25095, n25096,
         n25097, n25098, n25099, n25100, n25101, n25102, n25103, n25104,
         n25105, n25106, n25107, n25108, n25109, n25110, n25111, n25112,
         n25113, n25114, n25115, n25116, n25117, n25118, n25119, n25120,
         n25121, n25122, n25123, n25124, n25125, n25126, n25127, n25128,
         n25129, n25130, n25131, n25132, n25133, n25134, n25135, n25136,
         n25137, n25138, n25139, n25140, n25141, n25142, n25143, n25144,
         n25145, n25146, n25147, n25148, n25149, n25150, n25151, n25152,
         n25153, n25154, n25155, n25156, n25157, n25158, n25159, n25160,
         n25161, n25162, n25163, n25164, n25165, n25166, n25167, n25168,
         n25169, n25170, n25171, n25172, n25173, n25174, n25175, n25176,
         n25177, n25178, n25179, n25180, n25181, n25182, n25183, n25184,
         n25185, n25186, n25187, n25188, n25189, n25190, n25191, n25192,
         n25193, n25194, n25195, n25196, n25197, n25198, n25199, n25200,
         n25201, n25202, n25203, n25204, n25205, n25206, n25207, n25208,
         n25209, n25210, n25211, n25212, n25213, n25214, n25215, n25216,
         n25217, n25218, n25219, n25220, n25221, n25222, n25223, n25224,
         n25225, n25226, n25227, n25228, n25229, n25230, n25231, n25232,
         n25233, n25234, n25235, n25236, n25237, n25238, n25239, n25240,
         n25241, n25242, n25243, n25244, n25245, n25246, n25247, n25248,
         n25249, n25250, n25251, n25252, n25253, n25254, n25255, n25256,
         n25257, n25258, n25259, n25260, n25261, n25262, n25263, n25264,
         n25265, n25266, n25267, n25268, n25269, n25270, n25271, n25272,
         n25273, n25274, n25275, n25276, n25277, n25278, n25279, n25280,
         n25281, n25282, n25283, n25284, n25285, n25286, n25287, n25288,
         n25289, n25290, n25291, n25292, n25293, n25294, n25295, n25296,
         n25297, n25298, n25299, n25300, n25301, n25302, n25303, n25304,
         n25305, n25306, n25307, n25308, n25309, n25310, n25311, n25312,
         n25313, n25314, n25315, n25316, n25317, n25318, n25319, n25320,
         n25321, n25322, n25323, n25324, n25325, n25326, n25327, n25328,
         n25329, n25330, n25331, n25332, n25333, n25334, n25335, n25336,
         n25337, n25338, n25339, n25340, n25341, n25342, n25343, n25344,
         n25345, n25346, n25347, n25348, n25349, n25350, n25351, n25352,
         n25353, n25354, n25355, n25356, n25357, n25358, n25359, n25360,
         n25361, n25362, n25363, n25364, n25365, n25366, n25367, n25368,
         n25369, n25370, n25371, n25372, n25373, n25374, n25375, n25376,
         n25377, n25378, n25379, n25380, n25381, n25382, n25383, n25384,
         n25385, n25386, n25387, n25388, n25389, n25390, n25391, n25392,
         n25393, n25394, n25395, n25396, n25397, n25398, n25399, n25400,
         n25401, n25402, n25403, n25404, n25405, n25406, n25407, n25408,
         n25409, n25410, n25411, n25412, n25413, n25414, n25415, n25416,
         n25417, n25418, n25419, n25420, n25421, n25422, n25423, n25424,
         n25425, n25426, n25427, n25428, n25429, n25430, n25431, n25432,
         n25433, n25434, n25435, n25436, n25437, n25438, n25439, n25440,
         n25441, n25442, n25443, n25444, n25445, n25446, n25447, n25448,
         n25449, n25450, n25451, n25452, n25453, n25454, n25455, n25456,
         n25457, n25458, n25459, n25460, n25461, n25462, n25463, n25464,
         n25465, n25466, n25467, n25468, n25469, n25470, n25471, n25472,
         n25473, n25474, n25475, n25476, n25477, n25478, n25479, n25480,
         n25481, n25482, n25483, n25484, n25485, n25486, n25487, n25488,
         n25489, n25490, n25491, n25492, n25493, n25494, n25495, n25496,
         n25497, n25498, n25499, n25500, n25501, n25502, n25503, n25504,
         n25505, n25506, n25507, n25508, n25509, n25510, n25511, n25512,
         n25513, n25514, n25515, n25516, n25517, n25518, n25519, n25520,
         n25521, n25522, n25523, n25524, n25525, n25526, n25527, n25528,
         n25529, n25530, n25531, n25532, n25533, n25534, n25535, n25536,
         n25537, n25538, n25539, n25540, n25541, n25542, n25543, n25544,
         n25545, n25546, n25547, n25548, n25549, n25550, n25551, n25552,
         n25553, n25554, n25555, n25556, n25557, n25558, n25559, n25560,
         n25561, n25562, n25563, n25564, n25565, n25566, n25567, n25568,
         n25569, n25570, n25571, n25572, n25573, n25574, n25575, n25576,
         n25577, n25578, n25579, n25580, n25581, n25582, n25583, n25584,
         n25585, n25586, n25587, n25588, n25589, n25590, n25591, n25592,
         n25593, n25594, n25595, n25596, n25597, n25598, n25599, n25600,
         n25601, n25602, n25603, n25604, n25605, n25606, n25607, n25608,
         n25609, n25610, n25611, n25612, n25613, n25614, n25615, n25616,
         n25617, n25618, n25619, n25620, n25621, n25622, n25623, n25624,
         n25625, n25626, n25627, n25628, n25629, n25630, n25631, n25632,
         n25633, n25634, n25635, n25636, n25637, n25638, n25639, n25640,
         n25641, n25642, n25643, n25644, n25645, n25646, n25647, n25648,
         n25649, n25650, n25651, n25652, n25653, n25654, n25655, n25656,
         n25657, n25658, n25659, n25660, n25661, n25662, n25663, n25664,
         n25665, n25666, n25667, n25668, n25669, n25670, n25671, n25672,
         n25673, n25674, n25675, n25676, n25677, n25678, n25679, n25680,
         n25681, n25682, n25683, n25684, n25685, n25686, n25687, n25688,
         n25689, n25690, n25691, n25692, n25693, n25694, n25695, n25696,
         n25697, n25698, n25699, n25700, n25701, n25702, n25703, n25704,
         n25705, n25706, n25707, n25708, n25709, n25710, n25711, n25712,
         n25713, n25714, n25715, n25716, n25717, n25718, n25719, n25720,
         n25721, n25722, n25723, n25724, n25725, n25726, n25727, n25728,
         n25729, n25730, n25731, n25732, n25733, n25734, n25735, n25736,
         n25737, n25738, n25739, n25740, n25741, n25742, n25743, n25744,
         n25745, n25746, n25747, n25748, n25749, n25750, n25751, n25752,
         n25753, n25754, n25755, n25756, n25757, n25758, n25759, n25760,
         n25761, n25762, n25763, n25764, n25765, n25766, n25767, n25768,
         n25769, n25770, n25771, n25772, n25773, n25774, n25775, n25776,
         n25777, n25778, n25779, n25780, n25781, n25782, n25783, n25784,
         n25785, n25786, n25787, n25788, n25789, n25790, n25791, n25792,
         n25793, n25794, n25795, n25796, n25797, n25798, n25799, n25800,
         n25801, n25802, n25803, n25804, n25805, n25806, n25807, n25808,
         n25809, n25810, n25811, n25812, n25813, n25814, n25815, n25816,
         n25817, n25818, n25819, n25820, n25821, n25822, n25823, n25824,
         n25825, n25826, n25827, n25828, n25829, n25830, n25831, n25832,
         n25833, n25834, n25835, n25836, n25837, n25838, n25839, n25840,
         n25841, n25842, n25843, n25844, n25845, n25846, n25847, n25848,
         n25849, n25850, n25851, n25852, n25853, n25854, n25855, n25856,
         n25857, n25858, n25859, n25860, n25861, n25862, n25863, n25864,
         n25865, n25866, n25867, n25868, n25869, n25870, n25871, n25872,
         n25873, n25874, n25875, n25876, n25877, n25878, n25879, n25880,
         n25881, n25882, n25883, n25884, n25885, n25886, n25887, n25888,
         n25889, n25890, n25891, n25892, n25893, n25894, n25895, n25896,
         n25897, n25898, n25899, n25900, n25901, n25902, n25903, n25904,
         n25905, n25906, n25907, n25908, n25909, n25910, n25911, n25912,
         n25913, n25914, n25915, n25916, n25917, n25918, n25919, n25920,
         n25921, n25922, n25923, n25924, n25925, n25926, n25927, n25928,
         n25929, n25930, n25931, n25932, n25933, n25934, n25935, n25936,
         n25937, n25938, n25939, n25940, n25941, n25942, n25943, n25944,
         n25945, n25946, n25947, n25948, n25949, n25950, n25951, n25952,
         n25953, n25954, n25955, n25956, n25957, n25958, n25959, n25960,
         n25961, n25962, n25963, n25964, n25965, n25966, n25967, n25968,
         n25969, n25970, n25971, n25972, n25973, n25974, n25975, n25976,
         n25977, n25978, n25979, n25980, n25981, n25982, n25983, n25984,
         n25985, n25986, n25987, n25988, n25989, n25990, n25991, n25992,
         n25993, n25994, n25995, n25996, n25997, n25998, n25999, n26000,
         n26001, n26002, n26003, n26004, n26005, n26006, n26007, n26008,
         n26009, n26010, n26011, n26012, n26013, n26014, n26015, n26016,
         n26017, n26018, n26019, n26020, n26021, n26022, n26023, n26024,
         n26025, n26026, n26027, n26028, n26029, n26030, n26031, n26032,
         n26033, n26034, n26035, n26036, n26037, n26038, n26039, n26040,
         n26041, n26042, n26043, n26044, n26045, n26046, n26047, n26048,
         n26049, n26050, n26051, n26052, n26053, n26054, n26055, n26056,
         n26057, n26058, n26059, n26060, n26061, n26062, n26063, n26064,
         n26065, n26066, n26067, n26068, n26069, n26070, n26071, n26072,
         n26073, n26074, n26075, n26076, n26077, n26078, n26079, n26080,
         n26081, n26082, n26083, n26084, n26085, n26086, n26087, n26088,
         n26089, n26090, n26091, n26092, n26093, n26094, n26095, n26096,
         n26097, n26098, n26099, n26100, n26101, n26102, n26103, n26104,
         n26105, n26106, n26107, n26108, n26109, n26110, n26111, n26112,
         n26113, n26114, n26115, n26116, n26117, n26118, n26119, n26120,
         n26121, n26122, n26123, n26124, n26125, n26126, n26127, n26128,
         n26129, n26130, n26131, n26132, n26133, n26134, n26135, n26136,
         n26137, n26138, n26139, n26140, n26141, n26142, n26143, n26144,
         n26145, n26146, n26147, n26148, n26149, n26150, n26151, n26152,
         n26153, n26154, n26155, n26156, n26157, n26158, n26159, n26160,
         n26161, n26162, n26163, n26164, n26165, n26166, n26167, n26168,
         n26169, n26170, n26171, n26172, n26173, n26174, n26175, n26176,
         n26177, n26178, n26179, n26180, n26181, n26182, n26183, n26184,
         n26185, n26186, n26187, n26188, n26189, n26190, n26191, n26192,
         n26193, n26194, n26195, n26196, n26197, n26198, n26199, n26200,
         n26201, n26202, n26203, n26204, n26205, n26206, n26207, n26208,
         n26209, n26210, n26211, n26212, n26213, n26214, n26215, n26216,
         n26217, n26218, n26219, n26220, n26221, n26222, n26223, n26224,
         n26225, n26226, n26227, n26228, n26229, n26230, n26231, n26232,
         n26233, n26234, n26235, n26236, n26237, n26238, n26239, n26240,
         n26241, n26242, n26243, n26244, n26245, n26246, n26247, n26248,
         n26249, n26250, n26251, n26252, n26253, n26254, n26255, n26256,
         n26257, n26258, n26259, n26260, n26261, n26262, n26263, n26264,
         n26265, n26266, n26267, n26268, n26269, n26270, n26271, n26272,
         n26273, n26274, n26275, n26276, n26277, n26278, n26279, n26280,
         n26281, n26282, n26283, n26284, n26285, n26286, n26287, n26288,
         n26289, n26290, n26291, n26292, n26293, n26294, n26295, n26296,
         n26297, n26298, n26299, n26300, n26301, n26302, n26303, n26304,
         n26305, n26306, n26307, n26308, n26309, n26310, n26311, n26312,
         n26313, n26314, n26315, n26316, n26317, n26318, n26319, n26320,
         n26321, n26322, n26323, n26324, n26325, n26326, n26327, n26328,
         n26329, n26330, n26331, n26332, n26333, n26334, n26335, n26336,
         n26337, n26338, n26339, n26340, n26341, n26342, n26343, n26344,
         n26345, n26346, n26347, n26348, n26349, n26350, n26351, n26352,
         n26353, n26354, n26355, n26356, n26357, n26358, n26359, n26360,
         n26361, n26362, n26363, n26364, n26365, n26366, n26367, n26368,
         n26369, n26370, n26371, n26372, n26373, n26374, n26375, n26376,
         n26377, n26378, n26379, n26380, n26381, n26382, n26383, n26384,
         n26385, n26386, n26387, n26388, n26389, n26390, n26391, n26392,
         n26393, n26394, n26395, n26396, n26397, n26398, n26399, n26400,
         n26401, n26402, n26403, n26404, n26405, n26406, n26407, n26408,
         n26409, n26410, n26411, n26412, n26413, n26414, n26415, n26416,
         n26417, n26418, n26419, n26420, n26421, n26422, n26423, n26424,
         n26425, n26426, n26427, n26428, n26429, n26430, n26431, n26432,
         n26433, n26434, n26435, n26436, n26437, n26438, n26439, n26440,
         n26441, n26442, n26443, n26444, n26445, n26446, n26447, n26448,
         n26449, n26450, n26451, n26452, n26453, n26454, n26455, n26456,
         n26457, n26458, n26459, n26460, n26461, n26462, n26463, n26464,
         n26465, n26466, n26467, n26468, n26469, n26470, n26471, n26472,
         n26473, n26474, n26475, n26476, n26477, n26478, n26479, n26480,
         n26481, n26482, n26483, n26484, n26485, n26486, n26487, n26488,
         n26489, n26490, n26491, n26492, n26493, n26494, n26495, n26496,
         n26497, n26498, n26499, n26500, n26501, n26502, n26503, n26504,
         n26505, n26506, n26507, n26508, n26509, n26510, n26511, n26512,
         n26513, n26514, n26515, n26516, n26517, n26518, n26519, n26520,
         n26521, n26522, n26523, n26524, n26525, n26526, n26527, n26528,
         n26529, n26530, n26531, n26532, n26533, n26534, n26535, n26536,
         n26537, n26538, n26539, n26540, n26541, n26542, n26543, n26544,
         n26545, n26546, n26547, n26548, n26549, n26550, n26551, n26552,
         n26553, n26554, n26555, n26556, n26557, n26558, n26559, n26560,
         n26561, n26562, n26563, n26564, n26565, n26566, n26567, n26568,
         n26569, n26570, n26571, n26572, n26573, n26574, n26575, n26576,
         n26577, n26578, n26579, n26580, n26581, n26582, n26583, n26584,
         n26585, n26586, n26587, n26588, n26589, n26590, n26591, n26592,
         n26593, n26594, n26595, n26596, n26597, n26598, n26599, n26600,
         n26601, n26602, n26603, n26604, n26605, n26606, n26607, n26608,
         n26609, n26610, n26611, n26612, n26613, n26614, n26615, n26616,
         n26617, n26618, n26619, n26620, n26621, n26622, n26623, n26624,
         n26625, n26626, n26627, n26628, n26629, n26630, n26631, n26632,
         n26633, n26634, n26635, n26636, n26637, n26638, n26639, n26640,
         n26641, n26642, n26643, n26644, n26645, n26646, n26647, n26648,
         n26649, n26650, n26651, n26652, n26653, n26654, n26655, n26656,
         n26657, n26658, n26659, n26660, n26661, n26662, n26663, n26664,
         n26665, n26666, n26667, n26668, n26669, n26670, n26671, n26672,
         n26673, n26674, n26675, n26676, n26677, n26678, n26679, n26680,
         n26681, n26682, n26683, n26684, n26685, n26686, n26687, n26688,
         n26689, n26690, n26691, n26692, n26693, n26694, n26695, n26696,
         n26697, n26698, n26699, n26700, n26701, n26702, n26703, n26704,
         n26705, n26706, n26707, n26708, n26709, n26710, n26711, n26712,
         n26713, n26714, n26715, n26716, n26717, n26718, n26719, n26720,
         n26721, n26722, n26723, n26724, n26725, n26726, n26727, n26728,
         n26729, n26730, n26731, n26732, n26733, n26734, n26735, n26736,
         n26737, n26738, n26739, n26740, n26741, n26742, n26743, n26744,
         n26745, n26746, n26747, n26748, n26749, n26750, n26751, n26752,
         n26753, n26754, n26755, n26756, n26757, n26758, n26759, n26760,
         n26761, n26762, n26763, n26764, n26765, n26766, n26767, n26768,
         n26769, n26770, n26771, n26772, n26773, n26774, n26775, n26776,
         n26777, n26778, n26779, n26780, n26781, n26782, n26783, n26784,
         n26785, n26786, n26787, n26788, n26789, n26790, n26791, n26792,
         n26793, n26794, n26795, n26796, n26797, n26798, n26799, n26800,
         n26801, n26802, n26803, n26804, n26805, n26806, n26807, n26808,
         n26809, n26810, n26811, n26812, n26813, n26814, n26815, n26816,
         n26817, n26818, n26819, n26820, n26821, n26822, n26823, n26824,
         n26825, n26826, n26827, n26828, n26829, n26830, n26831, n26832,
         n26833, n26834, n26835, n26836, n26837, n26838, n26839, n26840,
         n26841, n26842, n26843, n26844, n26845, n26846, n26847, n26848,
         n26849, n26850, n26851, n26852, n26853, n26854, n26855, n26856,
         n26857, n26858, n26859, n26860, n26861, n26862, n26863, n26864,
         n26865, n26866, n26867, n26868, n26869, n26870, n26871, n26872,
         n26873, n26874, n26875, n26876, n26877, n26878, n26879, n26880,
         n26881, n26882, n26883, n26884, n26885, n26886, n26887, n26888,
         n26889, n26890, n26891, n26892, n26893, n26894, n26895, n26896,
         n26897, n26898, n26899, n26900, n26901, n26902, n26903, n26904,
         n26905, n26906, n26907, n26908, n26909, n26910, n26911, n26912,
         n26913, n26914, n26915, n26916, n26917, n26918, n26919, n26920,
         n26921, n26922, n26923, n26924, n26925, n26926, n26927, n26928,
         n26929, n26930, n26931, n26932, n26933, n26934, n26935, n26936,
         n26937, n26938, n26939, n26940, n26941, n26942, n26943, n26944,
         n26945, n26946, n26947, n26948, n26949, n26950, n26951, n26952,
         n26953, n26954, n26955, n26956, n26957, n26958, n26959, n26960,
         n26961, n26962, n26963, n26964, n26965, n26966, n26967, n26968,
         n26969, n26970, n26971, n26972, n26973, n26974, n26975, n26976,
         n26977, n26978, n26979, n26980, n26981, n26982, n26983, n26984,
         n26985, n26986, n26987, n26988, n26989, n26990, n26991, n26992,
         n26993, n26994, n26995, n26996, n26997, n26998, n26999, n27000,
         n27001, n27002, n27003, n27004, n27005, n27006, n27007, n27008,
         n27009, n27010, n27011, n27012, n27013, n27014, n27015, n27016,
         n27017, n27018, n27019, n27020, n27021, n27022, n27023, n27024,
         n27025, n27026, n27027, n27028, n27029, n27030, n27031, n27032,
         n27033, n27034, n27035, n27036, n27037, n27038, n27039, n27040,
         n27041, n27042, n27043, n27044, n27045, n27046, n27047, n27048,
         n27049, n27050, n27051, n27052, n27053, n27054, n27055, n27056,
         n27057, n27058, n27059, n27060, n27061, n27062, n27063, n27064,
         n27065, n27066, n27067, n27068, n27069, n27070, n27071, n27072,
         n27073, n27074, n27075, n27076, n27077, n27078, n27079, n27080,
         n27081, n27082, n27083, n27084, n27085, n27086, n27087, n27088,
         n27089, n27090, n27091, n27092, n27093, n27094, n27095, n27096,
         n27097, n27098, n27099, n27100, n27101, n27102, n27103, n27104,
         n27105, n27106, n27107, n27108, n27109, n27110, n27111, n27112,
         n27113, n27114, n27115, n27116, n27117, n27118, n27119, n27120,
         n27121, n27122, n27123, n27124, n27125, n27126, n27127, n27128,
         n27129, n27130, n27131, n27132, n27133, n27134, n27135, n27136,
         n27137, n27138, n27139, n27140, n27141, n27142, n27143, n27144,
         n27145, n27146, n27147, n27148, n27149, n27150, n27151, n27152,
         n27153, n27154, n27155, n27156, n27157, n27158, n27159, n27160,
         n27161, n27162, n27163, n27164, n27165, n27166, n27167, n27168,
         n27169, n27170, n27171, n27172, n27173;
  wire   [11:0] olocal;
  wire   [13:0] oglobal;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154, SYNOPSYS_UNCONNECTED__155, 
        SYNOPSYS_UNCONNECTED__156, SYNOPSYS_UNCONNECTED__157, 
        SYNOPSYS_UNCONNECTED__158, SYNOPSYS_UNCONNECTED__159, 
        SYNOPSYS_UNCONNECTED__160, SYNOPSYS_UNCONNECTED__161, 
        SYNOPSYS_UNCONNECTED__162, SYNOPSYS_UNCONNECTED__163, 
        SYNOPSYS_UNCONNECTED__164, SYNOPSYS_UNCONNECTED__165, 
        SYNOPSYS_UNCONNECTED__166, SYNOPSYS_UNCONNECTED__167, 
        SYNOPSYS_UNCONNECTED__168, SYNOPSYS_UNCONNECTED__169, 
        SYNOPSYS_UNCONNECTED__170, SYNOPSYS_UNCONNECTED__171, 
        SYNOPSYS_UNCONNECTED__172, SYNOPSYS_UNCONNECTED__173, 
        SYNOPSYS_UNCONNECTED__174, SYNOPSYS_UNCONNECTED__175, 
        SYNOPSYS_UNCONNECTED__176, SYNOPSYS_UNCONNECTED__177, 
        SYNOPSYS_UNCONNECTED__178, SYNOPSYS_UNCONNECTED__179, 
        SYNOPSYS_UNCONNECTED__180, SYNOPSYS_UNCONNECTED__181, 
        SYNOPSYS_UNCONNECTED__182, SYNOPSYS_UNCONNECTED__183, 
        SYNOPSYS_UNCONNECTED__184, SYNOPSYS_UNCONNECTED__185, 
        SYNOPSYS_UNCONNECTED__186, SYNOPSYS_UNCONNECTED__187, 
        SYNOPSYS_UNCONNECTED__188, SYNOPSYS_UNCONNECTED__189, 
        SYNOPSYS_UNCONNECTED__190, SYNOPSYS_UNCONNECTED__191, 
        SYNOPSYS_UNCONNECTED__192, SYNOPSYS_UNCONNECTED__193, 
        SYNOPSYS_UNCONNECTED__194, SYNOPSYS_UNCONNECTED__195, 
        SYNOPSYS_UNCONNECTED__196, SYNOPSYS_UNCONNECTED__197, 
        SYNOPSYS_UNCONNECTED__198, SYNOPSYS_UNCONNECTED__199, 
        SYNOPSYS_UNCONNECTED__200, SYNOPSYS_UNCONNECTED__201, 
        SYNOPSYS_UNCONNECTED__202, SYNOPSYS_UNCONNECTED__203, 
        SYNOPSYS_UNCONNECTED__204, SYNOPSYS_UNCONNECTED__205, 
        SYNOPSYS_UNCONNECTED__206, SYNOPSYS_UNCONNECTED__207, 
        SYNOPSYS_UNCONNECTED__208, SYNOPSYS_UNCONNECTED__209, 
        SYNOPSYS_UNCONNECTED__210, SYNOPSYS_UNCONNECTED__211, 
        SYNOPSYS_UNCONNECTED__212, SYNOPSYS_UNCONNECTED__213, 
        SYNOPSYS_UNCONNECTED__214, SYNOPSYS_UNCONNECTED__215, 
        SYNOPSYS_UNCONNECTED__216, SYNOPSYS_UNCONNECTED__217, 
        SYNOPSYS_UNCONNECTED__218, SYNOPSYS_UNCONNECTED__219, 
        SYNOPSYS_UNCONNECTED__220, SYNOPSYS_UNCONNECTED__221, 
        SYNOPSYS_UNCONNECTED__222, SYNOPSYS_UNCONNECTED__223, 
        SYNOPSYS_UNCONNECTED__224, SYNOPSYS_UNCONNECTED__225, 
        SYNOPSYS_UNCONNECTED__226, SYNOPSYS_UNCONNECTED__227, 
        SYNOPSYS_UNCONNECTED__228, SYNOPSYS_UNCONNECTED__229, 
        SYNOPSYS_UNCONNECTED__230, SYNOPSYS_UNCONNECTED__231, 
        SYNOPSYS_UNCONNECTED__232, SYNOPSYS_UNCONNECTED__233, 
        SYNOPSYS_UNCONNECTED__234, SYNOPSYS_UNCONNECTED__235, 
        SYNOPSYS_UNCONNECTED__236, SYNOPSYS_UNCONNECTED__237, 
        SYNOPSYS_UNCONNECTED__238, SYNOPSYS_UNCONNECTED__239, 
        SYNOPSYS_UNCONNECTED__240, SYNOPSYS_UNCONNECTED__241, 
        SYNOPSYS_UNCONNECTED__242, SYNOPSYS_UNCONNECTED__243, 
        SYNOPSYS_UNCONNECTED__244, SYNOPSYS_UNCONNECTED__245, 
        SYNOPSYS_UNCONNECTED__246, SYNOPSYS_UNCONNECTED__247, 
        SYNOPSYS_UNCONNECTED__248, SYNOPSYS_UNCONNECTED__249, 
        SYNOPSYS_UNCONNECTED__250, SYNOPSYS_UNCONNECTED__251, 
        SYNOPSYS_UNCONNECTED__252, SYNOPSYS_UNCONNECTED__253, 
        SYNOPSYS_UNCONNECTED__254, SYNOPSYS_UNCONNECTED__255, 
        SYNOPSYS_UNCONNECTED__256, SYNOPSYS_UNCONNECTED__257, 
        SYNOPSYS_UNCONNECTED__258, SYNOPSYS_UNCONNECTED__259, 
        SYNOPSYS_UNCONNECTED__260, SYNOPSYS_UNCONNECTED__261, 
        SYNOPSYS_UNCONNECTED__262, SYNOPSYS_UNCONNECTED__263, 
        SYNOPSYS_UNCONNECTED__264, SYNOPSYS_UNCONNECTED__265, 
        SYNOPSYS_UNCONNECTED__266, SYNOPSYS_UNCONNECTED__267, 
        SYNOPSYS_UNCONNECTED__268, SYNOPSYS_UNCONNECTED__269, 
        SYNOPSYS_UNCONNECTED__270, SYNOPSYS_UNCONNECTED__271, 
        SYNOPSYS_UNCONNECTED__272, SYNOPSYS_UNCONNECTED__273, 
        SYNOPSYS_UNCONNECTED__274, SYNOPSYS_UNCONNECTED__275, 
        SYNOPSYS_UNCONNECTED__276, SYNOPSYS_UNCONNECTED__277, 
        SYNOPSYS_UNCONNECTED__278, SYNOPSYS_UNCONNECTED__279, 
        SYNOPSYS_UNCONNECTED__280, SYNOPSYS_UNCONNECTED__281, 
        SYNOPSYS_UNCONNECTED__282, SYNOPSYS_UNCONNECTED__283, 
        SYNOPSYS_UNCONNECTED__284, SYNOPSYS_UNCONNECTED__285, 
        SYNOPSYS_UNCONNECTED__286, SYNOPSYS_UNCONNECTED__287, 
        SYNOPSYS_UNCONNECTED__288, SYNOPSYS_UNCONNECTED__289, 
        SYNOPSYS_UNCONNECTED__290, SYNOPSYS_UNCONNECTED__291, 
        SYNOPSYS_UNCONNECTED__292, SYNOPSYS_UNCONNECTED__293, 
        SYNOPSYS_UNCONNECTED__294, SYNOPSYS_UNCONNECTED__295, 
        SYNOPSYS_UNCONNECTED__296, SYNOPSYS_UNCONNECTED__297, 
        SYNOPSYS_UNCONNECTED__298, SYNOPSYS_UNCONNECTED__299, 
        SYNOPSYS_UNCONNECTED__300, SYNOPSYS_UNCONNECTED__301, 
        SYNOPSYS_UNCONNECTED__302, SYNOPSYS_UNCONNECTED__303, 
        SYNOPSYS_UNCONNECTED__304, SYNOPSYS_UNCONNECTED__305, 
        SYNOPSYS_UNCONNECTED__306, SYNOPSYS_UNCONNECTED__307, 
        SYNOPSYS_UNCONNECTED__308, SYNOPSYS_UNCONNECTED__309, 
        SYNOPSYS_UNCONNECTED__310, SYNOPSYS_UNCONNECTED__311, 
        SYNOPSYS_UNCONNECTED__312, SYNOPSYS_UNCONNECTED__313, 
        SYNOPSYS_UNCONNECTED__314, SYNOPSYS_UNCONNECTED__315, 
        SYNOPSYS_UNCONNECTED__316, SYNOPSYS_UNCONNECTED__317, 
        SYNOPSYS_UNCONNECTED__318, SYNOPSYS_UNCONNECTED__319, 
        SYNOPSYS_UNCONNECTED__320, SYNOPSYS_UNCONNECTED__321, 
        SYNOPSYS_UNCONNECTED__322, SYNOPSYS_UNCONNECTED__323, 
        SYNOPSYS_UNCONNECTED__324, SYNOPSYS_UNCONNECTED__325, 
        SYNOPSYS_UNCONNECTED__326, SYNOPSYS_UNCONNECTED__327, 
        SYNOPSYS_UNCONNECTED__328, SYNOPSYS_UNCONNECTED__329, 
        SYNOPSYS_UNCONNECTED__330, SYNOPSYS_UNCONNECTED__331, 
        SYNOPSYS_UNCONNECTED__332, SYNOPSYS_UNCONNECTED__333, 
        SYNOPSYS_UNCONNECTED__334, SYNOPSYS_UNCONNECTED__335, 
        SYNOPSYS_UNCONNECTED__336, SYNOPSYS_UNCONNECTED__337, 
        SYNOPSYS_UNCONNECTED__338, SYNOPSYS_UNCONNECTED__339, 
        SYNOPSYS_UNCONNECTED__340, SYNOPSYS_UNCONNECTED__341, 
        SYNOPSYS_UNCONNECTED__342, SYNOPSYS_UNCONNECTED__343, 
        SYNOPSYS_UNCONNECTED__344, SYNOPSYS_UNCONNECTED__345, 
        SYNOPSYS_UNCONNECTED__346, SYNOPSYS_UNCONNECTED__347, 
        SYNOPSYS_UNCONNECTED__348, SYNOPSYS_UNCONNECTED__349, 
        SYNOPSYS_UNCONNECTED__350, SYNOPSYS_UNCONNECTED__351, 
        SYNOPSYS_UNCONNECTED__352, SYNOPSYS_UNCONNECTED__353, 
        SYNOPSYS_UNCONNECTED__354, SYNOPSYS_UNCONNECTED__355, 
        SYNOPSYS_UNCONNECTED__356, SYNOPSYS_UNCONNECTED__357, 
        SYNOPSYS_UNCONNECTED__358, SYNOPSYS_UNCONNECTED__359, 
        SYNOPSYS_UNCONNECTED__360, SYNOPSYS_UNCONNECTED__361, 
        SYNOPSYS_UNCONNECTED__362, SYNOPSYS_UNCONNECTED__363, 
        SYNOPSYS_UNCONNECTED__364, SYNOPSYS_UNCONNECTED__365, 
        SYNOPSYS_UNCONNECTED__366, SYNOPSYS_UNCONNECTED__367, 
        SYNOPSYS_UNCONNECTED__368, SYNOPSYS_UNCONNECTED__369, 
        SYNOPSYS_UNCONNECTED__370, SYNOPSYS_UNCONNECTED__371, 
        SYNOPSYS_UNCONNECTED__372, SYNOPSYS_UNCONNECTED__373, 
        SYNOPSYS_UNCONNECTED__374, SYNOPSYS_UNCONNECTED__375, 
        SYNOPSYS_UNCONNECTED__376, SYNOPSYS_UNCONNECTED__377, 
        SYNOPSYS_UNCONNECTED__378, SYNOPSYS_UNCONNECTED__379, 
        SYNOPSYS_UNCONNECTED__380, SYNOPSYS_UNCONNECTED__381, 
        SYNOPSYS_UNCONNECTED__382, SYNOPSYS_UNCONNECTED__383, 
        SYNOPSYS_UNCONNECTED__384, SYNOPSYS_UNCONNECTED__385, 
        SYNOPSYS_UNCONNECTED__386, SYNOPSYS_UNCONNECTED__387, 
        SYNOPSYS_UNCONNECTED__388, SYNOPSYS_UNCONNECTED__389, 
        SYNOPSYS_UNCONNECTED__390, SYNOPSYS_UNCONNECTED__391, 
        SYNOPSYS_UNCONNECTED__392, SYNOPSYS_UNCONNECTED__393, 
        SYNOPSYS_UNCONNECTED__394, SYNOPSYS_UNCONNECTED__395, 
        SYNOPSYS_UNCONNECTED__396, SYNOPSYS_UNCONNECTED__397, 
        SYNOPSYS_UNCONNECTED__398, SYNOPSYS_UNCONNECTED__399, 
        SYNOPSYS_UNCONNECTED__400, SYNOPSYS_UNCONNECTED__401, 
        SYNOPSYS_UNCONNECTED__402, SYNOPSYS_UNCONNECTED__403, 
        SYNOPSYS_UNCONNECTED__404, SYNOPSYS_UNCONNECTED__405, 
        SYNOPSYS_UNCONNECTED__406, SYNOPSYS_UNCONNECTED__407, 
        SYNOPSYS_UNCONNECTED__408, SYNOPSYS_UNCONNECTED__409, 
        SYNOPSYS_UNCONNECTED__410, SYNOPSYS_UNCONNECTED__411, 
        SYNOPSYS_UNCONNECTED__412, SYNOPSYS_UNCONNECTED__413, 
        SYNOPSYS_UNCONNECTED__414, SYNOPSYS_UNCONNECTED__415, 
        SYNOPSYS_UNCONNECTED__416, SYNOPSYS_UNCONNECTED__417, 
        SYNOPSYS_UNCONNECTED__418, SYNOPSYS_UNCONNECTED__419, 
        SYNOPSYS_UNCONNECTED__420, SYNOPSYS_UNCONNECTED__421, 
        SYNOPSYS_UNCONNECTED__422, SYNOPSYS_UNCONNECTED__423, 
        SYNOPSYS_UNCONNECTED__424, SYNOPSYS_UNCONNECTED__425, 
        SYNOPSYS_UNCONNECTED__426, SYNOPSYS_UNCONNECTED__427, 
        SYNOPSYS_UNCONNECTED__428, SYNOPSYS_UNCONNECTED__429, 
        SYNOPSYS_UNCONNECTED__430, SYNOPSYS_UNCONNECTED__431, 
        SYNOPSYS_UNCONNECTED__432, SYNOPSYS_UNCONNECTED__433, 
        SYNOPSYS_UNCONNECTED__434, SYNOPSYS_UNCONNECTED__435, 
        SYNOPSYS_UNCONNECTED__436, SYNOPSYS_UNCONNECTED__437, 
        SYNOPSYS_UNCONNECTED__438, SYNOPSYS_UNCONNECTED__439, 
        SYNOPSYS_UNCONNECTED__440, SYNOPSYS_UNCONNECTED__441, 
        SYNOPSYS_UNCONNECTED__442, SYNOPSYS_UNCONNECTED__443, 
        SYNOPSYS_UNCONNECTED__444, SYNOPSYS_UNCONNECTED__445, 
        SYNOPSYS_UNCONNECTED__446, SYNOPSYS_UNCONNECTED__447, 
        SYNOPSYS_UNCONNECTED__448, SYNOPSYS_UNCONNECTED__449, 
        SYNOPSYS_UNCONNECTED__450, SYNOPSYS_UNCONNECTED__451, 
        SYNOPSYS_UNCONNECTED__452, SYNOPSYS_UNCONNECTED__453, 
        SYNOPSYS_UNCONNECTED__454, SYNOPSYS_UNCONNECTED__455, 
        SYNOPSYS_UNCONNECTED__456, SYNOPSYS_UNCONNECTED__457, 
        SYNOPSYS_UNCONNECTED__458, SYNOPSYS_UNCONNECTED__459, 
        SYNOPSYS_UNCONNECTED__460, SYNOPSYS_UNCONNECTED__461, 
        SYNOPSYS_UNCONNECTED__462, SYNOPSYS_UNCONNECTED__463, 
        SYNOPSYS_UNCONNECTED__464, SYNOPSYS_UNCONNECTED__465, 
        SYNOPSYS_UNCONNECTED__466, SYNOPSYS_UNCONNECTED__467, 
        SYNOPSYS_UNCONNECTED__468, SYNOPSYS_UNCONNECTED__469, 
        SYNOPSYS_UNCONNECTED__470, SYNOPSYS_UNCONNECTED__471, 
        SYNOPSYS_UNCONNECTED__472, SYNOPSYS_UNCONNECTED__473, 
        SYNOPSYS_UNCONNECTED__474, SYNOPSYS_UNCONNECTED__475, 
        SYNOPSYS_UNCONNECTED__476, SYNOPSYS_UNCONNECTED__477, 
        SYNOPSYS_UNCONNECTED__478, SYNOPSYS_UNCONNECTED__479, 
        SYNOPSYS_UNCONNECTED__480, SYNOPSYS_UNCONNECTED__481, 
        SYNOPSYS_UNCONNECTED__482, SYNOPSYS_UNCONNECTED__483, 
        SYNOPSYS_UNCONNECTED__484, SYNOPSYS_UNCONNECTED__485, 
        SYNOPSYS_UNCONNECTED__486, SYNOPSYS_UNCONNECTED__487, 
        SYNOPSYS_UNCONNECTED__488, SYNOPSYS_UNCONNECTED__489, 
        SYNOPSYS_UNCONNECTED__490, SYNOPSYS_UNCONNECTED__491, 
        SYNOPSYS_UNCONNECTED__492, SYNOPSYS_UNCONNECTED__493, 
        SYNOPSYS_UNCONNECTED__494, SYNOPSYS_UNCONNECTED__495, 
        SYNOPSYS_UNCONNECTED__496, SYNOPSYS_UNCONNECTED__497, 
        SYNOPSYS_UNCONNECTED__498, SYNOPSYS_UNCONNECTED__499, 
        SYNOPSYS_UNCONNECTED__500, SYNOPSYS_UNCONNECTED__501, 
        SYNOPSYS_UNCONNECTED__502, SYNOPSYS_UNCONNECTED__503, 
        SYNOPSYS_UNCONNECTED__504, SYNOPSYS_UNCONNECTED__505, 
        SYNOPSYS_UNCONNECTED__506, SYNOPSYS_UNCONNECTED__507, 
        SYNOPSYS_UNCONNECTED__508, SYNOPSYS_UNCONNECTED__509, 
        SYNOPSYS_UNCONNECTED__510, SYNOPSYS_UNCONNECTED__511, 
        SYNOPSYS_UNCONNECTED__512, SYNOPSYS_UNCONNECTED__513, 
        SYNOPSYS_UNCONNECTED__514, SYNOPSYS_UNCONNECTED__515, 
        SYNOPSYS_UNCONNECTED__516, SYNOPSYS_UNCONNECTED__517, 
        SYNOPSYS_UNCONNECTED__518, SYNOPSYS_UNCONNECTED__519, 
        SYNOPSYS_UNCONNECTED__520, SYNOPSYS_UNCONNECTED__521, 
        SYNOPSYS_UNCONNECTED__522, SYNOPSYS_UNCONNECTED__523, 
        SYNOPSYS_UNCONNECTED__524, SYNOPSYS_UNCONNECTED__525, 
        SYNOPSYS_UNCONNECTED__526, SYNOPSYS_UNCONNECTED__527, 
        SYNOPSYS_UNCONNECTED__528, SYNOPSYS_UNCONNECTED__529, 
        SYNOPSYS_UNCONNECTED__530, SYNOPSYS_UNCONNECTED__531, 
        SYNOPSYS_UNCONNECTED__532, SYNOPSYS_UNCONNECTED__533, 
        SYNOPSYS_UNCONNECTED__534, SYNOPSYS_UNCONNECTED__535, 
        SYNOPSYS_UNCONNECTED__536, SYNOPSYS_UNCONNECTED__537, 
        SYNOPSYS_UNCONNECTED__538, SYNOPSYS_UNCONNECTED__539, 
        SYNOPSYS_UNCONNECTED__540, SYNOPSYS_UNCONNECTED__541, 
        SYNOPSYS_UNCONNECTED__542, SYNOPSYS_UNCONNECTED__543, 
        SYNOPSYS_UNCONNECTED__544, SYNOPSYS_UNCONNECTED__545, 
        SYNOPSYS_UNCONNECTED__546, SYNOPSYS_UNCONNECTED__547, 
        SYNOPSYS_UNCONNECTED__548, SYNOPSYS_UNCONNECTED__549, 
        SYNOPSYS_UNCONNECTED__550, SYNOPSYS_UNCONNECTED__551, 
        SYNOPSYS_UNCONNECTED__552, SYNOPSYS_UNCONNECTED__553, 
        SYNOPSYS_UNCONNECTED__554, SYNOPSYS_UNCONNECTED__555, 
        SYNOPSYS_UNCONNECTED__556, SYNOPSYS_UNCONNECTED__557, 
        SYNOPSYS_UNCONNECTED__558, SYNOPSYS_UNCONNECTED__559, 
        SYNOPSYS_UNCONNECTED__560, SYNOPSYS_UNCONNECTED__561, 
        SYNOPSYS_UNCONNECTED__562, SYNOPSYS_UNCONNECTED__563, 
        SYNOPSYS_UNCONNECTED__564, SYNOPSYS_UNCONNECTED__565, 
        SYNOPSYS_UNCONNECTED__566, SYNOPSYS_UNCONNECTED__567, 
        SYNOPSYS_UNCONNECTED__568, SYNOPSYS_UNCONNECTED__569, 
        SYNOPSYS_UNCONNECTED__570, SYNOPSYS_UNCONNECTED__571, 
        SYNOPSYS_UNCONNECTED__572, SYNOPSYS_UNCONNECTED__573, 
        SYNOPSYS_UNCONNECTED__574, SYNOPSYS_UNCONNECTED__575, 
        SYNOPSYS_UNCONNECTED__576, SYNOPSYS_UNCONNECTED__577, 
        SYNOPSYS_UNCONNECTED__578, SYNOPSYS_UNCONNECTED__579, 
        SYNOPSYS_UNCONNECTED__580, SYNOPSYS_UNCONNECTED__581, 
        SYNOPSYS_UNCONNECTED__582, SYNOPSYS_UNCONNECTED__583, 
        SYNOPSYS_UNCONNECTED__584, SYNOPSYS_UNCONNECTED__585, 
        SYNOPSYS_UNCONNECTED__586, SYNOPSYS_UNCONNECTED__587, 
        SYNOPSYS_UNCONNECTED__588, SYNOPSYS_UNCONNECTED__589, 
        SYNOPSYS_UNCONNECTED__590, SYNOPSYS_UNCONNECTED__591, 
        SYNOPSYS_UNCONNECTED__592, SYNOPSYS_UNCONNECTED__593, 
        SYNOPSYS_UNCONNECTED__594, SYNOPSYS_UNCONNECTED__595, 
        SYNOPSYS_UNCONNECTED__596, SYNOPSYS_UNCONNECTED__597, 
        SYNOPSYS_UNCONNECTED__598, SYNOPSYS_UNCONNECTED__599, 
        SYNOPSYS_UNCONNECTED__600, SYNOPSYS_UNCONNECTED__601, 
        SYNOPSYS_UNCONNECTED__602, SYNOPSYS_UNCONNECTED__603, 
        SYNOPSYS_UNCONNECTED__604, SYNOPSYS_UNCONNECTED__605, 
        SYNOPSYS_UNCONNECTED__606, SYNOPSYS_UNCONNECTED__607, 
        SYNOPSYS_UNCONNECTED__608, SYNOPSYS_UNCONNECTED__609, 
        SYNOPSYS_UNCONNECTED__610, SYNOPSYS_UNCONNECTED__611, 
        SYNOPSYS_UNCONNECTED__612, SYNOPSYS_UNCONNECTED__613, 
        SYNOPSYS_UNCONNECTED__614, SYNOPSYS_UNCONNECTED__615, 
        SYNOPSYS_UNCONNECTED__616, SYNOPSYS_UNCONNECTED__617, 
        SYNOPSYS_UNCONNECTED__618, SYNOPSYS_UNCONNECTED__619, 
        SYNOPSYS_UNCONNECTED__620, SYNOPSYS_UNCONNECTED__621, 
        SYNOPSYS_UNCONNECTED__622, SYNOPSYS_UNCONNECTED__623, 
        SYNOPSYS_UNCONNECTED__624, SYNOPSYS_UNCONNECTED__625, 
        SYNOPSYS_UNCONNECTED__626, SYNOPSYS_UNCONNECTED__627, 
        SYNOPSYS_UNCONNECTED__628, SYNOPSYS_UNCONNECTED__629, 
        SYNOPSYS_UNCONNECTED__630, SYNOPSYS_UNCONNECTED__631, 
        SYNOPSYS_UNCONNECTED__632, SYNOPSYS_UNCONNECTED__633, 
        SYNOPSYS_UNCONNECTED__634, SYNOPSYS_UNCONNECTED__635, 
        SYNOPSYS_UNCONNECTED__636, SYNOPSYS_UNCONNECTED__637, 
        SYNOPSYS_UNCONNECTED__638, SYNOPSYS_UNCONNECTED__639, 
        SYNOPSYS_UNCONNECTED__640, SYNOPSYS_UNCONNECTED__641, 
        SYNOPSYS_UNCONNECTED__642, SYNOPSYS_UNCONNECTED__643, 
        SYNOPSYS_UNCONNECTED__644, SYNOPSYS_UNCONNECTED__645, 
        SYNOPSYS_UNCONNECTED__646, SYNOPSYS_UNCONNECTED__647, 
        SYNOPSYS_UNCONNECTED__648, SYNOPSYS_UNCONNECTED__649, 
        SYNOPSYS_UNCONNECTED__650, SYNOPSYS_UNCONNECTED__651, 
        SYNOPSYS_UNCONNECTED__652, SYNOPSYS_UNCONNECTED__653, 
        SYNOPSYS_UNCONNECTED__654, SYNOPSYS_UNCONNECTED__655, 
        SYNOPSYS_UNCONNECTED__656, SYNOPSYS_UNCONNECTED__657, 
        SYNOPSYS_UNCONNECTED__658, SYNOPSYS_UNCONNECTED__659, 
        SYNOPSYS_UNCONNECTED__660, SYNOPSYS_UNCONNECTED__661, 
        SYNOPSYS_UNCONNECTED__662, SYNOPSYS_UNCONNECTED__663, 
        SYNOPSYS_UNCONNECTED__664, SYNOPSYS_UNCONNECTED__665, 
        SYNOPSYS_UNCONNECTED__666, SYNOPSYS_UNCONNECTED__667, 
        SYNOPSYS_UNCONNECTED__668, SYNOPSYS_UNCONNECTED__669, 
        SYNOPSYS_UNCONNECTED__670, SYNOPSYS_UNCONNECTED__671, 
        SYNOPSYS_UNCONNECTED__672, SYNOPSYS_UNCONNECTED__673, 
        SYNOPSYS_UNCONNECTED__674, SYNOPSYS_UNCONNECTED__675, 
        SYNOPSYS_UNCONNECTED__676, SYNOPSYS_UNCONNECTED__677, 
        SYNOPSYS_UNCONNECTED__678, SYNOPSYS_UNCONNECTED__679, 
        SYNOPSYS_UNCONNECTED__680, SYNOPSYS_UNCONNECTED__681, 
        SYNOPSYS_UNCONNECTED__682, SYNOPSYS_UNCONNECTED__683, 
        SYNOPSYS_UNCONNECTED__684, SYNOPSYS_UNCONNECTED__685, 
        SYNOPSYS_UNCONNECTED__686, SYNOPSYS_UNCONNECTED__687, 
        SYNOPSYS_UNCONNECTED__688, SYNOPSYS_UNCONNECTED__689, 
        SYNOPSYS_UNCONNECTED__690, SYNOPSYS_UNCONNECTED__691, 
        SYNOPSYS_UNCONNECTED__692, SYNOPSYS_UNCONNECTED__693, 
        SYNOPSYS_UNCONNECTED__694, SYNOPSYS_UNCONNECTED__695, 
        SYNOPSYS_UNCONNECTED__696, SYNOPSYS_UNCONNECTED__697, 
        SYNOPSYS_UNCONNECTED__698, SYNOPSYS_UNCONNECTED__699, 
        SYNOPSYS_UNCONNECTED__700, SYNOPSYS_UNCONNECTED__701, 
        SYNOPSYS_UNCONNECTED__702, SYNOPSYS_UNCONNECTED__703, 
        SYNOPSYS_UNCONNECTED__704, SYNOPSYS_UNCONNECTED__705, 
        SYNOPSYS_UNCONNECTED__706, SYNOPSYS_UNCONNECTED__707, 
        SYNOPSYS_UNCONNECTED__708, SYNOPSYS_UNCONNECTED__709, 
        SYNOPSYS_UNCONNECTED__710, SYNOPSYS_UNCONNECTED__711, 
        SYNOPSYS_UNCONNECTED__712, SYNOPSYS_UNCONNECTED__713, 
        SYNOPSYS_UNCONNECTED__714, SYNOPSYS_UNCONNECTED__715, 
        SYNOPSYS_UNCONNECTED__716, SYNOPSYS_UNCONNECTED__717, 
        SYNOPSYS_UNCONNECTED__718, SYNOPSYS_UNCONNECTED__719, 
        SYNOPSYS_UNCONNECTED__720, SYNOPSYS_UNCONNECTED__721, 
        SYNOPSYS_UNCONNECTED__722, SYNOPSYS_UNCONNECTED__723, 
        SYNOPSYS_UNCONNECTED__724, SYNOPSYS_UNCONNECTED__725, 
        SYNOPSYS_UNCONNECTED__726, SYNOPSYS_UNCONNECTED__727, 
        SYNOPSYS_UNCONNECTED__728, SYNOPSYS_UNCONNECTED__729, 
        SYNOPSYS_UNCONNECTED__730, SYNOPSYS_UNCONNECTED__731, 
        SYNOPSYS_UNCONNECTED__732, SYNOPSYS_UNCONNECTED__733, 
        SYNOPSYS_UNCONNECTED__734, SYNOPSYS_UNCONNECTED__735, 
        SYNOPSYS_UNCONNECTED__736, SYNOPSYS_UNCONNECTED__737, 
        SYNOPSYS_UNCONNECTED__738, SYNOPSYS_UNCONNECTED__739, 
        SYNOPSYS_UNCONNECTED__740, SYNOPSYS_UNCONNECTED__741, 
        SYNOPSYS_UNCONNECTED__742, SYNOPSYS_UNCONNECTED__743, 
        SYNOPSYS_UNCONNECTED__744, SYNOPSYS_UNCONNECTED__745, 
        SYNOPSYS_UNCONNECTED__746, SYNOPSYS_UNCONNECTED__747, 
        SYNOPSYS_UNCONNECTED__748, SYNOPSYS_UNCONNECTED__749, 
        SYNOPSYS_UNCONNECTED__750, SYNOPSYS_UNCONNECTED__751, 
        SYNOPSYS_UNCONNECTED__752, SYNOPSYS_UNCONNECTED__753, 
        SYNOPSYS_UNCONNECTED__754, SYNOPSYS_UNCONNECTED__755, 
        SYNOPSYS_UNCONNECTED__756, SYNOPSYS_UNCONNECTED__757, 
        SYNOPSYS_UNCONNECTED__758, SYNOPSYS_UNCONNECTED__759, 
        SYNOPSYS_UNCONNECTED__760, SYNOPSYS_UNCONNECTED__761, 
        SYNOPSYS_UNCONNECTED__762, SYNOPSYS_UNCONNECTED__763, 
        SYNOPSYS_UNCONNECTED__764, SYNOPSYS_UNCONNECTED__765, 
        SYNOPSYS_UNCONNECTED__766, SYNOPSYS_UNCONNECTED__767, 
        SYNOPSYS_UNCONNECTED__768, SYNOPSYS_UNCONNECTED__769, 
        SYNOPSYS_UNCONNECTED__770, SYNOPSYS_UNCONNECTED__771, 
        SYNOPSYS_UNCONNECTED__772, SYNOPSYS_UNCONNECTED__773, 
        SYNOPSYS_UNCONNECTED__774, SYNOPSYS_UNCONNECTED__775, 
        SYNOPSYS_UNCONNECTED__776, SYNOPSYS_UNCONNECTED__777, 
        SYNOPSYS_UNCONNECTED__778, SYNOPSYS_UNCONNECTED__779, 
        SYNOPSYS_UNCONNECTED__780, SYNOPSYS_UNCONNECTED__781, 
        SYNOPSYS_UNCONNECTED__782, SYNOPSYS_UNCONNECTED__783, 
        SYNOPSYS_UNCONNECTED__784, SYNOPSYS_UNCONNECTED__785, 
        SYNOPSYS_UNCONNECTED__786, SYNOPSYS_UNCONNECTED__787, 
        SYNOPSYS_UNCONNECTED__788, SYNOPSYS_UNCONNECTED__789, 
        SYNOPSYS_UNCONNECTED__790, SYNOPSYS_UNCONNECTED__791, 
        SYNOPSYS_UNCONNECTED__792, SYNOPSYS_UNCONNECTED__793, 
        SYNOPSYS_UNCONNECTED__794, SYNOPSYS_UNCONNECTED__795, 
        SYNOPSYS_UNCONNECTED__796, SYNOPSYS_UNCONNECTED__797, 
        SYNOPSYS_UNCONNECTED__798, SYNOPSYS_UNCONNECTED__799, 
        SYNOPSYS_UNCONNECTED__800, SYNOPSYS_UNCONNECTED__801, 
        SYNOPSYS_UNCONNECTED__802, SYNOPSYS_UNCONNECTED__803, 
        SYNOPSYS_UNCONNECTED__804, SYNOPSYS_UNCONNECTED__805, 
        SYNOPSYS_UNCONNECTED__806, SYNOPSYS_UNCONNECTED__807, 
        SYNOPSYS_UNCONNECTED__808, SYNOPSYS_UNCONNECTED__809, 
        SYNOPSYS_UNCONNECTED__810, SYNOPSYS_UNCONNECTED__811, 
        SYNOPSYS_UNCONNECTED__812, SYNOPSYS_UNCONNECTED__813, 
        SYNOPSYS_UNCONNECTED__814, SYNOPSYS_UNCONNECTED__815, 
        SYNOPSYS_UNCONNECTED__816, SYNOPSYS_UNCONNECTED__817, 
        SYNOPSYS_UNCONNECTED__818, SYNOPSYS_UNCONNECTED__819, 
        SYNOPSYS_UNCONNECTED__820, SYNOPSYS_UNCONNECTED__821, 
        SYNOPSYS_UNCONNECTED__822, SYNOPSYS_UNCONNECTED__823, 
        SYNOPSYS_UNCONNECTED__824, SYNOPSYS_UNCONNECTED__825, 
        SYNOPSYS_UNCONNECTED__826, SYNOPSYS_UNCONNECTED__827, 
        SYNOPSYS_UNCONNECTED__828, SYNOPSYS_UNCONNECTED__829, 
        SYNOPSYS_UNCONNECTED__830, SYNOPSYS_UNCONNECTED__831, 
        SYNOPSYS_UNCONNECTED__832, SYNOPSYS_UNCONNECTED__833, 
        SYNOPSYS_UNCONNECTED__834;

  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(oglobal[0]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(oglobal[1]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(oglobal[2]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(oglobal[3]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(oglobal[4]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(oglobal[5]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(oglobal[6]) );
  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(oglobal[7]) );
  DFF \oglobal_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .Q(oglobal[8]) );
  DFF \oglobal_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .Q(oglobal[9]) );
  DFF \oglobal_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .Q(oglobal[10]) );
  DFF \oglobal_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .Q(oglobal[11]) );
  DFF \oglobal_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .Q(oglobal[12]) );
  DFF \oglobal_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .Q(oglobal[13]) );
  hamming_N16000_CC4_DW01_add_0 add_97 ( .A(oglobal), .B({1'b0, 1'b0, olocal}), 
        .CI(1'b0), .SUM(o) );
  hamming_N16000_CC4_DW01_add_1 add_1334_root_add_71_I928 ( .A({1'b0, N31899, 
        N31898, N31897, N31896, N31895, N31894, N31893, N31892, N31891, N31890, 
        N31889}), .B({N31912, N31911, N31910, N31909, N31908, N31907, N31906, 
        N31905, N31904, N31903, N31902, N31901}), .CI(1'b0), .SUM(olocal) );
  hamming_N16000_CC4_DW01_add_2 add_1335_root_add_71_I928 ( .A({1'b0, N31875, 
        N31874, N31873, N31872, N31871, N31870, N31869, N31868, N31867, N31866, 
        N31865}), .B({1'b0, N31887, N31886, N31885, N31884, N31883, N31882, 
        N31881, N31880, N31879, N31878, N31877}), .CI(1'b0), .SUM({N31912, 
        N31911, N31910, N31909, N31908, N31907, N31906, N31905, N31904, N31903, 
        N31902, N31901}) );
  hamming_N16000_CC4_DW01_add_3 add_1336_root_add_71_I928 ( .A({1'b0, 1'b0, 
        N31850, N31849, N31848, N31847, N31846, N31845, N31844, N31843, N31842, 
        N31841}), .B({1'b0, 1'b0, N31862, N31861, N31860, N31859, N31858, 
        N31857, N31856, N31855, N31854, N31853}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__0, N31899, N31898, N31897, N31896, N31895, 
        N31894, N31893, N31892, N31891, N31890, N31889}) );
  hamming_N16000_CC4_DW01_add_4 add_1337_root_add_71_I928 ( .A({1'b0, 1'b0, 
        N31826, N31825, N31824, N31823, N31822, N31821, N31820, N31819, N31818, 
        N31817}), .B({1'b0, 1'b0, N31838, N31837, N31836, N31835, N31834, 
        N31833, N31832, N31831, N31830, N31829}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1, N31887, N31886, N31885, N31884, N31883, 
        N31882, N31881, N31880, N31879, N31878, N31877}) );
  hamming_N16000_CC4_DW01_add_5 add_1338_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, N31801, N31800, N31799, N31798, N31797, N31796, N31795, N31794, 
        N31793}), .B({1'b0, 1'b0, N31814, N31813, N31812, N31811, N31810, 
        N31809, N31808, N31807, N31806, N31805}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__2, N31875, N31874, N31873, N31872, N31871, 
        N31870, N31869, N31868, N31867, N31866, N31865}) );
  hamming_N16000_CC4_DW01_add_6 add_1339_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, N31777, N31776, N31775, N31774, N31773, N31772, N31771, N31770, 
        N31769}), .B({1'b0, 1'b0, 1'b0, N31789, N31788, N31787, N31786, N31785, 
        N31784, N31783, N31782, N31781}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, N31862, N31861, 
        N31860, N31859, N31858, N31857, N31856, N31855, N31854, N31853}) );
  hamming_N16000_CC4_DW01_add_7 add_1340_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, N31753, N31752, N31751, N31750, N31749, N31748, N31747, N31746, 
        N31745}), .B({1'b0, 1'b0, 1'b0, N31765, N31764, N31763, N31762, N31761, 
        N31760, N31759, N31758, N31757}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, N31850, N31849, 
        N31848, N31847, N31846, N31845, N31844, N31843, N31842, N31841}) );
  hamming_N16000_CC4_DW01_add_8 add_1341_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, N31729, N31728, N31727, N31726, N31725, N31724, N31723, N31722, 
        N31721}), .B({1'b0, 1'b0, 1'b0, N31741, N31740, N31739, N31738, N31737, 
        N31736, N31735, N31734, N31733}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, N31838, N31837, 
        N31836, N31835, N31834, N31833, N31832, N31831, N31830, N31829}) );
  hamming_N16000_CC4_DW01_add_9 add_1342_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, N31705, N31704, N31703, N31702, N31701, N31700, N31699, N31698, 
        N31697}), .B({1'b0, 1'b0, 1'b0, N31717, N31716, N31715, N31714, N31713, 
        N31712, N31711, N31710, N31709}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, N31826, N31825, 
        N31824, N31823, N31822, N31821, N31820, N31819, N31818, N31817}) );
  hamming_N16000_CC4_DW01_add_10 add_1343_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N31680, N31679, N31678, N31677, N31676, N31675, N31674, 
        N31673}), .B({1'b0, 1'b0, 1'b0, N31693, N31692, N31691, N31690, N31689, 
        N31688, N31687, N31686, N31685}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, N31814, N31813, 
        N31812, N31811, N31810, N31809, N31808, N31807, N31806, N31805}) );
  hamming_N16000_CC4_DW01_add_11 add_1344_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N31656, N31655, N31654, N31653, N31652, N31651, N31650, 
        N31649}), .B({1'b0, 1'b0, 1'b0, 1'b0, N31668, N31667, N31666, N31665, 
        N31664, N31663, N31662, N31661}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N31801, N31800, N31799, N31798, N31797, 
        N31796, N31795, N31794, N31793}) );
  hamming_N16000_CC4_DW01_add_12 add_1345_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N31632, N31631, N31630, N31629, N31628, N31627, N31626, 
        N31625}), .B({1'b0, 1'b0, 1'b0, 1'b0, N31644, N31643, N31642, N31641, 
        N31640, N31639, N31638, N31637}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, N31789, N31788, N31787, N31786, N31785, 
        N31784, N31783, N31782, N31781}) );
  hamming_N16000_CC4_DW01_add_13 add_1346_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N31608, N31607, N31606, N31605, N31604, N31603, N31602, 
        N31601}), .B({1'b0, 1'b0, 1'b0, 1'b0, N31620, N31619, N31618, N31617, 
        N31616, N31615, N31614, N31613}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, N31777, N31776, N31775, N31774, N31773, 
        N31772, N31771, N31770, N31769}) );
  hamming_N16000_CC4_DW01_add_14 add_1347_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N31584, N31583, N31582, N31581, N31580, N31579, N31578, 
        N31577}), .B({1'b0, 1'b0, 1'b0, 1'b0, N31596, N31595, N31594, N31593, 
        N31592, N31591, N31590, N31589}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, N31765, N31764, N31763, N31762, N31761, 
        N31760, N31759, N31758, N31757}) );
  hamming_N16000_CC4_DW01_add_15 add_1348_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N31560, N31559, N31558, N31557, N31556, N31555, N31554, 
        N31553}), .B({1'b0, 1'b0, 1'b0, 1'b0, N31572, N31571, N31570, N31569, 
        N31568, N31567, N31566, N31565}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, N31753, N31752, N31751, N31750, N31749, 
        N31748, N31747, N31746, N31745}) );
  hamming_N16000_CC4_DW01_add_16 add_1349_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N31536, N31535, N31534, N31533, N31532, N31531, N31530, 
        N31529}), .B({1'b0, 1'b0, 1'b0, 1'b0, N31548, N31547, N31546, N31545, 
        N31544, N31543, N31542, N31541}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, N31741, N31740, N31739, N31738, N31737, 
        N31736, N31735, N31734, N31733}) );
  hamming_N16000_CC4_DW01_add_17 add_1350_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N31512, N31511, N31510, N31509, N31508, N31507, N31506, 
        N31505}), .B({1'b0, 1'b0, 1'b0, 1'b0, N31524, N31523, N31522, N31521, 
        N31520, N31519, N31518, N31517}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, N31729, N31728, N31727, N31726, N31725, 
        N31724, N31723, N31722, N31721}) );
  hamming_N16000_CC4_DW01_add_18 add_1351_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N31488, N31487, N31486, N31485, N31484, N31483, N31482, 
        N31481}), .B({1'b0, 1'b0, 1'b0, 1'b0, N31500, N31499, N31498, N31497, 
        N31496, N31495, N31494, N31493}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, N31717, N31716, N31715, N31714, N31713, 
        N31712, N31711, N31710, N31709}) );
  hamming_N16000_CC4_DW01_add_19 add_1352_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N31464, N31463, N31462, N31461, N31460, N31459, N31458, 
        N31457}), .B({1'b0, 1'b0, 1'b0, 1'b0, N31476, N31475, N31474, N31473, 
        N31472, N31471, N31470, N31469}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39, N31705, N31704, N31703, N31702, N31701, 
        N31700, N31699, N31698, N31697}) );
  hamming_N16000_CC4_DW01_add_20 add_1353_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N31440, N31439, N31438, N31437, N31436, N31435, N31434, 
        N31433}), .B({1'b0, 1'b0, 1'b0, 1'b0, N31452, N31451, N31450, N31449, 
        N31448, N31447, N31446, N31445}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, N31693, N31692, N31691, N31690, N31689, 
        N31688, N31687, N31686, N31685}) );
  hamming_N16000_CC4_DW01_add_21 add_1354_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31415, N31414, N31413, N31412, N31411, N31410, 
        N31409}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31427, N31426, N31425, 
        N31424, N31423, N31422, N31421}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44, 
        SYNOPSYS_UNCONNECTED__45, SYNOPSYS_UNCONNECTED__46, N31680, N31679, 
        N31678, N31677, N31676, N31675, N31674, N31673}) );
  hamming_N16000_CC4_DW01_add_22 add_1355_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31391, N31390, N31389, N31388, N31387, N31386, 
        N31385}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31403, N31402, N31401, 
        N31400, N31399, N31398, N31397}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__47, SYNOPSYS_UNCONNECTED__48, 
        SYNOPSYS_UNCONNECTED__49, SYNOPSYS_UNCONNECTED__50, N31668, N31667, 
        N31666, N31665, N31664, N31663, N31662, N31661}) );
  hamming_N16000_CC4_DW01_add_23 add_1356_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31367, N31366, N31365, N31364, N31363, N31362, 
        N31361}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31379, N31378, N31377, 
        N31376, N31375, N31374, N31373}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__51, SYNOPSYS_UNCONNECTED__52, 
        SYNOPSYS_UNCONNECTED__53, SYNOPSYS_UNCONNECTED__54, N31656, N31655, 
        N31654, N31653, N31652, N31651, N31650, N31649}) );
  hamming_N16000_CC4_DW01_add_24 add_1357_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31343, N31342, N31341, N31340, N31339, N31338, 
        N31337}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31355, N31354, N31353, 
        N31352, N31351, N31350, N31349}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__55, SYNOPSYS_UNCONNECTED__56, 
        SYNOPSYS_UNCONNECTED__57, SYNOPSYS_UNCONNECTED__58, N31644, N31643, 
        N31642, N31641, N31640, N31639, N31638, N31637}) );
  hamming_N16000_CC4_DW01_add_25 add_1358_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31319, N31318, N31317, N31316, N31315, N31314, 
        N31313}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31331, N31330, N31329, 
        N31328, N31327, N31326, N31325}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__59, SYNOPSYS_UNCONNECTED__60, 
        SYNOPSYS_UNCONNECTED__61, SYNOPSYS_UNCONNECTED__62, N31632, N31631, 
        N31630, N31629, N31628, N31627, N31626, N31625}) );
  hamming_N16000_CC4_DW01_add_26 add_1359_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31295, N31294, N31293, N31292, N31291, N31290, 
        N31289}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31307, N31306, N31305, 
        N31304, N31303, N31302, N31301}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__63, SYNOPSYS_UNCONNECTED__64, 
        SYNOPSYS_UNCONNECTED__65, SYNOPSYS_UNCONNECTED__66, N31620, N31619, 
        N31618, N31617, N31616, N31615, N31614, N31613}) );
  hamming_N16000_CC4_DW01_add_27 add_1360_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31271, N31270, N31269, N31268, N31267, N31266, 
        N31265}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31283, N31282, N31281, 
        N31280, N31279, N31278, N31277}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__67, SYNOPSYS_UNCONNECTED__68, 
        SYNOPSYS_UNCONNECTED__69, SYNOPSYS_UNCONNECTED__70, N31608, N31607, 
        N31606, N31605, N31604, N31603, N31602, N31601}) );
  hamming_N16000_CC4_DW01_add_28 add_1361_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31247, N31246, N31245, N31244, N31243, N31242, 
        N31241}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31259, N31258, N31257, 
        N31256, N31255, N31254, N31253}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__71, SYNOPSYS_UNCONNECTED__72, 
        SYNOPSYS_UNCONNECTED__73, SYNOPSYS_UNCONNECTED__74, N31596, N31595, 
        N31594, N31593, N31592, N31591, N31590, N31589}) );
  hamming_N16000_CC4_DW01_add_29 add_1362_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31223, N31222, N31221, N31220, N31219, N31218, 
        N31217}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31235, N31234, N31233, 
        N31232, N31231, N31230, N31229}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__75, SYNOPSYS_UNCONNECTED__76, 
        SYNOPSYS_UNCONNECTED__77, SYNOPSYS_UNCONNECTED__78, N31584, N31583, 
        N31582, N31581, N31580, N31579, N31578, N31577}) );
  hamming_N16000_CC4_DW01_add_30 add_1363_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31199, N31198, N31197, N31196, N31195, N31194, 
        N31193}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31211, N31210, N31209, 
        N31208, N31207, N31206, N31205}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__79, SYNOPSYS_UNCONNECTED__80, 
        SYNOPSYS_UNCONNECTED__81, SYNOPSYS_UNCONNECTED__82, N31572, N31571, 
        N31570, N31569, N31568, N31567, N31566, N31565}) );
  hamming_N16000_CC4_DW01_add_31 add_1364_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31175, N31174, N31173, N31172, N31171, N31170, 
        N31169}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31187, N31186, N31185, 
        N31184, N31183, N31182, N31181}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__83, SYNOPSYS_UNCONNECTED__84, 
        SYNOPSYS_UNCONNECTED__85, SYNOPSYS_UNCONNECTED__86, N31560, N31559, 
        N31558, N31557, N31556, N31555, N31554, N31553}) );
  hamming_N16000_CC4_DW01_add_32 add_1365_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31151, N31150, N31149, N31148, N31147, N31146, 
        N31145}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31163, N31162, N31161, 
        N31160, N31159, N31158, N31157}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__87, SYNOPSYS_UNCONNECTED__88, 
        SYNOPSYS_UNCONNECTED__89, SYNOPSYS_UNCONNECTED__90, N31548, N31547, 
        N31546, N31545, N31544, N31543, N31542, N31541}) );
  hamming_N16000_CC4_DW01_add_33 add_1366_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31127, N31126, N31125, N31124, N31123, N31122, 
        N31121}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31139, N31138, N31137, 
        N31136, N31135, N31134, N31133}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__91, SYNOPSYS_UNCONNECTED__92, 
        SYNOPSYS_UNCONNECTED__93, SYNOPSYS_UNCONNECTED__94, N31536, N31535, 
        N31534, N31533, N31532, N31531, N31530, N31529}) );
  hamming_N16000_CC4_DW01_add_34 add_1367_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31103, N31102, N31101, N31100, N31099, N31098, 
        N31097}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31115, N31114, N31113, 
        N31112, N31111, N31110, N31109}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__95, SYNOPSYS_UNCONNECTED__96, 
        SYNOPSYS_UNCONNECTED__97, SYNOPSYS_UNCONNECTED__98, N31524, N31523, 
        N31522, N31521, N31520, N31519, N31518, N31517}) );
  hamming_N16000_CC4_DW01_add_35 add_1368_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31079, N31078, N31077, N31076, N31075, N31074, 
        N31073}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31091, N31090, N31089, 
        N31088, N31087, N31086, N31085}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__99, SYNOPSYS_UNCONNECTED__100, 
        SYNOPSYS_UNCONNECTED__101, SYNOPSYS_UNCONNECTED__102, N31512, N31511, 
        N31510, N31509, N31508, N31507, N31506, N31505}) );
  hamming_N16000_CC4_DW01_add_36 add_1369_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31055, N31054, N31053, N31052, N31051, N31050, 
        N31049}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31067, N31066, N31065, 
        N31064, N31063, N31062, N31061}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__103, SYNOPSYS_UNCONNECTED__104, 
        SYNOPSYS_UNCONNECTED__105, SYNOPSYS_UNCONNECTED__106, N31500, N31499, 
        N31498, N31497, N31496, N31495, N31494, N31493}) );
  hamming_N16000_CC4_DW01_add_37 add_1370_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31031, N31030, N31029, N31028, N31027, N31026, 
        N31025}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31043, N31042, N31041, 
        N31040, N31039, N31038, N31037}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__107, SYNOPSYS_UNCONNECTED__108, 
        SYNOPSYS_UNCONNECTED__109, SYNOPSYS_UNCONNECTED__110, N31488, N31487, 
        N31486, N31485, N31484, N31483, N31482, N31481}) );
  hamming_N16000_CC4_DW01_add_38 add_1371_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31007, N31006, N31005, N31004, N31003, N31002, 
        N31001}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31019, N31018, N31017, 
        N31016, N31015, N31014, N31013}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__111, SYNOPSYS_UNCONNECTED__112, 
        SYNOPSYS_UNCONNECTED__113, SYNOPSYS_UNCONNECTED__114, N31476, N31475, 
        N31474, N31473, N31472, N31471, N31470, N31469}) );
  hamming_N16000_CC4_DW01_add_39 add_1372_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N30983, N30982, N30981, N30980, N30979, N30978, 
        N30977}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30995, N30994, N30993, 
        N30992, N30991, N30990, N30989}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__115, SYNOPSYS_UNCONNECTED__116, 
        SYNOPSYS_UNCONNECTED__117, SYNOPSYS_UNCONNECTED__118, N31464, N31463, 
        N31462, N31461, N31460, N31459, N31458, N31457}) );
  hamming_N16000_CC4_DW01_add_40 add_1373_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N30959, N30958, N30957, N30956, N30955, N30954, 
        N30953}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30971, N30970, N30969, 
        N30968, N30967, N30966, N30965}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__119, SYNOPSYS_UNCONNECTED__120, 
        SYNOPSYS_UNCONNECTED__121, SYNOPSYS_UNCONNECTED__122, N31452, N31451, 
        N31450, N31449, N31448, N31447, N31446, N31445}) );
  hamming_N16000_CC4_DW01_add_41 add_1374_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N30935, N30934, N30933, N30932, N30931, N30930, 
        N30929}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30947, N30946, N30945, 
        N30944, N30943, N30942, N30941}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__123, SYNOPSYS_UNCONNECTED__124, 
        SYNOPSYS_UNCONNECTED__125, SYNOPSYS_UNCONNECTED__126, N31440, N31439, 
        N31438, N31437, N31436, N31435, N31434, N31433}) );
  hamming_N16000_CC4_DW01_add_42 add_1375_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30910, N30909, N30908, N30907, N30906, N30905}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30922, N30921, N30920, N30919, 
        N30918, N30917}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, N31427, N31426, 
        N31425, N31424, N31423, N31422, N31421}) );
  hamming_N16000_CC4_DW01_add_43 add_1376_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30886, N30885, N30884, N30883, N30882, N30881}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30898, N30897, N30896, N30895, 
        N30894, N30893}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__132, 
        SYNOPSYS_UNCONNECTED__133, SYNOPSYS_UNCONNECTED__134, 
        SYNOPSYS_UNCONNECTED__135, SYNOPSYS_UNCONNECTED__136, N31415, N31414, 
        N31413, N31412, N31411, N31410, N31409}) );
  hamming_N16000_CC4_DW01_add_44 add_1377_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30862, N30861, N30860, N30859, N30858, N30857}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30874, N30873, N30872, N30871, 
        N30870, N30869}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, N31403, N31402, 
        N31401, N31400, N31399, N31398, N31397}) );
  hamming_N16000_CC4_DW01_add_45 add_1378_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30838, N30837, N30836, N30835, N30834, N30833}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30850, N30849, N30848, N30847, 
        N30846, N30845}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__142, 
        SYNOPSYS_UNCONNECTED__143, SYNOPSYS_UNCONNECTED__144, 
        SYNOPSYS_UNCONNECTED__145, SYNOPSYS_UNCONNECTED__146, N31391, N31390, 
        N31389, N31388, N31387, N31386, N31385}) );
  hamming_N16000_CC4_DW01_add_46 add_1379_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30814, N30813, N30812, N30811, N30810, N30809}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30826, N30825, N30824, N30823, 
        N30822, N30821}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, N31379, N31378, 
        N31377, N31376, N31375, N31374, N31373}) );
  hamming_N16000_CC4_DW01_add_47 add_1380_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30790, N30789, N30788, N30787, N30786, N30785}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30802, N30801, N30800, N30799, 
        N30798, N30797}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__152, 
        SYNOPSYS_UNCONNECTED__153, SYNOPSYS_UNCONNECTED__154, 
        SYNOPSYS_UNCONNECTED__155, SYNOPSYS_UNCONNECTED__156, N31367, N31366, 
        N31365, N31364, N31363, N31362, N31361}) );
  hamming_N16000_CC4_DW01_add_48 add_1381_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30766, N30765, N30764, N30763, N30762, N30761}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30778, N30777, N30776, N30775, 
        N30774, N30773}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__157, 
        SYNOPSYS_UNCONNECTED__158, SYNOPSYS_UNCONNECTED__159, 
        SYNOPSYS_UNCONNECTED__160, SYNOPSYS_UNCONNECTED__161, N31355, N31354, 
        N31353, N31352, N31351, N31350, N31349}) );
  hamming_N16000_CC4_DW01_add_49 add_1382_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30742, N30741, N30740, N30739, N30738, N30737}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30754, N30753, N30752, N30751, 
        N30750, N30749}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__162, 
        SYNOPSYS_UNCONNECTED__163, SYNOPSYS_UNCONNECTED__164, 
        SYNOPSYS_UNCONNECTED__165, SYNOPSYS_UNCONNECTED__166, N31343, N31342, 
        N31341, N31340, N31339, N31338, N31337}) );
  hamming_N16000_CC4_DW01_add_50 add_1383_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30718, N30717, N30716, N30715, N30714, N30713}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30730, N30729, N30728, N30727, 
        N30726, N30725}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__167, 
        SYNOPSYS_UNCONNECTED__168, SYNOPSYS_UNCONNECTED__169, 
        SYNOPSYS_UNCONNECTED__170, SYNOPSYS_UNCONNECTED__171, N31331, N31330, 
        N31329, N31328, N31327, N31326, N31325}) );
  hamming_N16000_CC4_DW01_add_51 add_1384_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30694, N30693, N30692, N30691, N30690, N30689}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30706, N30705, N30704, N30703, 
        N30702, N30701}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__172, 
        SYNOPSYS_UNCONNECTED__173, SYNOPSYS_UNCONNECTED__174, 
        SYNOPSYS_UNCONNECTED__175, SYNOPSYS_UNCONNECTED__176, N31319, N31318, 
        N31317, N31316, N31315, N31314, N31313}) );
  hamming_N16000_CC4_DW01_add_52 add_1385_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30670, N30669, N30668, N30667, N30666, N30665}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30682, N30681, N30680, N30679, 
        N30678, N30677}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__177, 
        SYNOPSYS_UNCONNECTED__178, SYNOPSYS_UNCONNECTED__179, 
        SYNOPSYS_UNCONNECTED__180, SYNOPSYS_UNCONNECTED__181, N31307, N31306, 
        N31305, N31304, N31303, N31302, N31301}) );
  hamming_N16000_CC4_DW01_add_53 add_1386_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30646, N30645, N30644, N30643, N30642, N30641}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30658, N30657, N30656, N30655, 
        N30654, N30653}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__182, 
        SYNOPSYS_UNCONNECTED__183, SYNOPSYS_UNCONNECTED__184, 
        SYNOPSYS_UNCONNECTED__185, SYNOPSYS_UNCONNECTED__186, N31295, N31294, 
        N31293, N31292, N31291, N31290, N31289}) );
  hamming_N16000_CC4_DW01_add_54 add_1387_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30622, N30621, N30620, N30619, N30618, N30617}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30634, N30633, N30632, N30631, 
        N30630, N30629}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__187, 
        SYNOPSYS_UNCONNECTED__188, SYNOPSYS_UNCONNECTED__189, 
        SYNOPSYS_UNCONNECTED__190, SYNOPSYS_UNCONNECTED__191, N31283, N31282, 
        N31281, N31280, N31279, N31278, N31277}) );
  hamming_N16000_CC4_DW01_add_55 add_1388_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30598, N30597, N30596, N30595, N30594, N30593}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30610, N30609, N30608, N30607, 
        N30606, N30605}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__192, 
        SYNOPSYS_UNCONNECTED__193, SYNOPSYS_UNCONNECTED__194, 
        SYNOPSYS_UNCONNECTED__195, SYNOPSYS_UNCONNECTED__196, N31271, N31270, 
        N31269, N31268, N31267, N31266, N31265}) );
  hamming_N16000_CC4_DW01_add_56 add_1389_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30574, N30573, N30572, N30571, N30570, N30569}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30586, N30585, N30584, N30583, 
        N30582, N30581}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__197, 
        SYNOPSYS_UNCONNECTED__198, SYNOPSYS_UNCONNECTED__199, 
        SYNOPSYS_UNCONNECTED__200, SYNOPSYS_UNCONNECTED__201, N31259, N31258, 
        N31257, N31256, N31255, N31254, N31253}) );
  hamming_N16000_CC4_DW01_add_57 add_1390_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30550, N30549, N30548, N30547, N30546, N30545}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30562, N30561, N30560, N30559, 
        N30558, N30557}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__202, 
        SYNOPSYS_UNCONNECTED__203, SYNOPSYS_UNCONNECTED__204, 
        SYNOPSYS_UNCONNECTED__205, SYNOPSYS_UNCONNECTED__206, N31247, N31246, 
        N31245, N31244, N31243, N31242, N31241}) );
  hamming_N16000_CC4_DW01_add_58 add_1391_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30526, N30525, N30524, N30523, N30522, N30521}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30538, N30537, N30536, N30535, 
        N30534, N30533}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__207, 
        SYNOPSYS_UNCONNECTED__208, SYNOPSYS_UNCONNECTED__209, 
        SYNOPSYS_UNCONNECTED__210, SYNOPSYS_UNCONNECTED__211, N31235, N31234, 
        N31233, N31232, N31231, N31230, N31229}) );
  hamming_N16000_CC4_DW01_add_59 add_1392_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30502, N30501, N30500, N30499, N30498, N30497}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30514, N30513, N30512, N30511, 
        N30510, N30509}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__212, 
        SYNOPSYS_UNCONNECTED__213, SYNOPSYS_UNCONNECTED__214, 
        SYNOPSYS_UNCONNECTED__215, SYNOPSYS_UNCONNECTED__216, N31223, N31222, 
        N31221, N31220, N31219, N31218, N31217}) );
  hamming_N16000_CC4_DW01_add_60 add_1393_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30478, N30477, N30476, N30475, N30474, N30473}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30490, N30489, N30488, N30487, 
        N30486, N30485}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__217, 
        SYNOPSYS_UNCONNECTED__218, SYNOPSYS_UNCONNECTED__219, 
        SYNOPSYS_UNCONNECTED__220, SYNOPSYS_UNCONNECTED__221, N31211, N31210, 
        N31209, N31208, N31207, N31206, N31205}) );
  hamming_N16000_CC4_DW01_add_61 add_1394_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30454, N30453, N30452, N30451, N30450, N30449}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30466, N30465, N30464, N30463, 
        N30462, N30461}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__222, 
        SYNOPSYS_UNCONNECTED__223, SYNOPSYS_UNCONNECTED__224, 
        SYNOPSYS_UNCONNECTED__225, SYNOPSYS_UNCONNECTED__226, N31199, N31198, 
        N31197, N31196, N31195, N31194, N31193}) );
  hamming_N16000_CC4_DW01_add_62 add_1395_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30430, N30429, N30428, N30427, N30426, N30425}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30442, N30441, N30440, N30439, 
        N30438, N30437}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__227, 
        SYNOPSYS_UNCONNECTED__228, SYNOPSYS_UNCONNECTED__229, 
        SYNOPSYS_UNCONNECTED__230, SYNOPSYS_UNCONNECTED__231, N31187, N31186, 
        N31185, N31184, N31183, N31182, N31181}) );
  hamming_N16000_CC4_DW01_add_63 add_1396_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30406, N30405, N30404, N30403, N30402, N30401}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30418, N30417, N30416, N30415, 
        N30414, N30413}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__232, 
        SYNOPSYS_UNCONNECTED__233, SYNOPSYS_UNCONNECTED__234, 
        SYNOPSYS_UNCONNECTED__235, SYNOPSYS_UNCONNECTED__236, N31175, N31174, 
        N31173, N31172, N31171, N31170, N31169}) );
  hamming_N16000_CC4_DW01_add_64 add_1397_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30382, N30381, N30380, N30379, N30378, N30377}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30394, N30393, N30392, N30391, 
        N30390, N30389}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__237, 
        SYNOPSYS_UNCONNECTED__238, SYNOPSYS_UNCONNECTED__239, 
        SYNOPSYS_UNCONNECTED__240, SYNOPSYS_UNCONNECTED__241, N31163, N31162, 
        N31161, N31160, N31159, N31158, N31157}) );
  hamming_N16000_CC4_DW01_add_65 add_1398_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30358, N30357, N30356, N30355, N30354, N30353}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30370, N30369, N30368, N30367, 
        N30366, N30365}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__242, 
        SYNOPSYS_UNCONNECTED__243, SYNOPSYS_UNCONNECTED__244, 
        SYNOPSYS_UNCONNECTED__245, SYNOPSYS_UNCONNECTED__246, N31151, N31150, 
        N31149, N31148, N31147, N31146, N31145}) );
  hamming_N16000_CC4_DW01_add_66 add_1399_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30334, N30333, N30332, N30331, N30330, N30329}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30346, N30345, N30344, N30343, 
        N30342, N30341}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__247, 
        SYNOPSYS_UNCONNECTED__248, SYNOPSYS_UNCONNECTED__249, 
        SYNOPSYS_UNCONNECTED__250, SYNOPSYS_UNCONNECTED__251, N31139, N31138, 
        N31137, N31136, N31135, N31134, N31133}) );
  hamming_N16000_CC4_DW01_add_67 add_1400_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30310, N30309, N30308, N30307, N30306, N30305}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30322, N30321, N30320, N30319, 
        N30318, N30317}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__252, 
        SYNOPSYS_UNCONNECTED__253, SYNOPSYS_UNCONNECTED__254, 
        SYNOPSYS_UNCONNECTED__255, SYNOPSYS_UNCONNECTED__256, N31127, N31126, 
        N31125, N31124, N31123, N31122, N31121}) );
  hamming_N16000_CC4_DW01_add_68 add_1401_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30286, N30285, N30284, N30283, N30282, N30281}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30298, N30297, N30296, N30295, 
        N30294, N30293}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__257, 
        SYNOPSYS_UNCONNECTED__258, SYNOPSYS_UNCONNECTED__259, 
        SYNOPSYS_UNCONNECTED__260, SYNOPSYS_UNCONNECTED__261, N31115, N31114, 
        N31113, N31112, N31111, N31110, N31109}) );
  hamming_N16000_CC4_DW01_add_69 add_1402_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30262, N30261, N30260, N30259, N30258, N30257}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30274, N30273, N30272, N30271, 
        N30270, N30269}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__262, 
        SYNOPSYS_UNCONNECTED__263, SYNOPSYS_UNCONNECTED__264, 
        SYNOPSYS_UNCONNECTED__265, SYNOPSYS_UNCONNECTED__266, N31103, N31102, 
        N31101, N31100, N31099, N31098, N31097}) );
  hamming_N16000_CC4_DW01_add_70 add_1403_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30238, N30237, N30236, N30235, N30234, N30233}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30250, N30249, N30248, N30247, 
        N30246, N30245}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__267, 
        SYNOPSYS_UNCONNECTED__268, SYNOPSYS_UNCONNECTED__269, 
        SYNOPSYS_UNCONNECTED__270, SYNOPSYS_UNCONNECTED__271, N31091, N31090, 
        N31089, N31088, N31087, N31086, N31085}) );
  hamming_N16000_CC4_DW01_add_71 add_1404_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30214, N30213, N30212, N30211, N30210, N30209}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30226, N30225, N30224, N30223, 
        N30222, N30221}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__272, 
        SYNOPSYS_UNCONNECTED__273, SYNOPSYS_UNCONNECTED__274, 
        SYNOPSYS_UNCONNECTED__275, SYNOPSYS_UNCONNECTED__276, N31079, N31078, 
        N31077, N31076, N31075, N31074, N31073}) );
  hamming_N16000_CC4_DW01_add_72 add_1405_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30190, N30189, N30188, N30187, N30186, N30185}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30202, N30201, N30200, N30199, 
        N30198, N30197}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__277, 
        SYNOPSYS_UNCONNECTED__278, SYNOPSYS_UNCONNECTED__279, 
        SYNOPSYS_UNCONNECTED__280, SYNOPSYS_UNCONNECTED__281, N31067, N31066, 
        N31065, N31064, N31063, N31062, N31061}) );
  hamming_N16000_CC4_DW01_add_73 add_1406_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30166, N30165, N30164, N30163, N30162, N30161}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30178, N30177, N30176, N30175, 
        N30174, N30173}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__282, 
        SYNOPSYS_UNCONNECTED__283, SYNOPSYS_UNCONNECTED__284, 
        SYNOPSYS_UNCONNECTED__285, SYNOPSYS_UNCONNECTED__286, N31055, N31054, 
        N31053, N31052, N31051, N31050, N31049}) );
  hamming_N16000_CC4_DW01_add_74 add_1407_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30142, N30141, N30140, N30139, N30138, N30137}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30154, N30153, N30152, N30151, 
        N30150, N30149}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__287, 
        SYNOPSYS_UNCONNECTED__288, SYNOPSYS_UNCONNECTED__289, 
        SYNOPSYS_UNCONNECTED__290, SYNOPSYS_UNCONNECTED__291, N31043, N31042, 
        N31041, N31040, N31039, N31038, N31037}) );
  hamming_N16000_CC4_DW01_add_75 add_1408_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30118, N30117, N30116, N30115, N30114, N30113}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30130, N30129, N30128, N30127, 
        N30126, N30125}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__292, 
        SYNOPSYS_UNCONNECTED__293, SYNOPSYS_UNCONNECTED__294, 
        SYNOPSYS_UNCONNECTED__295, SYNOPSYS_UNCONNECTED__296, N31031, N31030, 
        N31029, N31028, N31027, N31026, N31025}) );
  hamming_N16000_CC4_DW01_add_76 add_1409_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30094, N30093, N30092, N30091, N30090, N30089}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30106, N30105, N30104, N30103, 
        N30102, N30101}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__297, 
        SYNOPSYS_UNCONNECTED__298, SYNOPSYS_UNCONNECTED__299, 
        SYNOPSYS_UNCONNECTED__300, SYNOPSYS_UNCONNECTED__301, N31019, N31018, 
        N31017, N31016, N31015, N31014, N31013}) );
  hamming_N16000_CC4_DW01_add_77 add_1410_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30070, N30069, N30068, N30067, N30066, N30065}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30082, N30081, N30080, N30079, 
        N30078, N30077}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__302, 
        SYNOPSYS_UNCONNECTED__303, SYNOPSYS_UNCONNECTED__304, 
        SYNOPSYS_UNCONNECTED__305, SYNOPSYS_UNCONNECTED__306, N31007, N31006, 
        N31005, N31004, N31003, N31002, N31001}) );
  hamming_N16000_CC4_DW01_add_78 add_1411_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30046, N30045, N30044, N30043, N30042, N30041}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30058, N30057, N30056, N30055, 
        N30054, N30053}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__307, 
        SYNOPSYS_UNCONNECTED__308, SYNOPSYS_UNCONNECTED__309, 
        SYNOPSYS_UNCONNECTED__310, SYNOPSYS_UNCONNECTED__311, N30995, N30994, 
        N30993, N30992, N30991, N30990, N30989}) );
  hamming_N16000_CC4_DW01_add_79 add_1412_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30022, N30021, N30020, N30019, N30018, N30017}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30034, N30033, N30032, N30031, 
        N30030, N30029}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__312, 
        SYNOPSYS_UNCONNECTED__313, SYNOPSYS_UNCONNECTED__314, 
        SYNOPSYS_UNCONNECTED__315, SYNOPSYS_UNCONNECTED__316, N30983, N30982, 
        N30981, N30980, N30979, N30978, N30977}) );
  hamming_N16000_CC4_DW01_add_80 add_1413_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N29998, N29997, N29996, N29995, N29994, N29993}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30010, N30009, N30008, N30007, 
        N30006, N30005}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__317, 
        SYNOPSYS_UNCONNECTED__318, SYNOPSYS_UNCONNECTED__319, 
        SYNOPSYS_UNCONNECTED__320, SYNOPSYS_UNCONNECTED__321, N30971, N30970, 
        N30969, N30968, N30967, N30966, N30965}) );
  hamming_N16000_CC4_DW01_add_81 add_1414_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N29974, N29973, N29972, N29971, N29970, N29969}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29986, N29985, N29984, N29983, 
        N29982, N29981}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__322, 
        SYNOPSYS_UNCONNECTED__323, SYNOPSYS_UNCONNECTED__324, 
        SYNOPSYS_UNCONNECTED__325, SYNOPSYS_UNCONNECTED__326, N30959, N30958, 
        N30957, N30956, N30955, N30954, N30953}) );
  hamming_N16000_CC4_DW01_add_82 add_1415_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N29950, N29949, N29948, N29947, N29946, N29945}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29962, N29961, N29960, N29959, 
        N29958, N29957}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__327, 
        SYNOPSYS_UNCONNECTED__328, SYNOPSYS_UNCONNECTED__329, 
        SYNOPSYS_UNCONNECTED__330, SYNOPSYS_UNCONNECTED__331, N30947, N30946, 
        N30945, N30944, N30943, N30942, N30941}) );
  hamming_N16000_CC4_DW01_add_83 add_1416_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29925, N29924, N29923, N29922, N29921}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29938, N29937, N29936, N29935, 
        N29934, N29933}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__332, 
        SYNOPSYS_UNCONNECTED__333, SYNOPSYS_UNCONNECTED__334, 
        SYNOPSYS_UNCONNECTED__335, SYNOPSYS_UNCONNECTED__336, N30935, N30934, 
        N30933, N30932, N30931, N30930, N30929}) );
  hamming_N16000_CC4_DW01_add_84 add_1417_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29901, N29900, N29899, N29898, N29897}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29913, N29912, N29911, 
        N29910, N29909}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__337, 
        SYNOPSYS_UNCONNECTED__338, SYNOPSYS_UNCONNECTED__339, 
        SYNOPSYS_UNCONNECTED__340, SYNOPSYS_UNCONNECTED__341, 
        SYNOPSYS_UNCONNECTED__342, N30922, N30921, N30920, N30919, N30918, 
        N30917}) );
  hamming_N16000_CC4_DW01_add_85 add_1418_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29877, N29876, N29875, N29874, N29873}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29889, N29888, N29887, 
        N29886, N29885}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__343, 
        SYNOPSYS_UNCONNECTED__344, SYNOPSYS_UNCONNECTED__345, 
        SYNOPSYS_UNCONNECTED__346, SYNOPSYS_UNCONNECTED__347, 
        SYNOPSYS_UNCONNECTED__348, N30910, N30909, N30908, N30907, N30906, 
        N30905}) );
  hamming_N16000_CC4_DW01_add_86 add_1419_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29853, N29852, N29851, N29850, N29849}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29865, N29864, N29863, 
        N29862, N29861}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__349, 
        SYNOPSYS_UNCONNECTED__350, SYNOPSYS_UNCONNECTED__351, 
        SYNOPSYS_UNCONNECTED__352, SYNOPSYS_UNCONNECTED__353, 
        SYNOPSYS_UNCONNECTED__354, N30898, N30897, N30896, N30895, N30894, 
        N30893}) );
  hamming_N16000_CC4_DW01_add_87 add_1420_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29829, N29828, N29827, N29826, N29825}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29841, N29840, N29839, 
        N29838, N29837}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__355, 
        SYNOPSYS_UNCONNECTED__356, SYNOPSYS_UNCONNECTED__357, 
        SYNOPSYS_UNCONNECTED__358, SYNOPSYS_UNCONNECTED__359, 
        SYNOPSYS_UNCONNECTED__360, N30886, N30885, N30884, N30883, N30882, 
        N30881}) );
  hamming_N16000_CC4_DW01_add_88 add_1421_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29805, N29804, N29803, N29802, N29801}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29817, N29816, N29815, 
        N29814, N29813}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__361, 
        SYNOPSYS_UNCONNECTED__362, SYNOPSYS_UNCONNECTED__363, 
        SYNOPSYS_UNCONNECTED__364, SYNOPSYS_UNCONNECTED__365, 
        SYNOPSYS_UNCONNECTED__366, N30874, N30873, N30872, N30871, N30870, 
        N30869}) );
  hamming_N16000_CC4_DW01_add_89 add_1422_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29781, N29780, N29779, N29778, N29777}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29793, N29792, N29791, 
        N29790, N29789}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__367, 
        SYNOPSYS_UNCONNECTED__368, SYNOPSYS_UNCONNECTED__369, 
        SYNOPSYS_UNCONNECTED__370, SYNOPSYS_UNCONNECTED__371, 
        SYNOPSYS_UNCONNECTED__372, N30862, N30861, N30860, N30859, N30858, 
        N30857}) );
  hamming_N16000_CC4_DW01_add_90 add_1423_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29757, N29756, N29755, N29754, N29753}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29769, N29768, N29767, 
        N29766, N29765}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__373, 
        SYNOPSYS_UNCONNECTED__374, SYNOPSYS_UNCONNECTED__375, 
        SYNOPSYS_UNCONNECTED__376, SYNOPSYS_UNCONNECTED__377, 
        SYNOPSYS_UNCONNECTED__378, N30850, N30849, N30848, N30847, N30846, 
        N30845}) );
  hamming_N16000_CC4_DW01_add_91 add_1424_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29733, N29732, N29731, N29730, N29729}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29745, N29744, N29743, 
        N29742, N29741}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__379, 
        SYNOPSYS_UNCONNECTED__380, SYNOPSYS_UNCONNECTED__381, 
        SYNOPSYS_UNCONNECTED__382, SYNOPSYS_UNCONNECTED__383, 
        SYNOPSYS_UNCONNECTED__384, N30838, N30837, N30836, N30835, N30834, 
        N30833}) );
  hamming_N16000_CC4_DW01_add_92 add_1425_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29709, N29708, N29707, N29706, N29705}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29721, N29720, N29719, 
        N29718, N29717}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__385, 
        SYNOPSYS_UNCONNECTED__386, SYNOPSYS_UNCONNECTED__387, 
        SYNOPSYS_UNCONNECTED__388, SYNOPSYS_UNCONNECTED__389, 
        SYNOPSYS_UNCONNECTED__390, N30826, N30825, N30824, N30823, N30822, 
        N30821}) );
  hamming_N16000_CC4_DW01_add_93 add_1426_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29685, N29684, N29683, N29682, N29681}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29697, N29696, N29695, 
        N29694, N29693}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__391, 
        SYNOPSYS_UNCONNECTED__392, SYNOPSYS_UNCONNECTED__393, 
        SYNOPSYS_UNCONNECTED__394, SYNOPSYS_UNCONNECTED__395, 
        SYNOPSYS_UNCONNECTED__396, N30814, N30813, N30812, N30811, N30810, 
        N30809}) );
  hamming_N16000_CC4_DW01_add_94 add_1427_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29661, N29660, N29659, N29658, N29657}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29673, N29672, N29671, 
        N29670, N29669}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__397, 
        SYNOPSYS_UNCONNECTED__398, SYNOPSYS_UNCONNECTED__399, 
        SYNOPSYS_UNCONNECTED__400, SYNOPSYS_UNCONNECTED__401, 
        SYNOPSYS_UNCONNECTED__402, N30802, N30801, N30800, N30799, N30798, 
        N30797}) );
  hamming_N16000_CC4_DW01_add_95 add_1428_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29637, N29636, N29635, N29634, N29633}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29649, N29648, N29647, 
        N29646, N29645}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__403, 
        SYNOPSYS_UNCONNECTED__404, SYNOPSYS_UNCONNECTED__405, 
        SYNOPSYS_UNCONNECTED__406, SYNOPSYS_UNCONNECTED__407, 
        SYNOPSYS_UNCONNECTED__408, N30790, N30789, N30788, N30787, N30786, 
        N30785}) );
  hamming_N16000_CC4_DW01_add_96 add_1429_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29613, N29612, N29611, N29610, N29609}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29625, N29624, N29623, 
        N29622, N29621}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__409, 
        SYNOPSYS_UNCONNECTED__410, SYNOPSYS_UNCONNECTED__411, 
        SYNOPSYS_UNCONNECTED__412, SYNOPSYS_UNCONNECTED__413, 
        SYNOPSYS_UNCONNECTED__414, N30778, N30777, N30776, N30775, N30774, 
        N30773}) );
  hamming_N16000_CC4_DW01_add_97 add_1430_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29589, N29588, N29587, N29586, N29585}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29601, N29600, N29599, 
        N29598, N29597}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__415, 
        SYNOPSYS_UNCONNECTED__416, SYNOPSYS_UNCONNECTED__417, 
        SYNOPSYS_UNCONNECTED__418, SYNOPSYS_UNCONNECTED__419, 
        SYNOPSYS_UNCONNECTED__420, N30766, N30765, N30764, N30763, N30762, 
        N30761}) );
  hamming_N16000_CC4_DW01_add_98 add_1431_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29565, N29564, N29563, N29562, N29561}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29577, N29576, N29575, 
        N29574, N29573}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__421, 
        SYNOPSYS_UNCONNECTED__422, SYNOPSYS_UNCONNECTED__423, 
        SYNOPSYS_UNCONNECTED__424, SYNOPSYS_UNCONNECTED__425, 
        SYNOPSYS_UNCONNECTED__426, N30754, N30753, N30752, N30751, N30750, 
        N30749}) );
  hamming_N16000_CC4_DW01_add_99 add_1432_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29541, N29540, N29539, N29538, N29537}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29553, N29552, N29551, 
        N29550, N29549}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__427, 
        SYNOPSYS_UNCONNECTED__428, SYNOPSYS_UNCONNECTED__429, 
        SYNOPSYS_UNCONNECTED__430, SYNOPSYS_UNCONNECTED__431, 
        SYNOPSYS_UNCONNECTED__432, N30742, N30741, N30740, N30739, N30738, 
        N30737}) );
  hamming_N16000_CC4_DW01_add_100 add_1433_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29517, N29516, N29515, N29514, N29513}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29529, N29528, N29527, 
        N29526, N29525}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__433, 
        SYNOPSYS_UNCONNECTED__434, SYNOPSYS_UNCONNECTED__435, 
        SYNOPSYS_UNCONNECTED__436, SYNOPSYS_UNCONNECTED__437, 
        SYNOPSYS_UNCONNECTED__438, N30730, N30729, N30728, N30727, N30726, 
        N30725}) );
  hamming_N16000_CC4_DW01_add_101 add_1434_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29493, N29492, N29491, N29490, N29489}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29505, N29504, N29503, 
        N29502, N29501}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__439, 
        SYNOPSYS_UNCONNECTED__440, SYNOPSYS_UNCONNECTED__441, 
        SYNOPSYS_UNCONNECTED__442, SYNOPSYS_UNCONNECTED__443, 
        SYNOPSYS_UNCONNECTED__444, N30718, N30717, N30716, N30715, N30714, 
        N30713}) );
  hamming_N16000_CC4_DW01_add_102 add_1435_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29469, N29468, N29467, N29466, N29465}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29481, N29480, N29479, 
        N29478, N29477}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__445, 
        SYNOPSYS_UNCONNECTED__446, SYNOPSYS_UNCONNECTED__447, 
        SYNOPSYS_UNCONNECTED__448, SYNOPSYS_UNCONNECTED__449, 
        SYNOPSYS_UNCONNECTED__450, N30706, N30705, N30704, N30703, N30702, 
        N30701}) );
  hamming_N16000_CC4_DW01_add_103 add_1436_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29445, N29444, N29443, N29442, N29441}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29457, N29456, N29455, 
        N29454, N29453}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__451, 
        SYNOPSYS_UNCONNECTED__452, SYNOPSYS_UNCONNECTED__453, 
        SYNOPSYS_UNCONNECTED__454, SYNOPSYS_UNCONNECTED__455, 
        SYNOPSYS_UNCONNECTED__456, N30694, N30693, N30692, N30691, N30690, 
        N30689}) );
  hamming_N16000_CC4_DW01_add_104 add_1437_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29421, N29420, N29419, N29418, N29417}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29433, N29432, N29431, 
        N29430, N29429}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__457, 
        SYNOPSYS_UNCONNECTED__458, SYNOPSYS_UNCONNECTED__459, 
        SYNOPSYS_UNCONNECTED__460, SYNOPSYS_UNCONNECTED__461, 
        SYNOPSYS_UNCONNECTED__462, N30682, N30681, N30680, N30679, N30678, 
        N30677}) );
  hamming_N16000_CC4_DW01_add_105 add_1438_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29397, N29396, N29395, N29394, N29393}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29409, N29408, N29407, 
        N29406, N29405}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__463, 
        SYNOPSYS_UNCONNECTED__464, SYNOPSYS_UNCONNECTED__465, 
        SYNOPSYS_UNCONNECTED__466, SYNOPSYS_UNCONNECTED__467, 
        SYNOPSYS_UNCONNECTED__468, N30670, N30669, N30668, N30667, N30666, 
        N30665}) );
  hamming_N16000_CC4_DW01_add_106 add_1439_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29373, N29372, N29371, N29370, N29369}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29385, N29384, N29383, 
        N29382, N29381}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__469, 
        SYNOPSYS_UNCONNECTED__470, SYNOPSYS_UNCONNECTED__471, 
        SYNOPSYS_UNCONNECTED__472, SYNOPSYS_UNCONNECTED__473, 
        SYNOPSYS_UNCONNECTED__474, N30658, N30657, N30656, N30655, N30654, 
        N30653}) );
  hamming_N16000_CC4_DW01_add_107 add_1440_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29349, N29348, N29347, N29346, N29345}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29361, N29360, N29359, 
        N29358, N29357}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__475, 
        SYNOPSYS_UNCONNECTED__476, SYNOPSYS_UNCONNECTED__477, 
        SYNOPSYS_UNCONNECTED__478, SYNOPSYS_UNCONNECTED__479, 
        SYNOPSYS_UNCONNECTED__480, N30646, N30645, N30644, N30643, N30642, 
        N30641}) );
  hamming_N16000_CC4_DW01_add_108 add_1441_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29325, N29324, N29323, N29322, N29321}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29337, N29336, N29335, 
        N29334, N29333}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__481, 
        SYNOPSYS_UNCONNECTED__482, SYNOPSYS_UNCONNECTED__483, 
        SYNOPSYS_UNCONNECTED__484, SYNOPSYS_UNCONNECTED__485, 
        SYNOPSYS_UNCONNECTED__486, N30634, N30633, N30632, N30631, N30630, 
        N30629}) );
  hamming_N16000_CC4_DW01_add_109 add_1442_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29301, N29300, N29299, N29298, N29297}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29313, N29312, N29311, 
        N29310, N29309}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__487, 
        SYNOPSYS_UNCONNECTED__488, SYNOPSYS_UNCONNECTED__489, 
        SYNOPSYS_UNCONNECTED__490, SYNOPSYS_UNCONNECTED__491, 
        SYNOPSYS_UNCONNECTED__492, N30622, N30621, N30620, N30619, N30618, 
        N30617}) );
  hamming_N16000_CC4_DW01_add_110 add_1443_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29277, N29276, N29275, N29274, N29273}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29289, N29288, N29287, 
        N29286, N29285}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__493, 
        SYNOPSYS_UNCONNECTED__494, SYNOPSYS_UNCONNECTED__495, 
        SYNOPSYS_UNCONNECTED__496, SYNOPSYS_UNCONNECTED__497, 
        SYNOPSYS_UNCONNECTED__498, N30610, N30609, N30608, N30607, N30606, 
        N30605}) );
  hamming_N16000_CC4_DW01_add_111 add_1444_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29253, N29252, N29251, N29250, N29249}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29265, N29264, N29263, 
        N29262, N29261}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__499, 
        SYNOPSYS_UNCONNECTED__500, SYNOPSYS_UNCONNECTED__501, 
        SYNOPSYS_UNCONNECTED__502, SYNOPSYS_UNCONNECTED__503, 
        SYNOPSYS_UNCONNECTED__504, N30598, N30597, N30596, N30595, N30594, 
        N30593}) );
  hamming_N16000_CC4_DW01_add_112 add_1445_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29229, N29228, N29227, N29226, N29225}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29241, N29240, N29239, 
        N29238, N29237}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__505, 
        SYNOPSYS_UNCONNECTED__506, SYNOPSYS_UNCONNECTED__507, 
        SYNOPSYS_UNCONNECTED__508, SYNOPSYS_UNCONNECTED__509, 
        SYNOPSYS_UNCONNECTED__510, N30586, N30585, N30584, N30583, N30582, 
        N30581}) );
  hamming_N16000_CC4_DW01_add_113 add_1446_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29205, N29204, N29203, N29202, N29201}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29217, N29216, N29215, 
        N29214, N29213}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__511, 
        SYNOPSYS_UNCONNECTED__512, SYNOPSYS_UNCONNECTED__513, 
        SYNOPSYS_UNCONNECTED__514, SYNOPSYS_UNCONNECTED__515, 
        SYNOPSYS_UNCONNECTED__516, N30574, N30573, N30572, N30571, N30570, 
        N30569}) );
  hamming_N16000_CC4_DW01_add_114 add_1447_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29181, N29180, N29179, N29178, N29177}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29193, N29192, N29191, 
        N29190, N29189}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__517, 
        SYNOPSYS_UNCONNECTED__518, SYNOPSYS_UNCONNECTED__519, 
        SYNOPSYS_UNCONNECTED__520, SYNOPSYS_UNCONNECTED__521, 
        SYNOPSYS_UNCONNECTED__522, N30562, N30561, N30560, N30559, N30558, 
        N30557}) );
  hamming_N16000_CC4_DW01_add_115 add_1448_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29157, N29156, N29155, N29154, N29153}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29169, N29168, N29167, 
        N29166, N29165}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__523, 
        SYNOPSYS_UNCONNECTED__524, SYNOPSYS_UNCONNECTED__525, 
        SYNOPSYS_UNCONNECTED__526, SYNOPSYS_UNCONNECTED__527, 
        SYNOPSYS_UNCONNECTED__528, N30550, N30549, N30548, N30547, N30546, 
        N30545}) );
  hamming_N16000_CC4_DW01_add_116 add_1449_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29133, N29132, N29131, N29130, N29129}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29145, N29144, N29143, 
        N29142, N29141}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__529, 
        SYNOPSYS_UNCONNECTED__530, SYNOPSYS_UNCONNECTED__531, 
        SYNOPSYS_UNCONNECTED__532, SYNOPSYS_UNCONNECTED__533, 
        SYNOPSYS_UNCONNECTED__534, N30538, N30537, N30536, N30535, N30534, 
        N30533}) );
  hamming_N16000_CC4_DW01_add_117 add_1450_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29109, N29108, N29107, N29106, N29105}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29121, N29120, N29119, 
        N29118, N29117}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__535, 
        SYNOPSYS_UNCONNECTED__536, SYNOPSYS_UNCONNECTED__537, 
        SYNOPSYS_UNCONNECTED__538, SYNOPSYS_UNCONNECTED__539, 
        SYNOPSYS_UNCONNECTED__540, N30526, N30525, N30524, N30523, N30522, 
        N30521}) );
  hamming_N16000_CC4_DW01_add_118 add_1451_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29085, N29084, N29083, N29082, N29081}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29097, N29096, N29095, 
        N29094, N29093}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__541, 
        SYNOPSYS_UNCONNECTED__542, SYNOPSYS_UNCONNECTED__543, 
        SYNOPSYS_UNCONNECTED__544, SYNOPSYS_UNCONNECTED__545, 
        SYNOPSYS_UNCONNECTED__546, N30514, N30513, N30512, N30511, N30510, 
        N30509}) );
  hamming_N16000_CC4_DW01_add_119 add_1452_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29061, N29060, N29059, N29058, N29057}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29073, N29072, N29071, 
        N29070, N29069}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__547, 
        SYNOPSYS_UNCONNECTED__548, SYNOPSYS_UNCONNECTED__549, 
        SYNOPSYS_UNCONNECTED__550, SYNOPSYS_UNCONNECTED__551, 
        SYNOPSYS_UNCONNECTED__552, N30502, N30501, N30500, N30499, N30498, 
        N30497}) );
  hamming_N16000_CC4_DW01_add_120 add_1453_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29037, N29036, N29035, N29034, N29033}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29049, N29048, N29047, 
        N29046, N29045}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__553, 
        SYNOPSYS_UNCONNECTED__554, SYNOPSYS_UNCONNECTED__555, 
        SYNOPSYS_UNCONNECTED__556, SYNOPSYS_UNCONNECTED__557, 
        SYNOPSYS_UNCONNECTED__558, N30490, N30489, N30488, N30487, N30486, 
        N30485}) );
  hamming_N16000_CC4_DW01_add_121 add_1454_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29013, N29012, N29011, N29010, N29009}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29025, N29024, N29023, 
        N29022, N29021}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__559, 
        SYNOPSYS_UNCONNECTED__560, SYNOPSYS_UNCONNECTED__561, 
        SYNOPSYS_UNCONNECTED__562, SYNOPSYS_UNCONNECTED__563, 
        SYNOPSYS_UNCONNECTED__564, N30478, N30477, N30476, N30475, N30474, 
        N30473}) );
  hamming_N16000_CC4_DW01_add_122 add_1455_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28989, N28988, N28987, N28986, N28985}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29001, N29000, N28999, 
        N28998, N28997}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__565, 
        SYNOPSYS_UNCONNECTED__566, SYNOPSYS_UNCONNECTED__567, 
        SYNOPSYS_UNCONNECTED__568, SYNOPSYS_UNCONNECTED__569, 
        SYNOPSYS_UNCONNECTED__570, N30466, N30465, N30464, N30463, N30462, 
        N30461}) );
  hamming_N16000_CC4_DW01_add_123 add_1456_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28965, N28964, N28963, N28962, N28961}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28977, N28976, N28975, 
        N28974, N28973}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__571, 
        SYNOPSYS_UNCONNECTED__572, SYNOPSYS_UNCONNECTED__573, 
        SYNOPSYS_UNCONNECTED__574, SYNOPSYS_UNCONNECTED__575, 
        SYNOPSYS_UNCONNECTED__576, N30454, N30453, N30452, N30451, N30450, 
        N30449}) );
  hamming_N16000_CC4_DW01_add_124 add_1457_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28941, N28940, N28939, N28938, N28937}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28953, N28952, N28951, 
        N28950, N28949}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__577, 
        SYNOPSYS_UNCONNECTED__578, SYNOPSYS_UNCONNECTED__579, 
        SYNOPSYS_UNCONNECTED__580, SYNOPSYS_UNCONNECTED__581, 
        SYNOPSYS_UNCONNECTED__582, N30442, N30441, N30440, N30439, N30438, 
        N30437}) );
  hamming_N16000_CC4_DW01_add_125 add_1458_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28917, N28916, N28915, N28914, N28913}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28929, N28928, N28927, 
        N28926, N28925}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__583, 
        SYNOPSYS_UNCONNECTED__584, SYNOPSYS_UNCONNECTED__585, 
        SYNOPSYS_UNCONNECTED__586, SYNOPSYS_UNCONNECTED__587, 
        SYNOPSYS_UNCONNECTED__588, N30430, N30429, N30428, N30427, N30426, 
        N30425}) );
  hamming_N16000_CC4_DW01_add_126 add_1459_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28893, N28892, N28891, N28890, N28889}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28905, N28904, N28903, 
        N28902, N28901}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__589, 
        SYNOPSYS_UNCONNECTED__590, SYNOPSYS_UNCONNECTED__591, 
        SYNOPSYS_UNCONNECTED__592, SYNOPSYS_UNCONNECTED__593, 
        SYNOPSYS_UNCONNECTED__594, N30418, N30417, N30416, N30415, N30414, 
        N30413}) );
  hamming_N16000_CC4_DW01_add_127 add_1460_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28869, N28868, N28867, N28866, N28865}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28881, N28880, N28879, 
        N28878, N28877}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__595, 
        SYNOPSYS_UNCONNECTED__596, SYNOPSYS_UNCONNECTED__597, 
        SYNOPSYS_UNCONNECTED__598, SYNOPSYS_UNCONNECTED__599, 
        SYNOPSYS_UNCONNECTED__600, N30406, N30405, N30404, N30403, N30402, 
        N30401}) );
  hamming_N16000_CC4_DW01_add_128 add_1461_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28845, N28844, N28843, N28842, N28841}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28857, N28856, N28855, 
        N28854, N28853}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__601, 
        SYNOPSYS_UNCONNECTED__602, SYNOPSYS_UNCONNECTED__603, 
        SYNOPSYS_UNCONNECTED__604, SYNOPSYS_UNCONNECTED__605, 
        SYNOPSYS_UNCONNECTED__606, N30394, N30393, N30392, N30391, N30390, 
        N30389}) );
  hamming_N16000_CC4_DW01_add_129 add_1462_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28821, N28820, N28819, N28818, N28817}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28833, N28832, N28831, 
        N28830, N28829}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__607, 
        SYNOPSYS_UNCONNECTED__608, SYNOPSYS_UNCONNECTED__609, 
        SYNOPSYS_UNCONNECTED__610, SYNOPSYS_UNCONNECTED__611, 
        SYNOPSYS_UNCONNECTED__612, N30382, N30381, N30380, N30379, N30378, 
        N30377}) );
  hamming_N16000_CC4_DW01_add_130 add_1463_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28797, N28796, N28795, N28794, N28793}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28809, N28808, N28807, 
        N28806, N28805}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__613, 
        SYNOPSYS_UNCONNECTED__614, SYNOPSYS_UNCONNECTED__615, 
        SYNOPSYS_UNCONNECTED__616, SYNOPSYS_UNCONNECTED__617, 
        SYNOPSYS_UNCONNECTED__618, N30370, N30369, N30368, N30367, N30366, 
        N30365}) );
  hamming_N16000_CC4_DW01_add_131 add_1464_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28773, N28772, N28771, N28770, N28769}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28785, N28784, N28783, 
        N28782, N28781}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__619, 
        SYNOPSYS_UNCONNECTED__620, SYNOPSYS_UNCONNECTED__621, 
        SYNOPSYS_UNCONNECTED__622, SYNOPSYS_UNCONNECTED__623, 
        SYNOPSYS_UNCONNECTED__624, N30358, N30357, N30356, N30355, N30354, 
        N30353}) );
  hamming_N16000_CC4_DW01_add_132 add_1465_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28749, N28748, N28747, N28746, N28745}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28761, N28760, N28759, 
        N28758, N28757}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__625, 
        SYNOPSYS_UNCONNECTED__626, SYNOPSYS_UNCONNECTED__627, 
        SYNOPSYS_UNCONNECTED__628, SYNOPSYS_UNCONNECTED__629, 
        SYNOPSYS_UNCONNECTED__630, N30346, N30345, N30344, N30343, N30342, 
        N30341}) );
  hamming_N16000_CC4_DW01_add_133 add_1466_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28725, N28724, N28723, N28722, N28721}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28737, N28736, N28735, 
        N28734, N28733}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__631, 
        SYNOPSYS_UNCONNECTED__632, SYNOPSYS_UNCONNECTED__633, 
        SYNOPSYS_UNCONNECTED__634, SYNOPSYS_UNCONNECTED__635, 
        SYNOPSYS_UNCONNECTED__636, N30334, N30333, N30332, N30331, N30330, 
        N30329}) );
  hamming_N16000_CC4_DW01_add_134 add_1467_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28701, N28700, N28699, N28698, N28697}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28713, N28712, N28711, 
        N28710, N28709}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__637, 
        SYNOPSYS_UNCONNECTED__638, SYNOPSYS_UNCONNECTED__639, 
        SYNOPSYS_UNCONNECTED__640, SYNOPSYS_UNCONNECTED__641, 
        SYNOPSYS_UNCONNECTED__642, N30322, N30321, N30320, N30319, N30318, 
        N30317}) );
  hamming_N16000_CC4_DW01_add_135 add_1468_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28677, N28676, N28675, N28674, N28673}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28689, N28688, N28687, 
        N28686, N28685}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__643, 
        SYNOPSYS_UNCONNECTED__644, SYNOPSYS_UNCONNECTED__645, 
        SYNOPSYS_UNCONNECTED__646, SYNOPSYS_UNCONNECTED__647, 
        SYNOPSYS_UNCONNECTED__648, N30310, N30309, N30308, N30307, N30306, 
        N30305}) );
  hamming_N16000_CC4_DW01_add_136 add_1469_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28653, N28652, N28651, N28650, N28649}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28665, N28664, N28663, 
        N28662, N28661}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__649, 
        SYNOPSYS_UNCONNECTED__650, SYNOPSYS_UNCONNECTED__651, 
        SYNOPSYS_UNCONNECTED__652, SYNOPSYS_UNCONNECTED__653, 
        SYNOPSYS_UNCONNECTED__654, N30298, N30297, N30296, N30295, N30294, 
        N30293}) );
  hamming_N16000_CC4_DW01_add_137 add_1470_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28629, N28628, N28627, N28626, N28625}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28641, N28640, N28639, 
        N28638, N28637}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__655, 
        SYNOPSYS_UNCONNECTED__656, SYNOPSYS_UNCONNECTED__657, 
        SYNOPSYS_UNCONNECTED__658, SYNOPSYS_UNCONNECTED__659, 
        SYNOPSYS_UNCONNECTED__660, N30286, N30285, N30284, N30283, N30282, 
        N30281}) );
  hamming_N16000_CC4_DW01_add_138 add_1471_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28605, N28604, N28603, N28602, N28601}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28617, N28616, N28615, 
        N28614, N28613}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__661, 
        SYNOPSYS_UNCONNECTED__662, SYNOPSYS_UNCONNECTED__663, 
        SYNOPSYS_UNCONNECTED__664, SYNOPSYS_UNCONNECTED__665, 
        SYNOPSYS_UNCONNECTED__666, N30274, N30273, N30272, N30271, N30270, 
        N30269}) );
  hamming_N16000_CC4_DW01_add_139 add_1472_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28581, N28580, N28579, N28578, N28577}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28593, N28592, N28591, 
        N28590, N28589}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__667, 
        SYNOPSYS_UNCONNECTED__668, SYNOPSYS_UNCONNECTED__669, 
        SYNOPSYS_UNCONNECTED__670, SYNOPSYS_UNCONNECTED__671, 
        SYNOPSYS_UNCONNECTED__672, N30262, N30261, N30260, N30259, N30258, 
        N30257}) );
  hamming_N16000_CC4_DW01_add_140 add_1473_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28557, N28556, N28555, N28554, N28553}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28569, N28568, N28567, 
        N28566, N28565}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__673, 
        SYNOPSYS_UNCONNECTED__674, SYNOPSYS_UNCONNECTED__675, 
        SYNOPSYS_UNCONNECTED__676, SYNOPSYS_UNCONNECTED__677, 
        SYNOPSYS_UNCONNECTED__678, N30250, N30249, N30248, N30247, N30246, 
        N30245}) );
  hamming_N16000_CC4_DW01_add_141 add_1474_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28533, N28532, N28531, N28530, N28529}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28545, N28544, N28543, 
        N28542, N28541}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__679, 
        SYNOPSYS_UNCONNECTED__680, SYNOPSYS_UNCONNECTED__681, 
        SYNOPSYS_UNCONNECTED__682, SYNOPSYS_UNCONNECTED__683, 
        SYNOPSYS_UNCONNECTED__684, N30238, N30237, N30236, N30235, N30234, 
        N30233}) );
  hamming_N16000_CC4_DW01_add_142 add_1475_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28509, N28508, N28507, N28506, N28505}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28521, N28520, N28519, 
        N28518, N28517}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__685, 
        SYNOPSYS_UNCONNECTED__686, SYNOPSYS_UNCONNECTED__687, 
        SYNOPSYS_UNCONNECTED__688, SYNOPSYS_UNCONNECTED__689, 
        SYNOPSYS_UNCONNECTED__690, N30226, N30225, N30224, N30223, N30222, 
        N30221}) );
  hamming_N16000_CC4_DW01_add_143 add_1476_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28485, N28484, N28483, N28482, N28481}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28497, N28496, N28495, 
        N28494, N28493}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__691, 
        SYNOPSYS_UNCONNECTED__692, SYNOPSYS_UNCONNECTED__693, 
        SYNOPSYS_UNCONNECTED__694, SYNOPSYS_UNCONNECTED__695, 
        SYNOPSYS_UNCONNECTED__696, N30214, N30213, N30212, N30211, N30210, 
        N30209}) );
  hamming_N16000_CC4_DW01_add_144 add_1477_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28461, N28460, N28459, N28458, N28457}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28473, N28472, N28471, 
        N28470, N28469}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__697, 
        SYNOPSYS_UNCONNECTED__698, SYNOPSYS_UNCONNECTED__699, 
        SYNOPSYS_UNCONNECTED__700, SYNOPSYS_UNCONNECTED__701, 
        SYNOPSYS_UNCONNECTED__702, N30202, N30201, N30200, N30199, N30198, 
        N30197}) );
  hamming_N16000_CC4_DW01_add_145 add_1478_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28437, N28436, N28435, N28434, N28433}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28449, N28448, N28447, 
        N28446, N28445}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__703, 
        SYNOPSYS_UNCONNECTED__704, SYNOPSYS_UNCONNECTED__705, 
        SYNOPSYS_UNCONNECTED__706, SYNOPSYS_UNCONNECTED__707, 
        SYNOPSYS_UNCONNECTED__708, N30190, N30189, N30188, N30187, N30186, 
        N30185}) );
  hamming_N16000_CC4_DW01_add_146 add_1479_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28413, N28412, N28411, N28410, N28409}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28425, N28424, N28423, 
        N28422, N28421}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__709, 
        SYNOPSYS_UNCONNECTED__710, SYNOPSYS_UNCONNECTED__711, 
        SYNOPSYS_UNCONNECTED__712, SYNOPSYS_UNCONNECTED__713, 
        SYNOPSYS_UNCONNECTED__714, N30178, N30177, N30176, N30175, N30174, 
        N30173}) );
  hamming_N16000_CC4_DW01_add_147 add_1480_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28389, N28388, N28387, N28386, N28385}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28401, N28400, N28399, 
        N28398, N28397}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__715, 
        SYNOPSYS_UNCONNECTED__716, SYNOPSYS_UNCONNECTED__717, 
        SYNOPSYS_UNCONNECTED__718, SYNOPSYS_UNCONNECTED__719, 
        SYNOPSYS_UNCONNECTED__720, N30166, N30165, N30164, N30163, N30162, 
        N30161}) );
  hamming_N16000_CC4_DW01_add_148 add_1481_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28365, N28364, N28363, N28362, N28361}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28377, N28376, N28375, 
        N28374, N28373}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__721, 
        SYNOPSYS_UNCONNECTED__722, SYNOPSYS_UNCONNECTED__723, 
        SYNOPSYS_UNCONNECTED__724, SYNOPSYS_UNCONNECTED__725, 
        SYNOPSYS_UNCONNECTED__726, N30154, N30153, N30152, N30151, N30150, 
        N30149}) );
  hamming_N16000_CC4_DW01_add_149 add_1482_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28341, N28340, N28339, N28338, N28337}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28353, N28352, N28351, 
        N28350, N28349}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__727, 
        SYNOPSYS_UNCONNECTED__728, SYNOPSYS_UNCONNECTED__729, 
        SYNOPSYS_UNCONNECTED__730, SYNOPSYS_UNCONNECTED__731, 
        SYNOPSYS_UNCONNECTED__732, N30142, N30141, N30140, N30139, N30138, 
        N30137}) );
  hamming_N16000_CC4_DW01_add_150 add_1483_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28317, N28316, N28315, N28314, N28313}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28329, N28328, N28327, 
        N28326, N28325}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__733, 
        SYNOPSYS_UNCONNECTED__734, SYNOPSYS_UNCONNECTED__735, 
        SYNOPSYS_UNCONNECTED__736, SYNOPSYS_UNCONNECTED__737, 
        SYNOPSYS_UNCONNECTED__738, N30130, N30129, N30128, N30127, N30126, 
        N30125}) );
  hamming_N16000_CC4_DW01_add_151 add_1484_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28293, N28292, N28291, N28290, N28289}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28305, N28304, N28303, 
        N28302, N28301}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__739, 
        SYNOPSYS_UNCONNECTED__740, SYNOPSYS_UNCONNECTED__741, 
        SYNOPSYS_UNCONNECTED__742, SYNOPSYS_UNCONNECTED__743, 
        SYNOPSYS_UNCONNECTED__744, N30118, N30117, N30116, N30115, N30114, 
        N30113}) );
  hamming_N16000_CC4_DW01_add_152 add_1485_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28269, N28268, N28267, N28266, N28265}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28281, N28280, N28279, 
        N28278, N28277}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__745, 
        SYNOPSYS_UNCONNECTED__746, SYNOPSYS_UNCONNECTED__747, 
        SYNOPSYS_UNCONNECTED__748, SYNOPSYS_UNCONNECTED__749, 
        SYNOPSYS_UNCONNECTED__750, N30106, N30105, N30104, N30103, N30102, 
        N30101}) );
  hamming_N16000_CC4_DW01_add_153 add_1486_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28245, N28244, N28243, N28242, N28241}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28257, N28256, N28255, 
        N28254, N28253}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__751, 
        SYNOPSYS_UNCONNECTED__752, SYNOPSYS_UNCONNECTED__753, 
        SYNOPSYS_UNCONNECTED__754, SYNOPSYS_UNCONNECTED__755, 
        SYNOPSYS_UNCONNECTED__756, N30094, N30093, N30092, N30091, N30090, 
        N30089}) );
  hamming_N16000_CC4_DW01_add_154 add_1487_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28221, N28220, N28219, N28218, N28217}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28233, N28232, N28231, 
        N28230, N28229}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__757, 
        SYNOPSYS_UNCONNECTED__758, SYNOPSYS_UNCONNECTED__759, 
        SYNOPSYS_UNCONNECTED__760, SYNOPSYS_UNCONNECTED__761, 
        SYNOPSYS_UNCONNECTED__762, N30082, N30081, N30080, N30079, N30078, 
        N30077}) );
  hamming_N16000_CC4_DW01_add_155 add_1488_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28197, N28196, N28195, N28194, N28193}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28209, N28208, N28207, 
        N28206, N28205}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__763, 
        SYNOPSYS_UNCONNECTED__764, SYNOPSYS_UNCONNECTED__765, 
        SYNOPSYS_UNCONNECTED__766, SYNOPSYS_UNCONNECTED__767, 
        SYNOPSYS_UNCONNECTED__768, N30070, N30069, N30068, N30067, N30066, 
        N30065}) );
  hamming_N16000_CC4_DW01_add_156 add_1489_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28173, N28172, N28171, N28170, N28169}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28185, N28184, N28183, 
        N28182, N28181}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__769, 
        SYNOPSYS_UNCONNECTED__770, SYNOPSYS_UNCONNECTED__771, 
        SYNOPSYS_UNCONNECTED__772, SYNOPSYS_UNCONNECTED__773, 
        SYNOPSYS_UNCONNECTED__774, N30058, N30057, N30056, N30055, N30054, 
        N30053}) );
  hamming_N16000_CC4_DW01_add_157 add_1490_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28149, N28148, N28147, N28146, N28145}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28161, N28160, N28159, 
        N28158, N28157}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__775, 
        SYNOPSYS_UNCONNECTED__776, SYNOPSYS_UNCONNECTED__777, 
        SYNOPSYS_UNCONNECTED__778, SYNOPSYS_UNCONNECTED__779, 
        SYNOPSYS_UNCONNECTED__780, N30046, N30045, N30044, N30043, N30042, 
        N30041}) );
  hamming_N16000_CC4_DW01_add_158 add_1491_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28125, N28124, N28123, N28122, N28121}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28137, N28136, N28135, 
        N28134, N28133}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__781, 
        SYNOPSYS_UNCONNECTED__782, SYNOPSYS_UNCONNECTED__783, 
        SYNOPSYS_UNCONNECTED__784, SYNOPSYS_UNCONNECTED__785, 
        SYNOPSYS_UNCONNECTED__786, N30034, N30033, N30032, N30031, N30030, 
        N30029}) );
  hamming_N16000_CC4_DW01_add_159 add_1492_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28101, N28100, N28099, N28098, N28097}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28113, N28112, N28111, 
        N28110, N28109}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__787, 
        SYNOPSYS_UNCONNECTED__788, SYNOPSYS_UNCONNECTED__789, 
        SYNOPSYS_UNCONNECTED__790, SYNOPSYS_UNCONNECTED__791, 
        SYNOPSYS_UNCONNECTED__792, N30022, N30021, N30020, N30019, N30018, 
        N30017}) );
  hamming_N16000_CC4_DW01_add_160 add_1493_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28077, N28076, N28075, N28074, N28073}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28089, N28088, N28087, 
        N28086, N28085}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__793, 
        SYNOPSYS_UNCONNECTED__794, SYNOPSYS_UNCONNECTED__795, 
        SYNOPSYS_UNCONNECTED__796, SYNOPSYS_UNCONNECTED__797, 
        SYNOPSYS_UNCONNECTED__798, N30010, N30009, N30008, N30007, N30006, 
        N30005}) );
  hamming_N16000_CC4_DW01_add_161 add_1494_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28053, N28052, N28051, N28050, N28049}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28065, N28064, N28063, 
        N28062, N28061}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__799, 
        SYNOPSYS_UNCONNECTED__800, SYNOPSYS_UNCONNECTED__801, 
        SYNOPSYS_UNCONNECTED__802, SYNOPSYS_UNCONNECTED__803, 
        SYNOPSYS_UNCONNECTED__804, N29998, N29997, N29996, N29995, N29994, 
        N29993}) );
  hamming_N16000_CC4_DW01_add_162 add_1495_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28029, N28028, N28027, N28026, N28025}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28041, N28040, N28039, 
        N28038, N28037}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__805, 
        SYNOPSYS_UNCONNECTED__806, SYNOPSYS_UNCONNECTED__807, 
        SYNOPSYS_UNCONNECTED__808, SYNOPSYS_UNCONNECTED__809, 
        SYNOPSYS_UNCONNECTED__810, N29986, N29985, N29984, N29983, N29982, 
        N29981}) );
  hamming_N16000_CC4_DW01_add_163 add_1496_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28005, N28004, N28003, N28002, N28001}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28017, N28016, N28015, 
        N28014, N28013}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__811, 
        SYNOPSYS_UNCONNECTED__812, SYNOPSYS_UNCONNECTED__813, 
        SYNOPSYS_UNCONNECTED__814, SYNOPSYS_UNCONNECTED__815, 
        SYNOPSYS_UNCONNECTED__816, N29974, N29973, N29972, N29971, N29970, 
        N29969}) );
  hamming_N16000_CC4_DW01_add_164 add_1497_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N27981, N27980, N27979, N27978, N27977}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N27993, N27992, N27991, 
        N27990, N27989}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__817, 
        SYNOPSYS_UNCONNECTED__818, SYNOPSYS_UNCONNECTED__819, 
        SYNOPSYS_UNCONNECTED__820, SYNOPSYS_UNCONNECTED__821, 
        SYNOPSYS_UNCONNECTED__822, N29962, N29961, N29960, N29959, N29958, 
        N29957}) );
  hamming_N16000_CC4_DW01_add_165 add_1498_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N27957, N27956, N27955, N27954, N27953}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N27969, N27968, N27967, 
        N27966, N27965}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__823, 
        SYNOPSYS_UNCONNECTED__824, SYNOPSYS_UNCONNECTED__825, 
        SYNOPSYS_UNCONNECTED__826, SYNOPSYS_UNCONNECTED__827, 
        SYNOPSYS_UNCONNECTED__828, N29950, N29949, N29948, N29947, N29946, 
        N29945}) );
  hamming_N16000_CC4_DW01_add_166 add_1499_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N27933, N27932, N27931, N27930, N27929}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N27945, N27944, N27943, 
        N27942, N27941}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__829, 
        SYNOPSYS_UNCONNECTED__830, SYNOPSYS_UNCONNECTED__831, 
        SYNOPSYS_UNCONNECTED__832, SYNOPSYS_UNCONNECTED__833, 
        SYNOPSYS_UNCONNECTED__834, N29938, N29937, N29936, N29935, N29934, 
        N29933}) );
  NAND U6686 ( .A(n2687), .B(n2688), .Z(N29925) );
  NANDN U6687 ( .A(n2689), .B(n2690), .Z(n2688) );
  OR U6688 ( .A(n2691), .B(n2692), .Z(n2690) );
  NAND U6689 ( .A(n2691), .B(n2692), .Z(n2687) );
  XOR U6690 ( .A(n2691), .B(n2693), .Z(N29924) );
  XNOR U6691 ( .A(n2689), .B(n2692), .Z(n2693) );
  AND U6692 ( .A(n2694), .B(n2695), .Z(n2692) );
  NANDN U6693 ( .A(n2696), .B(n2697), .Z(n2695) );
  NANDN U6694 ( .A(n2698), .B(n2699), .Z(n2697) );
  NANDN U6695 ( .A(n2699), .B(n2698), .Z(n2694) );
  NAND U6696 ( .A(n2700), .B(n2701), .Z(n2689) );
  NANDN U6697 ( .A(n2702), .B(n2703), .Z(n2701) );
  OR U6698 ( .A(n2704), .B(n2705), .Z(n2703) );
  NAND U6699 ( .A(n2705), .B(n2704), .Z(n2700) );
  AND U6700 ( .A(n2706), .B(n2707), .Z(n2691) );
  NANDN U6701 ( .A(n2708), .B(n2709), .Z(n2707) );
  NANDN U6702 ( .A(n2710), .B(n2711), .Z(n2709) );
  NANDN U6703 ( .A(n2711), .B(n2710), .Z(n2706) );
  XOR U6704 ( .A(n2705), .B(n2712), .Z(N29923) );
  XOR U6705 ( .A(n2702), .B(n2704), .Z(n2712) );
  XNOR U6706 ( .A(n2698), .B(n2713), .Z(n2704) );
  XNOR U6707 ( .A(n2696), .B(n2699), .Z(n2713) );
  NAND U6708 ( .A(n2714), .B(n2715), .Z(n2699) );
  NAND U6709 ( .A(n2716), .B(n2717), .Z(n2715) );
  OR U6710 ( .A(n2718), .B(n2719), .Z(n2716) );
  NANDN U6711 ( .A(n2720), .B(n2718), .Z(n2714) );
  IV U6712 ( .A(n2719), .Z(n2720) );
  NAND U6713 ( .A(n2721), .B(n2722), .Z(n2696) );
  NAND U6714 ( .A(n2723), .B(n2724), .Z(n2722) );
  NANDN U6715 ( .A(n2725), .B(n2726), .Z(n2723) );
  NANDN U6716 ( .A(n2726), .B(n2725), .Z(n2721) );
  AND U6717 ( .A(n2727), .B(n2728), .Z(n2698) );
  NAND U6718 ( .A(n2729), .B(n2730), .Z(n2728) );
  OR U6719 ( .A(n2731), .B(n2732), .Z(n2729) );
  NANDN U6720 ( .A(n2733), .B(n2731), .Z(n2727) );
  NAND U6721 ( .A(n2734), .B(n2735), .Z(n2702) );
  NANDN U6722 ( .A(n2736), .B(n2737), .Z(n2735) );
  OR U6723 ( .A(n2738), .B(n2739), .Z(n2737) );
  NANDN U6724 ( .A(n2740), .B(n2738), .Z(n2734) );
  IV U6725 ( .A(n2739), .Z(n2740) );
  XNOR U6726 ( .A(n2710), .B(n2741), .Z(n2705) );
  XNOR U6727 ( .A(n2708), .B(n2711), .Z(n2741) );
  NAND U6728 ( .A(n2742), .B(n2743), .Z(n2711) );
  NAND U6729 ( .A(n2744), .B(n2745), .Z(n2743) );
  OR U6730 ( .A(n2746), .B(n2747), .Z(n2744) );
  NANDN U6731 ( .A(n2748), .B(n2746), .Z(n2742) );
  IV U6732 ( .A(n2747), .Z(n2748) );
  NAND U6733 ( .A(n2749), .B(n2750), .Z(n2708) );
  NAND U6734 ( .A(n2751), .B(n2752), .Z(n2750) );
  NANDN U6735 ( .A(n2753), .B(n2754), .Z(n2751) );
  NANDN U6736 ( .A(n2754), .B(n2753), .Z(n2749) );
  AND U6737 ( .A(n2755), .B(n2756), .Z(n2710) );
  NAND U6738 ( .A(n2757), .B(n2758), .Z(n2756) );
  OR U6739 ( .A(n2759), .B(n2760), .Z(n2757) );
  NANDN U6740 ( .A(n2761), .B(n2759), .Z(n2755) );
  XNOR U6741 ( .A(n2736), .B(n2762), .Z(N29922) );
  XOR U6742 ( .A(n2738), .B(n2739), .Z(n2762) );
  XNOR U6743 ( .A(n2752), .B(n2763), .Z(n2739) );
  XOR U6744 ( .A(n2753), .B(n2754), .Z(n2763) );
  XOR U6745 ( .A(n2759), .B(n2764), .Z(n2754) );
  XOR U6746 ( .A(n2758), .B(n2761), .Z(n2764) );
  IV U6747 ( .A(n2760), .Z(n2761) );
  NAND U6748 ( .A(n2765), .B(n2766), .Z(n2760) );
  OR U6749 ( .A(n2767), .B(n2768), .Z(n2766) );
  OR U6750 ( .A(n2769), .B(n2770), .Z(n2765) );
  NAND U6751 ( .A(n2771), .B(n2772), .Z(n2758) );
  OR U6752 ( .A(n2773), .B(n2774), .Z(n2772) );
  OR U6753 ( .A(n2775), .B(n2776), .Z(n2771) );
  NOR U6754 ( .A(n2777), .B(n2778), .Z(n2759) );
  ANDN U6755 ( .B(n2779), .A(n2780), .Z(n2753) );
  XNOR U6756 ( .A(n2746), .B(n2781), .Z(n2752) );
  XNOR U6757 ( .A(n2745), .B(n2747), .Z(n2781) );
  NAND U6758 ( .A(n2782), .B(n2783), .Z(n2747) );
  OR U6759 ( .A(n2784), .B(n2785), .Z(n2783) );
  OR U6760 ( .A(n2786), .B(n2787), .Z(n2782) );
  NAND U6761 ( .A(n2788), .B(n2789), .Z(n2745) );
  OR U6762 ( .A(n2790), .B(n2791), .Z(n2789) );
  OR U6763 ( .A(n2792), .B(n2793), .Z(n2788) );
  ANDN U6764 ( .B(n2794), .A(n2795), .Z(n2746) );
  IV U6765 ( .A(n2796), .Z(n2794) );
  ANDN U6766 ( .B(n2797), .A(n2798), .Z(n2738) );
  XOR U6767 ( .A(n2724), .B(n2799), .Z(n2736) );
  XOR U6768 ( .A(n2725), .B(n2726), .Z(n2799) );
  XOR U6769 ( .A(n2731), .B(n2800), .Z(n2726) );
  XOR U6770 ( .A(n2730), .B(n2733), .Z(n2800) );
  IV U6771 ( .A(n2732), .Z(n2733) );
  NAND U6772 ( .A(n2801), .B(n2802), .Z(n2732) );
  OR U6773 ( .A(n2803), .B(n2804), .Z(n2802) );
  OR U6774 ( .A(n2805), .B(n2806), .Z(n2801) );
  NAND U6775 ( .A(n2807), .B(n2808), .Z(n2730) );
  OR U6776 ( .A(n2809), .B(n2810), .Z(n2808) );
  OR U6777 ( .A(n2811), .B(n2812), .Z(n2807) );
  NOR U6778 ( .A(n2813), .B(n2814), .Z(n2731) );
  ANDN U6779 ( .B(n2815), .A(n2816), .Z(n2725) );
  IV U6780 ( .A(n2817), .Z(n2815) );
  XNOR U6781 ( .A(n2718), .B(n2818), .Z(n2724) );
  XNOR U6782 ( .A(n2717), .B(n2719), .Z(n2818) );
  NAND U6783 ( .A(n2819), .B(n2820), .Z(n2719) );
  OR U6784 ( .A(n2821), .B(n2822), .Z(n2820) );
  OR U6785 ( .A(n2823), .B(n2824), .Z(n2819) );
  NAND U6786 ( .A(n2825), .B(n2826), .Z(n2717) );
  OR U6787 ( .A(n2827), .B(n2828), .Z(n2826) );
  OR U6788 ( .A(n2829), .B(n2830), .Z(n2825) );
  ANDN U6789 ( .B(n2831), .A(n2832), .Z(n2718) );
  IV U6790 ( .A(n2833), .Z(n2831) );
  XNOR U6791 ( .A(n2798), .B(n2797), .Z(N29921) );
  XOR U6792 ( .A(n2817), .B(n2816), .Z(n2797) );
  XNOR U6793 ( .A(n2832), .B(n2833), .Z(n2816) );
  XNOR U6794 ( .A(n2827), .B(n2828), .Z(n2833) );
  XNOR U6795 ( .A(n2829), .B(n2830), .Z(n2828) );
  XNOR U6796 ( .A(y[3988]), .B(x[3988]), .Z(n2830) );
  XNOR U6797 ( .A(y[3989]), .B(x[3989]), .Z(n2829) );
  XNOR U6798 ( .A(y[3987]), .B(x[3987]), .Z(n2827) );
  XNOR U6799 ( .A(n2821), .B(n2822), .Z(n2832) );
  XNOR U6800 ( .A(y[3984]), .B(x[3984]), .Z(n2822) );
  XNOR U6801 ( .A(n2823), .B(n2824), .Z(n2821) );
  XNOR U6802 ( .A(y[3985]), .B(x[3985]), .Z(n2824) );
  XNOR U6803 ( .A(y[3986]), .B(x[3986]), .Z(n2823) );
  XNOR U6804 ( .A(n2814), .B(n2813), .Z(n2817) );
  XNOR U6805 ( .A(n2809), .B(n2810), .Z(n2813) );
  XNOR U6806 ( .A(y[3981]), .B(x[3981]), .Z(n2810) );
  XNOR U6807 ( .A(n2811), .B(n2812), .Z(n2809) );
  XNOR U6808 ( .A(y[3982]), .B(x[3982]), .Z(n2812) );
  XNOR U6809 ( .A(y[3983]), .B(x[3983]), .Z(n2811) );
  XNOR U6810 ( .A(n2803), .B(n2804), .Z(n2814) );
  XNOR U6811 ( .A(y[3978]), .B(x[3978]), .Z(n2804) );
  XNOR U6812 ( .A(n2805), .B(n2806), .Z(n2803) );
  XNOR U6813 ( .A(y[3979]), .B(x[3979]), .Z(n2806) );
  XNOR U6814 ( .A(y[3980]), .B(x[3980]), .Z(n2805) );
  XOR U6815 ( .A(n2779), .B(n2780), .Z(n2798) );
  XNOR U6816 ( .A(n2795), .B(n2796), .Z(n2780) );
  XNOR U6817 ( .A(n2790), .B(n2791), .Z(n2796) );
  XNOR U6818 ( .A(n2792), .B(n2793), .Z(n2791) );
  XNOR U6819 ( .A(y[3976]), .B(x[3976]), .Z(n2793) );
  XNOR U6820 ( .A(y[3977]), .B(x[3977]), .Z(n2792) );
  XNOR U6821 ( .A(y[3975]), .B(x[3975]), .Z(n2790) );
  XNOR U6822 ( .A(n2784), .B(n2785), .Z(n2795) );
  XNOR U6823 ( .A(y[3972]), .B(x[3972]), .Z(n2785) );
  XNOR U6824 ( .A(n2786), .B(n2787), .Z(n2784) );
  XNOR U6825 ( .A(y[3973]), .B(x[3973]), .Z(n2787) );
  XNOR U6826 ( .A(y[3974]), .B(x[3974]), .Z(n2786) );
  XOR U6827 ( .A(n2778), .B(n2777), .Z(n2779) );
  XNOR U6828 ( .A(n2773), .B(n2774), .Z(n2777) );
  XNOR U6829 ( .A(y[3969]), .B(x[3969]), .Z(n2774) );
  XNOR U6830 ( .A(n2775), .B(n2776), .Z(n2773) );
  XNOR U6831 ( .A(y[3970]), .B(x[3970]), .Z(n2776) );
  XNOR U6832 ( .A(y[3971]), .B(x[3971]), .Z(n2775) );
  XNOR U6833 ( .A(n2767), .B(n2768), .Z(n2778) );
  XNOR U6834 ( .A(y[3966]), .B(x[3966]), .Z(n2768) );
  XNOR U6835 ( .A(n2769), .B(n2770), .Z(n2767) );
  XNOR U6836 ( .A(y[3967]), .B(x[3967]), .Z(n2770) );
  XNOR U6837 ( .A(y[3968]), .B(x[3968]), .Z(n2769) );
  NAND U6838 ( .A(n2834), .B(n2835), .Z(N29913) );
  NANDN U6839 ( .A(n2836), .B(n2837), .Z(n2835) );
  OR U6840 ( .A(n2838), .B(n2839), .Z(n2837) );
  NAND U6841 ( .A(n2838), .B(n2839), .Z(n2834) );
  XOR U6842 ( .A(n2838), .B(n2840), .Z(N29912) );
  XNOR U6843 ( .A(n2836), .B(n2839), .Z(n2840) );
  AND U6844 ( .A(n2841), .B(n2842), .Z(n2839) );
  NANDN U6845 ( .A(n2843), .B(n2844), .Z(n2842) );
  NANDN U6846 ( .A(n2845), .B(n2846), .Z(n2844) );
  NANDN U6847 ( .A(n2846), .B(n2845), .Z(n2841) );
  NAND U6848 ( .A(n2847), .B(n2848), .Z(n2836) );
  NANDN U6849 ( .A(n2849), .B(n2850), .Z(n2848) );
  OR U6850 ( .A(n2851), .B(n2852), .Z(n2850) );
  NAND U6851 ( .A(n2852), .B(n2851), .Z(n2847) );
  AND U6852 ( .A(n2853), .B(n2854), .Z(n2838) );
  NANDN U6853 ( .A(n2855), .B(n2856), .Z(n2854) );
  NANDN U6854 ( .A(n2857), .B(n2858), .Z(n2856) );
  NANDN U6855 ( .A(n2858), .B(n2857), .Z(n2853) );
  XOR U6856 ( .A(n2852), .B(n2859), .Z(N29911) );
  XOR U6857 ( .A(n2849), .B(n2851), .Z(n2859) );
  XNOR U6858 ( .A(n2845), .B(n2860), .Z(n2851) );
  XNOR U6859 ( .A(n2843), .B(n2846), .Z(n2860) );
  NAND U6860 ( .A(n2861), .B(n2862), .Z(n2846) );
  NAND U6861 ( .A(n2863), .B(n2864), .Z(n2862) );
  OR U6862 ( .A(n2865), .B(n2866), .Z(n2863) );
  NANDN U6863 ( .A(n2867), .B(n2865), .Z(n2861) );
  IV U6864 ( .A(n2866), .Z(n2867) );
  NAND U6865 ( .A(n2868), .B(n2869), .Z(n2843) );
  NAND U6866 ( .A(n2870), .B(n2871), .Z(n2869) );
  NANDN U6867 ( .A(n2872), .B(n2873), .Z(n2870) );
  NANDN U6868 ( .A(n2873), .B(n2872), .Z(n2868) );
  AND U6869 ( .A(n2874), .B(n2875), .Z(n2845) );
  NAND U6870 ( .A(n2876), .B(n2877), .Z(n2875) );
  OR U6871 ( .A(n2878), .B(n2879), .Z(n2876) );
  NANDN U6872 ( .A(n2880), .B(n2878), .Z(n2874) );
  NAND U6873 ( .A(n2881), .B(n2882), .Z(n2849) );
  NANDN U6874 ( .A(n2883), .B(n2884), .Z(n2882) );
  OR U6875 ( .A(n2885), .B(n2886), .Z(n2884) );
  NANDN U6876 ( .A(n2887), .B(n2885), .Z(n2881) );
  IV U6877 ( .A(n2886), .Z(n2887) );
  XNOR U6878 ( .A(n2857), .B(n2888), .Z(n2852) );
  XNOR U6879 ( .A(n2855), .B(n2858), .Z(n2888) );
  NAND U6880 ( .A(n2889), .B(n2890), .Z(n2858) );
  NAND U6881 ( .A(n2891), .B(n2892), .Z(n2890) );
  OR U6882 ( .A(n2893), .B(n2894), .Z(n2891) );
  NANDN U6883 ( .A(n2895), .B(n2893), .Z(n2889) );
  IV U6884 ( .A(n2894), .Z(n2895) );
  NAND U6885 ( .A(n2896), .B(n2897), .Z(n2855) );
  NAND U6886 ( .A(n2898), .B(n2899), .Z(n2897) );
  NANDN U6887 ( .A(n2900), .B(n2901), .Z(n2898) );
  NANDN U6888 ( .A(n2901), .B(n2900), .Z(n2896) );
  AND U6889 ( .A(n2902), .B(n2903), .Z(n2857) );
  NAND U6890 ( .A(n2904), .B(n2905), .Z(n2903) );
  OR U6891 ( .A(n2906), .B(n2907), .Z(n2904) );
  NANDN U6892 ( .A(n2908), .B(n2906), .Z(n2902) );
  XNOR U6893 ( .A(n2883), .B(n2909), .Z(N29910) );
  XOR U6894 ( .A(n2885), .B(n2886), .Z(n2909) );
  XNOR U6895 ( .A(n2899), .B(n2910), .Z(n2886) );
  XOR U6896 ( .A(n2900), .B(n2901), .Z(n2910) );
  XOR U6897 ( .A(n2906), .B(n2911), .Z(n2901) );
  XOR U6898 ( .A(n2905), .B(n2908), .Z(n2911) );
  IV U6899 ( .A(n2907), .Z(n2908) );
  NAND U6900 ( .A(n2912), .B(n2913), .Z(n2907) );
  OR U6901 ( .A(n2914), .B(n2915), .Z(n2913) );
  OR U6902 ( .A(n2916), .B(n2917), .Z(n2912) );
  NAND U6903 ( .A(n2918), .B(n2919), .Z(n2905) );
  OR U6904 ( .A(n2920), .B(n2921), .Z(n2919) );
  OR U6905 ( .A(n2922), .B(n2923), .Z(n2918) );
  NOR U6906 ( .A(n2924), .B(n2925), .Z(n2906) );
  ANDN U6907 ( .B(n2926), .A(n2927), .Z(n2900) );
  XNOR U6908 ( .A(n2893), .B(n2928), .Z(n2899) );
  XNOR U6909 ( .A(n2892), .B(n2894), .Z(n2928) );
  NAND U6910 ( .A(n2929), .B(n2930), .Z(n2894) );
  OR U6911 ( .A(n2931), .B(n2932), .Z(n2930) );
  OR U6912 ( .A(n2933), .B(n2934), .Z(n2929) );
  NAND U6913 ( .A(n2935), .B(n2936), .Z(n2892) );
  OR U6914 ( .A(n2937), .B(n2938), .Z(n2936) );
  OR U6915 ( .A(n2939), .B(n2940), .Z(n2935) );
  ANDN U6916 ( .B(n2941), .A(n2942), .Z(n2893) );
  IV U6917 ( .A(n2943), .Z(n2941) );
  ANDN U6918 ( .B(n2944), .A(n2945), .Z(n2885) );
  XOR U6919 ( .A(n2871), .B(n2946), .Z(n2883) );
  XOR U6920 ( .A(n2872), .B(n2873), .Z(n2946) );
  XOR U6921 ( .A(n2878), .B(n2947), .Z(n2873) );
  XOR U6922 ( .A(n2877), .B(n2880), .Z(n2947) );
  IV U6923 ( .A(n2879), .Z(n2880) );
  NAND U6924 ( .A(n2948), .B(n2949), .Z(n2879) );
  OR U6925 ( .A(n2950), .B(n2951), .Z(n2949) );
  OR U6926 ( .A(n2952), .B(n2953), .Z(n2948) );
  NAND U6927 ( .A(n2954), .B(n2955), .Z(n2877) );
  OR U6928 ( .A(n2956), .B(n2957), .Z(n2955) );
  OR U6929 ( .A(n2958), .B(n2959), .Z(n2954) );
  NOR U6930 ( .A(n2960), .B(n2961), .Z(n2878) );
  ANDN U6931 ( .B(n2962), .A(n2963), .Z(n2872) );
  IV U6932 ( .A(n2964), .Z(n2962) );
  XNOR U6933 ( .A(n2865), .B(n2965), .Z(n2871) );
  XNOR U6934 ( .A(n2864), .B(n2866), .Z(n2965) );
  NAND U6935 ( .A(n2966), .B(n2967), .Z(n2866) );
  OR U6936 ( .A(n2968), .B(n2969), .Z(n2967) );
  OR U6937 ( .A(n2970), .B(n2971), .Z(n2966) );
  NAND U6938 ( .A(n2972), .B(n2973), .Z(n2864) );
  OR U6939 ( .A(n2974), .B(n2975), .Z(n2973) );
  OR U6940 ( .A(n2976), .B(n2977), .Z(n2972) );
  ANDN U6941 ( .B(n2978), .A(n2979), .Z(n2865) );
  IV U6942 ( .A(n2980), .Z(n2978) );
  XNOR U6943 ( .A(n2945), .B(n2944), .Z(N29909) );
  XOR U6944 ( .A(n2964), .B(n2963), .Z(n2944) );
  XNOR U6945 ( .A(n2979), .B(n2980), .Z(n2963) );
  XNOR U6946 ( .A(n2974), .B(n2975), .Z(n2980) );
  XNOR U6947 ( .A(n2976), .B(n2977), .Z(n2975) );
  XNOR U6948 ( .A(y[3964]), .B(x[3964]), .Z(n2977) );
  XNOR U6949 ( .A(y[3965]), .B(x[3965]), .Z(n2976) );
  XNOR U6950 ( .A(y[3963]), .B(x[3963]), .Z(n2974) );
  XNOR U6951 ( .A(n2968), .B(n2969), .Z(n2979) );
  XNOR U6952 ( .A(y[3960]), .B(x[3960]), .Z(n2969) );
  XNOR U6953 ( .A(n2970), .B(n2971), .Z(n2968) );
  XNOR U6954 ( .A(y[3961]), .B(x[3961]), .Z(n2971) );
  XNOR U6955 ( .A(y[3962]), .B(x[3962]), .Z(n2970) );
  XNOR U6956 ( .A(n2961), .B(n2960), .Z(n2964) );
  XNOR U6957 ( .A(n2956), .B(n2957), .Z(n2960) );
  XNOR U6958 ( .A(y[3957]), .B(x[3957]), .Z(n2957) );
  XNOR U6959 ( .A(n2958), .B(n2959), .Z(n2956) );
  XNOR U6960 ( .A(y[3958]), .B(x[3958]), .Z(n2959) );
  XNOR U6961 ( .A(y[3959]), .B(x[3959]), .Z(n2958) );
  XNOR U6962 ( .A(n2950), .B(n2951), .Z(n2961) );
  XNOR U6963 ( .A(y[3954]), .B(x[3954]), .Z(n2951) );
  XNOR U6964 ( .A(n2952), .B(n2953), .Z(n2950) );
  XNOR U6965 ( .A(y[3955]), .B(x[3955]), .Z(n2953) );
  XNOR U6966 ( .A(y[3956]), .B(x[3956]), .Z(n2952) );
  XOR U6967 ( .A(n2926), .B(n2927), .Z(n2945) );
  XNOR U6968 ( .A(n2942), .B(n2943), .Z(n2927) );
  XNOR U6969 ( .A(n2937), .B(n2938), .Z(n2943) );
  XNOR U6970 ( .A(n2939), .B(n2940), .Z(n2938) );
  XNOR U6971 ( .A(y[3952]), .B(x[3952]), .Z(n2940) );
  XNOR U6972 ( .A(y[3953]), .B(x[3953]), .Z(n2939) );
  XNOR U6973 ( .A(y[3951]), .B(x[3951]), .Z(n2937) );
  XNOR U6974 ( .A(n2931), .B(n2932), .Z(n2942) );
  XNOR U6975 ( .A(y[3948]), .B(x[3948]), .Z(n2932) );
  XNOR U6976 ( .A(n2933), .B(n2934), .Z(n2931) );
  XNOR U6977 ( .A(y[3949]), .B(x[3949]), .Z(n2934) );
  XNOR U6978 ( .A(y[3950]), .B(x[3950]), .Z(n2933) );
  XOR U6979 ( .A(n2925), .B(n2924), .Z(n2926) );
  XNOR U6980 ( .A(n2920), .B(n2921), .Z(n2924) );
  XNOR U6981 ( .A(y[3945]), .B(x[3945]), .Z(n2921) );
  XNOR U6982 ( .A(n2922), .B(n2923), .Z(n2920) );
  XNOR U6983 ( .A(y[3946]), .B(x[3946]), .Z(n2923) );
  XNOR U6984 ( .A(y[3947]), .B(x[3947]), .Z(n2922) );
  XNOR U6985 ( .A(n2914), .B(n2915), .Z(n2925) );
  XNOR U6986 ( .A(y[3942]), .B(x[3942]), .Z(n2915) );
  XNOR U6987 ( .A(n2916), .B(n2917), .Z(n2914) );
  XNOR U6988 ( .A(y[3943]), .B(x[3943]), .Z(n2917) );
  XNOR U6989 ( .A(y[3944]), .B(x[3944]), .Z(n2916) );
  NAND U6990 ( .A(n2981), .B(n2982), .Z(N29901) );
  NANDN U6991 ( .A(n2983), .B(n2984), .Z(n2982) );
  OR U6992 ( .A(n2985), .B(n2986), .Z(n2984) );
  NAND U6993 ( .A(n2985), .B(n2986), .Z(n2981) );
  XOR U6994 ( .A(n2985), .B(n2987), .Z(N29900) );
  XNOR U6995 ( .A(n2983), .B(n2986), .Z(n2987) );
  AND U6996 ( .A(n2988), .B(n2989), .Z(n2986) );
  NANDN U6997 ( .A(n2990), .B(n2991), .Z(n2989) );
  NANDN U6998 ( .A(n2992), .B(n2993), .Z(n2991) );
  NANDN U6999 ( .A(n2993), .B(n2992), .Z(n2988) );
  NAND U7000 ( .A(n2994), .B(n2995), .Z(n2983) );
  NANDN U7001 ( .A(n2996), .B(n2997), .Z(n2995) );
  OR U7002 ( .A(n2998), .B(n2999), .Z(n2997) );
  NAND U7003 ( .A(n2999), .B(n2998), .Z(n2994) );
  AND U7004 ( .A(n3000), .B(n3001), .Z(n2985) );
  NANDN U7005 ( .A(n3002), .B(n3003), .Z(n3001) );
  NANDN U7006 ( .A(n3004), .B(n3005), .Z(n3003) );
  NANDN U7007 ( .A(n3005), .B(n3004), .Z(n3000) );
  XOR U7008 ( .A(n2999), .B(n3006), .Z(N29899) );
  XOR U7009 ( .A(n2996), .B(n2998), .Z(n3006) );
  XNOR U7010 ( .A(n2992), .B(n3007), .Z(n2998) );
  XNOR U7011 ( .A(n2990), .B(n2993), .Z(n3007) );
  NAND U7012 ( .A(n3008), .B(n3009), .Z(n2993) );
  NAND U7013 ( .A(n3010), .B(n3011), .Z(n3009) );
  OR U7014 ( .A(n3012), .B(n3013), .Z(n3010) );
  NANDN U7015 ( .A(n3014), .B(n3012), .Z(n3008) );
  IV U7016 ( .A(n3013), .Z(n3014) );
  NAND U7017 ( .A(n3015), .B(n3016), .Z(n2990) );
  NAND U7018 ( .A(n3017), .B(n3018), .Z(n3016) );
  NANDN U7019 ( .A(n3019), .B(n3020), .Z(n3017) );
  NANDN U7020 ( .A(n3020), .B(n3019), .Z(n3015) );
  AND U7021 ( .A(n3021), .B(n3022), .Z(n2992) );
  NAND U7022 ( .A(n3023), .B(n3024), .Z(n3022) );
  OR U7023 ( .A(n3025), .B(n3026), .Z(n3023) );
  NANDN U7024 ( .A(n3027), .B(n3025), .Z(n3021) );
  NAND U7025 ( .A(n3028), .B(n3029), .Z(n2996) );
  NANDN U7026 ( .A(n3030), .B(n3031), .Z(n3029) );
  OR U7027 ( .A(n3032), .B(n3033), .Z(n3031) );
  NANDN U7028 ( .A(n3034), .B(n3032), .Z(n3028) );
  IV U7029 ( .A(n3033), .Z(n3034) );
  XNOR U7030 ( .A(n3004), .B(n3035), .Z(n2999) );
  XNOR U7031 ( .A(n3002), .B(n3005), .Z(n3035) );
  NAND U7032 ( .A(n3036), .B(n3037), .Z(n3005) );
  NAND U7033 ( .A(n3038), .B(n3039), .Z(n3037) );
  OR U7034 ( .A(n3040), .B(n3041), .Z(n3038) );
  NANDN U7035 ( .A(n3042), .B(n3040), .Z(n3036) );
  IV U7036 ( .A(n3041), .Z(n3042) );
  NAND U7037 ( .A(n3043), .B(n3044), .Z(n3002) );
  NAND U7038 ( .A(n3045), .B(n3046), .Z(n3044) );
  NANDN U7039 ( .A(n3047), .B(n3048), .Z(n3045) );
  NANDN U7040 ( .A(n3048), .B(n3047), .Z(n3043) );
  AND U7041 ( .A(n3049), .B(n3050), .Z(n3004) );
  NAND U7042 ( .A(n3051), .B(n3052), .Z(n3050) );
  OR U7043 ( .A(n3053), .B(n3054), .Z(n3051) );
  NANDN U7044 ( .A(n3055), .B(n3053), .Z(n3049) );
  XNOR U7045 ( .A(n3030), .B(n3056), .Z(N29898) );
  XOR U7046 ( .A(n3032), .B(n3033), .Z(n3056) );
  XNOR U7047 ( .A(n3046), .B(n3057), .Z(n3033) );
  XOR U7048 ( .A(n3047), .B(n3048), .Z(n3057) );
  XOR U7049 ( .A(n3053), .B(n3058), .Z(n3048) );
  XOR U7050 ( .A(n3052), .B(n3055), .Z(n3058) );
  IV U7051 ( .A(n3054), .Z(n3055) );
  NAND U7052 ( .A(n3059), .B(n3060), .Z(n3054) );
  OR U7053 ( .A(n3061), .B(n3062), .Z(n3060) );
  OR U7054 ( .A(n3063), .B(n3064), .Z(n3059) );
  NAND U7055 ( .A(n3065), .B(n3066), .Z(n3052) );
  OR U7056 ( .A(n3067), .B(n3068), .Z(n3066) );
  OR U7057 ( .A(n3069), .B(n3070), .Z(n3065) );
  NOR U7058 ( .A(n3071), .B(n3072), .Z(n3053) );
  ANDN U7059 ( .B(n3073), .A(n3074), .Z(n3047) );
  XNOR U7060 ( .A(n3040), .B(n3075), .Z(n3046) );
  XNOR U7061 ( .A(n3039), .B(n3041), .Z(n3075) );
  NAND U7062 ( .A(n3076), .B(n3077), .Z(n3041) );
  OR U7063 ( .A(n3078), .B(n3079), .Z(n3077) );
  OR U7064 ( .A(n3080), .B(n3081), .Z(n3076) );
  NAND U7065 ( .A(n3082), .B(n3083), .Z(n3039) );
  OR U7066 ( .A(n3084), .B(n3085), .Z(n3083) );
  OR U7067 ( .A(n3086), .B(n3087), .Z(n3082) );
  ANDN U7068 ( .B(n3088), .A(n3089), .Z(n3040) );
  IV U7069 ( .A(n3090), .Z(n3088) );
  ANDN U7070 ( .B(n3091), .A(n3092), .Z(n3032) );
  XOR U7071 ( .A(n3018), .B(n3093), .Z(n3030) );
  XOR U7072 ( .A(n3019), .B(n3020), .Z(n3093) );
  XOR U7073 ( .A(n3025), .B(n3094), .Z(n3020) );
  XOR U7074 ( .A(n3024), .B(n3027), .Z(n3094) );
  IV U7075 ( .A(n3026), .Z(n3027) );
  NAND U7076 ( .A(n3095), .B(n3096), .Z(n3026) );
  OR U7077 ( .A(n3097), .B(n3098), .Z(n3096) );
  OR U7078 ( .A(n3099), .B(n3100), .Z(n3095) );
  NAND U7079 ( .A(n3101), .B(n3102), .Z(n3024) );
  OR U7080 ( .A(n3103), .B(n3104), .Z(n3102) );
  OR U7081 ( .A(n3105), .B(n3106), .Z(n3101) );
  NOR U7082 ( .A(n3107), .B(n3108), .Z(n3025) );
  ANDN U7083 ( .B(n3109), .A(n3110), .Z(n3019) );
  IV U7084 ( .A(n3111), .Z(n3109) );
  XNOR U7085 ( .A(n3012), .B(n3112), .Z(n3018) );
  XNOR U7086 ( .A(n3011), .B(n3013), .Z(n3112) );
  NAND U7087 ( .A(n3113), .B(n3114), .Z(n3013) );
  OR U7088 ( .A(n3115), .B(n3116), .Z(n3114) );
  OR U7089 ( .A(n3117), .B(n3118), .Z(n3113) );
  NAND U7090 ( .A(n3119), .B(n3120), .Z(n3011) );
  OR U7091 ( .A(n3121), .B(n3122), .Z(n3120) );
  OR U7092 ( .A(n3123), .B(n3124), .Z(n3119) );
  ANDN U7093 ( .B(n3125), .A(n3126), .Z(n3012) );
  IV U7094 ( .A(n3127), .Z(n3125) );
  XNOR U7095 ( .A(n3092), .B(n3091), .Z(N29897) );
  XOR U7096 ( .A(n3111), .B(n3110), .Z(n3091) );
  XNOR U7097 ( .A(n3126), .B(n3127), .Z(n3110) );
  XNOR U7098 ( .A(n3121), .B(n3122), .Z(n3127) );
  XNOR U7099 ( .A(n3123), .B(n3124), .Z(n3122) );
  XNOR U7100 ( .A(y[3940]), .B(x[3940]), .Z(n3124) );
  XNOR U7101 ( .A(y[3941]), .B(x[3941]), .Z(n3123) );
  XNOR U7102 ( .A(y[3939]), .B(x[3939]), .Z(n3121) );
  XNOR U7103 ( .A(n3115), .B(n3116), .Z(n3126) );
  XNOR U7104 ( .A(y[3936]), .B(x[3936]), .Z(n3116) );
  XNOR U7105 ( .A(n3117), .B(n3118), .Z(n3115) );
  XNOR U7106 ( .A(y[3937]), .B(x[3937]), .Z(n3118) );
  XNOR U7107 ( .A(y[3938]), .B(x[3938]), .Z(n3117) );
  XNOR U7108 ( .A(n3108), .B(n3107), .Z(n3111) );
  XNOR U7109 ( .A(n3103), .B(n3104), .Z(n3107) );
  XNOR U7110 ( .A(y[3933]), .B(x[3933]), .Z(n3104) );
  XNOR U7111 ( .A(n3105), .B(n3106), .Z(n3103) );
  XNOR U7112 ( .A(y[3934]), .B(x[3934]), .Z(n3106) );
  XNOR U7113 ( .A(y[3935]), .B(x[3935]), .Z(n3105) );
  XNOR U7114 ( .A(n3097), .B(n3098), .Z(n3108) );
  XNOR U7115 ( .A(y[3930]), .B(x[3930]), .Z(n3098) );
  XNOR U7116 ( .A(n3099), .B(n3100), .Z(n3097) );
  XNOR U7117 ( .A(y[3931]), .B(x[3931]), .Z(n3100) );
  XNOR U7118 ( .A(y[3932]), .B(x[3932]), .Z(n3099) );
  XOR U7119 ( .A(n3073), .B(n3074), .Z(n3092) );
  XNOR U7120 ( .A(n3089), .B(n3090), .Z(n3074) );
  XNOR U7121 ( .A(n3084), .B(n3085), .Z(n3090) );
  XNOR U7122 ( .A(n3086), .B(n3087), .Z(n3085) );
  XNOR U7123 ( .A(y[3928]), .B(x[3928]), .Z(n3087) );
  XNOR U7124 ( .A(y[3929]), .B(x[3929]), .Z(n3086) );
  XNOR U7125 ( .A(y[3927]), .B(x[3927]), .Z(n3084) );
  XNOR U7126 ( .A(n3078), .B(n3079), .Z(n3089) );
  XNOR U7127 ( .A(y[3924]), .B(x[3924]), .Z(n3079) );
  XNOR U7128 ( .A(n3080), .B(n3081), .Z(n3078) );
  XNOR U7129 ( .A(y[3925]), .B(x[3925]), .Z(n3081) );
  XNOR U7130 ( .A(y[3926]), .B(x[3926]), .Z(n3080) );
  XOR U7131 ( .A(n3072), .B(n3071), .Z(n3073) );
  XNOR U7132 ( .A(n3067), .B(n3068), .Z(n3071) );
  XNOR U7133 ( .A(y[3921]), .B(x[3921]), .Z(n3068) );
  XNOR U7134 ( .A(n3069), .B(n3070), .Z(n3067) );
  XNOR U7135 ( .A(y[3922]), .B(x[3922]), .Z(n3070) );
  XNOR U7136 ( .A(y[3923]), .B(x[3923]), .Z(n3069) );
  XNOR U7137 ( .A(n3061), .B(n3062), .Z(n3072) );
  XNOR U7138 ( .A(y[3918]), .B(x[3918]), .Z(n3062) );
  XNOR U7139 ( .A(n3063), .B(n3064), .Z(n3061) );
  XNOR U7140 ( .A(y[3919]), .B(x[3919]), .Z(n3064) );
  XNOR U7141 ( .A(y[3920]), .B(x[3920]), .Z(n3063) );
  NAND U7142 ( .A(n3128), .B(n3129), .Z(N29889) );
  NANDN U7143 ( .A(n3130), .B(n3131), .Z(n3129) );
  OR U7144 ( .A(n3132), .B(n3133), .Z(n3131) );
  NAND U7145 ( .A(n3132), .B(n3133), .Z(n3128) );
  XOR U7146 ( .A(n3132), .B(n3134), .Z(N29888) );
  XNOR U7147 ( .A(n3130), .B(n3133), .Z(n3134) );
  AND U7148 ( .A(n3135), .B(n3136), .Z(n3133) );
  NANDN U7149 ( .A(n3137), .B(n3138), .Z(n3136) );
  NANDN U7150 ( .A(n3139), .B(n3140), .Z(n3138) );
  NANDN U7151 ( .A(n3140), .B(n3139), .Z(n3135) );
  NAND U7152 ( .A(n3141), .B(n3142), .Z(n3130) );
  NANDN U7153 ( .A(n3143), .B(n3144), .Z(n3142) );
  OR U7154 ( .A(n3145), .B(n3146), .Z(n3144) );
  NAND U7155 ( .A(n3146), .B(n3145), .Z(n3141) );
  AND U7156 ( .A(n3147), .B(n3148), .Z(n3132) );
  NANDN U7157 ( .A(n3149), .B(n3150), .Z(n3148) );
  NANDN U7158 ( .A(n3151), .B(n3152), .Z(n3150) );
  NANDN U7159 ( .A(n3152), .B(n3151), .Z(n3147) );
  XOR U7160 ( .A(n3146), .B(n3153), .Z(N29887) );
  XOR U7161 ( .A(n3143), .B(n3145), .Z(n3153) );
  XNOR U7162 ( .A(n3139), .B(n3154), .Z(n3145) );
  XNOR U7163 ( .A(n3137), .B(n3140), .Z(n3154) );
  NAND U7164 ( .A(n3155), .B(n3156), .Z(n3140) );
  NAND U7165 ( .A(n3157), .B(n3158), .Z(n3156) );
  OR U7166 ( .A(n3159), .B(n3160), .Z(n3157) );
  NANDN U7167 ( .A(n3161), .B(n3159), .Z(n3155) );
  IV U7168 ( .A(n3160), .Z(n3161) );
  NAND U7169 ( .A(n3162), .B(n3163), .Z(n3137) );
  NAND U7170 ( .A(n3164), .B(n3165), .Z(n3163) );
  NANDN U7171 ( .A(n3166), .B(n3167), .Z(n3164) );
  NANDN U7172 ( .A(n3167), .B(n3166), .Z(n3162) );
  AND U7173 ( .A(n3168), .B(n3169), .Z(n3139) );
  NAND U7174 ( .A(n3170), .B(n3171), .Z(n3169) );
  OR U7175 ( .A(n3172), .B(n3173), .Z(n3170) );
  NANDN U7176 ( .A(n3174), .B(n3172), .Z(n3168) );
  NAND U7177 ( .A(n3175), .B(n3176), .Z(n3143) );
  NANDN U7178 ( .A(n3177), .B(n3178), .Z(n3176) );
  OR U7179 ( .A(n3179), .B(n3180), .Z(n3178) );
  NANDN U7180 ( .A(n3181), .B(n3179), .Z(n3175) );
  IV U7181 ( .A(n3180), .Z(n3181) );
  XNOR U7182 ( .A(n3151), .B(n3182), .Z(n3146) );
  XNOR U7183 ( .A(n3149), .B(n3152), .Z(n3182) );
  NAND U7184 ( .A(n3183), .B(n3184), .Z(n3152) );
  NAND U7185 ( .A(n3185), .B(n3186), .Z(n3184) );
  OR U7186 ( .A(n3187), .B(n3188), .Z(n3185) );
  NANDN U7187 ( .A(n3189), .B(n3187), .Z(n3183) );
  IV U7188 ( .A(n3188), .Z(n3189) );
  NAND U7189 ( .A(n3190), .B(n3191), .Z(n3149) );
  NAND U7190 ( .A(n3192), .B(n3193), .Z(n3191) );
  NANDN U7191 ( .A(n3194), .B(n3195), .Z(n3192) );
  NANDN U7192 ( .A(n3195), .B(n3194), .Z(n3190) );
  AND U7193 ( .A(n3196), .B(n3197), .Z(n3151) );
  NAND U7194 ( .A(n3198), .B(n3199), .Z(n3197) );
  OR U7195 ( .A(n3200), .B(n3201), .Z(n3198) );
  NANDN U7196 ( .A(n3202), .B(n3200), .Z(n3196) );
  XNOR U7197 ( .A(n3177), .B(n3203), .Z(N29886) );
  XOR U7198 ( .A(n3179), .B(n3180), .Z(n3203) );
  XNOR U7199 ( .A(n3193), .B(n3204), .Z(n3180) );
  XOR U7200 ( .A(n3194), .B(n3195), .Z(n3204) );
  XOR U7201 ( .A(n3200), .B(n3205), .Z(n3195) );
  XOR U7202 ( .A(n3199), .B(n3202), .Z(n3205) );
  IV U7203 ( .A(n3201), .Z(n3202) );
  NAND U7204 ( .A(n3206), .B(n3207), .Z(n3201) );
  OR U7205 ( .A(n3208), .B(n3209), .Z(n3207) );
  OR U7206 ( .A(n3210), .B(n3211), .Z(n3206) );
  NAND U7207 ( .A(n3212), .B(n3213), .Z(n3199) );
  OR U7208 ( .A(n3214), .B(n3215), .Z(n3213) );
  OR U7209 ( .A(n3216), .B(n3217), .Z(n3212) );
  NOR U7210 ( .A(n3218), .B(n3219), .Z(n3200) );
  ANDN U7211 ( .B(n3220), .A(n3221), .Z(n3194) );
  XNOR U7212 ( .A(n3187), .B(n3222), .Z(n3193) );
  XNOR U7213 ( .A(n3186), .B(n3188), .Z(n3222) );
  NAND U7214 ( .A(n3223), .B(n3224), .Z(n3188) );
  OR U7215 ( .A(n3225), .B(n3226), .Z(n3224) );
  OR U7216 ( .A(n3227), .B(n3228), .Z(n3223) );
  NAND U7217 ( .A(n3229), .B(n3230), .Z(n3186) );
  OR U7218 ( .A(n3231), .B(n3232), .Z(n3230) );
  OR U7219 ( .A(n3233), .B(n3234), .Z(n3229) );
  ANDN U7220 ( .B(n3235), .A(n3236), .Z(n3187) );
  IV U7221 ( .A(n3237), .Z(n3235) );
  ANDN U7222 ( .B(n3238), .A(n3239), .Z(n3179) );
  XOR U7223 ( .A(n3165), .B(n3240), .Z(n3177) );
  XOR U7224 ( .A(n3166), .B(n3167), .Z(n3240) );
  XOR U7225 ( .A(n3172), .B(n3241), .Z(n3167) );
  XOR U7226 ( .A(n3171), .B(n3174), .Z(n3241) );
  IV U7227 ( .A(n3173), .Z(n3174) );
  NAND U7228 ( .A(n3242), .B(n3243), .Z(n3173) );
  OR U7229 ( .A(n3244), .B(n3245), .Z(n3243) );
  OR U7230 ( .A(n3246), .B(n3247), .Z(n3242) );
  NAND U7231 ( .A(n3248), .B(n3249), .Z(n3171) );
  OR U7232 ( .A(n3250), .B(n3251), .Z(n3249) );
  OR U7233 ( .A(n3252), .B(n3253), .Z(n3248) );
  NOR U7234 ( .A(n3254), .B(n3255), .Z(n3172) );
  ANDN U7235 ( .B(n3256), .A(n3257), .Z(n3166) );
  IV U7236 ( .A(n3258), .Z(n3256) );
  XNOR U7237 ( .A(n3159), .B(n3259), .Z(n3165) );
  XNOR U7238 ( .A(n3158), .B(n3160), .Z(n3259) );
  NAND U7239 ( .A(n3260), .B(n3261), .Z(n3160) );
  OR U7240 ( .A(n3262), .B(n3263), .Z(n3261) );
  OR U7241 ( .A(n3264), .B(n3265), .Z(n3260) );
  NAND U7242 ( .A(n3266), .B(n3267), .Z(n3158) );
  OR U7243 ( .A(n3268), .B(n3269), .Z(n3267) );
  OR U7244 ( .A(n3270), .B(n3271), .Z(n3266) );
  ANDN U7245 ( .B(n3272), .A(n3273), .Z(n3159) );
  IV U7246 ( .A(n3274), .Z(n3272) );
  XNOR U7247 ( .A(n3239), .B(n3238), .Z(N29885) );
  XOR U7248 ( .A(n3258), .B(n3257), .Z(n3238) );
  XNOR U7249 ( .A(n3273), .B(n3274), .Z(n3257) );
  XNOR U7250 ( .A(n3268), .B(n3269), .Z(n3274) );
  XNOR U7251 ( .A(n3270), .B(n3271), .Z(n3269) );
  XNOR U7252 ( .A(y[3916]), .B(x[3916]), .Z(n3271) );
  XNOR U7253 ( .A(y[3917]), .B(x[3917]), .Z(n3270) );
  XNOR U7254 ( .A(y[3915]), .B(x[3915]), .Z(n3268) );
  XNOR U7255 ( .A(n3262), .B(n3263), .Z(n3273) );
  XNOR U7256 ( .A(y[3912]), .B(x[3912]), .Z(n3263) );
  XNOR U7257 ( .A(n3264), .B(n3265), .Z(n3262) );
  XNOR U7258 ( .A(y[3913]), .B(x[3913]), .Z(n3265) );
  XNOR U7259 ( .A(y[3914]), .B(x[3914]), .Z(n3264) );
  XNOR U7260 ( .A(n3255), .B(n3254), .Z(n3258) );
  XNOR U7261 ( .A(n3250), .B(n3251), .Z(n3254) );
  XNOR U7262 ( .A(y[3909]), .B(x[3909]), .Z(n3251) );
  XNOR U7263 ( .A(n3252), .B(n3253), .Z(n3250) );
  XNOR U7264 ( .A(y[3910]), .B(x[3910]), .Z(n3253) );
  XNOR U7265 ( .A(y[3911]), .B(x[3911]), .Z(n3252) );
  XNOR U7266 ( .A(n3244), .B(n3245), .Z(n3255) );
  XNOR U7267 ( .A(y[3906]), .B(x[3906]), .Z(n3245) );
  XNOR U7268 ( .A(n3246), .B(n3247), .Z(n3244) );
  XNOR U7269 ( .A(y[3907]), .B(x[3907]), .Z(n3247) );
  XNOR U7270 ( .A(y[3908]), .B(x[3908]), .Z(n3246) );
  XOR U7271 ( .A(n3220), .B(n3221), .Z(n3239) );
  XNOR U7272 ( .A(n3236), .B(n3237), .Z(n3221) );
  XNOR U7273 ( .A(n3231), .B(n3232), .Z(n3237) );
  XNOR U7274 ( .A(n3233), .B(n3234), .Z(n3232) );
  XNOR U7275 ( .A(y[3904]), .B(x[3904]), .Z(n3234) );
  XNOR U7276 ( .A(y[3905]), .B(x[3905]), .Z(n3233) );
  XNOR U7277 ( .A(y[3903]), .B(x[3903]), .Z(n3231) );
  XNOR U7278 ( .A(n3225), .B(n3226), .Z(n3236) );
  XNOR U7279 ( .A(y[3900]), .B(x[3900]), .Z(n3226) );
  XNOR U7280 ( .A(n3227), .B(n3228), .Z(n3225) );
  XNOR U7281 ( .A(y[3901]), .B(x[3901]), .Z(n3228) );
  XNOR U7282 ( .A(y[3902]), .B(x[3902]), .Z(n3227) );
  XOR U7283 ( .A(n3219), .B(n3218), .Z(n3220) );
  XNOR U7284 ( .A(n3214), .B(n3215), .Z(n3218) );
  XNOR U7285 ( .A(y[3897]), .B(x[3897]), .Z(n3215) );
  XNOR U7286 ( .A(n3216), .B(n3217), .Z(n3214) );
  XNOR U7287 ( .A(y[3898]), .B(x[3898]), .Z(n3217) );
  XNOR U7288 ( .A(y[3899]), .B(x[3899]), .Z(n3216) );
  XNOR U7289 ( .A(n3208), .B(n3209), .Z(n3219) );
  XNOR U7290 ( .A(y[3894]), .B(x[3894]), .Z(n3209) );
  XNOR U7291 ( .A(n3210), .B(n3211), .Z(n3208) );
  XNOR U7292 ( .A(y[3895]), .B(x[3895]), .Z(n3211) );
  XNOR U7293 ( .A(y[3896]), .B(x[3896]), .Z(n3210) );
  NAND U7294 ( .A(n3275), .B(n3276), .Z(N29877) );
  NANDN U7295 ( .A(n3277), .B(n3278), .Z(n3276) );
  OR U7296 ( .A(n3279), .B(n3280), .Z(n3278) );
  NAND U7297 ( .A(n3279), .B(n3280), .Z(n3275) );
  XOR U7298 ( .A(n3279), .B(n3281), .Z(N29876) );
  XNOR U7299 ( .A(n3277), .B(n3280), .Z(n3281) );
  AND U7300 ( .A(n3282), .B(n3283), .Z(n3280) );
  NANDN U7301 ( .A(n3284), .B(n3285), .Z(n3283) );
  NANDN U7302 ( .A(n3286), .B(n3287), .Z(n3285) );
  NANDN U7303 ( .A(n3287), .B(n3286), .Z(n3282) );
  NAND U7304 ( .A(n3288), .B(n3289), .Z(n3277) );
  NANDN U7305 ( .A(n3290), .B(n3291), .Z(n3289) );
  OR U7306 ( .A(n3292), .B(n3293), .Z(n3291) );
  NAND U7307 ( .A(n3293), .B(n3292), .Z(n3288) );
  AND U7308 ( .A(n3294), .B(n3295), .Z(n3279) );
  NANDN U7309 ( .A(n3296), .B(n3297), .Z(n3295) );
  NANDN U7310 ( .A(n3298), .B(n3299), .Z(n3297) );
  NANDN U7311 ( .A(n3299), .B(n3298), .Z(n3294) );
  XOR U7312 ( .A(n3293), .B(n3300), .Z(N29875) );
  XOR U7313 ( .A(n3290), .B(n3292), .Z(n3300) );
  XNOR U7314 ( .A(n3286), .B(n3301), .Z(n3292) );
  XNOR U7315 ( .A(n3284), .B(n3287), .Z(n3301) );
  NAND U7316 ( .A(n3302), .B(n3303), .Z(n3287) );
  NAND U7317 ( .A(n3304), .B(n3305), .Z(n3303) );
  OR U7318 ( .A(n3306), .B(n3307), .Z(n3304) );
  NANDN U7319 ( .A(n3308), .B(n3306), .Z(n3302) );
  IV U7320 ( .A(n3307), .Z(n3308) );
  NAND U7321 ( .A(n3309), .B(n3310), .Z(n3284) );
  NAND U7322 ( .A(n3311), .B(n3312), .Z(n3310) );
  NANDN U7323 ( .A(n3313), .B(n3314), .Z(n3311) );
  NANDN U7324 ( .A(n3314), .B(n3313), .Z(n3309) );
  AND U7325 ( .A(n3315), .B(n3316), .Z(n3286) );
  NAND U7326 ( .A(n3317), .B(n3318), .Z(n3316) );
  OR U7327 ( .A(n3319), .B(n3320), .Z(n3317) );
  NANDN U7328 ( .A(n3321), .B(n3319), .Z(n3315) );
  NAND U7329 ( .A(n3322), .B(n3323), .Z(n3290) );
  NANDN U7330 ( .A(n3324), .B(n3325), .Z(n3323) );
  OR U7331 ( .A(n3326), .B(n3327), .Z(n3325) );
  NANDN U7332 ( .A(n3328), .B(n3326), .Z(n3322) );
  IV U7333 ( .A(n3327), .Z(n3328) );
  XNOR U7334 ( .A(n3298), .B(n3329), .Z(n3293) );
  XNOR U7335 ( .A(n3296), .B(n3299), .Z(n3329) );
  NAND U7336 ( .A(n3330), .B(n3331), .Z(n3299) );
  NAND U7337 ( .A(n3332), .B(n3333), .Z(n3331) );
  OR U7338 ( .A(n3334), .B(n3335), .Z(n3332) );
  NANDN U7339 ( .A(n3336), .B(n3334), .Z(n3330) );
  IV U7340 ( .A(n3335), .Z(n3336) );
  NAND U7341 ( .A(n3337), .B(n3338), .Z(n3296) );
  NAND U7342 ( .A(n3339), .B(n3340), .Z(n3338) );
  NANDN U7343 ( .A(n3341), .B(n3342), .Z(n3339) );
  NANDN U7344 ( .A(n3342), .B(n3341), .Z(n3337) );
  AND U7345 ( .A(n3343), .B(n3344), .Z(n3298) );
  NAND U7346 ( .A(n3345), .B(n3346), .Z(n3344) );
  OR U7347 ( .A(n3347), .B(n3348), .Z(n3345) );
  NANDN U7348 ( .A(n3349), .B(n3347), .Z(n3343) );
  XNOR U7349 ( .A(n3324), .B(n3350), .Z(N29874) );
  XOR U7350 ( .A(n3326), .B(n3327), .Z(n3350) );
  XNOR U7351 ( .A(n3340), .B(n3351), .Z(n3327) );
  XOR U7352 ( .A(n3341), .B(n3342), .Z(n3351) );
  XOR U7353 ( .A(n3347), .B(n3352), .Z(n3342) );
  XOR U7354 ( .A(n3346), .B(n3349), .Z(n3352) );
  IV U7355 ( .A(n3348), .Z(n3349) );
  NAND U7356 ( .A(n3353), .B(n3354), .Z(n3348) );
  OR U7357 ( .A(n3355), .B(n3356), .Z(n3354) );
  OR U7358 ( .A(n3357), .B(n3358), .Z(n3353) );
  NAND U7359 ( .A(n3359), .B(n3360), .Z(n3346) );
  OR U7360 ( .A(n3361), .B(n3362), .Z(n3360) );
  OR U7361 ( .A(n3363), .B(n3364), .Z(n3359) );
  NOR U7362 ( .A(n3365), .B(n3366), .Z(n3347) );
  ANDN U7363 ( .B(n3367), .A(n3368), .Z(n3341) );
  XNOR U7364 ( .A(n3334), .B(n3369), .Z(n3340) );
  XNOR U7365 ( .A(n3333), .B(n3335), .Z(n3369) );
  NAND U7366 ( .A(n3370), .B(n3371), .Z(n3335) );
  OR U7367 ( .A(n3372), .B(n3373), .Z(n3371) );
  OR U7368 ( .A(n3374), .B(n3375), .Z(n3370) );
  NAND U7369 ( .A(n3376), .B(n3377), .Z(n3333) );
  OR U7370 ( .A(n3378), .B(n3379), .Z(n3377) );
  OR U7371 ( .A(n3380), .B(n3381), .Z(n3376) );
  ANDN U7372 ( .B(n3382), .A(n3383), .Z(n3334) );
  IV U7373 ( .A(n3384), .Z(n3382) );
  ANDN U7374 ( .B(n3385), .A(n3386), .Z(n3326) );
  XOR U7375 ( .A(n3312), .B(n3387), .Z(n3324) );
  XOR U7376 ( .A(n3313), .B(n3314), .Z(n3387) );
  XOR U7377 ( .A(n3319), .B(n3388), .Z(n3314) );
  XOR U7378 ( .A(n3318), .B(n3321), .Z(n3388) );
  IV U7379 ( .A(n3320), .Z(n3321) );
  NAND U7380 ( .A(n3389), .B(n3390), .Z(n3320) );
  OR U7381 ( .A(n3391), .B(n3392), .Z(n3390) );
  OR U7382 ( .A(n3393), .B(n3394), .Z(n3389) );
  NAND U7383 ( .A(n3395), .B(n3396), .Z(n3318) );
  OR U7384 ( .A(n3397), .B(n3398), .Z(n3396) );
  OR U7385 ( .A(n3399), .B(n3400), .Z(n3395) );
  NOR U7386 ( .A(n3401), .B(n3402), .Z(n3319) );
  ANDN U7387 ( .B(n3403), .A(n3404), .Z(n3313) );
  IV U7388 ( .A(n3405), .Z(n3403) );
  XNOR U7389 ( .A(n3306), .B(n3406), .Z(n3312) );
  XNOR U7390 ( .A(n3305), .B(n3307), .Z(n3406) );
  NAND U7391 ( .A(n3407), .B(n3408), .Z(n3307) );
  OR U7392 ( .A(n3409), .B(n3410), .Z(n3408) );
  OR U7393 ( .A(n3411), .B(n3412), .Z(n3407) );
  NAND U7394 ( .A(n3413), .B(n3414), .Z(n3305) );
  OR U7395 ( .A(n3415), .B(n3416), .Z(n3414) );
  OR U7396 ( .A(n3417), .B(n3418), .Z(n3413) );
  ANDN U7397 ( .B(n3419), .A(n3420), .Z(n3306) );
  IV U7398 ( .A(n3421), .Z(n3419) );
  XNOR U7399 ( .A(n3386), .B(n3385), .Z(N29873) );
  XOR U7400 ( .A(n3405), .B(n3404), .Z(n3385) );
  XNOR U7401 ( .A(n3420), .B(n3421), .Z(n3404) );
  XNOR U7402 ( .A(n3415), .B(n3416), .Z(n3421) );
  XNOR U7403 ( .A(n3417), .B(n3418), .Z(n3416) );
  XNOR U7404 ( .A(y[3892]), .B(x[3892]), .Z(n3418) );
  XNOR U7405 ( .A(y[3893]), .B(x[3893]), .Z(n3417) );
  XNOR U7406 ( .A(y[3891]), .B(x[3891]), .Z(n3415) );
  XNOR U7407 ( .A(n3409), .B(n3410), .Z(n3420) );
  XNOR U7408 ( .A(y[3888]), .B(x[3888]), .Z(n3410) );
  XNOR U7409 ( .A(n3411), .B(n3412), .Z(n3409) );
  XNOR U7410 ( .A(y[3889]), .B(x[3889]), .Z(n3412) );
  XNOR U7411 ( .A(y[3890]), .B(x[3890]), .Z(n3411) );
  XNOR U7412 ( .A(n3402), .B(n3401), .Z(n3405) );
  XNOR U7413 ( .A(n3397), .B(n3398), .Z(n3401) );
  XNOR U7414 ( .A(y[3885]), .B(x[3885]), .Z(n3398) );
  XNOR U7415 ( .A(n3399), .B(n3400), .Z(n3397) );
  XNOR U7416 ( .A(y[3886]), .B(x[3886]), .Z(n3400) );
  XNOR U7417 ( .A(y[3887]), .B(x[3887]), .Z(n3399) );
  XNOR U7418 ( .A(n3391), .B(n3392), .Z(n3402) );
  XNOR U7419 ( .A(y[3882]), .B(x[3882]), .Z(n3392) );
  XNOR U7420 ( .A(n3393), .B(n3394), .Z(n3391) );
  XNOR U7421 ( .A(y[3883]), .B(x[3883]), .Z(n3394) );
  XNOR U7422 ( .A(y[3884]), .B(x[3884]), .Z(n3393) );
  XOR U7423 ( .A(n3367), .B(n3368), .Z(n3386) );
  XNOR U7424 ( .A(n3383), .B(n3384), .Z(n3368) );
  XNOR U7425 ( .A(n3378), .B(n3379), .Z(n3384) );
  XNOR U7426 ( .A(n3380), .B(n3381), .Z(n3379) );
  XNOR U7427 ( .A(y[3880]), .B(x[3880]), .Z(n3381) );
  XNOR U7428 ( .A(y[3881]), .B(x[3881]), .Z(n3380) );
  XNOR U7429 ( .A(y[3879]), .B(x[3879]), .Z(n3378) );
  XNOR U7430 ( .A(n3372), .B(n3373), .Z(n3383) );
  XNOR U7431 ( .A(y[3876]), .B(x[3876]), .Z(n3373) );
  XNOR U7432 ( .A(n3374), .B(n3375), .Z(n3372) );
  XNOR U7433 ( .A(y[3877]), .B(x[3877]), .Z(n3375) );
  XNOR U7434 ( .A(y[3878]), .B(x[3878]), .Z(n3374) );
  XOR U7435 ( .A(n3366), .B(n3365), .Z(n3367) );
  XNOR U7436 ( .A(n3361), .B(n3362), .Z(n3365) );
  XNOR U7437 ( .A(y[3873]), .B(x[3873]), .Z(n3362) );
  XNOR U7438 ( .A(n3363), .B(n3364), .Z(n3361) );
  XNOR U7439 ( .A(y[3874]), .B(x[3874]), .Z(n3364) );
  XNOR U7440 ( .A(y[3875]), .B(x[3875]), .Z(n3363) );
  XNOR U7441 ( .A(n3355), .B(n3356), .Z(n3366) );
  XNOR U7442 ( .A(y[3870]), .B(x[3870]), .Z(n3356) );
  XNOR U7443 ( .A(n3357), .B(n3358), .Z(n3355) );
  XNOR U7444 ( .A(y[3871]), .B(x[3871]), .Z(n3358) );
  XNOR U7445 ( .A(y[3872]), .B(x[3872]), .Z(n3357) );
  NAND U7446 ( .A(n3422), .B(n3423), .Z(N29865) );
  NANDN U7447 ( .A(n3424), .B(n3425), .Z(n3423) );
  OR U7448 ( .A(n3426), .B(n3427), .Z(n3425) );
  NAND U7449 ( .A(n3426), .B(n3427), .Z(n3422) );
  XOR U7450 ( .A(n3426), .B(n3428), .Z(N29864) );
  XNOR U7451 ( .A(n3424), .B(n3427), .Z(n3428) );
  AND U7452 ( .A(n3429), .B(n3430), .Z(n3427) );
  NANDN U7453 ( .A(n3431), .B(n3432), .Z(n3430) );
  NANDN U7454 ( .A(n3433), .B(n3434), .Z(n3432) );
  NANDN U7455 ( .A(n3434), .B(n3433), .Z(n3429) );
  NAND U7456 ( .A(n3435), .B(n3436), .Z(n3424) );
  NANDN U7457 ( .A(n3437), .B(n3438), .Z(n3436) );
  OR U7458 ( .A(n3439), .B(n3440), .Z(n3438) );
  NAND U7459 ( .A(n3440), .B(n3439), .Z(n3435) );
  AND U7460 ( .A(n3441), .B(n3442), .Z(n3426) );
  NANDN U7461 ( .A(n3443), .B(n3444), .Z(n3442) );
  NANDN U7462 ( .A(n3445), .B(n3446), .Z(n3444) );
  NANDN U7463 ( .A(n3446), .B(n3445), .Z(n3441) );
  XOR U7464 ( .A(n3440), .B(n3447), .Z(N29863) );
  XOR U7465 ( .A(n3437), .B(n3439), .Z(n3447) );
  XNOR U7466 ( .A(n3433), .B(n3448), .Z(n3439) );
  XNOR U7467 ( .A(n3431), .B(n3434), .Z(n3448) );
  NAND U7468 ( .A(n3449), .B(n3450), .Z(n3434) );
  NAND U7469 ( .A(n3451), .B(n3452), .Z(n3450) );
  OR U7470 ( .A(n3453), .B(n3454), .Z(n3451) );
  NANDN U7471 ( .A(n3455), .B(n3453), .Z(n3449) );
  IV U7472 ( .A(n3454), .Z(n3455) );
  NAND U7473 ( .A(n3456), .B(n3457), .Z(n3431) );
  NAND U7474 ( .A(n3458), .B(n3459), .Z(n3457) );
  NANDN U7475 ( .A(n3460), .B(n3461), .Z(n3458) );
  NANDN U7476 ( .A(n3461), .B(n3460), .Z(n3456) );
  AND U7477 ( .A(n3462), .B(n3463), .Z(n3433) );
  NAND U7478 ( .A(n3464), .B(n3465), .Z(n3463) );
  OR U7479 ( .A(n3466), .B(n3467), .Z(n3464) );
  NANDN U7480 ( .A(n3468), .B(n3466), .Z(n3462) );
  NAND U7481 ( .A(n3469), .B(n3470), .Z(n3437) );
  NANDN U7482 ( .A(n3471), .B(n3472), .Z(n3470) );
  OR U7483 ( .A(n3473), .B(n3474), .Z(n3472) );
  NANDN U7484 ( .A(n3475), .B(n3473), .Z(n3469) );
  IV U7485 ( .A(n3474), .Z(n3475) );
  XNOR U7486 ( .A(n3445), .B(n3476), .Z(n3440) );
  XNOR U7487 ( .A(n3443), .B(n3446), .Z(n3476) );
  NAND U7488 ( .A(n3477), .B(n3478), .Z(n3446) );
  NAND U7489 ( .A(n3479), .B(n3480), .Z(n3478) );
  OR U7490 ( .A(n3481), .B(n3482), .Z(n3479) );
  NANDN U7491 ( .A(n3483), .B(n3481), .Z(n3477) );
  IV U7492 ( .A(n3482), .Z(n3483) );
  NAND U7493 ( .A(n3484), .B(n3485), .Z(n3443) );
  NAND U7494 ( .A(n3486), .B(n3487), .Z(n3485) );
  NANDN U7495 ( .A(n3488), .B(n3489), .Z(n3486) );
  NANDN U7496 ( .A(n3489), .B(n3488), .Z(n3484) );
  AND U7497 ( .A(n3490), .B(n3491), .Z(n3445) );
  NAND U7498 ( .A(n3492), .B(n3493), .Z(n3491) );
  OR U7499 ( .A(n3494), .B(n3495), .Z(n3492) );
  NANDN U7500 ( .A(n3496), .B(n3494), .Z(n3490) );
  XNOR U7501 ( .A(n3471), .B(n3497), .Z(N29862) );
  XOR U7502 ( .A(n3473), .B(n3474), .Z(n3497) );
  XNOR U7503 ( .A(n3487), .B(n3498), .Z(n3474) );
  XOR U7504 ( .A(n3488), .B(n3489), .Z(n3498) );
  XOR U7505 ( .A(n3494), .B(n3499), .Z(n3489) );
  XOR U7506 ( .A(n3493), .B(n3496), .Z(n3499) );
  IV U7507 ( .A(n3495), .Z(n3496) );
  NAND U7508 ( .A(n3500), .B(n3501), .Z(n3495) );
  OR U7509 ( .A(n3502), .B(n3503), .Z(n3501) );
  OR U7510 ( .A(n3504), .B(n3505), .Z(n3500) );
  NAND U7511 ( .A(n3506), .B(n3507), .Z(n3493) );
  OR U7512 ( .A(n3508), .B(n3509), .Z(n3507) );
  OR U7513 ( .A(n3510), .B(n3511), .Z(n3506) );
  NOR U7514 ( .A(n3512), .B(n3513), .Z(n3494) );
  ANDN U7515 ( .B(n3514), .A(n3515), .Z(n3488) );
  XNOR U7516 ( .A(n3481), .B(n3516), .Z(n3487) );
  XNOR U7517 ( .A(n3480), .B(n3482), .Z(n3516) );
  NAND U7518 ( .A(n3517), .B(n3518), .Z(n3482) );
  OR U7519 ( .A(n3519), .B(n3520), .Z(n3518) );
  OR U7520 ( .A(n3521), .B(n3522), .Z(n3517) );
  NAND U7521 ( .A(n3523), .B(n3524), .Z(n3480) );
  OR U7522 ( .A(n3525), .B(n3526), .Z(n3524) );
  OR U7523 ( .A(n3527), .B(n3528), .Z(n3523) );
  ANDN U7524 ( .B(n3529), .A(n3530), .Z(n3481) );
  IV U7525 ( .A(n3531), .Z(n3529) );
  ANDN U7526 ( .B(n3532), .A(n3533), .Z(n3473) );
  XOR U7527 ( .A(n3459), .B(n3534), .Z(n3471) );
  XOR U7528 ( .A(n3460), .B(n3461), .Z(n3534) );
  XOR U7529 ( .A(n3466), .B(n3535), .Z(n3461) );
  XOR U7530 ( .A(n3465), .B(n3468), .Z(n3535) );
  IV U7531 ( .A(n3467), .Z(n3468) );
  NAND U7532 ( .A(n3536), .B(n3537), .Z(n3467) );
  OR U7533 ( .A(n3538), .B(n3539), .Z(n3537) );
  OR U7534 ( .A(n3540), .B(n3541), .Z(n3536) );
  NAND U7535 ( .A(n3542), .B(n3543), .Z(n3465) );
  OR U7536 ( .A(n3544), .B(n3545), .Z(n3543) );
  OR U7537 ( .A(n3546), .B(n3547), .Z(n3542) );
  NOR U7538 ( .A(n3548), .B(n3549), .Z(n3466) );
  ANDN U7539 ( .B(n3550), .A(n3551), .Z(n3460) );
  IV U7540 ( .A(n3552), .Z(n3550) );
  XNOR U7541 ( .A(n3453), .B(n3553), .Z(n3459) );
  XNOR U7542 ( .A(n3452), .B(n3454), .Z(n3553) );
  NAND U7543 ( .A(n3554), .B(n3555), .Z(n3454) );
  OR U7544 ( .A(n3556), .B(n3557), .Z(n3555) );
  OR U7545 ( .A(n3558), .B(n3559), .Z(n3554) );
  NAND U7546 ( .A(n3560), .B(n3561), .Z(n3452) );
  OR U7547 ( .A(n3562), .B(n3563), .Z(n3561) );
  OR U7548 ( .A(n3564), .B(n3565), .Z(n3560) );
  ANDN U7549 ( .B(n3566), .A(n3567), .Z(n3453) );
  IV U7550 ( .A(n3568), .Z(n3566) );
  XNOR U7551 ( .A(n3533), .B(n3532), .Z(N29861) );
  XOR U7552 ( .A(n3552), .B(n3551), .Z(n3532) );
  XNOR U7553 ( .A(n3567), .B(n3568), .Z(n3551) );
  XNOR U7554 ( .A(n3562), .B(n3563), .Z(n3568) );
  XNOR U7555 ( .A(n3564), .B(n3565), .Z(n3563) );
  XNOR U7556 ( .A(y[3868]), .B(x[3868]), .Z(n3565) );
  XNOR U7557 ( .A(y[3869]), .B(x[3869]), .Z(n3564) );
  XNOR U7558 ( .A(y[3867]), .B(x[3867]), .Z(n3562) );
  XNOR U7559 ( .A(n3556), .B(n3557), .Z(n3567) );
  XNOR U7560 ( .A(y[3864]), .B(x[3864]), .Z(n3557) );
  XNOR U7561 ( .A(n3558), .B(n3559), .Z(n3556) );
  XNOR U7562 ( .A(y[3865]), .B(x[3865]), .Z(n3559) );
  XNOR U7563 ( .A(y[3866]), .B(x[3866]), .Z(n3558) );
  XNOR U7564 ( .A(n3549), .B(n3548), .Z(n3552) );
  XNOR U7565 ( .A(n3544), .B(n3545), .Z(n3548) );
  XNOR U7566 ( .A(y[3861]), .B(x[3861]), .Z(n3545) );
  XNOR U7567 ( .A(n3546), .B(n3547), .Z(n3544) );
  XNOR U7568 ( .A(y[3862]), .B(x[3862]), .Z(n3547) );
  XNOR U7569 ( .A(y[3863]), .B(x[3863]), .Z(n3546) );
  XNOR U7570 ( .A(n3538), .B(n3539), .Z(n3549) );
  XNOR U7571 ( .A(y[3858]), .B(x[3858]), .Z(n3539) );
  XNOR U7572 ( .A(n3540), .B(n3541), .Z(n3538) );
  XNOR U7573 ( .A(y[3859]), .B(x[3859]), .Z(n3541) );
  XNOR U7574 ( .A(y[3860]), .B(x[3860]), .Z(n3540) );
  XOR U7575 ( .A(n3514), .B(n3515), .Z(n3533) );
  XNOR U7576 ( .A(n3530), .B(n3531), .Z(n3515) );
  XNOR U7577 ( .A(n3525), .B(n3526), .Z(n3531) );
  XNOR U7578 ( .A(n3527), .B(n3528), .Z(n3526) );
  XNOR U7579 ( .A(y[3856]), .B(x[3856]), .Z(n3528) );
  XNOR U7580 ( .A(y[3857]), .B(x[3857]), .Z(n3527) );
  XNOR U7581 ( .A(y[3855]), .B(x[3855]), .Z(n3525) );
  XNOR U7582 ( .A(n3519), .B(n3520), .Z(n3530) );
  XNOR U7583 ( .A(y[3852]), .B(x[3852]), .Z(n3520) );
  XNOR U7584 ( .A(n3521), .B(n3522), .Z(n3519) );
  XNOR U7585 ( .A(y[3853]), .B(x[3853]), .Z(n3522) );
  XNOR U7586 ( .A(y[3854]), .B(x[3854]), .Z(n3521) );
  XOR U7587 ( .A(n3513), .B(n3512), .Z(n3514) );
  XNOR U7588 ( .A(n3508), .B(n3509), .Z(n3512) );
  XNOR U7589 ( .A(y[3849]), .B(x[3849]), .Z(n3509) );
  XNOR U7590 ( .A(n3510), .B(n3511), .Z(n3508) );
  XNOR U7591 ( .A(y[3850]), .B(x[3850]), .Z(n3511) );
  XNOR U7592 ( .A(y[3851]), .B(x[3851]), .Z(n3510) );
  XNOR U7593 ( .A(n3502), .B(n3503), .Z(n3513) );
  XNOR U7594 ( .A(y[3846]), .B(x[3846]), .Z(n3503) );
  XNOR U7595 ( .A(n3504), .B(n3505), .Z(n3502) );
  XNOR U7596 ( .A(y[3847]), .B(x[3847]), .Z(n3505) );
  XNOR U7597 ( .A(y[3848]), .B(x[3848]), .Z(n3504) );
  NAND U7598 ( .A(n3569), .B(n3570), .Z(N29853) );
  NANDN U7599 ( .A(n3571), .B(n3572), .Z(n3570) );
  OR U7600 ( .A(n3573), .B(n3574), .Z(n3572) );
  NAND U7601 ( .A(n3573), .B(n3574), .Z(n3569) );
  XOR U7602 ( .A(n3573), .B(n3575), .Z(N29852) );
  XNOR U7603 ( .A(n3571), .B(n3574), .Z(n3575) );
  AND U7604 ( .A(n3576), .B(n3577), .Z(n3574) );
  NANDN U7605 ( .A(n3578), .B(n3579), .Z(n3577) );
  NANDN U7606 ( .A(n3580), .B(n3581), .Z(n3579) );
  NANDN U7607 ( .A(n3581), .B(n3580), .Z(n3576) );
  NAND U7608 ( .A(n3582), .B(n3583), .Z(n3571) );
  NANDN U7609 ( .A(n3584), .B(n3585), .Z(n3583) );
  OR U7610 ( .A(n3586), .B(n3587), .Z(n3585) );
  NAND U7611 ( .A(n3587), .B(n3586), .Z(n3582) );
  AND U7612 ( .A(n3588), .B(n3589), .Z(n3573) );
  NANDN U7613 ( .A(n3590), .B(n3591), .Z(n3589) );
  NANDN U7614 ( .A(n3592), .B(n3593), .Z(n3591) );
  NANDN U7615 ( .A(n3593), .B(n3592), .Z(n3588) );
  XOR U7616 ( .A(n3587), .B(n3594), .Z(N29851) );
  XOR U7617 ( .A(n3584), .B(n3586), .Z(n3594) );
  XNOR U7618 ( .A(n3580), .B(n3595), .Z(n3586) );
  XNOR U7619 ( .A(n3578), .B(n3581), .Z(n3595) );
  NAND U7620 ( .A(n3596), .B(n3597), .Z(n3581) );
  NAND U7621 ( .A(n3598), .B(n3599), .Z(n3597) );
  OR U7622 ( .A(n3600), .B(n3601), .Z(n3598) );
  NANDN U7623 ( .A(n3602), .B(n3600), .Z(n3596) );
  IV U7624 ( .A(n3601), .Z(n3602) );
  NAND U7625 ( .A(n3603), .B(n3604), .Z(n3578) );
  NAND U7626 ( .A(n3605), .B(n3606), .Z(n3604) );
  NANDN U7627 ( .A(n3607), .B(n3608), .Z(n3605) );
  NANDN U7628 ( .A(n3608), .B(n3607), .Z(n3603) );
  AND U7629 ( .A(n3609), .B(n3610), .Z(n3580) );
  NAND U7630 ( .A(n3611), .B(n3612), .Z(n3610) );
  OR U7631 ( .A(n3613), .B(n3614), .Z(n3611) );
  NANDN U7632 ( .A(n3615), .B(n3613), .Z(n3609) );
  NAND U7633 ( .A(n3616), .B(n3617), .Z(n3584) );
  NANDN U7634 ( .A(n3618), .B(n3619), .Z(n3617) );
  OR U7635 ( .A(n3620), .B(n3621), .Z(n3619) );
  NANDN U7636 ( .A(n3622), .B(n3620), .Z(n3616) );
  IV U7637 ( .A(n3621), .Z(n3622) );
  XNOR U7638 ( .A(n3592), .B(n3623), .Z(n3587) );
  XNOR U7639 ( .A(n3590), .B(n3593), .Z(n3623) );
  NAND U7640 ( .A(n3624), .B(n3625), .Z(n3593) );
  NAND U7641 ( .A(n3626), .B(n3627), .Z(n3625) );
  OR U7642 ( .A(n3628), .B(n3629), .Z(n3626) );
  NANDN U7643 ( .A(n3630), .B(n3628), .Z(n3624) );
  IV U7644 ( .A(n3629), .Z(n3630) );
  NAND U7645 ( .A(n3631), .B(n3632), .Z(n3590) );
  NAND U7646 ( .A(n3633), .B(n3634), .Z(n3632) );
  NANDN U7647 ( .A(n3635), .B(n3636), .Z(n3633) );
  NANDN U7648 ( .A(n3636), .B(n3635), .Z(n3631) );
  AND U7649 ( .A(n3637), .B(n3638), .Z(n3592) );
  NAND U7650 ( .A(n3639), .B(n3640), .Z(n3638) );
  OR U7651 ( .A(n3641), .B(n3642), .Z(n3639) );
  NANDN U7652 ( .A(n3643), .B(n3641), .Z(n3637) );
  XNOR U7653 ( .A(n3618), .B(n3644), .Z(N29850) );
  XOR U7654 ( .A(n3620), .B(n3621), .Z(n3644) );
  XNOR U7655 ( .A(n3634), .B(n3645), .Z(n3621) );
  XOR U7656 ( .A(n3635), .B(n3636), .Z(n3645) );
  XOR U7657 ( .A(n3641), .B(n3646), .Z(n3636) );
  XOR U7658 ( .A(n3640), .B(n3643), .Z(n3646) );
  IV U7659 ( .A(n3642), .Z(n3643) );
  NAND U7660 ( .A(n3647), .B(n3648), .Z(n3642) );
  OR U7661 ( .A(n3649), .B(n3650), .Z(n3648) );
  OR U7662 ( .A(n3651), .B(n3652), .Z(n3647) );
  NAND U7663 ( .A(n3653), .B(n3654), .Z(n3640) );
  OR U7664 ( .A(n3655), .B(n3656), .Z(n3654) );
  OR U7665 ( .A(n3657), .B(n3658), .Z(n3653) );
  NOR U7666 ( .A(n3659), .B(n3660), .Z(n3641) );
  ANDN U7667 ( .B(n3661), .A(n3662), .Z(n3635) );
  XNOR U7668 ( .A(n3628), .B(n3663), .Z(n3634) );
  XNOR U7669 ( .A(n3627), .B(n3629), .Z(n3663) );
  NAND U7670 ( .A(n3664), .B(n3665), .Z(n3629) );
  OR U7671 ( .A(n3666), .B(n3667), .Z(n3665) );
  OR U7672 ( .A(n3668), .B(n3669), .Z(n3664) );
  NAND U7673 ( .A(n3670), .B(n3671), .Z(n3627) );
  OR U7674 ( .A(n3672), .B(n3673), .Z(n3671) );
  OR U7675 ( .A(n3674), .B(n3675), .Z(n3670) );
  ANDN U7676 ( .B(n3676), .A(n3677), .Z(n3628) );
  IV U7677 ( .A(n3678), .Z(n3676) );
  ANDN U7678 ( .B(n3679), .A(n3680), .Z(n3620) );
  XOR U7679 ( .A(n3606), .B(n3681), .Z(n3618) );
  XOR U7680 ( .A(n3607), .B(n3608), .Z(n3681) );
  XOR U7681 ( .A(n3613), .B(n3682), .Z(n3608) );
  XOR U7682 ( .A(n3612), .B(n3615), .Z(n3682) );
  IV U7683 ( .A(n3614), .Z(n3615) );
  NAND U7684 ( .A(n3683), .B(n3684), .Z(n3614) );
  OR U7685 ( .A(n3685), .B(n3686), .Z(n3684) );
  OR U7686 ( .A(n3687), .B(n3688), .Z(n3683) );
  NAND U7687 ( .A(n3689), .B(n3690), .Z(n3612) );
  OR U7688 ( .A(n3691), .B(n3692), .Z(n3690) );
  OR U7689 ( .A(n3693), .B(n3694), .Z(n3689) );
  NOR U7690 ( .A(n3695), .B(n3696), .Z(n3613) );
  ANDN U7691 ( .B(n3697), .A(n3698), .Z(n3607) );
  IV U7692 ( .A(n3699), .Z(n3697) );
  XNOR U7693 ( .A(n3600), .B(n3700), .Z(n3606) );
  XNOR U7694 ( .A(n3599), .B(n3601), .Z(n3700) );
  NAND U7695 ( .A(n3701), .B(n3702), .Z(n3601) );
  OR U7696 ( .A(n3703), .B(n3704), .Z(n3702) );
  OR U7697 ( .A(n3705), .B(n3706), .Z(n3701) );
  NAND U7698 ( .A(n3707), .B(n3708), .Z(n3599) );
  OR U7699 ( .A(n3709), .B(n3710), .Z(n3708) );
  OR U7700 ( .A(n3711), .B(n3712), .Z(n3707) );
  ANDN U7701 ( .B(n3713), .A(n3714), .Z(n3600) );
  IV U7702 ( .A(n3715), .Z(n3713) );
  XNOR U7703 ( .A(n3680), .B(n3679), .Z(N29849) );
  XOR U7704 ( .A(n3699), .B(n3698), .Z(n3679) );
  XNOR U7705 ( .A(n3714), .B(n3715), .Z(n3698) );
  XNOR U7706 ( .A(n3709), .B(n3710), .Z(n3715) );
  XNOR U7707 ( .A(n3711), .B(n3712), .Z(n3710) );
  XNOR U7708 ( .A(y[3844]), .B(x[3844]), .Z(n3712) );
  XNOR U7709 ( .A(y[3845]), .B(x[3845]), .Z(n3711) );
  XNOR U7710 ( .A(y[3843]), .B(x[3843]), .Z(n3709) );
  XNOR U7711 ( .A(n3703), .B(n3704), .Z(n3714) );
  XNOR U7712 ( .A(y[3840]), .B(x[3840]), .Z(n3704) );
  XNOR U7713 ( .A(n3705), .B(n3706), .Z(n3703) );
  XNOR U7714 ( .A(y[3841]), .B(x[3841]), .Z(n3706) );
  XNOR U7715 ( .A(y[3842]), .B(x[3842]), .Z(n3705) );
  XNOR U7716 ( .A(n3696), .B(n3695), .Z(n3699) );
  XNOR U7717 ( .A(n3691), .B(n3692), .Z(n3695) );
  XNOR U7718 ( .A(y[3837]), .B(x[3837]), .Z(n3692) );
  XNOR U7719 ( .A(n3693), .B(n3694), .Z(n3691) );
  XNOR U7720 ( .A(y[3838]), .B(x[3838]), .Z(n3694) );
  XNOR U7721 ( .A(y[3839]), .B(x[3839]), .Z(n3693) );
  XNOR U7722 ( .A(n3685), .B(n3686), .Z(n3696) );
  XNOR U7723 ( .A(y[3834]), .B(x[3834]), .Z(n3686) );
  XNOR U7724 ( .A(n3687), .B(n3688), .Z(n3685) );
  XNOR U7725 ( .A(y[3835]), .B(x[3835]), .Z(n3688) );
  XNOR U7726 ( .A(y[3836]), .B(x[3836]), .Z(n3687) );
  XOR U7727 ( .A(n3661), .B(n3662), .Z(n3680) );
  XNOR U7728 ( .A(n3677), .B(n3678), .Z(n3662) );
  XNOR U7729 ( .A(n3672), .B(n3673), .Z(n3678) );
  XNOR U7730 ( .A(n3674), .B(n3675), .Z(n3673) );
  XNOR U7731 ( .A(y[3832]), .B(x[3832]), .Z(n3675) );
  XNOR U7732 ( .A(y[3833]), .B(x[3833]), .Z(n3674) );
  XNOR U7733 ( .A(y[3831]), .B(x[3831]), .Z(n3672) );
  XNOR U7734 ( .A(n3666), .B(n3667), .Z(n3677) );
  XNOR U7735 ( .A(y[3828]), .B(x[3828]), .Z(n3667) );
  XNOR U7736 ( .A(n3668), .B(n3669), .Z(n3666) );
  XNOR U7737 ( .A(y[3829]), .B(x[3829]), .Z(n3669) );
  XNOR U7738 ( .A(y[3830]), .B(x[3830]), .Z(n3668) );
  XOR U7739 ( .A(n3660), .B(n3659), .Z(n3661) );
  XNOR U7740 ( .A(n3655), .B(n3656), .Z(n3659) );
  XNOR U7741 ( .A(y[3825]), .B(x[3825]), .Z(n3656) );
  XNOR U7742 ( .A(n3657), .B(n3658), .Z(n3655) );
  XNOR U7743 ( .A(y[3826]), .B(x[3826]), .Z(n3658) );
  XNOR U7744 ( .A(y[3827]), .B(x[3827]), .Z(n3657) );
  XNOR U7745 ( .A(n3649), .B(n3650), .Z(n3660) );
  XNOR U7746 ( .A(y[3822]), .B(x[3822]), .Z(n3650) );
  XNOR U7747 ( .A(n3651), .B(n3652), .Z(n3649) );
  XNOR U7748 ( .A(y[3823]), .B(x[3823]), .Z(n3652) );
  XNOR U7749 ( .A(y[3824]), .B(x[3824]), .Z(n3651) );
  NAND U7750 ( .A(n3716), .B(n3717), .Z(N29841) );
  NANDN U7751 ( .A(n3718), .B(n3719), .Z(n3717) );
  OR U7752 ( .A(n3720), .B(n3721), .Z(n3719) );
  NAND U7753 ( .A(n3720), .B(n3721), .Z(n3716) );
  XOR U7754 ( .A(n3720), .B(n3722), .Z(N29840) );
  XNOR U7755 ( .A(n3718), .B(n3721), .Z(n3722) );
  AND U7756 ( .A(n3723), .B(n3724), .Z(n3721) );
  NANDN U7757 ( .A(n3725), .B(n3726), .Z(n3724) );
  NANDN U7758 ( .A(n3727), .B(n3728), .Z(n3726) );
  NANDN U7759 ( .A(n3728), .B(n3727), .Z(n3723) );
  NAND U7760 ( .A(n3729), .B(n3730), .Z(n3718) );
  NANDN U7761 ( .A(n3731), .B(n3732), .Z(n3730) );
  OR U7762 ( .A(n3733), .B(n3734), .Z(n3732) );
  NAND U7763 ( .A(n3734), .B(n3733), .Z(n3729) );
  AND U7764 ( .A(n3735), .B(n3736), .Z(n3720) );
  NANDN U7765 ( .A(n3737), .B(n3738), .Z(n3736) );
  NANDN U7766 ( .A(n3739), .B(n3740), .Z(n3738) );
  NANDN U7767 ( .A(n3740), .B(n3739), .Z(n3735) );
  XOR U7768 ( .A(n3734), .B(n3741), .Z(N29839) );
  XOR U7769 ( .A(n3731), .B(n3733), .Z(n3741) );
  XNOR U7770 ( .A(n3727), .B(n3742), .Z(n3733) );
  XNOR U7771 ( .A(n3725), .B(n3728), .Z(n3742) );
  NAND U7772 ( .A(n3743), .B(n3744), .Z(n3728) );
  NAND U7773 ( .A(n3745), .B(n3746), .Z(n3744) );
  OR U7774 ( .A(n3747), .B(n3748), .Z(n3745) );
  NANDN U7775 ( .A(n3749), .B(n3747), .Z(n3743) );
  IV U7776 ( .A(n3748), .Z(n3749) );
  NAND U7777 ( .A(n3750), .B(n3751), .Z(n3725) );
  NAND U7778 ( .A(n3752), .B(n3753), .Z(n3751) );
  NANDN U7779 ( .A(n3754), .B(n3755), .Z(n3752) );
  NANDN U7780 ( .A(n3755), .B(n3754), .Z(n3750) );
  AND U7781 ( .A(n3756), .B(n3757), .Z(n3727) );
  NAND U7782 ( .A(n3758), .B(n3759), .Z(n3757) );
  OR U7783 ( .A(n3760), .B(n3761), .Z(n3758) );
  NANDN U7784 ( .A(n3762), .B(n3760), .Z(n3756) );
  NAND U7785 ( .A(n3763), .B(n3764), .Z(n3731) );
  NANDN U7786 ( .A(n3765), .B(n3766), .Z(n3764) );
  OR U7787 ( .A(n3767), .B(n3768), .Z(n3766) );
  NANDN U7788 ( .A(n3769), .B(n3767), .Z(n3763) );
  IV U7789 ( .A(n3768), .Z(n3769) );
  XNOR U7790 ( .A(n3739), .B(n3770), .Z(n3734) );
  XNOR U7791 ( .A(n3737), .B(n3740), .Z(n3770) );
  NAND U7792 ( .A(n3771), .B(n3772), .Z(n3740) );
  NAND U7793 ( .A(n3773), .B(n3774), .Z(n3772) );
  OR U7794 ( .A(n3775), .B(n3776), .Z(n3773) );
  NANDN U7795 ( .A(n3777), .B(n3775), .Z(n3771) );
  IV U7796 ( .A(n3776), .Z(n3777) );
  NAND U7797 ( .A(n3778), .B(n3779), .Z(n3737) );
  NAND U7798 ( .A(n3780), .B(n3781), .Z(n3779) );
  NANDN U7799 ( .A(n3782), .B(n3783), .Z(n3780) );
  NANDN U7800 ( .A(n3783), .B(n3782), .Z(n3778) );
  AND U7801 ( .A(n3784), .B(n3785), .Z(n3739) );
  NAND U7802 ( .A(n3786), .B(n3787), .Z(n3785) );
  OR U7803 ( .A(n3788), .B(n3789), .Z(n3786) );
  NANDN U7804 ( .A(n3790), .B(n3788), .Z(n3784) );
  XNOR U7805 ( .A(n3765), .B(n3791), .Z(N29838) );
  XOR U7806 ( .A(n3767), .B(n3768), .Z(n3791) );
  XNOR U7807 ( .A(n3781), .B(n3792), .Z(n3768) );
  XOR U7808 ( .A(n3782), .B(n3783), .Z(n3792) );
  XOR U7809 ( .A(n3788), .B(n3793), .Z(n3783) );
  XOR U7810 ( .A(n3787), .B(n3790), .Z(n3793) );
  IV U7811 ( .A(n3789), .Z(n3790) );
  NAND U7812 ( .A(n3794), .B(n3795), .Z(n3789) );
  OR U7813 ( .A(n3796), .B(n3797), .Z(n3795) );
  OR U7814 ( .A(n3798), .B(n3799), .Z(n3794) );
  NAND U7815 ( .A(n3800), .B(n3801), .Z(n3787) );
  OR U7816 ( .A(n3802), .B(n3803), .Z(n3801) );
  OR U7817 ( .A(n3804), .B(n3805), .Z(n3800) );
  NOR U7818 ( .A(n3806), .B(n3807), .Z(n3788) );
  ANDN U7819 ( .B(n3808), .A(n3809), .Z(n3782) );
  XNOR U7820 ( .A(n3775), .B(n3810), .Z(n3781) );
  XNOR U7821 ( .A(n3774), .B(n3776), .Z(n3810) );
  NAND U7822 ( .A(n3811), .B(n3812), .Z(n3776) );
  OR U7823 ( .A(n3813), .B(n3814), .Z(n3812) );
  OR U7824 ( .A(n3815), .B(n3816), .Z(n3811) );
  NAND U7825 ( .A(n3817), .B(n3818), .Z(n3774) );
  OR U7826 ( .A(n3819), .B(n3820), .Z(n3818) );
  OR U7827 ( .A(n3821), .B(n3822), .Z(n3817) );
  ANDN U7828 ( .B(n3823), .A(n3824), .Z(n3775) );
  IV U7829 ( .A(n3825), .Z(n3823) );
  ANDN U7830 ( .B(n3826), .A(n3827), .Z(n3767) );
  XOR U7831 ( .A(n3753), .B(n3828), .Z(n3765) );
  XOR U7832 ( .A(n3754), .B(n3755), .Z(n3828) );
  XOR U7833 ( .A(n3760), .B(n3829), .Z(n3755) );
  XOR U7834 ( .A(n3759), .B(n3762), .Z(n3829) );
  IV U7835 ( .A(n3761), .Z(n3762) );
  NAND U7836 ( .A(n3830), .B(n3831), .Z(n3761) );
  OR U7837 ( .A(n3832), .B(n3833), .Z(n3831) );
  OR U7838 ( .A(n3834), .B(n3835), .Z(n3830) );
  NAND U7839 ( .A(n3836), .B(n3837), .Z(n3759) );
  OR U7840 ( .A(n3838), .B(n3839), .Z(n3837) );
  OR U7841 ( .A(n3840), .B(n3841), .Z(n3836) );
  NOR U7842 ( .A(n3842), .B(n3843), .Z(n3760) );
  ANDN U7843 ( .B(n3844), .A(n3845), .Z(n3754) );
  IV U7844 ( .A(n3846), .Z(n3844) );
  XNOR U7845 ( .A(n3747), .B(n3847), .Z(n3753) );
  XNOR U7846 ( .A(n3746), .B(n3748), .Z(n3847) );
  NAND U7847 ( .A(n3848), .B(n3849), .Z(n3748) );
  OR U7848 ( .A(n3850), .B(n3851), .Z(n3849) );
  OR U7849 ( .A(n3852), .B(n3853), .Z(n3848) );
  NAND U7850 ( .A(n3854), .B(n3855), .Z(n3746) );
  OR U7851 ( .A(n3856), .B(n3857), .Z(n3855) );
  OR U7852 ( .A(n3858), .B(n3859), .Z(n3854) );
  ANDN U7853 ( .B(n3860), .A(n3861), .Z(n3747) );
  IV U7854 ( .A(n3862), .Z(n3860) );
  XNOR U7855 ( .A(n3827), .B(n3826), .Z(N29837) );
  XOR U7856 ( .A(n3846), .B(n3845), .Z(n3826) );
  XNOR U7857 ( .A(n3861), .B(n3862), .Z(n3845) );
  XNOR U7858 ( .A(n3856), .B(n3857), .Z(n3862) );
  XNOR U7859 ( .A(n3858), .B(n3859), .Z(n3857) );
  XNOR U7860 ( .A(y[3820]), .B(x[3820]), .Z(n3859) );
  XNOR U7861 ( .A(y[3821]), .B(x[3821]), .Z(n3858) );
  XNOR U7862 ( .A(y[3819]), .B(x[3819]), .Z(n3856) );
  XNOR U7863 ( .A(n3850), .B(n3851), .Z(n3861) );
  XNOR U7864 ( .A(y[3816]), .B(x[3816]), .Z(n3851) );
  XNOR U7865 ( .A(n3852), .B(n3853), .Z(n3850) );
  XNOR U7866 ( .A(y[3817]), .B(x[3817]), .Z(n3853) );
  XNOR U7867 ( .A(y[3818]), .B(x[3818]), .Z(n3852) );
  XNOR U7868 ( .A(n3843), .B(n3842), .Z(n3846) );
  XNOR U7869 ( .A(n3838), .B(n3839), .Z(n3842) );
  XNOR U7870 ( .A(y[3813]), .B(x[3813]), .Z(n3839) );
  XNOR U7871 ( .A(n3840), .B(n3841), .Z(n3838) );
  XNOR U7872 ( .A(y[3814]), .B(x[3814]), .Z(n3841) );
  XNOR U7873 ( .A(y[3815]), .B(x[3815]), .Z(n3840) );
  XNOR U7874 ( .A(n3832), .B(n3833), .Z(n3843) );
  XNOR U7875 ( .A(y[3810]), .B(x[3810]), .Z(n3833) );
  XNOR U7876 ( .A(n3834), .B(n3835), .Z(n3832) );
  XNOR U7877 ( .A(y[3811]), .B(x[3811]), .Z(n3835) );
  XNOR U7878 ( .A(y[3812]), .B(x[3812]), .Z(n3834) );
  XOR U7879 ( .A(n3808), .B(n3809), .Z(n3827) );
  XNOR U7880 ( .A(n3824), .B(n3825), .Z(n3809) );
  XNOR U7881 ( .A(n3819), .B(n3820), .Z(n3825) );
  XNOR U7882 ( .A(n3821), .B(n3822), .Z(n3820) );
  XNOR U7883 ( .A(y[3808]), .B(x[3808]), .Z(n3822) );
  XNOR U7884 ( .A(y[3809]), .B(x[3809]), .Z(n3821) );
  XNOR U7885 ( .A(y[3807]), .B(x[3807]), .Z(n3819) );
  XNOR U7886 ( .A(n3813), .B(n3814), .Z(n3824) );
  XNOR U7887 ( .A(y[3804]), .B(x[3804]), .Z(n3814) );
  XNOR U7888 ( .A(n3815), .B(n3816), .Z(n3813) );
  XNOR U7889 ( .A(y[3805]), .B(x[3805]), .Z(n3816) );
  XNOR U7890 ( .A(y[3806]), .B(x[3806]), .Z(n3815) );
  XOR U7891 ( .A(n3807), .B(n3806), .Z(n3808) );
  XNOR U7892 ( .A(n3802), .B(n3803), .Z(n3806) );
  XNOR U7893 ( .A(y[3801]), .B(x[3801]), .Z(n3803) );
  XNOR U7894 ( .A(n3804), .B(n3805), .Z(n3802) );
  XNOR U7895 ( .A(y[3802]), .B(x[3802]), .Z(n3805) );
  XNOR U7896 ( .A(y[3803]), .B(x[3803]), .Z(n3804) );
  XNOR U7897 ( .A(n3796), .B(n3797), .Z(n3807) );
  XNOR U7898 ( .A(y[3798]), .B(x[3798]), .Z(n3797) );
  XNOR U7899 ( .A(n3798), .B(n3799), .Z(n3796) );
  XNOR U7900 ( .A(y[3799]), .B(x[3799]), .Z(n3799) );
  XNOR U7901 ( .A(y[3800]), .B(x[3800]), .Z(n3798) );
  NAND U7902 ( .A(n3863), .B(n3864), .Z(N29829) );
  NANDN U7903 ( .A(n3865), .B(n3866), .Z(n3864) );
  OR U7904 ( .A(n3867), .B(n3868), .Z(n3866) );
  NAND U7905 ( .A(n3867), .B(n3868), .Z(n3863) );
  XOR U7906 ( .A(n3867), .B(n3869), .Z(N29828) );
  XNOR U7907 ( .A(n3865), .B(n3868), .Z(n3869) );
  AND U7908 ( .A(n3870), .B(n3871), .Z(n3868) );
  NANDN U7909 ( .A(n3872), .B(n3873), .Z(n3871) );
  NANDN U7910 ( .A(n3874), .B(n3875), .Z(n3873) );
  NANDN U7911 ( .A(n3875), .B(n3874), .Z(n3870) );
  NAND U7912 ( .A(n3876), .B(n3877), .Z(n3865) );
  NANDN U7913 ( .A(n3878), .B(n3879), .Z(n3877) );
  OR U7914 ( .A(n3880), .B(n3881), .Z(n3879) );
  NAND U7915 ( .A(n3881), .B(n3880), .Z(n3876) );
  AND U7916 ( .A(n3882), .B(n3883), .Z(n3867) );
  NANDN U7917 ( .A(n3884), .B(n3885), .Z(n3883) );
  NANDN U7918 ( .A(n3886), .B(n3887), .Z(n3885) );
  NANDN U7919 ( .A(n3887), .B(n3886), .Z(n3882) );
  XOR U7920 ( .A(n3881), .B(n3888), .Z(N29827) );
  XOR U7921 ( .A(n3878), .B(n3880), .Z(n3888) );
  XNOR U7922 ( .A(n3874), .B(n3889), .Z(n3880) );
  XNOR U7923 ( .A(n3872), .B(n3875), .Z(n3889) );
  NAND U7924 ( .A(n3890), .B(n3891), .Z(n3875) );
  NAND U7925 ( .A(n3892), .B(n3893), .Z(n3891) );
  OR U7926 ( .A(n3894), .B(n3895), .Z(n3892) );
  NANDN U7927 ( .A(n3896), .B(n3894), .Z(n3890) );
  IV U7928 ( .A(n3895), .Z(n3896) );
  NAND U7929 ( .A(n3897), .B(n3898), .Z(n3872) );
  NAND U7930 ( .A(n3899), .B(n3900), .Z(n3898) );
  NANDN U7931 ( .A(n3901), .B(n3902), .Z(n3899) );
  NANDN U7932 ( .A(n3902), .B(n3901), .Z(n3897) );
  AND U7933 ( .A(n3903), .B(n3904), .Z(n3874) );
  NAND U7934 ( .A(n3905), .B(n3906), .Z(n3904) );
  OR U7935 ( .A(n3907), .B(n3908), .Z(n3905) );
  NANDN U7936 ( .A(n3909), .B(n3907), .Z(n3903) );
  NAND U7937 ( .A(n3910), .B(n3911), .Z(n3878) );
  NANDN U7938 ( .A(n3912), .B(n3913), .Z(n3911) );
  OR U7939 ( .A(n3914), .B(n3915), .Z(n3913) );
  NANDN U7940 ( .A(n3916), .B(n3914), .Z(n3910) );
  IV U7941 ( .A(n3915), .Z(n3916) );
  XNOR U7942 ( .A(n3886), .B(n3917), .Z(n3881) );
  XNOR U7943 ( .A(n3884), .B(n3887), .Z(n3917) );
  NAND U7944 ( .A(n3918), .B(n3919), .Z(n3887) );
  NAND U7945 ( .A(n3920), .B(n3921), .Z(n3919) );
  OR U7946 ( .A(n3922), .B(n3923), .Z(n3920) );
  NANDN U7947 ( .A(n3924), .B(n3922), .Z(n3918) );
  IV U7948 ( .A(n3923), .Z(n3924) );
  NAND U7949 ( .A(n3925), .B(n3926), .Z(n3884) );
  NAND U7950 ( .A(n3927), .B(n3928), .Z(n3926) );
  NANDN U7951 ( .A(n3929), .B(n3930), .Z(n3927) );
  NANDN U7952 ( .A(n3930), .B(n3929), .Z(n3925) );
  AND U7953 ( .A(n3931), .B(n3932), .Z(n3886) );
  NAND U7954 ( .A(n3933), .B(n3934), .Z(n3932) );
  OR U7955 ( .A(n3935), .B(n3936), .Z(n3933) );
  NANDN U7956 ( .A(n3937), .B(n3935), .Z(n3931) );
  XNOR U7957 ( .A(n3912), .B(n3938), .Z(N29826) );
  XOR U7958 ( .A(n3914), .B(n3915), .Z(n3938) );
  XNOR U7959 ( .A(n3928), .B(n3939), .Z(n3915) );
  XOR U7960 ( .A(n3929), .B(n3930), .Z(n3939) );
  XOR U7961 ( .A(n3935), .B(n3940), .Z(n3930) );
  XOR U7962 ( .A(n3934), .B(n3937), .Z(n3940) );
  IV U7963 ( .A(n3936), .Z(n3937) );
  NAND U7964 ( .A(n3941), .B(n3942), .Z(n3936) );
  OR U7965 ( .A(n3943), .B(n3944), .Z(n3942) );
  OR U7966 ( .A(n3945), .B(n3946), .Z(n3941) );
  NAND U7967 ( .A(n3947), .B(n3948), .Z(n3934) );
  OR U7968 ( .A(n3949), .B(n3950), .Z(n3948) );
  OR U7969 ( .A(n3951), .B(n3952), .Z(n3947) );
  NOR U7970 ( .A(n3953), .B(n3954), .Z(n3935) );
  ANDN U7971 ( .B(n3955), .A(n3956), .Z(n3929) );
  XNOR U7972 ( .A(n3922), .B(n3957), .Z(n3928) );
  XNOR U7973 ( .A(n3921), .B(n3923), .Z(n3957) );
  NAND U7974 ( .A(n3958), .B(n3959), .Z(n3923) );
  OR U7975 ( .A(n3960), .B(n3961), .Z(n3959) );
  OR U7976 ( .A(n3962), .B(n3963), .Z(n3958) );
  NAND U7977 ( .A(n3964), .B(n3965), .Z(n3921) );
  OR U7978 ( .A(n3966), .B(n3967), .Z(n3965) );
  OR U7979 ( .A(n3968), .B(n3969), .Z(n3964) );
  ANDN U7980 ( .B(n3970), .A(n3971), .Z(n3922) );
  IV U7981 ( .A(n3972), .Z(n3970) );
  ANDN U7982 ( .B(n3973), .A(n3974), .Z(n3914) );
  XOR U7983 ( .A(n3900), .B(n3975), .Z(n3912) );
  XOR U7984 ( .A(n3901), .B(n3902), .Z(n3975) );
  XOR U7985 ( .A(n3907), .B(n3976), .Z(n3902) );
  XOR U7986 ( .A(n3906), .B(n3909), .Z(n3976) );
  IV U7987 ( .A(n3908), .Z(n3909) );
  NAND U7988 ( .A(n3977), .B(n3978), .Z(n3908) );
  OR U7989 ( .A(n3979), .B(n3980), .Z(n3978) );
  OR U7990 ( .A(n3981), .B(n3982), .Z(n3977) );
  NAND U7991 ( .A(n3983), .B(n3984), .Z(n3906) );
  OR U7992 ( .A(n3985), .B(n3986), .Z(n3984) );
  OR U7993 ( .A(n3987), .B(n3988), .Z(n3983) );
  NOR U7994 ( .A(n3989), .B(n3990), .Z(n3907) );
  ANDN U7995 ( .B(n3991), .A(n3992), .Z(n3901) );
  IV U7996 ( .A(n3993), .Z(n3991) );
  XNOR U7997 ( .A(n3894), .B(n3994), .Z(n3900) );
  XNOR U7998 ( .A(n3893), .B(n3895), .Z(n3994) );
  NAND U7999 ( .A(n3995), .B(n3996), .Z(n3895) );
  OR U8000 ( .A(n3997), .B(n3998), .Z(n3996) );
  OR U8001 ( .A(n3999), .B(n4000), .Z(n3995) );
  NAND U8002 ( .A(n4001), .B(n4002), .Z(n3893) );
  OR U8003 ( .A(n4003), .B(n4004), .Z(n4002) );
  OR U8004 ( .A(n4005), .B(n4006), .Z(n4001) );
  ANDN U8005 ( .B(n4007), .A(n4008), .Z(n3894) );
  IV U8006 ( .A(n4009), .Z(n4007) );
  XNOR U8007 ( .A(n3974), .B(n3973), .Z(N29825) );
  XOR U8008 ( .A(n3993), .B(n3992), .Z(n3973) );
  XNOR U8009 ( .A(n4008), .B(n4009), .Z(n3992) );
  XNOR U8010 ( .A(n4003), .B(n4004), .Z(n4009) );
  XNOR U8011 ( .A(n4005), .B(n4006), .Z(n4004) );
  XNOR U8012 ( .A(y[3796]), .B(x[3796]), .Z(n4006) );
  XNOR U8013 ( .A(y[3797]), .B(x[3797]), .Z(n4005) );
  XNOR U8014 ( .A(y[3795]), .B(x[3795]), .Z(n4003) );
  XNOR U8015 ( .A(n3997), .B(n3998), .Z(n4008) );
  XNOR U8016 ( .A(y[3792]), .B(x[3792]), .Z(n3998) );
  XNOR U8017 ( .A(n3999), .B(n4000), .Z(n3997) );
  XNOR U8018 ( .A(y[3793]), .B(x[3793]), .Z(n4000) );
  XNOR U8019 ( .A(y[3794]), .B(x[3794]), .Z(n3999) );
  XNOR U8020 ( .A(n3990), .B(n3989), .Z(n3993) );
  XNOR U8021 ( .A(n3985), .B(n3986), .Z(n3989) );
  XNOR U8022 ( .A(y[3789]), .B(x[3789]), .Z(n3986) );
  XNOR U8023 ( .A(n3987), .B(n3988), .Z(n3985) );
  XNOR U8024 ( .A(y[3790]), .B(x[3790]), .Z(n3988) );
  XNOR U8025 ( .A(y[3791]), .B(x[3791]), .Z(n3987) );
  XNOR U8026 ( .A(n3979), .B(n3980), .Z(n3990) );
  XNOR U8027 ( .A(y[3786]), .B(x[3786]), .Z(n3980) );
  XNOR U8028 ( .A(n3981), .B(n3982), .Z(n3979) );
  XNOR U8029 ( .A(y[3787]), .B(x[3787]), .Z(n3982) );
  XNOR U8030 ( .A(y[3788]), .B(x[3788]), .Z(n3981) );
  XOR U8031 ( .A(n3955), .B(n3956), .Z(n3974) );
  XNOR U8032 ( .A(n3971), .B(n3972), .Z(n3956) );
  XNOR U8033 ( .A(n3966), .B(n3967), .Z(n3972) );
  XNOR U8034 ( .A(n3968), .B(n3969), .Z(n3967) );
  XNOR U8035 ( .A(y[3784]), .B(x[3784]), .Z(n3969) );
  XNOR U8036 ( .A(y[3785]), .B(x[3785]), .Z(n3968) );
  XNOR U8037 ( .A(y[3783]), .B(x[3783]), .Z(n3966) );
  XNOR U8038 ( .A(n3960), .B(n3961), .Z(n3971) );
  XNOR U8039 ( .A(y[3780]), .B(x[3780]), .Z(n3961) );
  XNOR U8040 ( .A(n3962), .B(n3963), .Z(n3960) );
  XNOR U8041 ( .A(y[3781]), .B(x[3781]), .Z(n3963) );
  XNOR U8042 ( .A(y[3782]), .B(x[3782]), .Z(n3962) );
  XOR U8043 ( .A(n3954), .B(n3953), .Z(n3955) );
  XNOR U8044 ( .A(n3949), .B(n3950), .Z(n3953) );
  XNOR U8045 ( .A(y[3777]), .B(x[3777]), .Z(n3950) );
  XNOR U8046 ( .A(n3951), .B(n3952), .Z(n3949) );
  XNOR U8047 ( .A(y[3778]), .B(x[3778]), .Z(n3952) );
  XNOR U8048 ( .A(y[3779]), .B(x[3779]), .Z(n3951) );
  XNOR U8049 ( .A(n3943), .B(n3944), .Z(n3954) );
  XNOR U8050 ( .A(y[3774]), .B(x[3774]), .Z(n3944) );
  XNOR U8051 ( .A(n3945), .B(n3946), .Z(n3943) );
  XNOR U8052 ( .A(y[3775]), .B(x[3775]), .Z(n3946) );
  XNOR U8053 ( .A(y[3776]), .B(x[3776]), .Z(n3945) );
  NAND U8054 ( .A(n4010), .B(n4011), .Z(N29817) );
  NANDN U8055 ( .A(n4012), .B(n4013), .Z(n4011) );
  OR U8056 ( .A(n4014), .B(n4015), .Z(n4013) );
  NAND U8057 ( .A(n4014), .B(n4015), .Z(n4010) );
  XOR U8058 ( .A(n4014), .B(n4016), .Z(N29816) );
  XNOR U8059 ( .A(n4012), .B(n4015), .Z(n4016) );
  AND U8060 ( .A(n4017), .B(n4018), .Z(n4015) );
  NANDN U8061 ( .A(n4019), .B(n4020), .Z(n4018) );
  NANDN U8062 ( .A(n4021), .B(n4022), .Z(n4020) );
  NANDN U8063 ( .A(n4022), .B(n4021), .Z(n4017) );
  NAND U8064 ( .A(n4023), .B(n4024), .Z(n4012) );
  NANDN U8065 ( .A(n4025), .B(n4026), .Z(n4024) );
  OR U8066 ( .A(n4027), .B(n4028), .Z(n4026) );
  NAND U8067 ( .A(n4028), .B(n4027), .Z(n4023) );
  AND U8068 ( .A(n4029), .B(n4030), .Z(n4014) );
  NANDN U8069 ( .A(n4031), .B(n4032), .Z(n4030) );
  NANDN U8070 ( .A(n4033), .B(n4034), .Z(n4032) );
  NANDN U8071 ( .A(n4034), .B(n4033), .Z(n4029) );
  XOR U8072 ( .A(n4028), .B(n4035), .Z(N29815) );
  XOR U8073 ( .A(n4025), .B(n4027), .Z(n4035) );
  XNOR U8074 ( .A(n4021), .B(n4036), .Z(n4027) );
  XNOR U8075 ( .A(n4019), .B(n4022), .Z(n4036) );
  NAND U8076 ( .A(n4037), .B(n4038), .Z(n4022) );
  NAND U8077 ( .A(n4039), .B(n4040), .Z(n4038) );
  OR U8078 ( .A(n4041), .B(n4042), .Z(n4039) );
  NANDN U8079 ( .A(n4043), .B(n4041), .Z(n4037) );
  IV U8080 ( .A(n4042), .Z(n4043) );
  NAND U8081 ( .A(n4044), .B(n4045), .Z(n4019) );
  NAND U8082 ( .A(n4046), .B(n4047), .Z(n4045) );
  NANDN U8083 ( .A(n4048), .B(n4049), .Z(n4046) );
  NANDN U8084 ( .A(n4049), .B(n4048), .Z(n4044) );
  AND U8085 ( .A(n4050), .B(n4051), .Z(n4021) );
  NAND U8086 ( .A(n4052), .B(n4053), .Z(n4051) );
  OR U8087 ( .A(n4054), .B(n4055), .Z(n4052) );
  NANDN U8088 ( .A(n4056), .B(n4054), .Z(n4050) );
  NAND U8089 ( .A(n4057), .B(n4058), .Z(n4025) );
  NANDN U8090 ( .A(n4059), .B(n4060), .Z(n4058) );
  OR U8091 ( .A(n4061), .B(n4062), .Z(n4060) );
  NANDN U8092 ( .A(n4063), .B(n4061), .Z(n4057) );
  IV U8093 ( .A(n4062), .Z(n4063) );
  XNOR U8094 ( .A(n4033), .B(n4064), .Z(n4028) );
  XNOR U8095 ( .A(n4031), .B(n4034), .Z(n4064) );
  NAND U8096 ( .A(n4065), .B(n4066), .Z(n4034) );
  NAND U8097 ( .A(n4067), .B(n4068), .Z(n4066) );
  OR U8098 ( .A(n4069), .B(n4070), .Z(n4067) );
  NANDN U8099 ( .A(n4071), .B(n4069), .Z(n4065) );
  IV U8100 ( .A(n4070), .Z(n4071) );
  NAND U8101 ( .A(n4072), .B(n4073), .Z(n4031) );
  NAND U8102 ( .A(n4074), .B(n4075), .Z(n4073) );
  NANDN U8103 ( .A(n4076), .B(n4077), .Z(n4074) );
  NANDN U8104 ( .A(n4077), .B(n4076), .Z(n4072) );
  AND U8105 ( .A(n4078), .B(n4079), .Z(n4033) );
  NAND U8106 ( .A(n4080), .B(n4081), .Z(n4079) );
  OR U8107 ( .A(n4082), .B(n4083), .Z(n4080) );
  NANDN U8108 ( .A(n4084), .B(n4082), .Z(n4078) );
  XNOR U8109 ( .A(n4059), .B(n4085), .Z(N29814) );
  XOR U8110 ( .A(n4061), .B(n4062), .Z(n4085) );
  XNOR U8111 ( .A(n4075), .B(n4086), .Z(n4062) );
  XOR U8112 ( .A(n4076), .B(n4077), .Z(n4086) );
  XOR U8113 ( .A(n4082), .B(n4087), .Z(n4077) );
  XOR U8114 ( .A(n4081), .B(n4084), .Z(n4087) );
  IV U8115 ( .A(n4083), .Z(n4084) );
  NAND U8116 ( .A(n4088), .B(n4089), .Z(n4083) );
  OR U8117 ( .A(n4090), .B(n4091), .Z(n4089) );
  OR U8118 ( .A(n4092), .B(n4093), .Z(n4088) );
  NAND U8119 ( .A(n4094), .B(n4095), .Z(n4081) );
  OR U8120 ( .A(n4096), .B(n4097), .Z(n4095) );
  OR U8121 ( .A(n4098), .B(n4099), .Z(n4094) );
  NOR U8122 ( .A(n4100), .B(n4101), .Z(n4082) );
  ANDN U8123 ( .B(n4102), .A(n4103), .Z(n4076) );
  XNOR U8124 ( .A(n4069), .B(n4104), .Z(n4075) );
  XNOR U8125 ( .A(n4068), .B(n4070), .Z(n4104) );
  NAND U8126 ( .A(n4105), .B(n4106), .Z(n4070) );
  OR U8127 ( .A(n4107), .B(n4108), .Z(n4106) );
  OR U8128 ( .A(n4109), .B(n4110), .Z(n4105) );
  NAND U8129 ( .A(n4111), .B(n4112), .Z(n4068) );
  OR U8130 ( .A(n4113), .B(n4114), .Z(n4112) );
  OR U8131 ( .A(n4115), .B(n4116), .Z(n4111) );
  ANDN U8132 ( .B(n4117), .A(n4118), .Z(n4069) );
  IV U8133 ( .A(n4119), .Z(n4117) );
  ANDN U8134 ( .B(n4120), .A(n4121), .Z(n4061) );
  XOR U8135 ( .A(n4047), .B(n4122), .Z(n4059) );
  XOR U8136 ( .A(n4048), .B(n4049), .Z(n4122) );
  XOR U8137 ( .A(n4054), .B(n4123), .Z(n4049) );
  XOR U8138 ( .A(n4053), .B(n4056), .Z(n4123) );
  IV U8139 ( .A(n4055), .Z(n4056) );
  NAND U8140 ( .A(n4124), .B(n4125), .Z(n4055) );
  OR U8141 ( .A(n4126), .B(n4127), .Z(n4125) );
  OR U8142 ( .A(n4128), .B(n4129), .Z(n4124) );
  NAND U8143 ( .A(n4130), .B(n4131), .Z(n4053) );
  OR U8144 ( .A(n4132), .B(n4133), .Z(n4131) );
  OR U8145 ( .A(n4134), .B(n4135), .Z(n4130) );
  NOR U8146 ( .A(n4136), .B(n4137), .Z(n4054) );
  ANDN U8147 ( .B(n4138), .A(n4139), .Z(n4048) );
  IV U8148 ( .A(n4140), .Z(n4138) );
  XNOR U8149 ( .A(n4041), .B(n4141), .Z(n4047) );
  XNOR U8150 ( .A(n4040), .B(n4042), .Z(n4141) );
  NAND U8151 ( .A(n4142), .B(n4143), .Z(n4042) );
  OR U8152 ( .A(n4144), .B(n4145), .Z(n4143) );
  OR U8153 ( .A(n4146), .B(n4147), .Z(n4142) );
  NAND U8154 ( .A(n4148), .B(n4149), .Z(n4040) );
  OR U8155 ( .A(n4150), .B(n4151), .Z(n4149) );
  OR U8156 ( .A(n4152), .B(n4153), .Z(n4148) );
  ANDN U8157 ( .B(n4154), .A(n4155), .Z(n4041) );
  IV U8158 ( .A(n4156), .Z(n4154) );
  XNOR U8159 ( .A(n4121), .B(n4120), .Z(N29813) );
  XOR U8160 ( .A(n4140), .B(n4139), .Z(n4120) );
  XNOR U8161 ( .A(n4155), .B(n4156), .Z(n4139) );
  XNOR U8162 ( .A(n4150), .B(n4151), .Z(n4156) );
  XNOR U8163 ( .A(n4152), .B(n4153), .Z(n4151) );
  XNOR U8164 ( .A(y[3772]), .B(x[3772]), .Z(n4153) );
  XNOR U8165 ( .A(y[3773]), .B(x[3773]), .Z(n4152) );
  XNOR U8166 ( .A(y[3771]), .B(x[3771]), .Z(n4150) );
  XNOR U8167 ( .A(n4144), .B(n4145), .Z(n4155) );
  XNOR U8168 ( .A(y[3768]), .B(x[3768]), .Z(n4145) );
  XNOR U8169 ( .A(n4146), .B(n4147), .Z(n4144) );
  XNOR U8170 ( .A(y[3769]), .B(x[3769]), .Z(n4147) );
  XNOR U8171 ( .A(y[3770]), .B(x[3770]), .Z(n4146) );
  XNOR U8172 ( .A(n4137), .B(n4136), .Z(n4140) );
  XNOR U8173 ( .A(n4132), .B(n4133), .Z(n4136) );
  XNOR U8174 ( .A(y[3765]), .B(x[3765]), .Z(n4133) );
  XNOR U8175 ( .A(n4134), .B(n4135), .Z(n4132) );
  XNOR U8176 ( .A(y[3766]), .B(x[3766]), .Z(n4135) );
  XNOR U8177 ( .A(y[3767]), .B(x[3767]), .Z(n4134) );
  XNOR U8178 ( .A(n4126), .B(n4127), .Z(n4137) );
  XNOR U8179 ( .A(y[3762]), .B(x[3762]), .Z(n4127) );
  XNOR U8180 ( .A(n4128), .B(n4129), .Z(n4126) );
  XNOR U8181 ( .A(y[3763]), .B(x[3763]), .Z(n4129) );
  XNOR U8182 ( .A(y[3764]), .B(x[3764]), .Z(n4128) );
  XOR U8183 ( .A(n4102), .B(n4103), .Z(n4121) );
  XNOR U8184 ( .A(n4118), .B(n4119), .Z(n4103) );
  XNOR U8185 ( .A(n4113), .B(n4114), .Z(n4119) );
  XNOR U8186 ( .A(n4115), .B(n4116), .Z(n4114) );
  XNOR U8187 ( .A(y[3760]), .B(x[3760]), .Z(n4116) );
  XNOR U8188 ( .A(y[3761]), .B(x[3761]), .Z(n4115) );
  XNOR U8189 ( .A(y[3759]), .B(x[3759]), .Z(n4113) );
  XNOR U8190 ( .A(n4107), .B(n4108), .Z(n4118) );
  XNOR U8191 ( .A(y[3756]), .B(x[3756]), .Z(n4108) );
  XNOR U8192 ( .A(n4109), .B(n4110), .Z(n4107) );
  XNOR U8193 ( .A(y[3757]), .B(x[3757]), .Z(n4110) );
  XNOR U8194 ( .A(y[3758]), .B(x[3758]), .Z(n4109) );
  XOR U8195 ( .A(n4101), .B(n4100), .Z(n4102) );
  XNOR U8196 ( .A(n4096), .B(n4097), .Z(n4100) );
  XNOR U8197 ( .A(y[3753]), .B(x[3753]), .Z(n4097) );
  XNOR U8198 ( .A(n4098), .B(n4099), .Z(n4096) );
  XNOR U8199 ( .A(y[3754]), .B(x[3754]), .Z(n4099) );
  XNOR U8200 ( .A(y[3755]), .B(x[3755]), .Z(n4098) );
  XNOR U8201 ( .A(n4090), .B(n4091), .Z(n4101) );
  XNOR U8202 ( .A(y[3750]), .B(x[3750]), .Z(n4091) );
  XNOR U8203 ( .A(n4092), .B(n4093), .Z(n4090) );
  XNOR U8204 ( .A(y[3751]), .B(x[3751]), .Z(n4093) );
  XNOR U8205 ( .A(y[3752]), .B(x[3752]), .Z(n4092) );
  NAND U8206 ( .A(n4157), .B(n4158), .Z(N29805) );
  NANDN U8207 ( .A(n4159), .B(n4160), .Z(n4158) );
  OR U8208 ( .A(n4161), .B(n4162), .Z(n4160) );
  NAND U8209 ( .A(n4161), .B(n4162), .Z(n4157) );
  XOR U8210 ( .A(n4161), .B(n4163), .Z(N29804) );
  XNOR U8211 ( .A(n4159), .B(n4162), .Z(n4163) );
  AND U8212 ( .A(n4164), .B(n4165), .Z(n4162) );
  NANDN U8213 ( .A(n4166), .B(n4167), .Z(n4165) );
  NANDN U8214 ( .A(n4168), .B(n4169), .Z(n4167) );
  NANDN U8215 ( .A(n4169), .B(n4168), .Z(n4164) );
  NAND U8216 ( .A(n4170), .B(n4171), .Z(n4159) );
  NANDN U8217 ( .A(n4172), .B(n4173), .Z(n4171) );
  OR U8218 ( .A(n4174), .B(n4175), .Z(n4173) );
  NAND U8219 ( .A(n4175), .B(n4174), .Z(n4170) );
  AND U8220 ( .A(n4176), .B(n4177), .Z(n4161) );
  NANDN U8221 ( .A(n4178), .B(n4179), .Z(n4177) );
  NANDN U8222 ( .A(n4180), .B(n4181), .Z(n4179) );
  NANDN U8223 ( .A(n4181), .B(n4180), .Z(n4176) );
  XOR U8224 ( .A(n4175), .B(n4182), .Z(N29803) );
  XOR U8225 ( .A(n4172), .B(n4174), .Z(n4182) );
  XNOR U8226 ( .A(n4168), .B(n4183), .Z(n4174) );
  XNOR U8227 ( .A(n4166), .B(n4169), .Z(n4183) );
  NAND U8228 ( .A(n4184), .B(n4185), .Z(n4169) );
  NAND U8229 ( .A(n4186), .B(n4187), .Z(n4185) );
  OR U8230 ( .A(n4188), .B(n4189), .Z(n4186) );
  NANDN U8231 ( .A(n4190), .B(n4188), .Z(n4184) );
  IV U8232 ( .A(n4189), .Z(n4190) );
  NAND U8233 ( .A(n4191), .B(n4192), .Z(n4166) );
  NAND U8234 ( .A(n4193), .B(n4194), .Z(n4192) );
  NANDN U8235 ( .A(n4195), .B(n4196), .Z(n4193) );
  NANDN U8236 ( .A(n4196), .B(n4195), .Z(n4191) );
  AND U8237 ( .A(n4197), .B(n4198), .Z(n4168) );
  NAND U8238 ( .A(n4199), .B(n4200), .Z(n4198) );
  OR U8239 ( .A(n4201), .B(n4202), .Z(n4199) );
  NANDN U8240 ( .A(n4203), .B(n4201), .Z(n4197) );
  NAND U8241 ( .A(n4204), .B(n4205), .Z(n4172) );
  NANDN U8242 ( .A(n4206), .B(n4207), .Z(n4205) );
  OR U8243 ( .A(n4208), .B(n4209), .Z(n4207) );
  NANDN U8244 ( .A(n4210), .B(n4208), .Z(n4204) );
  IV U8245 ( .A(n4209), .Z(n4210) );
  XNOR U8246 ( .A(n4180), .B(n4211), .Z(n4175) );
  XNOR U8247 ( .A(n4178), .B(n4181), .Z(n4211) );
  NAND U8248 ( .A(n4212), .B(n4213), .Z(n4181) );
  NAND U8249 ( .A(n4214), .B(n4215), .Z(n4213) );
  OR U8250 ( .A(n4216), .B(n4217), .Z(n4214) );
  NANDN U8251 ( .A(n4218), .B(n4216), .Z(n4212) );
  IV U8252 ( .A(n4217), .Z(n4218) );
  NAND U8253 ( .A(n4219), .B(n4220), .Z(n4178) );
  NAND U8254 ( .A(n4221), .B(n4222), .Z(n4220) );
  NANDN U8255 ( .A(n4223), .B(n4224), .Z(n4221) );
  NANDN U8256 ( .A(n4224), .B(n4223), .Z(n4219) );
  AND U8257 ( .A(n4225), .B(n4226), .Z(n4180) );
  NAND U8258 ( .A(n4227), .B(n4228), .Z(n4226) );
  OR U8259 ( .A(n4229), .B(n4230), .Z(n4227) );
  NANDN U8260 ( .A(n4231), .B(n4229), .Z(n4225) );
  XNOR U8261 ( .A(n4206), .B(n4232), .Z(N29802) );
  XOR U8262 ( .A(n4208), .B(n4209), .Z(n4232) );
  XNOR U8263 ( .A(n4222), .B(n4233), .Z(n4209) );
  XOR U8264 ( .A(n4223), .B(n4224), .Z(n4233) );
  XOR U8265 ( .A(n4229), .B(n4234), .Z(n4224) );
  XOR U8266 ( .A(n4228), .B(n4231), .Z(n4234) );
  IV U8267 ( .A(n4230), .Z(n4231) );
  NAND U8268 ( .A(n4235), .B(n4236), .Z(n4230) );
  OR U8269 ( .A(n4237), .B(n4238), .Z(n4236) );
  OR U8270 ( .A(n4239), .B(n4240), .Z(n4235) );
  NAND U8271 ( .A(n4241), .B(n4242), .Z(n4228) );
  OR U8272 ( .A(n4243), .B(n4244), .Z(n4242) );
  OR U8273 ( .A(n4245), .B(n4246), .Z(n4241) );
  NOR U8274 ( .A(n4247), .B(n4248), .Z(n4229) );
  ANDN U8275 ( .B(n4249), .A(n4250), .Z(n4223) );
  XNOR U8276 ( .A(n4216), .B(n4251), .Z(n4222) );
  XNOR U8277 ( .A(n4215), .B(n4217), .Z(n4251) );
  NAND U8278 ( .A(n4252), .B(n4253), .Z(n4217) );
  OR U8279 ( .A(n4254), .B(n4255), .Z(n4253) );
  OR U8280 ( .A(n4256), .B(n4257), .Z(n4252) );
  NAND U8281 ( .A(n4258), .B(n4259), .Z(n4215) );
  OR U8282 ( .A(n4260), .B(n4261), .Z(n4259) );
  OR U8283 ( .A(n4262), .B(n4263), .Z(n4258) );
  ANDN U8284 ( .B(n4264), .A(n4265), .Z(n4216) );
  IV U8285 ( .A(n4266), .Z(n4264) );
  ANDN U8286 ( .B(n4267), .A(n4268), .Z(n4208) );
  XOR U8287 ( .A(n4194), .B(n4269), .Z(n4206) );
  XOR U8288 ( .A(n4195), .B(n4196), .Z(n4269) );
  XOR U8289 ( .A(n4201), .B(n4270), .Z(n4196) );
  XOR U8290 ( .A(n4200), .B(n4203), .Z(n4270) );
  IV U8291 ( .A(n4202), .Z(n4203) );
  NAND U8292 ( .A(n4271), .B(n4272), .Z(n4202) );
  OR U8293 ( .A(n4273), .B(n4274), .Z(n4272) );
  OR U8294 ( .A(n4275), .B(n4276), .Z(n4271) );
  NAND U8295 ( .A(n4277), .B(n4278), .Z(n4200) );
  OR U8296 ( .A(n4279), .B(n4280), .Z(n4278) );
  OR U8297 ( .A(n4281), .B(n4282), .Z(n4277) );
  NOR U8298 ( .A(n4283), .B(n4284), .Z(n4201) );
  ANDN U8299 ( .B(n4285), .A(n4286), .Z(n4195) );
  IV U8300 ( .A(n4287), .Z(n4285) );
  XNOR U8301 ( .A(n4188), .B(n4288), .Z(n4194) );
  XNOR U8302 ( .A(n4187), .B(n4189), .Z(n4288) );
  NAND U8303 ( .A(n4289), .B(n4290), .Z(n4189) );
  OR U8304 ( .A(n4291), .B(n4292), .Z(n4290) );
  OR U8305 ( .A(n4293), .B(n4294), .Z(n4289) );
  NAND U8306 ( .A(n4295), .B(n4296), .Z(n4187) );
  OR U8307 ( .A(n4297), .B(n4298), .Z(n4296) );
  OR U8308 ( .A(n4299), .B(n4300), .Z(n4295) );
  ANDN U8309 ( .B(n4301), .A(n4302), .Z(n4188) );
  IV U8310 ( .A(n4303), .Z(n4301) );
  XNOR U8311 ( .A(n4268), .B(n4267), .Z(N29801) );
  XOR U8312 ( .A(n4287), .B(n4286), .Z(n4267) );
  XNOR U8313 ( .A(n4302), .B(n4303), .Z(n4286) );
  XNOR U8314 ( .A(n4297), .B(n4298), .Z(n4303) );
  XNOR U8315 ( .A(n4299), .B(n4300), .Z(n4298) );
  XNOR U8316 ( .A(y[3748]), .B(x[3748]), .Z(n4300) );
  XNOR U8317 ( .A(y[3749]), .B(x[3749]), .Z(n4299) );
  XNOR U8318 ( .A(y[3747]), .B(x[3747]), .Z(n4297) );
  XNOR U8319 ( .A(n4291), .B(n4292), .Z(n4302) );
  XNOR U8320 ( .A(y[3744]), .B(x[3744]), .Z(n4292) );
  XNOR U8321 ( .A(n4293), .B(n4294), .Z(n4291) );
  XNOR U8322 ( .A(y[3745]), .B(x[3745]), .Z(n4294) );
  XNOR U8323 ( .A(y[3746]), .B(x[3746]), .Z(n4293) );
  XNOR U8324 ( .A(n4284), .B(n4283), .Z(n4287) );
  XNOR U8325 ( .A(n4279), .B(n4280), .Z(n4283) );
  XNOR U8326 ( .A(y[3741]), .B(x[3741]), .Z(n4280) );
  XNOR U8327 ( .A(n4281), .B(n4282), .Z(n4279) );
  XNOR U8328 ( .A(y[3742]), .B(x[3742]), .Z(n4282) );
  XNOR U8329 ( .A(y[3743]), .B(x[3743]), .Z(n4281) );
  XNOR U8330 ( .A(n4273), .B(n4274), .Z(n4284) );
  XNOR U8331 ( .A(y[3738]), .B(x[3738]), .Z(n4274) );
  XNOR U8332 ( .A(n4275), .B(n4276), .Z(n4273) );
  XNOR U8333 ( .A(y[3739]), .B(x[3739]), .Z(n4276) );
  XNOR U8334 ( .A(y[3740]), .B(x[3740]), .Z(n4275) );
  XOR U8335 ( .A(n4249), .B(n4250), .Z(n4268) );
  XNOR U8336 ( .A(n4265), .B(n4266), .Z(n4250) );
  XNOR U8337 ( .A(n4260), .B(n4261), .Z(n4266) );
  XNOR U8338 ( .A(n4262), .B(n4263), .Z(n4261) );
  XNOR U8339 ( .A(y[3736]), .B(x[3736]), .Z(n4263) );
  XNOR U8340 ( .A(y[3737]), .B(x[3737]), .Z(n4262) );
  XNOR U8341 ( .A(y[3735]), .B(x[3735]), .Z(n4260) );
  XNOR U8342 ( .A(n4254), .B(n4255), .Z(n4265) );
  XNOR U8343 ( .A(y[3732]), .B(x[3732]), .Z(n4255) );
  XNOR U8344 ( .A(n4256), .B(n4257), .Z(n4254) );
  XNOR U8345 ( .A(y[3733]), .B(x[3733]), .Z(n4257) );
  XNOR U8346 ( .A(y[3734]), .B(x[3734]), .Z(n4256) );
  XOR U8347 ( .A(n4248), .B(n4247), .Z(n4249) );
  XNOR U8348 ( .A(n4243), .B(n4244), .Z(n4247) );
  XNOR U8349 ( .A(y[3729]), .B(x[3729]), .Z(n4244) );
  XNOR U8350 ( .A(n4245), .B(n4246), .Z(n4243) );
  XNOR U8351 ( .A(y[3730]), .B(x[3730]), .Z(n4246) );
  XNOR U8352 ( .A(y[3731]), .B(x[3731]), .Z(n4245) );
  XNOR U8353 ( .A(n4237), .B(n4238), .Z(n4248) );
  XNOR U8354 ( .A(y[3726]), .B(x[3726]), .Z(n4238) );
  XNOR U8355 ( .A(n4239), .B(n4240), .Z(n4237) );
  XNOR U8356 ( .A(y[3727]), .B(x[3727]), .Z(n4240) );
  XNOR U8357 ( .A(y[3728]), .B(x[3728]), .Z(n4239) );
  NAND U8358 ( .A(n4304), .B(n4305), .Z(N29793) );
  NANDN U8359 ( .A(n4306), .B(n4307), .Z(n4305) );
  OR U8360 ( .A(n4308), .B(n4309), .Z(n4307) );
  NAND U8361 ( .A(n4308), .B(n4309), .Z(n4304) );
  XOR U8362 ( .A(n4308), .B(n4310), .Z(N29792) );
  XNOR U8363 ( .A(n4306), .B(n4309), .Z(n4310) );
  AND U8364 ( .A(n4311), .B(n4312), .Z(n4309) );
  NANDN U8365 ( .A(n4313), .B(n4314), .Z(n4312) );
  NANDN U8366 ( .A(n4315), .B(n4316), .Z(n4314) );
  NANDN U8367 ( .A(n4316), .B(n4315), .Z(n4311) );
  NAND U8368 ( .A(n4317), .B(n4318), .Z(n4306) );
  NANDN U8369 ( .A(n4319), .B(n4320), .Z(n4318) );
  OR U8370 ( .A(n4321), .B(n4322), .Z(n4320) );
  NAND U8371 ( .A(n4322), .B(n4321), .Z(n4317) );
  AND U8372 ( .A(n4323), .B(n4324), .Z(n4308) );
  NANDN U8373 ( .A(n4325), .B(n4326), .Z(n4324) );
  NANDN U8374 ( .A(n4327), .B(n4328), .Z(n4326) );
  NANDN U8375 ( .A(n4328), .B(n4327), .Z(n4323) );
  XOR U8376 ( .A(n4322), .B(n4329), .Z(N29791) );
  XOR U8377 ( .A(n4319), .B(n4321), .Z(n4329) );
  XNOR U8378 ( .A(n4315), .B(n4330), .Z(n4321) );
  XNOR U8379 ( .A(n4313), .B(n4316), .Z(n4330) );
  NAND U8380 ( .A(n4331), .B(n4332), .Z(n4316) );
  NAND U8381 ( .A(n4333), .B(n4334), .Z(n4332) );
  OR U8382 ( .A(n4335), .B(n4336), .Z(n4333) );
  NANDN U8383 ( .A(n4337), .B(n4335), .Z(n4331) );
  IV U8384 ( .A(n4336), .Z(n4337) );
  NAND U8385 ( .A(n4338), .B(n4339), .Z(n4313) );
  NAND U8386 ( .A(n4340), .B(n4341), .Z(n4339) );
  NANDN U8387 ( .A(n4342), .B(n4343), .Z(n4340) );
  NANDN U8388 ( .A(n4343), .B(n4342), .Z(n4338) );
  AND U8389 ( .A(n4344), .B(n4345), .Z(n4315) );
  NAND U8390 ( .A(n4346), .B(n4347), .Z(n4345) );
  OR U8391 ( .A(n4348), .B(n4349), .Z(n4346) );
  NANDN U8392 ( .A(n4350), .B(n4348), .Z(n4344) );
  NAND U8393 ( .A(n4351), .B(n4352), .Z(n4319) );
  NANDN U8394 ( .A(n4353), .B(n4354), .Z(n4352) );
  OR U8395 ( .A(n4355), .B(n4356), .Z(n4354) );
  NANDN U8396 ( .A(n4357), .B(n4355), .Z(n4351) );
  IV U8397 ( .A(n4356), .Z(n4357) );
  XNOR U8398 ( .A(n4327), .B(n4358), .Z(n4322) );
  XNOR U8399 ( .A(n4325), .B(n4328), .Z(n4358) );
  NAND U8400 ( .A(n4359), .B(n4360), .Z(n4328) );
  NAND U8401 ( .A(n4361), .B(n4362), .Z(n4360) );
  OR U8402 ( .A(n4363), .B(n4364), .Z(n4361) );
  NANDN U8403 ( .A(n4365), .B(n4363), .Z(n4359) );
  IV U8404 ( .A(n4364), .Z(n4365) );
  NAND U8405 ( .A(n4366), .B(n4367), .Z(n4325) );
  NAND U8406 ( .A(n4368), .B(n4369), .Z(n4367) );
  NANDN U8407 ( .A(n4370), .B(n4371), .Z(n4368) );
  NANDN U8408 ( .A(n4371), .B(n4370), .Z(n4366) );
  AND U8409 ( .A(n4372), .B(n4373), .Z(n4327) );
  NAND U8410 ( .A(n4374), .B(n4375), .Z(n4373) );
  OR U8411 ( .A(n4376), .B(n4377), .Z(n4374) );
  NANDN U8412 ( .A(n4378), .B(n4376), .Z(n4372) );
  XNOR U8413 ( .A(n4353), .B(n4379), .Z(N29790) );
  XOR U8414 ( .A(n4355), .B(n4356), .Z(n4379) );
  XNOR U8415 ( .A(n4369), .B(n4380), .Z(n4356) );
  XOR U8416 ( .A(n4370), .B(n4371), .Z(n4380) );
  XOR U8417 ( .A(n4376), .B(n4381), .Z(n4371) );
  XOR U8418 ( .A(n4375), .B(n4378), .Z(n4381) );
  IV U8419 ( .A(n4377), .Z(n4378) );
  NAND U8420 ( .A(n4382), .B(n4383), .Z(n4377) );
  OR U8421 ( .A(n4384), .B(n4385), .Z(n4383) );
  OR U8422 ( .A(n4386), .B(n4387), .Z(n4382) );
  NAND U8423 ( .A(n4388), .B(n4389), .Z(n4375) );
  OR U8424 ( .A(n4390), .B(n4391), .Z(n4389) );
  OR U8425 ( .A(n4392), .B(n4393), .Z(n4388) );
  NOR U8426 ( .A(n4394), .B(n4395), .Z(n4376) );
  ANDN U8427 ( .B(n4396), .A(n4397), .Z(n4370) );
  XNOR U8428 ( .A(n4363), .B(n4398), .Z(n4369) );
  XNOR U8429 ( .A(n4362), .B(n4364), .Z(n4398) );
  NAND U8430 ( .A(n4399), .B(n4400), .Z(n4364) );
  OR U8431 ( .A(n4401), .B(n4402), .Z(n4400) );
  OR U8432 ( .A(n4403), .B(n4404), .Z(n4399) );
  NAND U8433 ( .A(n4405), .B(n4406), .Z(n4362) );
  OR U8434 ( .A(n4407), .B(n4408), .Z(n4406) );
  OR U8435 ( .A(n4409), .B(n4410), .Z(n4405) );
  ANDN U8436 ( .B(n4411), .A(n4412), .Z(n4363) );
  IV U8437 ( .A(n4413), .Z(n4411) );
  ANDN U8438 ( .B(n4414), .A(n4415), .Z(n4355) );
  XOR U8439 ( .A(n4341), .B(n4416), .Z(n4353) );
  XOR U8440 ( .A(n4342), .B(n4343), .Z(n4416) );
  XOR U8441 ( .A(n4348), .B(n4417), .Z(n4343) );
  XOR U8442 ( .A(n4347), .B(n4350), .Z(n4417) );
  IV U8443 ( .A(n4349), .Z(n4350) );
  NAND U8444 ( .A(n4418), .B(n4419), .Z(n4349) );
  OR U8445 ( .A(n4420), .B(n4421), .Z(n4419) );
  OR U8446 ( .A(n4422), .B(n4423), .Z(n4418) );
  NAND U8447 ( .A(n4424), .B(n4425), .Z(n4347) );
  OR U8448 ( .A(n4426), .B(n4427), .Z(n4425) );
  OR U8449 ( .A(n4428), .B(n4429), .Z(n4424) );
  NOR U8450 ( .A(n4430), .B(n4431), .Z(n4348) );
  ANDN U8451 ( .B(n4432), .A(n4433), .Z(n4342) );
  IV U8452 ( .A(n4434), .Z(n4432) );
  XNOR U8453 ( .A(n4335), .B(n4435), .Z(n4341) );
  XNOR U8454 ( .A(n4334), .B(n4336), .Z(n4435) );
  NAND U8455 ( .A(n4436), .B(n4437), .Z(n4336) );
  OR U8456 ( .A(n4438), .B(n4439), .Z(n4437) );
  OR U8457 ( .A(n4440), .B(n4441), .Z(n4436) );
  NAND U8458 ( .A(n4442), .B(n4443), .Z(n4334) );
  OR U8459 ( .A(n4444), .B(n4445), .Z(n4443) );
  OR U8460 ( .A(n4446), .B(n4447), .Z(n4442) );
  ANDN U8461 ( .B(n4448), .A(n4449), .Z(n4335) );
  IV U8462 ( .A(n4450), .Z(n4448) );
  XNOR U8463 ( .A(n4415), .B(n4414), .Z(N29789) );
  XOR U8464 ( .A(n4434), .B(n4433), .Z(n4414) );
  XNOR U8465 ( .A(n4449), .B(n4450), .Z(n4433) );
  XNOR U8466 ( .A(n4444), .B(n4445), .Z(n4450) );
  XNOR U8467 ( .A(n4446), .B(n4447), .Z(n4445) );
  XNOR U8468 ( .A(y[3724]), .B(x[3724]), .Z(n4447) );
  XNOR U8469 ( .A(y[3725]), .B(x[3725]), .Z(n4446) );
  XNOR U8470 ( .A(y[3723]), .B(x[3723]), .Z(n4444) );
  XNOR U8471 ( .A(n4438), .B(n4439), .Z(n4449) );
  XNOR U8472 ( .A(y[3720]), .B(x[3720]), .Z(n4439) );
  XNOR U8473 ( .A(n4440), .B(n4441), .Z(n4438) );
  XNOR U8474 ( .A(y[3721]), .B(x[3721]), .Z(n4441) );
  XNOR U8475 ( .A(y[3722]), .B(x[3722]), .Z(n4440) );
  XNOR U8476 ( .A(n4431), .B(n4430), .Z(n4434) );
  XNOR U8477 ( .A(n4426), .B(n4427), .Z(n4430) );
  XNOR U8478 ( .A(y[3717]), .B(x[3717]), .Z(n4427) );
  XNOR U8479 ( .A(n4428), .B(n4429), .Z(n4426) );
  XNOR U8480 ( .A(y[3718]), .B(x[3718]), .Z(n4429) );
  XNOR U8481 ( .A(y[3719]), .B(x[3719]), .Z(n4428) );
  XNOR U8482 ( .A(n4420), .B(n4421), .Z(n4431) );
  XNOR U8483 ( .A(y[3714]), .B(x[3714]), .Z(n4421) );
  XNOR U8484 ( .A(n4422), .B(n4423), .Z(n4420) );
  XNOR U8485 ( .A(y[3715]), .B(x[3715]), .Z(n4423) );
  XNOR U8486 ( .A(y[3716]), .B(x[3716]), .Z(n4422) );
  XOR U8487 ( .A(n4396), .B(n4397), .Z(n4415) );
  XNOR U8488 ( .A(n4412), .B(n4413), .Z(n4397) );
  XNOR U8489 ( .A(n4407), .B(n4408), .Z(n4413) );
  XNOR U8490 ( .A(n4409), .B(n4410), .Z(n4408) );
  XNOR U8491 ( .A(y[3712]), .B(x[3712]), .Z(n4410) );
  XNOR U8492 ( .A(y[3713]), .B(x[3713]), .Z(n4409) );
  XNOR U8493 ( .A(y[3711]), .B(x[3711]), .Z(n4407) );
  XNOR U8494 ( .A(n4401), .B(n4402), .Z(n4412) );
  XNOR U8495 ( .A(y[3708]), .B(x[3708]), .Z(n4402) );
  XNOR U8496 ( .A(n4403), .B(n4404), .Z(n4401) );
  XNOR U8497 ( .A(y[3709]), .B(x[3709]), .Z(n4404) );
  XNOR U8498 ( .A(y[3710]), .B(x[3710]), .Z(n4403) );
  XOR U8499 ( .A(n4395), .B(n4394), .Z(n4396) );
  XNOR U8500 ( .A(n4390), .B(n4391), .Z(n4394) );
  XNOR U8501 ( .A(y[3705]), .B(x[3705]), .Z(n4391) );
  XNOR U8502 ( .A(n4392), .B(n4393), .Z(n4390) );
  XNOR U8503 ( .A(y[3706]), .B(x[3706]), .Z(n4393) );
  XNOR U8504 ( .A(y[3707]), .B(x[3707]), .Z(n4392) );
  XNOR U8505 ( .A(n4384), .B(n4385), .Z(n4395) );
  XNOR U8506 ( .A(y[3702]), .B(x[3702]), .Z(n4385) );
  XNOR U8507 ( .A(n4386), .B(n4387), .Z(n4384) );
  XNOR U8508 ( .A(y[3703]), .B(x[3703]), .Z(n4387) );
  XNOR U8509 ( .A(y[3704]), .B(x[3704]), .Z(n4386) );
  NAND U8510 ( .A(n4451), .B(n4452), .Z(N29781) );
  NANDN U8511 ( .A(n4453), .B(n4454), .Z(n4452) );
  OR U8512 ( .A(n4455), .B(n4456), .Z(n4454) );
  NAND U8513 ( .A(n4455), .B(n4456), .Z(n4451) );
  XOR U8514 ( .A(n4455), .B(n4457), .Z(N29780) );
  XNOR U8515 ( .A(n4453), .B(n4456), .Z(n4457) );
  AND U8516 ( .A(n4458), .B(n4459), .Z(n4456) );
  NANDN U8517 ( .A(n4460), .B(n4461), .Z(n4459) );
  NANDN U8518 ( .A(n4462), .B(n4463), .Z(n4461) );
  NANDN U8519 ( .A(n4463), .B(n4462), .Z(n4458) );
  NAND U8520 ( .A(n4464), .B(n4465), .Z(n4453) );
  NANDN U8521 ( .A(n4466), .B(n4467), .Z(n4465) );
  OR U8522 ( .A(n4468), .B(n4469), .Z(n4467) );
  NAND U8523 ( .A(n4469), .B(n4468), .Z(n4464) );
  AND U8524 ( .A(n4470), .B(n4471), .Z(n4455) );
  NANDN U8525 ( .A(n4472), .B(n4473), .Z(n4471) );
  NANDN U8526 ( .A(n4474), .B(n4475), .Z(n4473) );
  NANDN U8527 ( .A(n4475), .B(n4474), .Z(n4470) );
  XOR U8528 ( .A(n4469), .B(n4476), .Z(N29779) );
  XOR U8529 ( .A(n4466), .B(n4468), .Z(n4476) );
  XNOR U8530 ( .A(n4462), .B(n4477), .Z(n4468) );
  XNOR U8531 ( .A(n4460), .B(n4463), .Z(n4477) );
  NAND U8532 ( .A(n4478), .B(n4479), .Z(n4463) );
  NAND U8533 ( .A(n4480), .B(n4481), .Z(n4479) );
  OR U8534 ( .A(n4482), .B(n4483), .Z(n4480) );
  NANDN U8535 ( .A(n4484), .B(n4482), .Z(n4478) );
  IV U8536 ( .A(n4483), .Z(n4484) );
  NAND U8537 ( .A(n4485), .B(n4486), .Z(n4460) );
  NAND U8538 ( .A(n4487), .B(n4488), .Z(n4486) );
  NANDN U8539 ( .A(n4489), .B(n4490), .Z(n4487) );
  NANDN U8540 ( .A(n4490), .B(n4489), .Z(n4485) );
  AND U8541 ( .A(n4491), .B(n4492), .Z(n4462) );
  NAND U8542 ( .A(n4493), .B(n4494), .Z(n4492) );
  OR U8543 ( .A(n4495), .B(n4496), .Z(n4493) );
  NANDN U8544 ( .A(n4497), .B(n4495), .Z(n4491) );
  NAND U8545 ( .A(n4498), .B(n4499), .Z(n4466) );
  NANDN U8546 ( .A(n4500), .B(n4501), .Z(n4499) );
  OR U8547 ( .A(n4502), .B(n4503), .Z(n4501) );
  NANDN U8548 ( .A(n4504), .B(n4502), .Z(n4498) );
  IV U8549 ( .A(n4503), .Z(n4504) );
  XNOR U8550 ( .A(n4474), .B(n4505), .Z(n4469) );
  XNOR U8551 ( .A(n4472), .B(n4475), .Z(n4505) );
  NAND U8552 ( .A(n4506), .B(n4507), .Z(n4475) );
  NAND U8553 ( .A(n4508), .B(n4509), .Z(n4507) );
  OR U8554 ( .A(n4510), .B(n4511), .Z(n4508) );
  NANDN U8555 ( .A(n4512), .B(n4510), .Z(n4506) );
  IV U8556 ( .A(n4511), .Z(n4512) );
  NAND U8557 ( .A(n4513), .B(n4514), .Z(n4472) );
  NAND U8558 ( .A(n4515), .B(n4516), .Z(n4514) );
  NANDN U8559 ( .A(n4517), .B(n4518), .Z(n4515) );
  NANDN U8560 ( .A(n4518), .B(n4517), .Z(n4513) );
  AND U8561 ( .A(n4519), .B(n4520), .Z(n4474) );
  NAND U8562 ( .A(n4521), .B(n4522), .Z(n4520) );
  OR U8563 ( .A(n4523), .B(n4524), .Z(n4521) );
  NANDN U8564 ( .A(n4525), .B(n4523), .Z(n4519) );
  XNOR U8565 ( .A(n4500), .B(n4526), .Z(N29778) );
  XOR U8566 ( .A(n4502), .B(n4503), .Z(n4526) );
  XNOR U8567 ( .A(n4516), .B(n4527), .Z(n4503) );
  XOR U8568 ( .A(n4517), .B(n4518), .Z(n4527) );
  XOR U8569 ( .A(n4523), .B(n4528), .Z(n4518) );
  XOR U8570 ( .A(n4522), .B(n4525), .Z(n4528) );
  IV U8571 ( .A(n4524), .Z(n4525) );
  NAND U8572 ( .A(n4529), .B(n4530), .Z(n4524) );
  OR U8573 ( .A(n4531), .B(n4532), .Z(n4530) );
  OR U8574 ( .A(n4533), .B(n4534), .Z(n4529) );
  NAND U8575 ( .A(n4535), .B(n4536), .Z(n4522) );
  OR U8576 ( .A(n4537), .B(n4538), .Z(n4536) );
  OR U8577 ( .A(n4539), .B(n4540), .Z(n4535) );
  NOR U8578 ( .A(n4541), .B(n4542), .Z(n4523) );
  ANDN U8579 ( .B(n4543), .A(n4544), .Z(n4517) );
  XNOR U8580 ( .A(n4510), .B(n4545), .Z(n4516) );
  XNOR U8581 ( .A(n4509), .B(n4511), .Z(n4545) );
  NAND U8582 ( .A(n4546), .B(n4547), .Z(n4511) );
  OR U8583 ( .A(n4548), .B(n4549), .Z(n4547) );
  OR U8584 ( .A(n4550), .B(n4551), .Z(n4546) );
  NAND U8585 ( .A(n4552), .B(n4553), .Z(n4509) );
  OR U8586 ( .A(n4554), .B(n4555), .Z(n4553) );
  OR U8587 ( .A(n4556), .B(n4557), .Z(n4552) );
  ANDN U8588 ( .B(n4558), .A(n4559), .Z(n4510) );
  IV U8589 ( .A(n4560), .Z(n4558) );
  ANDN U8590 ( .B(n4561), .A(n4562), .Z(n4502) );
  XOR U8591 ( .A(n4488), .B(n4563), .Z(n4500) );
  XOR U8592 ( .A(n4489), .B(n4490), .Z(n4563) );
  XOR U8593 ( .A(n4495), .B(n4564), .Z(n4490) );
  XOR U8594 ( .A(n4494), .B(n4497), .Z(n4564) );
  IV U8595 ( .A(n4496), .Z(n4497) );
  NAND U8596 ( .A(n4565), .B(n4566), .Z(n4496) );
  OR U8597 ( .A(n4567), .B(n4568), .Z(n4566) );
  OR U8598 ( .A(n4569), .B(n4570), .Z(n4565) );
  NAND U8599 ( .A(n4571), .B(n4572), .Z(n4494) );
  OR U8600 ( .A(n4573), .B(n4574), .Z(n4572) );
  OR U8601 ( .A(n4575), .B(n4576), .Z(n4571) );
  NOR U8602 ( .A(n4577), .B(n4578), .Z(n4495) );
  ANDN U8603 ( .B(n4579), .A(n4580), .Z(n4489) );
  IV U8604 ( .A(n4581), .Z(n4579) );
  XNOR U8605 ( .A(n4482), .B(n4582), .Z(n4488) );
  XNOR U8606 ( .A(n4481), .B(n4483), .Z(n4582) );
  NAND U8607 ( .A(n4583), .B(n4584), .Z(n4483) );
  OR U8608 ( .A(n4585), .B(n4586), .Z(n4584) );
  OR U8609 ( .A(n4587), .B(n4588), .Z(n4583) );
  NAND U8610 ( .A(n4589), .B(n4590), .Z(n4481) );
  OR U8611 ( .A(n4591), .B(n4592), .Z(n4590) );
  OR U8612 ( .A(n4593), .B(n4594), .Z(n4589) );
  ANDN U8613 ( .B(n4595), .A(n4596), .Z(n4482) );
  IV U8614 ( .A(n4597), .Z(n4595) );
  XNOR U8615 ( .A(n4562), .B(n4561), .Z(N29777) );
  XOR U8616 ( .A(n4581), .B(n4580), .Z(n4561) );
  XNOR U8617 ( .A(n4596), .B(n4597), .Z(n4580) );
  XNOR U8618 ( .A(n4591), .B(n4592), .Z(n4597) );
  XNOR U8619 ( .A(n4593), .B(n4594), .Z(n4592) );
  XNOR U8620 ( .A(y[3700]), .B(x[3700]), .Z(n4594) );
  XNOR U8621 ( .A(y[3701]), .B(x[3701]), .Z(n4593) );
  XNOR U8622 ( .A(y[3699]), .B(x[3699]), .Z(n4591) );
  XNOR U8623 ( .A(n4585), .B(n4586), .Z(n4596) );
  XNOR U8624 ( .A(y[3696]), .B(x[3696]), .Z(n4586) );
  XNOR U8625 ( .A(n4587), .B(n4588), .Z(n4585) );
  XNOR U8626 ( .A(y[3697]), .B(x[3697]), .Z(n4588) );
  XNOR U8627 ( .A(y[3698]), .B(x[3698]), .Z(n4587) );
  XNOR U8628 ( .A(n4578), .B(n4577), .Z(n4581) );
  XNOR U8629 ( .A(n4573), .B(n4574), .Z(n4577) );
  XNOR U8630 ( .A(y[3693]), .B(x[3693]), .Z(n4574) );
  XNOR U8631 ( .A(n4575), .B(n4576), .Z(n4573) );
  XNOR U8632 ( .A(y[3694]), .B(x[3694]), .Z(n4576) );
  XNOR U8633 ( .A(y[3695]), .B(x[3695]), .Z(n4575) );
  XNOR U8634 ( .A(n4567), .B(n4568), .Z(n4578) );
  XNOR U8635 ( .A(y[3690]), .B(x[3690]), .Z(n4568) );
  XNOR U8636 ( .A(n4569), .B(n4570), .Z(n4567) );
  XNOR U8637 ( .A(y[3691]), .B(x[3691]), .Z(n4570) );
  XNOR U8638 ( .A(y[3692]), .B(x[3692]), .Z(n4569) );
  XOR U8639 ( .A(n4543), .B(n4544), .Z(n4562) );
  XNOR U8640 ( .A(n4559), .B(n4560), .Z(n4544) );
  XNOR U8641 ( .A(n4554), .B(n4555), .Z(n4560) );
  XNOR U8642 ( .A(n4556), .B(n4557), .Z(n4555) );
  XNOR U8643 ( .A(y[3688]), .B(x[3688]), .Z(n4557) );
  XNOR U8644 ( .A(y[3689]), .B(x[3689]), .Z(n4556) );
  XNOR U8645 ( .A(y[3687]), .B(x[3687]), .Z(n4554) );
  XNOR U8646 ( .A(n4548), .B(n4549), .Z(n4559) );
  XNOR U8647 ( .A(y[3684]), .B(x[3684]), .Z(n4549) );
  XNOR U8648 ( .A(n4550), .B(n4551), .Z(n4548) );
  XNOR U8649 ( .A(y[3685]), .B(x[3685]), .Z(n4551) );
  XNOR U8650 ( .A(y[3686]), .B(x[3686]), .Z(n4550) );
  XOR U8651 ( .A(n4542), .B(n4541), .Z(n4543) );
  XNOR U8652 ( .A(n4537), .B(n4538), .Z(n4541) );
  XNOR U8653 ( .A(y[3681]), .B(x[3681]), .Z(n4538) );
  XNOR U8654 ( .A(n4539), .B(n4540), .Z(n4537) );
  XNOR U8655 ( .A(y[3682]), .B(x[3682]), .Z(n4540) );
  XNOR U8656 ( .A(y[3683]), .B(x[3683]), .Z(n4539) );
  XNOR U8657 ( .A(n4531), .B(n4532), .Z(n4542) );
  XNOR U8658 ( .A(y[3678]), .B(x[3678]), .Z(n4532) );
  XNOR U8659 ( .A(n4533), .B(n4534), .Z(n4531) );
  XNOR U8660 ( .A(y[3679]), .B(x[3679]), .Z(n4534) );
  XNOR U8661 ( .A(y[3680]), .B(x[3680]), .Z(n4533) );
  NAND U8662 ( .A(n4598), .B(n4599), .Z(N29769) );
  NANDN U8663 ( .A(n4600), .B(n4601), .Z(n4599) );
  OR U8664 ( .A(n4602), .B(n4603), .Z(n4601) );
  NAND U8665 ( .A(n4602), .B(n4603), .Z(n4598) );
  XOR U8666 ( .A(n4602), .B(n4604), .Z(N29768) );
  XNOR U8667 ( .A(n4600), .B(n4603), .Z(n4604) );
  AND U8668 ( .A(n4605), .B(n4606), .Z(n4603) );
  NANDN U8669 ( .A(n4607), .B(n4608), .Z(n4606) );
  NANDN U8670 ( .A(n4609), .B(n4610), .Z(n4608) );
  NANDN U8671 ( .A(n4610), .B(n4609), .Z(n4605) );
  NAND U8672 ( .A(n4611), .B(n4612), .Z(n4600) );
  NANDN U8673 ( .A(n4613), .B(n4614), .Z(n4612) );
  OR U8674 ( .A(n4615), .B(n4616), .Z(n4614) );
  NAND U8675 ( .A(n4616), .B(n4615), .Z(n4611) );
  AND U8676 ( .A(n4617), .B(n4618), .Z(n4602) );
  NANDN U8677 ( .A(n4619), .B(n4620), .Z(n4618) );
  NANDN U8678 ( .A(n4621), .B(n4622), .Z(n4620) );
  NANDN U8679 ( .A(n4622), .B(n4621), .Z(n4617) );
  XOR U8680 ( .A(n4616), .B(n4623), .Z(N29767) );
  XOR U8681 ( .A(n4613), .B(n4615), .Z(n4623) );
  XNOR U8682 ( .A(n4609), .B(n4624), .Z(n4615) );
  XNOR U8683 ( .A(n4607), .B(n4610), .Z(n4624) );
  NAND U8684 ( .A(n4625), .B(n4626), .Z(n4610) );
  NAND U8685 ( .A(n4627), .B(n4628), .Z(n4626) );
  OR U8686 ( .A(n4629), .B(n4630), .Z(n4627) );
  NANDN U8687 ( .A(n4631), .B(n4629), .Z(n4625) );
  IV U8688 ( .A(n4630), .Z(n4631) );
  NAND U8689 ( .A(n4632), .B(n4633), .Z(n4607) );
  NAND U8690 ( .A(n4634), .B(n4635), .Z(n4633) );
  NANDN U8691 ( .A(n4636), .B(n4637), .Z(n4634) );
  NANDN U8692 ( .A(n4637), .B(n4636), .Z(n4632) );
  AND U8693 ( .A(n4638), .B(n4639), .Z(n4609) );
  NAND U8694 ( .A(n4640), .B(n4641), .Z(n4639) );
  OR U8695 ( .A(n4642), .B(n4643), .Z(n4640) );
  NANDN U8696 ( .A(n4644), .B(n4642), .Z(n4638) );
  NAND U8697 ( .A(n4645), .B(n4646), .Z(n4613) );
  NANDN U8698 ( .A(n4647), .B(n4648), .Z(n4646) );
  OR U8699 ( .A(n4649), .B(n4650), .Z(n4648) );
  NANDN U8700 ( .A(n4651), .B(n4649), .Z(n4645) );
  IV U8701 ( .A(n4650), .Z(n4651) );
  XNOR U8702 ( .A(n4621), .B(n4652), .Z(n4616) );
  XNOR U8703 ( .A(n4619), .B(n4622), .Z(n4652) );
  NAND U8704 ( .A(n4653), .B(n4654), .Z(n4622) );
  NAND U8705 ( .A(n4655), .B(n4656), .Z(n4654) );
  OR U8706 ( .A(n4657), .B(n4658), .Z(n4655) );
  NANDN U8707 ( .A(n4659), .B(n4657), .Z(n4653) );
  IV U8708 ( .A(n4658), .Z(n4659) );
  NAND U8709 ( .A(n4660), .B(n4661), .Z(n4619) );
  NAND U8710 ( .A(n4662), .B(n4663), .Z(n4661) );
  NANDN U8711 ( .A(n4664), .B(n4665), .Z(n4662) );
  NANDN U8712 ( .A(n4665), .B(n4664), .Z(n4660) );
  AND U8713 ( .A(n4666), .B(n4667), .Z(n4621) );
  NAND U8714 ( .A(n4668), .B(n4669), .Z(n4667) );
  OR U8715 ( .A(n4670), .B(n4671), .Z(n4668) );
  NANDN U8716 ( .A(n4672), .B(n4670), .Z(n4666) );
  XNOR U8717 ( .A(n4647), .B(n4673), .Z(N29766) );
  XOR U8718 ( .A(n4649), .B(n4650), .Z(n4673) );
  XNOR U8719 ( .A(n4663), .B(n4674), .Z(n4650) );
  XOR U8720 ( .A(n4664), .B(n4665), .Z(n4674) );
  XOR U8721 ( .A(n4670), .B(n4675), .Z(n4665) );
  XOR U8722 ( .A(n4669), .B(n4672), .Z(n4675) );
  IV U8723 ( .A(n4671), .Z(n4672) );
  NAND U8724 ( .A(n4676), .B(n4677), .Z(n4671) );
  OR U8725 ( .A(n4678), .B(n4679), .Z(n4677) );
  OR U8726 ( .A(n4680), .B(n4681), .Z(n4676) );
  NAND U8727 ( .A(n4682), .B(n4683), .Z(n4669) );
  OR U8728 ( .A(n4684), .B(n4685), .Z(n4683) );
  OR U8729 ( .A(n4686), .B(n4687), .Z(n4682) );
  NOR U8730 ( .A(n4688), .B(n4689), .Z(n4670) );
  ANDN U8731 ( .B(n4690), .A(n4691), .Z(n4664) );
  XNOR U8732 ( .A(n4657), .B(n4692), .Z(n4663) );
  XNOR U8733 ( .A(n4656), .B(n4658), .Z(n4692) );
  NAND U8734 ( .A(n4693), .B(n4694), .Z(n4658) );
  OR U8735 ( .A(n4695), .B(n4696), .Z(n4694) );
  OR U8736 ( .A(n4697), .B(n4698), .Z(n4693) );
  NAND U8737 ( .A(n4699), .B(n4700), .Z(n4656) );
  OR U8738 ( .A(n4701), .B(n4702), .Z(n4700) );
  OR U8739 ( .A(n4703), .B(n4704), .Z(n4699) );
  ANDN U8740 ( .B(n4705), .A(n4706), .Z(n4657) );
  IV U8741 ( .A(n4707), .Z(n4705) );
  ANDN U8742 ( .B(n4708), .A(n4709), .Z(n4649) );
  XOR U8743 ( .A(n4635), .B(n4710), .Z(n4647) );
  XOR U8744 ( .A(n4636), .B(n4637), .Z(n4710) );
  XOR U8745 ( .A(n4642), .B(n4711), .Z(n4637) );
  XOR U8746 ( .A(n4641), .B(n4644), .Z(n4711) );
  IV U8747 ( .A(n4643), .Z(n4644) );
  NAND U8748 ( .A(n4712), .B(n4713), .Z(n4643) );
  OR U8749 ( .A(n4714), .B(n4715), .Z(n4713) );
  OR U8750 ( .A(n4716), .B(n4717), .Z(n4712) );
  NAND U8751 ( .A(n4718), .B(n4719), .Z(n4641) );
  OR U8752 ( .A(n4720), .B(n4721), .Z(n4719) );
  OR U8753 ( .A(n4722), .B(n4723), .Z(n4718) );
  NOR U8754 ( .A(n4724), .B(n4725), .Z(n4642) );
  ANDN U8755 ( .B(n4726), .A(n4727), .Z(n4636) );
  IV U8756 ( .A(n4728), .Z(n4726) );
  XNOR U8757 ( .A(n4629), .B(n4729), .Z(n4635) );
  XNOR U8758 ( .A(n4628), .B(n4630), .Z(n4729) );
  NAND U8759 ( .A(n4730), .B(n4731), .Z(n4630) );
  OR U8760 ( .A(n4732), .B(n4733), .Z(n4731) );
  OR U8761 ( .A(n4734), .B(n4735), .Z(n4730) );
  NAND U8762 ( .A(n4736), .B(n4737), .Z(n4628) );
  OR U8763 ( .A(n4738), .B(n4739), .Z(n4737) );
  OR U8764 ( .A(n4740), .B(n4741), .Z(n4736) );
  ANDN U8765 ( .B(n4742), .A(n4743), .Z(n4629) );
  IV U8766 ( .A(n4744), .Z(n4742) );
  XNOR U8767 ( .A(n4709), .B(n4708), .Z(N29765) );
  XOR U8768 ( .A(n4728), .B(n4727), .Z(n4708) );
  XNOR U8769 ( .A(n4743), .B(n4744), .Z(n4727) );
  XNOR U8770 ( .A(n4738), .B(n4739), .Z(n4744) );
  XNOR U8771 ( .A(n4740), .B(n4741), .Z(n4739) );
  XNOR U8772 ( .A(y[3676]), .B(x[3676]), .Z(n4741) );
  XNOR U8773 ( .A(y[3677]), .B(x[3677]), .Z(n4740) );
  XNOR U8774 ( .A(y[3675]), .B(x[3675]), .Z(n4738) );
  XNOR U8775 ( .A(n4732), .B(n4733), .Z(n4743) );
  XNOR U8776 ( .A(y[3672]), .B(x[3672]), .Z(n4733) );
  XNOR U8777 ( .A(n4734), .B(n4735), .Z(n4732) );
  XNOR U8778 ( .A(y[3673]), .B(x[3673]), .Z(n4735) );
  XNOR U8779 ( .A(y[3674]), .B(x[3674]), .Z(n4734) );
  XNOR U8780 ( .A(n4725), .B(n4724), .Z(n4728) );
  XNOR U8781 ( .A(n4720), .B(n4721), .Z(n4724) );
  XNOR U8782 ( .A(y[3669]), .B(x[3669]), .Z(n4721) );
  XNOR U8783 ( .A(n4722), .B(n4723), .Z(n4720) );
  XNOR U8784 ( .A(y[3670]), .B(x[3670]), .Z(n4723) );
  XNOR U8785 ( .A(y[3671]), .B(x[3671]), .Z(n4722) );
  XNOR U8786 ( .A(n4714), .B(n4715), .Z(n4725) );
  XNOR U8787 ( .A(y[3666]), .B(x[3666]), .Z(n4715) );
  XNOR U8788 ( .A(n4716), .B(n4717), .Z(n4714) );
  XNOR U8789 ( .A(y[3667]), .B(x[3667]), .Z(n4717) );
  XNOR U8790 ( .A(y[3668]), .B(x[3668]), .Z(n4716) );
  XOR U8791 ( .A(n4690), .B(n4691), .Z(n4709) );
  XNOR U8792 ( .A(n4706), .B(n4707), .Z(n4691) );
  XNOR U8793 ( .A(n4701), .B(n4702), .Z(n4707) );
  XNOR U8794 ( .A(n4703), .B(n4704), .Z(n4702) );
  XNOR U8795 ( .A(y[3664]), .B(x[3664]), .Z(n4704) );
  XNOR U8796 ( .A(y[3665]), .B(x[3665]), .Z(n4703) );
  XNOR U8797 ( .A(y[3663]), .B(x[3663]), .Z(n4701) );
  XNOR U8798 ( .A(n4695), .B(n4696), .Z(n4706) );
  XNOR U8799 ( .A(y[3660]), .B(x[3660]), .Z(n4696) );
  XNOR U8800 ( .A(n4697), .B(n4698), .Z(n4695) );
  XNOR U8801 ( .A(y[3661]), .B(x[3661]), .Z(n4698) );
  XNOR U8802 ( .A(y[3662]), .B(x[3662]), .Z(n4697) );
  XOR U8803 ( .A(n4689), .B(n4688), .Z(n4690) );
  XNOR U8804 ( .A(n4684), .B(n4685), .Z(n4688) );
  XNOR U8805 ( .A(y[3657]), .B(x[3657]), .Z(n4685) );
  XNOR U8806 ( .A(n4686), .B(n4687), .Z(n4684) );
  XNOR U8807 ( .A(y[3658]), .B(x[3658]), .Z(n4687) );
  XNOR U8808 ( .A(y[3659]), .B(x[3659]), .Z(n4686) );
  XNOR U8809 ( .A(n4678), .B(n4679), .Z(n4689) );
  XNOR U8810 ( .A(y[3654]), .B(x[3654]), .Z(n4679) );
  XNOR U8811 ( .A(n4680), .B(n4681), .Z(n4678) );
  XNOR U8812 ( .A(y[3655]), .B(x[3655]), .Z(n4681) );
  XNOR U8813 ( .A(y[3656]), .B(x[3656]), .Z(n4680) );
  NAND U8814 ( .A(n4745), .B(n4746), .Z(N29757) );
  NANDN U8815 ( .A(n4747), .B(n4748), .Z(n4746) );
  OR U8816 ( .A(n4749), .B(n4750), .Z(n4748) );
  NAND U8817 ( .A(n4749), .B(n4750), .Z(n4745) );
  XOR U8818 ( .A(n4749), .B(n4751), .Z(N29756) );
  XNOR U8819 ( .A(n4747), .B(n4750), .Z(n4751) );
  AND U8820 ( .A(n4752), .B(n4753), .Z(n4750) );
  NANDN U8821 ( .A(n4754), .B(n4755), .Z(n4753) );
  NANDN U8822 ( .A(n4756), .B(n4757), .Z(n4755) );
  NANDN U8823 ( .A(n4757), .B(n4756), .Z(n4752) );
  NAND U8824 ( .A(n4758), .B(n4759), .Z(n4747) );
  NANDN U8825 ( .A(n4760), .B(n4761), .Z(n4759) );
  OR U8826 ( .A(n4762), .B(n4763), .Z(n4761) );
  NAND U8827 ( .A(n4763), .B(n4762), .Z(n4758) );
  AND U8828 ( .A(n4764), .B(n4765), .Z(n4749) );
  NANDN U8829 ( .A(n4766), .B(n4767), .Z(n4765) );
  NANDN U8830 ( .A(n4768), .B(n4769), .Z(n4767) );
  NANDN U8831 ( .A(n4769), .B(n4768), .Z(n4764) );
  XOR U8832 ( .A(n4763), .B(n4770), .Z(N29755) );
  XOR U8833 ( .A(n4760), .B(n4762), .Z(n4770) );
  XNOR U8834 ( .A(n4756), .B(n4771), .Z(n4762) );
  XNOR U8835 ( .A(n4754), .B(n4757), .Z(n4771) );
  NAND U8836 ( .A(n4772), .B(n4773), .Z(n4757) );
  NAND U8837 ( .A(n4774), .B(n4775), .Z(n4773) );
  OR U8838 ( .A(n4776), .B(n4777), .Z(n4774) );
  NANDN U8839 ( .A(n4778), .B(n4776), .Z(n4772) );
  IV U8840 ( .A(n4777), .Z(n4778) );
  NAND U8841 ( .A(n4779), .B(n4780), .Z(n4754) );
  NAND U8842 ( .A(n4781), .B(n4782), .Z(n4780) );
  NANDN U8843 ( .A(n4783), .B(n4784), .Z(n4781) );
  NANDN U8844 ( .A(n4784), .B(n4783), .Z(n4779) );
  AND U8845 ( .A(n4785), .B(n4786), .Z(n4756) );
  NAND U8846 ( .A(n4787), .B(n4788), .Z(n4786) );
  OR U8847 ( .A(n4789), .B(n4790), .Z(n4787) );
  NANDN U8848 ( .A(n4791), .B(n4789), .Z(n4785) );
  NAND U8849 ( .A(n4792), .B(n4793), .Z(n4760) );
  NANDN U8850 ( .A(n4794), .B(n4795), .Z(n4793) );
  OR U8851 ( .A(n4796), .B(n4797), .Z(n4795) );
  NANDN U8852 ( .A(n4798), .B(n4796), .Z(n4792) );
  IV U8853 ( .A(n4797), .Z(n4798) );
  XNOR U8854 ( .A(n4768), .B(n4799), .Z(n4763) );
  XNOR U8855 ( .A(n4766), .B(n4769), .Z(n4799) );
  NAND U8856 ( .A(n4800), .B(n4801), .Z(n4769) );
  NAND U8857 ( .A(n4802), .B(n4803), .Z(n4801) );
  OR U8858 ( .A(n4804), .B(n4805), .Z(n4802) );
  NANDN U8859 ( .A(n4806), .B(n4804), .Z(n4800) );
  IV U8860 ( .A(n4805), .Z(n4806) );
  NAND U8861 ( .A(n4807), .B(n4808), .Z(n4766) );
  NAND U8862 ( .A(n4809), .B(n4810), .Z(n4808) );
  NANDN U8863 ( .A(n4811), .B(n4812), .Z(n4809) );
  NANDN U8864 ( .A(n4812), .B(n4811), .Z(n4807) );
  AND U8865 ( .A(n4813), .B(n4814), .Z(n4768) );
  NAND U8866 ( .A(n4815), .B(n4816), .Z(n4814) );
  OR U8867 ( .A(n4817), .B(n4818), .Z(n4815) );
  NANDN U8868 ( .A(n4819), .B(n4817), .Z(n4813) );
  XNOR U8869 ( .A(n4794), .B(n4820), .Z(N29754) );
  XOR U8870 ( .A(n4796), .B(n4797), .Z(n4820) );
  XNOR U8871 ( .A(n4810), .B(n4821), .Z(n4797) );
  XOR U8872 ( .A(n4811), .B(n4812), .Z(n4821) );
  XOR U8873 ( .A(n4817), .B(n4822), .Z(n4812) );
  XOR U8874 ( .A(n4816), .B(n4819), .Z(n4822) );
  IV U8875 ( .A(n4818), .Z(n4819) );
  NAND U8876 ( .A(n4823), .B(n4824), .Z(n4818) );
  OR U8877 ( .A(n4825), .B(n4826), .Z(n4824) );
  OR U8878 ( .A(n4827), .B(n4828), .Z(n4823) );
  NAND U8879 ( .A(n4829), .B(n4830), .Z(n4816) );
  OR U8880 ( .A(n4831), .B(n4832), .Z(n4830) );
  OR U8881 ( .A(n4833), .B(n4834), .Z(n4829) );
  NOR U8882 ( .A(n4835), .B(n4836), .Z(n4817) );
  ANDN U8883 ( .B(n4837), .A(n4838), .Z(n4811) );
  XNOR U8884 ( .A(n4804), .B(n4839), .Z(n4810) );
  XNOR U8885 ( .A(n4803), .B(n4805), .Z(n4839) );
  NAND U8886 ( .A(n4840), .B(n4841), .Z(n4805) );
  OR U8887 ( .A(n4842), .B(n4843), .Z(n4841) );
  OR U8888 ( .A(n4844), .B(n4845), .Z(n4840) );
  NAND U8889 ( .A(n4846), .B(n4847), .Z(n4803) );
  OR U8890 ( .A(n4848), .B(n4849), .Z(n4847) );
  OR U8891 ( .A(n4850), .B(n4851), .Z(n4846) );
  ANDN U8892 ( .B(n4852), .A(n4853), .Z(n4804) );
  IV U8893 ( .A(n4854), .Z(n4852) );
  ANDN U8894 ( .B(n4855), .A(n4856), .Z(n4796) );
  XOR U8895 ( .A(n4782), .B(n4857), .Z(n4794) );
  XOR U8896 ( .A(n4783), .B(n4784), .Z(n4857) );
  XOR U8897 ( .A(n4789), .B(n4858), .Z(n4784) );
  XOR U8898 ( .A(n4788), .B(n4791), .Z(n4858) );
  IV U8899 ( .A(n4790), .Z(n4791) );
  NAND U8900 ( .A(n4859), .B(n4860), .Z(n4790) );
  OR U8901 ( .A(n4861), .B(n4862), .Z(n4860) );
  OR U8902 ( .A(n4863), .B(n4864), .Z(n4859) );
  NAND U8903 ( .A(n4865), .B(n4866), .Z(n4788) );
  OR U8904 ( .A(n4867), .B(n4868), .Z(n4866) );
  OR U8905 ( .A(n4869), .B(n4870), .Z(n4865) );
  NOR U8906 ( .A(n4871), .B(n4872), .Z(n4789) );
  ANDN U8907 ( .B(n4873), .A(n4874), .Z(n4783) );
  IV U8908 ( .A(n4875), .Z(n4873) );
  XNOR U8909 ( .A(n4776), .B(n4876), .Z(n4782) );
  XNOR U8910 ( .A(n4775), .B(n4777), .Z(n4876) );
  NAND U8911 ( .A(n4877), .B(n4878), .Z(n4777) );
  OR U8912 ( .A(n4879), .B(n4880), .Z(n4878) );
  OR U8913 ( .A(n4881), .B(n4882), .Z(n4877) );
  NAND U8914 ( .A(n4883), .B(n4884), .Z(n4775) );
  OR U8915 ( .A(n4885), .B(n4886), .Z(n4884) );
  OR U8916 ( .A(n4887), .B(n4888), .Z(n4883) );
  ANDN U8917 ( .B(n4889), .A(n4890), .Z(n4776) );
  IV U8918 ( .A(n4891), .Z(n4889) );
  XNOR U8919 ( .A(n4856), .B(n4855), .Z(N29753) );
  XOR U8920 ( .A(n4875), .B(n4874), .Z(n4855) );
  XNOR U8921 ( .A(n4890), .B(n4891), .Z(n4874) );
  XNOR U8922 ( .A(n4885), .B(n4886), .Z(n4891) );
  XNOR U8923 ( .A(n4887), .B(n4888), .Z(n4886) );
  XNOR U8924 ( .A(y[3652]), .B(x[3652]), .Z(n4888) );
  XNOR U8925 ( .A(y[3653]), .B(x[3653]), .Z(n4887) );
  XNOR U8926 ( .A(y[3651]), .B(x[3651]), .Z(n4885) );
  XNOR U8927 ( .A(n4879), .B(n4880), .Z(n4890) );
  XNOR U8928 ( .A(y[3648]), .B(x[3648]), .Z(n4880) );
  XNOR U8929 ( .A(n4881), .B(n4882), .Z(n4879) );
  XNOR U8930 ( .A(y[3649]), .B(x[3649]), .Z(n4882) );
  XNOR U8931 ( .A(y[3650]), .B(x[3650]), .Z(n4881) );
  XNOR U8932 ( .A(n4872), .B(n4871), .Z(n4875) );
  XNOR U8933 ( .A(n4867), .B(n4868), .Z(n4871) );
  XNOR U8934 ( .A(y[3645]), .B(x[3645]), .Z(n4868) );
  XNOR U8935 ( .A(n4869), .B(n4870), .Z(n4867) );
  XNOR U8936 ( .A(y[3646]), .B(x[3646]), .Z(n4870) );
  XNOR U8937 ( .A(y[3647]), .B(x[3647]), .Z(n4869) );
  XNOR U8938 ( .A(n4861), .B(n4862), .Z(n4872) );
  XNOR U8939 ( .A(y[3642]), .B(x[3642]), .Z(n4862) );
  XNOR U8940 ( .A(n4863), .B(n4864), .Z(n4861) );
  XNOR U8941 ( .A(y[3643]), .B(x[3643]), .Z(n4864) );
  XNOR U8942 ( .A(y[3644]), .B(x[3644]), .Z(n4863) );
  XOR U8943 ( .A(n4837), .B(n4838), .Z(n4856) );
  XNOR U8944 ( .A(n4853), .B(n4854), .Z(n4838) );
  XNOR U8945 ( .A(n4848), .B(n4849), .Z(n4854) );
  XNOR U8946 ( .A(n4850), .B(n4851), .Z(n4849) );
  XNOR U8947 ( .A(y[3640]), .B(x[3640]), .Z(n4851) );
  XNOR U8948 ( .A(y[3641]), .B(x[3641]), .Z(n4850) );
  XNOR U8949 ( .A(y[3639]), .B(x[3639]), .Z(n4848) );
  XNOR U8950 ( .A(n4842), .B(n4843), .Z(n4853) );
  XNOR U8951 ( .A(y[3636]), .B(x[3636]), .Z(n4843) );
  XNOR U8952 ( .A(n4844), .B(n4845), .Z(n4842) );
  XNOR U8953 ( .A(y[3637]), .B(x[3637]), .Z(n4845) );
  XNOR U8954 ( .A(y[3638]), .B(x[3638]), .Z(n4844) );
  XOR U8955 ( .A(n4836), .B(n4835), .Z(n4837) );
  XNOR U8956 ( .A(n4831), .B(n4832), .Z(n4835) );
  XNOR U8957 ( .A(y[3633]), .B(x[3633]), .Z(n4832) );
  XNOR U8958 ( .A(n4833), .B(n4834), .Z(n4831) );
  XNOR U8959 ( .A(y[3634]), .B(x[3634]), .Z(n4834) );
  XNOR U8960 ( .A(y[3635]), .B(x[3635]), .Z(n4833) );
  XNOR U8961 ( .A(n4825), .B(n4826), .Z(n4836) );
  XNOR U8962 ( .A(y[3630]), .B(x[3630]), .Z(n4826) );
  XNOR U8963 ( .A(n4827), .B(n4828), .Z(n4825) );
  XNOR U8964 ( .A(y[3631]), .B(x[3631]), .Z(n4828) );
  XNOR U8965 ( .A(y[3632]), .B(x[3632]), .Z(n4827) );
  NAND U8966 ( .A(n4892), .B(n4893), .Z(N29745) );
  NANDN U8967 ( .A(n4894), .B(n4895), .Z(n4893) );
  OR U8968 ( .A(n4896), .B(n4897), .Z(n4895) );
  NAND U8969 ( .A(n4896), .B(n4897), .Z(n4892) );
  XOR U8970 ( .A(n4896), .B(n4898), .Z(N29744) );
  XNOR U8971 ( .A(n4894), .B(n4897), .Z(n4898) );
  AND U8972 ( .A(n4899), .B(n4900), .Z(n4897) );
  NANDN U8973 ( .A(n4901), .B(n4902), .Z(n4900) );
  NANDN U8974 ( .A(n4903), .B(n4904), .Z(n4902) );
  NANDN U8975 ( .A(n4904), .B(n4903), .Z(n4899) );
  NAND U8976 ( .A(n4905), .B(n4906), .Z(n4894) );
  NANDN U8977 ( .A(n4907), .B(n4908), .Z(n4906) );
  OR U8978 ( .A(n4909), .B(n4910), .Z(n4908) );
  NAND U8979 ( .A(n4910), .B(n4909), .Z(n4905) );
  AND U8980 ( .A(n4911), .B(n4912), .Z(n4896) );
  NANDN U8981 ( .A(n4913), .B(n4914), .Z(n4912) );
  NANDN U8982 ( .A(n4915), .B(n4916), .Z(n4914) );
  NANDN U8983 ( .A(n4916), .B(n4915), .Z(n4911) );
  XOR U8984 ( .A(n4910), .B(n4917), .Z(N29743) );
  XOR U8985 ( .A(n4907), .B(n4909), .Z(n4917) );
  XNOR U8986 ( .A(n4903), .B(n4918), .Z(n4909) );
  XNOR U8987 ( .A(n4901), .B(n4904), .Z(n4918) );
  NAND U8988 ( .A(n4919), .B(n4920), .Z(n4904) );
  NAND U8989 ( .A(n4921), .B(n4922), .Z(n4920) );
  OR U8990 ( .A(n4923), .B(n4924), .Z(n4921) );
  NANDN U8991 ( .A(n4925), .B(n4923), .Z(n4919) );
  IV U8992 ( .A(n4924), .Z(n4925) );
  NAND U8993 ( .A(n4926), .B(n4927), .Z(n4901) );
  NAND U8994 ( .A(n4928), .B(n4929), .Z(n4927) );
  NANDN U8995 ( .A(n4930), .B(n4931), .Z(n4928) );
  NANDN U8996 ( .A(n4931), .B(n4930), .Z(n4926) );
  AND U8997 ( .A(n4932), .B(n4933), .Z(n4903) );
  NAND U8998 ( .A(n4934), .B(n4935), .Z(n4933) );
  OR U8999 ( .A(n4936), .B(n4937), .Z(n4934) );
  NANDN U9000 ( .A(n4938), .B(n4936), .Z(n4932) );
  NAND U9001 ( .A(n4939), .B(n4940), .Z(n4907) );
  NANDN U9002 ( .A(n4941), .B(n4942), .Z(n4940) );
  OR U9003 ( .A(n4943), .B(n4944), .Z(n4942) );
  NANDN U9004 ( .A(n4945), .B(n4943), .Z(n4939) );
  IV U9005 ( .A(n4944), .Z(n4945) );
  XNOR U9006 ( .A(n4915), .B(n4946), .Z(n4910) );
  XNOR U9007 ( .A(n4913), .B(n4916), .Z(n4946) );
  NAND U9008 ( .A(n4947), .B(n4948), .Z(n4916) );
  NAND U9009 ( .A(n4949), .B(n4950), .Z(n4948) );
  OR U9010 ( .A(n4951), .B(n4952), .Z(n4949) );
  NANDN U9011 ( .A(n4953), .B(n4951), .Z(n4947) );
  IV U9012 ( .A(n4952), .Z(n4953) );
  NAND U9013 ( .A(n4954), .B(n4955), .Z(n4913) );
  NAND U9014 ( .A(n4956), .B(n4957), .Z(n4955) );
  NANDN U9015 ( .A(n4958), .B(n4959), .Z(n4956) );
  NANDN U9016 ( .A(n4959), .B(n4958), .Z(n4954) );
  AND U9017 ( .A(n4960), .B(n4961), .Z(n4915) );
  NAND U9018 ( .A(n4962), .B(n4963), .Z(n4961) );
  OR U9019 ( .A(n4964), .B(n4965), .Z(n4962) );
  NANDN U9020 ( .A(n4966), .B(n4964), .Z(n4960) );
  XNOR U9021 ( .A(n4941), .B(n4967), .Z(N29742) );
  XOR U9022 ( .A(n4943), .B(n4944), .Z(n4967) );
  XNOR U9023 ( .A(n4957), .B(n4968), .Z(n4944) );
  XOR U9024 ( .A(n4958), .B(n4959), .Z(n4968) );
  XOR U9025 ( .A(n4964), .B(n4969), .Z(n4959) );
  XOR U9026 ( .A(n4963), .B(n4966), .Z(n4969) );
  IV U9027 ( .A(n4965), .Z(n4966) );
  NAND U9028 ( .A(n4970), .B(n4971), .Z(n4965) );
  OR U9029 ( .A(n4972), .B(n4973), .Z(n4971) );
  OR U9030 ( .A(n4974), .B(n4975), .Z(n4970) );
  NAND U9031 ( .A(n4976), .B(n4977), .Z(n4963) );
  OR U9032 ( .A(n4978), .B(n4979), .Z(n4977) );
  OR U9033 ( .A(n4980), .B(n4981), .Z(n4976) );
  NOR U9034 ( .A(n4982), .B(n4983), .Z(n4964) );
  ANDN U9035 ( .B(n4984), .A(n4985), .Z(n4958) );
  XNOR U9036 ( .A(n4951), .B(n4986), .Z(n4957) );
  XNOR U9037 ( .A(n4950), .B(n4952), .Z(n4986) );
  NAND U9038 ( .A(n4987), .B(n4988), .Z(n4952) );
  OR U9039 ( .A(n4989), .B(n4990), .Z(n4988) );
  OR U9040 ( .A(n4991), .B(n4992), .Z(n4987) );
  NAND U9041 ( .A(n4993), .B(n4994), .Z(n4950) );
  OR U9042 ( .A(n4995), .B(n4996), .Z(n4994) );
  OR U9043 ( .A(n4997), .B(n4998), .Z(n4993) );
  ANDN U9044 ( .B(n4999), .A(n5000), .Z(n4951) );
  IV U9045 ( .A(n5001), .Z(n4999) );
  ANDN U9046 ( .B(n5002), .A(n5003), .Z(n4943) );
  XOR U9047 ( .A(n4929), .B(n5004), .Z(n4941) );
  XOR U9048 ( .A(n4930), .B(n4931), .Z(n5004) );
  XOR U9049 ( .A(n4936), .B(n5005), .Z(n4931) );
  XOR U9050 ( .A(n4935), .B(n4938), .Z(n5005) );
  IV U9051 ( .A(n4937), .Z(n4938) );
  NAND U9052 ( .A(n5006), .B(n5007), .Z(n4937) );
  OR U9053 ( .A(n5008), .B(n5009), .Z(n5007) );
  OR U9054 ( .A(n5010), .B(n5011), .Z(n5006) );
  NAND U9055 ( .A(n5012), .B(n5013), .Z(n4935) );
  OR U9056 ( .A(n5014), .B(n5015), .Z(n5013) );
  OR U9057 ( .A(n5016), .B(n5017), .Z(n5012) );
  NOR U9058 ( .A(n5018), .B(n5019), .Z(n4936) );
  ANDN U9059 ( .B(n5020), .A(n5021), .Z(n4930) );
  IV U9060 ( .A(n5022), .Z(n5020) );
  XNOR U9061 ( .A(n4923), .B(n5023), .Z(n4929) );
  XNOR U9062 ( .A(n4922), .B(n4924), .Z(n5023) );
  NAND U9063 ( .A(n5024), .B(n5025), .Z(n4924) );
  OR U9064 ( .A(n5026), .B(n5027), .Z(n5025) );
  OR U9065 ( .A(n5028), .B(n5029), .Z(n5024) );
  NAND U9066 ( .A(n5030), .B(n5031), .Z(n4922) );
  OR U9067 ( .A(n5032), .B(n5033), .Z(n5031) );
  OR U9068 ( .A(n5034), .B(n5035), .Z(n5030) );
  ANDN U9069 ( .B(n5036), .A(n5037), .Z(n4923) );
  IV U9070 ( .A(n5038), .Z(n5036) );
  XNOR U9071 ( .A(n5003), .B(n5002), .Z(N29741) );
  XOR U9072 ( .A(n5022), .B(n5021), .Z(n5002) );
  XNOR U9073 ( .A(n5037), .B(n5038), .Z(n5021) );
  XNOR U9074 ( .A(n5032), .B(n5033), .Z(n5038) );
  XNOR U9075 ( .A(n5034), .B(n5035), .Z(n5033) );
  XNOR U9076 ( .A(y[3628]), .B(x[3628]), .Z(n5035) );
  XNOR U9077 ( .A(y[3629]), .B(x[3629]), .Z(n5034) );
  XNOR U9078 ( .A(y[3627]), .B(x[3627]), .Z(n5032) );
  XNOR U9079 ( .A(n5026), .B(n5027), .Z(n5037) );
  XNOR U9080 ( .A(y[3624]), .B(x[3624]), .Z(n5027) );
  XNOR U9081 ( .A(n5028), .B(n5029), .Z(n5026) );
  XNOR U9082 ( .A(y[3625]), .B(x[3625]), .Z(n5029) );
  XNOR U9083 ( .A(y[3626]), .B(x[3626]), .Z(n5028) );
  XNOR U9084 ( .A(n5019), .B(n5018), .Z(n5022) );
  XNOR U9085 ( .A(n5014), .B(n5015), .Z(n5018) );
  XNOR U9086 ( .A(y[3621]), .B(x[3621]), .Z(n5015) );
  XNOR U9087 ( .A(n5016), .B(n5017), .Z(n5014) );
  XNOR U9088 ( .A(y[3622]), .B(x[3622]), .Z(n5017) );
  XNOR U9089 ( .A(y[3623]), .B(x[3623]), .Z(n5016) );
  XNOR U9090 ( .A(n5008), .B(n5009), .Z(n5019) );
  XNOR U9091 ( .A(y[3618]), .B(x[3618]), .Z(n5009) );
  XNOR U9092 ( .A(n5010), .B(n5011), .Z(n5008) );
  XNOR U9093 ( .A(y[3619]), .B(x[3619]), .Z(n5011) );
  XNOR U9094 ( .A(y[3620]), .B(x[3620]), .Z(n5010) );
  XOR U9095 ( .A(n4984), .B(n4985), .Z(n5003) );
  XNOR U9096 ( .A(n5000), .B(n5001), .Z(n4985) );
  XNOR U9097 ( .A(n4995), .B(n4996), .Z(n5001) );
  XNOR U9098 ( .A(n4997), .B(n4998), .Z(n4996) );
  XNOR U9099 ( .A(y[3616]), .B(x[3616]), .Z(n4998) );
  XNOR U9100 ( .A(y[3617]), .B(x[3617]), .Z(n4997) );
  XNOR U9101 ( .A(y[3615]), .B(x[3615]), .Z(n4995) );
  XNOR U9102 ( .A(n4989), .B(n4990), .Z(n5000) );
  XNOR U9103 ( .A(y[3612]), .B(x[3612]), .Z(n4990) );
  XNOR U9104 ( .A(n4991), .B(n4992), .Z(n4989) );
  XNOR U9105 ( .A(y[3613]), .B(x[3613]), .Z(n4992) );
  XNOR U9106 ( .A(y[3614]), .B(x[3614]), .Z(n4991) );
  XOR U9107 ( .A(n4983), .B(n4982), .Z(n4984) );
  XNOR U9108 ( .A(n4978), .B(n4979), .Z(n4982) );
  XNOR U9109 ( .A(y[3609]), .B(x[3609]), .Z(n4979) );
  XNOR U9110 ( .A(n4980), .B(n4981), .Z(n4978) );
  XNOR U9111 ( .A(y[3610]), .B(x[3610]), .Z(n4981) );
  XNOR U9112 ( .A(y[3611]), .B(x[3611]), .Z(n4980) );
  XNOR U9113 ( .A(n4972), .B(n4973), .Z(n4983) );
  XNOR U9114 ( .A(y[3606]), .B(x[3606]), .Z(n4973) );
  XNOR U9115 ( .A(n4974), .B(n4975), .Z(n4972) );
  XNOR U9116 ( .A(y[3607]), .B(x[3607]), .Z(n4975) );
  XNOR U9117 ( .A(y[3608]), .B(x[3608]), .Z(n4974) );
  NAND U9118 ( .A(n5039), .B(n5040), .Z(N29733) );
  NANDN U9119 ( .A(n5041), .B(n5042), .Z(n5040) );
  OR U9120 ( .A(n5043), .B(n5044), .Z(n5042) );
  NAND U9121 ( .A(n5043), .B(n5044), .Z(n5039) );
  XOR U9122 ( .A(n5043), .B(n5045), .Z(N29732) );
  XNOR U9123 ( .A(n5041), .B(n5044), .Z(n5045) );
  AND U9124 ( .A(n5046), .B(n5047), .Z(n5044) );
  NANDN U9125 ( .A(n5048), .B(n5049), .Z(n5047) );
  NANDN U9126 ( .A(n5050), .B(n5051), .Z(n5049) );
  NANDN U9127 ( .A(n5051), .B(n5050), .Z(n5046) );
  NAND U9128 ( .A(n5052), .B(n5053), .Z(n5041) );
  NANDN U9129 ( .A(n5054), .B(n5055), .Z(n5053) );
  OR U9130 ( .A(n5056), .B(n5057), .Z(n5055) );
  NAND U9131 ( .A(n5057), .B(n5056), .Z(n5052) );
  AND U9132 ( .A(n5058), .B(n5059), .Z(n5043) );
  NANDN U9133 ( .A(n5060), .B(n5061), .Z(n5059) );
  NANDN U9134 ( .A(n5062), .B(n5063), .Z(n5061) );
  NANDN U9135 ( .A(n5063), .B(n5062), .Z(n5058) );
  XOR U9136 ( .A(n5057), .B(n5064), .Z(N29731) );
  XOR U9137 ( .A(n5054), .B(n5056), .Z(n5064) );
  XNOR U9138 ( .A(n5050), .B(n5065), .Z(n5056) );
  XNOR U9139 ( .A(n5048), .B(n5051), .Z(n5065) );
  NAND U9140 ( .A(n5066), .B(n5067), .Z(n5051) );
  NAND U9141 ( .A(n5068), .B(n5069), .Z(n5067) );
  OR U9142 ( .A(n5070), .B(n5071), .Z(n5068) );
  NANDN U9143 ( .A(n5072), .B(n5070), .Z(n5066) );
  IV U9144 ( .A(n5071), .Z(n5072) );
  NAND U9145 ( .A(n5073), .B(n5074), .Z(n5048) );
  NAND U9146 ( .A(n5075), .B(n5076), .Z(n5074) );
  NANDN U9147 ( .A(n5077), .B(n5078), .Z(n5075) );
  NANDN U9148 ( .A(n5078), .B(n5077), .Z(n5073) );
  AND U9149 ( .A(n5079), .B(n5080), .Z(n5050) );
  NAND U9150 ( .A(n5081), .B(n5082), .Z(n5080) );
  OR U9151 ( .A(n5083), .B(n5084), .Z(n5081) );
  NANDN U9152 ( .A(n5085), .B(n5083), .Z(n5079) );
  NAND U9153 ( .A(n5086), .B(n5087), .Z(n5054) );
  NANDN U9154 ( .A(n5088), .B(n5089), .Z(n5087) );
  OR U9155 ( .A(n5090), .B(n5091), .Z(n5089) );
  NANDN U9156 ( .A(n5092), .B(n5090), .Z(n5086) );
  IV U9157 ( .A(n5091), .Z(n5092) );
  XNOR U9158 ( .A(n5062), .B(n5093), .Z(n5057) );
  XNOR U9159 ( .A(n5060), .B(n5063), .Z(n5093) );
  NAND U9160 ( .A(n5094), .B(n5095), .Z(n5063) );
  NAND U9161 ( .A(n5096), .B(n5097), .Z(n5095) );
  OR U9162 ( .A(n5098), .B(n5099), .Z(n5096) );
  NANDN U9163 ( .A(n5100), .B(n5098), .Z(n5094) );
  IV U9164 ( .A(n5099), .Z(n5100) );
  NAND U9165 ( .A(n5101), .B(n5102), .Z(n5060) );
  NAND U9166 ( .A(n5103), .B(n5104), .Z(n5102) );
  NANDN U9167 ( .A(n5105), .B(n5106), .Z(n5103) );
  NANDN U9168 ( .A(n5106), .B(n5105), .Z(n5101) );
  AND U9169 ( .A(n5107), .B(n5108), .Z(n5062) );
  NAND U9170 ( .A(n5109), .B(n5110), .Z(n5108) );
  OR U9171 ( .A(n5111), .B(n5112), .Z(n5109) );
  NANDN U9172 ( .A(n5113), .B(n5111), .Z(n5107) );
  XNOR U9173 ( .A(n5088), .B(n5114), .Z(N29730) );
  XOR U9174 ( .A(n5090), .B(n5091), .Z(n5114) );
  XNOR U9175 ( .A(n5104), .B(n5115), .Z(n5091) );
  XOR U9176 ( .A(n5105), .B(n5106), .Z(n5115) );
  XOR U9177 ( .A(n5111), .B(n5116), .Z(n5106) );
  XOR U9178 ( .A(n5110), .B(n5113), .Z(n5116) );
  IV U9179 ( .A(n5112), .Z(n5113) );
  NAND U9180 ( .A(n5117), .B(n5118), .Z(n5112) );
  OR U9181 ( .A(n5119), .B(n5120), .Z(n5118) );
  OR U9182 ( .A(n5121), .B(n5122), .Z(n5117) );
  NAND U9183 ( .A(n5123), .B(n5124), .Z(n5110) );
  OR U9184 ( .A(n5125), .B(n5126), .Z(n5124) );
  OR U9185 ( .A(n5127), .B(n5128), .Z(n5123) );
  NOR U9186 ( .A(n5129), .B(n5130), .Z(n5111) );
  ANDN U9187 ( .B(n5131), .A(n5132), .Z(n5105) );
  XNOR U9188 ( .A(n5098), .B(n5133), .Z(n5104) );
  XNOR U9189 ( .A(n5097), .B(n5099), .Z(n5133) );
  NAND U9190 ( .A(n5134), .B(n5135), .Z(n5099) );
  OR U9191 ( .A(n5136), .B(n5137), .Z(n5135) );
  OR U9192 ( .A(n5138), .B(n5139), .Z(n5134) );
  NAND U9193 ( .A(n5140), .B(n5141), .Z(n5097) );
  OR U9194 ( .A(n5142), .B(n5143), .Z(n5141) );
  OR U9195 ( .A(n5144), .B(n5145), .Z(n5140) );
  ANDN U9196 ( .B(n5146), .A(n5147), .Z(n5098) );
  IV U9197 ( .A(n5148), .Z(n5146) );
  ANDN U9198 ( .B(n5149), .A(n5150), .Z(n5090) );
  XOR U9199 ( .A(n5076), .B(n5151), .Z(n5088) );
  XOR U9200 ( .A(n5077), .B(n5078), .Z(n5151) );
  XOR U9201 ( .A(n5083), .B(n5152), .Z(n5078) );
  XOR U9202 ( .A(n5082), .B(n5085), .Z(n5152) );
  IV U9203 ( .A(n5084), .Z(n5085) );
  NAND U9204 ( .A(n5153), .B(n5154), .Z(n5084) );
  OR U9205 ( .A(n5155), .B(n5156), .Z(n5154) );
  OR U9206 ( .A(n5157), .B(n5158), .Z(n5153) );
  NAND U9207 ( .A(n5159), .B(n5160), .Z(n5082) );
  OR U9208 ( .A(n5161), .B(n5162), .Z(n5160) );
  OR U9209 ( .A(n5163), .B(n5164), .Z(n5159) );
  NOR U9210 ( .A(n5165), .B(n5166), .Z(n5083) );
  ANDN U9211 ( .B(n5167), .A(n5168), .Z(n5077) );
  IV U9212 ( .A(n5169), .Z(n5167) );
  XNOR U9213 ( .A(n5070), .B(n5170), .Z(n5076) );
  XNOR U9214 ( .A(n5069), .B(n5071), .Z(n5170) );
  NAND U9215 ( .A(n5171), .B(n5172), .Z(n5071) );
  OR U9216 ( .A(n5173), .B(n5174), .Z(n5172) );
  OR U9217 ( .A(n5175), .B(n5176), .Z(n5171) );
  NAND U9218 ( .A(n5177), .B(n5178), .Z(n5069) );
  OR U9219 ( .A(n5179), .B(n5180), .Z(n5178) );
  OR U9220 ( .A(n5181), .B(n5182), .Z(n5177) );
  ANDN U9221 ( .B(n5183), .A(n5184), .Z(n5070) );
  IV U9222 ( .A(n5185), .Z(n5183) );
  XNOR U9223 ( .A(n5150), .B(n5149), .Z(N29729) );
  XOR U9224 ( .A(n5169), .B(n5168), .Z(n5149) );
  XNOR U9225 ( .A(n5184), .B(n5185), .Z(n5168) );
  XNOR U9226 ( .A(n5179), .B(n5180), .Z(n5185) );
  XNOR U9227 ( .A(n5181), .B(n5182), .Z(n5180) );
  XNOR U9228 ( .A(y[3604]), .B(x[3604]), .Z(n5182) );
  XNOR U9229 ( .A(y[3605]), .B(x[3605]), .Z(n5181) );
  XNOR U9230 ( .A(y[3603]), .B(x[3603]), .Z(n5179) );
  XNOR U9231 ( .A(n5173), .B(n5174), .Z(n5184) );
  XNOR U9232 ( .A(y[3600]), .B(x[3600]), .Z(n5174) );
  XNOR U9233 ( .A(n5175), .B(n5176), .Z(n5173) );
  XNOR U9234 ( .A(y[3601]), .B(x[3601]), .Z(n5176) );
  XNOR U9235 ( .A(y[3602]), .B(x[3602]), .Z(n5175) );
  XNOR U9236 ( .A(n5166), .B(n5165), .Z(n5169) );
  XNOR U9237 ( .A(n5161), .B(n5162), .Z(n5165) );
  XNOR U9238 ( .A(y[3597]), .B(x[3597]), .Z(n5162) );
  XNOR U9239 ( .A(n5163), .B(n5164), .Z(n5161) );
  XNOR U9240 ( .A(y[3598]), .B(x[3598]), .Z(n5164) );
  XNOR U9241 ( .A(y[3599]), .B(x[3599]), .Z(n5163) );
  XNOR U9242 ( .A(n5155), .B(n5156), .Z(n5166) );
  XNOR U9243 ( .A(y[3594]), .B(x[3594]), .Z(n5156) );
  XNOR U9244 ( .A(n5157), .B(n5158), .Z(n5155) );
  XNOR U9245 ( .A(y[3595]), .B(x[3595]), .Z(n5158) );
  XNOR U9246 ( .A(y[3596]), .B(x[3596]), .Z(n5157) );
  XOR U9247 ( .A(n5131), .B(n5132), .Z(n5150) );
  XNOR U9248 ( .A(n5147), .B(n5148), .Z(n5132) );
  XNOR U9249 ( .A(n5142), .B(n5143), .Z(n5148) );
  XNOR U9250 ( .A(n5144), .B(n5145), .Z(n5143) );
  XNOR U9251 ( .A(y[3592]), .B(x[3592]), .Z(n5145) );
  XNOR U9252 ( .A(y[3593]), .B(x[3593]), .Z(n5144) );
  XNOR U9253 ( .A(y[3591]), .B(x[3591]), .Z(n5142) );
  XNOR U9254 ( .A(n5136), .B(n5137), .Z(n5147) );
  XNOR U9255 ( .A(y[3588]), .B(x[3588]), .Z(n5137) );
  XNOR U9256 ( .A(n5138), .B(n5139), .Z(n5136) );
  XNOR U9257 ( .A(y[3589]), .B(x[3589]), .Z(n5139) );
  XNOR U9258 ( .A(y[3590]), .B(x[3590]), .Z(n5138) );
  XOR U9259 ( .A(n5130), .B(n5129), .Z(n5131) );
  XNOR U9260 ( .A(n5125), .B(n5126), .Z(n5129) );
  XNOR U9261 ( .A(y[3585]), .B(x[3585]), .Z(n5126) );
  XNOR U9262 ( .A(n5127), .B(n5128), .Z(n5125) );
  XNOR U9263 ( .A(y[3586]), .B(x[3586]), .Z(n5128) );
  XNOR U9264 ( .A(y[3587]), .B(x[3587]), .Z(n5127) );
  XNOR U9265 ( .A(n5119), .B(n5120), .Z(n5130) );
  XNOR U9266 ( .A(y[3582]), .B(x[3582]), .Z(n5120) );
  XNOR U9267 ( .A(n5121), .B(n5122), .Z(n5119) );
  XNOR U9268 ( .A(y[3583]), .B(x[3583]), .Z(n5122) );
  XNOR U9269 ( .A(y[3584]), .B(x[3584]), .Z(n5121) );
  NAND U9270 ( .A(n5186), .B(n5187), .Z(N29721) );
  NANDN U9271 ( .A(n5188), .B(n5189), .Z(n5187) );
  OR U9272 ( .A(n5190), .B(n5191), .Z(n5189) );
  NAND U9273 ( .A(n5190), .B(n5191), .Z(n5186) );
  XOR U9274 ( .A(n5190), .B(n5192), .Z(N29720) );
  XNOR U9275 ( .A(n5188), .B(n5191), .Z(n5192) );
  AND U9276 ( .A(n5193), .B(n5194), .Z(n5191) );
  NANDN U9277 ( .A(n5195), .B(n5196), .Z(n5194) );
  NANDN U9278 ( .A(n5197), .B(n5198), .Z(n5196) );
  NANDN U9279 ( .A(n5198), .B(n5197), .Z(n5193) );
  NAND U9280 ( .A(n5199), .B(n5200), .Z(n5188) );
  NANDN U9281 ( .A(n5201), .B(n5202), .Z(n5200) );
  OR U9282 ( .A(n5203), .B(n5204), .Z(n5202) );
  NAND U9283 ( .A(n5204), .B(n5203), .Z(n5199) );
  AND U9284 ( .A(n5205), .B(n5206), .Z(n5190) );
  NANDN U9285 ( .A(n5207), .B(n5208), .Z(n5206) );
  NANDN U9286 ( .A(n5209), .B(n5210), .Z(n5208) );
  NANDN U9287 ( .A(n5210), .B(n5209), .Z(n5205) );
  XOR U9288 ( .A(n5204), .B(n5211), .Z(N29719) );
  XOR U9289 ( .A(n5201), .B(n5203), .Z(n5211) );
  XNOR U9290 ( .A(n5197), .B(n5212), .Z(n5203) );
  XNOR U9291 ( .A(n5195), .B(n5198), .Z(n5212) );
  NAND U9292 ( .A(n5213), .B(n5214), .Z(n5198) );
  NAND U9293 ( .A(n5215), .B(n5216), .Z(n5214) );
  OR U9294 ( .A(n5217), .B(n5218), .Z(n5215) );
  NANDN U9295 ( .A(n5219), .B(n5217), .Z(n5213) );
  IV U9296 ( .A(n5218), .Z(n5219) );
  NAND U9297 ( .A(n5220), .B(n5221), .Z(n5195) );
  NAND U9298 ( .A(n5222), .B(n5223), .Z(n5221) );
  NANDN U9299 ( .A(n5224), .B(n5225), .Z(n5222) );
  NANDN U9300 ( .A(n5225), .B(n5224), .Z(n5220) );
  AND U9301 ( .A(n5226), .B(n5227), .Z(n5197) );
  NAND U9302 ( .A(n5228), .B(n5229), .Z(n5227) );
  OR U9303 ( .A(n5230), .B(n5231), .Z(n5228) );
  NANDN U9304 ( .A(n5232), .B(n5230), .Z(n5226) );
  NAND U9305 ( .A(n5233), .B(n5234), .Z(n5201) );
  NANDN U9306 ( .A(n5235), .B(n5236), .Z(n5234) );
  OR U9307 ( .A(n5237), .B(n5238), .Z(n5236) );
  NANDN U9308 ( .A(n5239), .B(n5237), .Z(n5233) );
  IV U9309 ( .A(n5238), .Z(n5239) );
  XNOR U9310 ( .A(n5209), .B(n5240), .Z(n5204) );
  XNOR U9311 ( .A(n5207), .B(n5210), .Z(n5240) );
  NAND U9312 ( .A(n5241), .B(n5242), .Z(n5210) );
  NAND U9313 ( .A(n5243), .B(n5244), .Z(n5242) );
  OR U9314 ( .A(n5245), .B(n5246), .Z(n5243) );
  NANDN U9315 ( .A(n5247), .B(n5245), .Z(n5241) );
  IV U9316 ( .A(n5246), .Z(n5247) );
  NAND U9317 ( .A(n5248), .B(n5249), .Z(n5207) );
  NAND U9318 ( .A(n5250), .B(n5251), .Z(n5249) );
  NANDN U9319 ( .A(n5252), .B(n5253), .Z(n5250) );
  NANDN U9320 ( .A(n5253), .B(n5252), .Z(n5248) );
  AND U9321 ( .A(n5254), .B(n5255), .Z(n5209) );
  NAND U9322 ( .A(n5256), .B(n5257), .Z(n5255) );
  OR U9323 ( .A(n5258), .B(n5259), .Z(n5256) );
  NANDN U9324 ( .A(n5260), .B(n5258), .Z(n5254) );
  XNOR U9325 ( .A(n5235), .B(n5261), .Z(N29718) );
  XOR U9326 ( .A(n5237), .B(n5238), .Z(n5261) );
  XNOR U9327 ( .A(n5251), .B(n5262), .Z(n5238) );
  XOR U9328 ( .A(n5252), .B(n5253), .Z(n5262) );
  XOR U9329 ( .A(n5258), .B(n5263), .Z(n5253) );
  XOR U9330 ( .A(n5257), .B(n5260), .Z(n5263) );
  IV U9331 ( .A(n5259), .Z(n5260) );
  NAND U9332 ( .A(n5264), .B(n5265), .Z(n5259) );
  OR U9333 ( .A(n5266), .B(n5267), .Z(n5265) );
  OR U9334 ( .A(n5268), .B(n5269), .Z(n5264) );
  NAND U9335 ( .A(n5270), .B(n5271), .Z(n5257) );
  OR U9336 ( .A(n5272), .B(n5273), .Z(n5271) );
  OR U9337 ( .A(n5274), .B(n5275), .Z(n5270) );
  NOR U9338 ( .A(n5276), .B(n5277), .Z(n5258) );
  ANDN U9339 ( .B(n5278), .A(n5279), .Z(n5252) );
  XNOR U9340 ( .A(n5245), .B(n5280), .Z(n5251) );
  XNOR U9341 ( .A(n5244), .B(n5246), .Z(n5280) );
  NAND U9342 ( .A(n5281), .B(n5282), .Z(n5246) );
  OR U9343 ( .A(n5283), .B(n5284), .Z(n5282) );
  OR U9344 ( .A(n5285), .B(n5286), .Z(n5281) );
  NAND U9345 ( .A(n5287), .B(n5288), .Z(n5244) );
  OR U9346 ( .A(n5289), .B(n5290), .Z(n5288) );
  OR U9347 ( .A(n5291), .B(n5292), .Z(n5287) );
  ANDN U9348 ( .B(n5293), .A(n5294), .Z(n5245) );
  IV U9349 ( .A(n5295), .Z(n5293) );
  ANDN U9350 ( .B(n5296), .A(n5297), .Z(n5237) );
  XOR U9351 ( .A(n5223), .B(n5298), .Z(n5235) );
  XOR U9352 ( .A(n5224), .B(n5225), .Z(n5298) );
  XOR U9353 ( .A(n5230), .B(n5299), .Z(n5225) );
  XOR U9354 ( .A(n5229), .B(n5232), .Z(n5299) );
  IV U9355 ( .A(n5231), .Z(n5232) );
  NAND U9356 ( .A(n5300), .B(n5301), .Z(n5231) );
  OR U9357 ( .A(n5302), .B(n5303), .Z(n5301) );
  OR U9358 ( .A(n5304), .B(n5305), .Z(n5300) );
  NAND U9359 ( .A(n5306), .B(n5307), .Z(n5229) );
  OR U9360 ( .A(n5308), .B(n5309), .Z(n5307) );
  OR U9361 ( .A(n5310), .B(n5311), .Z(n5306) );
  NOR U9362 ( .A(n5312), .B(n5313), .Z(n5230) );
  ANDN U9363 ( .B(n5314), .A(n5315), .Z(n5224) );
  IV U9364 ( .A(n5316), .Z(n5314) );
  XNOR U9365 ( .A(n5217), .B(n5317), .Z(n5223) );
  XNOR U9366 ( .A(n5216), .B(n5218), .Z(n5317) );
  NAND U9367 ( .A(n5318), .B(n5319), .Z(n5218) );
  OR U9368 ( .A(n5320), .B(n5321), .Z(n5319) );
  OR U9369 ( .A(n5322), .B(n5323), .Z(n5318) );
  NAND U9370 ( .A(n5324), .B(n5325), .Z(n5216) );
  OR U9371 ( .A(n5326), .B(n5327), .Z(n5325) );
  OR U9372 ( .A(n5328), .B(n5329), .Z(n5324) );
  ANDN U9373 ( .B(n5330), .A(n5331), .Z(n5217) );
  IV U9374 ( .A(n5332), .Z(n5330) );
  XNOR U9375 ( .A(n5297), .B(n5296), .Z(N29717) );
  XOR U9376 ( .A(n5316), .B(n5315), .Z(n5296) );
  XNOR U9377 ( .A(n5331), .B(n5332), .Z(n5315) );
  XNOR U9378 ( .A(n5326), .B(n5327), .Z(n5332) );
  XNOR U9379 ( .A(n5328), .B(n5329), .Z(n5327) );
  XNOR U9380 ( .A(y[3580]), .B(x[3580]), .Z(n5329) );
  XNOR U9381 ( .A(y[3581]), .B(x[3581]), .Z(n5328) );
  XNOR U9382 ( .A(y[3579]), .B(x[3579]), .Z(n5326) );
  XNOR U9383 ( .A(n5320), .B(n5321), .Z(n5331) );
  XNOR U9384 ( .A(y[3576]), .B(x[3576]), .Z(n5321) );
  XNOR U9385 ( .A(n5322), .B(n5323), .Z(n5320) );
  XNOR U9386 ( .A(y[3577]), .B(x[3577]), .Z(n5323) );
  XNOR U9387 ( .A(y[3578]), .B(x[3578]), .Z(n5322) );
  XNOR U9388 ( .A(n5313), .B(n5312), .Z(n5316) );
  XNOR U9389 ( .A(n5308), .B(n5309), .Z(n5312) );
  XNOR U9390 ( .A(y[3573]), .B(x[3573]), .Z(n5309) );
  XNOR U9391 ( .A(n5310), .B(n5311), .Z(n5308) );
  XNOR U9392 ( .A(y[3574]), .B(x[3574]), .Z(n5311) );
  XNOR U9393 ( .A(y[3575]), .B(x[3575]), .Z(n5310) );
  XNOR U9394 ( .A(n5302), .B(n5303), .Z(n5313) );
  XNOR U9395 ( .A(y[3570]), .B(x[3570]), .Z(n5303) );
  XNOR U9396 ( .A(n5304), .B(n5305), .Z(n5302) );
  XNOR U9397 ( .A(y[3571]), .B(x[3571]), .Z(n5305) );
  XNOR U9398 ( .A(y[3572]), .B(x[3572]), .Z(n5304) );
  XOR U9399 ( .A(n5278), .B(n5279), .Z(n5297) );
  XNOR U9400 ( .A(n5294), .B(n5295), .Z(n5279) );
  XNOR U9401 ( .A(n5289), .B(n5290), .Z(n5295) );
  XNOR U9402 ( .A(n5291), .B(n5292), .Z(n5290) );
  XNOR U9403 ( .A(y[3568]), .B(x[3568]), .Z(n5292) );
  XNOR U9404 ( .A(y[3569]), .B(x[3569]), .Z(n5291) );
  XNOR U9405 ( .A(y[3567]), .B(x[3567]), .Z(n5289) );
  XNOR U9406 ( .A(n5283), .B(n5284), .Z(n5294) );
  XNOR U9407 ( .A(y[3564]), .B(x[3564]), .Z(n5284) );
  XNOR U9408 ( .A(n5285), .B(n5286), .Z(n5283) );
  XNOR U9409 ( .A(y[3565]), .B(x[3565]), .Z(n5286) );
  XNOR U9410 ( .A(y[3566]), .B(x[3566]), .Z(n5285) );
  XOR U9411 ( .A(n5277), .B(n5276), .Z(n5278) );
  XNOR U9412 ( .A(n5272), .B(n5273), .Z(n5276) );
  XNOR U9413 ( .A(y[3561]), .B(x[3561]), .Z(n5273) );
  XNOR U9414 ( .A(n5274), .B(n5275), .Z(n5272) );
  XNOR U9415 ( .A(y[3562]), .B(x[3562]), .Z(n5275) );
  XNOR U9416 ( .A(y[3563]), .B(x[3563]), .Z(n5274) );
  XNOR U9417 ( .A(n5266), .B(n5267), .Z(n5277) );
  XNOR U9418 ( .A(y[3558]), .B(x[3558]), .Z(n5267) );
  XNOR U9419 ( .A(n5268), .B(n5269), .Z(n5266) );
  XNOR U9420 ( .A(y[3559]), .B(x[3559]), .Z(n5269) );
  XNOR U9421 ( .A(y[3560]), .B(x[3560]), .Z(n5268) );
  NAND U9422 ( .A(n5333), .B(n5334), .Z(N29709) );
  NANDN U9423 ( .A(n5335), .B(n5336), .Z(n5334) );
  OR U9424 ( .A(n5337), .B(n5338), .Z(n5336) );
  NAND U9425 ( .A(n5337), .B(n5338), .Z(n5333) );
  XOR U9426 ( .A(n5337), .B(n5339), .Z(N29708) );
  XNOR U9427 ( .A(n5335), .B(n5338), .Z(n5339) );
  AND U9428 ( .A(n5340), .B(n5341), .Z(n5338) );
  NANDN U9429 ( .A(n5342), .B(n5343), .Z(n5341) );
  NANDN U9430 ( .A(n5344), .B(n5345), .Z(n5343) );
  NANDN U9431 ( .A(n5345), .B(n5344), .Z(n5340) );
  NAND U9432 ( .A(n5346), .B(n5347), .Z(n5335) );
  NANDN U9433 ( .A(n5348), .B(n5349), .Z(n5347) );
  OR U9434 ( .A(n5350), .B(n5351), .Z(n5349) );
  NAND U9435 ( .A(n5351), .B(n5350), .Z(n5346) );
  AND U9436 ( .A(n5352), .B(n5353), .Z(n5337) );
  NANDN U9437 ( .A(n5354), .B(n5355), .Z(n5353) );
  NANDN U9438 ( .A(n5356), .B(n5357), .Z(n5355) );
  NANDN U9439 ( .A(n5357), .B(n5356), .Z(n5352) );
  XOR U9440 ( .A(n5351), .B(n5358), .Z(N29707) );
  XOR U9441 ( .A(n5348), .B(n5350), .Z(n5358) );
  XNOR U9442 ( .A(n5344), .B(n5359), .Z(n5350) );
  XNOR U9443 ( .A(n5342), .B(n5345), .Z(n5359) );
  NAND U9444 ( .A(n5360), .B(n5361), .Z(n5345) );
  NAND U9445 ( .A(n5362), .B(n5363), .Z(n5361) );
  OR U9446 ( .A(n5364), .B(n5365), .Z(n5362) );
  NANDN U9447 ( .A(n5366), .B(n5364), .Z(n5360) );
  IV U9448 ( .A(n5365), .Z(n5366) );
  NAND U9449 ( .A(n5367), .B(n5368), .Z(n5342) );
  NAND U9450 ( .A(n5369), .B(n5370), .Z(n5368) );
  NANDN U9451 ( .A(n5371), .B(n5372), .Z(n5369) );
  NANDN U9452 ( .A(n5372), .B(n5371), .Z(n5367) );
  AND U9453 ( .A(n5373), .B(n5374), .Z(n5344) );
  NAND U9454 ( .A(n5375), .B(n5376), .Z(n5374) );
  OR U9455 ( .A(n5377), .B(n5378), .Z(n5375) );
  NANDN U9456 ( .A(n5379), .B(n5377), .Z(n5373) );
  NAND U9457 ( .A(n5380), .B(n5381), .Z(n5348) );
  NANDN U9458 ( .A(n5382), .B(n5383), .Z(n5381) );
  OR U9459 ( .A(n5384), .B(n5385), .Z(n5383) );
  NANDN U9460 ( .A(n5386), .B(n5384), .Z(n5380) );
  IV U9461 ( .A(n5385), .Z(n5386) );
  XNOR U9462 ( .A(n5356), .B(n5387), .Z(n5351) );
  XNOR U9463 ( .A(n5354), .B(n5357), .Z(n5387) );
  NAND U9464 ( .A(n5388), .B(n5389), .Z(n5357) );
  NAND U9465 ( .A(n5390), .B(n5391), .Z(n5389) );
  OR U9466 ( .A(n5392), .B(n5393), .Z(n5390) );
  NANDN U9467 ( .A(n5394), .B(n5392), .Z(n5388) );
  IV U9468 ( .A(n5393), .Z(n5394) );
  NAND U9469 ( .A(n5395), .B(n5396), .Z(n5354) );
  NAND U9470 ( .A(n5397), .B(n5398), .Z(n5396) );
  NANDN U9471 ( .A(n5399), .B(n5400), .Z(n5397) );
  NANDN U9472 ( .A(n5400), .B(n5399), .Z(n5395) );
  AND U9473 ( .A(n5401), .B(n5402), .Z(n5356) );
  NAND U9474 ( .A(n5403), .B(n5404), .Z(n5402) );
  OR U9475 ( .A(n5405), .B(n5406), .Z(n5403) );
  NANDN U9476 ( .A(n5407), .B(n5405), .Z(n5401) );
  XNOR U9477 ( .A(n5382), .B(n5408), .Z(N29706) );
  XOR U9478 ( .A(n5384), .B(n5385), .Z(n5408) );
  XNOR U9479 ( .A(n5398), .B(n5409), .Z(n5385) );
  XOR U9480 ( .A(n5399), .B(n5400), .Z(n5409) );
  XOR U9481 ( .A(n5405), .B(n5410), .Z(n5400) );
  XOR U9482 ( .A(n5404), .B(n5407), .Z(n5410) );
  IV U9483 ( .A(n5406), .Z(n5407) );
  NAND U9484 ( .A(n5411), .B(n5412), .Z(n5406) );
  OR U9485 ( .A(n5413), .B(n5414), .Z(n5412) );
  OR U9486 ( .A(n5415), .B(n5416), .Z(n5411) );
  NAND U9487 ( .A(n5417), .B(n5418), .Z(n5404) );
  OR U9488 ( .A(n5419), .B(n5420), .Z(n5418) );
  OR U9489 ( .A(n5421), .B(n5422), .Z(n5417) );
  NOR U9490 ( .A(n5423), .B(n5424), .Z(n5405) );
  ANDN U9491 ( .B(n5425), .A(n5426), .Z(n5399) );
  XNOR U9492 ( .A(n5392), .B(n5427), .Z(n5398) );
  XNOR U9493 ( .A(n5391), .B(n5393), .Z(n5427) );
  NAND U9494 ( .A(n5428), .B(n5429), .Z(n5393) );
  OR U9495 ( .A(n5430), .B(n5431), .Z(n5429) );
  OR U9496 ( .A(n5432), .B(n5433), .Z(n5428) );
  NAND U9497 ( .A(n5434), .B(n5435), .Z(n5391) );
  OR U9498 ( .A(n5436), .B(n5437), .Z(n5435) );
  OR U9499 ( .A(n5438), .B(n5439), .Z(n5434) );
  ANDN U9500 ( .B(n5440), .A(n5441), .Z(n5392) );
  IV U9501 ( .A(n5442), .Z(n5440) );
  ANDN U9502 ( .B(n5443), .A(n5444), .Z(n5384) );
  XOR U9503 ( .A(n5370), .B(n5445), .Z(n5382) );
  XOR U9504 ( .A(n5371), .B(n5372), .Z(n5445) );
  XOR U9505 ( .A(n5377), .B(n5446), .Z(n5372) );
  XOR U9506 ( .A(n5376), .B(n5379), .Z(n5446) );
  IV U9507 ( .A(n5378), .Z(n5379) );
  NAND U9508 ( .A(n5447), .B(n5448), .Z(n5378) );
  OR U9509 ( .A(n5449), .B(n5450), .Z(n5448) );
  OR U9510 ( .A(n5451), .B(n5452), .Z(n5447) );
  NAND U9511 ( .A(n5453), .B(n5454), .Z(n5376) );
  OR U9512 ( .A(n5455), .B(n5456), .Z(n5454) );
  OR U9513 ( .A(n5457), .B(n5458), .Z(n5453) );
  NOR U9514 ( .A(n5459), .B(n5460), .Z(n5377) );
  ANDN U9515 ( .B(n5461), .A(n5462), .Z(n5371) );
  IV U9516 ( .A(n5463), .Z(n5461) );
  XNOR U9517 ( .A(n5364), .B(n5464), .Z(n5370) );
  XNOR U9518 ( .A(n5363), .B(n5365), .Z(n5464) );
  NAND U9519 ( .A(n5465), .B(n5466), .Z(n5365) );
  OR U9520 ( .A(n5467), .B(n5468), .Z(n5466) );
  OR U9521 ( .A(n5469), .B(n5470), .Z(n5465) );
  NAND U9522 ( .A(n5471), .B(n5472), .Z(n5363) );
  OR U9523 ( .A(n5473), .B(n5474), .Z(n5472) );
  OR U9524 ( .A(n5475), .B(n5476), .Z(n5471) );
  ANDN U9525 ( .B(n5477), .A(n5478), .Z(n5364) );
  IV U9526 ( .A(n5479), .Z(n5477) );
  XNOR U9527 ( .A(n5444), .B(n5443), .Z(N29705) );
  XOR U9528 ( .A(n5463), .B(n5462), .Z(n5443) );
  XNOR U9529 ( .A(n5478), .B(n5479), .Z(n5462) );
  XNOR U9530 ( .A(n5473), .B(n5474), .Z(n5479) );
  XNOR U9531 ( .A(n5475), .B(n5476), .Z(n5474) );
  XNOR U9532 ( .A(y[3556]), .B(x[3556]), .Z(n5476) );
  XNOR U9533 ( .A(y[3557]), .B(x[3557]), .Z(n5475) );
  XNOR U9534 ( .A(y[3555]), .B(x[3555]), .Z(n5473) );
  XNOR U9535 ( .A(n5467), .B(n5468), .Z(n5478) );
  XNOR U9536 ( .A(y[3552]), .B(x[3552]), .Z(n5468) );
  XNOR U9537 ( .A(n5469), .B(n5470), .Z(n5467) );
  XNOR U9538 ( .A(y[3553]), .B(x[3553]), .Z(n5470) );
  XNOR U9539 ( .A(y[3554]), .B(x[3554]), .Z(n5469) );
  XNOR U9540 ( .A(n5460), .B(n5459), .Z(n5463) );
  XNOR U9541 ( .A(n5455), .B(n5456), .Z(n5459) );
  XNOR U9542 ( .A(y[3549]), .B(x[3549]), .Z(n5456) );
  XNOR U9543 ( .A(n5457), .B(n5458), .Z(n5455) );
  XNOR U9544 ( .A(y[3550]), .B(x[3550]), .Z(n5458) );
  XNOR U9545 ( .A(y[3551]), .B(x[3551]), .Z(n5457) );
  XNOR U9546 ( .A(n5449), .B(n5450), .Z(n5460) );
  XNOR U9547 ( .A(y[3546]), .B(x[3546]), .Z(n5450) );
  XNOR U9548 ( .A(n5451), .B(n5452), .Z(n5449) );
  XNOR U9549 ( .A(y[3547]), .B(x[3547]), .Z(n5452) );
  XNOR U9550 ( .A(y[3548]), .B(x[3548]), .Z(n5451) );
  XOR U9551 ( .A(n5425), .B(n5426), .Z(n5444) );
  XNOR U9552 ( .A(n5441), .B(n5442), .Z(n5426) );
  XNOR U9553 ( .A(n5436), .B(n5437), .Z(n5442) );
  XNOR U9554 ( .A(n5438), .B(n5439), .Z(n5437) );
  XNOR U9555 ( .A(y[3544]), .B(x[3544]), .Z(n5439) );
  XNOR U9556 ( .A(y[3545]), .B(x[3545]), .Z(n5438) );
  XNOR U9557 ( .A(y[3543]), .B(x[3543]), .Z(n5436) );
  XNOR U9558 ( .A(n5430), .B(n5431), .Z(n5441) );
  XNOR U9559 ( .A(y[3540]), .B(x[3540]), .Z(n5431) );
  XNOR U9560 ( .A(n5432), .B(n5433), .Z(n5430) );
  XNOR U9561 ( .A(y[3541]), .B(x[3541]), .Z(n5433) );
  XNOR U9562 ( .A(y[3542]), .B(x[3542]), .Z(n5432) );
  XOR U9563 ( .A(n5424), .B(n5423), .Z(n5425) );
  XNOR U9564 ( .A(n5419), .B(n5420), .Z(n5423) );
  XNOR U9565 ( .A(y[3537]), .B(x[3537]), .Z(n5420) );
  XNOR U9566 ( .A(n5421), .B(n5422), .Z(n5419) );
  XNOR U9567 ( .A(y[3538]), .B(x[3538]), .Z(n5422) );
  XNOR U9568 ( .A(y[3539]), .B(x[3539]), .Z(n5421) );
  XNOR U9569 ( .A(n5413), .B(n5414), .Z(n5424) );
  XNOR U9570 ( .A(y[3534]), .B(x[3534]), .Z(n5414) );
  XNOR U9571 ( .A(n5415), .B(n5416), .Z(n5413) );
  XNOR U9572 ( .A(y[3535]), .B(x[3535]), .Z(n5416) );
  XNOR U9573 ( .A(y[3536]), .B(x[3536]), .Z(n5415) );
  NAND U9574 ( .A(n5480), .B(n5481), .Z(N29697) );
  NANDN U9575 ( .A(n5482), .B(n5483), .Z(n5481) );
  OR U9576 ( .A(n5484), .B(n5485), .Z(n5483) );
  NAND U9577 ( .A(n5484), .B(n5485), .Z(n5480) );
  XOR U9578 ( .A(n5484), .B(n5486), .Z(N29696) );
  XNOR U9579 ( .A(n5482), .B(n5485), .Z(n5486) );
  AND U9580 ( .A(n5487), .B(n5488), .Z(n5485) );
  NANDN U9581 ( .A(n5489), .B(n5490), .Z(n5488) );
  NANDN U9582 ( .A(n5491), .B(n5492), .Z(n5490) );
  NANDN U9583 ( .A(n5492), .B(n5491), .Z(n5487) );
  NAND U9584 ( .A(n5493), .B(n5494), .Z(n5482) );
  NANDN U9585 ( .A(n5495), .B(n5496), .Z(n5494) );
  OR U9586 ( .A(n5497), .B(n5498), .Z(n5496) );
  NAND U9587 ( .A(n5498), .B(n5497), .Z(n5493) );
  AND U9588 ( .A(n5499), .B(n5500), .Z(n5484) );
  NANDN U9589 ( .A(n5501), .B(n5502), .Z(n5500) );
  NANDN U9590 ( .A(n5503), .B(n5504), .Z(n5502) );
  NANDN U9591 ( .A(n5504), .B(n5503), .Z(n5499) );
  XOR U9592 ( .A(n5498), .B(n5505), .Z(N29695) );
  XOR U9593 ( .A(n5495), .B(n5497), .Z(n5505) );
  XNOR U9594 ( .A(n5491), .B(n5506), .Z(n5497) );
  XNOR U9595 ( .A(n5489), .B(n5492), .Z(n5506) );
  NAND U9596 ( .A(n5507), .B(n5508), .Z(n5492) );
  NAND U9597 ( .A(n5509), .B(n5510), .Z(n5508) );
  OR U9598 ( .A(n5511), .B(n5512), .Z(n5509) );
  NANDN U9599 ( .A(n5513), .B(n5511), .Z(n5507) );
  IV U9600 ( .A(n5512), .Z(n5513) );
  NAND U9601 ( .A(n5514), .B(n5515), .Z(n5489) );
  NAND U9602 ( .A(n5516), .B(n5517), .Z(n5515) );
  NANDN U9603 ( .A(n5518), .B(n5519), .Z(n5516) );
  NANDN U9604 ( .A(n5519), .B(n5518), .Z(n5514) );
  AND U9605 ( .A(n5520), .B(n5521), .Z(n5491) );
  NAND U9606 ( .A(n5522), .B(n5523), .Z(n5521) );
  OR U9607 ( .A(n5524), .B(n5525), .Z(n5522) );
  NANDN U9608 ( .A(n5526), .B(n5524), .Z(n5520) );
  NAND U9609 ( .A(n5527), .B(n5528), .Z(n5495) );
  NANDN U9610 ( .A(n5529), .B(n5530), .Z(n5528) );
  OR U9611 ( .A(n5531), .B(n5532), .Z(n5530) );
  NANDN U9612 ( .A(n5533), .B(n5531), .Z(n5527) );
  IV U9613 ( .A(n5532), .Z(n5533) );
  XNOR U9614 ( .A(n5503), .B(n5534), .Z(n5498) );
  XNOR U9615 ( .A(n5501), .B(n5504), .Z(n5534) );
  NAND U9616 ( .A(n5535), .B(n5536), .Z(n5504) );
  NAND U9617 ( .A(n5537), .B(n5538), .Z(n5536) );
  OR U9618 ( .A(n5539), .B(n5540), .Z(n5537) );
  NANDN U9619 ( .A(n5541), .B(n5539), .Z(n5535) );
  IV U9620 ( .A(n5540), .Z(n5541) );
  NAND U9621 ( .A(n5542), .B(n5543), .Z(n5501) );
  NAND U9622 ( .A(n5544), .B(n5545), .Z(n5543) );
  NANDN U9623 ( .A(n5546), .B(n5547), .Z(n5544) );
  NANDN U9624 ( .A(n5547), .B(n5546), .Z(n5542) );
  AND U9625 ( .A(n5548), .B(n5549), .Z(n5503) );
  NAND U9626 ( .A(n5550), .B(n5551), .Z(n5549) );
  OR U9627 ( .A(n5552), .B(n5553), .Z(n5550) );
  NANDN U9628 ( .A(n5554), .B(n5552), .Z(n5548) );
  XNOR U9629 ( .A(n5529), .B(n5555), .Z(N29694) );
  XOR U9630 ( .A(n5531), .B(n5532), .Z(n5555) );
  XNOR U9631 ( .A(n5545), .B(n5556), .Z(n5532) );
  XOR U9632 ( .A(n5546), .B(n5547), .Z(n5556) );
  XOR U9633 ( .A(n5552), .B(n5557), .Z(n5547) );
  XOR U9634 ( .A(n5551), .B(n5554), .Z(n5557) );
  IV U9635 ( .A(n5553), .Z(n5554) );
  NAND U9636 ( .A(n5558), .B(n5559), .Z(n5553) );
  OR U9637 ( .A(n5560), .B(n5561), .Z(n5559) );
  OR U9638 ( .A(n5562), .B(n5563), .Z(n5558) );
  NAND U9639 ( .A(n5564), .B(n5565), .Z(n5551) );
  OR U9640 ( .A(n5566), .B(n5567), .Z(n5565) );
  OR U9641 ( .A(n5568), .B(n5569), .Z(n5564) );
  NOR U9642 ( .A(n5570), .B(n5571), .Z(n5552) );
  ANDN U9643 ( .B(n5572), .A(n5573), .Z(n5546) );
  XNOR U9644 ( .A(n5539), .B(n5574), .Z(n5545) );
  XNOR U9645 ( .A(n5538), .B(n5540), .Z(n5574) );
  NAND U9646 ( .A(n5575), .B(n5576), .Z(n5540) );
  OR U9647 ( .A(n5577), .B(n5578), .Z(n5576) );
  OR U9648 ( .A(n5579), .B(n5580), .Z(n5575) );
  NAND U9649 ( .A(n5581), .B(n5582), .Z(n5538) );
  OR U9650 ( .A(n5583), .B(n5584), .Z(n5582) );
  OR U9651 ( .A(n5585), .B(n5586), .Z(n5581) );
  ANDN U9652 ( .B(n5587), .A(n5588), .Z(n5539) );
  IV U9653 ( .A(n5589), .Z(n5587) );
  ANDN U9654 ( .B(n5590), .A(n5591), .Z(n5531) );
  XOR U9655 ( .A(n5517), .B(n5592), .Z(n5529) );
  XOR U9656 ( .A(n5518), .B(n5519), .Z(n5592) );
  XOR U9657 ( .A(n5524), .B(n5593), .Z(n5519) );
  XOR U9658 ( .A(n5523), .B(n5526), .Z(n5593) );
  IV U9659 ( .A(n5525), .Z(n5526) );
  NAND U9660 ( .A(n5594), .B(n5595), .Z(n5525) );
  OR U9661 ( .A(n5596), .B(n5597), .Z(n5595) );
  OR U9662 ( .A(n5598), .B(n5599), .Z(n5594) );
  NAND U9663 ( .A(n5600), .B(n5601), .Z(n5523) );
  OR U9664 ( .A(n5602), .B(n5603), .Z(n5601) );
  OR U9665 ( .A(n5604), .B(n5605), .Z(n5600) );
  NOR U9666 ( .A(n5606), .B(n5607), .Z(n5524) );
  ANDN U9667 ( .B(n5608), .A(n5609), .Z(n5518) );
  IV U9668 ( .A(n5610), .Z(n5608) );
  XNOR U9669 ( .A(n5511), .B(n5611), .Z(n5517) );
  XNOR U9670 ( .A(n5510), .B(n5512), .Z(n5611) );
  NAND U9671 ( .A(n5612), .B(n5613), .Z(n5512) );
  OR U9672 ( .A(n5614), .B(n5615), .Z(n5613) );
  OR U9673 ( .A(n5616), .B(n5617), .Z(n5612) );
  NAND U9674 ( .A(n5618), .B(n5619), .Z(n5510) );
  OR U9675 ( .A(n5620), .B(n5621), .Z(n5619) );
  OR U9676 ( .A(n5622), .B(n5623), .Z(n5618) );
  ANDN U9677 ( .B(n5624), .A(n5625), .Z(n5511) );
  IV U9678 ( .A(n5626), .Z(n5624) );
  XNOR U9679 ( .A(n5591), .B(n5590), .Z(N29693) );
  XOR U9680 ( .A(n5610), .B(n5609), .Z(n5590) );
  XNOR U9681 ( .A(n5625), .B(n5626), .Z(n5609) );
  XNOR U9682 ( .A(n5620), .B(n5621), .Z(n5626) );
  XNOR U9683 ( .A(n5622), .B(n5623), .Z(n5621) );
  XNOR U9684 ( .A(y[3532]), .B(x[3532]), .Z(n5623) );
  XNOR U9685 ( .A(y[3533]), .B(x[3533]), .Z(n5622) );
  XNOR U9686 ( .A(y[3531]), .B(x[3531]), .Z(n5620) );
  XNOR U9687 ( .A(n5614), .B(n5615), .Z(n5625) );
  XNOR U9688 ( .A(y[3528]), .B(x[3528]), .Z(n5615) );
  XNOR U9689 ( .A(n5616), .B(n5617), .Z(n5614) );
  XNOR U9690 ( .A(y[3529]), .B(x[3529]), .Z(n5617) );
  XNOR U9691 ( .A(y[3530]), .B(x[3530]), .Z(n5616) );
  XNOR U9692 ( .A(n5607), .B(n5606), .Z(n5610) );
  XNOR U9693 ( .A(n5602), .B(n5603), .Z(n5606) );
  XNOR U9694 ( .A(y[3525]), .B(x[3525]), .Z(n5603) );
  XNOR U9695 ( .A(n5604), .B(n5605), .Z(n5602) );
  XNOR U9696 ( .A(y[3526]), .B(x[3526]), .Z(n5605) );
  XNOR U9697 ( .A(y[3527]), .B(x[3527]), .Z(n5604) );
  XNOR U9698 ( .A(n5596), .B(n5597), .Z(n5607) );
  XNOR U9699 ( .A(y[3522]), .B(x[3522]), .Z(n5597) );
  XNOR U9700 ( .A(n5598), .B(n5599), .Z(n5596) );
  XNOR U9701 ( .A(y[3523]), .B(x[3523]), .Z(n5599) );
  XNOR U9702 ( .A(y[3524]), .B(x[3524]), .Z(n5598) );
  XOR U9703 ( .A(n5572), .B(n5573), .Z(n5591) );
  XNOR U9704 ( .A(n5588), .B(n5589), .Z(n5573) );
  XNOR U9705 ( .A(n5583), .B(n5584), .Z(n5589) );
  XNOR U9706 ( .A(n5585), .B(n5586), .Z(n5584) );
  XNOR U9707 ( .A(y[3520]), .B(x[3520]), .Z(n5586) );
  XNOR U9708 ( .A(y[3521]), .B(x[3521]), .Z(n5585) );
  XNOR U9709 ( .A(y[3519]), .B(x[3519]), .Z(n5583) );
  XNOR U9710 ( .A(n5577), .B(n5578), .Z(n5588) );
  XNOR U9711 ( .A(y[3516]), .B(x[3516]), .Z(n5578) );
  XNOR U9712 ( .A(n5579), .B(n5580), .Z(n5577) );
  XNOR U9713 ( .A(y[3517]), .B(x[3517]), .Z(n5580) );
  XNOR U9714 ( .A(y[3518]), .B(x[3518]), .Z(n5579) );
  XOR U9715 ( .A(n5571), .B(n5570), .Z(n5572) );
  XNOR U9716 ( .A(n5566), .B(n5567), .Z(n5570) );
  XNOR U9717 ( .A(y[3513]), .B(x[3513]), .Z(n5567) );
  XNOR U9718 ( .A(n5568), .B(n5569), .Z(n5566) );
  XNOR U9719 ( .A(y[3514]), .B(x[3514]), .Z(n5569) );
  XNOR U9720 ( .A(y[3515]), .B(x[3515]), .Z(n5568) );
  XNOR U9721 ( .A(n5560), .B(n5561), .Z(n5571) );
  XNOR U9722 ( .A(y[3510]), .B(x[3510]), .Z(n5561) );
  XNOR U9723 ( .A(n5562), .B(n5563), .Z(n5560) );
  XNOR U9724 ( .A(y[3511]), .B(x[3511]), .Z(n5563) );
  XNOR U9725 ( .A(y[3512]), .B(x[3512]), .Z(n5562) );
  NAND U9726 ( .A(n5627), .B(n5628), .Z(N29685) );
  NANDN U9727 ( .A(n5629), .B(n5630), .Z(n5628) );
  OR U9728 ( .A(n5631), .B(n5632), .Z(n5630) );
  NAND U9729 ( .A(n5631), .B(n5632), .Z(n5627) );
  XOR U9730 ( .A(n5631), .B(n5633), .Z(N29684) );
  XNOR U9731 ( .A(n5629), .B(n5632), .Z(n5633) );
  AND U9732 ( .A(n5634), .B(n5635), .Z(n5632) );
  NANDN U9733 ( .A(n5636), .B(n5637), .Z(n5635) );
  NANDN U9734 ( .A(n5638), .B(n5639), .Z(n5637) );
  NANDN U9735 ( .A(n5639), .B(n5638), .Z(n5634) );
  NAND U9736 ( .A(n5640), .B(n5641), .Z(n5629) );
  NANDN U9737 ( .A(n5642), .B(n5643), .Z(n5641) );
  OR U9738 ( .A(n5644), .B(n5645), .Z(n5643) );
  NAND U9739 ( .A(n5645), .B(n5644), .Z(n5640) );
  AND U9740 ( .A(n5646), .B(n5647), .Z(n5631) );
  NANDN U9741 ( .A(n5648), .B(n5649), .Z(n5647) );
  NANDN U9742 ( .A(n5650), .B(n5651), .Z(n5649) );
  NANDN U9743 ( .A(n5651), .B(n5650), .Z(n5646) );
  XOR U9744 ( .A(n5645), .B(n5652), .Z(N29683) );
  XOR U9745 ( .A(n5642), .B(n5644), .Z(n5652) );
  XNOR U9746 ( .A(n5638), .B(n5653), .Z(n5644) );
  XNOR U9747 ( .A(n5636), .B(n5639), .Z(n5653) );
  NAND U9748 ( .A(n5654), .B(n5655), .Z(n5639) );
  NAND U9749 ( .A(n5656), .B(n5657), .Z(n5655) );
  OR U9750 ( .A(n5658), .B(n5659), .Z(n5656) );
  NANDN U9751 ( .A(n5660), .B(n5658), .Z(n5654) );
  IV U9752 ( .A(n5659), .Z(n5660) );
  NAND U9753 ( .A(n5661), .B(n5662), .Z(n5636) );
  NAND U9754 ( .A(n5663), .B(n5664), .Z(n5662) );
  NANDN U9755 ( .A(n5665), .B(n5666), .Z(n5663) );
  NANDN U9756 ( .A(n5666), .B(n5665), .Z(n5661) );
  AND U9757 ( .A(n5667), .B(n5668), .Z(n5638) );
  NAND U9758 ( .A(n5669), .B(n5670), .Z(n5668) );
  OR U9759 ( .A(n5671), .B(n5672), .Z(n5669) );
  NANDN U9760 ( .A(n5673), .B(n5671), .Z(n5667) );
  NAND U9761 ( .A(n5674), .B(n5675), .Z(n5642) );
  NANDN U9762 ( .A(n5676), .B(n5677), .Z(n5675) );
  OR U9763 ( .A(n5678), .B(n5679), .Z(n5677) );
  NANDN U9764 ( .A(n5680), .B(n5678), .Z(n5674) );
  IV U9765 ( .A(n5679), .Z(n5680) );
  XNOR U9766 ( .A(n5650), .B(n5681), .Z(n5645) );
  XNOR U9767 ( .A(n5648), .B(n5651), .Z(n5681) );
  NAND U9768 ( .A(n5682), .B(n5683), .Z(n5651) );
  NAND U9769 ( .A(n5684), .B(n5685), .Z(n5683) );
  OR U9770 ( .A(n5686), .B(n5687), .Z(n5684) );
  NANDN U9771 ( .A(n5688), .B(n5686), .Z(n5682) );
  IV U9772 ( .A(n5687), .Z(n5688) );
  NAND U9773 ( .A(n5689), .B(n5690), .Z(n5648) );
  NAND U9774 ( .A(n5691), .B(n5692), .Z(n5690) );
  NANDN U9775 ( .A(n5693), .B(n5694), .Z(n5691) );
  NANDN U9776 ( .A(n5694), .B(n5693), .Z(n5689) );
  AND U9777 ( .A(n5695), .B(n5696), .Z(n5650) );
  NAND U9778 ( .A(n5697), .B(n5698), .Z(n5696) );
  OR U9779 ( .A(n5699), .B(n5700), .Z(n5697) );
  NANDN U9780 ( .A(n5701), .B(n5699), .Z(n5695) );
  XNOR U9781 ( .A(n5676), .B(n5702), .Z(N29682) );
  XOR U9782 ( .A(n5678), .B(n5679), .Z(n5702) );
  XNOR U9783 ( .A(n5692), .B(n5703), .Z(n5679) );
  XOR U9784 ( .A(n5693), .B(n5694), .Z(n5703) );
  XOR U9785 ( .A(n5699), .B(n5704), .Z(n5694) );
  XOR U9786 ( .A(n5698), .B(n5701), .Z(n5704) );
  IV U9787 ( .A(n5700), .Z(n5701) );
  NAND U9788 ( .A(n5705), .B(n5706), .Z(n5700) );
  OR U9789 ( .A(n5707), .B(n5708), .Z(n5706) );
  OR U9790 ( .A(n5709), .B(n5710), .Z(n5705) );
  NAND U9791 ( .A(n5711), .B(n5712), .Z(n5698) );
  OR U9792 ( .A(n5713), .B(n5714), .Z(n5712) );
  OR U9793 ( .A(n5715), .B(n5716), .Z(n5711) );
  NOR U9794 ( .A(n5717), .B(n5718), .Z(n5699) );
  ANDN U9795 ( .B(n5719), .A(n5720), .Z(n5693) );
  XNOR U9796 ( .A(n5686), .B(n5721), .Z(n5692) );
  XNOR U9797 ( .A(n5685), .B(n5687), .Z(n5721) );
  NAND U9798 ( .A(n5722), .B(n5723), .Z(n5687) );
  OR U9799 ( .A(n5724), .B(n5725), .Z(n5723) );
  OR U9800 ( .A(n5726), .B(n5727), .Z(n5722) );
  NAND U9801 ( .A(n5728), .B(n5729), .Z(n5685) );
  OR U9802 ( .A(n5730), .B(n5731), .Z(n5729) );
  OR U9803 ( .A(n5732), .B(n5733), .Z(n5728) );
  ANDN U9804 ( .B(n5734), .A(n5735), .Z(n5686) );
  IV U9805 ( .A(n5736), .Z(n5734) );
  ANDN U9806 ( .B(n5737), .A(n5738), .Z(n5678) );
  XOR U9807 ( .A(n5664), .B(n5739), .Z(n5676) );
  XOR U9808 ( .A(n5665), .B(n5666), .Z(n5739) );
  XOR U9809 ( .A(n5671), .B(n5740), .Z(n5666) );
  XOR U9810 ( .A(n5670), .B(n5673), .Z(n5740) );
  IV U9811 ( .A(n5672), .Z(n5673) );
  NAND U9812 ( .A(n5741), .B(n5742), .Z(n5672) );
  OR U9813 ( .A(n5743), .B(n5744), .Z(n5742) );
  OR U9814 ( .A(n5745), .B(n5746), .Z(n5741) );
  NAND U9815 ( .A(n5747), .B(n5748), .Z(n5670) );
  OR U9816 ( .A(n5749), .B(n5750), .Z(n5748) );
  OR U9817 ( .A(n5751), .B(n5752), .Z(n5747) );
  NOR U9818 ( .A(n5753), .B(n5754), .Z(n5671) );
  ANDN U9819 ( .B(n5755), .A(n5756), .Z(n5665) );
  IV U9820 ( .A(n5757), .Z(n5755) );
  XNOR U9821 ( .A(n5658), .B(n5758), .Z(n5664) );
  XNOR U9822 ( .A(n5657), .B(n5659), .Z(n5758) );
  NAND U9823 ( .A(n5759), .B(n5760), .Z(n5659) );
  OR U9824 ( .A(n5761), .B(n5762), .Z(n5760) );
  OR U9825 ( .A(n5763), .B(n5764), .Z(n5759) );
  NAND U9826 ( .A(n5765), .B(n5766), .Z(n5657) );
  OR U9827 ( .A(n5767), .B(n5768), .Z(n5766) );
  OR U9828 ( .A(n5769), .B(n5770), .Z(n5765) );
  ANDN U9829 ( .B(n5771), .A(n5772), .Z(n5658) );
  IV U9830 ( .A(n5773), .Z(n5771) );
  XNOR U9831 ( .A(n5738), .B(n5737), .Z(N29681) );
  XOR U9832 ( .A(n5757), .B(n5756), .Z(n5737) );
  XNOR U9833 ( .A(n5772), .B(n5773), .Z(n5756) );
  XNOR U9834 ( .A(n5767), .B(n5768), .Z(n5773) );
  XNOR U9835 ( .A(n5769), .B(n5770), .Z(n5768) );
  XNOR U9836 ( .A(y[3508]), .B(x[3508]), .Z(n5770) );
  XNOR U9837 ( .A(y[3509]), .B(x[3509]), .Z(n5769) );
  XNOR U9838 ( .A(y[3507]), .B(x[3507]), .Z(n5767) );
  XNOR U9839 ( .A(n5761), .B(n5762), .Z(n5772) );
  XNOR U9840 ( .A(y[3504]), .B(x[3504]), .Z(n5762) );
  XNOR U9841 ( .A(n5763), .B(n5764), .Z(n5761) );
  XNOR U9842 ( .A(y[3505]), .B(x[3505]), .Z(n5764) );
  XNOR U9843 ( .A(y[3506]), .B(x[3506]), .Z(n5763) );
  XNOR U9844 ( .A(n5754), .B(n5753), .Z(n5757) );
  XNOR U9845 ( .A(n5749), .B(n5750), .Z(n5753) );
  XNOR U9846 ( .A(y[3501]), .B(x[3501]), .Z(n5750) );
  XNOR U9847 ( .A(n5751), .B(n5752), .Z(n5749) );
  XNOR U9848 ( .A(y[3502]), .B(x[3502]), .Z(n5752) );
  XNOR U9849 ( .A(y[3503]), .B(x[3503]), .Z(n5751) );
  XNOR U9850 ( .A(n5743), .B(n5744), .Z(n5754) );
  XNOR U9851 ( .A(y[3498]), .B(x[3498]), .Z(n5744) );
  XNOR U9852 ( .A(n5745), .B(n5746), .Z(n5743) );
  XNOR U9853 ( .A(y[3499]), .B(x[3499]), .Z(n5746) );
  XNOR U9854 ( .A(y[3500]), .B(x[3500]), .Z(n5745) );
  XOR U9855 ( .A(n5719), .B(n5720), .Z(n5738) );
  XNOR U9856 ( .A(n5735), .B(n5736), .Z(n5720) );
  XNOR U9857 ( .A(n5730), .B(n5731), .Z(n5736) );
  XNOR U9858 ( .A(n5732), .B(n5733), .Z(n5731) );
  XNOR U9859 ( .A(y[3496]), .B(x[3496]), .Z(n5733) );
  XNOR U9860 ( .A(y[3497]), .B(x[3497]), .Z(n5732) );
  XNOR U9861 ( .A(y[3495]), .B(x[3495]), .Z(n5730) );
  XNOR U9862 ( .A(n5724), .B(n5725), .Z(n5735) );
  XNOR U9863 ( .A(y[3492]), .B(x[3492]), .Z(n5725) );
  XNOR U9864 ( .A(n5726), .B(n5727), .Z(n5724) );
  XNOR U9865 ( .A(y[3493]), .B(x[3493]), .Z(n5727) );
  XNOR U9866 ( .A(y[3494]), .B(x[3494]), .Z(n5726) );
  XOR U9867 ( .A(n5718), .B(n5717), .Z(n5719) );
  XNOR U9868 ( .A(n5713), .B(n5714), .Z(n5717) );
  XNOR U9869 ( .A(y[3489]), .B(x[3489]), .Z(n5714) );
  XNOR U9870 ( .A(n5715), .B(n5716), .Z(n5713) );
  XNOR U9871 ( .A(y[3490]), .B(x[3490]), .Z(n5716) );
  XNOR U9872 ( .A(y[3491]), .B(x[3491]), .Z(n5715) );
  XNOR U9873 ( .A(n5707), .B(n5708), .Z(n5718) );
  XNOR U9874 ( .A(y[3486]), .B(x[3486]), .Z(n5708) );
  XNOR U9875 ( .A(n5709), .B(n5710), .Z(n5707) );
  XNOR U9876 ( .A(y[3487]), .B(x[3487]), .Z(n5710) );
  XNOR U9877 ( .A(y[3488]), .B(x[3488]), .Z(n5709) );
  NAND U9878 ( .A(n5774), .B(n5775), .Z(N29673) );
  NANDN U9879 ( .A(n5776), .B(n5777), .Z(n5775) );
  OR U9880 ( .A(n5778), .B(n5779), .Z(n5777) );
  NAND U9881 ( .A(n5778), .B(n5779), .Z(n5774) );
  XOR U9882 ( .A(n5778), .B(n5780), .Z(N29672) );
  XNOR U9883 ( .A(n5776), .B(n5779), .Z(n5780) );
  AND U9884 ( .A(n5781), .B(n5782), .Z(n5779) );
  NANDN U9885 ( .A(n5783), .B(n5784), .Z(n5782) );
  NANDN U9886 ( .A(n5785), .B(n5786), .Z(n5784) );
  NANDN U9887 ( .A(n5786), .B(n5785), .Z(n5781) );
  NAND U9888 ( .A(n5787), .B(n5788), .Z(n5776) );
  NANDN U9889 ( .A(n5789), .B(n5790), .Z(n5788) );
  OR U9890 ( .A(n5791), .B(n5792), .Z(n5790) );
  NAND U9891 ( .A(n5792), .B(n5791), .Z(n5787) );
  AND U9892 ( .A(n5793), .B(n5794), .Z(n5778) );
  NANDN U9893 ( .A(n5795), .B(n5796), .Z(n5794) );
  NANDN U9894 ( .A(n5797), .B(n5798), .Z(n5796) );
  NANDN U9895 ( .A(n5798), .B(n5797), .Z(n5793) );
  XOR U9896 ( .A(n5792), .B(n5799), .Z(N29671) );
  XOR U9897 ( .A(n5789), .B(n5791), .Z(n5799) );
  XNOR U9898 ( .A(n5785), .B(n5800), .Z(n5791) );
  XNOR U9899 ( .A(n5783), .B(n5786), .Z(n5800) );
  NAND U9900 ( .A(n5801), .B(n5802), .Z(n5786) );
  NAND U9901 ( .A(n5803), .B(n5804), .Z(n5802) );
  OR U9902 ( .A(n5805), .B(n5806), .Z(n5803) );
  NANDN U9903 ( .A(n5807), .B(n5805), .Z(n5801) );
  IV U9904 ( .A(n5806), .Z(n5807) );
  NAND U9905 ( .A(n5808), .B(n5809), .Z(n5783) );
  NAND U9906 ( .A(n5810), .B(n5811), .Z(n5809) );
  NANDN U9907 ( .A(n5812), .B(n5813), .Z(n5810) );
  NANDN U9908 ( .A(n5813), .B(n5812), .Z(n5808) );
  AND U9909 ( .A(n5814), .B(n5815), .Z(n5785) );
  NAND U9910 ( .A(n5816), .B(n5817), .Z(n5815) );
  OR U9911 ( .A(n5818), .B(n5819), .Z(n5816) );
  NANDN U9912 ( .A(n5820), .B(n5818), .Z(n5814) );
  NAND U9913 ( .A(n5821), .B(n5822), .Z(n5789) );
  NANDN U9914 ( .A(n5823), .B(n5824), .Z(n5822) );
  OR U9915 ( .A(n5825), .B(n5826), .Z(n5824) );
  NANDN U9916 ( .A(n5827), .B(n5825), .Z(n5821) );
  IV U9917 ( .A(n5826), .Z(n5827) );
  XNOR U9918 ( .A(n5797), .B(n5828), .Z(n5792) );
  XNOR U9919 ( .A(n5795), .B(n5798), .Z(n5828) );
  NAND U9920 ( .A(n5829), .B(n5830), .Z(n5798) );
  NAND U9921 ( .A(n5831), .B(n5832), .Z(n5830) );
  OR U9922 ( .A(n5833), .B(n5834), .Z(n5831) );
  NANDN U9923 ( .A(n5835), .B(n5833), .Z(n5829) );
  IV U9924 ( .A(n5834), .Z(n5835) );
  NAND U9925 ( .A(n5836), .B(n5837), .Z(n5795) );
  NAND U9926 ( .A(n5838), .B(n5839), .Z(n5837) );
  NANDN U9927 ( .A(n5840), .B(n5841), .Z(n5838) );
  NANDN U9928 ( .A(n5841), .B(n5840), .Z(n5836) );
  AND U9929 ( .A(n5842), .B(n5843), .Z(n5797) );
  NAND U9930 ( .A(n5844), .B(n5845), .Z(n5843) );
  OR U9931 ( .A(n5846), .B(n5847), .Z(n5844) );
  NANDN U9932 ( .A(n5848), .B(n5846), .Z(n5842) );
  XNOR U9933 ( .A(n5823), .B(n5849), .Z(N29670) );
  XOR U9934 ( .A(n5825), .B(n5826), .Z(n5849) );
  XNOR U9935 ( .A(n5839), .B(n5850), .Z(n5826) );
  XOR U9936 ( .A(n5840), .B(n5841), .Z(n5850) );
  XOR U9937 ( .A(n5846), .B(n5851), .Z(n5841) );
  XOR U9938 ( .A(n5845), .B(n5848), .Z(n5851) );
  IV U9939 ( .A(n5847), .Z(n5848) );
  NAND U9940 ( .A(n5852), .B(n5853), .Z(n5847) );
  OR U9941 ( .A(n5854), .B(n5855), .Z(n5853) );
  OR U9942 ( .A(n5856), .B(n5857), .Z(n5852) );
  NAND U9943 ( .A(n5858), .B(n5859), .Z(n5845) );
  OR U9944 ( .A(n5860), .B(n5861), .Z(n5859) );
  OR U9945 ( .A(n5862), .B(n5863), .Z(n5858) );
  NOR U9946 ( .A(n5864), .B(n5865), .Z(n5846) );
  ANDN U9947 ( .B(n5866), .A(n5867), .Z(n5840) );
  XNOR U9948 ( .A(n5833), .B(n5868), .Z(n5839) );
  XNOR U9949 ( .A(n5832), .B(n5834), .Z(n5868) );
  NAND U9950 ( .A(n5869), .B(n5870), .Z(n5834) );
  OR U9951 ( .A(n5871), .B(n5872), .Z(n5870) );
  OR U9952 ( .A(n5873), .B(n5874), .Z(n5869) );
  NAND U9953 ( .A(n5875), .B(n5876), .Z(n5832) );
  OR U9954 ( .A(n5877), .B(n5878), .Z(n5876) );
  OR U9955 ( .A(n5879), .B(n5880), .Z(n5875) );
  ANDN U9956 ( .B(n5881), .A(n5882), .Z(n5833) );
  IV U9957 ( .A(n5883), .Z(n5881) );
  ANDN U9958 ( .B(n5884), .A(n5885), .Z(n5825) );
  XOR U9959 ( .A(n5811), .B(n5886), .Z(n5823) );
  XOR U9960 ( .A(n5812), .B(n5813), .Z(n5886) );
  XOR U9961 ( .A(n5818), .B(n5887), .Z(n5813) );
  XOR U9962 ( .A(n5817), .B(n5820), .Z(n5887) );
  IV U9963 ( .A(n5819), .Z(n5820) );
  NAND U9964 ( .A(n5888), .B(n5889), .Z(n5819) );
  OR U9965 ( .A(n5890), .B(n5891), .Z(n5889) );
  OR U9966 ( .A(n5892), .B(n5893), .Z(n5888) );
  NAND U9967 ( .A(n5894), .B(n5895), .Z(n5817) );
  OR U9968 ( .A(n5896), .B(n5897), .Z(n5895) );
  OR U9969 ( .A(n5898), .B(n5899), .Z(n5894) );
  NOR U9970 ( .A(n5900), .B(n5901), .Z(n5818) );
  ANDN U9971 ( .B(n5902), .A(n5903), .Z(n5812) );
  IV U9972 ( .A(n5904), .Z(n5902) );
  XNOR U9973 ( .A(n5805), .B(n5905), .Z(n5811) );
  XNOR U9974 ( .A(n5804), .B(n5806), .Z(n5905) );
  NAND U9975 ( .A(n5906), .B(n5907), .Z(n5806) );
  OR U9976 ( .A(n5908), .B(n5909), .Z(n5907) );
  OR U9977 ( .A(n5910), .B(n5911), .Z(n5906) );
  NAND U9978 ( .A(n5912), .B(n5913), .Z(n5804) );
  OR U9979 ( .A(n5914), .B(n5915), .Z(n5913) );
  OR U9980 ( .A(n5916), .B(n5917), .Z(n5912) );
  ANDN U9981 ( .B(n5918), .A(n5919), .Z(n5805) );
  IV U9982 ( .A(n5920), .Z(n5918) );
  XNOR U9983 ( .A(n5885), .B(n5884), .Z(N29669) );
  XOR U9984 ( .A(n5904), .B(n5903), .Z(n5884) );
  XNOR U9985 ( .A(n5919), .B(n5920), .Z(n5903) );
  XNOR U9986 ( .A(n5914), .B(n5915), .Z(n5920) );
  XNOR U9987 ( .A(n5916), .B(n5917), .Z(n5915) );
  XNOR U9988 ( .A(y[3484]), .B(x[3484]), .Z(n5917) );
  XNOR U9989 ( .A(y[3485]), .B(x[3485]), .Z(n5916) );
  XNOR U9990 ( .A(y[3483]), .B(x[3483]), .Z(n5914) );
  XNOR U9991 ( .A(n5908), .B(n5909), .Z(n5919) );
  XNOR U9992 ( .A(y[3480]), .B(x[3480]), .Z(n5909) );
  XNOR U9993 ( .A(n5910), .B(n5911), .Z(n5908) );
  XNOR U9994 ( .A(y[3481]), .B(x[3481]), .Z(n5911) );
  XNOR U9995 ( .A(y[3482]), .B(x[3482]), .Z(n5910) );
  XNOR U9996 ( .A(n5901), .B(n5900), .Z(n5904) );
  XNOR U9997 ( .A(n5896), .B(n5897), .Z(n5900) );
  XNOR U9998 ( .A(y[3477]), .B(x[3477]), .Z(n5897) );
  XNOR U9999 ( .A(n5898), .B(n5899), .Z(n5896) );
  XNOR U10000 ( .A(y[3478]), .B(x[3478]), .Z(n5899) );
  XNOR U10001 ( .A(y[3479]), .B(x[3479]), .Z(n5898) );
  XNOR U10002 ( .A(n5890), .B(n5891), .Z(n5901) );
  XNOR U10003 ( .A(y[3474]), .B(x[3474]), .Z(n5891) );
  XNOR U10004 ( .A(n5892), .B(n5893), .Z(n5890) );
  XNOR U10005 ( .A(y[3475]), .B(x[3475]), .Z(n5893) );
  XNOR U10006 ( .A(y[3476]), .B(x[3476]), .Z(n5892) );
  XOR U10007 ( .A(n5866), .B(n5867), .Z(n5885) );
  XNOR U10008 ( .A(n5882), .B(n5883), .Z(n5867) );
  XNOR U10009 ( .A(n5877), .B(n5878), .Z(n5883) );
  XNOR U10010 ( .A(n5879), .B(n5880), .Z(n5878) );
  XNOR U10011 ( .A(y[3472]), .B(x[3472]), .Z(n5880) );
  XNOR U10012 ( .A(y[3473]), .B(x[3473]), .Z(n5879) );
  XNOR U10013 ( .A(y[3471]), .B(x[3471]), .Z(n5877) );
  XNOR U10014 ( .A(n5871), .B(n5872), .Z(n5882) );
  XNOR U10015 ( .A(y[3468]), .B(x[3468]), .Z(n5872) );
  XNOR U10016 ( .A(n5873), .B(n5874), .Z(n5871) );
  XNOR U10017 ( .A(y[3469]), .B(x[3469]), .Z(n5874) );
  XNOR U10018 ( .A(y[3470]), .B(x[3470]), .Z(n5873) );
  XOR U10019 ( .A(n5865), .B(n5864), .Z(n5866) );
  XNOR U10020 ( .A(n5860), .B(n5861), .Z(n5864) );
  XNOR U10021 ( .A(y[3465]), .B(x[3465]), .Z(n5861) );
  XNOR U10022 ( .A(n5862), .B(n5863), .Z(n5860) );
  XNOR U10023 ( .A(y[3466]), .B(x[3466]), .Z(n5863) );
  XNOR U10024 ( .A(y[3467]), .B(x[3467]), .Z(n5862) );
  XNOR U10025 ( .A(n5854), .B(n5855), .Z(n5865) );
  XNOR U10026 ( .A(y[3462]), .B(x[3462]), .Z(n5855) );
  XNOR U10027 ( .A(n5856), .B(n5857), .Z(n5854) );
  XNOR U10028 ( .A(y[3463]), .B(x[3463]), .Z(n5857) );
  XNOR U10029 ( .A(y[3464]), .B(x[3464]), .Z(n5856) );
  NAND U10030 ( .A(n5921), .B(n5922), .Z(N29661) );
  NANDN U10031 ( .A(n5923), .B(n5924), .Z(n5922) );
  OR U10032 ( .A(n5925), .B(n5926), .Z(n5924) );
  NAND U10033 ( .A(n5925), .B(n5926), .Z(n5921) );
  XOR U10034 ( .A(n5925), .B(n5927), .Z(N29660) );
  XNOR U10035 ( .A(n5923), .B(n5926), .Z(n5927) );
  AND U10036 ( .A(n5928), .B(n5929), .Z(n5926) );
  NANDN U10037 ( .A(n5930), .B(n5931), .Z(n5929) );
  NANDN U10038 ( .A(n5932), .B(n5933), .Z(n5931) );
  NANDN U10039 ( .A(n5933), .B(n5932), .Z(n5928) );
  NAND U10040 ( .A(n5934), .B(n5935), .Z(n5923) );
  NANDN U10041 ( .A(n5936), .B(n5937), .Z(n5935) );
  OR U10042 ( .A(n5938), .B(n5939), .Z(n5937) );
  NAND U10043 ( .A(n5939), .B(n5938), .Z(n5934) );
  AND U10044 ( .A(n5940), .B(n5941), .Z(n5925) );
  NANDN U10045 ( .A(n5942), .B(n5943), .Z(n5941) );
  NANDN U10046 ( .A(n5944), .B(n5945), .Z(n5943) );
  NANDN U10047 ( .A(n5945), .B(n5944), .Z(n5940) );
  XOR U10048 ( .A(n5939), .B(n5946), .Z(N29659) );
  XOR U10049 ( .A(n5936), .B(n5938), .Z(n5946) );
  XNOR U10050 ( .A(n5932), .B(n5947), .Z(n5938) );
  XNOR U10051 ( .A(n5930), .B(n5933), .Z(n5947) );
  NAND U10052 ( .A(n5948), .B(n5949), .Z(n5933) );
  NAND U10053 ( .A(n5950), .B(n5951), .Z(n5949) );
  OR U10054 ( .A(n5952), .B(n5953), .Z(n5950) );
  NANDN U10055 ( .A(n5954), .B(n5952), .Z(n5948) );
  IV U10056 ( .A(n5953), .Z(n5954) );
  NAND U10057 ( .A(n5955), .B(n5956), .Z(n5930) );
  NAND U10058 ( .A(n5957), .B(n5958), .Z(n5956) );
  NANDN U10059 ( .A(n5959), .B(n5960), .Z(n5957) );
  NANDN U10060 ( .A(n5960), .B(n5959), .Z(n5955) );
  AND U10061 ( .A(n5961), .B(n5962), .Z(n5932) );
  NAND U10062 ( .A(n5963), .B(n5964), .Z(n5962) );
  OR U10063 ( .A(n5965), .B(n5966), .Z(n5963) );
  NANDN U10064 ( .A(n5967), .B(n5965), .Z(n5961) );
  NAND U10065 ( .A(n5968), .B(n5969), .Z(n5936) );
  NANDN U10066 ( .A(n5970), .B(n5971), .Z(n5969) );
  OR U10067 ( .A(n5972), .B(n5973), .Z(n5971) );
  NANDN U10068 ( .A(n5974), .B(n5972), .Z(n5968) );
  IV U10069 ( .A(n5973), .Z(n5974) );
  XNOR U10070 ( .A(n5944), .B(n5975), .Z(n5939) );
  XNOR U10071 ( .A(n5942), .B(n5945), .Z(n5975) );
  NAND U10072 ( .A(n5976), .B(n5977), .Z(n5945) );
  NAND U10073 ( .A(n5978), .B(n5979), .Z(n5977) );
  OR U10074 ( .A(n5980), .B(n5981), .Z(n5978) );
  NANDN U10075 ( .A(n5982), .B(n5980), .Z(n5976) );
  IV U10076 ( .A(n5981), .Z(n5982) );
  NAND U10077 ( .A(n5983), .B(n5984), .Z(n5942) );
  NAND U10078 ( .A(n5985), .B(n5986), .Z(n5984) );
  NANDN U10079 ( .A(n5987), .B(n5988), .Z(n5985) );
  NANDN U10080 ( .A(n5988), .B(n5987), .Z(n5983) );
  AND U10081 ( .A(n5989), .B(n5990), .Z(n5944) );
  NAND U10082 ( .A(n5991), .B(n5992), .Z(n5990) );
  OR U10083 ( .A(n5993), .B(n5994), .Z(n5991) );
  NANDN U10084 ( .A(n5995), .B(n5993), .Z(n5989) );
  XNOR U10085 ( .A(n5970), .B(n5996), .Z(N29658) );
  XOR U10086 ( .A(n5972), .B(n5973), .Z(n5996) );
  XNOR U10087 ( .A(n5986), .B(n5997), .Z(n5973) );
  XOR U10088 ( .A(n5987), .B(n5988), .Z(n5997) );
  XOR U10089 ( .A(n5993), .B(n5998), .Z(n5988) );
  XOR U10090 ( .A(n5992), .B(n5995), .Z(n5998) );
  IV U10091 ( .A(n5994), .Z(n5995) );
  NAND U10092 ( .A(n5999), .B(n6000), .Z(n5994) );
  OR U10093 ( .A(n6001), .B(n6002), .Z(n6000) );
  OR U10094 ( .A(n6003), .B(n6004), .Z(n5999) );
  NAND U10095 ( .A(n6005), .B(n6006), .Z(n5992) );
  OR U10096 ( .A(n6007), .B(n6008), .Z(n6006) );
  OR U10097 ( .A(n6009), .B(n6010), .Z(n6005) );
  NOR U10098 ( .A(n6011), .B(n6012), .Z(n5993) );
  ANDN U10099 ( .B(n6013), .A(n6014), .Z(n5987) );
  XNOR U10100 ( .A(n5980), .B(n6015), .Z(n5986) );
  XNOR U10101 ( .A(n5979), .B(n5981), .Z(n6015) );
  NAND U10102 ( .A(n6016), .B(n6017), .Z(n5981) );
  OR U10103 ( .A(n6018), .B(n6019), .Z(n6017) );
  OR U10104 ( .A(n6020), .B(n6021), .Z(n6016) );
  NAND U10105 ( .A(n6022), .B(n6023), .Z(n5979) );
  OR U10106 ( .A(n6024), .B(n6025), .Z(n6023) );
  OR U10107 ( .A(n6026), .B(n6027), .Z(n6022) );
  ANDN U10108 ( .B(n6028), .A(n6029), .Z(n5980) );
  IV U10109 ( .A(n6030), .Z(n6028) );
  ANDN U10110 ( .B(n6031), .A(n6032), .Z(n5972) );
  XOR U10111 ( .A(n5958), .B(n6033), .Z(n5970) );
  XOR U10112 ( .A(n5959), .B(n5960), .Z(n6033) );
  XOR U10113 ( .A(n5965), .B(n6034), .Z(n5960) );
  XOR U10114 ( .A(n5964), .B(n5967), .Z(n6034) );
  IV U10115 ( .A(n5966), .Z(n5967) );
  NAND U10116 ( .A(n6035), .B(n6036), .Z(n5966) );
  OR U10117 ( .A(n6037), .B(n6038), .Z(n6036) );
  OR U10118 ( .A(n6039), .B(n6040), .Z(n6035) );
  NAND U10119 ( .A(n6041), .B(n6042), .Z(n5964) );
  OR U10120 ( .A(n6043), .B(n6044), .Z(n6042) );
  OR U10121 ( .A(n6045), .B(n6046), .Z(n6041) );
  NOR U10122 ( .A(n6047), .B(n6048), .Z(n5965) );
  ANDN U10123 ( .B(n6049), .A(n6050), .Z(n5959) );
  IV U10124 ( .A(n6051), .Z(n6049) );
  XNOR U10125 ( .A(n5952), .B(n6052), .Z(n5958) );
  XNOR U10126 ( .A(n5951), .B(n5953), .Z(n6052) );
  NAND U10127 ( .A(n6053), .B(n6054), .Z(n5953) );
  OR U10128 ( .A(n6055), .B(n6056), .Z(n6054) );
  OR U10129 ( .A(n6057), .B(n6058), .Z(n6053) );
  NAND U10130 ( .A(n6059), .B(n6060), .Z(n5951) );
  OR U10131 ( .A(n6061), .B(n6062), .Z(n6060) );
  OR U10132 ( .A(n6063), .B(n6064), .Z(n6059) );
  ANDN U10133 ( .B(n6065), .A(n6066), .Z(n5952) );
  IV U10134 ( .A(n6067), .Z(n6065) );
  XNOR U10135 ( .A(n6032), .B(n6031), .Z(N29657) );
  XOR U10136 ( .A(n6051), .B(n6050), .Z(n6031) );
  XNOR U10137 ( .A(n6066), .B(n6067), .Z(n6050) );
  XNOR U10138 ( .A(n6061), .B(n6062), .Z(n6067) );
  XNOR U10139 ( .A(n6063), .B(n6064), .Z(n6062) );
  XNOR U10140 ( .A(y[3460]), .B(x[3460]), .Z(n6064) );
  XNOR U10141 ( .A(y[3461]), .B(x[3461]), .Z(n6063) );
  XNOR U10142 ( .A(y[3459]), .B(x[3459]), .Z(n6061) );
  XNOR U10143 ( .A(n6055), .B(n6056), .Z(n6066) );
  XNOR U10144 ( .A(y[3456]), .B(x[3456]), .Z(n6056) );
  XNOR U10145 ( .A(n6057), .B(n6058), .Z(n6055) );
  XNOR U10146 ( .A(y[3457]), .B(x[3457]), .Z(n6058) );
  XNOR U10147 ( .A(y[3458]), .B(x[3458]), .Z(n6057) );
  XNOR U10148 ( .A(n6048), .B(n6047), .Z(n6051) );
  XNOR U10149 ( .A(n6043), .B(n6044), .Z(n6047) );
  XNOR U10150 ( .A(y[3453]), .B(x[3453]), .Z(n6044) );
  XNOR U10151 ( .A(n6045), .B(n6046), .Z(n6043) );
  XNOR U10152 ( .A(y[3454]), .B(x[3454]), .Z(n6046) );
  XNOR U10153 ( .A(y[3455]), .B(x[3455]), .Z(n6045) );
  XNOR U10154 ( .A(n6037), .B(n6038), .Z(n6048) );
  XNOR U10155 ( .A(y[3450]), .B(x[3450]), .Z(n6038) );
  XNOR U10156 ( .A(n6039), .B(n6040), .Z(n6037) );
  XNOR U10157 ( .A(y[3451]), .B(x[3451]), .Z(n6040) );
  XNOR U10158 ( .A(y[3452]), .B(x[3452]), .Z(n6039) );
  XOR U10159 ( .A(n6013), .B(n6014), .Z(n6032) );
  XNOR U10160 ( .A(n6029), .B(n6030), .Z(n6014) );
  XNOR U10161 ( .A(n6024), .B(n6025), .Z(n6030) );
  XNOR U10162 ( .A(n6026), .B(n6027), .Z(n6025) );
  XNOR U10163 ( .A(y[3448]), .B(x[3448]), .Z(n6027) );
  XNOR U10164 ( .A(y[3449]), .B(x[3449]), .Z(n6026) );
  XNOR U10165 ( .A(y[3447]), .B(x[3447]), .Z(n6024) );
  XNOR U10166 ( .A(n6018), .B(n6019), .Z(n6029) );
  XNOR U10167 ( .A(y[3444]), .B(x[3444]), .Z(n6019) );
  XNOR U10168 ( .A(n6020), .B(n6021), .Z(n6018) );
  XNOR U10169 ( .A(y[3445]), .B(x[3445]), .Z(n6021) );
  XNOR U10170 ( .A(y[3446]), .B(x[3446]), .Z(n6020) );
  XOR U10171 ( .A(n6012), .B(n6011), .Z(n6013) );
  XNOR U10172 ( .A(n6007), .B(n6008), .Z(n6011) );
  XNOR U10173 ( .A(y[3441]), .B(x[3441]), .Z(n6008) );
  XNOR U10174 ( .A(n6009), .B(n6010), .Z(n6007) );
  XNOR U10175 ( .A(y[3442]), .B(x[3442]), .Z(n6010) );
  XNOR U10176 ( .A(y[3443]), .B(x[3443]), .Z(n6009) );
  XNOR U10177 ( .A(n6001), .B(n6002), .Z(n6012) );
  XNOR U10178 ( .A(y[3438]), .B(x[3438]), .Z(n6002) );
  XNOR U10179 ( .A(n6003), .B(n6004), .Z(n6001) );
  XNOR U10180 ( .A(y[3439]), .B(x[3439]), .Z(n6004) );
  XNOR U10181 ( .A(y[3440]), .B(x[3440]), .Z(n6003) );
  NAND U10182 ( .A(n6068), .B(n6069), .Z(N29649) );
  NANDN U10183 ( .A(n6070), .B(n6071), .Z(n6069) );
  OR U10184 ( .A(n6072), .B(n6073), .Z(n6071) );
  NAND U10185 ( .A(n6072), .B(n6073), .Z(n6068) );
  XOR U10186 ( .A(n6072), .B(n6074), .Z(N29648) );
  XNOR U10187 ( .A(n6070), .B(n6073), .Z(n6074) );
  AND U10188 ( .A(n6075), .B(n6076), .Z(n6073) );
  NANDN U10189 ( .A(n6077), .B(n6078), .Z(n6076) );
  NANDN U10190 ( .A(n6079), .B(n6080), .Z(n6078) );
  NANDN U10191 ( .A(n6080), .B(n6079), .Z(n6075) );
  NAND U10192 ( .A(n6081), .B(n6082), .Z(n6070) );
  NANDN U10193 ( .A(n6083), .B(n6084), .Z(n6082) );
  OR U10194 ( .A(n6085), .B(n6086), .Z(n6084) );
  NAND U10195 ( .A(n6086), .B(n6085), .Z(n6081) );
  AND U10196 ( .A(n6087), .B(n6088), .Z(n6072) );
  NANDN U10197 ( .A(n6089), .B(n6090), .Z(n6088) );
  NANDN U10198 ( .A(n6091), .B(n6092), .Z(n6090) );
  NANDN U10199 ( .A(n6092), .B(n6091), .Z(n6087) );
  XOR U10200 ( .A(n6086), .B(n6093), .Z(N29647) );
  XOR U10201 ( .A(n6083), .B(n6085), .Z(n6093) );
  XNOR U10202 ( .A(n6079), .B(n6094), .Z(n6085) );
  XNOR U10203 ( .A(n6077), .B(n6080), .Z(n6094) );
  NAND U10204 ( .A(n6095), .B(n6096), .Z(n6080) );
  NAND U10205 ( .A(n6097), .B(n6098), .Z(n6096) );
  OR U10206 ( .A(n6099), .B(n6100), .Z(n6097) );
  NANDN U10207 ( .A(n6101), .B(n6099), .Z(n6095) );
  IV U10208 ( .A(n6100), .Z(n6101) );
  NAND U10209 ( .A(n6102), .B(n6103), .Z(n6077) );
  NAND U10210 ( .A(n6104), .B(n6105), .Z(n6103) );
  NANDN U10211 ( .A(n6106), .B(n6107), .Z(n6104) );
  NANDN U10212 ( .A(n6107), .B(n6106), .Z(n6102) );
  AND U10213 ( .A(n6108), .B(n6109), .Z(n6079) );
  NAND U10214 ( .A(n6110), .B(n6111), .Z(n6109) );
  OR U10215 ( .A(n6112), .B(n6113), .Z(n6110) );
  NANDN U10216 ( .A(n6114), .B(n6112), .Z(n6108) );
  NAND U10217 ( .A(n6115), .B(n6116), .Z(n6083) );
  NANDN U10218 ( .A(n6117), .B(n6118), .Z(n6116) );
  OR U10219 ( .A(n6119), .B(n6120), .Z(n6118) );
  NANDN U10220 ( .A(n6121), .B(n6119), .Z(n6115) );
  IV U10221 ( .A(n6120), .Z(n6121) );
  XNOR U10222 ( .A(n6091), .B(n6122), .Z(n6086) );
  XNOR U10223 ( .A(n6089), .B(n6092), .Z(n6122) );
  NAND U10224 ( .A(n6123), .B(n6124), .Z(n6092) );
  NAND U10225 ( .A(n6125), .B(n6126), .Z(n6124) );
  OR U10226 ( .A(n6127), .B(n6128), .Z(n6125) );
  NANDN U10227 ( .A(n6129), .B(n6127), .Z(n6123) );
  IV U10228 ( .A(n6128), .Z(n6129) );
  NAND U10229 ( .A(n6130), .B(n6131), .Z(n6089) );
  NAND U10230 ( .A(n6132), .B(n6133), .Z(n6131) );
  NANDN U10231 ( .A(n6134), .B(n6135), .Z(n6132) );
  NANDN U10232 ( .A(n6135), .B(n6134), .Z(n6130) );
  AND U10233 ( .A(n6136), .B(n6137), .Z(n6091) );
  NAND U10234 ( .A(n6138), .B(n6139), .Z(n6137) );
  OR U10235 ( .A(n6140), .B(n6141), .Z(n6138) );
  NANDN U10236 ( .A(n6142), .B(n6140), .Z(n6136) );
  XNOR U10237 ( .A(n6117), .B(n6143), .Z(N29646) );
  XOR U10238 ( .A(n6119), .B(n6120), .Z(n6143) );
  XNOR U10239 ( .A(n6133), .B(n6144), .Z(n6120) );
  XOR U10240 ( .A(n6134), .B(n6135), .Z(n6144) );
  XOR U10241 ( .A(n6140), .B(n6145), .Z(n6135) );
  XOR U10242 ( .A(n6139), .B(n6142), .Z(n6145) );
  IV U10243 ( .A(n6141), .Z(n6142) );
  NAND U10244 ( .A(n6146), .B(n6147), .Z(n6141) );
  OR U10245 ( .A(n6148), .B(n6149), .Z(n6147) );
  OR U10246 ( .A(n6150), .B(n6151), .Z(n6146) );
  NAND U10247 ( .A(n6152), .B(n6153), .Z(n6139) );
  OR U10248 ( .A(n6154), .B(n6155), .Z(n6153) );
  OR U10249 ( .A(n6156), .B(n6157), .Z(n6152) );
  NOR U10250 ( .A(n6158), .B(n6159), .Z(n6140) );
  ANDN U10251 ( .B(n6160), .A(n6161), .Z(n6134) );
  XNOR U10252 ( .A(n6127), .B(n6162), .Z(n6133) );
  XNOR U10253 ( .A(n6126), .B(n6128), .Z(n6162) );
  NAND U10254 ( .A(n6163), .B(n6164), .Z(n6128) );
  OR U10255 ( .A(n6165), .B(n6166), .Z(n6164) );
  OR U10256 ( .A(n6167), .B(n6168), .Z(n6163) );
  NAND U10257 ( .A(n6169), .B(n6170), .Z(n6126) );
  OR U10258 ( .A(n6171), .B(n6172), .Z(n6170) );
  OR U10259 ( .A(n6173), .B(n6174), .Z(n6169) );
  ANDN U10260 ( .B(n6175), .A(n6176), .Z(n6127) );
  IV U10261 ( .A(n6177), .Z(n6175) );
  ANDN U10262 ( .B(n6178), .A(n6179), .Z(n6119) );
  XOR U10263 ( .A(n6105), .B(n6180), .Z(n6117) );
  XOR U10264 ( .A(n6106), .B(n6107), .Z(n6180) );
  XOR U10265 ( .A(n6112), .B(n6181), .Z(n6107) );
  XOR U10266 ( .A(n6111), .B(n6114), .Z(n6181) );
  IV U10267 ( .A(n6113), .Z(n6114) );
  NAND U10268 ( .A(n6182), .B(n6183), .Z(n6113) );
  OR U10269 ( .A(n6184), .B(n6185), .Z(n6183) );
  OR U10270 ( .A(n6186), .B(n6187), .Z(n6182) );
  NAND U10271 ( .A(n6188), .B(n6189), .Z(n6111) );
  OR U10272 ( .A(n6190), .B(n6191), .Z(n6189) );
  OR U10273 ( .A(n6192), .B(n6193), .Z(n6188) );
  NOR U10274 ( .A(n6194), .B(n6195), .Z(n6112) );
  ANDN U10275 ( .B(n6196), .A(n6197), .Z(n6106) );
  IV U10276 ( .A(n6198), .Z(n6196) );
  XNOR U10277 ( .A(n6099), .B(n6199), .Z(n6105) );
  XNOR U10278 ( .A(n6098), .B(n6100), .Z(n6199) );
  NAND U10279 ( .A(n6200), .B(n6201), .Z(n6100) );
  OR U10280 ( .A(n6202), .B(n6203), .Z(n6201) );
  OR U10281 ( .A(n6204), .B(n6205), .Z(n6200) );
  NAND U10282 ( .A(n6206), .B(n6207), .Z(n6098) );
  OR U10283 ( .A(n6208), .B(n6209), .Z(n6207) );
  OR U10284 ( .A(n6210), .B(n6211), .Z(n6206) );
  ANDN U10285 ( .B(n6212), .A(n6213), .Z(n6099) );
  IV U10286 ( .A(n6214), .Z(n6212) );
  XNOR U10287 ( .A(n6179), .B(n6178), .Z(N29645) );
  XOR U10288 ( .A(n6198), .B(n6197), .Z(n6178) );
  XNOR U10289 ( .A(n6213), .B(n6214), .Z(n6197) );
  XNOR U10290 ( .A(n6208), .B(n6209), .Z(n6214) );
  XNOR U10291 ( .A(n6210), .B(n6211), .Z(n6209) );
  XNOR U10292 ( .A(y[3436]), .B(x[3436]), .Z(n6211) );
  XNOR U10293 ( .A(y[3437]), .B(x[3437]), .Z(n6210) );
  XNOR U10294 ( .A(y[3435]), .B(x[3435]), .Z(n6208) );
  XNOR U10295 ( .A(n6202), .B(n6203), .Z(n6213) );
  XNOR U10296 ( .A(y[3432]), .B(x[3432]), .Z(n6203) );
  XNOR U10297 ( .A(n6204), .B(n6205), .Z(n6202) );
  XNOR U10298 ( .A(y[3433]), .B(x[3433]), .Z(n6205) );
  XNOR U10299 ( .A(y[3434]), .B(x[3434]), .Z(n6204) );
  XNOR U10300 ( .A(n6195), .B(n6194), .Z(n6198) );
  XNOR U10301 ( .A(n6190), .B(n6191), .Z(n6194) );
  XNOR U10302 ( .A(y[3429]), .B(x[3429]), .Z(n6191) );
  XNOR U10303 ( .A(n6192), .B(n6193), .Z(n6190) );
  XNOR U10304 ( .A(y[3430]), .B(x[3430]), .Z(n6193) );
  XNOR U10305 ( .A(y[3431]), .B(x[3431]), .Z(n6192) );
  XNOR U10306 ( .A(n6184), .B(n6185), .Z(n6195) );
  XNOR U10307 ( .A(y[3426]), .B(x[3426]), .Z(n6185) );
  XNOR U10308 ( .A(n6186), .B(n6187), .Z(n6184) );
  XNOR U10309 ( .A(y[3427]), .B(x[3427]), .Z(n6187) );
  XNOR U10310 ( .A(y[3428]), .B(x[3428]), .Z(n6186) );
  XOR U10311 ( .A(n6160), .B(n6161), .Z(n6179) );
  XNOR U10312 ( .A(n6176), .B(n6177), .Z(n6161) );
  XNOR U10313 ( .A(n6171), .B(n6172), .Z(n6177) );
  XNOR U10314 ( .A(n6173), .B(n6174), .Z(n6172) );
  XNOR U10315 ( .A(y[3424]), .B(x[3424]), .Z(n6174) );
  XNOR U10316 ( .A(y[3425]), .B(x[3425]), .Z(n6173) );
  XNOR U10317 ( .A(y[3423]), .B(x[3423]), .Z(n6171) );
  XNOR U10318 ( .A(n6165), .B(n6166), .Z(n6176) );
  XNOR U10319 ( .A(y[3420]), .B(x[3420]), .Z(n6166) );
  XNOR U10320 ( .A(n6167), .B(n6168), .Z(n6165) );
  XNOR U10321 ( .A(y[3421]), .B(x[3421]), .Z(n6168) );
  XNOR U10322 ( .A(y[3422]), .B(x[3422]), .Z(n6167) );
  XOR U10323 ( .A(n6159), .B(n6158), .Z(n6160) );
  XNOR U10324 ( .A(n6154), .B(n6155), .Z(n6158) );
  XNOR U10325 ( .A(y[3417]), .B(x[3417]), .Z(n6155) );
  XNOR U10326 ( .A(n6156), .B(n6157), .Z(n6154) );
  XNOR U10327 ( .A(y[3418]), .B(x[3418]), .Z(n6157) );
  XNOR U10328 ( .A(y[3419]), .B(x[3419]), .Z(n6156) );
  XNOR U10329 ( .A(n6148), .B(n6149), .Z(n6159) );
  XNOR U10330 ( .A(y[3414]), .B(x[3414]), .Z(n6149) );
  XNOR U10331 ( .A(n6150), .B(n6151), .Z(n6148) );
  XNOR U10332 ( .A(y[3415]), .B(x[3415]), .Z(n6151) );
  XNOR U10333 ( .A(y[3416]), .B(x[3416]), .Z(n6150) );
  NAND U10334 ( .A(n6215), .B(n6216), .Z(N29637) );
  NANDN U10335 ( .A(n6217), .B(n6218), .Z(n6216) );
  OR U10336 ( .A(n6219), .B(n6220), .Z(n6218) );
  NAND U10337 ( .A(n6219), .B(n6220), .Z(n6215) );
  XOR U10338 ( .A(n6219), .B(n6221), .Z(N29636) );
  XNOR U10339 ( .A(n6217), .B(n6220), .Z(n6221) );
  AND U10340 ( .A(n6222), .B(n6223), .Z(n6220) );
  NANDN U10341 ( .A(n6224), .B(n6225), .Z(n6223) );
  NANDN U10342 ( .A(n6226), .B(n6227), .Z(n6225) );
  NANDN U10343 ( .A(n6227), .B(n6226), .Z(n6222) );
  NAND U10344 ( .A(n6228), .B(n6229), .Z(n6217) );
  NANDN U10345 ( .A(n6230), .B(n6231), .Z(n6229) );
  OR U10346 ( .A(n6232), .B(n6233), .Z(n6231) );
  NAND U10347 ( .A(n6233), .B(n6232), .Z(n6228) );
  AND U10348 ( .A(n6234), .B(n6235), .Z(n6219) );
  NANDN U10349 ( .A(n6236), .B(n6237), .Z(n6235) );
  NANDN U10350 ( .A(n6238), .B(n6239), .Z(n6237) );
  NANDN U10351 ( .A(n6239), .B(n6238), .Z(n6234) );
  XOR U10352 ( .A(n6233), .B(n6240), .Z(N29635) );
  XOR U10353 ( .A(n6230), .B(n6232), .Z(n6240) );
  XNOR U10354 ( .A(n6226), .B(n6241), .Z(n6232) );
  XNOR U10355 ( .A(n6224), .B(n6227), .Z(n6241) );
  NAND U10356 ( .A(n6242), .B(n6243), .Z(n6227) );
  NAND U10357 ( .A(n6244), .B(n6245), .Z(n6243) );
  OR U10358 ( .A(n6246), .B(n6247), .Z(n6244) );
  NANDN U10359 ( .A(n6248), .B(n6246), .Z(n6242) );
  IV U10360 ( .A(n6247), .Z(n6248) );
  NAND U10361 ( .A(n6249), .B(n6250), .Z(n6224) );
  NAND U10362 ( .A(n6251), .B(n6252), .Z(n6250) );
  NANDN U10363 ( .A(n6253), .B(n6254), .Z(n6251) );
  NANDN U10364 ( .A(n6254), .B(n6253), .Z(n6249) );
  AND U10365 ( .A(n6255), .B(n6256), .Z(n6226) );
  NAND U10366 ( .A(n6257), .B(n6258), .Z(n6256) );
  OR U10367 ( .A(n6259), .B(n6260), .Z(n6257) );
  NANDN U10368 ( .A(n6261), .B(n6259), .Z(n6255) );
  NAND U10369 ( .A(n6262), .B(n6263), .Z(n6230) );
  NANDN U10370 ( .A(n6264), .B(n6265), .Z(n6263) );
  OR U10371 ( .A(n6266), .B(n6267), .Z(n6265) );
  NANDN U10372 ( .A(n6268), .B(n6266), .Z(n6262) );
  IV U10373 ( .A(n6267), .Z(n6268) );
  XNOR U10374 ( .A(n6238), .B(n6269), .Z(n6233) );
  XNOR U10375 ( .A(n6236), .B(n6239), .Z(n6269) );
  NAND U10376 ( .A(n6270), .B(n6271), .Z(n6239) );
  NAND U10377 ( .A(n6272), .B(n6273), .Z(n6271) );
  OR U10378 ( .A(n6274), .B(n6275), .Z(n6272) );
  NANDN U10379 ( .A(n6276), .B(n6274), .Z(n6270) );
  IV U10380 ( .A(n6275), .Z(n6276) );
  NAND U10381 ( .A(n6277), .B(n6278), .Z(n6236) );
  NAND U10382 ( .A(n6279), .B(n6280), .Z(n6278) );
  NANDN U10383 ( .A(n6281), .B(n6282), .Z(n6279) );
  NANDN U10384 ( .A(n6282), .B(n6281), .Z(n6277) );
  AND U10385 ( .A(n6283), .B(n6284), .Z(n6238) );
  NAND U10386 ( .A(n6285), .B(n6286), .Z(n6284) );
  OR U10387 ( .A(n6287), .B(n6288), .Z(n6285) );
  NANDN U10388 ( .A(n6289), .B(n6287), .Z(n6283) );
  XNOR U10389 ( .A(n6264), .B(n6290), .Z(N29634) );
  XOR U10390 ( .A(n6266), .B(n6267), .Z(n6290) );
  XNOR U10391 ( .A(n6280), .B(n6291), .Z(n6267) );
  XOR U10392 ( .A(n6281), .B(n6282), .Z(n6291) );
  XOR U10393 ( .A(n6287), .B(n6292), .Z(n6282) );
  XOR U10394 ( .A(n6286), .B(n6289), .Z(n6292) );
  IV U10395 ( .A(n6288), .Z(n6289) );
  NAND U10396 ( .A(n6293), .B(n6294), .Z(n6288) );
  OR U10397 ( .A(n6295), .B(n6296), .Z(n6294) );
  OR U10398 ( .A(n6297), .B(n6298), .Z(n6293) );
  NAND U10399 ( .A(n6299), .B(n6300), .Z(n6286) );
  OR U10400 ( .A(n6301), .B(n6302), .Z(n6300) );
  OR U10401 ( .A(n6303), .B(n6304), .Z(n6299) );
  NOR U10402 ( .A(n6305), .B(n6306), .Z(n6287) );
  ANDN U10403 ( .B(n6307), .A(n6308), .Z(n6281) );
  XNOR U10404 ( .A(n6274), .B(n6309), .Z(n6280) );
  XNOR U10405 ( .A(n6273), .B(n6275), .Z(n6309) );
  NAND U10406 ( .A(n6310), .B(n6311), .Z(n6275) );
  OR U10407 ( .A(n6312), .B(n6313), .Z(n6311) );
  OR U10408 ( .A(n6314), .B(n6315), .Z(n6310) );
  NAND U10409 ( .A(n6316), .B(n6317), .Z(n6273) );
  OR U10410 ( .A(n6318), .B(n6319), .Z(n6317) );
  OR U10411 ( .A(n6320), .B(n6321), .Z(n6316) );
  ANDN U10412 ( .B(n6322), .A(n6323), .Z(n6274) );
  IV U10413 ( .A(n6324), .Z(n6322) );
  ANDN U10414 ( .B(n6325), .A(n6326), .Z(n6266) );
  XOR U10415 ( .A(n6252), .B(n6327), .Z(n6264) );
  XOR U10416 ( .A(n6253), .B(n6254), .Z(n6327) );
  XOR U10417 ( .A(n6259), .B(n6328), .Z(n6254) );
  XOR U10418 ( .A(n6258), .B(n6261), .Z(n6328) );
  IV U10419 ( .A(n6260), .Z(n6261) );
  NAND U10420 ( .A(n6329), .B(n6330), .Z(n6260) );
  OR U10421 ( .A(n6331), .B(n6332), .Z(n6330) );
  OR U10422 ( .A(n6333), .B(n6334), .Z(n6329) );
  NAND U10423 ( .A(n6335), .B(n6336), .Z(n6258) );
  OR U10424 ( .A(n6337), .B(n6338), .Z(n6336) );
  OR U10425 ( .A(n6339), .B(n6340), .Z(n6335) );
  NOR U10426 ( .A(n6341), .B(n6342), .Z(n6259) );
  ANDN U10427 ( .B(n6343), .A(n6344), .Z(n6253) );
  IV U10428 ( .A(n6345), .Z(n6343) );
  XNOR U10429 ( .A(n6246), .B(n6346), .Z(n6252) );
  XNOR U10430 ( .A(n6245), .B(n6247), .Z(n6346) );
  NAND U10431 ( .A(n6347), .B(n6348), .Z(n6247) );
  OR U10432 ( .A(n6349), .B(n6350), .Z(n6348) );
  OR U10433 ( .A(n6351), .B(n6352), .Z(n6347) );
  NAND U10434 ( .A(n6353), .B(n6354), .Z(n6245) );
  OR U10435 ( .A(n6355), .B(n6356), .Z(n6354) );
  OR U10436 ( .A(n6357), .B(n6358), .Z(n6353) );
  ANDN U10437 ( .B(n6359), .A(n6360), .Z(n6246) );
  IV U10438 ( .A(n6361), .Z(n6359) );
  XNOR U10439 ( .A(n6326), .B(n6325), .Z(N29633) );
  XOR U10440 ( .A(n6345), .B(n6344), .Z(n6325) );
  XNOR U10441 ( .A(n6360), .B(n6361), .Z(n6344) );
  XNOR U10442 ( .A(n6355), .B(n6356), .Z(n6361) );
  XNOR U10443 ( .A(n6357), .B(n6358), .Z(n6356) );
  XNOR U10444 ( .A(y[3412]), .B(x[3412]), .Z(n6358) );
  XNOR U10445 ( .A(y[3413]), .B(x[3413]), .Z(n6357) );
  XNOR U10446 ( .A(y[3411]), .B(x[3411]), .Z(n6355) );
  XNOR U10447 ( .A(n6349), .B(n6350), .Z(n6360) );
  XNOR U10448 ( .A(y[3408]), .B(x[3408]), .Z(n6350) );
  XNOR U10449 ( .A(n6351), .B(n6352), .Z(n6349) );
  XNOR U10450 ( .A(y[3409]), .B(x[3409]), .Z(n6352) );
  XNOR U10451 ( .A(y[3410]), .B(x[3410]), .Z(n6351) );
  XNOR U10452 ( .A(n6342), .B(n6341), .Z(n6345) );
  XNOR U10453 ( .A(n6337), .B(n6338), .Z(n6341) );
  XNOR U10454 ( .A(y[3405]), .B(x[3405]), .Z(n6338) );
  XNOR U10455 ( .A(n6339), .B(n6340), .Z(n6337) );
  XNOR U10456 ( .A(y[3406]), .B(x[3406]), .Z(n6340) );
  XNOR U10457 ( .A(y[3407]), .B(x[3407]), .Z(n6339) );
  XNOR U10458 ( .A(n6331), .B(n6332), .Z(n6342) );
  XNOR U10459 ( .A(y[3402]), .B(x[3402]), .Z(n6332) );
  XNOR U10460 ( .A(n6333), .B(n6334), .Z(n6331) );
  XNOR U10461 ( .A(y[3403]), .B(x[3403]), .Z(n6334) );
  XNOR U10462 ( .A(y[3404]), .B(x[3404]), .Z(n6333) );
  XOR U10463 ( .A(n6307), .B(n6308), .Z(n6326) );
  XNOR U10464 ( .A(n6323), .B(n6324), .Z(n6308) );
  XNOR U10465 ( .A(n6318), .B(n6319), .Z(n6324) );
  XNOR U10466 ( .A(n6320), .B(n6321), .Z(n6319) );
  XNOR U10467 ( .A(y[3400]), .B(x[3400]), .Z(n6321) );
  XNOR U10468 ( .A(y[3401]), .B(x[3401]), .Z(n6320) );
  XNOR U10469 ( .A(y[3399]), .B(x[3399]), .Z(n6318) );
  XNOR U10470 ( .A(n6312), .B(n6313), .Z(n6323) );
  XNOR U10471 ( .A(y[3396]), .B(x[3396]), .Z(n6313) );
  XNOR U10472 ( .A(n6314), .B(n6315), .Z(n6312) );
  XNOR U10473 ( .A(y[3397]), .B(x[3397]), .Z(n6315) );
  XNOR U10474 ( .A(y[3398]), .B(x[3398]), .Z(n6314) );
  XOR U10475 ( .A(n6306), .B(n6305), .Z(n6307) );
  XNOR U10476 ( .A(n6301), .B(n6302), .Z(n6305) );
  XNOR U10477 ( .A(y[3393]), .B(x[3393]), .Z(n6302) );
  XNOR U10478 ( .A(n6303), .B(n6304), .Z(n6301) );
  XNOR U10479 ( .A(y[3394]), .B(x[3394]), .Z(n6304) );
  XNOR U10480 ( .A(y[3395]), .B(x[3395]), .Z(n6303) );
  XNOR U10481 ( .A(n6295), .B(n6296), .Z(n6306) );
  XNOR U10482 ( .A(y[3390]), .B(x[3390]), .Z(n6296) );
  XNOR U10483 ( .A(n6297), .B(n6298), .Z(n6295) );
  XNOR U10484 ( .A(y[3391]), .B(x[3391]), .Z(n6298) );
  XNOR U10485 ( .A(y[3392]), .B(x[3392]), .Z(n6297) );
  NAND U10486 ( .A(n6362), .B(n6363), .Z(N29625) );
  NANDN U10487 ( .A(n6364), .B(n6365), .Z(n6363) );
  OR U10488 ( .A(n6366), .B(n6367), .Z(n6365) );
  NAND U10489 ( .A(n6366), .B(n6367), .Z(n6362) );
  XOR U10490 ( .A(n6366), .B(n6368), .Z(N29624) );
  XNOR U10491 ( .A(n6364), .B(n6367), .Z(n6368) );
  AND U10492 ( .A(n6369), .B(n6370), .Z(n6367) );
  NANDN U10493 ( .A(n6371), .B(n6372), .Z(n6370) );
  NANDN U10494 ( .A(n6373), .B(n6374), .Z(n6372) );
  NANDN U10495 ( .A(n6374), .B(n6373), .Z(n6369) );
  NAND U10496 ( .A(n6375), .B(n6376), .Z(n6364) );
  NANDN U10497 ( .A(n6377), .B(n6378), .Z(n6376) );
  OR U10498 ( .A(n6379), .B(n6380), .Z(n6378) );
  NAND U10499 ( .A(n6380), .B(n6379), .Z(n6375) );
  AND U10500 ( .A(n6381), .B(n6382), .Z(n6366) );
  NANDN U10501 ( .A(n6383), .B(n6384), .Z(n6382) );
  NANDN U10502 ( .A(n6385), .B(n6386), .Z(n6384) );
  NANDN U10503 ( .A(n6386), .B(n6385), .Z(n6381) );
  XOR U10504 ( .A(n6380), .B(n6387), .Z(N29623) );
  XOR U10505 ( .A(n6377), .B(n6379), .Z(n6387) );
  XNOR U10506 ( .A(n6373), .B(n6388), .Z(n6379) );
  XNOR U10507 ( .A(n6371), .B(n6374), .Z(n6388) );
  NAND U10508 ( .A(n6389), .B(n6390), .Z(n6374) );
  NAND U10509 ( .A(n6391), .B(n6392), .Z(n6390) );
  OR U10510 ( .A(n6393), .B(n6394), .Z(n6391) );
  NANDN U10511 ( .A(n6395), .B(n6393), .Z(n6389) );
  IV U10512 ( .A(n6394), .Z(n6395) );
  NAND U10513 ( .A(n6396), .B(n6397), .Z(n6371) );
  NAND U10514 ( .A(n6398), .B(n6399), .Z(n6397) );
  NANDN U10515 ( .A(n6400), .B(n6401), .Z(n6398) );
  NANDN U10516 ( .A(n6401), .B(n6400), .Z(n6396) );
  AND U10517 ( .A(n6402), .B(n6403), .Z(n6373) );
  NAND U10518 ( .A(n6404), .B(n6405), .Z(n6403) );
  OR U10519 ( .A(n6406), .B(n6407), .Z(n6404) );
  NANDN U10520 ( .A(n6408), .B(n6406), .Z(n6402) );
  NAND U10521 ( .A(n6409), .B(n6410), .Z(n6377) );
  NANDN U10522 ( .A(n6411), .B(n6412), .Z(n6410) );
  OR U10523 ( .A(n6413), .B(n6414), .Z(n6412) );
  NANDN U10524 ( .A(n6415), .B(n6413), .Z(n6409) );
  IV U10525 ( .A(n6414), .Z(n6415) );
  XNOR U10526 ( .A(n6385), .B(n6416), .Z(n6380) );
  XNOR U10527 ( .A(n6383), .B(n6386), .Z(n6416) );
  NAND U10528 ( .A(n6417), .B(n6418), .Z(n6386) );
  NAND U10529 ( .A(n6419), .B(n6420), .Z(n6418) );
  OR U10530 ( .A(n6421), .B(n6422), .Z(n6419) );
  NANDN U10531 ( .A(n6423), .B(n6421), .Z(n6417) );
  IV U10532 ( .A(n6422), .Z(n6423) );
  NAND U10533 ( .A(n6424), .B(n6425), .Z(n6383) );
  NAND U10534 ( .A(n6426), .B(n6427), .Z(n6425) );
  NANDN U10535 ( .A(n6428), .B(n6429), .Z(n6426) );
  NANDN U10536 ( .A(n6429), .B(n6428), .Z(n6424) );
  AND U10537 ( .A(n6430), .B(n6431), .Z(n6385) );
  NAND U10538 ( .A(n6432), .B(n6433), .Z(n6431) );
  OR U10539 ( .A(n6434), .B(n6435), .Z(n6432) );
  NANDN U10540 ( .A(n6436), .B(n6434), .Z(n6430) );
  XNOR U10541 ( .A(n6411), .B(n6437), .Z(N29622) );
  XOR U10542 ( .A(n6413), .B(n6414), .Z(n6437) );
  XNOR U10543 ( .A(n6427), .B(n6438), .Z(n6414) );
  XOR U10544 ( .A(n6428), .B(n6429), .Z(n6438) );
  XOR U10545 ( .A(n6434), .B(n6439), .Z(n6429) );
  XOR U10546 ( .A(n6433), .B(n6436), .Z(n6439) );
  IV U10547 ( .A(n6435), .Z(n6436) );
  NAND U10548 ( .A(n6440), .B(n6441), .Z(n6435) );
  OR U10549 ( .A(n6442), .B(n6443), .Z(n6441) );
  OR U10550 ( .A(n6444), .B(n6445), .Z(n6440) );
  NAND U10551 ( .A(n6446), .B(n6447), .Z(n6433) );
  OR U10552 ( .A(n6448), .B(n6449), .Z(n6447) );
  OR U10553 ( .A(n6450), .B(n6451), .Z(n6446) );
  NOR U10554 ( .A(n6452), .B(n6453), .Z(n6434) );
  ANDN U10555 ( .B(n6454), .A(n6455), .Z(n6428) );
  XNOR U10556 ( .A(n6421), .B(n6456), .Z(n6427) );
  XNOR U10557 ( .A(n6420), .B(n6422), .Z(n6456) );
  NAND U10558 ( .A(n6457), .B(n6458), .Z(n6422) );
  OR U10559 ( .A(n6459), .B(n6460), .Z(n6458) );
  OR U10560 ( .A(n6461), .B(n6462), .Z(n6457) );
  NAND U10561 ( .A(n6463), .B(n6464), .Z(n6420) );
  OR U10562 ( .A(n6465), .B(n6466), .Z(n6464) );
  OR U10563 ( .A(n6467), .B(n6468), .Z(n6463) );
  ANDN U10564 ( .B(n6469), .A(n6470), .Z(n6421) );
  IV U10565 ( .A(n6471), .Z(n6469) );
  ANDN U10566 ( .B(n6472), .A(n6473), .Z(n6413) );
  XOR U10567 ( .A(n6399), .B(n6474), .Z(n6411) );
  XOR U10568 ( .A(n6400), .B(n6401), .Z(n6474) );
  XOR U10569 ( .A(n6406), .B(n6475), .Z(n6401) );
  XOR U10570 ( .A(n6405), .B(n6408), .Z(n6475) );
  IV U10571 ( .A(n6407), .Z(n6408) );
  NAND U10572 ( .A(n6476), .B(n6477), .Z(n6407) );
  OR U10573 ( .A(n6478), .B(n6479), .Z(n6477) );
  OR U10574 ( .A(n6480), .B(n6481), .Z(n6476) );
  NAND U10575 ( .A(n6482), .B(n6483), .Z(n6405) );
  OR U10576 ( .A(n6484), .B(n6485), .Z(n6483) );
  OR U10577 ( .A(n6486), .B(n6487), .Z(n6482) );
  NOR U10578 ( .A(n6488), .B(n6489), .Z(n6406) );
  ANDN U10579 ( .B(n6490), .A(n6491), .Z(n6400) );
  IV U10580 ( .A(n6492), .Z(n6490) );
  XNOR U10581 ( .A(n6393), .B(n6493), .Z(n6399) );
  XNOR U10582 ( .A(n6392), .B(n6394), .Z(n6493) );
  NAND U10583 ( .A(n6494), .B(n6495), .Z(n6394) );
  OR U10584 ( .A(n6496), .B(n6497), .Z(n6495) );
  OR U10585 ( .A(n6498), .B(n6499), .Z(n6494) );
  NAND U10586 ( .A(n6500), .B(n6501), .Z(n6392) );
  OR U10587 ( .A(n6502), .B(n6503), .Z(n6501) );
  OR U10588 ( .A(n6504), .B(n6505), .Z(n6500) );
  ANDN U10589 ( .B(n6506), .A(n6507), .Z(n6393) );
  IV U10590 ( .A(n6508), .Z(n6506) );
  XNOR U10591 ( .A(n6473), .B(n6472), .Z(N29621) );
  XOR U10592 ( .A(n6492), .B(n6491), .Z(n6472) );
  XNOR U10593 ( .A(n6507), .B(n6508), .Z(n6491) );
  XNOR U10594 ( .A(n6502), .B(n6503), .Z(n6508) );
  XNOR U10595 ( .A(n6504), .B(n6505), .Z(n6503) );
  XNOR U10596 ( .A(y[3388]), .B(x[3388]), .Z(n6505) );
  XNOR U10597 ( .A(y[3389]), .B(x[3389]), .Z(n6504) );
  XNOR U10598 ( .A(y[3387]), .B(x[3387]), .Z(n6502) );
  XNOR U10599 ( .A(n6496), .B(n6497), .Z(n6507) );
  XNOR U10600 ( .A(y[3384]), .B(x[3384]), .Z(n6497) );
  XNOR U10601 ( .A(n6498), .B(n6499), .Z(n6496) );
  XNOR U10602 ( .A(y[3385]), .B(x[3385]), .Z(n6499) );
  XNOR U10603 ( .A(y[3386]), .B(x[3386]), .Z(n6498) );
  XNOR U10604 ( .A(n6489), .B(n6488), .Z(n6492) );
  XNOR U10605 ( .A(n6484), .B(n6485), .Z(n6488) );
  XNOR U10606 ( .A(y[3381]), .B(x[3381]), .Z(n6485) );
  XNOR U10607 ( .A(n6486), .B(n6487), .Z(n6484) );
  XNOR U10608 ( .A(y[3382]), .B(x[3382]), .Z(n6487) );
  XNOR U10609 ( .A(y[3383]), .B(x[3383]), .Z(n6486) );
  XNOR U10610 ( .A(n6478), .B(n6479), .Z(n6489) );
  XNOR U10611 ( .A(y[3378]), .B(x[3378]), .Z(n6479) );
  XNOR U10612 ( .A(n6480), .B(n6481), .Z(n6478) );
  XNOR U10613 ( .A(y[3379]), .B(x[3379]), .Z(n6481) );
  XNOR U10614 ( .A(y[3380]), .B(x[3380]), .Z(n6480) );
  XOR U10615 ( .A(n6454), .B(n6455), .Z(n6473) );
  XNOR U10616 ( .A(n6470), .B(n6471), .Z(n6455) );
  XNOR U10617 ( .A(n6465), .B(n6466), .Z(n6471) );
  XNOR U10618 ( .A(n6467), .B(n6468), .Z(n6466) );
  XNOR U10619 ( .A(y[3376]), .B(x[3376]), .Z(n6468) );
  XNOR U10620 ( .A(y[3377]), .B(x[3377]), .Z(n6467) );
  XNOR U10621 ( .A(y[3375]), .B(x[3375]), .Z(n6465) );
  XNOR U10622 ( .A(n6459), .B(n6460), .Z(n6470) );
  XNOR U10623 ( .A(y[3372]), .B(x[3372]), .Z(n6460) );
  XNOR U10624 ( .A(n6461), .B(n6462), .Z(n6459) );
  XNOR U10625 ( .A(y[3373]), .B(x[3373]), .Z(n6462) );
  XNOR U10626 ( .A(y[3374]), .B(x[3374]), .Z(n6461) );
  XOR U10627 ( .A(n6453), .B(n6452), .Z(n6454) );
  XNOR U10628 ( .A(n6448), .B(n6449), .Z(n6452) );
  XNOR U10629 ( .A(y[3369]), .B(x[3369]), .Z(n6449) );
  XNOR U10630 ( .A(n6450), .B(n6451), .Z(n6448) );
  XNOR U10631 ( .A(y[3370]), .B(x[3370]), .Z(n6451) );
  XNOR U10632 ( .A(y[3371]), .B(x[3371]), .Z(n6450) );
  XNOR U10633 ( .A(n6442), .B(n6443), .Z(n6453) );
  XNOR U10634 ( .A(y[3366]), .B(x[3366]), .Z(n6443) );
  XNOR U10635 ( .A(n6444), .B(n6445), .Z(n6442) );
  XNOR U10636 ( .A(y[3367]), .B(x[3367]), .Z(n6445) );
  XNOR U10637 ( .A(y[3368]), .B(x[3368]), .Z(n6444) );
  NAND U10638 ( .A(n6509), .B(n6510), .Z(N29613) );
  NANDN U10639 ( .A(n6511), .B(n6512), .Z(n6510) );
  OR U10640 ( .A(n6513), .B(n6514), .Z(n6512) );
  NAND U10641 ( .A(n6513), .B(n6514), .Z(n6509) );
  XOR U10642 ( .A(n6513), .B(n6515), .Z(N29612) );
  XNOR U10643 ( .A(n6511), .B(n6514), .Z(n6515) );
  AND U10644 ( .A(n6516), .B(n6517), .Z(n6514) );
  NANDN U10645 ( .A(n6518), .B(n6519), .Z(n6517) );
  NANDN U10646 ( .A(n6520), .B(n6521), .Z(n6519) );
  NANDN U10647 ( .A(n6521), .B(n6520), .Z(n6516) );
  NAND U10648 ( .A(n6522), .B(n6523), .Z(n6511) );
  NANDN U10649 ( .A(n6524), .B(n6525), .Z(n6523) );
  OR U10650 ( .A(n6526), .B(n6527), .Z(n6525) );
  NAND U10651 ( .A(n6527), .B(n6526), .Z(n6522) );
  AND U10652 ( .A(n6528), .B(n6529), .Z(n6513) );
  NANDN U10653 ( .A(n6530), .B(n6531), .Z(n6529) );
  NANDN U10654 ( .A(n6532), .B(n6533), .Z(n6531) );
  NANDN U10655 ( .A(n6533), .B(n6532), .Z(n6528) );
  XOR U10656 ( .A(n6527), .B(n6534), .Z(N29611) );
  XOR U10657 ( .A(n6524), .B(n6526), .Z(n6534) );
  XNOR U10658 ( .A(n6520), .B(n6535), .Z(n6526) );
  XNOR U10659 ( .A(n6518), .B(n6521), .Z(n6535) );
  NAND U10660 ( .A(n6536), .B(n6537), .Z(n6521) );
  NAND U10661 ( .A(n6538), .B(n6539), .Z(n6537) );
  OR U10662 ( .A(n6540), .B(n6541), .Z(n6538) );
  NANDN U10663 ( .A(n6542), .B(n6540), .Z(n6536) );
  IV U10664 ( .A(n6541), .Z(n6542) );
  NAND U10665 ( .A(n6543), .B(n6544), .Z(n6518) );
  NAND U10666 ( .A(n6545), .B(n6546), .Z(n6544) );
  NANDN U10667 ( .A(n6547), .B(n6548), .Z(n6545) );
  NANDN U10668 ( .A(n6548), .B(n6547), .Z(n6543) );
  AND U10669 ( .A(n6549), .B(n6550), .Z(n6520) );
  NAND U10670 ( .A(n6551), .B(n6552), .Z(n6550) );
  OR U10671 ( .A(n6553), .B(n6554), .Z(n6551) );
  NANDN U10672 ( .A(n6555), .B(n6553), .Z(n6549) );
  NAND U10673 ( .A(n6556), .B(n6557), .Z(n6524) );
  NANDN U10674 ( .A(n6558), .B(n6559), .Z(n6557) );
  OR U10675 ( .A(n6560), .B(n6561), .Z(n6559) );
  NANDN U10676 ( .A(n6562), .B(n6560), .Z(n6556) );
  IV U10677 ( .A(n6561), .Z(n6562) );
  XNOR U10678 ( .A(n6532), .B(n6563), .Z(n6527) );
  XNOR U10679 ( .A(n6530), .B(n6533), .Z(n6563) );
  NAND U10680 ( .A(n6564), .B(n6565), .Z(n6533) );
  NAND U10681 ( .A(n6566), .B(n6567), .Z(n6565) );
  OR U10682 ( .A(n6568), .B(n6569), .Z(n6566) );
  NANDN U10683 ( .A(n6570), .B(n6568), .Z(n6564) );
  IV U10684 ( .A(n6569), .Z(n6570) );
  NAND U10685 ( .A(n6571), .B(n6572), .Z(n6530) );
  NAND U10686 ( .A(n6573), .B(n6574), .Z(n6572) );
  NANDN U10687 ( .A(n6575), .B(n6576), .Z(n6573) );
  NANDN U10688 ( .A(n6576), .B(n6575), .Z(n6571) );
  AND U10689 ( .A(n6577), .B(n6578), .Z(n6532) );
  NAND U10690 ( .A(n6579), .B(n6580), .Z(n6578) );
  OR U10691 ( .A(n6581), .B(n6582), .Z(n6579) );
  NANDN U10692 ( .A(n6583), .B(n6581), .Z(n6577) );
  XNOR U10693 ( .A(n6558), .B(n6584), .Z(N29610) );
  XOR U10694 ( .A(n6560), .B(n6561), .Z(n6584) );
  XNOR U10695 ( .A(n6574), .B(n6585), .Z(n6561) );
  XOR U10696 ( .A(n6575), .B(n6576), .Z(n6585) );
  XOR U10697 ( .A(n6581), .B(n6586), .Z(n6576) );
  XOR U10698 ( .A(n6580), .B(n6583), .Z(n6586) );
  IV U10699 ( .A(n6582), .Z(n6583) );
  NAND U10700 ( .A(n6587), .B(n6588), .Z(n6582) );
  OR U10701 ( .A(n6589), .B(n6590), .Z(n6588) );
  OR U10702 ( .A(n6591), .B(n6592), .Z(n6587) );
  NAND U10703 ( .A(n6593), .B(n6594), .Z(n6580) );
  OR U10704 ( .A(n6595), .B(n6596), .Z(n6594) );
  OR U10705 ( .A(n6597), .B(n6598), .Z(n6593) );
  NOR U10706 ( .A(n6599), .B(n6600), .Z(n6581) );
  ANDN U10707 ( .B(n6601), .A(n6602), .Z(n6575) );
  XNOR U10708 ( .A(n6568), .B(n6603), .Z(n6574) );
  XNOR U10709 ( .A(n6567), .B(n6569), .Z(n6603) );
  NAND U10710 ( .A(n6604), .B(n6605), .Z(n6569) );
  OR U10711 ( .A(n6606), .B(n6607), .Z(n6605) );
  OR U10712 ( .A(n6608), .B(n6609), .Z(n6604) );
  NAND U10713 ( .A(n6610), .B(n6611), .Z(n6567) );
  OR U10714 ( .A(n6612), .B(n6613), .Z(n6611) );
  OR U10715 ( .A(n6614), .B(n6615), .Z(n6610) );
  ANDN U10716 ( .B(n6616), .A(n6617), .Z(n6568) );
  IV U10717 ( .A(n6618), .Z(n6616) );
  ANDN U10718 ( .B(n6619), .A(n6620), .Z(n6560) );
  XOR U10719 ( .A(n6546), .B(n6621), .Z(n6558) );
  XOR U10720 ( .A(n6547), .B(n6548), .Z(n6621) );
  XOR U10721 ( .A(n6553), .B(n6622), .Z(n6548) );
  XOR U10722 ( .A(n6552), .B(n6555), .Z(n6622) );
  IV U10723 ( .A(n6554), .Z(n6555) );
  NAND U10724 ( .A(n6623), .B(n6624), .Z(n6554) );
  OR U10725 ( .A(n6625), .B(n6626), .Z(n6624) );
  OR U10726 ( .A(n6627), .B(n6628), .Z(n6623) );
  NAND U10727 ( .A(n6629), .B(n6630), .Z(n6552) );
  OR U10728 ( .A(n6631), .B(n6632), .Z(n6630) );
  OR U10729 ( .A(n6633), .B(n6634), .Z(n6629) );
  NOR U10730 ( .A(n6635), .B(n6636), .Z(n6553) );
  ANDN U10731 ( .B(n6637), .A(n6638), .Z(n6547) );
  IV U10732 ( .A(n6639), .Z(n6637) );
  XNOR U10733 ( .A(n6540), .B(n6640), .Z(n6546) );
  XNOR U10734 ( .A(n6539), .B(n6541), .Z(n6640) );
  NAND U10735 ( .A(n6641), .B(n6642), .Z(n6541) );
  OR U10736 ( .A(n6643), .B(n6644), .Z(n6642) );
  OR U10737 ( .A(n6645), .B(n6646), .Z(n6641) );
  NAND U10738 ( .A(n6647), .B(n6648), .Z(n6539) );
  OR U10739 ( .A(n6649), .B(n6650), .Z(n6648) );
  OR U10740 ( .A(n6651), .B(n6652), .Z(n6647) );
  ANDN U10741 ( .B(n6653), .A(n6654), .Z(n6540) );
  IV U10742 ( .A(n6655), .Z(n6653) );
  XNOR U10743 ( .A(n6620), .B(n6619), .Z(N29609) );
  XOR U10744 ( .A(n6639), .B(n6638), .Z(n6619) );
  XNOR U10745 ( .A(n6654), .B(n6655), .Z(n6638) );
  XNOR U10746 ( .A(n6649), .B(n6650), .Z(n6655) );
  XNOR U10747 ( .A(n6651), .B(n6652), .Z(n6650) );
  XNOR U10748 ( .A(y[3364]), .B(x[3364]), .Z(n6652) );
  XNOR U10749 ( .A(y[3365]), .B(x[3365]), .Z(n6651) );
  XNOR U10750 ( .A(y[3363]), .B(x[3363]), .Z(n6649) );
  XNOR U10751 ( .A(n6643), .B(n6644), .Z(n6654) );
  XNOR U10752 ( .A(y[3360]), .B(x[3360]), .Z(n6644) );
  XNOR U10753 ( .A(n6645), .B(n6646), .Z(n6643) );
  XNOR U10754 ( .A(y[3361]), .B(x[3361]), .Z(n6646) );
  XNOR U10755 ( .A(y[3362]), .B(x[3362]), .Z(n6645) );
  XNOR U10756 ( .A(n6636), .B(n6635), .Z(n6639) );
  XNOR U10757 ( .A(n6631), .B(n6632), .Z(n6635) );
  XNOR U10758 ( .A(y[3357]), .B(x[3357]), .Z(n6632) );
  XNOR U10759 ( .A(n6633), .B(n6634), .Z(n6631) );
  XNOR U10760 ( .A(y[3358]), .B(x[3358]), .Z(n6634) );
  XNOR U10761 ( .A(y[3359]), .B(x[3359]), .Z(n6633) );
  XNOR U10762 ( .A(n6625), .B(n6626), .Z(n6636) );
  XNOR U10763 ( .A(y[3354]), .B(x[3354]), .Z(n6626) );
  XNOR U10764 ( .A(n6627), .B(n6628), .Z(n6625) );
  XNOR U10765 ( .A(y[3355]), .B(x[3355]), .Z(n6628) );
  XNOR U10766 ( .A(y[3356]), .B(x[3356]), .Z(n6627) );
  XOR U10767 ( .A(n6601), .B(n6602), .Z(n6620) );
  XNOR U10768 ( .A(n6617), .B(n6618), .Z(n6602) );
  XNOR U10769 ( .A(n6612), .B(n6613), .Z(n6618) );
  XNOR U10770 ( .A(n6614), .B(n6615), .Z(n6613) );
  XNOR U10771 ( .A(y[3352]), .B(x[3352]), .Z(n6615) );
  XNOR U10772 ( .A(y[3353]), .B(x[3353]), .Z(n6614) );
  XNOR U10773 ( .A(y[3351]), .B(x[3351]), .Z(n6612) );
  XNOR U10774 ( .A(n6606), .B(n6607), .Z(n6617) );
  XNOR U10775 ( .A(y[3348]), .B(x[3348]), .Z(n6607) );
  XNOR U10776 ( .A(n6608), .B(n6609), .Z(n6606) );
  XNOR U10777 ( .A(y[3349]), .B(x[3349]), .Z(n6609) );
  XNOR U10778 ( .A(y[3350]), .B(x[3350]), .Z(n6608) );
  XOR U10779 ( .A(n6600), .B(n6599), .Z(n6601) );
  XNOR U10780 ( .A(n6595), .B(n6596), .Z(n6599) );
  XNOR U10781 ( .A(y[3345]), .B(x[3345]), .Z(n6596) );
  XNOR U10782 ( .A(n6597), .B(n6598), .Z(n6595) );
  XNOR U10783 ( .A(y[3346]), .B(x[3346]), .Z(n6598) );
  XNOR U10784 ( .A(y[3347]), .B(x[3347]), .Z(n6597) );
  XNOR U10785 ( .A(n6589), .B(n6590), .Z(n6600) );
  XNOR U10786 ( .A(y[3342]), .B(x[3342]), .Z(n6590) );
  XNOR U10787 ( .A(n6591), .B(n6592), .Z(n6589) );
  XNOR U10788 ( .A(y[3343]), .B(x[3343]), .Z(n6592) );
  XNOR U10789 ( .A(y[3344]), .B(x[3344]), .Z(n6591) );
  NAND U10790 ( .A(n6656), .B(n6657), .Z(N29601) );
  NANDN U10791 ( .A(n6658), .B(n6659), .Z(n6657) );
  OR U10792 ( .A(n6660), .B(n6661), .Z(n6659) );
  NAND U10793 ( .A(n6660), .B(n6661), .Z(n6656) );
  XOR U10794 ( .A(n6660), .B(n6662), .Z(N29600) );
  XNOR U10795 ( .A(n6658), .B(n6661), .Z(n6662) );
  AND U10796 ( .A(n6663), .B(n6664), .Z(n6661) );
  NANDN U10797 ( .A(n6665), .B(n6666), .Z(n6664) );
  NANDN U10798 ( .A(n6667), .B(n6668), .Z(n6666) );
  NANDN U10799 ( .A(n6668), .B(n6667), .Z(n6663) );
  NAND U10800 ( .A(n6669), .B(n6670), .Z(n6658) );
  NANDN U10801 ( .A(n6671), .B(n6672), .Z(n6670) );
  OR U10802 ( .A(n6673), .B(n6674), .Z(n6672) );
  NAND U10803 ( .A(n6674), .B(n6673), .Z(n6669) );
  AND U10804 ( .A(n6675), .B(n6676), .Z(n6660) );
  NANDN U10805 ( .A(n6677), .B(n6678), .Z(n6676) );
  NANDN U10806 ( .A(n6679), .B(n6680), .Z(n6678) );
  NANDN U10807 ( .A(n6680), .B(n6679), .Z(n6675) );
  XOR U10808 ( .A(n6674), .B(n6681), .Z(N29599) );
  XOR U10809 ( .A(n6671), .B(n6673), .Z(n6681) );
  XNOR U10810 ( .A(n6667), .B(n6682), .Z(n6673) );
  XNOR U10811 ( .A(n6665), .B(n6668), .Z(n6682) );
  NAND U10812 ( .A(n6683), .B(n6684), .Z(n6668) );
  NAND U10813 ( .A(n6685), .B(n6686), .Z(n6684) );
  OR U10814 ( .A(n6687), .B(n6688), .Z(n6685) );
  NANDN U10815 ( .A(n6689), .B(n6687), .Z(n6683) );
  IV U10816 ( .A(n6688), .Z(n6689) );
  NAND U10817 ( .A(n6690), .B(n6691), .Z(n6665) );
  NAND U10818 ( .A(n6692), .B(n6693), .Z(n6691) );
  NANDN U10819 ( .A(n6694), .B(n6695), .Z(n6692) );
  NANDN U10820 ( .A(n6695), .B(n6694), .Z(n6690) );
  AND U10821 ( .A(n6696), .B(n6697), .Z(n6667) );
  NAND U10822 ( .A(n6698), .B(n6699), .Z(n6697) );
  OR U10823 ( .A(n6700), .B(n6701), .Z(n6698) );
  NANDN U10824 ( .A(n6702), .B(n6700), .Z(n6696) );
  NAND U10825 ( .A(n6703), .B(n6704), .Z(n6671) );
  NANDN U10826 ( .A(n6705), .B(n6706), .Z(n6704) );
  OR U10827 ( .A(n6707), .B(n6708), .Z(n6706) );
  NANDN U10828 ( .A(n6709), .B(n6707), .Z(n6703) );
  IV U10829 ( .A(n6708), .Z(n6709) );
  XNOR U10830 ( .A(n6679), .B(n6710), .Z(n6674) );
  XNOR U10831 ( .A(n6677), .B(n6680), .Z(n6710) );
  NAND U10832 ( .A(n6711), .B(n6712), .Z(n6680) );
  NAND U10833 ( .A(n6713), .B(n6714), .Z(n6712) );
  OR U10834 ( .A(n6715), .B(n6716), .Z(n6713) );
  NANDN U10835 ( .A(n6717), .B(n6715), .Z(n6711) );
  IV U10836 ( .A(n6716), .Z(n6717) );
  NAND U10837 ( .A(n6718), .B(n6719), .Z(n6677) );
  NAND U10838 ( .A(n6720), .B(n6721), .Z(n6719) );
  NANDN U10839 ( .A(n6722), .B(n6723), .Z(n6720) );
  NANDN U10840 ( .A(n6723), .B(n6722), .Z(n6718) );
  AND U10841 ( .A(n6724), .B(n6725), .Z(n6679) );
  NAND U10842 ( .A(n6726), .B(n6727), .Z(n6725) );
  OR U10843 ( .A(n6728), .B(n6729), .Z(n6726) );
  NANDN U10844 ( .A(n6730), .B(n6728), .Z(n6724) );
  XNOR U10845 ( .A(n6705), .B(n6731), .Z(N29598) );
  XOR U10846 ( .A(n6707), .B(n6708), .Z(n6731) );
  XNOR U10847 ( .A(n6721), .B(n6732), .Z(n6708) );
  XOR U10848 ( .A(n6722), .B(n6723), .Z(n6732) );
  XOR U10849 ( .A(n6728), .B(n6733), .Z(n6723) );
  XOR U10850 ( .A(n6727), .B(n6730), .Z(n6733) );
  IV U10851 ( .A(n6729), .Z(n6730) );
  NAND U10852 ( .A(n6734), .B(n6735), .Z(n6729) );
  OR U10853 ( .A(n6736), .B(n6737), .Z(n6735) );
  OR U10854 ( .A(n6738), .B(n6739), .Z(n6734) );
  NAND U10855 ( .A(n6740), .B(n6741), .Z(n6727) );
  OR U10856 ( .A(n6742), .B(n6743), .Z(n6741) );
  OR U10857 ( .A(n6744), .B(n6745), .Z(n6740) );
  NOR U10858 ( .A(n6746), .B(n6747), .Z(n6728) );
  ANDN U10859 ( .B(n6748), .A(n6749), .Z(n6722) );
  XNOR U10860 ( .A(n6715), .B(n6750), .Z(n6721) );
  XNOR U10861 ( .A(n6714), .B(n6716), .Z(n6750) );
  NAND U10862 ( .A(n6751), .B(n6752), .Z(n6716) );
  OR U10863 ( .A(n6753), .B(n6754), .Z(n6752) );
  OR U10864 ( .A(n6755), .B(n6756), .Z(n6751) );
  NAND U10865 ( .A(n6757), .B(n6758), .Z(n6714) );
  OR U10866 ( .A(n6759), .B(n6760), .Z(n6758) );
  OR U10867 ( .A(n6761), .B(n6762), .Z(n6757) );
  ANDN U10868 ( .B(n6763), .A(n6764), .Z(n6715) );
  IV U10869 ( .A(n6765), .Z(n6763) );
  ANDN U10870 ( .B(n6766), .A(n6767), .Z(n6707) );
  XOR U10871 ( .A(n6693), .B(n6768), .Z(n6705) );
  XOR U10872 ( .A(n6694), .B(n6695), .Z(n6768) );
  XOR U10873 ( .A(n6700), .B(n6769), .Z(n6695) );
  XOR U10874 ( .A(n6699), .B(n6702), .Z(n6769) );
  IV U10875 ( .A(n6701), .Z(n6702) );
  NAND U10876 ( .A(n6770), .B(n6771), .Z(n6701) );
  OR U10877 ( .A(n6772), .B(n6773), .Z(n6771) );
  OR U10878 ( .A(n6774), .B(n6775), .Z(n6770) );
  NAND U10879 ( .A(n6776), .B(n6777), .Z(n6699) );
  OR U10880 ( .A(n6778), .B(n6779), .Z(n6777) );
  OR U10881 ( .A(n6780), .B(n6781), .Z(n6776) );
  NOR U10882 ( .A(n6782), .B(n6783), .Z(n6700) );
  ANDN U10883 ( .B(n6784), .A(n6785), .Z(n6694) );
  IV U10884 ( .A(n6786), .Z(n6784) );
  XNOR U10885 ( .A(n6687), .B(n6787), .Z(n6693) );
  XNOR U10886 ( .A(n6686), .B(n6688), .Z(n6787) );
  NAND U10887 ( .A(n6788), .B(n6789), .Z(n6688) );
  OR U10888 ( .A(n6790), .B(n6791), .Z(n6789) );
  OR U10889 ( .A(n6792), .B(n6793), .Z(n6788) );
  NAND U10890 ( .A(n6794), .B(n6795), .Z(n6686) );
  OR U10891 ( .A(n6796), .B(n6797), .Z(n6795) );
  OR U10892 ( .A(n6798), .B(n6799), .Z(n6794) );
  ANDN U10893 ( .B(n6800), .A(n6801), .Z(n6687) );
  IV U10894 ( .A(n6802), .Z(n6800) );
  XNOR U10895 ( .A(n6767), .B(n6766), .Z(N29597) );
  XOR U10896 ( .A(n6786), .B(n6785), .Z(n6766) );
  XNOR U10897 ( .A(n6801), .B(n6802), .Z(n6785) );
  XNOR U10898 ( .A(n6796), .B(n6797), .Z(n6802) );
  XNOR U10899 ( .A(n6798), .B(n6799), .Z(n6797) );
  XNOR U10900 ( .A(y[3340]), .B(x[3340]), .Z(n6799) );
  XNOR U10901 ( .A(y[3341]), .B(x[3341]), .Z(n6798) );
  XNOR U10902 ( .A(y[3339]), .B(x[3339]), .Z(n6796) );
  XNOR U10903 ( .A(n6790), .B(n6791), .Z(n6801) );
  XNOR U10904 ( .A(y[3336]), .B(x[3336]), .Z(n6791) );
  XNOR U10905 ( .A(n6792), .B(n6793), .Z(n6790) );
  XNOR U10906 ( .A(y[3337]), .B(x[3337]), .Z(n6793) );
  XNOR U10907 ( .A(y[3338]), .B(x[3338]), .Z(n6792) );
  XNOR U10908 ( .A(n6783), .B(n6782), .Z(n6786) );
  XNOR U10909 ( .A(n6778), .B(n6779), .Z(n6782) );
  XNOR U10910 ( .A(y[3333]), .B(x[3333]), .Z(n6779) );
  XNOR U10911 ( .A(n6780), .B(n6781), .Z(n6778) );
  XNOR U10912 ( .A(y[3334]), .B(x[3334]), .Z(n6781) );
  XNOR U10913 ( .A(y[3335]), .B(x[3335]), .Z(n6780) );
  XNOR U10914 ( .A(n6772), .B(n6773), .Z(n6783) );
  XNOR U10915 ( .A(y[3330]), .B(x[3330]), .Z(n6773) );
  XNOR U10916 ( .A(n6774), .B(n6775), .Z(n6772) );
  XNOR U10917 ( .A(y[3331]), .B(x[3331]), .Z(n6775) );
  XNOR U10918 ( .A(y[3332]), .B(x[3332]), .Z(n6774) );
  XOR U10919 ( .A(n6748), .B(n6749), .Z(n6767) );
  XNOR U10920 ( .A(n6764), .B(n6765), .Z(n6749) );
  XNOR U10921 ( .A(n6759), .B(n6760), .Z(n6765) );
  XNOR U10922 ( .A(n6761), .B(n6762), .Z(n6760) );
  XNOR U10923 ( .A(y[3328]), .B(x[3328]), .Z(n6762) );
  XNOR U10924 ( .A(y[3329]), .B(x[3329]), .Z(n6761) );
  XNOR U10925 ( .A(y[3327]), .B(x[3327]), .Z(n6759) );
  XNOR U10926 ( .A(n6753), .B(n6754), .Z(n6764) );
  XNOR U10927 ( .A(y[3324]), .B(x[3324]), .Z(n6754) );
  XNOR U10928 ( .A(n6755), .B(n6756), .Z(n6753) );
  XNOR U10929 ( .A(y[3325]), .B(x[3325]), .Z(n6756) );
  XNOR U10930 ( .A(y[3326]), .B(x[3326]), .Z(n6755) );
  XOR U10931 ( .A(n6747), .B(n6746), .Z(n6748) );
  XNOR U10932 ( .A(n6742), .B(n6743), .Z(n6746) );
  XNOR U10933 ( .A(y[3321]), .B(x[3321]), .Z(n6743) );
  XNOR U10934 ( .A(n6744), .B(n6745), .Z(n6742) );
  XNOR U10935 ( .A(y[3322]), .B(x[3322]), .Z(n6745) );
  XNOR U10936 ( .A(y[3323]), .B(x[3323]), .Z(n6744) );
  XNOR U10937 ( .A(n6736), .B(n6737), .Z(n6747) );
  XNOR U10938 ( .A(y[3318]), .B(x[3318]), .Z(n6737) );
  XNOR U10939 ( .A(n6738), .B(n6739), .Z(n6736) );
  XNOR U10940 ( .A(y[3319]), .B(x[3319]), .Z(n6739) );
  XNOR U10941 ( .A(y[3320]), .B(x[3320]), .Z(n6738) );
  NAND U10942 ( .A(n6803), .B(n6804), .Z(N29589) );
  NANDN U10943 ( .A(n6805), .B(n6806), .Z(n6804) );
  OR U10944 ( .A(n6807), .B(n6808), .Z(n6806) );
  NAND U10945 ( .A(n6807), .B(n6808), .Z(n6803) );
  XOR U10946 ( .A(n6807), .B(n6809), .Z(N29588) );
  XNOR U10947 ( .A(n6805), .B(n6808), .Z(n6809) );
  AND U10948 ( .A(n6810), .B(n6811), .Z(n6808) );
  NANDN U10949 ( .A(n6812), .B(n6813), .Z(n6811) );
  NANDN U10950 ( .A(n6814), .B(n6815), .Z(n6813) );
  NANDN U10951 ( .A(n6815), .B(n6814), .Z(n6810) );
  NAND U10952 ( .A(n6816), .B(n6817), .Z(n6805) );
  NANDN U10953 ( .A(n6818), .B(n6819), .Z(n6817) );
  OR U10954 ( .A(n6820), .B(n6821), .Z(n6819) );
  NAND U10955 ( .A(n6821), .B(n6820), .Z(n6816) );
  AND U10956 ( .A(n6822), .B(n6823), .Z(n6807) );
  NANDN U10957 ( .A(n6824), .B(n6825), .Z(n6823) );
  NANDN U10958 ( .A(n6826), .B(n6827), .Z(n6825) );
  NANDN U10959 ( .A(n6827), .B(n6826), .Z(n6822) );
  XOR U10960 ( .A(n6821), .B(n6828), .Z(N29587) );
  XOR U10961 ( .A(n6818), .B(n6820), .Z(n6828) );
  XNOR U10962 ( .A(n6814), .B(n6829), .Z(n6820) );
  XNOR U10963 ( .A(n6812), .B(n6815), .Z(n6829) );
  NAND U10964 ( .A(n6830), .B(n6831), .Z(n6815) );
  NAND U10965 ( .A(n6832), .B(n6833), .Z(n6831) );
  OR U10966 ( .A(n6834), .B(n6835), .Z(n6832) );
  NANDN U10967 ( .A(n6836), .B(n6834), .Z(n6830) );
  IV U10968 ( .A(n6835), .Z(n6836) );
  NAND U10969 ( .A(n6837), .B(n6838), .Z(n6812) );
  NAND U10970 ( .A(n6839), .B(n6840), .Z(n6838) );
  NANDN U10971 ( .A(n6841), .B(n6842), .Z(n6839) );
  NANDN U10972 ( .A(n6842), .B(n6841), .Z(n6837) );
  AND U10973 ( .A(n6843), .B(n6844), .Z(n6814) );
  NAND U10974 ( .A(n6845), .B(n6846), .Z(n6844) );
  OR U10975 ( .A(n6847), .B(n6848), .Z(n6845) );
  NANDN U10976 ( .A(n6849), .B(n6847), .Z(n6843) );
  NAND U10977 ( .A(n6850), .B(n6851), .Z(n6818) );
  NANDN U10978 ( .A(n6852), .B(n6853), .Z(n6851) );
  OR U10979 ( .A(n6854), .B(n6855), .Z(n6853) );
  NANDN U10980 ( .A(n6856), .B(n6854), .Z(n6850) );
  IV U10981 ( .A(n6855), .Z(n6856) );
  XNOR U10982 ( .A(n6826), .B(n6857), .Z(n6821) );
  XNOR U10983 ( .A(n6824), .B(n6827), .Z(n6857) );
  NAND U10984 ( .A(n6858), .B(n6859), .Z(n6827) );
  NAND U10985 ( .A(n6860), .B(n6861), .Z(n6859) );
  OR U10986 ( .A(n6862), .B(n6863), .Z(n6860) );
  NANDN U10987 ( .A(n6864), .B(n6862), .Z(n6858) );
  IV U10988 ( .A(n6863), .Z(n6864) );
  NAND U10989 ( .A(n6865), .B(n6866), .Z(n6824) );
  NAND U10990 ( .A(n6867), .B(n6868), .Z(n6866) );
  NANDN U10991 ( .A(n6869), .B(n6870), .Z(n6867) );
  NANDN U10992 ( .A(n6870), .B(n6869), .Z(n6865) );
  AND U10993 ( .A(n6871), .B(n6872), .Z(n6826) );
  NAND U10994 ( .A(n6873), .B(n6874), .Z(n6872) );
  OR U10995 ( .A(n6875), .B(n6876), .Z(n6873) );
  NANDN U10996 ( .A(n6877), .B(n6875), .Z(n6871) );
  XNOR U10997 ( .A(n6852), .B(n6878), .Z(N29586) );
  XOR U10998 ( .A(n6854), .B(n6855), .Z(n6878) );
  XNOR U10999 ( .A(n6868), .B(n6879), .Z(n6855) );
  XOR U11000 ( .A(n6869), .B(n6870), .Z(n6879) );
  XOR U11001 ( .A(n6875), .B(n6880), .Z(n6870) );
  XOR U11002 ( .A(n6874), .B(n6877), .Z(n6880) );
  IV U11003 ( .A(n6876), .Z(n6877) );
  NAND U11004 ( .A(n6881), .B(n6882), .Z(n6876) );
  OR U11005 ( .A(n6883), .B(n6884), .Z(n6882) );
  OR U11006 ( .A(n6885), .B(n6886), .Z(n6881) );
  NAND U11007 ( .A(n6887), .B(n6888), .Z(n6874) );
  OR U11008 ( .A(n6889), .B(n6890), .Z(n6888) );
  OR U11009 ( .A(n6891), .B(n6892), .Z(n6887) );
  NOR U11010 ( .A(n6893), .B(n6894), .Z(n6875) );
  ANDN U11011 ( .B(n6895), .A(n6896), .Z(n6869) );
  XNOR U11012 ( .A(n6862), .B(n6897), .Z(n6868) );
  XNOR U11013 ( .A(n6861), .B(n6863), .Z(n6897) );
  NAND U11014 ( .A(n6898), .B(n6899), .Z(n6863) );
  OR U11015 ( .A(n6900), .B(n6901), .Z(n6899) );
  OR U11016 ( .A(n6902), .B(n6903), .Z(n6898) );
  NAND U11017 ( .A(n6904), .B(n6905), .Z(n6861) );
  OR U11018 ( .A(n6906), .B(n6907), .Z(n6905) );
  OR U11019 ( .A(n6908), .B(n6909), .Z(n6904) );
  ANDN U11020 ( .B(n6910), .A(n6911), .Z(n6862) );
  IV U11021 ( .A(n6912), .Z(n6910) );
  ANDN U11022 ( .B(n6913), .A(n6914), .Z(n6854) );
  XOR U11023 ( .A(n6840), .B(n6915), .Z(n6852) );
  XOR U11024 ( .A(n6841), .B(n6842), .Z(n6915) );
  XOR U11025 ( .A(n6847), .B(n6916), .Z(n6842) );
  XOR U11026 ( .A(n6846), .B(n6849), .Z(n6916) );
  IV U11027 ( .A(n6848), .Z(n6849) );
  NAND U11028 ( .A(n6917), .B(n6918), .Z(n6848) );
  OR U11029 ( .A(n6919), .B(n6920), .Z(n6918) );
  OR U11030 ( .A(n6921), .B(n6922), .Z(n6917) );
  NAND U11031 ( .A(n6923), .B(n6924), .Z(n6846) );
  OR U11032 ( .A(n6925), .B(n6926), .Z(n6924) );
  OR U11033 ( .A(n6927), .B(n6928), .Z(n6923) );
  NOR U11034 ( .A(n6929), .B(n6930), .Z(n6847) );
  ANDN U11035 ( .B(n6931), .A(n6932), .Z(n6841) );
  IV U11036 ( .A(n6933), .Z(n6931) );
  XNOR U11037 ( .A(n6834), .B(n6934), .Z(n6840) );
  XNOR U11038 ( .A(n6833), .B(n6835), .Z(n6934) );
  NAND U11039 ( .A(n6935), .B(n6936), .Z(n6835) );
  OR U11040 ( .A(n6937), .B(n6938), .Z(n6936) );
  OR U11041 ( .A(n6939), .B(n6940), .Z(n6935) );
  NAND U11042 ( .A(n6941), .B(n6942), .Z(n6833) );
  OR U11043 ( .A(n6943), .B(n6944), .Z(n6942) );
  OR U11044 ( .A(n6945), .B(n6946), .Z(n6941) );
  ANDN U11045 ( .B(n6947), .A(n6948), .Z(n6834) );
  IV U11046 ( .A(n6949), .Z(n6947) );
  XNOR U11047 ( .A(n6914), .B(n6913), .Z(N29585) );
  XOR U11048 ( .A(n6933), .B(n6932), .Z(n6913) );
  XNOR U11049 ( .A(n6948), .B(n6949), .Z(n6932) );
  XNOR U11050 ( .A(n6943), .B(n6944), .Z(n6949) );
  XNOR U11051 ( .A(n6945), .B(n6946), .Z(n6944) );
  XNOR U11052 ( .A(y[3316]), .B(x[3316]), .Z(n6946) );
  XNOR U11053 ( .A(y[3317]), .B(x[3317]), .Z(n6945) );
  XNOR U11054 ( .A(y[3315]), .B(x[3315]), .Z(n6943) );
  XNOR U11055 ( .A(n6937), .B(n6938), .Z(n6948) );
  XNOR U11056 ( .A(y[3312]), .B(x[3312]), .Z(n6938) );
  XNOR U11057 ( .A(n6939), .B(n6940), .Z(n6937) );
  XNOR U11058 ( .A(y[3313]), .B(x[3313]), .Z(n6940) );
  XNOR U11059 ( .A(y[3314]), .B(x[3314]), .Z(n6939) );
  XNOR U11060 ( .A(n6930), .B(n6929), .Z(n6933) );
  XNOR U11061 ( .A(n6925), .B(n6926), .Z(n6929) );
  XNOR U11062 ( .A(y[3309]), .B(x[3309]), .Z(n6926) );
  XNOR U11063 ( .A(n6927), .B(n6928), .Z(n6925) );
  XNOR U11064 ( .A(y[3310]), .B(x[3310]), .Z(n6928) );
  XNOR U11065 ( .A(y[3311]), .B(x[3311]), .Z(n6927) );
  XNOR U11066 ( .A(n6919), .B(n6920), .Z(n6930) );
  XNOR U11067 ( .A(y[3306]), .B(x[3306]), .Z(n6920) );
  XNOR U11068 ( .A(n6921), .B(n6922), .Z(n6919) );
  XNOR U11069 ( .A(y[3307]), .B(x[3307]), .Z(n6922) );
  XNOR U11070 ( .A(y[3308]), .B(x[3308]), .Z(n6921) );
  XOR U11071 ( .A(n6895), .B(n6896), .Z(n6914) );
  XNOR U11072 ( .A(n6911), .B(n6912), .Z(n6896) );
  XNOR U11073 ( .A(n6906), .B(n6907), .Z(n6912) );
  XNOR U11074 ( .A(n6908), .B(n6909), .Z(n6907) );
  XNOR U11075 ( .A(y[3304]), .B(x[3304]), .Z(n6909) );
  XNOR U11076 ( .A(y[3305]), .B(x[3305]), .Z(n6908) );
  XNOR U11077 ( .A(y[3303]), .B(x[3303]), .Z(n6906) );
  XNOR U11078 ( .A(n6900), .B(n6901), .Z(n6911) );
  XNOR U11079 ( .A(y[3300]), .B(x[3300]), .Z(n6901) );
  XNOR U11080 ( .A(n6902), .B(n6903), .Z(n6900) );
  XNOR U11081 ( .A(y[3301]), .B(x[3301]), .Z(n6903) );
  XNOR U11082 ( .A(y[3302]), .B(x[3302]), .Z(n6902) );
  XOR U11083 ( .A(n6894), .B(n6893), .Z(n6895) );
  XNOR U11084 ( .A(n6889), .B(n6890), .Z(n6893) );
  XNOR U11085 ( .A(y[3297]), .B(x[3297]), .Z(n6890) );
  XNOR U11086 ( .A(n6891), .B(n6892), .Z(n6889) );
  XNOR U11087 ( .A(y[3298]), .B(x[3298]), .Z(n6892) );
  XNOR U11088 ( .A(y[3299]), .B(x[3299]), .Z(n6891) );
  XNOR U11089 ( .A(n6883), .B(n6884), .Z(n6894) );
  XNOR U11090 ( .A(y[3294]), .B(x[3294]), .Z(n6884) );
  XNOR U11091 ( .A(n6885), .B(n6886), .Z(n6883) );
  XNOR U11092 ( .A(y[3295]), .B(x[3295]), .Z(n6886) );
  XNOR U11093 ( .A(y[3296]), .B(x[3296]), .Z(n6885) );
  NAND U11094 ( .A(n6950), .B(n6951), .Z(N29577) );
  NANDN U11095 ( .A(n6952), .B(n6953), .Z(n6951) );
  OR U11096 ( .A(n6954), .B(n6955), .Z(n6953) );
  NAND U11097 ( .A(n6954), .B(n6955), .Z(n6950) );
  XOR U11098 ( .A(n6954), .B(n6956), .Z(N29576) );
  XNOR U11099 ( .A(n6952), .B(n6955), .Z(n6956) );
  AND U11100 ( .A(n6957), .B(n6958), .Z(n6955) );
  NANDN U11101 ( .A(n6959), .B(n6960), .Z(n6958) );
  NANDN U11102 ( .A(n6961), .B(n6962), .Z(n6960) );
  NANDN U11103 ( .A(n6962), .B(n6961), .Z(n6957) );
  NAND U11104 ( .A(n6963), .B(n6964), .Z(n6952) );
  NANDN U11105 ( .A(n6965), .B(n6966), .Z(n6964) );
  OR U11106 ( .A(n6967), .B(n6968), .Z(n6966) );
  NAND U11107 ( .A(n6968), .B(n6967), .Z(n6963) );
  AND U11108 ( .A(n6969), .B(n6970), .Z(n6954) );
  NANDN U11109 ( .A(n6971), .B(n6972), .Z(n6970) );
  NANDN U11110 ( .A(n6973), .B(n6974), .Z(n6972) );
  NANDN U11111 ( .A(n6974), .B(n6973), .Z(n6969) );
  XOR U11112 ( .A(n6968), .B(n6975), .Z(N29575) );
  XOR U11113 ( .A(n6965), .B(n6967), .Z(n6975) );
  XNOR U11114 ( .A(n6961), .B(n6976), .Z(n6967) );
  XNOR U11115 ( .A(n6959), .B(n6962), .Z(n6976) );
  NAND U11116 ( .A(n6977), .B(n6978), .Z(n6962) );
  NAND U11117 ( .A(n6979), .B(n6980), .Z(n6978) );
  OR U11118 ( .A(n6981), .B(n6982), .Z(n6979) );
  NANDN U11119 ( .A(n6983), .B(n6981), .Z(n6977) );
  IV U11120 ( .A(n6982), .Z(n6983) );
  NAND U11121 ( .A(n6984), .B(n6985), .Z(n6959) );
  NAND U11122 ( .A(n6986), .B(n6987), .Z(n6985) );
  NANDN U11123 ( .A(n6988), .B(n6989), .Z(n6986) );
  NANDN U11124 ( .A(n6989), .B(n6988), .Z(n6984) );
  AND U11125 ( .A(n6990), .B(n6991), .Z(n6961) );
  NAND U11126 ( .A(n6992), .B(n6993), .Z(n6991) );
  OR U11127 ( .A(n6994), .B(n6995), .Z(n6992) );
  NANDN U11128 ( .A(n6996), .B(n6994), .Z(n6990) );
  NAND U11129 ( .A(n6997), .B(n6998), .Z(n6965) );
  NANDN U11130 ( .A(n6999), .B(n7000), .Z(n6998) );
  OR U11131 ( .A(n7001), .B(n7002), .Z(n7000) );
  NANDN U11132 ( .A(n7003), .B(n7001), .Z(n6997) );
  IV U11133 ( .A(n7002), .Z(n7003) );
  XNOR U11134 ( .A(n6973), .B(n7004), .Z(n6968) );
  XNOR U11135 ( .A(n6971), .B(n6974), .Z(n7004) );
  NAND U11136 ( .A(n7005), .B(n7006), .Z(n6974) );
  NAND U11137 ( .A(n7007), .B(n7008), .Z(n7006) );
  OR U11138 ( .A(n7009), .B(n7010), .Z(n7007) );
  NANDN U11139 ( .A(n7011), .B(n7009), .Z(n7005) );
  IV U11140 ( .A(n7010), .Z(n7011) );
  NAND U11141 ( .A(n7012), .B(n7013), .Z(n6971) );
  NAND U11142 ( .A(n7014), .B(n7015), .Z(n7013) );
  NANDN U11143 ( .A(n7016), .B(n7017), .Z(n7014) );
  NANDN U11144 ( .A(n7017), .B(n7016), .Z(n7012) );
  AND U11145 ( .A(n7018), .B(n7019), .Z(n6973) );
  NAND U11146 ( .A(n7020), .B(n7021), .Z(n7019) );
  OR U11147 ( .A(n7022), .B(n7023), .Z(n7020) );
  NANDN U11148 ( .A(n7024), .B(n7022), .Z(n7018) );
  XNOR U11149 ( .A(n6999), .B(n7025), .Z(N29574) );
  XOR U11150 ( .A(n7001), .B(n7002), .Z(n7025) );
  XNOR U11151 ( .A(n7015), .B(n7026), .Z(n7002) );
  XOR U11152 ( .A(n7016), .B(n7017), .Z(n7026) );
  XOR U11153 ( .A(n7022), .B(n7027), .Z(n7017) );
  XOR U11154 ( .A(n7021), .B(n7024), .Z(n7027) );
  IV U11155 ( .A(n7023), .Z(n7024) );
  NAND U11156 ( .A(n7028), .B(n7029), .Z(n7023) );
  OR U11157 ( .A(n7030), .B(n7031), .Z(n7029) );
  OR U11158 ( .A(n7032), .B(n7033), .Z(n7028) );
  NAND U11159 ( .A(n7034), .B(n7035), .Z(n7021) );
  OR U11160 ( .A(n7036), .B(n7037), .Z(n7035) );
  OR U11161 ( .A(n7038), .B(n7039), .Z(n7034) );
  NOR U11162 ( .A(n7040), .B(n7041), .Z(n7022) );
  ANDN U11163 ( .B(n7042), .A(n7043), .Z(n7016) );
  XNOR U11164 ( .A(n7009), .B(n7044), .Z(n7015) );
  XNOR U11165 ( .A(n7008), .B(n7010), .Z(n7044) );
  NAND U11166 ( .A(n7045), .B(n7046), .Z(n7010) );
  OR U11167 ( .A(n7047), .B(n7048), .Z(n7046) );
  OR U11168 ( .A(n7049), .B(n7050), .Z(n7045) );
  NAND U11169 ( .A(n7051), .B(n7052), .Z(n7008) );
  OR U11170 ( .A(n7053), .B(n7054), .Z(n7052) );
  OR U11171 ( .A(n7055), .B(n7056), .Z(n7051) );
  ANDN U11172 ( .B(n7057), .A(n7058), .Z(n7009) );
  IV U11173 ( .A(n7059), .Z(n7057) );
  ANDN U11174 ( .B(n7060), .A(n7061), .Z(n7001) );
  XOR U11175 ( .A(n6987), .B(n7062), .Z(n6999) );
  XOR U11176 ( .A(n6988), .B(n6989), .Z(n7062) );
  XOR U11177 ( .A(n6994), .B(n7063), .Z(n6989) );
  XOR U11178 ( .A(n6993), .B(n6996), .Z(n7063) );
  IV U11179 ( .A(n6995), .Z(n6996) );
  NAND U11180 ( .A(n7064), .B(n7065), .Z(n6995) );
  OR U11181 ( .A(n7066), .B(n7067), .Z(n7065) );
  OR U11182 ( .A(n7068), .B(n7069), .Z(n7064) );
  NAND U11183 ( .A(n7070), .B(n7071), .Z(n6993) );
  OR U11184 ( .A(n7072), .B(n7073), .Z(n7071) );
  OR U11185 ( .A(n7074), .B(n7075), .Z(n7070) );
  NOR U11186 ( .A(n7076), .B(n7077), .Z(n6994) );
  ANDN U11187 ( .B(n7078), .A(n7079), .Z(n6988) );
  IV U11188 ( .A(n7080), .Z(n7078) );
  XNOR U11189 ( .A(n6981), .B(n7081), .Z(n6987) );
  XNOR U11190 ( .A(n6980), .B(n6982), .Z(n7081) );
  NAND U11191 ( .A(n7082), .B(n7083), .Z(n6982) );
  OR U11192 ( .A(n7084), .B(n7085), .Z(n7083) );
  OR U11193 ( .A(n7086), .B(n7087), .Z(n7082) );
  NAND U11194 ( .A(n7088), .B(n7089), .Z(n6980) );
  OR U11195 ( .A(n7090), .B(n7091), .Z(n7089) );
  OR U11196 ( .A(n7092), .B(n7093), .Z(n7088) );
  ANDN U11197 ( .B(n7094), .A(n7095), .Z(n6981) );
  IV U11198 ( .A(n7096), .Z(n7094) );
  XNOR U11199 ( .A(n7061), .B(n7060), .Z(N29573) );
  XOR U11200 ( .A(n7080), .B(n7079), .Z(n7060) );
  XNOR U11201 ( .A(n7095), .B(n7096), .Z(n7079) );
  XNOR U11202 ( .A(n7090), .B(n7091), .Z(n7096) );
  XNOR U11203 ( .A(n7092), .B(n7093), .Z(n7091) );
  XNOR U11204 ( .A(y[3292]), .B(x[3292]), .Z(n7093) );
  XNOR U11205 ( .A(y[3293]), .B(x[3293]), .Z(n7092) );
  XNOR U11206 ( .A(y[3291]), .B(x[3291]), .Z(n7090) );
  XNOR U11207 ( .A(n7084), .B(n7085), .Z(n7095) );
  XNOR U11208 ( .A(y[3288]), .B(x[3288]), .Z(n7085) );
  XNOR U11209 ( .A(n7086), .B(n7087), .Z(n7084) );
  XNOR U11210 ( .A(y[3289]), .B(x[3289]), .Z(n7087) );
  XNOR U11211 ( .A(y[3290]), .B(x[3290]), .Z(n7086) );
  XNOR U11212 ( .A(n7077), .B(n7076), .Z(n7080) );
  XNOR U11213 ( .A(n7072), .B(n7073), .Z(n7076) );
  XNOR U11214 ( .A(y[3285]), .B(x[3285]), .Z(n7073) );
  XNOR U11215 ( .A(n7074), .B(n7075), .Z(n7072) );
  XNOR U11216 ( .A(y[3286]), .B(x[3286]), .Z(n7075) );
  XNOR U11217 ( .A(y[3287]), .B(x[3287]), .Z(n7074) );
  XNOR U11218 ( .A(n7066), .B(n7067), .Z(n7077) );
  XNOR U11219 ( .A(y[3282]), .B(x[3282]), .Z(n7067) );
  XNOR U11220 ( .A(n7068), .B(n7069), .Z(n7066) );
  XNOR U11221 ( .A(y[3283]), .B(x[3283]), .Z(n7069) );
  XNOR U11222 ( .A(y[3284]), .B(x[3284]), .Z(n7068) );
  XOR U11223 ( .A(n7042), .B(n7043), .Z(n7061) );
  XNOR U11224 ( .A(n7058), .B(n7059), .Z(n7043) );
  XNOR U11225 ( .A(n7053), .B(n7054), .Z(n7059) );
  XNOR U11226 ( .A(n7055), .B(n7056), .Z(n7054) );
  XNOR U11227 ( .A(y[3280]), .B(x[3280]), .Z(n7056) );
  XNOR U11228 ( .A(y[3281]), .B(x[3281]), .Z(n7055) );
  XNOR U11229 ( .A(y[3279]), .B(x[3279]), .Z(n7053) );
  XNOR U11230 ( .A(n7047), .B(n7048), .Z(n7058) );
  XNOR U11231 ( .A(y[3276]), .B(x[3276]), .Z(n7048) );
  XNOR U11232 ( .A(n7049), .B(n7050), .Z(n7047) );
  XNOR U11233 ( .A(y[3277]), .B(x[3277]), .Z(n7050) );
  XNOR U11234 ( .A(y[3278]), .B(x[3278]), .Z(n7049) );
  XOR U11235 ( .A(n7041), .B(n7040), .Z(n7042) );
  XNOR U11236 ( .A(n7036), .B(n7037), .Z(n7040) );
  XNOR U11237 ( .A(y[3273]), .B(x[3273]), .Z(n7037) );
  XNOR U11238 ( .A(n7038), .B(n7039), .Z(n7036) );
  XNOR U11239 ( .A(y[3274]), .B(x[3274]), .Z(n7039) );
  XNOR U11240 ( .A(y[3275]), .B(x[3275]), .Z(n7038) );
  XNOR U11241 ( .A(n7030), .B(n7031), .Z(n7041) );
  XNOR U11242 ( .A(y[3270]), .B(x[3270]), .Z(n7031) );
  XNOR U11243 ( .A(n7032), .B(n7033), .Z(n7030) );
  XNOR U11244 ( .A(y[3271]), .B(x[3271]), .Z(n7033) );
  XNOR U11245 ( .A(y[3272]), .B(x[3272]), .Z(n7032) );
  NAND U11246 ( .A(n7097), .B(n7098), .Z(N29565) );
  NANDN U11247 ( .A(n7099), .B(n7100), .Z(n7098) );
  OR U11248 ( .A(n7101), .B(n7102), .Z(n7100) );
  NAND U11249 ( .A(n7101), .B(n7102), .Z(n7097) );
  XOR U11250 ( .A(n7101), .B(n7103), .Z(N29564) );
  XNOR U11251 ( .A(n7099), .B(n7102), .Z(n7103) );
  AND U11252 ( .A(n7104), .B(n7105), .Z(n7102) );
  NANDN U11253 ( .A(n7106), .B(n7107), .Z(n7105) );
  NANDN U11254 ( .A(n7108), .B(n7109), .Z(n7107) );
  NANDN U11255 ( .A(n7109), .B(n7108), .Z(n7104) );
  NAND U11256 ( .A(n7110), .B(n7111), .Z(n7099) );
  NANDN U11257 ( .A(n7112), .B(n7113), .Z(n7111) );
  OR U11258 ( .A(n7114), .B(n7115), .Z(n7113) );
  NAND U11259 ( .A(n7115), .B(n7114), .Z(n7110) );
  AND U11260 ( .A(n7116), .B(n7117), .Z(n7101) );
  NANDN U11261 ( .A(n7118), .B(n7119), .Z(n7117) );
  NANDN U11262 ( .A(n7120), .B(n7121), .Z(n7119) );
  NANDN U11263 ( .A(n7121), .B(n7120), .Z(n7116) );
  XOR U11264 ( .A(n7115), .B(n7122), .Z(N29563) );
  XOR U11265 ( .A(n7112), .B(n7114), .Z(n7122) );
  XNOR U11266 ( .A(n7108), .B(n7123), .Z(n7114) );
  XNOR U11267 ( .A(n7106), .B(n7109), .Z(n7123) );
  NAND U11268 ( .A(n7124), .B(n7125), .Z(n7109) );
  NAND U11269 ( .A(n7126), .B(n7127), .Z(n7125) );
  OR U11270 ( .A(n7128), .B(n7129), .Z(n7126) );
  NANDN U11271 ( .A(n7130), .B(n7128), .Z(n7124) );
  IV U11272 ( .A(n7129), .Z(n7130) );
  NAND U11273 ( .A(n7131), .B(n7132), .Z(n7106) );
  NAND U11274 ( .A(n7133), .B(n7134), .Z(n7132) );
  NANDN U11275 ( .A(n7135), .B(n7136), .Z(n7133) );
  NANDN U11276 ( .A(n7136), .B(n7135), .Z(n7131) );
  AND U11277 ( .A(n7137), .B(n7138), .Z(n7108) );
  NAND U11278 ( .A(n7139), .B(n7140), .Z(n7138) );
  OR U11279 ( .A(n7141), .B(n7142), .Z(n7139) );
  NANDN U11280 ( .A(n7143), .B(n7141), .Z(n7137) );
  NAND U11281 ( .A(n7144), .B(n7145), .Z(n7112) );
  NANDN U11282 ( .A(n7146), .B(n7147), .Z(n7145) );
  OR U11283 ( .A(n7148), .B(n7149), .Z(n7147) );
  NANDN U11284 ( .A(n7150), .B(n7148), .Z(n7144) );
  IV U11285 ( .A(n7149), .Z(n7150) );
  XNOR U11286 ( .A(n7120), .B(n7151), .Z(n7115) );
  XNOR U11287 ( .A(n7118), .B(n7121), .Z(n7151) );
  NAND U11288 ( .A(n7152), .B(n7153), .Z(n7121) );
  NAND U11289 ( .A(n7154), .B(n7155), .Z(n7153) );
  OR U11290 ( .A(n7156), .B(n7157), .Z(n7154) );
  NANDN U11291 ( .A(n7158), .B(n7156), .Z(n7152) );
  IV U11292 ( .A(n7157), .Z(n7158) );
  NAND U11293 ( .A(n7159), .B(n7160), .Z(n7118) );
  NAND U11294 ( .A(n7161), .B(n7162), .Z(n7160) );
  NANDN U11295 ( .A(n7163), .B(n7164), .Z(n7161) );
  NANDN U11296 ( .A(n7164), .B(n7163), .Z(n7159) );
  AND U11297 ( .A(n7165), .B(n7166), .Z(n7120) );
  NAND U11298 ( .A(n7167), .B(n7168), .Z(n7166) );
  OR U11299 ( .A(n7169), .B(n7170), .Z(n7167) );
  NANDN U11300 ( .A(n7171), .B(n7169), .Z(n7165) );
  XNOR U11301 ( .A(n7146), .B(n7172), .Z(N29562) );
  XOR U11302 ( .A(n7148), .B(n7149), .Z(n7172) );
  XNOR U11303 ( .A(n7162), .B(n7173), .Z(n7149) );
  XOR U11304 ( .A(n7163), .B(n7164), .Z(n7173) );
  XOR U11305 ( .A(n7169), .B(n7174), .Z(n7164) );
  XOR U11306 ( .A(n7168), .B(n7171), .Z(n7174) );
  IV U11307 ( .A(n7170), .Z(n7171) );
  NAND U11308 ( .A(n7175), .B(n7176), .Z(n7170) );
  OR U11309 ( .A(n7177), .B(n7178), .Z(n7176) );
  OR U11310 ( .A(n7179), .B(n7180), .Z(n7175) );
  NAND U11311 ( .A(n7181), .B(n7182), .Z(n7168) );
  OR U11312 ( .A(n7183), .B(n7184), .Z(n7182) );
  OR U11313 ( .A(n7185), .B(n7186), .Z(n7181) );
  NOR U11314 ( .A(n7187), .B(n7188), .Z(n7169) );
  ANDN U11315 ( .B(n7189), .A(n7190), .Z(n7163) );
  XNOR U11316 ( .A(n7156), .B(n7191), .Z(n7162) );
  XNOR U11317 ( .A(n7155), .B(n7157), .Z(n7191) );
  NAND U11318 ( .A(n7192), .B(n7193), .Z(n7157) );
  OR U11319 ( .A(n7194), .B(n7195), .Z(n7193) );
  OR U11320 ( .A(n7196), .B(n7197), .Z(n7192) );
  NAND U11321 ( .A(n7198), .B(n7199), .Z(n7155) );
  OR U11322 ( .A(n7200), .B(n7201), .Z(n7199) );
  OR U11323 ( .A(n7202), .B(n7203), .Z(n7198) );
  ANDN U11324 ( .B(n7204), .A(n7205), .Z(n7156) );
  IV U11325 ( .A(n7206), .Z(n7204) );
  ANDN U11326 ( .B(n7207), .A(n7208), .Z(n7148) );
  XOR U11327 ( .A(n7134), .B(n7209), .Z(n7146) );
  XOR U11328 ( .A(n7135), .B(n7136), .Z(n7209) );
  XOR U11329 ( .A(n7141), .B(n7210), .Z(n7136) );
  XOR U11330 ( .A(n7140), .B(n7143), .Z(n7210) );
  IV U11331 ( .A(n7142), .Z(n7143) );
  NAND U11332 ( .A(n7211), .B(n7212), .Z(n7142) );
  OR U11333 ( .A(n7213), .B(n7214), .Z(n7212) );
  OR U11334 ( .A(n7215), .B(n7216), .Z(n7211) );
  NAND U11335 ( .A(n7217), .B(n7218), .Z(n7140) );
  OR U11336 ( .A(n7219), .B(n7220), .Z(n7218) );
  OR U11337 ( .A(n7221), .B(n7222), .Z(n7217) );
  NOR U11338 ( .A(n7223), .B(n7224), .Z(n7141) );
  ANDN U11339 ( .B(n7225), .A(n7226), .Z(n7135) );
  IV U11340 ( .A(n7227), .Z(n7225) );
  XNOR U11341 ( .A(n7128), .B(n7228), .Z(n7134) );
  XNOR U11342 ( .A(n7127), .B(n7129), .Z(n7228) );
  NAND U11343 ( .A(n7229), .B(n7230), .Z(n7129) );
  OR U11344 ( .A(n7231), .B(n7232), .Z(n7230) );
  OR U11345 ( .A(n7233), .B(n7234), .Z(n7229) );
  NAND U11346 ( .A(n7235), .B(n7236), .Z(n7127) );
  OR U11347 ( .A(n7237), .B(n7238), .Z(n7236) );
  OR U11348 ( .A(n7239), .B(n7240), .Z(n7235) );
  ANDN U11349 ( .B(n7241), .A(n7242), .Z(n7128) );
  IV U11350 ( .A(n7243), .Z(n7241) );
  XNOR U11351 ( .A(n7208), .B(n7207), .Z(N29561) );
  XOR U11352 ( .A(n7227), .B(n7226), .Z(n7207) );
  XNOR U11353 ( .A(n7242), .B(n7243), .Z(n7226) );
  XNOR U11354 ( .A(n7237), .B(n7238), .Z(n7243) );
  XNOR U11355 ( .A(n7239), .B(n7240), .Z(n7238) );
  XNOR U11356 ( .A(y[3268]), .B(x[3268]), .Z(n7240) );
  XNOR U11357 ( .A(y[3269]), .B(x[3269]), .Z(n7239) );
  XNOR U11358 ( .A(y[3267]), .B(x[3267]), .Z(n7237) );
  XNOR U11359 ( .A(n7231), .B(n7232), .Z(n7242) );
  XNOR U11360 ( .A(y[3264]), .B(x[3264]), .Z(n7232) );
  XNOR U11361 ( .A(n7233), .B(n7234), .Z(n7231) );
  XNOR U11362 ( .A(y[3265]), .B(x[3265]), .Z(n7234) );
  XNOR U11363 ( .A(y[3266]), .B(x[3266]), .Z(n7233) );
  XNOR U11364 ( .A(n7224), .B(n7223), .Z(n7227) );
  XNOR U11365 ( .A(n7219), .B(n7220), .Z(n7223) );
  XNOR U11366 ( .A(y[3261]), .B(x[3261]), .Z(n7220) );
  XNOR U11367 ( .A(n7221), .B(n7222), .Z(n7219) );
  XNOR U11368 ( .A(y[3262]), .B(x[3262]), .Z(n7222) );
  XNOR U11369 ( .A(y[3263]), .B(x[3263]), .Z(n7221) );
  XNOR U11370 ( .A(n7213), .B(n7214), .Z(n7224) );
  XNOR U11371 ( .A(y[3258]), .B(x[3258]), .Z(n7214) );
  XNOR U11372 ( .A(n7215), .B(n7216), .Z(n7213) );
  XNOR U11373 ( .A(y[3259]), .B(x[3259]), .Z(n7216) );
  XNOR U11374 ( .A(y[3260]), .B(x[3260]), .Z(n7215) );
  XOR U11375 ( .A(n7189), .B(n7190), .Z(n7208) );
  XNOR U11376 ( .A(n7205), .B(n7206), .Z(n7190) );
  XNOR U11377 ( .A(n7200), .B(n7201), .Z(n7206) );
  XNOR U11378 ( .A(n7202), .B(n7203), .Z(n7201) );
  XNOR U11379 ( .A(y[3256]), .B(x[3256]), .Z(n7203) );
  XNOR U11380 ( .A(y[3257]), .B(x[3257]), .Z(n7202) );
  XNOR U11381 ( .A(y[3255]), .B(x[3255]), .Z(n7200) );
  XNOR U11382 ( .A(n7194), .B(n7195), .Z(n7205) );
  XNOR U11383 ( .A(y[3252]), .B(x[3252]), .Z(n7195) );
  XNOR U11384 ( .A(n7196), .B(n7197), .Z(n7194) );
  XNOR U11385 ( .A(y[3253]), .B(x[3253]), .Z(n7197) );
  XNOR U11386 ( .A(y[3254]), .B(x[3254]), .Z(n7196) );
  XOR U11387 ( .A(n7188), .B(n7187), .Z(n7189) );
  XNOR U11388 ( .A(n7183), .B(n7184), .Z(n7187) );
  XNOR U11389 ( .A(y[3249]), .B(x[3249]), .Z(n7184) );
  XNOR U11390 ( .A(n7185), .B(n7186), .Z(n7183) );
  XNOR U11391 ( .A(y[3250]), .B(x[3250]), .Z(n7186) );
  XNOR U11392 ( .A(y[3251]), .B(x[3251]), .Z(n7185) );
  XNOR U11393 ( .A(n7177), .B(n7178), .Z(n7188) );
  XNOR U11394 ( .A(y[3246]), .B(x[3246]), .Z(n7178) );
  XNOR U11395 ( .A(n7179), .B(n7180), .Z(n7177) );
  XNOR U11396 ( .A(y[3247]), .B(x[3247]), .Z(n7180) );
  XNOR U11397 ( .A(y[3248]), .B(x[3248]), .Z(n7179) );
  NAND U11398 ( .A(n7244), .B(n7245), .Z(N29553) );
  NANDN U11399 ( .A(n7246), .B(n7247), .Z(n7245) );
  OR U11400 ( .A(n7248), .B(n7249), .Z(n7247) );
  NAND U11401 ( .A(n7248), .B(n7249), .Z(n7244) );
  XOR U11402 ( .A(n7248), .B(n7250), .Z(N29552) );
  XNOR U11403 ( .A(n7246), .B(n7249), .Z(n7250) );
  AND U11404 ( .A(n7251), .B(n7252), .Z(n7249) );
  NANDN U11405 ( .A(n7253), .B(n7254), .Z(n7252) );
  NANDN U11406 ( .A(n7255), .B(n7256), .Z(n7254) );
  NANDN U11407 ( .A(n7256), .B(n7255), .Z(n7251) );
  NAND U11408 ( .A(n7257), .B(n7258), .Z(n7246) );
  NANDN U11409 ( .A(n7259), .B(n7260), .Z(n7258) );
  OR U11410 ( .A(n7261), .B(n7262), .Z(n7260) );
  NAND U11411 ( .A(n7262), .B(n7261), .Z(n7257) );
  AND U11412 ( .A(n7263), .B(n7264), .Z(n7248) );
  NANDN U11413 ( .A(n7265), .B(n7266), .Z(n7264) );
  NANDN U11414 ( .A(n7267), .B(n7268), .Z(n7266) );
  NANDN U11415 ( .A(n7268), .B(n7267), .Z(n7263) );
  XOR U11416 ( .A(n7262), .B(n7269), .Z(N29551) );
  XOR U11417 ( .A(n7259), .B(n7261), .Z(n7269) );
  XNOR U11418 ( .A(n7255), .B(n7270), .Z(n7261) );
  XNOR U11419 ( .A(n7253), .B(n7256), .Z(n7270) );
  NAND U11420 ( .A(n7271), .B(n7272), .Z(n7256) );
  NAND U11421 ( .A(n7273), .B(n7274), .Z(n7272) );
  OR U11422 ( .A(n7275), .B(n7276), .Z(n7273) );
  NANDN U11423 ( .A(n7277), .B(n7275), .Z(n7271) );
  IV U11424 ( .A(n7276), .Z(n7277) );
  NAND U11425 ( .A(n7278), .B(n7279), .Z(n7253) );
  NAND U11426 ( .A(n7280), .B(n7281), .Z(n7279) );
  NANDN U11427 ( .A(n7282), .B(n7283), .Z(n7280) );
  NANDN U11428 ( .A(n7283), .B(n7282), .Z(n7278) );
  AND U11429 ( .A(n7284), .B(n7285), .Z(n7255) );
  NAND U11430 ( .A(n7286), .B(n7287), .Z(n7285) );
  OR U11431 ( .A(n7288), .B(n7289), .Z(n7286) );
  NANDN U11432 ( .A(n7290), .B(n7288), .Z(n7284) );
  NAND U11433 ( .A(n7291), .B(n7292), .Z(n7259) );
  NANDN U11434 ( .A(n7293), .B(n7294), .Z(n7292) );
  OR U11435 ( .A(n7295), .B(n7296), .Z(n7294) );
  NANDN U11436 ( .A(n7297), .B(n7295), .Z(n7291) );
  IV U11437 ( .A(n7296), .Z(n7297) );
  XNOR U11438 ( .A(n7267), .B(n7298), .Z(n7262) );
  XNOR U11439 ( .A(n7265), .B(n7268), .Z(n7298) );
  NAND U11440 ( .A(n7299), .B(n7300), .Z(n7268) );
  NAND U11441 ( .A(n7301), .B(n7302), .Z(n7300) );
  OR U11442 ( .A(n7303), .B(n7304), .Z(n7301) );
  NANDN U11443 ( .A(n7305), .B(n7303), .Z(n7299) );
  IV U11444 ( .A(n7304), .Z(n7305) );
  NAND U11445 ( .A(n7306), .B(n7307), .Z(n7265) );
  NAND U11446 ( .A(n7308), .B(n7309), .Z(n7307) );
  NANDN U11447 ( .A(n7310), .B(n7311), .Z(n7308) );
  NANDN U11448 ( .A(n7311), .B(n7310), .Z(n7306) );
  AND U11449 ( .A(n7312), .B(n7313), .Z(n7267) );
  NAND U11450 ( .A(n7314), .B(n7315), .Z(n7313) );
  OR U11451 ( .A(n7316), .B(n7317), .Z(n7314) );
  NANDN U11452 ( .A(n7318), .B(n7316), .Z(n7312) );
  XNOR U11453 ( .A(n7293), .B(n7319), .Z(N29550) );
  XOR U11454 ( .A(n7295), .B(n7296), .Z(n7319) );
  XNOR U11455 ( .A(n7309), .B(n7320), .Z(n7296) );
  XOR U11456 ( .A(n7310), .B(n7311), .Z(n7320) );
  XOR U11457 ( .A(n7316), .B(n7321), .Z(n7311) );
  XOR U11458 ( .A(n7315), .B(n7318), .Z(n7321) );
  IV U11459 ( .A(n7317), .Z(n7318) );
  NAND U11460 ( .A(n7322), .B(n7323), .Z(n7317) );
  OR U11461 ( .A(n7324), .B(n7325), .Z(n7323) );
  OR U11462 ( .A(n7326), .B(n7327), .Z(n7322) );
  NAND U11463 ( .A(n7328), .B(n7329), .Z(n7315) );
  OR U11464 ( .A(n7330), .B(n7331), .Z(n7329) );
  OR U11465 ( .A(n7332), .B(n7333), .Z(n7328) );
  NOR U11466 ( .A(n7334), .B(n7335), .Z(n7316) );
  ANDN U11467 ( .B(n7336), .A(n7337), .Z(n7310) );
  XNOR U11468 ( .A(n7303), .B(n7338), .Z(n7309) );
  XNOR U11469 ( .A(n7302), .B(n7304), .Z(n7338) );
  NAND U11470 ( .A(n7339), .B(n7340), .Z(n7304) );
  OR U11471 ( .A(n7341), .B(n7342), .Z(n7340) );
  OR U11472 ( .A(n7343), .B(n7344), .Z(n7339) );
  NAND U11473 ( .A(n7345), .B(n7346), .Z(n7302) );
  OR U11474 ( .A(n7347), .B(n7348), .Z(n7346) );
  OR U11475 ( .A(n7349), .B(n7350), .Z(n7345) );
  ANDN U11476 ( .B(n7351), .A(n7352), .Z(n7303) );
  IV U11477 ( .A(n7353), .Z(n7351) );
  ANDN U11478 ( .B(n7354), .A(n7355), .Z(n7295) );
  XOR U11479 ( .A(n7281), .B(n7356), .Z(n7293) );
  XOR U11480 ( .A(n7282), .B(n7283), .Z(n7356) );
  XOR U11481 ( .A(n7288), .B(n7357), .Z(n7283) );
  XOR U11482 ( .A(n7287), .B(n7290), .Z(n7357) );
  IV U11483 ( .A(n7289), .Z(n7290) );
  NAND U11484 ( .A(n7358), .B(n7359), .Z(n7289) );
  OR U11485 ( .A(n7360), .B(n7361), .Z(n7359) );
  OR U11486 ( .A(n7362), .B(n7363), .Z(n7358) );
  NAND U11487 ( .A(n7364), .B(n7365), .Z(n7287) );
  OR U11488 ( .A(n7366), .B(n7367), .Z(n7365) );
  OR U11489 ( .A(n7368), .B(n7369), .Z(n7364) );
  NOR U11490 ( .A(n7370), .B(n7371), .Z(n7288) );
  ANDN U11491 ( .B(n7372), .A(n7373), .Z(n7282) );
  IV U11492 ( .A(n7374), .Z(n7372) );
  XNOR U11493 ( .A(n7275), .B(n7375), .Z(n7281) );
  XNOR U11494 ( .A(n7274), .B(n7276), .Z(n7375) );
  NAND U11495 ( .A(n7376), .B(n7377), .Z(n7276) );
  OR U11496 ( .A(n7378), .B(n7379), .Z(n7377) );
  OR U11497 ( .A(n7380), .B(n7381), .Z(n7376) );
  NAND U11498 ( .A(n7382), .B(n7383), .Z(n7274) );
  OR U11499 ( .A(n7384), .B(n7385), .Z(n7383) );
  OR U11500 ( .A(n7386), .B(n7387), .Z(n7382) );
  ANDN U11501 ( .B(n7388), .A(n7389), .Z(n7275) );
  IV U11502 ( .A(n7390), .Z(n7388) );
  XNOR U11503 ( .A(n7355), .B(n7354), .Z(N29549) );
  XOR U11504 ( .A(n7374), .B(n7373), .Z(n7354) );
  XNOR U11505 ( .A(n7389), .B(n7390), .Z(n7373) );
  XNOR U11506 ( .A(n7384), .B(n7385), .Z(n7390) );
  XNOR U11507 ( .A(n7386), .B(n7387), .Z(n7385) );
  XNOR U11508 ( .A(y[3244]), .B(x[3244]), .Z(n7387) );
  XNOR U11509 ( .A(y[3245]), .B(x[3245]), .Z(n7386) );
  XNOR U11510 ( .A(y[3243]), .B(x[3243]), .Z(n7384) );
  XNOR U11511 ( .A(n7378), .B(n7379), .Z(n7389) );
  XNOR U11512 ( .A(y[3240]), .B(x[3240]), .Z(n7379) );
  XNOR U11513 ( .A(n7380), .B(n7381), .Z(n7378) );
  XNOR U11514 ( .A(y[3241]), .B(x[3241]), .Z(n7381) );
  XNOR U11515 ( .A(y[3242]), .B(x[3242]), .Z(n7380) );
  XNOR U11516 ( .A(n7371), .B(n7370), .Z(n7374) );
  XNOR U11517 ( .A(n7366), .B(n7367), .Z(n7370) );
  XNOR U11518 ( .A(y[3237]), .B(x[3237]), .Z(n7367) );
  XNOR U11519 ( .A(n7368), .B(n7369), .Z(n7366) );
  XNOR U11520 ( .A(y[3238]), .B(x[3238]), .Z(n7369) );
  XNOR U11521 ( .A(y[3239]), .B(x[3239]), .Z(n7368) );
  XNOR U11522 ( .A(n7360), .B(n7361), .Z(n7371) );
  XNOR U11523 ( .A(y[3234]), .B(x[3234]), .Z(n7361) );
  XNOR U11524 ( .A(n7362), .B(n7363), .Z(n7360) );
  XNOR U11525 ( .A(y[3235]), .B(x[3235]), .Z(n7363) );
  XNOR U11526 ( .A(y[3236]), .B(x[3236]), .Z(n7362) );
  XOR U11527 ( .A(n7336), .B(n7337), .Z(n7355) );
  XNOR U11528 ( .A(n7352), .B(n7353), .Z(n7337) );
  XNOR U11529 ( .A(n7347), .B(n7348), .Z(n7353) );
  XNOR U11530 ( .A(n7349), .B(n7350), .Z(n7348) );
  XNOR U11531 ( .A(y[3232]), .B(x[3232]), .Z(n7350) );
  XNOR U11532 ( .A(y[3233]), .B(x[3233]), .Z(n7349) );
  XNOR U11533 ( .A(y[3231]), .B(x[3231]), .Z(n7347) );
  XNOR U11534 ( .A(n7341), .B(n7342), .Z(n7352) );
  XNOR U11535 ( .A(y[3228]), .B(x[3228]), .Z(n7342) );
  XNOR U11536 ( .A(n7343), .B(n7344), .Z(n7341) );
  XNOR U11537 ( .A(y[3229]), .B(x[3229]), .Z(n7344) );
  XNOR U11538 ( .A(y[3230]), .B(x[3230]), .Z(n7343) );
  XOR U11539 ( .A(n7335), .B(n7334), .Z(n7336) );
  XNOR U11540 ( .A(n7330), .B(n7331), .Z(n7334) );
  XNOR U11541 ( .A(y[3225]), .B(x[3225]), .Z(n7331) );
  XNOR U11542 ( .A(n7332), .B(n7333), .Z(n7330) );
  XNOR U11543 ( .A(y[3226]), .B(x[3226]), .Z(n7333) );
  XNOR U11544 ( .A(y[3227]), .B(x[3227]), .Z(n7332) );
  XNOR U11545 ( .A(n7324), .B(n7325), .Z(n7335) );
  XNOR U11546 ( .A(y[3222]), .B(x[3222]), .Z(n7325) );
  XNOR U11547 ( .A(n7326), .B(n7327), .Z(n7324) );
  XNOR U11548 ( .A(y[3223]), .B(x[3223]), .Z(n7327) );
  XNOR U11549 ( .A(y[3224]), .B(x[3224]), .Z(n7326) );
  NAND U11550 ( .A(n7391), .B(n7392), .Z(N29541) );
  NANDN U11551 ( .A(n7393), .B(n7394), .Z(n7392) );
  OR U11552 ( .A(n7395), .B(n7396), .Z(n7394) );
  NAND U11553 ( .A(n7395), .B(n7396), .Z(n7391) );
  XOR U11554 ( .A(n7395), .B(n7397), .Z(N29540) );
  XNOR U11555 ( .A(n7393), .B(n7396), .Z(n7397) );
  AND U11556 ( .A(n7398), .B(n7399), .Z(n7396) );
  NANDN U11557 ( .A(n7400), .B(n7401), .Z(n7399) );
  NANDN U11558 ( .A(n7402), .B(n7403), .Z(n7401) );
  NANDN U11559 ( .A(n7403), .B(n7402), .Z(n7398) );
  NAND U11560 ( .A(n7404), .B(n7405), .Z(n7393) );
  NANDN U11561 ( .A(n7406), .B(n7407), .Z(n7405) );
  OR U11562 ( .A(n7408), .B(n7409), .Z(n7407) );
  NAND U11563 ( .A(n7409), .B(n7408), .Z(n7404) );
  AND U11564 ( .A(n7410), .B(n7411), .Z(n7395) );
  NANDN U11565 ( .A(n7412), .B(n7413), .Z(n7411) );
  NANDN U11566 ( .A(n7414), .B(n7415), .Z(n7413) );
  NANDN U11567 ( .A(n7415), .B(n7414), .Z(n7410) );
  XOR U11568 ( .A(n7409), .B(n7416), .Z(N29539) );
  XOR U11569 ( .A(n7406), .B(n7408), .Z(n7416) );
  XNOR U11570 ( .A(n7402), .B(n7417), .Z(n7408) );
  XNOR U11571 ( .A(n7400), .B(n7403), .Z(n7417) );
  NAND U11572 ( .A(n7418), .B(n7419), .Z(n7403) );
  NAND U11573 ( .A(n7420), .B(n7421), .Z(n7419) );
  OR U11574 ( .A(n7422), .B(n7423), .Z(n7420) );
  NANDN U11575 ( .A(n7424), .B(n7422), .Z(n7418) );
  IV U11576 ( .A(n7423), .Z(n7424) );
  NAND U11577 ( .A(n7425), .B(n7426), .Z(n7400) );
  NAND U11578 ( .A(n7427), .B(n7428), .Z(n7426) );
  NANDN U11579 ( .A(n7429), .B(n7430), .Z(n7427) );
  NANDN U11580 ( .A(n7430), .B(n7429), .Z(n7425) );
  AND U11581 ( .A(n7431), .B(n7432), .Z(n7402) );
  NAND U11582 ( .A(n7433), .B(n7434), .Z(n7432) );
  OR U11583 ( .A(n7435), .B(n7436), .Z(n7433) );
  NANDN U11584 ( .A(n7437), .B(n7435), .Z(n7431) );
  NAND U11585 ( .A(n7438), .B(n7439), .Z(n7406) );
  NANDN U11586 ( .A(n7440), .B(n7441), .Z(n7439) );
  OR U11587 ( .A(n7442), .B(n7443), .Z(n7441) );
  NANDN U11588 ( .A(n7444), .B(n7442), .Z(n7438) );
  IV U11589 ( .A(n7443), .Z(n7444) );
  XNOR U11590 ( .A(n7414), .B(n7445), .Z(n7409) );
  XNOR U11591 ( .A(n7412), .B(n7415), .Z(n7445) );
  NAND U11592 ( .A(n7446), .B(n7447), .Z(n7415) );
  NAND U11593 ( .A(n7448), .B(n7449), .Z(n7447) );
  OR U11594 ( .A(n7450), .B(n7451), .Z(n7448) );
  NANDN U11595 ( .A(n7452), .B(n7450), .Z(n7446) );
  IV U11596 ( .A(n7451), .Z(n7452) );
  NAND U11597 ( .A(n7453), .B(n7454), .Z(n7412) );
  NAND U11598 ( .A(n7455), .B(n7456), .Z(n7454) );
  NANDN U11599 ( .A(n7457), .B(n7458), .Z(n7455) );
  NANDN U11600 ( .A(n7458), .B(n7457), .Z(n7453) );
  AND U11601 ( .A(n7459), .B(n7460), .Z(n7414) );
  NAND U11602 ( .A(n7461), .B(n7462), .Z(n7460) );
  OR U11603 ( .A(n7463), .B(n7464), .Z(n7461) );
  NANDN U11604 ( .A(n7465), .B(n7463), .Z(n7459) );
  XNOR U11605 ( .A(n7440), .B(n7466), .Z(N29538) );
  XOR U11606 ( .A(n7442), .B(n7443), .Z(n7466) );
  XNOR U11607 ( .A(n7456), .B(n7467), .Z(n7443) );
  XOR U11608 ( .A(n7457), .B(n7458), .Z(n7467) );
  XOR U11609 ( .A(n7463), .B(n7468), .Z(n7458) );
  XOR U11610 ( .A(n7462), .B(n7465), .Z(n7468) );
  IV U11611 ( .A(n7464), .Z(n7465) );
  NAND U11612 ( .A(n7469), .B(n7470), .Z(n7464) );
  OR U11613 ( .A(n7471), .B(n7472), .Z(n7470) );
  OR U11614 ( .A(n7473), .B(n7474), .Z(n7469) );
  NAND U11615 ( .A(n7475), .B(n7476), .Z(n7462) );
  OR U11616 ( .A(n7477), .B(n7478), .Z(n7476) );
  OR U11617 ( .A(n7479), .B(n7480), .Z(n7475) );
  NOR U11618 ( .A(n7481), .B(n7482), .Z(n7463) );
  ANDN U11619 ( .B(n7483), .A(n7484), .Z(n7457) );
  XNOR U11620 ( .A(n7450), .B(n7485), .Z(n7456) );
  XNOR U11621 ( .A(n7449), .B(n7451), .Z(n7485) );
  NAND U11622 ( .A(n7486), .B(n7487), .Z(n7451) );
  OR U11623 ( .A(n7488), .B(n7489), .Z(n7487) );
  OR U11624 ( .A(n7490), .B(n7491), .Z(n7486) );
  NAND U11625 ( .A(n7492), .B(n7493), .Z(n7449) );
  OR U11626 ( .A(n7494), .B(n7495), .Z(n7493) );
  OR U11627 ( .A(n7496), .B(n7497), .Z(n7492) );
  ANDN U11628 ( .B(n7498), .A(n7499), .Z(n7450) );
  IV U11629 ( .A(n7500), .Z(n7498) );
  ANDN U11630 ( .B(n7501), .A(n7502), .Z(n7442) );
  XOR U11631 ( .A(n7428), .B(n7503), .Z(n7440) );
  XOR U11632 ( .A(n7429), .B(n7430), .Z(n7503) );
  XOR U11633 ( .A(n7435), .B(n7504), .Z(n7430) );
  XOR U11634 ( .A(n7434), .B(n7437), .Z(n7504) );
  IV U11635 ( .A(n7436), .Z(n7437) );
  NAND U11636 ( .A(n7505), .B(n7506), .Z(n7436) );
  OR U11637 ( .A(n7507), .B(n7508), .Z(n7506) );
  OR U11638 ( .A(n7509), .B(n7510), .Z(n7505) );
  NAND U11639 ( .A(n7511), .B(n7512), .Z(n7434) );
  OR U11640 ( .A(n7513), .B(n7514), .Z(n7512) );
  OR U11641 ( .A(n7515), .B(n7516), .Z(n7511) );
  NOR U11642 ( .A(n7517), .B(n7518), .Z(n7435) );
  ANDN U11643 ( .B(n7519), .A(n7520), .Z(n7429) );
  IV U11644 ( .A(n7521), .Z(n7519) );
  XNOR U11645 ( .A(n7422), .B(n7522), .Z(n7428) );
  XNOR U11646 ( .A(n7421), .B(n7423), .Z(n7522) );
  NAND U11647 ( .A(n7523), .B(n7524), .Z(n7423) );
  OR U11648 ( .A(n7525), .B(n7526), .Z(n7524) );
  OR U11649 ( .A(n7527), .B(n7528), .Z(n7523) );
  NAND U11650 ( .A(n7529), .B(n7530), .Z(n7421) );
  OR U11651 ( .A(n7531), .B(n7532), .Z(n7530) );
  OR U11652 ( .A(n7533), .B(n7534), .Z(n7529) );
  ANDN U11653 ( .B(n7535), .A(n7536), .Z(n7422) );
  IV U11654 ( .A(n7537), .Z(n7535) );
  XNOR U11655 ( .A(n7502), .B(n7501), .Z(N29537) );
  XOR U11656 ( .A(n7521), .B(n7520), .Z(n7501) );
  XNOR U11657 ( .A(n7536), .B(n7537), .Z(n7520) );
  XNOR U11658 ( .A(n7531), .B(n7532), .Z(n7537) );
  XNOR U11659 ( .A(n7533), .B(n7534), .Z(n7532) );
  XNOR U11660 ( .A(y[3220]), .B(x[3220]), .Z(n7534) );
  XNOR U11661 ( .A(y[3221]), .B(x[3221]), .Z(n7533) );
  XNOR U11662 ( .A(y[3219]), .B(x[3219]), .Z(n7531) );
  XNOR U11663 ( .A(n7525), .B(n7526), .Z(n7536) );
  XNOR U11664 ( .A(y[3216]), .B(x[3216]), .Z(n7526) );
  XNOR U11665 ( .A(n7527), .B(n7528), .Z(n7525) );
  XNOR U11666 ( .A(y[3217]), .B(x[3217]), .Z(n7528) );
  XNOR U11667 ( .A(y[3218]), .B(x[3218]), .Z(n7527) );
  XNOR U11668 ( .A(n7518), .B(n7517), .Z(n7521) );
  XNOR U11669 ( .A(n7513), .B(n7514), .Z(n7517) );
  XNOR U11670 ( .A(y[3213]), .B(x[3213]), .Z(n7514) );
  XNOR U11671 ( .A(n7515), .B(n7516), .Z(n7513) );
  XNOR U11672 ( .A(y[3214]), .B(x[3214]), .Z(n7516) );
  XNOR U11673 ( .A(y[3215]), .B(x[3215]), .Z(n7515) );
  XNOR U11674 ( .A(n7507), .B(n7508), .Z(n7518) );
  XNOR U11675 ( .A(y[3210]), .B(x[3210]), .Z(n7508) );
  XNOR U11676 ( .A(n7509), .B(n7510), .Z(n7507) );
  XNOR U11677 ( .A(y[3211]), .B(x[3211]), .Z(n7510) );
  XNOR U11678 ( .A(y[3212]), .B(x[3212]), .Z(n7509) );
  XOR U11679 ( .A(n7483), .B(n7484), .Z(n7502) );
  XNOR U11680 ( .A(n7499), .B(n7500), .Z(n7484) );
  XNOR U11681 ( .A(n7494), .B(n7495), .Z(n7500) );
  XNOR U11682 ( .A(n7496), .B(n7497), .Z(n7495) );
  XNOR U11683 ( .A(y[3208]), .B(x[3208]), .Z(n7497) );
  XNOR U11684 ( .A(y[3209]), .B(x[3209]), .Z(n7496) );
  XNOR U11685 ( .A(y[3207]), .B(x[3207]), .Z(n7494) );
  XNOR U11686 ( .A(n7488), .B(n7489), .Z(n7499) );
  XNOR U11687 ( .A(y[3204]), .B(x[3204]), .Z(n7489) );
  XNOR U11688 ( .A(n7490), .B(n7491), .Z(n7488) );
  XNOR U11689 ( .A(y[3205]), .B(x[3205]), .Z(n7491) );
  XNOR U11690 ( .A(y[3206]), .B(x[3206]), .Z(n7490) );
  XOR U11691 ( .A(n7482), .B(n7481), .Z(n7483) );
  XNOR U11692 ( .A(n7477), .B(n7478), .Z(n7481) );
  XNOR U11693 ( .A(y[3201]), .B(x[3201]), .Z(n7478) );
  XNOR U11694 ( .A(n7479), .B(n7480), .Z(n7477) );
  XNOR U11695 ( .A(y[3202]), .B(x[3202]), .Z(n7480) );
  XNOR U11696 ( .A(y[3203]), .B(x[3203]), .Z(n7479) );
  XNOR U11697 ( .A(n7471), .B(n7472), .Z(n7482) );
  XNOR U11698 ( .A(y[3198]), .B(x[3198]), .Z(n7472) );
  XNOR U11699 ( .A(n7473), .B(n7474), .Z(n7471) );
  XNOR U11700 ( .A(y[3199]), .B(x[3199]), .Z(n7474) );
  XNOR U11701 ( .A(y[3200]), .B(x[3200]), .Z(n7473) );
  NAND U11702 ( .A(n7538), .B(n7539), .Z(N29529) );
  NANDN U11703 ( .A(n7540), .B(n7541), .Z(n7539) );
  OR U11704 ( .A(n7542), .B(n7543), .Z(n7541) );
  NAND U11705 ( .A(n7542), .B(n7543), .Z(n7538) );
  XOR U11706 ( .A(n7542), .B(n7544), .Z(N29528) );
  XNOR U11707 ( .A(n7540), .B(n7543), .Z(n7544) );
  AND U11708 ( .A(n7545), .B(n7546), .Z(n7543) );
  NANDN U11709 ( .A(n7547), .B(n7548), .Z(n7546) );
  NANDN U11710 ( .A(n7549), .B(n7550), .Z(n7548) );
  NANDN U11711 ( .A(n7550), .B(n7549), .Z(n7545) );
  NAND U11712 ( .A(n7551), .B(n7552), .Z(n7540) );
  NANDN U11713 ( .A(n7553), .B(n7554), .Z(n7552) );
  OR U11714 ( .A(n7555), .B(n7556), .Z(n7554) );
  NAND U11715 ( .A(n7556), .B(n7555), .Z(n7551) );
  AND U11716 ( .A(n7557), .B(n7558), .Z(n7542) );
  NANDN U11717 ( .A(n7559), .B(n7560), .Z(n7558) );
  NANDN U11718 ( .A(n7561), .B(n7562), .Z(n7560) );
  NANDN U11719 ( .A(n7562), .B(n7561), .Z(n7557) );
  XOR U11720 ( .A(n7556), .B(n7563), .Z(N29527) );
  XOR U11721 ( .A(n7553), .B(n7555), .Z(n7563) );
  XNOR U11722 ( .A(n7549), .B(n7564), .Z(n7555) );
  XNOR U11723 ( .A(n7547), .B(n7550), .Z(n7564) );
  NAND U11724 ( .A(n7565), .B(n7566), .Z(n7550) );
  NAND U11725 ( .A(n7567), .B(n7568), .Z(n7566) );
  OR U11726 ( .A(n7569), .B(n7570), .Z(n7567) );
  NANDN U11727 ( .A(n7571), .B(n7569), .Z(n7565) );
  IV U11728 ( .A(n7570), .Z(n7571) );
  NAND U11729 ( .A(n7572), .B(n7573), .Z(n7547) );
  NAND U11730 ( .A(n7574), .B(n7575), .Z(n7573) );
  NANDN U11731 ( .A(n7576), .B(n7577), .Z(n7574) );
  NANDN U11732 ( .A(n7577), .B(n7576), .Z(n7572) );
  AND U11733 ( .A(n7578), .B(n7579), .Z(n7549) );
  NAND U11734 ( .A(n7580), .B(n7581), .Z(n7579) );
  OR U11735 ( .A(n7582), .B(n7583), .Z(n7580) );
  NANDN U11736 ( .A(n7584), .B(n7582), .Z(n7578) );
  NAND U11737 ( .A(n7585), .B(n7586), .Z(n7553) );
  NANDN U11738 ( .A(n7587), .B(n7588), .Z(n7586) );
  OR U11739 ( .A(n7589), .B(n7590), .Z(n7588) );
  NANDN U11740 ( .A(n7591), .B(n7589), .Z(n7585) );
  IV U11741 ( .A(n7590), .Z(n7591) );
  XNOR U11742 ( .A(n7561), .B(n7592), .Z(n7556) );
  XNOR U11743 ( .A(n7559), .B(n7562), .Z(n7592) );
  NAND U11744 ( .A(n7593), .B(n7594), .Z(n7562) );
  NAND U11745 ( .A(n7595), .B(n7596), .Z(n7594) );
  OR U11746 ( .A(n7597), .B(n7598), .Z(n7595) );
  NANDN U11747 ( .A(n7599), .B(n7597), .Z(n7593) );
  IV U11748 ( .A(n7598), .Z(n7599) );
  NAND U11749 ( .A(n7600), .B(n7601), .Z(n7559) );
  NAND U11750 ( .A(n7602), .B(n7603), .Z(n7601) );
  NANDN U11751 ( .A(n7604), .B(n7605), .Z(n7602) );
  NANDN U11752 ( .A(n7605), .B(n7604), .Z(n7600) );
  AND U11753 ( .A(n7606), .B(n7607), .Z(n7561) );
  NAND U11754 ( .A(n7608), .B(n7609), .Z(n7607) );
  OR U11755 ( .A(n7610), .B(n7611), .Z(n7608) );
  NANDN U11756 ( .A(n7612), .B(n7610), .Z(n7606) );
  XNOR U11757 ( .A(n7587), .B(n7613), .Z(N29526) );
  XOR U11758 ( .A(n7589), .B(n7590), .Z(n7613) );
  XNOR U11759 ( .A(n7603), .B(n7614), .Z(n7590) );
  XOR U11760 ( .A(n7604), .B(n7605), .Z(n7614) );
  XOR U11761 ( .A(n7610), .B(n7615), .Z(n7605) );
  XOR U11762 ( .A(n7609), .B(n7612), .Z(n7615) );
  IV U11763 ( .A(n7611), .Z(n7612) );
  NAND U11764 ( .A(n7616), .B(n7617), .Z(n7611) );
  OR U11765 ( .A(n7618), .B(n7619), .Z(n7617) );
  OR U11766 ( .A(n7620), .B(n7621), .Z(n7616) );
  NAND U11767 ( .A(n7622), .B(n7623), .Z(n7609) );
  OR U11768 ( .A(n7624), .B(n7625), .Z(n7623) );
  OR U11769 ( .A(n7626), .B(n7627), .Z(n7622) );
  NOR U11770 ( .A(n7628), .B(n7629), .Z(n7610) );
  ANDN U11771 ( .B(n7630), .A(n7631), .Z(n7604) );
  XNOR U11772 ( .A(n7597), .B(n7632), .Z(n7603) );
  XNOR U11773 ( .A(n7596), .B(n7598), .Z(n7632) );
  NAND U11774 ( .A(n7633), .B(n7634), .Z(n7598) );
  OR U11775 ( .A(n7635), .B(n7636), .Z(n7634) );
  OR U11776 ( .A(n7637), .B(n7638), .Z(n7633) );
  NAND U11777 ( .A(n7639), .B(n7640), .Z(n7596) );
  OR U11778 ( .A(n7641), .B(n7642), .Z(n7640) );
  OR U11779 ( .A(n7643), .B(n7644), .Z(n7639) );
  ANDN U11780 ( .B(n7645), .A(n7646), .Z(n7597) );
  IV U11781 ( .A(n7647), .Z(n7645) );
  ANDN U11782 ( .B(n7648), .A(n7649), .Z(n7589) );
  XOR U11783 ( .A(n7575), .B(n7650), .Z(n7587) );
  XOR U11784 ( .A(n7576), .B(n7577), .Z(n7650) );
  XOR U11785 ( .A(n7582), .B(n7651), .Z(n7577) );
  XOR U11786 ( .A(n7581), .B(n7584), .Z(n7651) );
  IV U11787 ( .A(n7583), .Z(n7584) );
  NAND U11788 ( .A(n7652), .B(n7653), .Z(n7583) );
  OR U11789 ( .A(n7654), .B(n7655), .Z(n7653) );
  OR U11790 ( .A(n7656), .B(n7657), .Z(n7652) );
  NAND U11791 ( .A(n7658), .B(n7659), .Z(n7581) );
  OR U11792 ( .A(n7660), .B(n7661), .Z(n7659) );
  OR U11793 ( .A(n7662), .B(n7663), .Z(n7658) );
  NOR U11794 ( .A(n7664), .B(n7665), .Z(n7582) );
  ANDN U11795 ( .B(n7666), .A(n7667), .Z(n7576) );
  IV U11796 ( .A(n7668), .Z(n7666) );
  XNOR U11797 ( .A(n7569), .B(n7669), .Z(n7575) );
  XNOR U11798 ( .A(n7568), .B(n7570), .Z(n7669) );
  NAND U11799 ( .A(n7670), .B(n7671), .Z(n7570) );
  OR U11800 ( .A(n7672), .B(n7673), .Z(n7671) );
  OR U11801 ( .A(n7674), .B(n7675), .Z(n7670) );
  NAND U11802 ( .A(n7676), .B(n7677), .Z(n7568) );
  OR U11803 ( .A(n7678), .B(n7679), .Z(n7677) );
  OR U11804 ( .A(n7680), .B(n7681), .Z(n7676) );
  ANDN U11805 ( .B(n7682), .A(n7683), .Z(n7569) );
  IV U11806 ( .A(n7684), .Z(n7682) );
  XNOR U11807 ( .A(n7649), .B(n7648), .Z(N29525) );
  XOR U11808 ( .A(n7668), .B(n7667), .Z(n7648) );
  XNOR U11809 ( .A(n7683), .B(n7684), .Z(n7667) );
  XNOR U11810 ( .A(n7678), .B(n7679), .Z(n7684) );
  XNOR U11811 ( .A(n7680), .B(n7681), .Z(n7679) );
  XNOR U11812 ( .A(y[3196]), .B(x[3196]), .Z(n7681) );
  XNOR U11813 ( .A(y[3197]), .B(x[3197]), .Z(n7680) );
  XNOR U11814 ( .A(y[3195]), .B(x[3195]), .Z(n7678) );
  XNOR U11815 ( .A(n7672), .B(n7673), .Z(n7683) );
  XNOR U11816 ( .A(y[3192]), .B(x[3192]), .Z(n7673) );
  XNOR U11817 ( .A(n7674), .B(n7675), .Z(n7672) );
  XNOR U11818 ( .A(y[3193]), .B(x[3193]), .Z(n7675) );
  XNOR U11819 ( .A(y[3194]), .B(x[3194]), .Z(n7674) );
  XNOR U11820 ( .A(n7665), .B(n7664), .Z(n7668) );
  XNOR U11821 ( .A(n7660), .B(n7661), .Z(n7664) );
  XNOR U11822 ( .A(y[3189]), .B(x[3189]), .Z(n7661) );
  XNOR U11823 ( .A(n7662), .B(n7663), .Z(n7660) );
  XNOR U11824 ( .A(y[3190]), .B(x[3190]), .Z(n7663) );
  XNOR U11825 ( .A(y[3191]), .B(x[3191]), .Z(n7662) );
  XNOR U11826 ( .A(n7654), .B(n7655), .Z(n7665) );
  XNOR U11827 ( .A(y[3186]), .B(x[3186]), .Z(n7655) );
  XNOR U11828 ( .A(n7656), .B(n7657), .Z(n7654) );
  XNOR U11829 ( .A(y[3187]), .B(x[3187]), .Z(n7657) );
  XNOR U11830 ( .A(y[3188]), .B(x[3188]), .Z(n7656) );
  XOR U11831 ( .A(n7630), .B(n7631), .Z(n7649) );
  XNOR U11832 ( .A(n7646), .B(n7647), .Z(n7631) );
  XNOR U11833 ( .A(n7641), .B(n7642), .Z(n7647) );
  XNOR U11834 ( .A(n7643), .B(n7644), .Z(n7642) );
  XNOR U11835 ( .A(y[3184]), .B(x[3184]), .Z(n7644) );
  XNOR U11836 ( .A(y[3185]), .B(x[3185]), .Z(n7643) );
  XNOR U11837 ( .A(y[3183]), .B(x[3183]), .Z(n7641) );
  XNOR U11838 ( .A(n7635), .B(n7636), .Z(n7646) );
  XNOR U11839 ( .A(y[3180]), .B(x[3180]), .Z(n7636) );
  XNOR U11840 ( .A(n7637), .B(n7638), .Z(n7635) );
  XNOR U11841 ( .A(y[3181]), .B(x[3181]), .Z(n7638) );
  XNOR U11842 ( .A(y[3182]), .B(x[3182]), .Z(n7637) );
  XOR U11843 ( .A(n7629), .B(n7628), .Z(n7630) );
  XNOR U11844 ( .A(n7624), .B(n7625), .Z(n7628) );
  XNOR U11845 ( .A(y[3177]), .B(x[3177]), .Z(n7625) );
  XNOR U11846 ( .A(n7626), .B(n7627), .Z(n7624) );
  XNOR U11847 ( .A(y[3178]), .B(x[3178]), .Z(n7627) );
  XNOR U11848 ( .A(y[3179]), .B(x[3179]), .Z(n7626) );
  XNOR U11849 ( .A(n7618), .B(n7619), .Z(n7629) );
  XNOR U11850 ( .A(y[3174]), .B(x[3174]), .Z(n7619) );
  XNOR U11851 ( .A(n7620), .B(n7621), .Z(n7618) );
  XNOR U11852 ( .A(y[3175]), .B(x[3175]), .Z(n7621) );
  XNOR U11853 ( .A(y[3176]), .B(x[3176]), .Z(n7620) );
  NAND U11854 ( .A(n7685), .B(n7686), .Z(N29517) );
  NANDN U11855 ( .A(n7687), .B(n7688), .Z(n7686) );
  OR U11856 ( .A(n7689), .B(n7690), .Z(n7688) );
  NAND U11857 ( .A(n7689), .B(n7690), .Z(n7685) );
  XOR U11858 ( .A(n7689), .B(n7691), .Z(N29516) );
  XNOR U11859 ( .A(n7687), .B(n7690), .Z(n7691) );
  AND U11860 ( .A(n7692), .B(n7693), .Z(n7690) );
  NANDN U11861 ( .A(n7694), .B(n7695), .Z(n7693) );
  NANDN U11862 ( .A(n7696), .B(n7697), .Z(n7695) );
  NANDN U11863 ( .A(n7697), .B(n7696), .Z(n7692) );
  NAND U11864 ( .A(n7698), .B(n7699), .Z(n7687) );
  NANDN U11865 ( .A(n7700), .B(n7701), .Z(n7699) );
  OR U11866 ( .A(n7702), .B(n7703), .Z(n7701) );
  NAND U11867 ( .A(n7703), .B(n7702), .Z(n7698) );
  AND U11868 ( .A(n7704), .B(n7705), .Z(n7689) );
  NANDN U11869 ( .A(n7706), .B(n7707), .Z(n7705) );
  NANDN U11870 ( .A(n7708), .B(n7709), .Z(n7707) );
  NANDN U11871 ( .A(n7709), .B(n7708), .Z(n7704) );
  XOR U11872 ( .A(n7703), .B(n7710), .Z(N29515) );
  XOR U11873 ( .A(n7700), .B(n7702), .Z(n7710) );
  XNOR U11874 ( .A(n7696), .B(n7711), .Z(n7702) );
  XNOR U11875 ( .A(n7694), .B(n7697), .Z(n7711) );
  NAND U11876 ( .A(n7712), .B(n7713), .Z(n7697) );
  NAND U11877 ( .A(n7714), .B(n7715), .Z(n7713) );
  OR U11878 ( .A(n7716), .B(n7717), .Z(n7714) );
  NANDN U11879 ( .A(n7718), .B(n7716), .Z(n7712) );
  IV U11880 ( .A(n7717), .Z(n7718) );
  NAND U11881 ( .A(n7719), .B(n7720), .Z(n7694) );
  NAND U11882 ( .A(n7721), .B(n7722), .Z(n7720) );
  NANDN U11883 ( .A(n7723), .B(n7724), .Z(n7721) );
  NANDN U11884 ( .A(n7724), .B(n7723), .Z(n7719) );
  AND U11885 ( .A(n7725), .B(n7726), .Z(n7696) );
  NAND U11886 ( .A(n7727), .B(n7728), .Z(n7726) );
  OR U11887 ( .A(n7729), .B(n7730), .Z(n7727) );
  NANDN U11888 ( .A(n7731), .B(n7729), .Z(n7725) );
  NAND U11889 ( .A(n7732), .B(n7733), .Z(n7700) );
  NANDN U11890 ( .A(n7734), .B(n7735), .Z(n7733) );
  OR U11891 ( .A(n7736), .B(n7737), .Z(n7735) );
  NANDN U11892 ( .A(n7738), .B(n7736), .Z(n7732) );
  IV U11893 ( .A(n7737), .Z(n7738) );
  XNOR U11894 ( .A(n7708), .B(n7739), .Z(n7703) );
  XNOR U11895 ( .A(n7706), .B(n7709), .Z(n7739) );
  NAND U11896 ( .A(n7740), .B(n7741), .Z(n7709) );
  NAND U11897 ( .A(n7742), .B(n7743), .Z(n7741) );
  OR U11898 ( .A(n7744), .B(n7745), .Z(n7742) );
  NANDN U11899 ( .A(n7746), .B(n7744), .Z(n7740) );
  IV U11900 ( .A(n7745), .Z(n7746) );
  NAND U11901 ( .A(n7747), .B(n7748), .Z(n7706) );
  NAND U11902 ( .A(n7749), .B(n7750), .Z(n7748) );
  NANDN U11903 ( .A(n7751), .B(n7752), .Z(n7749) );
  NANDN U11904 ( .A(n7752), .B(n7751), .Z(n7747) );
  AND U11905 ( .A(n7753), .B(n7754), .Z(n7708) );
  NAND U11906 ( .A(n7755), .B(n7756), .Z(n7754) );
  OR U11907 ( .A(n7757), .B(n7758), .Z(n7755) );
  NANDN U11908 ( .A(n7759), .B(n7757), .Z(n7753) );
  XNOR U11909 ( .A(n7734), .B(n7760), .Z(N29514) );
  XOR U11910 ( .A(n7736), .B(n7737), .Z(n7760) );
  XNOR U11911 ( .A(n7750), .B(n7761), .Z(n7737) );
  XOR U11912 ( .A(n7751), .B(n7752), .Z(n7761) );
  XOR U11913 ( .A(n7757), .B(n7762), .Z(n7752) );
  XOR U11914 ( .A(n7756), .B(n7759), .Z(n7762) );
  IV U11915 ( .A(n7758), .Z(n7759) );
  NAND U11916 ( .A(n7763), .B(n7764), .Z(n7758) );
  OR U11917 ( .A(n7765), .B(n7766), .Z(n7764) );
  OR U11918 ( .A(n7767), .B(n7768), .Z(n7763) );
  NAND U11919 ( .A(n7769), .B(n7770), .Z(n7756) );
  OR U11920 ( .A(n7771), .B(n7772), .Z(n7770) );
  OR U11921 ( .A(n7773), .B(n7774), .Z(n7769) );
  NOR U11922 ( .A(n7775), .B(n7776), .Z(n7757) );
  ANDN U11923 ( .B(n7777), .A(n7778), .Z(n7751) );
  XNOR U11924 ( .A(n7744), .B(n7779), .Z(n7750) );
  XNOR U11925 ( .A(n7743), .B(n7745), .Z(n7779) );
  NAND U11926 ( .A(n7780), .B(n7781), .Z(n7745) );
  OR U11927 ( .A(n7782), .B(n7783), .Z(n7781) );
  OR U11928 ( .A(n7784), .B(n7785), .Z(n7780) );
  NAND U11929 ( .A(n7786), .B(n7787), .Z(n7743) );
  OR U11930 ( .A(n7788), .B(n7789), .Z(n7787) );
  OR U11931 ( .A(n7790), .B(n7791), .Z(n7786) );
  ANDN U11932 ( .B(n7792), .A(n7793), .Z(n7744) );
  IV U11933 ( .A(n7794), .Z(n7792) );
  ANDN U11934 ( .B(n7795), .A(n7796), .Z(n7736) );
  XOR U11935 ( .A(n7722), .B(n7797), .Z(n7734) );
  XOR U11936 ( .A(n7723), .B(n7724), .Z(n7797) );
  XOR U11937 ( .A(n7729), .B(n7798), .Z(n7724) );
  XOR U11938 ( .A(n7728), .B(n7731), .Z(n7798) );
  IV U11939 ( .A(n7730), .Z(n7731) );
  NAND U11940 ( .A(n7799), .B(n7800), .Z(n7730) );
  OR U11941 ( .A(n7801), .B(n7802), .Z(n7800) );
  OR U11942 ( .A(n7803), .B(n7804), .Z(n7799) );
  NAND U11943 ( .A(n7805), .B(n7806), .Z(n7728) );
  OR U11944 ( .A(n7807), .B(n7808), .Z(n7806) );
  OR U11945 ( .A(n7809), .B(n7810), .Z(n7805) );
  NOR U11946 ( .A(n7811), .B(n7812), .Z(n7729) );
  ANDN U11947 ( .B(n7813), .A(n7814), .Z(n7723) );
  IV U11948 ( .A(n7815), .Z(n7813) );
  XNOR U11949 ( .A(n7716), .B(n7816), .Z(n7722) );
  XNOR U11950 ( .A(n7715), .B(n7717), .Z(n7816) );
  NAND U11951 ( .A(n7817), .B(n7818), .Z(n7717) );
  OR U11952 ( .A(n7819), .B(n7820), .Z(n7818) );
  OR U11953 ( .A(n7821), .B(n7822), .Z(n7817) );
  NAND U11954 ( .A(n7823), .B(n7824), .Z(n7715) );
  OR U11955 ( .A(n7825), .B(n7826), .Z(n7824) );
  OR U11956 ( .A(n7827), .B(n7828), .Z(n7823) );
  ANDN U11957 ( .B(n7829), .A(n7830), .Z(n7716) );
  IV U11958 ( .A(n7831), .Z(n7829) );
  XNOR U11959 ( .A(n7796), .B(n7795), .Z(N29513) );
  XOR U11960 ( .A(n7815), .B(n7814), .Z(n7795) );
  XNOR U11961 ( .A(n7830), .B(n7831), .Z(n7814) );
  XNOR U11962 ( .A(n7825), .B(n7826), .Z(n7831) );
  XNOR U11963 ( .A(n7827), .B(n7828), .Z(n7826) );
  XNOR U11964 ( .A(y[3172]), .B(x[3172]), .Z(n7828) );
  XNOR U11965 ( .A(y[3173]), .B(x[3173]), .Z(n7827) );
  XNOR U11966 ( .A(y[3171]), .B(x[3171]), .Z(n7825) );
  XNOR U11967 ( .A(n7819), .B(n7820), .Z(n7830) );
  XNOR U11968 ( .A(y[3168]), .B(x[3168]), .Z(n7820) );
  XNOR U11969 ( .A(n7821), .B(n7822), .Z(n7819) );
  XNOR U11970 ( .A(y[3169]), .B(x[3169]), .Z(n7822) );
  XNOR U11971 ( .A(y[3170]), .B(x[3170]), .Z(n7821) );
  XNOR U11972 ( .A(n7812), .B(n7811), .Z(n7815) );
  XNOR U11973 ( .A(n7807), .B(n7808), .Z(n7811) );
  XNOR U11974 ( .A(y[3165]), .B(x[3165]), .Z(n7808) );
  XNOR U11975 ( .A(n7809), .B(n7810), .Z(n7807) );
  XNOR U11976 ( .A(y[3166]), .B(x[3166]), .Z(n7810) );
  XNOR U11977 ( .A(y[3167]), .B(x[3167]), .Z(n7809) );
  XNOR U11978 ( .A(n7801), .B(n7802), .Z(n7812) );
  XNOR U11979 ( .A(y[3162]), .B(x[3162]), .Z(n7802) );
  XNOR U11980 ( .A(n7803), .B(n7804), .Z(n7801) );
  XNOR U11981 ( .A(y[3163]), .B(x[3163]), .Z(n7804) );
  XNOR U11982 ( .A(y[3164]), .B(x[3164]), .Z(n7803) );
  XOR U11983 ( .A(n7777), .B(n7778), .Z(n7796) );
  XNOR U11984 ( .A(n7793), .B(n7794), .Z(n7778) );
  XNOR U11985 ( .A(n7788), .B(n7789), .Z(n7794) );
  XNOR U11986 ( .A(n7790), .B(n7791), .Z(n7789) );
  XNOR U11987 ( .A(y[3160]), .B(x[3160]), .Z(n7791) );
  XNOR U11988 ( .A(y[3161]), .B(x[3161]), .Z(n7790) );
  XNOR U11989 ( .A(y[3159]), .B(x[3159]), .Z(n7788) );
  XNOR U11990 ( .A(n7782), .B(n7783), .Z(n7793) );
  XNOR U11991 ( .A(y[3156]), .B(x[3156]), .Z(n7783) );
  XNOR U11992 ( .A(n7784), .B(n7785), .Z(n7782) );
  XNOR U11993 ( .A(y[3157]), .B(x[3157]), .Z(n7785) );
  XNOR U11994 ( .A(y[3158]), .B(x[3158]), .Z(n7784) );
  XOR U11995 ( .A(n7776), .B(n7775), .Z(n7777) );
  XNOR U11996 ( .A(n7771), .B(n7772), .Z(n7775) );
  XNOR U11997 ( .A(y[3153]), .B(x[3153]), .Z(n7772) );
  XNOR U11998 ( .A(n7773), .B(n7774), .Z(n7771) );
  XNOR U11999 ( .A(y[3154]), .B(x[3154]), .Z(n7774) );
  XNOR U12000 ( .A(y[3155]), .B(x[3155]), .Z(n7773) );
  XNOR U12001 ( .A(n7765), .B(n7766), .Z(n7776) );
  XNOR U12002 ( .A(y[3150]), .B(x[3150]), .Z(n7766) );
  XNOR U12003 ( .A(n7767), .B(n7768), .Z(n7765) );
  XNOR U12004 ( .A(y[3151]), .B(x[3151]), .Z(n7768) );
  XNOR U12005 ( .A(y[3152]), .B(x[3152]), .Z(n7767) );
  NAND U12006 ( .A(n7832), .B(n7833), .Z(N29505) );
  NANDN U12007 ( .A(n7834), .B(n7835), .Z(n7833) );
  OR U12008 ( .A(n7836), .B(n7837), .Z(n7835) );
  NAND U12009 ( .A(n7836), .B(n7837), .Z(n7832) );
  XOR U12010 ( .A(n7836), .B(n7838), .Z(N29504) );
  XNOR U12011 ( .A(n7834), .B(n7837), .Z(n7838) );
  AND U12012 ( .A(n7839), .B(n7840), .Z(n7837) );
  NANDN U12013 ( .A(n7841), .B(n7842), .Z(n7840) );
  NANDN U12014 ( .A(n7843), .B(n7844), .Z(n7842) );
  NANDN U12015 ( .A(n7844), .B(n7843), .Z(n7839) );
  NAND U12016 ( .A(n7845), .B(n7846), .Z(n7834) );
  NANDN U12017 ( .A(n7847), .B(n7848), .Z(n7846) );
  OR U12018 ( .A(n7849), .B(n7850), .Z(n7848) );
  NAND U12019 ( .A(n7850), .B(n7849), .Z(n7845) );
  AND U12020 ( .A(n7851), .B(n7852), .Z(n7836) );
  NANDN U12021 ( .A(n7853), .B(n7854), .Z(n7852) );
  NANDN U12022 ( .A(n7855), .B(n7856), .Z(n7854) );
  NANDN U12023 ( .A(n7856), .B(n7855), .Z(n7851) );
  XOR U12024 ( .A(n7850), .B(n7857), .Z(N29503) );
  XOR U12025 ( .A(n7847), .B(n7849), .Z(n7857) );
  XNOR U12026 ( .A(n7843), .B(n7858), .Z(n7849) );
  XNOR U12027 ( .A(n7841), .B(n7844), .Z(n7858) );
  NAND U12028 ( .A(n7859), .B(n7860), .Z(n7844) );
  NAND U12029 ( .A(n7861), .B(n7862), .Z(n7860) );
  OR U12030 ( .A(n7863), .B(n7864), .Z(n7861) );
  NANDN U12031 ( .A(n7865), .B(n7863), .Z(n7859) );
  IV U12032 ( .A(n7864), .Z(n7865) );
  NAND U12033 ( .A(n7866), .B(n7867), .Z(n7841) );
  NAND U12034 ( .A(n7868), .B(n7869), .Z(n7867) );
  NANDN U12035 ( .A(n7870), .B(n7871), .Z(n7868) );
  NANDN U12036 ( .A(n7871), .B(n7870), .Z(n7866) );
  AND U12037 ( .A(n7872), .B(n7873), .Z(n7843) );
  NAND U12038 ( .A(n7874), .B(n7875), .Z(n7873) );
  OR U12039 ( .A(n7876), .B(n7877), .Z(n7874) );
  NANDN U12040 ( .A(n7878), .B(n7876), .Z(n7872) );
  NAND U12041 ( .A(n7879), .B(n7880), .Z(n7847) );
  NANDN U12042 ( .A(n7881), .B(n7882), .Z(n7880) );
  OR U12043 ( .A(n7883), .B(n7884), .Z(n7882) );
  NANDN U12044 ( .A(n7885), .B(n7883), .Z(n7879) );
  IV U12045 ( .A(n7884), .Z(n7885) );
  XNOR U12046 ( .A(n7855), .B(n7886), .Z(n7850) );
  XNOR U12047 ( .A(n7853), .B(n7856), .Z(n7886) );
  NAND U12048 ( .A(n7887), .B(n7888), .Z(n7856) );
  NAND U12049 ( .A(n7889), .B(n7890), .Z(n7888) );
  OR U12050 ( .A(n7891), .B(n7892), .Z(n7889) );
  NANDN U12051 ( .A(n7893), .B(n7891), .Z(n7887) );
  IV U12052 ( .A(n7892), .Z(n7893) );
  NAND U12053 ( .A(n7894), .B(n7895), .Z(n7853) );
  NAND U12054 ( .A(n7896), .B(n7897), .Z(n7895) );
  NANDN U12055 ( .A(n7898), .B(n7899), .Z(n7896) );
  NANDN U12056 ( .A(n7899), .B(n7898), .Z(n7894) );
  AND U12057 ( .A(n7900), .B(n7901), .Z(n7855) );
  NAND U12058 ( .A(n7902), .B(n7903), .Z(n7901) );
  OR U12059 ( .A(n7904), .B(n7905), .Z(n7902) );
  NANDN U12060 ( .A(n7906), .B(n7904), .Z(n7900) );
  XNOR U12061 ( .A(n7881), .B(n7907), .Z(N29502) );
  XOR U12062 ( .A(n7883), .B(n7884), .Z(n7907) );
  XNOR U12063 ( .A(n7897), .B(n7908), .Z(n7884) );
  XOR U12064 ( .A(n7898), .B(n7899), .Z(n7908) );
  XOR U12065 ( .A(n7904), .B(n7909), .Z(n7899) );
  XOR U12066 ( .A(n7903), .B(n7906), .Z(n7909) );
  IV U12067 ( .A(n7905), .Z(n7906) );
  NAND U12068 ( .A(n7910), .B(n7911), .Z(n7905) );
  OR U12069 ( .A(n7912), .B(n7913), .Z(n7911) );
  OR U12070 ( .A(n7914), .B(n7915), .Z(n7910) );
  NAND U12071 ( .A(n7916), .B(n7917), .Z(n7903) );
  OR U12072 ( .A(n7918), .B(n7919), .Z(n7917) );
  OR U12073 ( .A(n7920), .B(n7921), .Z(n7916) );
  NOR U12074 ( .A(n7922), .B(n7923), .Z(n7904) );
  ANDN U12075 ( .B(n7924), .A(n7925), .Z(n7898) );
  XNOR U12076 ( .A(n7891), .B(n7926), .Z(n7897) );
  XNOR U12077 ( .A(n7890), .B(n7892), .Z(n7926) );
  NAND U12078 ( .A(n7927), .B(n7928), .Z(n7892) );
  OR U12079 ( .A(n7929), .B(n7930), .Z(n7928) );
  OR U12080 ( .A(n7931), .B(n7932), .Z(n7927) );
  NAND U12081 ( .A(n7933), .B(n7934), .Z(n7890) );
  OR U12082 ( .A(n7935), .B(n7936), .Z(n7934) );
  OR U12083 ( .A(n7937), .B(n7938), .Z(n7933) );
  ANDN U12084 ( .B(n7939), .A(n7940), .Z(n7891) );
  IV U12085 ( .A(n7941), .Z(n7939) );
  ANDN U12086 ( .B(n7942), .A(n7943), .Z(n7883) );
  XOR U12087 ( .A(n7869), .B(n7944), .Z(n7881) );
  XOR U12088 ( .A(n7870), .B(n7871), .Z(n7944) );
  XOR U12089 ( .A(n7876), .B(n7945), .Z(n7871) );
  XOR U12090 ( .A(n7875), .B(n7878), .Z(n7945) );
  IV U12091 ( .A(n7877), .Z(n7878) );
  NAND U12092 ( .A(n7946), .B(n7947), .Z(n7877) );
  OR U12093 ( .A(n7948), .B(n7949), .Z(n7947) );
  OR U12094 ( .A(n7950), .B(n7951), .Z(n7946) );
  NAND U12095 ( .A(n7952), .B(n7953), .Z(n7875) );
  OR U12096 ( .A(n7954), .B(n7955), .Z(n7953) );
  OR U12097 ( .A(n7956), .B(n7957), .Z(n7952) );
  NOR U12098 ( .A(n7958), .B(n7959), .Z(n7876) );
  ANDN U12099 ( .B(n7960), .A(n7961), .Z(n7870) );
  IV U12100 ( .A(n7962), .Z(n7960) );
  XNOR U12101 ( .A(n7863), .B(n7963), .Z(n7869) );
  XNOR U12102 ( .A(n7862), .B(n7864), .Z(n7963) );
  NAND U12103 ( .A(n7964), .B(n7965), .Z(n7864) );
  OR U12104 ( .A(n7966), .B(n7967), .Z(n7965) );
  OR U12105 ( .A(n7968), .B(n7969), .Z(n7964) );
  NAND U12106 ( .A(n7970), .B(n7971), .Z(n7862) );
  OR U12107 ( .A(n7972), .B(n7973), .Z(n7971) );
  OR U12108 ( .A(n7974), .B(n7975), .Z(n7970) );
  ANDN U12109 ( .B(n7976), .A(n7977), .Z(n7863) );
  IV U12110 ( .A(n7978), .Z(n7976) );
  XNOR U12111 ( .A(n7943), .B(n7942), .Z(N29501) );
  XOR U12112 ( .A(n7962), .B(n7961), .Z(n7942) );
  XNOR U12113 ( .A(n7977), .B(n7978), .Z(n7961) );
  XNOR U12114 ( .A(n7972), .B(n7973), .Z(n7978) );
  XNOR U12115 ( .A(n7974), .B(n7975), .Z(n7973) );
  XNOR U12116 ( .A(y[3148]), .B(x[3148]), .Z(n7975) );
  XNOR U12117 ( .A(y[3149]), .B(x[3149]), .Z(n7974) );
  XNOR U12118 ( .A(y[3147]), .B(x[3147]), .Z(n7972) );
  XNOR U12119 ( .A(n7966), .B(n7967), .Z(n7977) );
  XNOR U12120 ( .A(y[3144]), .B(x[3144]), .Z(n7967) );
  XNOR U12121 ( .A(n7968), .B(n7969), .Z(n7966) );
  XNOR U12122 ( .A(y[3145]), .B(x[3145]), .Z(n7969) );
  XNOR U12123 ( .A(y[3146]), .B(x[3146]), .Z(n7968) );
  XNOR U12124 ( .A(n7959), .B(n7958), .Z(n7962) );
  XNOR U12125 ( .A(n7954), .B(n7955), .Z(n7958) );
  XNOR U12126 ( .A(y[3141]), .B(x[3141]), .Z(n7955) );
  XNOR U12127 ( .A(n7956), .B(n7957), .Z(n7954) );
  XNOR U12128 ( .A(y[3142]), .B(x[3142]), .Z(n7957) );
  XNOR U12129 ( .A(y[3143]), .B(x[3143]), .Z(n7956) );
  XNOR U12130 ( .A(n7948), .B(n7949), .Z(n7959) );
  XNOR U12131 ( .A(y[3138]), .B(x[3138]), .Z(n7949) );
  XNOR U12132 ( .A(n7950), .B(n7951), .Z(n7948) );
  XNOR U12133 ( .A(y[3139]), .B(x[3139]), .Z(n7951) );
  XNOR U12134 ( .A(y[3140]), .B(x[3140]), .Z(n7950) );
  XOR U12135 ( .A(n7924), .B(n7925), .Z(n7943) );
  XNOR U12136 ( .A(n7940), .B(n7941), .Z(n7925) );
  XNOR U12137 ( .A(n7935), .B(n7936), .Z(n7941) );
  XNOR U12138 ( .A(n7937), .B(n7938), .Z(n7936) );
  XNOR U12139 ( .A(y[3136]), .B(x[3136]), .Z(n7938) );
  XNOR U12140 ( .A(y[3137]), .B(x[3137]), .Z(n7937) );
  XNOR U12141 ( .A(y[3135]), .B(x[3135]), .Z(n7935) );
  XNOR U12142 ( .A(n7929), .B(n7930), .Z(n7940) );
  XNOR U12143 ( .A(y[3132]), .B(x[3132]), .Z(n7930) );
  XNOR U12144 ( .A(n7931), .B(n7932), .Z(n7929) );
  XNOR U12145 ( .A(y[3133]), .B(x[3133]), .Z(n7932) );
  XNOR U12146 ( .A(y[3134]), .B(x[3134]), .Z(n7931) );
  XOR U12147 ( .A(n7923), .B(n7922), .Z(n7924) );
  XNOR U12148 ( .A(n7918), .B(n7919), .Z(n7922) );
  XNOR U12149 ( .A(y[3129]), .B(x[3129]), .Z(n7919) );
  XNOR U12150 ( .A(n7920), .B(n7921), .Z(n7918) );
  XNOR U12151 ( .A(y[3130]), .B(x[3130]), .Z(n7921) );
  XNOR U12152 ( .A(y[3131]), .B(x[3131]), .Z(n7920) );
  XNOR U12153 ( .A(n7912), .B(n7913), .Z(n7923) );
  XNOR U12154 ( .A(y[3126]), .B(x[3126]), .Z(n7913) );
  XNOR U12155 ( .A(n7914), .B(n7915), .Z(n7912) );
  XNOR U12156 ( .A(y[3127]), .B(x[3127]), .Z(n7915) );
  XNOR U12157 ( .A(y[3128]), .B(x[3128]), .Z(n7914) );
  NAND U12158 ( .A(n7979), .B(n7980), .Z(N29493) );
  NANDN U12159 ( .A(n7981), .B(n7982), .Z(n7980) );
  OR U12160 ( .A(n7983), .B(n7984), .Z(n7982) );
  NAND U12161 ( .A(n7983), .B(n7984), .Z(n7979) );
  XOR U12162 ( .A(n7983), .B(n7985), .Z(N29492) );
  XNOR U12163 ( .A(n7981), .B(n7984), .Z(n7985) );
  AND U12164 ( .A(n7986), .B(n7987), .Z(n7984) );
  NANDN U12165 ( .A(n7988), .B(n7989), .Z(n7987) );
  NANDN U12166 ( .A(n7990), .B(n7991), .Z(n7989) );
  NANDN U12167 ( .A(n7991), .B(n7990), .Z(n7986) );
  NAND U12168 ( .A(n7992), .B(n7993), .Z(n7981) );
  NANDN U12169 ( .A(n7994), .B(n7995), .Z(n7993) );
  OR U12170 ( .A(n7996), .B(n7997), .Z(n7995) );
  NAND U12171 ( .A(n7997), .B(n7996), .Z(n7992) );
  AND U12172 ( .A(n7998), .B(n7999), .Z(n7983) );
  NANDN U12173 ( .A(n8000), .B(n8001), .Z(n7999) );
  NANDN U12174 ( .A(n8002), .B(n8003), .Z(n8001) );
  NANDN U12175 ( .A(n8003), .B(n8002), .Z(n7998) );
  XOR U12176 ( .A(n7997), .B(n8004), .Z(N29491) );
  XOR U12177 ( .A(n7994), .B(n7996), .Z(n8004) );
  XNOR U12178 ( .A(n7990), .B(n8005), .Z(n7996) );
  XNOR U12179 ( .A(n7988), .B(n7991), .Z(n8005) );
  NAND U12180 ( .A(n8006), .B(n8007), .Z(n7991) );
  NAND U12181 ( .A(n8008), .B(n8009), .Z(n8007) );
  OR U12182 ( .A(n8010), .B(n8011), .Z(n8008) );
  NANDN U12183 ( .A(n8012), .B(n8010), .Z(n8006) );
  IV U12184 ( .A(n8011), .Z(n8012) );
  NAND U12185 ( .A(n8013), .B(n8014), .Z(n7988) );
  NAND U12186 ( .A(n8015), .B(n8016), .Z(n8014) );
  NANDN U12187 ( .A(n8017), .B(n8018), .Z(n8015) );
  NANDN U12188 ( .A(n8018), .B(n8017), .Z(n8013) );
  AND U12189 ( .A(n8019), .B(n8020), .Z(n7990) );
  NAND U12190 ( .A(n8021), .B(n8022), .Z(n8020) );
  OR U12191 ( .A(n8023), .B(n8024), .Z(n8021) );
  NANDN U12192 ( .A(n8025), .B(n8023), .Z(n8019) );
  NAND U12193 ( .A(n8026), .B(n8027), .Z(n7994) );
  NANDN U12194 ( .A(n8028), .B(n8029), .Z(n8027) );
  OR U12195 ( .A(n8030), .B(n8031), .Z(n8029) );
  NANDN U12196 ( .A(n8032), .B(n8030), .Z(n8026) );
  IV U12197 ( .A(n8031), .Z(n8032) );
  XNOR U12198 ( .A(n8002), .B(n8033), .Z(n7997) );
  XNOR U12199 ( .A(n8000), .B(n8003), .Z(n8033) );
  NAND U12200 ( .A(n8034), .B(n8035), .Z(n8003) );
  NAND U12201 ( .A(n8036), .B(n8037), .Z(n8035) );
  OR U12202 ( .A(n8038), .B(n8039), .Z(n8036) );
  NANDN U12203 ( .A(n8040), .B(n8038), .Z(n8034) );
  IV U12204 ( .A(n8039), .Z(n8040) );
  NAND U12205 ( .A(n8041), .B(n8042), .Z(n8000) );
  NAND U12206 ( .A(n8043), .B(n8044), .Z(n8042) );
  NANDN U12207 ( .A(n8045), .B(n8046), .Z(n8043) );
  NANDN U12208 ( .A(n8046), .B(n8045), .Z(n8041) );
  AND U12209 ( .A(n8047), .B(n8048), .Z(n8002) );
  NAND U12210 ( .A(n8049), .B(n8050), .Z(n8048) );
  OR U12211 ( .A(n8051), .B(n8052), .Z(n8049) );
  NANDN U12212 ( .A(n8053), .B(n8051), .Z(n8047) );
  XNOR U12213 ( .A(n8028), .B(n8054), .Z(N29490) );
  XOR U12214 ( .A(n8030), .B(n8031), .Z(n8054) );
  XNOR U12215 ( .A(n8044), .B(n8055), .Z(n8031) );
  XOR U12216 ( .A(n8045), .B(n8046), .Z(n8055) );
  XOR U12217 ( .A(n8051), .B(n8056), .Z(n8046) );
  XOR U12218 ( .A(n8050), .B(n8053), .Z(n8056) );
  IV U12219 ( .A(n8052), .Z(n8053) );
  NAND U12220 ( .A(n8057), .B(n8058), .Z(n8052) );
  OR U12221 ( .A(n8059), .B(n8060), .Z(n8058) );
  OR U12222 ( .A(n8061), .B(n8062), .Z(n8057) );
  NAND U12223 ( .A(n8063), .B(n8064), .Z(n8050) );
  OR U12224 ( .A(n8065), .B(n8066), .Z(n8064) );
  OR U12225 ( .A(n8067), .B(n8068), .Z(n8063) );
  NOR U12226 ( .A(n8069), .B(n8070), .Z(n8051) );
  ANDN U12227 ( .B(n8071), .A(n8072), .Z(n8045) );
  XNOR U12228 ( .A(n8038), .B(n8073), .Z(n8044) );
  XNOR U12229 ( .A(n8037), .B(n8039), .Z(n8073) );
  NAND U12230 ( .A(n8074), .B(n8075), .Z(n8039) );
  OR U12231 ( .A(n8076), .B(n8077), .Z(n8075) );
  OR U12232 ( .A(n8078), .B(n8079), .Z(n8074) );
  NAND U12233 ( .A(n8080), .B(n8081), .Z(n8037) );
  OR U12234 ( .A(n8082), .B(n8083), .Z(n8081) );
  OR U12235 ( .A(n8084), .B(n8085), .Z(n8080) );
  ANDN U12236 ( .B(n8086), .A(n8087), .Z(n8038) );
  IV U12237 ( .A(n8088), .Z(n8086) );
  ANDN U12238 ( .B(n8089), .A(n8090), .Z(n8030) );
  XOR U12239 ( .A(n8016), .B(n8091), .Z(n8028) );
  XOR U12240 ( .A(n8017), .B(n8018), .Z(n8091) );
  XOR U12241 ( .A(n8023), .B(n8092), .Z(n8018) );
  XOR U12242 ( .A(n8022), .B(n8025), .Z(n8092) );
  IV U12243 ( .A(n8024), .Z(n8025) );
  NAND U12244 ( .A(n8093), .B(n8094), .Z(n8024) );
  OR U12245 ( .A(n8095), .B(n8096), .Z(n8094) );
  OR U12246 ( .A(n8097), .B(n8098), .Z(n8093) );
  NAND U12247 ( .A(n8099), .B(n8100), .Z(n8022) );
  OR U12248 ( .A(n8101), .B(n8102), .Z(n8100) );
  OR U12249 ( .A(n8103), .B(n8104), .Z(n8099) );
  NOR U12250 ( .A(n8105), .B(n8106), .Z(n8023) );
  ANDN U12251 ( .B(n8107), .A(n8108), .Z(n8017) );
  IV U12252 ( .A(n8109), .Z(n8107) );
  XNOR U12253 ( .A(n8010), .B(n8110), .Z(n8016) );
  XNOR U12254 ( .A(n8009), .B(n8011), .Z(n8110) );
  NAND U12255 ( .A(n8111), .B(n8112), .Z(n8011) );
  OR U12256 ( .A(n8113), .B(n8114), .Z(n8112) );
  OR U12257 ( .A(n8115), .B(n8116), .Z(n8111) );
  NAND U12258 ( .A(n8117), .B(n8118), .Z(n8009) );
  OR U12259 ( .A(n8119), .B(n8120), .Z(n8118) );
  OR U12260 ( .A(n8121), .B(n8122), .Z(n8117) );
  ANDN U12261 ( .B(n8123), .A(n8124), .Z(n8010) );
  IV U12262 ( .A(n8125), .Z(n8123) );
  XNOR U12263 ( .A(n8090), .B(n8089), .Z(N29489) );
  XOR U12264 ( .A(n8109), .B(n8108), .Z(n8089) );
  XNOR U12265 ( .A(n8124), .B(n8125), .Z(n8108) );
  XNOR U12266 ( .A(n8119), .B(n8120), .Z(n8125) );
  XNOR U12267 ( .A(n8121), .B(n8122), .Z(n8120) );
  XNOR U12268 ( .A(y[3124]), .B(x[3124]), .Z(n8122) );
  XNOR U12269 ( .A(y[3125]), .B(x[3125]), .Z(n8121) );
  XNOR U12270 ( .A(y[3123]), .B(x[3123]), .Z(n8119) );
  XNOR U12271 ( .A(n8113), .B(n8114), .Z(n8124) );
  XNOR U12272 ( .A(y[3120]), .B(x[3120]), .Z(n8114) );
  XNOR U12273 ( .A(n8115), .B(n8116), .Z(n8113) );
  XNOR U12274 ( .A(y[3121]), .B(x[3121]), .Z(n8116) );
  XNOR U12275 ( .A(y[3122]), .B(x[3122]), .Z(n8115) );
  XNOR U12276 ( .A(n8106), .B(n8105), .Z(n8109) );
  XNOR U12277 ( .A(n8101), .B(n8102), .Z(n8105) );
  XNOR U12278 ( .A(y[3117]), .B(x[3117]), .Z(n8102) );
  XNOR U12279 ( .A(n8103), .B(n8104), .Z(n8101) );
  XNOR U12280 ( .A(y[3118]), .B(x[3118]), .Z(n8104) );
  XNOR U12281 ( .A(y[3119]), .B(x[3119]), .Z(n8103) );
  XNOR U12282 ( .A(n8095), .B(n8096), .Z(n8106) );
  XNOR U12283 ( .A(y[3114]), .B(x[3114]), .Z(n8096) );
  XNOR U12284 ( .A(n8097), .B(n8098), .Z(n8095) );
  XNOR U12285 ( .A(y[3115]), .B(x[3115]), .Z(n8098) );
  XNOR U12286 ( .A(y[3116]), .B(x[3116]), .Z(n8097) );
  XOR U12287 ( .A(n8071), .B(n8072), .Z(n8090) );
  XNOR U12288 ( .A(n8087), .B(n8088), .Z(n8072) );
  XNOR U12289 ( .A(n8082), .B(n8083), .Z(n8088) );
  XNOR U12290 ( .A(n8084), .B(n8085), .Z(n8083) );
  XNOR U12291 ( .A(y[3112]), .B(x[3112]), .Z(n8085) );
  XNOR U12292 ( .A(y[3113]), .B(x[3113]), .Z(n8084) );
  XNOR U12293 ( .A(y[3111]), .B(x[3111]), .Z(n8082) );
  XNOR U12294 ( .A(n8076), .B(n8077), .Z(n8087) );
  XNOR U12295 ( .A(y[3108]), .B(x[3108]), .Z(n8077) );
  XNOR U12296 ( .A(n8078), .B(n8079), .Z(n8076) );
  XNOR U12297 ( .A(y[3109]), .B(x[3109]), .Z(n8079) );
  XNOR U12298 ( .A(y[3110]), .B(x[3110]), .Z(n8078) );
  XOR U12299 ( .A(n8070), .B(n8069), .Z(n8071) );
  XNOR U12300 ( .A(n8065), .B(n8066), .Z(n8069) );
  XNOR U12301 ( .A(y[3105]), .B(x[3105]), .Z(n8066) );
  XNOR U12302 ( .A(n8067), .B(n8068), .Z(n8065) );
  XNOR U12303 ( .A(y[3106]), .B(x[3106]), .Z(n8068) );
  XNOR U12304 ( .A(y[3107]), .B(x[3107]), .Z(n8067) );
  XNOR U12305 ( .A(n8059), .B(n8060), .Z(n8070) );
  XNOR U12306 ( .A(y[3102]), .B(x[3102]), .Z(n8060) );
  XNOR U12307 ( .A(n8061), .B(n8062), .Z(n8059) );
  XNOR U12308 ( .A(y[3103]), .B(x[3103]), .Z(n8062) );
  XNOR U12309 ( .A(y[3104]), .B(x[3104]), .Z(n8061) );
  NAND U12310 ( .A(n8126), .B(n8127), .Z(N29481) );
  NANDN U12311 ( .A(n8128), .B(n8129), .Z(n8127) );
  OR U12312 ( .A(n8130), .B(n8131), .Z(n8129) );
  NAND U12313 ( .A(n8130), .B(n8131), .Z(n8126) );
  XOR U12314 ( .A(n8130), .B(n8132), .Z(N29480) );
  XNOR U12315 ( .A(n8128), .B(n8131), .Z(n8132) );
  AND U12316 ( .A(n8133), .B(n8134), .Z(n8131) );
  NANDN U12317 ( .A(n8135), .B(n8136), .Z(n8134) );
  NANDN U12318 ( .A(n8137), .B(n8138), .Z(n8136) );
  NANDN U12319 ( .A(n8138), .B(n8137), .Z(n8133) );
  NAND U12320 ( .A(n8139), .B(n8140), .Z(n8128) );
  NANDN U12321 ( .A(n8141), .B(n8142), .Z(n8140) );
  OR U12322 ( .A(n8143), .B(n8144), .Z(n8142) );
  NAND U12323 ( .A(n8144), .B(n8143), .Z(n8139) );
  AND U12324 ( .A(n8145), .B(n8146), .Z(n8130) );
  NANDN U12325 ( .A(n8147), .B(n8148), .Z(n8146) );
  NANDN U12326 ( .A(n8149), .B(n8150), .Z(n8148) );
  NANDN U12327 ( .A(n8150), .B(n8149), .Z(n8145) );
  XOR U12328 ( .A(n8144), .B(n8151), .Z(N29479) );
  XOR U12329 ( .A(n8141), .B(n8143), .Z(n8151) );
  XNOR U12330 ( .A(n8137), .B(n8152), .Z(n8143) );
  XNOR U12331 ( .A(n8135), .B(n8138), .Z(n8152) );
  NAND U12332 ( .A(n8153), .B(n8154), .Z(n8138) );
  NAND U12333 ( .A(n8155), .B(n8156), .Z(n8154) );
  OR U12334 ( .A(n8157), .B(n8158), .Z(n8155) );
  NANDN U12335 ( .A(n8159), .B(n8157), .Z(n8153) );
  IV U12336 ( .A(n8158), .Z(n8159) );
  NAND U12337 ( .A(n8160), .B(n8161), .Z(n8135) );
  NAND U12338 ( .A(n8162), .B(n8163), .Z(n8161) );
  NANDN U12339 ( .A(n8164), .B(n8165), .Z(n8162) );
  NANDN U12340 ( .A(n8165), .B(n8164), .Z(n8160) );
  AND U12341 ( .A(n8166), .B(n8167), .Z(n8137) );
  NAND U12342 ( .A(n8168), .B(n8169), .Z(n8167) );
  OR U12343 ( .A(n8170), .B(n8171), .Z(n8168) );
  NANDN U12344 ( .A(n8172), .B(n8170), .Z(n8166) );
  NAND U12345 ( .A(n8173), .B(n8174), .Z(n8141) );
  NANDN U12346 ( .A(n8175), .B(n8176), .Z(n8174) );
  OR U12347 ( .A(n8177), .B(n8178), .Z(n8176) );
  NANDN U12348 ( .A(n8179), .B(n8177), .Z(n8173) );
  IV U12349 ( .A(n8178), .Z(n8179) );
  XNOR U12350 ( .A(n8149), .B(n8180), .Z(n8144) );
  XNOR U12351 ( .A(n8147), .B(n8150), .Z(n8180) );
  NAND U12352 ( .A(n8181), .B(n8182), .Z(n8150) );
  NAND U12353 ( .A(n8183), .B(n8184), .Z(n8182) );
  OR U12354 ( .A(n8185), .B(n8186), .Z(n8183) );
  NANDN U12355 ( .A(n8187), .B(n8185), .Z(n8181) );
  IV U12356 ( .A(n8186), .Z(n8187) );
  NAND U12357 ( .A(n8188), .B(n8189), .Z(n8147) );
  NAND U12358 ( .A(n8190), .B(n8191), .Z(n8189) );
  NANDN U12359 ( .A(n8192), .B(n8193), .Z(n8190) );
  NANDN U12360 ( .A(n8193), .B(n8192), .Z(n8188) );
  AND U12361 ( .A(n8194), .B(n8195), .Z(n8149) );
  NAND U12362 ( .A(n8196), .B(n8197), .Z(n8195) );
  OR U12363 ( .A(n8198), .B(n8199), .Z(n8196) );
  NANDN U12364 ( .A(n8200), .B(n8198), .Z(n8194) );
  XNOR U12365 ( .A(n8175), .B(n8201), .Z(N29478) );
  XOR U12366 ( .A(n8177), .B(n8178), .Z(n8201) );
  XNOR U12367 ( .A(n8191), .B(n8202), .Z(n8178) );
  XOR U12368 ( .A(n8192), .B(n8193), .Z(n8202) );
  XOR U12369 ( .A(n8198), .B(n8203), .Z(n8193) );
  XOR U12370 ( .A(n8197), .B(n8200), .Z(n8203) );
  IV U12371 ( .A(n8199), .Z(n8200) );
  NAND U12372 ( .A(n8204), .B(n8205), .Z(n8199) );
  OR U12373 ( .A(n8206), .B(n8207), .Z(n8205) );
  OR U12374 ( .A(n8208), .B(n8209), .Z(n8204) );
  NAND U12375 ( .A(n8210), .B(n8211), .Z(n8197) );
  OR U12376 ( .A(n8212), .B(n8213), .Z(n8211) );
  OR U12377 ( .A(n8214), .B(n8215), .Z(n8210) );
  NOR U12378 ( .A(n8216), .B(n8217), .Z(n8198) );
  ANDN U12379 ( .B(n8218), .A(n8219), .Z(n8192) );
  XNOR U12380 ( .A(n8185), .B(n8220), .Z(n8191) );
  XNOR U12381 ( .A(n8184), .B(n8186), .Z(n8220) );
  NAND U12382 ( .A(n8221), .B(n8222), .Z(n8186) );
  OR U12383 ( .A(n8223), .B(n8224), .Z(n8222) );
  OR U12384 ( .A(n8225), .B(n8226), .Z(n8221) );
  NAND U12385 ( .A(n8227), .B(n8228), .Z(n8184) );
  OR U12386 ( .A(n8229), .B(n8230), .Z(n8228) );
  OR U12387 ( .A(n8231), .B(n8232), .Z(n8227) );
  ANDN U12388 ( .B(n8233), .A(n8234), .Z(n8185) );
  IV U12389 ( .A(n8235), .Z(n8233) );
  ANDN U12390 ( .B(n8236), .A(n8237), .Z(n8177) );
  XOR U12391 ( .A(n8163), .B(n8238), .Z(n8175) );
  XOR U12392 ( .A(n8164), .B(n8165), .Z(n8238) );
  XOR U12393 ( .A(n8170), .B(n8239), .Z(n8165) );
  XOR U12394 ( .A(n8169), .B(n8172), .Z(n8239) );
  IV U12395 ( .A(n8171), .Z(n8172) );
  NAND U12396 ( .A(n8240), .B(n8241), .Z(n8171) );
  OR U12397 ( .A(n8242), .B(n8243), .Z(n8241) );
  OR U12398 ( .A(n8244), .B(n8245), .Z(n8240) );
  NAND U12399 ( .A(n8246), .B(n8247), .Z(n8169) );
  OR U12400 ( .A(n8248), .B(n8249), .Z(n8247) );
  OR U12401 ( .A(n8250), .B(n8251), .Z(n8246) );
  NOR U12402 ( .A(n8252), .B(n8253), .Z(n8170) );
  ANDN U12403 ( .B(n8254), .A(n8255), .Z(n8164) );
  IV U12404 ( .A(n8256), .Z(n8254) );
  XNOR U12405 ( .A(n8157), .B(n8257), .Z(n8163) );
  XNOR U12406 ( .A(n8156), .B(n8158), .Z(n8257) );
  NAND U12407 ( .A(n8258), .B(n8259), .Z(n8158) );
  OR U12408 ( .A(n8260), .B(n8261), .Z(n8259) );
  OR U12409 ( .A(n8262), .B(n8263), .Z(n8258) );
  NAND U12410 ( .A(n8264), .B(n8265), .Z(n8156) );
  OR U12411 ( .A(n8266), .B(n8267), .Z(n8265) );
  OR U12412 ( .A(n8268), .B(n8269), .Z(n8264) );
  ANDN U12413 ( .B(n8270), .A(n8271), .Z(n8157) );
  IV U12414 ( .A(n8272), .Z(n8270) );
  XNOR U12415 ( .A(n8237), .B(n8236), .Z(N29477) );
  XOR U12416 ( .A(n8256), .B(n8255), .Z(n8236) );
  XNOR U12417 ( .A(n8271), .B(n8272), .Z(n8255) );
  XNOR U12418 ( .A(n8266), .B(n8267), .Z(n8272) );
  XNOR U12419 ( .A(n8268), .B(n8269), .Z(n8267) );
  XNOR U12420 ( .A(y[3100]), .B(x[3100]), .Z(n8269) );
  XNOR U12421 ( .A(y[3101]), .B(x[3101]), .Z(n8268) );
  XNOR U12422 ( .A(y[3099]), .B(x[3099]), .Z(n8266) );
  XNOR U12423 ( .A(n8260), .B(n8261), .Z(n8271) );
  XNOR U12424 ( .A(y[3096]), .B(x[3096]), .Z(n8261) );
  XNOR U12425 ( .A(n8262), .B(n8263), .Z(n8260) );
  XNOR U12426 ( .A(y[3097]), .B(x[3097]), .Z(n8263) );
  XNOR U12427 ( .A(y[3098]), .B(x[3098]), .Z(n8262) );
  XNOR U12428 ( .A(n8253), .B(n8252), .Z(n8256) );
  XNOR U12429 ( .A(n8248), .B(n8249), .Z(n8252) );
  XNOR U12430 ( .A(y[3093]), .B(x[3093]), .Z(n8249) );
  XNOR U12431 ( .A(n8250), .B(n8251), .Z(n8248) );
  XNOR U12432 ( .A(y[3094]), .B(x[3094]), .Z(n8251) );
  XNOR U12433 ( .A(y[3095]), .B(x[3095]), .Z(n8250) );
  XNOR U12434 ( .A(n8242), .B(n8243), .Z(n8253) );
  XNOR U12435 ( .A(y[3090]), .B(x[3090]), .Z(n8243) );
  XNOR U12436 ( .A(n8244), .B(n8245), .Z(n8242) );
  XNOR U12437 ( .A(y[3091]), .B(x[3091]), .Z(n8245) );
  XNOR U12438 ( .A(y[3092]), .B(x[3092]), .Z(n8244) );
  XOR U12439 ( .A(n8218), .B(n8219), .Z(n8237) );
  XNOR U12440 ( .A(n8234), .B(n8235), .Z(n8219) );
  XNOR U12441 ( .A(n8229), .B(n8230), .Z(n8235) );
  XNOR U12442 ( .A(n8231), .B(n8232), .Z(n8230) );
  XNOR U12443 ( .A(y[3088]), .B(x[3088]), .Z(n8232) );
  XNOR U12444 ( .A(y[3089]), .B(x[3089]), .Z(n8231) );
  XNOR U12445 ( .A(y[3087]), .B(x[3087]), .Z(n8229) );
  XNOR U12446 ( .A(n8223), .B(n8224), .Z(n8234) );
  XNOR U12447 ( .A(y[3084]), .B(x[3084]), .Z(n8224) );
  XNOR U12448 ( .A(n8225), .B(n8226), .Z(n8223) );
  XNOR U12449 ( .A(y[3085]), .B(x[3085]), .Z(n8226) );
  XNOR U12450 ( .A(y[3086]), .B(x[3086]), .Z(n8225) );
  XOR U12451 ( .A(n8217), .B(n8216), .Z(n8218) );
  XNOR U12452 ( .A(n8212), .B(n8213), .Z(n8216) );
  XNOR U12453 ( .A(y[3081]), .B(x[3081]), .Z(n8213) );
  XNOR U12454 ( .A(n8214), .B(n8215), .Z(n8212) );
  XNOR U12455 ( .A(y[3082]), .B(x[3082]), .Z(n8215) );
  XNOR U12456 ( .A(y[3083]), .B(x[3083]), .Z(n8214) );
  XNOR U12457 ( .A(n8206), .B(n8207), .Z(n8217) );
  XNOR U12458 ( .A(y[3078]), .B(x[3078]), .Z(n8207) );
  XNOR U12459 ( .A(n8208), .B(n8209), .Z(n8206) );
  XNOR U12460 ( .A(y[3079]), .B(x[3079]), .Z(n8209) );
  XNOR U12461 ( .A(y[3080]), .B(x[3080]), .Z(n8208) );
  NAND U12462 ( .A(n8273), .B(n8274), .Z(N29469) );
  NANDN U12463 ( .A(n8275), .B(n8276), .Z(n8274) );
  OR U12464 ( .A(n8277), .B(n8278), .Z(n8276) );
  NAND U12465 ( .A(n8277), .B(n8278), .Z(n8273) );
  XOR U12466 ( .A(n8277), .B(n8279), .Z(N29468) );
  XNOR U12467 ( .A(n8275), .B(n8278), .Z(n8279) );
  AND U12468 ( .A(n8280), .B(n8281), .Z(n8278) );
  NANDN U12469 ( .A(n8282), .B(n8283), .Z(n8281) );
  NANDN U12470 ( .A(n8284), .B(n8285), .Z(n8283) );
  NANDN U12471 ( .A(n8285), .B(n8284), .Z(n8280) );
  NAND U12472 ( .A(n8286), .B(n8287), .Z(n8275) );
  NANDN U12473 ( .A(n8288), .B(n8289), .Z(n8287) );
  OR U12474 ( .A(n8290), .B(n8291), .Z(n8289) );
  NAND U12475 ( .A(n8291), .B(n8290), .Z(n8286) );
  AND U12476 ( .A(n8292), .B(n8293), .Z(n8277) );
  NANDN U12477 ( .A(n8294), .B(n8295), .Z(n8293) );
  NANDN U12478 ( .A(n8296), .B(n8297), .Z(n8295) );
  NANDN U12479 ( .A(n8297), .B(n8296), .Z(n8292) );
  XOR U12480 ( .A(n8291), .B(n8298), .Z(N29467) );
  XOR U12481 ( .A(n8288), .B(n8290), .Z(n8298) );
  XNOR U12482 ( .A(n8284), .B(n8299), .Z(n8290) );
  XNOR U12483 ( .A(n8282), .B(n8285), .Z(n8299) );
  NAND U12484 ( .A(n8300), .B(n8301), .Z(n8285) );
  NAND U12485 ( .A(n8302), .B(n8303), .Z(n8301) );
  OR U12486 ( .A(n8304), .B(n8305), .Z(n8302) );
  NANDN U12487 ( .A(n8306), .B(n8304), .Z(n8300) );
  IV U12488 ( .A(n8305), .Z(n8306) );
  NAND U12489 ( .A(n8307), .B(n8308), .Z(n8282) );
  NAND U12490 ( .A(n8309), .B(n8310), .Z(n8308) );
  NANDN U12491 ( .A(n8311), .B(n8312), .Z(n8309) );
  NANDN U12492 ( .A(n8312), .B(n8311), .Z(n8307) );
  AND U12493 ( .A(n8313), .B(n8314), .Z(n8284) );
  NAND U12494 ( .A(n8315), .B(n8316), .Z(n8314) );
  OR U12495 ( .A(n8317), .B(n8318), .Z(n8315) );
  NANDN U12496 ( .A(n8319), .B(n8317), .Z(n8313) );
  NAND U12497 ( .A(n8320), .B(n8321), .Z(n8288) );
  NANDN U12498 ( .A(n8322), .B(n8323), .Z(n8321) );
  OR U12499 ( .A(n8324), .B(n8325), .Z(n8323) );
  NANDN U12500 ( .A(n8326), .B(n8324), .Z(n8320) );
  IV U12501 ( .A(n8325), .Z(n8326) );
  XNOR U12502 ( .A(n8296), .B(n8327), .Z(n8291) );
  XNOR U12503 ( .A(n8294), .B(n8297), .Z(n8327) );
  NAND U12504 ( .A(n8328), .B(n8329), .Z(n8297) );
  NAND U12505 ( .A(n8330), .B(n8331), .Z(n8329) );
  OR U12506 ( .A(n8332), .B(n8333), .Z(n8330) );
  NANDN U12507 ( .A(n8334), .B(n8332), .Z(n8328) );
  IV U12508 ( .A(n8333), .Z(n8334) );
  NAND U12509 ( .A(n8335), .B(n8336), .Z(n8294) );
  NAND U12510 ( .A(n8337), .B(n8338), .Z(n8336) );
  NANDN U12511 ( .A(n8339), .B(n8340), .Z(n8337) );
  NANDN U12512 ( .A(n8340), .B(n8339), .Z(n8335) );
  AND U12513 ( .A(n8341), .B(n8342), .Z(n8296) );
  NAND U12514 ( .A(n8343), .B(n8344), .Z(n8342) );
  OR U12515 ( .A(n8345), .B(n8346), .Z(n8343) );
  NANDN U12516 ( .A(n8347), .B(n8345), .Z(n8341) );
  XNOR U12517 ( .A(n8322), .B(n8348), .Z(N29466) );
  XOR U12518 ( .A(n8324), .B(n8325), .Z(n8348) );
  XNOR U12519 ( .A(n8338), .B(n8349), .Z(n8325) );
  XOR U12520 ( .A(n8339), .B(n8340), .Z(n8349) );
  XOR U12521 ( .A(n8345), .B(n8350), .Z(n8340) );
  XOR U12522 ( .A(n8344), .B(n8347), .Z(n8350) );
  IV U12523 ( .A(n8346), .Z(n8347) );
  NAND U12524 ( .A(n8351), .B(n8352), .Z(n8346) );
  OR U12525 ( .A(n8353), .B(n8354), .Z(n8352) );
  OR U12526 ( .A(n8355), .B(n8356), .Z(n8351) );
  NAND U12527 ( .A(n8357), .B(n8358), .Z(n8344) );
  OR U12528 ( .A(n8359), .B(n8360), .Z(n8358) );
  OR U12529 ( .A(n8361), .B(n8362), .Z(n8357) );
  NOR U12530 ( .A(n8363), .B(n8364), .Z(n8345) );
  ANDN U12531 ( .B(n8365), .A(n8366), .Z(n8339) );
  XNOR U12532 ( .A(n8332), .B(n8367), .Z(n8338) );
  XNOR U12533 ( .A(n8331), .B(n8333), .Z(n8367) );
  NAND U12534 ( .A(n8368), .B(n8369), .Z(n8333) );
  OR U12535 ( .A(n8370), .B(n8371), .Z(n8369) );
  OR U12536 ( .A(n8372), .B(n8373), .Z(n8368) );
  NAND U12537 ( .A(n8374), .B(n8375), .Z(n8331) );
  OR U12538 ( .A(n8376), .B(n8377), .Z(n8375) );
  OR U12539 ( .A(n8378), .B(n8379), .Z(n8374) );
  ANDN U12540 ( .B(n8380), .A(n8381), .Z(n8332) );
  IV U12541 ( .A(n8382), .Z(n8380) );
  ANDN U12542 ( .B(n8383), .A(n8384), .Z(n8324) );
  XOR U12543 ( .A(n8310), .B(n8385), .Z(n8322) );
  XOR U12544 ( .A(n8311), .B(n8312), .Z(n8385) );
  XOR U12545 ( .A(n8317), .B(n8386), .Z(n8312) );
  XOR U12546 ( .A(n8316), .B(n8319), .Z(n8386) );
  IV U12547 ( .A(n8318), .Z(n8319) );
  NAND U12548 ( .A(n8387), .B(n8388), .Z(n8318) );
  OR U12549 ( .A(n8389), .B(n8390), .Z(n8388) );
  OR U12550 ( .A(n8391), .B(n8392), .Z(n8387) );
  NAND U12551 ( .A(n8393), .B(n8394), .Z(n8316) );
  OR U12552 ( .A(n8395), .B(n8396), .Z(n8394) );
  OR U12553 ( .A(n8397), .B(n8398), .Z(n8393) );
  NOR U12554 ( .A(n8399), .B(n8400), .Z(n8317) );
  ANDN U12555 ( .B(n8401), .A(n8402), .Z(n8311) );
  IV U12556 ( .A(n8403), .Z(n8401) );
  XNOR U12557 ( .A(n8304), .B(n8404), .Z(n8310) );
  XNOR U12558 ( .A(n8303), .B(n8305), .Z(n8404) );
  NAND U12559 ( .A(n8405), .B(n8406), .Z(n8305) );
  OR U12560 ( .A(n8407), .B(n8408), .Z(n8406) );
  OR U12561 ( .A(n8409), .B(n8410), .Z(n8405) );
  NAND U12562 ( .A(n8411), .B(n8412), .Z(n8303) );
  OR U12563 ( .A(n8413), .B(n8414), .Z(n8412) );
  OR U12564 ( .A(n8415), .B(n8416), .Z(n8411) );
  ANDN U12565 ( .B(n8417), .A(n8418), .Z(n8304) );
  IV U12566 ( .A(n8419), .Z(n8417) );
  XNOR U12567 ( .A(n8384), .B(n8383), .Z(N29465) );
  XOR U12568 ( .A(n8403), .B(n8402), .Z(n8383) );
  XNOR U12569 ( .A(n8418), .B(n8419), .Z(n8402) );
  XNOR U12570 ( .A(n8413), .B(n8414), .Z(n8419) );
  XNOR U12571 ( .A(n8415), .B(n8416), .Z(n8414) );
  XNOR U12572 ( .A(y[3076]), .B(x[3076]), .Z(n8416) );
  XNOR U12573 ( .A(y[3077]), .B(x[3077]), .Z(n8415) );
  XNOR U12574 ( .A(y[3075]), .B(x[3075]), .Z(n8413) );
  XNOR U12575 ( .A(n8407), .B(n8408), .Z(n8418) );
  XNOR U12576 ( .A(y[3072]), .B(x[3072]), .Z(n8408) );
  XNOR U12577 ( .A(n8409), .B(n8410), .Z(n8407) );
  XNOR U12578 ( .A(y[3073]), .B(x[3073]), .Z(n8410) );
  XNOR U12579 ( .A(y[3074]), .B(x[3074]), .Z(n8409) );
  XNOR U12580 ( .A(n8400), .B(n8399), .Z(n8403) );
  XNOR U12581 ( .A(n8395), .B(n8396), .Z(n8399) );
  XNOR U12582 ( .A(y[3069]), .B(x[3069]), .Z(n8396) );
  XNOR U12583 ( .A(n8397), .B(n8398), .Z(n8395) );
  XNOR U12584 ( .A(y[3070]), .B(x[3070]), .Z(n8398) );
  XNOR U12585 ( .A(y[3071]), .B(x[3071]), .Z(n8397) );
  XNOR U12586 ( .A(n8389), .B(n8390), .Z(n8400) );
  XNOR U12587 ( .A(y[3066]), .B(x[3066]), .Z(n8390) );
  XNOR U12588 ( .A(n8391), .B(n8392), .Z(n8389) );
  XNOR U12589 ( .A(y[3067]), .B(x[3067]), .Z(n8392) );
  XNOR U12590 ( .A(y[3068]), .B(x[3068]), .Z(n8391) );
  XOR U12591 ( .A(n8365), .B(n8366), .Z(n8384) );
  XNOR U12592 ( .A(n8381), .B(n8382), .Z(n8366) );
  XNOR U12593 ( .A(n8376), .B(n8377), .Z(n8382) );
  XNOR U12594 ( .A(n8378), .B(n8379), .Z(n8377) );
  XNOR U12595 ( .A(y[3064]), .B(x[3064]), .Z(n8379) );
  XNOR U12596 ( .A(y[3065]), .B(x[3065]), .Z(n8378) );
  XNOR U12597 ( .A(y[3063]), .B(x[3063]), .Z(n8376) );
  XNOR U12598 ( .A(n8370), .B(n8371), .Z(n8381) );
  XNOR U12599 ( .A(y[3060]), .B(x[3060]), .Z(n8371) );
  XNOR U12600 ( .A(n8372), .B(n8373), .Z(n8370) );
  XNOR U12601 ( .A(y[3061]), .B(x[3061]), .Z(n8373) );
  XNOR U12602 ( .A(y[3062]), .B(x[3062]), .Z(n8372) );
  XOR U12603 ( .A(n8364), .B(n8363), .Z(n8365) );
  XNOR U12604 ( .A(n8359), .B(n8360), .Z(n8363) );
  XNOR U12605 ( .A(y[3057]), .B(x[3057]), .Z(n8360) );
  XNOR U12606 ( .A(n8361), .B(n8362), .Z(n8359) );
  XNOR U12607 ( .A(y[3058]), .B(x[3058]), .Z(n8362) );
  XNOR U12608 ( .A(y[3059]), .B(x[3059]), .Z(n8361) );
  XNOR U12609 ( .A(n8353), .B(n8354), .Z(n8364) );
  XNOR U12610 ( .A(y[3054]), .B(x[3054]), .Z(n8354) );
  XNOR U12611 ( .A(n8355), .B(n8356), .Z(n8353) );
  XNOR U12612 ( .A(y[3055]), .B(x[3055]), .Z(n8356) );
  XNOR U12613 ( .A(y[3056]), .B(x[3056]), .Z(n8355) );
  NAND U12614 ( .A(n8420), .B(n8421), .Z(N29457) );
  NANDN U12615 ( .A(n8422), .B(n8423), .Z(n8421) );
  OR U12616 ( .A(n8424), .B(n8425), .Z(n8423) );
  NAND U12617 ( .A(n8424), .B(n8425), .Z(n8420) );
  XOR U12618 ( .A(n8424), .B(n8426), .Z(N29456) );
  XNOR U12619 ( .A(n8422), .B(n8425), .Z(n8426) );
  AND U12620 ( .A(n8427), .B(n8428), .Z(n8425) );
  NANDN U12621 ( .A(n8429), .B(n8430), .Z(n8428) );
  NANDN U12622 ( .A(n8431), .B(n8432), .Z(n8430) );
  NANDN U12623 ( .A(n8432), .B(n8431), .Z(n8427) );
  NAND U12624 ( .A(n8433), .B(n8434), .Z(n8422) );
  NANDN U12625 ( .A(n8435), .B(n8436), .Z(n8434) );
  OR U12626 ( .A(n8437), .B(n8438), .Z(n8436) );
  NAND U12627 ( .A(n8438), .B(n8437), .Z(n8433) );
  AND U12628 ( .A(n8439), .B(n8440), .Z(n8424) );
  NANDN U12629 ( .A(n8441), .B(n8442), .Z(n8440) );
  NANDN U12630 ( .A(n8443), .B(n8444), .Z(n8442) );
  NANDN U12631 ( .A(n8444), .B(n8443), .Z(n8439) );
  XOR U12632 ( .A(n8438), .B(n8445), .Z(N29455) );
  XOR U12633 ( .A(n8435), .B(n8437), .Z(n8445) );
  XNOR U12634 ( .A(n8431), .B(n8446), .Z(n8437) );
  XNOR U12635 ( .A(n8429), .B(n8432), .Z(n8446) );
  NAND U12636 ( .A(n8447), .B(n8448), .Z(n8432) );
  NAND U12637 ( .A(n8449), .B(n8450), .Z(n8448) );
  OR U12638 ( .A(n8451), .B(n8452), .Z(n8449) );
  NANDN U12639 ( .A(n8453), .B(n8451), .Z(n8447) );
  IV U12640 ( .A(n8452), .Z(n8453) );
  NAND U12641 ( .A(n8454), .B(n8455), .Z(n8429) );
  NAND U12642 ( .A(n8456), .B(n8457), .Z(n8455) );
  NANDN U12643 ( .A(n8458), .B(n8459), .Z(n8456) );
  NANDN U12644 ( .A(n8459), .B(n8458), .Z(n8454) );
  AND U12645 ( .A(n8460), .B(n8461), .Z(n8431) );
  NAND U12646 ( .A(n8462), .B(n8463), .Z(n8461) );
  OR U12647 ( .A(n8464), .B(n8465), .Z(n8462) );
  NANDN U12648 ( .A(n8466), .B(n8464), .Z(n8460) );
  NAND U12649 ( .A(n8467), .B(n8468), .Z(n8435) );
  NANDN U12650 ( .A(n8469), .B(n8470), .Z(n8468) );
  OR U12651 ( .A(n8471), .B(n8472), .Z(n8470) );
  NANDN U12652 ( .A(n8473), .B(n8471), .Z(n8467) );
  IV U12653 ( .A(n8472), .Z(n8473) );
  XNOR U12654 ( .A(n8443), .B(n8474), .Z(n8438) );
  XNOR U12655 ( .A(n8441), .B(n8444), .Z(n8474) );
  NAND U12656 ( .A(n8475), .B(n8476), .Z(n8444) );
  NAND U12657 ( .A(n8477), .B(n8478), .Z(n8476) );
  OR U12658 ( .A(n8479), .B(n8480), .Z(n8477) );
  NANDN U12659 ( .A(n8481), .B(n8479), .Z(n8475) );
  IV U12660 ( .A(n8480), .Z(n8481) );
  NAND U12661 ( .A(n8482), .B(n8483), .Z(n8441) );
  NAND U12662 ( .A(n8484), .B(n8485), .Z(n8483) );
  NANDN U12663 ( .A(n8486), .B(n8487), .Z(n8484) );
  NANDN U12664 ( .A(n8487), .B(n8486), .Z(n8482) );
  AND U12665 ( .A(n8488), .B(n8489), .Z(n8443) );
  NAND U12666 ( .A(n8490), .B(n8491), .Z(n8489) );
  OR U12667 ( .A(n8492), .B(n8493), .Z(n8490) );
  NANDN U12668 ( .A(n8494), .B(n8492), .Z(n8488) );
  XNOR U12669 ( .A(n8469), .B(n8495), .Z(N29454) );
  XOR U12670 ( .A(n8471), .B(n8472), .Z(n8495) );
  XNOR U12671 ( .A(n8485), .B(n8496), .Z(n8472) );
  XOR U12672 ( .A(n8486), .B(n8487), .Z(n8496) );
  XOR U12673 ( .A(n8492), .B(n8497), .Z(n8487) );
  XOR U12674 ( .A(n8491), .B(n8494), .Z(n8497) );
  IV U12675 ( .A(n8493), .Z(n8494) );
  NAND U12676 ( .A(n8498), .B(n8499), .Z(n8493) );
  OR U12677 ( .A(n8500), .B(n8501), .Z(n8499) );
  OR U12678 ( .A(n8502), .B(n8503), .Z(n8498) );
  NAND U12679 ( .A(n8504), .B(n8505), .Z(n8491) );
  OR U12680 ( .A(n8506), .B(n8507), .Z(n8505) );
  OR U12681 ( .A(n8508), .B(n8509), .Z(n8504) );
  NOR U12682 ( .A(n8510), .B(n8511), .Z(n8492) );
  ANDN U12683 ( .B(n8512), .A(n8513), .Z(n8486) );
  XNOR U12684 ( .A(n8479), .B(n8514), .Z(n8485) );
  XNOR U12685 ( .A(n8478), .B(n8480), .Z(n8514) );
  NAND U12686 ( .A(n8515), .B(n8516), .Z(n8480) );
  OR U12687 ( .A(n8517), .B(n8518), .Z(n8516) );
  OR U12688 ( .A(n8519), .B(n8520), .Z(n8515) );
  NAND U12689 ( .A(n8521), .B(n8522), .Z(n8478) );
  OR U12690 ( .A(n8523), .B(n8524), .Z(n8522) );
  OR U12691 ( .A(n8525), .B(n8526), .Z(n8521) );
  ANDN U12692 ( .B(n8527), .A(n8528), .Z(n8479) );
  IV U12693 ( .A(n8529), .Z(n8527) );
  ANDN U12694 ( .B(n8530), .A(n8531), .Z(n8471) );
  XOR U12695 ( .A(n8457), .B(n8532), .Z(n8469) );
  XOR U12696 ( .A(n8458), .B(n8459), .Z(n8532) );
  XOR U12697 ( .A(n8464), .B(n8533), .Z(n8459) );
  XOR U12698 ( .A(n8463), .B(n8466), .Z(n8533) );
  IV U12699 ( .A(n8465), .Z(n8466) );
  NAND U12700 ( .A(n8534), .B(n8535), .Z(n8465) );
  OR U12701 ( .A(n8536), .B(n8537), .Z(n8535) );
  OR U12702 ( .A(n8538), .B(n8539), .Z(n8534) );
  NAND U12703 ( .A(n8540), .B(n8541), .Z(n8463) );
  OR U12704 ( .A(n8542), .B(n8543), .Z(n8541) );
  OR U12705 ( .A(n8544), .B(n8545), .Z(n8540) );
  NOR U12706 ( .A(n8546), .B(n8547), .Z(n8464) );
  ANDN U12707 ( .B(n8548), .A(n8549), .Z(n8458) );
  IV U12708 ( .A(n8550), .Z(n8548) );
  XNOR U12709 ( .A(n8451), .B(n8551), .Z(n8457) );
  XNOR U12710 ( .A(n8450), .B(n8452), .Z(n8551) );
  NAND U12711 ( .A(n8552), .B(n8553), .Z(n8452) );
  OR U12712 ( .A(n8554), .B(n8555), .Z(n8553) );
  OR U12713 ( .A(n8556), .B(n8557), .Z(n8552) );
  NAND U12714 ( .A(n8558), .B(n8559), .Z(n8450) );
  OR U12715 ( .A(n8560), .B(n8561), .Z(n8559) );
  OR U12716 ( .A(n8562), .B(n8563), .Z(n8558) );
  ANDN U12717 ( .B(n8564), .A(n8565), .Z(n8451) );
  IV U12718 ( .A(n8566), .Z(n8564) );
  XNOR U12719 ( .A(n8531), .B(n8530), .Z(N29453) );
  XOR U12720 ( .A(n8550), .B(n8549), .Z(n8530) );
  XNOR U12721 ( .A(n8565), .B(n8566), .Z(n8549) );
  XNOR U12722 ( .A(n8560), .B(n8561), .Z(n8566) );
  XNOR U12723 ( .A(n8562), .B(n8563), .Z(n8561) );
  XNOR U12724 ( .A(y[3052]), .B(x[3052]), .Z(n8563) );
  XNOR U12725 ( .A(y[3053]), .B(x[3053]), .Z(n8562) );
  XNOR U12726 ( .A(y[3051]), .B(x[3051]), .Z(n8560) );
  XNOR U12727 ( .A(n8554), .B(n8555), .Z(n8565) );
  XNOR U12728 ( .A(y[3048]), .B(x[3048]), .Z(n8555) );
  XNOR U12729 ( .A(n8556), .B(n8557), .Z(n8554) );
  XNOR U12730 ( .A(y[3049]), .B(x[3049]), .Z(n8557) );
  XNOR U12731 ( .A(y[3050]), .B(x[3050]), .Z(n8556) );
  XNOR U12732 ( .A(n8547), .B(n8546), .Z(n8550) );
  XNOR U12733 ( .A(n8542), .B(n8543), .Z(n8546) );
  XNOR U12734 ( .A(y[3045]), .B(x[3045]), .Z(n8543) );
  XNOR U12735 ( .A(n8544), .B(n8545), .Z(n8542) );
  XNOR U12736 ( .A(y[3046]), .B(x[3046]), .Z(n8545) );
  XNOR U12737 ( .A(y[3047]), .B(x[3047]), .Z(n8544) );
  XNOR U12738 ( .A(n8536), .B(n8537), .Z(n8547) );
  XNOR U12739 ( .A(y[3042]), .B(x[3042]), .Z(n8537) );
  XNOR U12740 ( .A(n8538), .B(n8539), .Z(n8536) );
  XNOR U12741 ( .A(y[3043]), .B(x[3043]), .Z(n8539) );
  XNOR U12742 ( .A(y[3044]), .B(x[3044]), .Z(n8538) );
  XOR U12743 ( .A(n8512), .B(n8513), .Z(n8531) );
  XNOR U12744 ( .A(n8528), .B(n8529), .Z(n8513) );
  XNOR U12745 ( .A(n8523), .B(n8524), .Z(n8529) );
  XNOR U12746 ( .A(n8525), .B(n8526), .Z(n8524) );
  XNOR U12747 ( .A(y[3040]), .B(x[3040]), .Z(n8526) );
  XNOR U12748 ( .A(y[3041]), .B(x[3041]), .Z(n8525) );
  XNOR U12749 ( .A(y[3039]), .B(x[3039]), .Z(n8523) );
  XNOR U12750 ( .A(n8517), .B(n8518), .Z(n8528) );
  XNOR U12751 ( .A(y[3036]), .B(x[3036]), .Z(n8518) );
  XNOR U12752 ( .A(n8519), .B(n8520), .Z(n8517) );
  XNOR U12753 ( .A(y[3037]), .B(x[3037]), .Z(n8520) );
  XNOR U12754 ( .A(y[3038]), .B(x[3038]), .Z(n8519) );
  XOR U12755 ( .A(n8511), .B(n8510), .Z(n8512) );
  XNOR U12756 ( .A(n8506), .B(n8507), .Z(n8510) );
  XNOR U12757 ( .A(y[3033]), .B(x[3033]), .Z(n8507) );
  XNOR U12758 ( .A(n8508), .B(n8509), .Z(n8506) );
  XNOR U12759 ( .A(y[3034]), .B(x[3034]), .Z(n8509) );
  XNOR U12760 ( .A(y[3035]), .B(x[3035]), .Z(n8508) );
  XNOR U12761 ( .A(n8500), .B(n8501), .Z(n8511) );
  XNOR U12762 ( .A(y[3030]), .B(x[3030]), .Z(n8501) );
  XNOR U12763 ( .A(n8502), .B(n8503), .Z(n8500) );
  XNOR U12764 ( .A(y[3031]), .B(x[3031]), .Z(n8503) );
  XNOR U12765 ( .A(y[3032]), .B(x[3032]), .Z(n8502) );
  NAND U12766 ( .A(n8567), .B(n8568), .Z(N29445) );
  NANDN U12767 ( .A(n8569), .B(n8570), .Z(n8568) );
  OR U12768 ( .A(n8571), .B(n8572), .Z(n8570) );
  NAND U12769 ( .A(n8571), .B(n8572), .Z(n8567) );
  XOR U12770 ( .A(n8571), .B(n8573), .Z(N29444) );
  XNOR U12771 ( .A(n8569), .B(n8572), .Z(n8573) );
  AND U12772 ( .A(n8574), .B(n8575), .Z(n8572) );
  NANDN U12773 ( .A(n8576), .B(n8577), .Z(n8575) );
  NANDN U12774 ( .A(n8578), .B(n8579), .Z(n8577) );
  NANDN U12775 ( .A(n8579), .B(n8578), .Z(n8574) );
  NAND U12776 ( .A(n8580), .B(n8581), .Z(n8569) );
  NANDN U12777 ( .A(n8582), .B(n8583), .Z(n8581) );
  OR U12778 ( .A(n8584), .B(n8585), .Z(n8583) );
  NAND U12779 ( .A(n8585), .B(n8584), .Z(n8580) );
  AND U12780 ( .A(n8586), .B(n8587), .Z(n8571) );
  NANDN U12781 ( .A(n8588), .B(n8589), .Z(n8587) );
  NANDN U12782 ( .A(n8590), .B(n8591), .Z(n8589) );
  NANDN U12783 ( .A(n8591), .B(n8590), .Z(n8586) );
  XOR U12784 ( .A(n8585), .B(n8592), .Z(N29443) );
  XOR U12785 ( .A(n8582), .B(n8584), .Z(n8592) );
  XNOR U12786 ( .A(n8578), .B(n8593), .Z(n8584) );
  XNOR U12787 ( .A(n8576), .B(n8579), .Z(n8593) );
  NAND U12788 ( .A(n8594), .B(n8595), .Z(n8579) );
  NAND U12789 ( .A(n8596), .B(n8597), .Z(n8595) );
  OR U12790 ( .A(n8598), .B(n8599), .Z(n8596) );
  NANDN U12791 ( .A(n8600), .B(n8598), .Z(n8594) );
  IV U12792 ( .A(n8599), .Z(n8600) );
  NAND U12793 ( .A(n8601), .B(n8602), .Z(n8576) );
  NAND U12794 ( .A(n8603), .B(n8604), .Z(n8602) );
  NANDN U12795 ( .A(n8605), .B(n8606), .Z(n8603) );
  NANDN U12796 ( .A(n8606), .B(n8605), .Z(n8601) );
  AND U12797 ( .A(n8607), .B(n8608), .Z(n8578) );
  NAND U12798 ( .A(n8609), .B(n8610), .Z(n8608) );
  OR U12799 ( .A(n8611), .B(n8612), .Z(n8609) );
  NANDN U12800 ( .A(n8613), .B(n8611), .Z(n8607) );
  NAND U12801 ( .A(n8614), .B(n8615), .Z(n8582) );
  NANDN U12802 ( .A(n8616), .B(n8617), .Z(n8615) );
  OR U12803 ( .A(n8618), .B(n8619), .Z(n8617) );
  NANDN U12804 ( .A(n8620), .B(n8618), .Z(n8614) );
  IV U12805 ( .A(n8619), .Z(n8620) );
  XNOR U12806 ( .A(n8590), .B(n8621), .Z(n8585) );
  XNOR U12807 ( .A(n8588), .B(n8591), .Z(n8621) );
  NAND U12808 ( .A(n8622), .B(n8623), .Z(n8591) );
  NAND U12809 ( .A(n8624), .B(n8625), .Z(n8623) );
  OR U12810 ( .A(n8626), .B(n8627), .Z(n8624) );
  NANDN U12811 ( .A(n8628), .B(n8626), .Z(n8622) );
  IV U12812 ( .A(n8627), .Z(n8628) );
  NAND U12813 ( .A(n8629), .B(n8630), .Z(n8588) );
  NAND U12814 ( .A(n8631), .B(n8632), .Z(n8630) );
  NANDN U12815 ( .A(n8633), .B(n8634), .Z(n8631) );
  NANDN U12816 ( .A(n8634), .B(n8633), .Z(n8629) );
  AND U12817 ( .A(n8635), .B(n8636), .Z(n8590) );
  NAND U12818 ( .A(n8637), .B(n8638), .Z(n8636) );
  OR U12819 ( .A(n8639), .B(n8640), .Z(n8637) );
  NANDN U12820 ( .A(n8641), .B(n8639), .Z(n8635) );
  XNOR U12821 ( .A(n8616), .B(n8642), .Z(N29442) );
  XOR U12822 ( .A(n8618), .B(n8619), .Z(n8642) );
  XNOR U12823 ( .A(n8632), .B(n8643), .Z(n8619) );
  XOR U12824 ( .A(n8633), .B(n8634), .Z(n8643) );
  XOR U12825 ( .A(n8639), .B(n8644), .Z(n8634) );
  XOR U12826 ( .A(n8638), .B(n8641), .Z(n8644) );
  IV U12827 ( .A(n8640), .Z(n8641) );
  NAND U12828 ( .A(n8645), .B(n8646), .Z(n8640) );
  OR U12829 ( .A(n8647), .B(n8648), .Z(n8646) );
  OR U12830 ( .A(n8649), .B(n8650), .Z(n8645) );
  NAND U12831 ( .A(n8651), .B(n8652), .Z(n8638) );
  OR U12832 ( .A(n8653), .B(n8654), .Z(n8652) );
  OR U12833 ( .A(n8655), .B(n8656), .Z(n8651) );
  NOR U12834 ( .A(n8657), .B(n8658), .Z(n8639) );
  ANDN U12835 ( .B(n8659), .A(n8660), .Z(n8633) );
  XNOR U12836 ( .A(n8626), .B(n8661), .Z(n8632) );
  XNOR U12837 ( .A(n8625), .B(n8627), .Z(n8661) );
  NAND U12838 ( .A(n8662), .B(n8663), .Z(n8627) );
  OR U12839 ( .A(n8664), .B(n8665), .Z(n8663) );
  OR U12840 ( .A(n8666), .B(n8667), .Z(n8662) );
  NAND U12841 ( .A(n8668), .B(n8669), .Z(n8625) );
  OR U12842 ( .A(n8670), .B(n8671), .Z(n8669) );
  OR U12843 ( .A(n8672), .B(n8673), .Z(n8668) );
  ANDN U12844 ( .B(n8674), .A(n8675), .Z(n8626) );
  IV U12845 ( .A(n8676), .Z(n8674) );
  ANDN U12846 ( .B(n8677), .A(n8678), .Z(n8618) );
  XOR U12847 ( .A(n8604), .B(n8679), .Z(n8616) );
  XOR U12848 ( .A(n8605), .B(n8606), .Z(n8679) );
  XOR U12849 ( .A(n8611), .B(n8680), .Z(n8606) );
  XOR U12850 ( .A(n8610), .B(n8613), .Z(n8680) );
  IV U12851 ( .A(n8612), .Z(n8613) );
  NAND U12852 ( .A(n8681), .B(n8682), .Z(n8612) );
  OR U12853 ( .A(n8683), .B(n8684), .Z(n8682) );
  OR U12854 ( .A(n8685), .B(n8686), .Z(n8681) );
  NAND U12855 ( .A(n8687), .B(n8688), .Z(n8610) );
  OR U12856 ( .A(n8689), .B(n8690), .Z(n8688) );
  OR U12857 ( .A(n8691), .B(n8692), .Z(n8687) );
  NOR U12858 ( .A(n8693), .B(n8694), .Z(n8611) );
  ANDN U12859 ( .B(n8695), .A(n8696), .Z(n8605) );
  IV U12860 ( .A(n8697), .Z(n8695) );
  XNOR U12861 ( .A(n8598), .B(n8698), .Z(n8604) );
  XNOR U12862 ( .A(n8597), .B(n8599), .Z(n8698) );
  NAND U12863 ( .A(n8699), .B(n8700), .Z(n8599) );
  OR U12864 ( .A(n8701), .B(n8702), .Z(n8700) );
  OR U12865 ( .A(n8703), .B(n8704), .Z(n8699) );
  NAND U12866 ( .A(n8705), .B(n8706), .Z(n8597) );
  OR U12867 ( .A(n8707), .B(n8708), .Z(n8706) );
  OR U12868 ( .A(n8709), .B(n8710), .Z(n8705) );
  ANDN U12869 ( .B(n8711), .A(n8712), .Z(n8598) );
  IV U12870 ( .A(n8713), .Z(n8711) );
  XNOR U12871 ( .A(n8678), .B(n8677), .Z(N29441) );
  XOR U12872 ( .A(n8697), .B(n8696), .Z(n8677) );
  XNOR U12873 ( .A(n8712), .B(n8713), .Z(n8696) );
  XNOR U12874 ( .A(n8707), .B(n8708), .Z(n8713) );
  XNOR U12875 ( .A(n8709), .B(n8710), .Z(n8708) );
  XNOR U12876 ( .A(y[3028]), .B(x[3028]), .Z(n8710) );
  XNOR U12877 ( .A(y[3029]), .B(x[3029]), .Z(n8709) );
  XNOR U12878 ( .A(y[3027]), .B(x[3027]), .Z(n8707) );
  XNOR U12879 ( .A(n8701), .B(n8702), .Z(n8712) );
  XNOR U12880 ( .A(y[3024]), .B(x[3024]), .Z(n8702) );
  XNOR U12881 ( .A(n8703), .B(n8704), .Z(n8701) );
  XNOR U12882 ( .A(y[3025]), .B(x[3025]), .Z(n8704) );
  XNOR U12883 ( .A(y[3026]), .B(x[3026]), .Z(n8703) );
  XNOR U12884 ( .A(n8694), .B(n8693), .Z(n8697) );
  XNOR U12885 ( .A(n8689), .B(n8690), .Z(n8693) );
  XNOR U12886 ( .A(y[3021]), .B(x[3021]), .Z(n8690) );
  XNOR U12887 ( .A(n8691), .B(n8692), .Z(n8689) );
  XNOR U12888 ( .A(y[3022]), .B(x[3022]), .Z(n8692) );
  XNOR U12889 ( .A(y[3023]), .B(x[3023]), .Z(n8691) );
  XNOR U12890 ( .A(n8683), .B(n8684), .Z(n8694) );
  XNOR U12891 ( .A(y[3018]), .B(x[3018]), .Z(n8684) );
  XNOR U12892 ( .A(n8685), .B(n8686), .Z(n8683) );
  XNOR U12893 ( .A(y[3019]), .B(x[3019]), .Z(n8686) );
  XNOR U12894 ( .A(y[3020]), .B(x[3020]), .Z(n8685) );
  XOR U12895 ( .A(n8659), .B(n8660), .Z(n8678) );
  XNOR U12896 ( .A(n8675), .B(n8676), .Z(n8660) );
  XNOR U12897 ( .A(n8670), .B(n8671), .Z(n8676) );
  XNOR U12898 ( .A(n8672), .B(n8673), .Z(n8671) );
  XNOR U12899 ( .A(y[3016]), .B(x[3016]), .Z(n8673) );
  XNOR U12900 ( .A(y[3017]), .B(x[3017]), .Z(n8672) );
  XNOR U12901 ( .A(y[3015]), .B(x[3015]), .Z(n8670) );
  XNOR U12902 ( .A(n8664), .B(n8665), .Z(n8675) );
  XNOR U12903 ( .A(y[3012]), .B(x[3012]), .Z(n8665) );
  XNOR U12904 ( .A(n8666), .B(n8667), .Z(n8664) );
  XNOR U12905 ( .A(y[3013]), .B(x[3013]), .Z(n8667) );
  XNOR U12906 ( .A(y[3014]), .B(x[3014]), .Z(n8666) );
  XOR U12907 ( .A(n8658), .B(n8657), .Z(n8659) );
  XNOR U12908 ( .A(n8653), .B(n8654), .Z(n8657) );
  XNOR U12909 ( .A(y[3009]), .B(x[3009]), .Z(n8654) );
  XNOR U12910 ( .A(n8655), .B(n8656), .Z(n8653) );
  XNOR U12911 ( .A(y[3010]), .B(x[3010]), .Z(n8656) );
  XNOR U12912 ( .A(y[3011]), .B(x[3011]), .Z(n8655) );
  XNOR U12913 ( .A(n8647), .B(n8648), .Z(n8658) );
  XNOR U12914 ( .A(y[3006]), .B(x[3006]), .Z(n8648) );
  XNOR U12915 ( .A(n8649), .B(n8650), .Z(n8647) );
  XNOR U12916 ( .A(y[3007]), .B(x[3007]), .Z(n8650) );
  XNOR U12917 ( .A(y[3008]), .B(x[3008]), .Z(n8649) );
  NAND U12918 ( .A(n8714), .B(n8715), .Z(N29433) );
  NANDN U12919 ( .A(n8716), .B(n8717), .Z(n8715) );
  OR U12920 ( .A(n8718), .B(n8719), .Z(n8717) );
  NAND U12921 ( .A(n8718), .B(n8719), .Z(n8714) );
  XOR U12922 ( .A(n8718), .B(n8720), .Z(N29432) );
  XNOR U12923 ( .A(n8716), .B(n8719), .Z(n8720) );
  AND U12924 ( .A(n8721), .B(n8722), .Z(n8719) );
  NANDN U12925 ( .A(n8723), .B(n8724), .Z(n8722) );
  NANDN U12926 ( .A(n8725), .B(n8726), .Z(n8724) );
  NANDN U12927 ( .A(n8726), .B(n8725), .Z(n8721) );
  NAND U12928 ( .A(n8727), .B(n8728), .Z(n8716) );
  NANDN U12929 ( .A(n8729), .B(n8730), .Z(n8728) );
  OR U12930 ( .A(n8731), .B(n8732), .Z(n8730) );
  NAND U12931 ( .A(n8732), .B(n8731), .Z(n8727) );
  AND U12932 ( .A(n8733), .B(n8734), .Z(n8718) );
  NANDN U12933 ( .A(n8735), .B(n8736), .Z(n8734) );
  NANDN U12934 ( .A(n8737), .B(n8738), .Z(n8736) );
  NANDN U12935 ( .A(n8738), .B(n8737), .Z(n8733) );
  XOR U12936 ( .A(n8732), .B(n8739), .Z(N29431) );
  XOR U12937 ( .A(n8729), .B(n8731), .Z(n8739) );
  XNOR U12938 ( .A(n8725), .B(n8740), .Z(n8731) );
  XNOR U12939 ( .A(n8723), .B(n8726), .Z(n8740) );
  NAND U12940 ( .A(n8741), .B(n8742), .Z(n8726) );
  NAND U12941 ( .A(n8743), .B(n8744), .Z(n8742) );
  OR U12942 ( .A(n8745), .B(n8746), .Z(n8743) );
  NANDN U12943 ( .A(n8747), .B(n8745), .Z(n8741) );
  IV U12944 ( .A(n8746), .Z(n8747) );
  NAND U12945 ( .A(n8748), .B(n8749), .Z(n8723) );
  NAND U12946 ( .A(n8750), .B(n8751), .Z(n8749) );
  NANDN U12947 ( .A(n8752), .B(n8753), .Z(n8750) );
  NANDN U12948 ( .A(n8753), .B(n8752), .Z(n8748) );
  AND U12949 ( .A(n8754), .B(n8755), .Z(n8725) );
  NAND U12950 ( .A(n8756), .B(n8757), .Z(n8755) );
  OR U12951 ( .A(n8758), .B(n8759), .Z(n8756) );
  NANDN U12952 ( .A(n8760), .B(n8758), .Z(n8754) );
  NAND U12953 ( .A(n8761), .B(n8762), .Z(n8729) );
  NANDN U12954 ( .A(n8763), .B(n8764), .Z(n8762) );
  OR U12955 ( .A(n8765), .B(n8766), .Z(n8764) );
  NANDN U12956 ( .A(n8767), .B(n8765), .Z(n8761) );
  IV U12957 ( .A(n8766), .Z(n8767) );
  XNOR U12958 ( .A(n8737), .B(n8768), .Z(n8732) );
  XNOR U12959 ( .A(n8735), .B(n8738), .Z(n8768) );
  NAND U12960 ( .A(n8769), .B(n8770), .Z(n8738) );
  NAND U12961 ( .A(n8771), .B(n8772), .Z(n8770) );
  OR U12962 ( .A(n8773), .B(n8774), .Z(n8771) );
  NANDN U12963 ( .A(n8775), .B(n8773), .Z(n8769) );
  IV U12964 ( .A(n8774), .Z(n8775) );
  NAND U12965 ( .A(n8776), .B(n8777), .Z(n8735) );
  NAND U12966 ( .A(n8778), .B(n8779), .Z(n8777) );
  NANDN U12967 ( .A(n8780), .B(n8781), .Z(n8778) );
  NANDN U12968 ( .A(n8781), .B(n8780), .Z(n8776) );
  AND U12969 ( .A(n8782), .B(n8783), .Z(n8737) );
  NAND U12970 ( .A(n8784), .B(n8785), .Z(n8783) );
  OR U12971 ( .A(n8786), .B(n8787), .Z(n8784) );
  NANDN U12972 ( .A(n8788), .B(n8786), .Z(n8782) );
  XNOR U12973 ( .A(n8763), .B(n8789), .Z(N29430) );
  XOR U12974 ( .A(n8765), .B(n8766), .Z(n8789) );
  XNOR U12975 ( .A(n8779), .B(n8790), .Z(n8766) );
  XOR U12976 ( .A(n8780), .B(n8781), .Z(n8790) );
  XOR U12977 ( .A(n8786), .B(n8791), .Z(n8781) );
  XOR U12978 ( .A(n8785), .B(n8788), .Z(n8791) );
  IV U12979 ( .A(n8787), .Z(n8788) );
  NAND U12980 ( .A(n8792), .B(n8793), .Z(n8787) );
  OR U12981 ( .A(n8794), .B(n8795), .Z(n8793) );
  OR U12982 ( .A(n8796), .B(n8797), .Z(n8792) );
  NAND U12983 ( .A(n8798), .B(n8799), .Z(n8785) );
  OR U12984 ( .A(n8800), .B(n8801), .Z(n8799) );
  OR U12985 ( .A(n8802), .B(n8803), .Z(n8798) );
  NOR U12986 ( .A(n8804), .B(n8805), .Z(n8786) );
  ANDN U12987 ( .B(n8806), .A(n8807), .Z(n8780) );
  XNOR U12988 ( .A(n8773), .B(n8808), .Z(n8779) );
  XNOR U12989 ( .A(n8772), .B(n8774), .Z(n8808) );
  NAND U12990 ( .A(n8809), .B(n8810), .Z(n8774) );
  OR U12991 ( .A(n8811), .B(n8812), .Z(n8810) );
  OR U12992 ( .A(n8813), .B(n8814), .Z(n8809) );
  NAND U12993 ( .A(n8815), .B(n8816), .Z(n8772) );
  OR U12994 ( .A(n8817), .B(n8818), .Z(n8816) );
  OR U12995 ( .A(n8819), .B(n8820), .Z(n8815) );
  ANDN U12996 ( .B(n8821), .A(n8822), .Z(n8773) );
  IV U12997 ( .A(n8823), .Z(n8821) );
  ANDN U12998 ( .B(n8824), .A(n8825), .Z(n8765) );
  XOR U12999 ( .A(n8751), .B(n8826), .Z(n8763) );
  XOR U13000 ( .A(n8752), .B(n8753), .Z(n8826) );
  XOR U13001 ( .A(n8758), .B(n8827), .Z(n8753) );
  XOR U13002 ( .A(n8757), .B(n8760), .Z(n8827) );
  IV U13003 ( .A(n8759), .Z(n8760) );
  NAND U13004 ( .A(n8828), .B(n8829), .Z(n8759) );
  OR U13005 ( .A(n8830), .B(n8831), .Z(n8829) );
  OR U13006 ( .A(n8832), .B(n8833), .Z(n8828) );
  NAND U13007 ( .A(n8834), .B(n8835), .Z(n8757) );
  OR U13008 ( .A(n8836), .B(n8837), .Z(n8835) );
  OR U13009 ( .A(n8838), .B(n8839), .Z(n8834) );
  NOR U13010 ( .A(n8840), .B(n8841), .Z(n8758) );
  ANDN U13011 ( .B(n8842), .A(n8843), .Z(n8752) );
  IV U13012 ( .A(n8844), .Z(n8842) );
  XNOR U13013 ( .A(n8745), .B(n8845), .Z(n8751) );
  XNOR U13014 ( .A(n8744), .B(n8746), .Z(n8845) );
  NAND U13015 ( .A(n8846), .B(n8847), .Z(n8746) );
  OR U13016 ( .A(n8848), .B(n8849), .Z(n8847) );
  OR U13017 ( .A(n8850), .B(n8851), .Z(n8846) );
  NAND U13018 ( .A(n8852), .B(n8853), .Z(n8744) );
  OR U13019 ( .A(n8854), .B(n8855), .Z(n8853) );
  OR U13020 ( .A(n8856), .B(n8857), .Z(n8852) );
  ANDN U13021 ( .B(n8858), .A(n8859), .Z(n8745) );
  IV U13022 ( .A(n8860), .Z(n8858) );
  XNOR U13023 ( .A(n8825), .B(n8824), .Z(N29429) );
  XOR U13024 ( .A(n8844), .B(n8843), .Z(n8824) );
  XNOR U13025 ( .A(n8859), .B(n8860), .Z(n8843) );
  XNOR U13026 ( .A(n8854), .B(n8855), .Z(n8860) );
  XNOR U13027 ( .A(n8856), .B(n8857), .Z(n8855) );
  XNOR U13028 ( .A(y[3004]), .B(x[3004]), .Z(n8857) );
  XNOR U13029 ( .A(y[3005]), .B(x[3005]), .Z(n8856) );
  XNOR U13030 ( .A(y[3003]), .B(x[3003]), .Z(n8854) );
  XNOR U13031 ( .A(n8848), .B(n8849), .Z(n8859) );
  XNOR U13032 ( .A(y[3000]), .B(x[3000]), .Z(n8849) );
  XNOR U13033 ( .A(n8850), .B(n8851), .Z(n8848) );
  XNOR U13034 ( .A(y[3001]), .B(x[3001]), .Z(n8851) );
  XNOR U13035 ( .A(y[3002]), .B(x[3002]), .Z(n8850) );
  XNOR U13036 ( .A(n8841), .B(n8840), .Z(n8844) );
  XNOR U13037 ( .A(n8836), .B(n8837), .Z(n8840) );
  XNOR U13038 ( .A(y[2997]), .B(x[2997]), .Z(n8837) );
  XNOR U13039 ( .A(n8838), .B(n8839), .Z(n8836) );
  XNOR U13040 ( .A(y[2998]), .B(x[2998]), .Z(n8839) );
  XNOR U13041 ( .A(y[2999]), .B(x[2999]), .Z(n8838) );
  XNOR U13042 ( .A(n8830), .B(n8831), .Z(n8841) );
  XNOR U13043 ( .A(y[2994]), .B(x[2994]), .Z(n8831) );
  XNOR U13044 ( .A(n8832), .B(n8833), .Z(n8830) );
  XNOR U13045 ( .A(y[2995]), .B(x[2995]), .Z(n8833) );
  XNOR U13046 ( .A(y[2996]), .B(x[2996]), .Z(n8832) );
  XOR U13047 ( .A(n8806), .B(n8807), .Z(n8825) );
  XNOR U13048 ( .A(n8822), .B(n8823), .Z(n8807) );
  XNOR U13049 ( .A(n8817), .B(n8818), .Z(n8823) );
  XNOR U13050 ( .A(n8819), .B(n8820), .Z(n8818) );
  XNOR U13051 ( .A(y[2992]), .B(x[2992]), .Z(n8820) );
  XNOR U13052 ( .A(y[2993]), .B(x[2993]), .Z(n8819) );
  XNOR U13053 ( .A(y[2991]), .B(x[2991]), .Z(n8817) );
  XNOR U13054 ( .A(n8811), .B(n8812), .Z(n8822) );
  XNOR U13055 ( .A(y[2988]), .B(x[2988]), .Z(n8812) );
  XNOR U13056 ( .A(n8813), .B(n8814), .Z(n8811) );
  XNOR U13057 ( .A(y[2989]), .B(x[2989]), .Z(n8814) );
  XNOR U13058 ( .A(y[2990]), .B(x[2990]), .Z(n8813) );
  XOR U13059 ( .A(n8805), .B(n8804), .Z(n8806) );
  XNOR U13060 ( .A(n8800), .B(n8801), .Z(n8804) );
  XNOR U13061 ( .A(y[2985]), .B(x[2985]), .Z(n8801) );
  XNOR U13062 ( .A(n8802), .B(n8803), .Z(n8800) );
  XNOR U13063 ( .A(y[2986]), .B(x[2986]), .Z(n8803) );
  XNOR U13064 ( .A(y[2987]), .B(x[2987]), .Z(n8802) );
  XNOR U13065 ( .A(n8794), .B(n8795), .Z(n8805) );
  XNOR U13066 ( .A(y[2982]), .B(x[2982]), .Z(n8795) );
  XNOR U13067 ( .A(n8796), .B(n8797), .Z(n8794) );
  XNOR U13068 ( .A(y[2983]), .B(x[2983]), .Z(n8797) );
  XNOR U13069 ( .A(y[2984]), .B(x[2984]), .Z(n8796) );
  NAND U13070 ( .A(n8861), .B(n8862), .Z(N29421) );
  NANDN U13071 ( .A(n8863), .B(n8864), .Z(n8862) );
  OR U13072 ( .A(n8865), .B(n8866), .Z(n8864) );
  NAND U13073 ( .A(n8865), .B(n8866), .Z(n8861) );
  XOR U13074 ( .A(n8865), .B(n8867), .Z(N29420) );
  XNOR U13075 ( .A(n8863), .B(n8866), .Z(n8867) );
  AND U13076 ( .A(n8868), .B(n8869), .Z(n8866) );
  NANDN U13077 ( .A(n8870), .B(n8871), .Z(n8869) );
  NANDN U13078 ( .A(n8872), .B(n8873), .Z(n8871) );
  NANDN U13079 ( .A(n8873), .B(n8872), .Z(n8868) );
  NAND U13080 ( .A(n8874), .B(n8875), .Z(n8863) );
  NANDN U13081 ( .A(n8876), .B(n8877), .Z(n8875) );
  OR U13082 ( .A(n8878), .B(n8879), .Z(n8877) );
  NAND U13083 ( .A(n8879), .B(n8878), .Z(n8874) );
  AND U13084 ( .A(n8880), .B(n8881), .Z(n8865) );
  NANDN U13085 ( .A(n8882), .B(n8883), .Z(n8881) );
  NANDN U13086 ( .A(n8884), .B(n8885), .Z(n8883) );
  NANDN U13087 ( .A(n8885), .B(n8884), .Z(n8880) );
  XOR U13088 ( .A(n8879), .B(n8886), .Z(N29419) );
  XOR U13089 ( .A(n8876), .B(n8878), .Z(n8886) );
  XNOR U13090 ( .A(n8872), .B(n8887), .Z(n8878) );
  XNOR U13091 ( .A(n8870), .B(n8873), .Z(n8887) );
  NAND U13092 ( .A(n8888), .B(n8889), .Z(n8873) );
  NAND U13093 ( .A(n8890), .B(n8891), .Z(n8889) );
  OR U13094 ( .A(n8892), .B(n8893), .Z(n8890) );
  NANDN U13095 ( .A(n8894), .B(n8892), .Z(n8888) );
  IV U13096 ( .A(n8893), .Z(n8894) );
  NAND U13097 ( .A(n8895), .B(n8896), .Z(n8870) );
  NAND U13098 ( .A(n8897), .B(n8898), .Z(n8896) );
  NANDN U13099 ( .A(n8899), .B(n8900), .Z(n8897) );
  NANDN U13100 ( .A(n8900), .B(n8899), .Z(n8895) );
  AND U13101 ( .A(n8901), .B(n8902), .Z(n8872) );
  NAND U13102 ( .A(n8903), .B(n8904), .Z(n8902) );
  OR U13103 ( .A(n8905), .B(n8906), .Z(n8903) );
  NANDN U13104 ( .A(n8907), .B(n8905), .Z(n8901) );
  NAND U13105 ( .A(n8908), .B(n8909), .Z(n8876) );
  NANDN U13106 ( .A(n8910), .B(n8911), .Z(n8909) );
  OR U13107 ( .A(n8912), .B(n8913), .Z(n8911) );
  NANDN U13108 ( .A(n8914), .B(n8912), .Z(n8908) );
  IV U13109 ( .A(n8913), .Z(n8914) );
  XNOR U13110 ( .A(n8884), .B(n8915), .Z(n8879) );
  XNOR U13111 ( .A(n8882), .B(n8885), .Z(n8915) );
  NAND U13112 ( .A(n8916), .B(n8917), .Z(n8885) );
  NAND U13113 ( .A(n8918), .B(n8919), .Z(n8917) );
  OR U13114 ( .A(n8920), .B(n8921), .Z(n8918) );
  NANDN U13115 ( .A(n8922), .B(n8920), .Z(n8916) );
  IV U13116 ( .A(n8921), .Z(n8922) );
  NAND U13117 ( .A(n8923), .B(n8924), .Z(n8882) );
  NAND U13118 ( .A(n8925), .B(n8926), .Z(n8924) );
  NANDN U13119 ( .A(n8927), .B(n8928), .Z(n8925) );
  NANDN U13120 ( .A(n8928), .B(n8927), .Z(n8923) );
  AND U13121 ( .A(n8929), .B(n8930), .Z(n8884) );
  NAND U13122 ( .A(n8931), .B(n8932), .Z(n8930) );
  OR U13123 ( .A(n8933), .B(n8934), .Z(n8931) );
  NANDN U13124 ( .A(n8935), .B(n8933), .Z(n8929) );
  XNOR U13125 ( .A(n8910), .B(n8936), .Z(N29418) );
  XOR U13126 ( .A(n8912), .B(n8913), .Z(n8936) );
  XNOR U13127 ( .A(n8926), .B(n8937), .Z(n8913) );
  XOR U13128 ( .A(n8927), .B(n8928), .Z(n8937) );
  XOR U13129 ( .A(n8933), .B(n8938), .Z(n8928) );
  XOR U13130 ( .A(n8932), .B(n8935), .Z(n8938) );
  IV U13131 ( .A(n8934), .Z(n8935) );
  NAND U13132 ( .A(n8939), .B(n8940), .Z(n8934) );
  OR U13133 ( .A(n8941), .B(n8942), .Z(n8940) );
  OR U13134 ( .A(n8943), .B(n8944), .Z(n8939) );
  NAND U13135 ( .A(n8945), .B(n8946), .Z(n8932) );
  OR U13136 ( .A(n8947), .B(n8948), .Z(n8946) );
  OR U13137 ( .A(n8949), .B(n8950), .Z(n8945) );
  NOR U13138 ( .A(n8951), .B(n8952), .Z(n8933) );
  ANDN U13139 ( .B(n8953), .A(n8954), .Z(n8927) );
  XNOR U13140 ( .A(n8920), .B(n8955), .Z(n8926) );
  XNOR U13141 ( .A(n8919), .B(n8921), .Z(n8955) );
  NAND U13142 ( .A(n8956), .B(n8957), .Z(n8921) );
  OR U13143 ( .A(n8958), .B(n8959), .Z(n8957) );
  OR U13144 ( .A(n8960), .B(n8961), .Z(n8956) );
  NAND U13145 ( .A(n8962), .B(n8963), .Z(n8919) );
  OR U13146 ( .A(n8964), .B(n8965), .Z(n8963) );
  OR U13147 ( .A(n8966), .B(n8967), .Z(n8962) );
  ANDN U13148 ( .B(n8968), .A(n8969), .Z(n8920) );
  IV U13149 ( .A(n8970), .Z(n8968) );
  ANDN U13150 ( .B(n8971), .A(n8972), .Z(n8912) );
  XOR U13151 ( .A(n8898), .B(n8973), .Z(n8910) );
  XOR U13152 ( .A(n8899), .B(n8900), .Z(n8973) );
  XOR U13153 ( .A(n8905), .B(n8974), .Z(n8900) );
  XOR U13154 ( .A(n8904), .B(n8907), .Z(n8974) );
  IV U13155 ( .A(n8906), .Z(n8907) );
  NAND U13156 ( .A(n8975), .B(n8976), .Z(n8906) );
  OR U13157 ( .A(n8977), .B(n8978), .Z(n8976) );
  OR U13158 ( .A(n8979), .B(n8980), .Z(n8975) );
  NAND U13159 ( .A(n8981), .B(n8982), .Z(n8904) );
  OR U13160 ( .A(n8983), .B(n8984), .Z(n8982) );
  OR U13161 ( .A(n8985), .B(n8986), .Z(n8981) );
  NOR U13162 ( .A(n8987), .B(n8988), .Z(n8905) );
  ANDN U13163 ( .B(n8989), .A(n8990), .Z(n8899) );
  IV U13164 ( .A(n8991), .Z(n8989) );
  XNOR U13165 ( .A(n8892), .B(n8992), .Z(n8898) );
  XNOR U13166 ( .A(n8891), .B(n8893), .Z(n8992) );
  NAND U13167 ( .A(n8993), .B(n8994), .Z(n8893) );
  OR U13168 ( .A(n8995), .B(n8996), .Z(n8994) );
  OR U13169 ( .A(n8997), .B(n8998), .Z(n8993) );
  NAND U13170 ( .A(n8999), .B(n9000), .Z(n8891) );
  OR U13171 ( .A(n9001), .B(n9002), .Z(n9000) );
  OR U13172 ( .A(n9003), .B(n9004), .Z(n8999) );
  ANDN U13173 ( .B(n9005), .A(n9006), .Z(n8892) );
  IV U13174 ( .A(n9007), .Z(n9005) );
  XNOR U13175 ( .A(n8972), .B(n8971), .Z(N29417) );
  XOR U13176 ( .A(n8991), .B(n8990), .Z(n8971) );
  XNOR U13177 ( .A(n9006), .B(n9007), .Z(n8990) );
  XNOR U13178 ( .A(n9001), .B(n9002), .Z(n9007) );
  XNOR U13179 ( .A(n9003), .B(n9004), .Z(n9002) );
  XNOR U13180 ( .A(y[2980]), .B(x[2980]), .Z(n9004) );
  XNOR U13181 ( .A(y[2981]), .B(x[2981]), .Z(n9003) );
  XNOR U13182 ( .A(y[2979]), .B(x[2979]), .Z(n9001) );
  XNOR U13183 ( .A(n8995), .B(n8996), .Z(n9006) );
  XNOR U13184 ( .A(y[2976]), .B(x[2976]), .Z(n8996) );
  XNOR U13185 ( .A(n8997), .B(n8998), .Z(n8995) );
  XNOR U13186 ( .A(y[2977]), .B(x[2977]), .Z(n8998) );
  XNOR U13187 ( .A(y[2978]), .B(x[2978]), .Z(n8997) );
  XNOR U13188 ( .A(n8988), .B(n8987), .Z(n8991) );
  XNOR U13189 ( .A(n8983), .B(n8984), .Z(n8987) );
  XNOR U13190 ( .A(y[2973]), .B(x[2973]), .Z(n8984) );
  XNOR U13191 ( .A(n8985), .B(n8986), .Z(n8983) );
  XNOR U13192 ( .A(y[2974]), .B(x[2974]), .Z(n8986) );
  XNOR U13193 ( .A(y[2975]), .B(x[2975]), .Z(n8985) );
  XNOR U13194 ( .A(n8977), .B(n8978), .Z(n8988) );
  XNOR U13195 ( .A(y[2970]), .B(x[2970]), .Z(n8978) );
  XNOR U13196 ( .A(n8979), .B(n8980), .Z(n8977) );
  XNOR U13197 ( .A(y[2971]), .B(x[2971]), .Z(n8980) );
  XNOR U13198 ( .A(y[2972]), .B(x[2972]), .Z(n8979) );
  XOR U13199 ( .A(n8953), .B(n8954), .Z(n8972) );
  XNOR U13200 ( .A(n8969), .B(n8970), .Z(n8954) );
  XNOR U13201 ( .A(n8964), .B(n8965), .Z(n8970) );
  XNOR U13202 ( .A(n8966), .B(n8967), .Z(n8965) );
  XNOR U13203 ( .A(y[2968]), .B(x[2968]), .Z(n8967) );
  XNOR U13204 ( .A(y[2969]), .B(x[2969]), .Z(n8966) );
  XNOR U13205 ( .A(y[2967]), .B(x[2967]), .Z(n8964) );
  XNOR U13206 ( .A(n8958), .B(n8959), .Z(n8969) );
  XNOR U13207 ( .A(y[2964]), .B(x[2964]), .Z(n8959) );
  XNOR U13208 ( .A(n8960), .B(n8961), .Z(n8958) );
  XNOR U13209 ( .A(y[2965]), .B(x[2965]), .Z(n8961) );
  XNOR U13210 ( .A(y[2966]), .B(x[2966]), .Z(n8960) );
  XOR U13211 ( .A(n8952), .B(n8951), .Z(n8953) );
  XNOR U13212 ( .A(n8947), .B(n8948), .Z(n8951) );
  XNOR U13213 ( .A(y[2961]), .B(x[2961]), .Z(n8948) );
  XNOR U13214 ( .A(n8949), .B(n8950), .Z(n8947) );
  XNOR U13215 ( .A(y[2962]), .B(x[2962]), .Z(n8950) );
  XNOR U13216 ( .A(y[2963]), .B(x[2963]), .Z(n8949) );
  XNOR U13217 ( .A(n8941), .B(n8942), .Z(n8952) );
  XNOR U13218 ( .A(y[2958]), .B(x[2958]), .Z(n8942) );
  XNOR U13219 ( .A(n8943), .B(n8944), .Z(n8941) );
  XNOR U13220 ( .A(y[2959]), .B(x[2959]), .Z(n8944) );
  XNOR U13221 ( .A(y[2960]), .B(x[2960]), .Z(n8943) );
  NAND U13222 ( .A(n9008), .B(n9009), .Z(N29409) );
  NANDN U13223 ( .A(n9010), .B(n9011), .Z(n9009) );
  OR U13224 ( .A(n9012), .B(n9013), .Z(n9011) );
  NAND U13225 ( .A(n9012), .B(n9013), .Z(n9008) );
  XOR U13226 ( .A(n9012), .B(n9014), .Z(N29408) );
  XNOR U13227 ( .A(n9010), .B(n9013), .Z(n9014) );
  AND U13228 ( .A(n9015), .B(n9016), .Z(n9013) );
  NANDN U13229 ( .A(n9017), .B(n9018), .Z(n9016) );
  NANDN U13230 ( .A(n9019), .B(n9020), .Z(n9018) );
  NANDN U13231 ( .A(n9020), .B(n9019), .Z(n9015) );
  NAND U13232 ( .A(n9021), .B(n9022), .Z(n9010) );
  NANDN U13233 ( .A(n9023), .B(n9024), .Z(n9022) );
  OR U13234 ( .A(n9025), .B(n9026), .Z(n9024) );
  NAND U13235 ( .A(n9026), .B(n9025), .Z(n9021) );
  AND U13236 ( .A(n9027), .B(n9028), .Z(n9012) );
  NANDN U13237 ( .A(n9029), .B(n9030), .Z(n9028) );
  NANDN U13238 ( .A(n9031), .B(n9032), .Z(n9030) );
  NANDN U13239 ( .A(n9032), .B(n9031), .Z(n9027) );
  XOR U13240 ( .A(n9026), .B(n9033), .Z(N29407) );
  XOR U13241 ( .A(n9023), .B(n9025), .Z(n9033) );
  XNOR U13242 ( .A(n9019), .B(n9034), .Z(n9025) );
  XNOR U13243 ( .A(n9017), .B(n9020), .Z(n9034) );
  NAND U13244 ( .A(n9035), .B(n9036), .Z(n9020) );
  NAND U13245 ( .A(n9037), .B(n9038), .Z(n9036) );
  OR U13246 ( .A(n9039), .B(n9040), .Z(n9037) );
  NANDN U13247 ( .A(n9041), .B(n9039), .Z(n9035) );
  IV U13248 ( .A(n9040), .Z(n9041) );
  NAND U13249 ( .A(n9042), .B(n9043), .Z(n9017) );
  NAND U13250 ( .A(n9044), .B(n9045), .Z(n9043) );
  NANDN U13251 ( .A(n9046), .B(n9047), .Z(n9044) );
  NANDN U13252 ( .A(n9047), .B(n9046), .Z(n9042) );
  AND U13253 ( .A(n9048), .B(n9049), .Z(n9019) );
  NAND U13254 ( .A(n9050), .B(n9051), .Z(n9049) );
  OR U13255 ( .A(n9052), .B(n9053), .Z(n9050) );
  NANDN U13256 ( .A(n9054), .B(n9052), .Z(n9048) );
  NAND U13257 ( .A(n9055), .B(n9056), .Z(n9023) );
  NANDN U13258 ( .A(n9057), .B(n9058), .Z(n9056) );
  OR U13259 ( .A(n9059), .B(n9060), .Z(n9058) );
  NANDN U13260 ( .A(n9061), .B(n9059), .Z(n9055) );
  IV U13261 ( .A(n9060), .Z(n9061) );
  XNOR U13262 ( .A(n9031), .B(n9062), .Z(n9026) );
  XNOR U13263 ( .A(n9029), .B(n9032), .Z(n9062) );
  NAND U13264 ( .A(n9063), .B(n9064), .Z(n9032) );
  NAND U13265 ( .A(n9065), .B(n9066), .Z(n9064) );
  OR U13266 ( .A(n9067), .B(n9068), .Z(n9065) );
  NANDN U13267 ( .A(n9069), .B(n9067), .Z(n9063) );
  IV U13268 ( .A(n9068), .Z(n9069) );
  NAND U13269 ( .A(n9070), .B(n9071), .Z(n9029) );
  NAND U13270 ( .A(n9072), .B(n9073), .Z(n9071) );
  NANDN U13271 ( .A(n9074), .B(n9075), .Z(n9072) );
  NANDN U13272 ( .A(n9075), .B(n9074), .Z(n9070) );
  AND U13273 ( .A(n9076), .B(n9077), .Z(n9031) );
  NAND U13274 ( .A(n9078), .B(n9079), .Z(n9077) );
  OR U13275 ( .A(n9080), .B(n9081), .Z(n9078) );
  NANDN U13276 ( .A(n9082), .B(n9080), .Z(n9076) );
  XNOR U13277 ( .A(n9057), .B(n9083), .Z(N29406) );
  XOR U13278 ( .A(n9059), .B(n9060), .Z(n9083) );
  XNOR U13279 ( .A(n9073), .B(n9084), .Z(n9060) );
  XOR U13280 ( .A(n9074), .B(n9075), .Z(n9084) );
  XOR U13281 ( .A(n9080), .B(n9085), .Z(n9075) );
  XOR U13282 ( .A(n9079), .B(n9082), .Z(n9085) );
  IV U13283 ( .A(n9081), .Z(n9082) );
  NAND U13284 ( .A(n9086), .B(n9087), .Z(n9081) );
  OR U13285 ( .A(n9088), .B(n9089), .Z(n9087) );
  OR U13286 ( .A(n9090), .B(n9091), .Z(n9086) );
  NAND U13287 ( .A(n9092), .B(n9093), .Z(n9079) );
  OR U13288 ( .A(n9094), .B(n9095), .Z(n9093) );
  OR U13289 ( .A(n9096), .B(n9097), .Z(n9092) );
  NOR U13290 ( .A(n9098), .B(n9099), .Z(n9080) );
  ANDN U13291 ( .B(n9100), .A(n9101), .Z(n9074) );
  XNOR U13292 ( .A(n9067), .B(n9102), .Z(n9073) );
  XNOR U13293 ( .A(n9066), .B(n9068), .Z(n9102) );
  NAND U13294 ( .A(n9103), .B(n9104), .Z(n9068) );
  OR U13295 ( .A(n9105), .B(n9106), .Z(n9104) );
  OR U13296 ( .A(n9107), .B(n9108), .Z(n9103) );
  NAND U13297 ( .A(n9109), .B(n9110), .Z(n9066) );
  OR U13298 ( .A(n9111), .B(n9112), .Z(n9110) );
  OR U13299 ( .A(n9113), .B(n9114), .Z(n9109) );
  ANDN U13300 ( .B(n9115), .A(n9116), .Z(n9067) );
  IV U13301 ( .A(n9117), .Z(n9115) );
  ANDN U13302 ( .B(n9118), .A(n9119), .Z(n9059) );
  XOR U13303 ( .A(n9045), .B(n9120), .Z(n9057) );
  XOR U13304 ( .A(n9046), .B(n9047), .Z(n9120) );
  XOR U13305 ( .A(n9052), .B(n9121), .Z(n9047) );
  XOR U13306 ( .A(n9051), .B(n9054), .Z(n9121) );
  IV U13307 ( .A(n9053), .Z(n9054) );
  NAND U13308 ( .A(n9122), .B(n9123), .Z(n9053) );
  OR U13309 ( .A(n9124), .B(n9125), .Z(n9123) );
  OR U13310 ( .A(n9126), .B(n9127), .Z(n9122) );
  NAND U13311 ( .A(n9128), .B(n9129), .Z(n9051) );
  OR U13312 ( .A(n9130), .B(n9131), .Z(n9129) );
  OR U13313 ( .A(n9132), .B(n9133), .Z(n9128) );
  NOR U13314 ( .A(n9134), .B(n9135), .Z(n9052) );
  ANDN U13315 ( .B(n9136), .A(n9137), .Z(n9046) );
  IV U13316 ( .A(n9138), .Z(n9136) );
  XNOR U13317 ( .A(n9039), .B(n9139), .Z(n9045) );
  XNOR U13318 ( .A(n9038), .B(n9040), .Z(n9139) );
  NAND U13319 ( .A(n9140), .B(n9141), .Z(n9040) );
  OR U13320 ( .A(n9142), .B(n9143), .Z(n9141) );
  OR U13321 ( .A(n9144), .B(n9145), .Z(n9140) );
  NAND U13322 ( .A(n9146), .B(n9147), .Z(n9038) );
  OR U13323 ( .A(n9148), .B(n9149), .Z(n9147) );
  OR U13324 ( .A(n9150), .B(n9151), .Z(n9146) );
  ANDN U13325 ( .B(n9152), .A(n9153), .Z(n9039) );
  IV U13326 ( .A(n9154), .Z(n9152) );
  XNOR U13327 ( .A(n9119), .B(n9118), .Z(N29405) );
  XOR U13328 ( .A(n9138), .B(n9137), .Z(n9118) );
  XNOR U13329 ( .A(n9153), .B(n9154), .Z(n9137) );
  XNOR U13330 ( .A(n9148), .B(n9149), .Z(n9154) );
  XNOR U13331 ( .A(n9150), .B(n9151), .Z(n9149) );
  XNOR U13332 ( .A(y[2956]), .B(x[2956]), .Z(n9151) );
  XNOR U13333 ( .A(y[2957]), .B(x[2957]), .Z(n9150) );
  XNOR U13334 ( .A(y[2955]), .B(x[2955]), .Z(n9148) );
  XNOR U13335 ( .A(n9142), .B(n9143), .Z(n9153) );
  XNOR U13336 ( .A(y[2952]), .B(x[2952]), .Z(n9143) );
  XNOR U13337 ( .A(n9144), .B(n9145), .Z(n9142) );
  XNOR U13338 ( .A(y[2953]), .B(x[2953]), .Z(n9145) );
  XNOR U13339 ( .A(y[2954]), .B(x[2954]), .Z(n9144) );
  XNOR U13340 ( .A(n9135), .B(n9134), .Z(n9138) );
  XNOR U13341 ( .A(n9130), .B(n9131), .Z(n9134) );
  XNOR U13342 ( .A(y[2949]), .B(x[2949]), .Z(n9131) );
  XNOR U13343 ( .A(n9132), .B(n9133), .Z(n9130) );
  XNOR U13344 ( .A(y[2950]), .B(x[2950]), .Z(n9133) );
  XNOR U13345 ( .A(y[2951]), .B(x[2951]), .Z(n9132) );
  XNOR U13346 ( .A(n9124), .B(n9125), .Z(n9135) );
  XNOR U13347 ( .A(y[2946]), .B(x[2946]), .Z(n9125) );
  XNOR U13348 ( .A(n9126), .B(n9127), .Z(n9124) );
  XNOR U13349 ( .A(y[2947]), .B(x[2947]), .Z(n9127) );
  XNOR U13350 ( .A(y[2948]), .B(x[2948]), .Z(n9126) );
  XOR U13351 ( .A(n9100), .B(n9101), .Z(n9119) );
  XNOR U13352 ( .A(n9116), .B(n9117), .Z(n9101) );
  XNOR U13353 ( .A(n9111), .B(n9112), .Z(n9117) );
  XNOR U13354 ( .A(n9113), .B(n9114), .Z(n9112) );
  XNOR U13355 ( .A(y[2944]), .B(x[2944]), .Z(n9114) );
  XNOR U13356 ( .A(y[2945]), .B(x[2945]), .Z(n9113) );
  XNOR U13357 ( .A(y[2943]), .B(x[2943]), .Z(n9111) );
  XNOR U13358 ( .A(n9105), .B(n9106), .Z(n9116) );
  XNOR U13359 ( .A(y[2940]), .B(x[2940]), .Z(n9106) );
  XNOR U13360 ( .A(n9107), .B(n9108), .Z(n9105) );
  XNOR U13361 ( .A(y[2941]), .B(x[2941]), .Z(n9108) );
  XNOR U13362 ( .A(y[2942]), .B(x[2942]), .Z(n9107) );
  XOR U13363 ( .A(n9099), .B(n9098), .Z(n9100) );
  XNOR U13364 ( .A(n9094), .B(n9095), .Z(n9098) );
  XNOR U13365 ( .A(y[2937]), .B(x[2937]), .Z(n9095) );
  XNOR U13366 ( .A(n9096), .B(n9097), .Z(n9094) );
  XNOR U13367 ( .A(y[2938]), .B(x[2938]), .Z(n9097) );
  XNOR U13368 ( .A(y[2939]), .B(x[2939]), .Z(n9096) );
  XNOR U13369 ( .A(n9088), .B(n9089), .Z(n9099) );
  XNOR U13370 ( .A(y[2934]), .B(x[2934]), .Z(n9089) );
  XNOR U13371 ( .A(n9090), .B(n9091), .Z(n9088) );
  XNOR U13372 ( .A(y[2935]), .B(x[2935]), .Z(n9091) );
  XNOR U13373 ( .A(y[2936]), .B(x[2936]), .Z(n9090) );
  NAND U13374 ( .A(n9155), .B(n9156), .Z(N29397) );
  NANDN U13375 ( .A(n9157), .B(n9158), .Z(n9156) );
  OR U13376 ( .A(n9159), .B(n9160), .Z(n9158) );
  NAND U13377 ( .A(n9159), .B(n9160), .Z(n9155) );
  XOR U13378 ( .A(n9159), .B(n9161), .Z(N29396) );
  XNOR U13379 ( .A(n9157), .B(n9160), .Z(n9161) );
  AND U13380 ( .A(n9162), .B(n9163), .Z(n9160) );
  NANDN U13381 ( .A(n9164), .B(n9165), .Z(n9163) );
  NANDN U13382 ( .A(n9166), .B(n9167), .Z(n9165) );
  NANDN U13383 ( .A(n9167), .B(n9166), .Z(n9162) );
  NAND U13384 ( .A(n9168), .B(n9169), .Z(n9157) );
  NANDN U13385 ( .A(n9170), .B(n9171), .Z(n9169) );
  OR U13386 ( .A(n9172), .B(n9173), .Z(n9171) );
  NAND U13387 ( .A(n9173), .B(n9172), .Z(n9168) );
  AND U13388 ( .A(n9174), .B(n9175), .Z(n9159) );
  NANDN U13389 ( .A(n9176), .B(n9177), .Z(n9175) );
  NANDN U13390 ( .A(n9178), .B(n9179), .Z(n9177) );
  NANDN U13391 ( .A(n9179), .B(n9178), .Z(n9174) );
  XOR U13392 ( .A(n9173), .B(n9180), .Z(N29395) );
  XOR U13393 ( .A(n9170), .B(n9172), .Z(n9180) );
  XNOR U13394 ( .A(n9166), .B(n9181), .Z(n9172) );
  XNOR U13395 ( .A(n9164), .B(n9167), .Z(n9181) );
  NAND U13396 ( .A(n9182), .B(n9183), .Z(n9167) );
  NAND U13397 ( .A(n9184), .B(n9185), .Z(n9183) );
  OR U13398 ( .A(n9186), .B(n9187), .Z(n9184) );
  NANDN U13399 ( .A(n9188), .B(n9186), .Z(n9182) );
  IV U13400 ( .A(n9187), .Z(n9188) );
  NAND U13401 ( .A(n9189), .B(n9190), .Z(n9164) );
  NAND U13402 ( .A(n9191), .B(n9192), .Z(n9190) );
  NANDN U13403 ( .A(n9193), .B(n9194), .Z(n9191) );
  NANDN U13404 ( .A(n9194), .B(n9193), .Z(n9189) );
  AND U13405 ( .A(n9195), .B(n9196), .Z(n9166) );
  NAND U13406 ( .A(n9197), .B(n9198), .Z(n9196) );
  OR U13407 ( .A(n9199), .B(n9200), .Z(n9197) );
  NANDN U13408 ( .A(n9201), .B(n9199), .Z(n9195) );
  NAND U13409 ( .A(n9202), .B(n9203), .Z(n9170) );
  NANDN U13410 ( .A(n9204), .B(n9205), .Z(n9203) );
  OR U13411 ( .A(n9206), .B(n9207), .Z(n9205) );
  NANDN U13412 ( .A(n9208), .B(n9206), .Z(n9202) );
  IV U13413 ( .A(n9207), .Z(n9208) );
  XNOR U13414 ( .A(n9178), .B(n9209), .Z(n9173) );
  XNOR U13415 ( .A(n9176), .B(n9179), .Z(n9209) );
  NAND U13416 ( .A(n9210), .B(n9211), .Z(n9179) );
  NAND U13417 ( .A(n9212), .B(n9213), .Z(n9211) );
  OR U13418 ( .A(n9214), .B(n9215), .Z(n9212) );
  NANDN U13419 ( .A(n9216), .B(n9214), .Z(n9210) );
  IV U13420 ( .A(n9215), .Z(n9216) );
  NAND U13421 ( .A(n9217), .B(n9218), .Z(n9176) );
  NAND U13422 ( .A(n9219), .B(n9220), .Z(n9218) );
  NANDN U13423 ( .A(n9221), .B(n9222), .Z(n9219) );
  NANDN U13424 ( .A(n9222), .B(n9221), .Z(n9217) );
  AND U13425 ( .A(n9223), .B(n9224), .Z(n9178) );
  NAND U13426 ( .A(n9225), .B(n9226), .Z(n9224) );
  OR U13427 ( .A(n9227), .B(n9228), .Z(n9225) );
  NANDN U13428 ( .A(n9229), .B(n9227), .Z(n9223) );
  XNOR U13429 ( .A(n9204), .B(n9230), .Z(N29394) );
  XOR U13430 ( .A(n9206), .B(n9207), .Z(n9230) );
  XNOR U13431 ( .A(n9220), .B(n9231), .Z(n9207) );
  XOR U13432 ( .A(n9221), .B(n9222), .Z(n9231) );
  XOR U13433 ( .A(n9227), .B(n9232), .Z(n9222) );
  XOR U13434 ( .A(n9226), .B(n9229), .Z(n9232) );
  IV U13435 ( .A(n9228), .Z(n9229) );
  NAND U13436 ( .A(n9233), .B(n9234), .Z(n9228) );
  OR U13437 ( .A(n9235), .B(n9236), .Z(n9234) );
  OR U13438 ( .A(n9237), .B(n9238), .Z(n9233) );
  NAND U13439 ( .A(n9239), .B(n9240), .Z(n9226) );
  OR U13440 ( .A(n9241), .B(n9242), .Z(n9240) );
  OR U13441 ( .A(n9243), .B(n9244), .Z(n9239) );
  NOR U13442 ( .A(n9245), .B(n9246), .Z(n9227) );
  ANDN U13443 ( .B(n9247), .A(n9248), .Z(n9221) );
  XNOR U13444 ( .A(n9214), .B(n9249), .Z(n9220) );
  XNOR U13445 ( .A(n9213), .B(n9215), .Z(n9249) );
  NAND U13446 ( .A(n9250), .B(n9251), .Z(n9215) );
  OR U13447 ( .A(n9252), .B(n9253), .Z(n9251) );
  OR U13448 ( .A(n9254), .B(n9255), .Z(n9250) );
  NAND U13449 ( .A(n9256), .B(n9257), .Z(n9213) );
  OR U13450 ( .A(n9258), .B(n9259), .Z(n9257) );
  OR U13451 ( .A(n9260), .B(n9261), .Z(n9256) );
  ANDN U13452 ( .B(n9262), .A(n9263), .Z(n9214) );
  IV U13453 ( .A(n9264), .Z(n9262) );
  ANDN U13454 ( .B(n9265), .A(n9266), .Z(n9206) );
  XOR U13455 ( .A(n9192), .B(n9267), .Z(n9204) );
  XOR U13456 ( .A(n9193), .B(n9194), .Z(n9267) );
  XOR U13457 ( .A(n9199), .B(n9268), .Z(n9194) );
  XOR U13458 ( .A(n9198), .B(n9201), .Z(n9268) );
  IV U13459 ( .A(n9200), .Z(n9201) );
  NAND U13460 ( .A(n9269), .B(n9270), .Z(n9200) );
  OR U13461 ( .A(n9271), .B(n9272), .Z(n9270) );
  OR U13462 ( .A(n9273), .B(n9274), .Z(n9269) );
  NAND U13463 ( .A(n9275), .B(n9276), .Z(n9198) );
  OR U13464 ( .A(n9277), .B(n9278), .Z(n9276) );
  OR U13465 ( .A(n9279), .B(n9280), .Z(n9275) );
  NOR U13466 ( .A(n9281), .B(n9282), .Z(n9199) );
  ANDN U13467 ( .B(n9283), .A(n9284), .Z(n9193) );
  IV U13468 ( .A(n9285), .Z(n9283) );
  XNOR U13469 ( .A(n9186), .B(n9286), .Z(n9192) );
  XNOR U13470 ( .A(n9185), .B(n9187), .Z(n9286) );
  NAND U13471 ( .A(n9287), .B(n9288), .Z(n9187) );
  OR U13472 ( .A(n9289), .B(n9290), .Z(n9288) );
  OR U13473 ( .A(n9291), .B(n9292), .Z(n9287) );
  NAND U13474 ( .A(n9293), .B(n9294), .Z(n9185) );
  OR U13475 ( .A(n9295), .B(n9296), .Z(n9294) );
  OR U13476 ( .A(n9297), .B(n9298), .Z(n9293) );
  ANDN U13477 ( .B(n9299), .A(n9300), .Z(n9186) );
  IV U13478 ( .A(n9301), .Z(n9299) );
  XNOR U13479 ( .A(n9266), .B(n9265), .Z(N29393) );
  XOR U13480 ( .A(n9285), .B(n9284), .Z(n9265) );
  XNOR U13481 ( .A(n9300), .B(n9301), .Z(n9284) );
  XNOR U13482 ( .A(n9295), .B(n9296), .Z(n9301) );
  XNOR U13483 ( .A(n9297), .B(n9298), .Z(n9296) );
  XNOR U13484 ( .A(y[2932]), .B(x[2932]), .Z(n9298) );
  XNOR U13485 ( .A(y[2933]), .B(x[2933]), .Z(n9297) );
  XNOR U13486 ( .A(y[2931]), .B(x[2931]), .Z(n9295) );
  XNOR U13487 ( .A(n9289), .B(n9290), .Z(n9300) );
  XNOR U13488 ( .A(y[2928]), .B(x[2928]), .Z(n9290) );
  XNOR U13489 ( .A(n9291), .B(n9292), .Z(n9289) );
  XNOR U13490 ( .A(y[2929]), .B(x[2929]), .Z(n9292) );
  XNOR U13491 ( .A(y[2930]), .B(x[2930]), .Z(n9291) );
  XNOR U13492 ( .A(n9282), .B(n9281), .Z(n9285) );
  XNOR U13493 ( .A(n9277), .B(n9278), .Z(n9281) );
  XNOR U13494 ( .A(y[2925]), .B(x[2925]), .Z(n9278) );
  XNOR U13495 ( .A(n9279), .B(n9280), .Z(n9277) );
  XNOR U13496 ( .A(y[2926]), .B(x[2926]), .Z(n9280) );
  XNOR U13497 ( .A(y[2927]), .B(x[2927]), .Z(n9279) );
  XNOR U13498 ( .A(n9271), .B(n9272), .Z(n9282) );
  XNOR U13499 ( .A(y[2922]), .B(x[2922]), .Z(n9272) );
  XNOR U13500 ( .A(n9273), .B(n9274), .Z(n9271) );
  XNOR U13501 ( .A(y[2923]), .B(x[2923]), .Z(n9274) );
  XNOR U13502 ( .A(y[2924]), .B(x[2924]), .Z(n9273) );
  XOR U13503 ( .A(n9247), .B(n9248), .Z(n9266) );
  XNOR U13504 ( .A(n9263), .B(n9264), .Z(n9248) );
  XNOR U13505 ( .A(n9258), .B(n9259), .Z(n9264) );
  XNOR U13506 ( .A(n9260), .B(n9261), .Z(n9259) );
  XNOR U13507 ( .A(y[2920]), .B(x[2920]), .Z(n9261) );
  XNOR U13508 ( .A(y[2921]), .B(x[2921]), .Z(n9260) );
  XNOR U13509 ( .A(y[2919]), .B(x[2919]), .Z(n9258) );
  XNOR U13510 ( .A(n9252), .B(n9253), .Z(n9263) );
  XNOR U13511 ( .A(y[2916]), .B(x[2916]), .Z(n9253) );
  XNOR U13512 ( .A(n9254), .B(n9255), .Z(n9252) );
  XNOR U13513 ( .A(y[2917]), .B(x[2917]), .Z(n9255) );
  XNOR U13514 ( .A(y[2918]), .B(x[2918]), .Z(n9254) );
  XOR U13515 ( .A(n9246), .B(n9245), .Z(n9247) );
  XNOR U13516 ( .A(n9241), .B(n9242), .Z(n9245) );
  XNOR U13517 ( .A(y[2913]), .B(x[2913]), .Z(n9242) );
  XNOR U13518 ( .A(n9243), .B(n9244), .Z(n9241) );
  XNOR U13519 ( .A(y[2914]), .B(x[2914]), .Z(n9244) );
  XNOR U13520 ( .A(y[2915]), .B(x[2915]), .Z(n9243) );
  XNOR U13521 ( .A(n9235), .B(n9236), .Z(n9246) );
  XNOR U13522 ( .A(y[2910]), .B(x[2910]), .Z(n9236) );
  XNOR U13523 ( .A(n9237), .B(n9238), .Z(n9235) );
  XNOR U13524 ( .A(y[2911]), .B(x[2911]), .Z(n9238) );
  XNOR U13525 ( .A(y[2912]), .B(x[2912]), .Z(n9237) );
  NAND U13526 ( .A(n9302), .B(n9303), .Z(N29385) );
  NANDN U13527 ( .A(n9304), .B(n9305), .Z(n9303) );
  OR U13528 ( .A(n9306), .B(n9307), .Z(n9305) );
  NAND U13529 ( .A(n9306), .B(n9307), .Z(n9302) );
  XOR U13530 ( .A(n9306), .B(n9308), .Z(N29384) );
  XNOR U13531 ( .A(n9304), .B(n9307), .Z(n9308) );
  AND U13532 ( .A(n9309), .B(n9310), .Z(n9307) );
  NANDN U13533 ( .A(n9311), .B(n9312), .Z(n9310) );
  NANDN U13534 ( .A(n9313), .B(n9314), .Z(n9312) );
  NANDN U13535 ( .A(n9314), .B(n9313), .Z(n9309) );
  NAND U13536 ( .A(n9315), .B(n9316), .Z(n9304) );
  NANDN U13537 ( .A(n9317), .B(n9318), .Z(n9316) );
  OR U13538 ( .A(n9319), .B(n9320), .Z(n9318) );
  NAND U13539 ( .A(n9320), .B(n9319), .Z(n9315) );
  AND U13540 ( .A(n9321), .B(n9322), .Z(n9306) );
  NANDN U13541 ( .A(n9323), .B(n9324), .Z(n9322) );
  NANDN U13542 ( .A(n9325), .B(n9326), .Z(n9324) );
  NANDN U13543 ( .A(n9326), .B(n9325), .Z(n9321) );
  XOR U13544 ( .A(n9320), .B(n9327), .Z(N29383) );
  XOR U13545 ( .A(n9317), .B(n9319), .Z(n9327) );
  XNOR U13546 ( .A(n9313), .B(n9328), .Z(n9319) );
  XNOR U13547 ( .A(n9311), .B(n9314), .Z(n9328) );
  NAND U13548 ( .A(n9329), .B(n9330), .Z(n9314) );
  NAND U13549 ( .A(n9331), .B(n9332), .Z(n9330) );
  OR U13550 ( .A(n9333), .B(n9334), .Z(n9331) );
  NANDN U13551 ( .A(n9335), .B(n9333), .Z(n9329) );
  IV U13552 ( .A(n9334), .Z(n9335) );
  NAND U13553 ( .A(n9336), .B(n9337), .Z(n9311) );
  NAND U13554 ( .A(n9338), .B(n9339), .Z(n9337) );
  NANDN U13555 ( .A(n9340), .B(n9341), .Z(n9338) );
  NANDN U13556 ( .A(n9341), .B(n9340), .Z(n9336) );
  AND U13557 ( .A(n9342), .B(n9343), .Z(n9313) );
  NAND U13558 ( .A(n9344), .B(n9345), .Z(n9343) );
  OR U13559 ( .A(n9346), .B(n9347), .Z(n9344) );
  NANDN U13560 ( .A(n9348), .B(n9346), .Z(n9342) );
  NAND U13561 ( .A(n9349), .B(n9350), .Z(n9317) );
  NANDN U13562 ( .A(n9351), .B(n9352), .Z(n9350) );
  OR U13563 ( .A(n9353), .B(n9354), .Z(n9352) );
  NANDN U13564 ( .A(n9355), .B(n9353), .Z(n9349) );
  IV U13565 ( .A(n9354), .Z(n9355) );
  XNOR U13566 ( .A(n9325), .B(n9356), .Z(n9320) );
  XNOR U13567 ( .A(n9323), .B(n9326), .Z(n9356) );
  NAND U13568 ( .A(n9357), .B(n9358), .Z(n9326) );
  NAND U13569 ( .A(n9359), .B(n9360), .Z(n9358) );
  OR U13570 ( .A(n9361), .B(n9362), .Z(n9359) );
  NANDN U13571 ( .A(n9363), .B(n9361), .Z(n9357) );
  IV U13572 ( .A(n9362), .Z(n9363) );
  NAND U13573 ( .A(n9364), .B(n9365), .Z(n9323) );
  NAND U13574 ( .A(n9366), .B(n9367), .Z(n9365) );
  NANDN U13575 ( .A(n9368), .B(n9369), .Z(n9366) );
  NANDN U13576 ( .A(n9369), .B(n9368), .Z(n9364) );
  AND U13577 ( .A(n9370), .B(n9371), .Z(n9325) );
  NAND U13578 ( .A(n9372), .B(n9373), .Z(n9371) );
  OR U13579 ( .A(n9374), .B(n9375), .Z(n9372) );
  NANDN U13580 ( .A(n9376), .B(n9374), .Z(n9370) );
  XNOR U13581 ( .A(n9351), .B(n9377), .Z(N29382) );
  XOR U13582 ( .A(n9353), .B(n9354), .Z(n9377) );
  XNOR U13583 ( .A(n9367), .B(n9378), .Z(n9354) );
  XOR U13584 ( .A(n9368), .B(n9369), .Z(n9378) );
  XOR U13585 ( .A(n9374), .B(n9379), .Z(n9369) );
  XOR U13586 ( .A(n9373), .B(n9376), .Z(n9379) );
  IV U13587 ( .A(n9375), .Z(n9376) );
  NAND U13588 ( .A(n9380), .B(n9381), .Z(n9375) );
  OR U13589 ( .A(n9382), .B(n9383), .Z(n9381) );
  OR U13590 ( .A(n9384), .B(n9385), .Z(n9380) );
  NAND U13591 ( .A(n9386), .B(n9387), .Z(n9373) );
  OR U13592 ( .A(n9388), .B(n9389), .Z(n9387) );
  OR U13593 ( .A(n9390), .B(n9391), .Z(n9386) );
  NOR U13594 ( .A(n9392), .B(n9393), .Z(n9374) );
  ANDN U13595 ( .B(n9394), .A(n9395), .Z(n9368) );
  XNOR U13596 ( .A(n9361), .B(n9396), .Z(n9367) );
  XNOR U13597 ( .A(n9360), .B(n9362), .Z(n9396) );
  NAND U13598 ( .A(n9397), .B(n9398), .Z(n9362) );
  OR U13599 ( .A(n9399), .B(n9400), .Z(n9398) );
  OR U13600 ( .A(n9401), .B(n9402), .Z(n9397) );
  NAND U13601 ( .A(n9403), .B(n9404), .Z(n9360) );
  OR U13602 ( .A(n9405), .B(n9406), .Z(n9404) );
  OR U13603 ( .A(n9407), .B(n9408), .Z(n9403) );
  ANDN U13604 ( .B(n9409), .A(n9410), .Z(n9361) );
  IV U13605 ( .A(n9411), .Z(n9409) );
  ANDN U13606 ( .B(n9412), .A(n9413), .Z(n9353) );
  XOR U13607 ( .A(n9339), .B(n9414), .Z(n9351) );
  XOR U13608 ( .A(n9340), .B(n9341), .Z(n9414) );
  XOR U13609 ( .A(n9346), .B(n9415), .Z(n9341) );
  XOR U13610 ( .A(n9345), .B(n9348), .Z(n9415) );
  IV U13611 ( .A(n9347), .Z(n9348) );
  NAND U13612 ( .A(n9416), .B(n9417), .Z(n9347) );
  OR U13613 ( .A(n9418), .B(n9419), .Z(n9417) );
  OR U13614 ( .A(n9420), .B(n9421), .Z(n9416) );
  NAND U13615 ( .A(n9422), .B(n9423), .Z(n9345) );
  OR U13616 ( .A(n9424), .B(n9425), .Z(n9423) );
  OR U13617 ( .A(n9426), .B(n9427), .Z(n9422) );
  NOR U13618 ( .A(n9428), .B(n9429), .Z(n9346) );
  ANDN U13619 ( .B(n9430), .A(n9431), .Z(n9340) );
  IV U13620 ( .A(n9432), .Z(n9430) );
  XNOR U13621 ( .A(n9333), .B(n9433), .Z(n9339) );
  XNOR U13622 ( .A(n9332), .B(n9334), .Z(n9433) );
  NAND U13623 ( .A(n9434), .B(n9435), .Z(n9334) );
  OR U13624 ( .A(n9436), .B(n9437), .Z(n9435) );
  OR U13625 ( .A(n9438), .B(n9439), .Z(n9434) );
  NAND U13626 ( .A(n9440), .B(n9441), .Z(n9332) );
  OR U13627 ( .A(n9442), .B(n9443), .Z(n9441) );
  OR U13628 ( .A(n9444), .B(n9445), .Z(n9440) );
  ANDN U13629 ( .B(n9446), .A(n9447), .Z(n9333) );
  IV U13630 ( .A(n9448), .Z(n9446) );
  XNOR U13631 ( .A(n9413), .B(n9412), .Z(N29381) );
  XOR U13632 ( .A(n9432), .B(n9431), .Z(n9412) );
  XNOR U13633 ( .A(n9447), .B(n9448), .Z(n9431) );
  XNOR U13634 ( .A(n9442), .B(n9443), .Z(n9448) );
  XNOR U13635 ( .A(n9444), .B(n9445), .Z(n9443) );
  XNOR U13636 ( .A(y[2908]), .B(x[2908]), .Z(n9445) );
  XNOR U13637 ( .A(y[2909]), .B(x[2909]), .Z(n9444) );
  XNOR U13638 ( .A(y[2907]), .B(x[2907]), .Z(n9442) );
  XNOR U13639 ( .A(n9436), .B(n9437), .Z(n9447) );
  XNOR U13640 ( .A(y[2904]), .B(x[2904]), .Z(n9437) );
  XNOR U13641 ( .A(n9438), .B(n9439), .Z(n9436) );
  XNOR U13642 ( .A(y[2905]), .B(x[2905]), .Z(n9439) );
  XNOR U13643 ( .A(y[2906]), .B(x[2906]), .Z(n9438) );
  XNOR U13644 ( .A(n9429), .B(n9428), .Z(n9432) );
  XNOR U13645 ( .A(n9424), .B(n9425), .Z(n9428) );
  XNOR U13646 ( .A(y[2901]), .B(x[2901]), .Z(n9425) );
  XNOR U13647 ( .A(n9426), .B(n9427), .Z(n9424) );
  XNOR U13648 ( .A(y[2902]), .B(x[2902]), .Z(n9427) );
  XNOR U13649 ( .A(y[2903]), .B(x[2903]), .Z(n9426) );
  XNOR U13650 ( .A(n9418), .B(n9419), .Z(n9429) );
  XNOR U13651 ( .A(y[2898]), .B(x[2898]), .Z(n9419) );
  XNOR U13652 ( .A(n9420), .B(n9421), .Z(n9418) );
  XNOR U13653 ( .A(y[2899]), .B(x[2899]), .Z(n9421) );
  XNOR U13654 ( .A(y[2900]), .B(x[2900]), .Z(n9420) );
  XOR U13655 ( .A(n9394), .B(n9395), .Z(n9413) );
  XNOR U13656 ( .A(n9410), .B(n9411), .Z(n9395) );
  XNOR U13657 ( .A(n9405), .B(n9406), .Z(n9411) );
  XNOR U13658 ( .A(n9407), .B(n9408), .Z(n9406) );
  XNOR U13659 ( .A(y[2896]), .B(x[2896]), .Z(n9408) );
  XNOR U13660 ( .A(y[2897]), .B(x[2897]), .Z(n9407) );
  XNOR U13661 ( .A(y[2895]), .B(x[2895]), .Z(n9405) );
  XNOR U13662 ( .A(n9399), .B(n9400), .Z(n9410) );
  XNOR U13663 ( .A(y[2892]), .B(x[2892]), .Z(n9400) );
  XNOR U13664 ( .A(n9401), .B(n9402), .Z(n9399) );
  XNOR U13665 ( .A(y[2893]), .B(x[2893]), .Z(n9402) );
  XNOR U13666 ( .A(y[2894]), .B(x[2894]), .Z(n9401) );
  XOR U13667 ( .A(n9393), .B(n9392), .Z(n9394) );
  XNOR U13668 ( .A(n9388), .B(n9389), .Z(n9392) );
  XNOR U13669 ( .A(y[2889]), .B(x[2889]), .Z(n9389) );
  XNOR U13670 ( .A(n9390), .B(n9391), .Z(n9388) );
  XNOR U13671 ( .A(y[2890]), .B(x[2890]), .Z(n9391) );
  XNOR U13672 ( .A(y[2891]), .B(x[2891]), .Z(n9390) );
  XNOR U13673 ( .A(n9382), .B(n9383), .Z(n9393) );
  XNOR U13674 ( .A(y[2886]), .B(x[2886]), .Z(n9383) );
  XNOR U13675 ( .A(n9384), .B(n9385), .Z(n9382) );
  XNOR U13676 ( .A(y[2887]), .B(x[2887]), .Z(n9385) );
  XNOR U13677 ( .A(y[2888]), .B(x[2888]), .Z(n9384) );
  NAND U13678 ( .A(n9449), .B(n9450), .Z(N29373) );
  NANDN U13679 ( .A(n9451), .B(n9452), .Z(n9450) );
  OR U13680 ( .A(n9453), .B(n9454), .Z(n9452) );
  NAND U13681 ( .A(n9453), .B(n9454), .Z(n9449) );
  XOR U13682 ( .A(n9453), .B(n9455), .Z(N29372) );
  XNOR U13683 ( .A(n9451), .B(n9454), .Z(n9455) );
  AND U13684 ( .A(n9456), .B(n9457), .Z(n9454) );
  NANDN U13685 ( .A(n9458), .B(n9459), .Z(n9457) );
  NANDN U13686 ( .A(n9460), .B(n9461), .Z(n9459) );
  NANDN U13687 ( .A(n9461), .B(n9460), .Z(n9456) );
  NAND U13688 ( .A(n9462), .B(n9463), .Z(n9451) );
  NANDN U13689 ( .A(n9464), .B(n9465), .Z(n9463) );
  OR U13690 ( .A(n9466), .B(n9467), .Z(n9465) );
  NAND U13691 ( .A(n9467), .B(n9466), .Z(n9462) );
  AND U13692 ( .A(n9468), .B(n9469), .Z(n9453) );
  NANDN U13693 ( .A(n9470), .B(n9471), .Z(n9469) );
  NANDN U13694 ( .A(n9472), .B(n9473), .Z(n9471) );
  NANDN U13695 ( .A(n9473), .B(n9472), .Z(n9468) );
  XOR U13696 ( .A(n9467), .B(n9474), .Z(N29371) );
  XOR U13697 ( .A(n9464), .B(n9466), .Z(n9474) );
  XNOR U13698 ( .A(n9460), .B(n9475), .Z(n9466) );
  XNOR U13699 ( .A(n9458), .B(n9461), .Z(n9475) );
  NAND U13700 ( .A(n9476), .B(n9477), .Z(n9461) );
  NAND U13701 ( .A(n9478), .B(n9479), .Z(n9477) );
  OR U13702 ( .A(n9480), .B(n9481), .Z(n9478) );
  NANDN U13703 ( .A(n9482), .B(n9480), .Z(n9476) );
  IV U13704 ( .A(n9481), .Z(n9482) );
  NAND U13705 ( .A(n9483), .B(n9484), .Z(n9458) );
  NAND U13706 ( .A(n9485), .B(n9486), .Z(n9484) );
  NANDN U13707 ( .A(n9487), .B(n9488), .Z(n9485) );
  NANDN U13708 ( .A(n9488), .B(n9487), .Z(n9483) );
  AND U13709 ( .A(n9489), .B(n9490), .Z(n9460) );
  NAND U13710 ( .A(n9491), .B(n9492), .Z(n9490) );
  OR U13711 ( .A(n9493), .B(n9494), .Z(n9491) );
  NANDN U13712 ( .A(n9495), .B(n9493), .Z(n9489) );
  NAND U13713 ( .A(n9496), .B(n9497), .Z(n9464) );
  NANDN U13714 ( .A(n9498), .B(n9499), .Z(n9497) );
  OR U13715 ( .A(n9500), .B(n9501), .Z(n9499) );
  NANDN U13716 ( .A(n9502), .B(n9500), .Z(n9496) );
  IV U13717 ( .A(n9501), .Z(n9502) );
  XNOR U13718 ( .A(n9472), .B(n9503), .Z(n9467) );
  XNOR U13719 ( .A(n9470), .B(n9473), .Z(n9503) );
  NAND U13720 ( .A(n9504), .B(n9505), .Z(n9473) );
  NAND U13721 ( .A(n9506), .B(n9507), .Z(n9505) );
  OR U13722 ( .A(n9508), .B(n9509), .Z(n9506) );
  NANDN U13723 ( .A(n9510), .B(n9508), .Z(n9504) );
  IV U13724 ( .A(n9509), .Z(n9510) );
  NAND U13725 ( .A(n9511), .B(n9512), .Z(n9470) );
  NAND U13726 ( .A(n9513), .B(n9514), .Z(n9512) );
  NANDN U13727 ( .A(n9515), .B(n9516), .Z(n9513) );
  NANDN U13728 ( .A(n9516), .B(n9515), .Z(n9511) );
  AND U13729 ( .A(n9517), .B(n9518), .Z(n9472) );
  NAND U13730 ( .A(n9519), .B(n9520), .Z(n9518) );
  OR U13731 ( .A(n9521), .B(n9522), .Z(n9519) );
  NANDN U13732 ( .A(n9523), .B(n9521), .Z(n9517) );
  XNOR U13733 ( .A(n9498), .B(n9524), .Z(N29370) );
  XOR U13734 ( .A(n9500), .B(n9501), .Z(n9524) );
  XNOR U13735 ( .A(n9514), .B(n9525), .Z(n9501) );
  XOR U13736 ( .A(n9515), .B(n9516), .Z(n9525) );
  XOR U13737 ( .A(n9521), .B(n9526), .Z(n9516) );
  XOR U13738 ( .A(n9520), .B(n9523), .Z(n9526) );
  IV U13739 ( .A(n9522), .Z(n9523) );
  NAND U13740 ( .A(n9527), .B(n9528), .Z(n9522) );
  OR U13741 ( .A(n9529), .B(n9530), .Z(n9528) );
  OR U13742 ( .A(n9531), .B(n9532), .Z(n9527) );
  NAND U13743 ( .A(n9533), .B(n9534), .Z(n9520) );
  OR U13744 ( .A(n9535), .B(n9536), .Z(n9534) );
  OR U13745 ( .A(n9537), .B(n9538), .Z(n9533) );
  NOR U13746 ( .A(n9539), .B(n9540), .Z(n9521) );
  ANDN U13747 ( .B(n9541), .A(n9542), .Z(n9515) );
  XNOR U13748 ( .A(n9508), .B(n9543), .Z(n9514) );
  XNOR U13749 ( .A(n9507), .B(n9509), .Z(n9543) );
  NAND U13750 ( .A(n9544), .B(n9545), .Z(n9509) );
  OR U13751 ( .A(n9546), .B(n9547), .Z(n9545) );
  OR U13752 ( .A(n9548), .B(n9549), .Z(n9544) );
  NAND U13753 ( .A(n9550), .B(n9551), .Z(n9507) );
  OR U13754 ( .A(n9552), .B(n9553), .Z(n9551) );
  OR U13755 ( .A(n9554), .B(n9555), .Z(n9550) );
  ANDN U13756 ( .B(n9556), .A(n9557), .Z(n9508) );
  IV U13757 ( .A(n9558), .Z(n9556) );
  ANDN U13758 ( .B(n9559), .A(n9560), .Z(n9500) );
  XOR U13759 ( .A(n9486), .B(n9561), .Z(n9498) );
  XOR U13760 ( .A(n9487), .B(n9488), .Z(n9561) );
  XOR U13761 ( .A(n9493), .B(n9562), .Z(n9488) );
  XOR U13762 ( .A(n9492), .B(n9495), .Z(n9562) );
  IV U13763 ( .A(n9494), .Z(n9495) );
  NAND U13764 ( .A(n9563), .B(n9564), .Z(n9494) );
  OR U13765 ( .A(n9565), .B(n9566), .Z(n9564) );
  OR U13766 ( .A(n9567), .B(n9568), .Z(n9563) );
  NAND U13767 ( .A(n9569), .B(n9570), .Z(n9492) );
  OR U13768 ( .A(n9571), .B(n9572), .Z(n9570) );
  OR U13769 ( .A(n9573), .B(n9574), .Z(n9569) );
  NOR U13770 ( .A(n9575), .B(n9576), .Z(n9493) );
  ANDN U13771 ( .B(n9577), .A(n9578), .Z(n9487) );
  IV U13772 ( .A(n9579), .Z(n9577) );
  XNOR U13773 ( .A(n9480), .B(n9580), .Z(n9486) );
  XNOR U13774 ( .A(n9479), .B(n9481), .Z(n9580) );
  NAND U13775 ( .A(n9581), .B(n9582), .Z(n9481) );
  OR U13776 ( .A(n9583), .B(n9584), .Z(n9582) );
  OR U13777 ( .A(n9585), .B(n9586), .Z(n9581) );
  NAND U13778 ( .A(n9587), .B(n9588), .Z(n9479) );
  OR U13779 ( .A(n9589), .B(n9590), .Z(n9588) );
  OR U13780 ( .A(n9591), .B(n9592), .Z(n9587) );
  ANDN U13781 ( .B(n9593), .A(n9594), .Z(n9480) );
  IV U13782 ( .A(n9595), .Z(n9593) );
  XNOR U13783 ( .A(n9560), .B(n9559), .Z(N29369) );
  XOR U13784 ( .A(n9579), .B(n9578), .Z(n9559) );
  XNOR U13785 ( .A(n9594), .B(n9595), .Z(n9578) );
  XNOR U13786 ( .A(n9589), .B(n9590), .Z(n9595) );
  XNOR U13787 ( .A(n9591), .B(n9592), .Z(n9590) );
  XNOR U13788 ( .A(y[2884]), .B(x[2884]), .Z(n9592) );
  XNOR U13789 ( .A(y[2885]), .B(x[2885]), .Z(n9591) );
  XNOR U13790 ( .A(y[2883]), .B(x[2883]), .Z(n9589) );
  XNOR U13791 ( .A(n9583), .B(n9584), .Z(n9594) );
  XNOR U13792 ( .A(y[2880]), .B(x[2880]), .Z(n9584) );
  XNOR U13793 ( .A(n9585), .B(n9586), .Z(n9583) );
  XNOR U13794 ( .A(y[2881]), .B(x[2881]), .Z(n9586) );
  XNOR U13795 ( .A(y[2882]), .B(x[2882]), .Z(n9585) );
  XNOR U13796 ( .A(n9576), .B(n9575), .Z(n9579) );
  XNOR U13797 ( .A(n9571), .B(n9572), .Z(n9575) );
  XNOR U13798 ( .A(y[2877]), .B(x[2877]), .Z(n9572) );
  XNOR U13799 ( .A(n9573), .B(n9574), .Z(n9571) );
  XNOR U13800 ( .A(y[2878]), .B(x[2878]), .Z(n9574) );
  XNOR U13801 ( .A(y[2879]), .B(x[2879]), .Z(n9573) );
  XNOR U13802 ( .A(n9565), .B(n9566), .Z(n9576) );
  XNOR U13803 ( .A(y[2874]), .B(x[2874]), .Z(n9566) );
  XNOR U13804 ( .A(n9567), .B(n9568), .Z(n9565) );
  XNOR U13805 ( .A(y[2875]), .B(x[2875]), .Z(n9568) );
  XNOR U13806 ( .A(y[2876]), .B(x[2876]), .Z(n9567) );
  XOR U13807 ( .A(n9541), .B(n9542), .Z(n9560) );
  XNOR U13808 ( .A(n9557), .B(n9558), .Z(n9542) );
  XNOR U13809 ( .A(n9552), .B(n9553), .Z(n9558) );
  XNOR U13810 ( .A(n9554), .B(n9555), .Z(n9553) );
  XNOR U13811 ( .A(y[2872]), .B(x[2872]), .Z(n9555) );
  XNOR U13812 ( .A(y[2873]), .B(x[2873]), .Z(n9554) );
  XNOR U13813 ( .A(y[2871]), .B(x[2871]), .Z(n9552) );
  XNOR U13814 ( .A(n9546), .B(n9547), .Z(n9557) );
  XNOR U13815 ( .A(y[2868]), .B(x[2868]), .Z(n9547) );
  XNOR U13816 ( .A(n9548), .B(n9549), .Z(n9546) );
  XNOR U13817 ( .A(y[2869]), .B(x[2869]), .Z(n9549) );
  XNOR U13818 ( .A(y[2870]), .B(x[2870]), .Z(n9548) );
  XOR U13819 ( .A(n9540), .B(n9539), .Z(n9541) );
  XNOR U13820 ( .A(n9535), .B(n9536), .Z(n9539) );
  XNOR U13821 ( .A(y[2865]), .B(x[2865]), .Z(n9536) );
  XNOR U13822 ( .A(n9537), .B(n9538), .Z(n9535) );
  XNOR U13823 ( .A(y[2866]), .B(x[2866]), .Z(n9538) );
  XNOR U13824 ( .A(y[2867]), .B(x[2867]), .Z(n9537) );
  XNOR U13825 ( .A(n9529), .B(n9530), .Z(n9540) );
  XNOR U13826 ( .A(y[2862]), .B(x[2862]), .Z(n9530) );
  XNOR U13827 ( .A(n9531), .B(n9532), .Z(n9529) );
  XNOR U13828 ( .A(y[2863]), .B(x[2863]), .Z(n9532) );
  XNOR U13829 ( .A(y[2864]), .B(x[2864]), .Z(n9531) );
  NAND U13830 ( .A(n9596), .B(n9597), .Z(N29361) );
  NANDN U13831 ( .A(n9598), .B(n9599), .Z(n9597) );
  OR U13832 ( .A(n9600), .B(n9601), .Z(n9599) );
  NAND U13833 ( .A(n9600), .B(n9601), .Z(n9596) );
  XOR U13834 ( .A(n9600), .B(n9602), .Z(N29360) );
  XNOR U13835 ( .A(n9598), .B(n9601), .Z(n9602) );
  AND U13836 ( .A(n9603), .B(n9604), .Z(n9601) );
  NANDN U13837 ( .A(n9605), .B(n9606), .Z(n9604) );
  NANDN U13838 ( .A(n9607), .B(n9608), .Z(n9606) );
  NANDN U13839 ( .A(n9608), .B(n9607), .Z(n9603) );
  NAND U13840 ( .A(n9609), .B(n9610), .Z(n9598) );
  NANDN U13841 ( .A(n9611), .B(n9612), .Z(n9610) );
  OR U13842 ( .A(n9613), .B(n9614), .Z(n9612) );
  NAND U13843 ( .A(n9614), .B(n9613), .Z(n9609) );
  AND U13844 ( .A(n9615), .B(n9616), .Z(n9600) );
  NANDN U13845 ( .A(n9617), .B(n9618), .Z(n9616) );
  NANDN U13846 ( .A(n9619), .B(n9620), .Z(n9618) );
  NANDN U13847 ( .A(n9620), .B(n9619), .Z(n9615) );
  XOR U13848 ( .A(n9614), .B(n9621), .Z(N29359) );
  XOR U13849 ( .A(n9611), .B(n9613), .Z(n9621) );
  XNOR U13850 ( .A(n9607), .B(n9622), .Z(n9613) );
  XNOR U13851 ( .A(n9605), .B(n9608), .Z(n9622) );
  NAND U13852 ( .A(n9623), .B(n9624), .Z(n9608) );
  NAND U13853 ( .A(n9625), .B(n9626), .Z(n9624) );
  OR U13854 ( .A(n9627), .B(n9628), .Z(n9625) );
  NANDN U13855 ( .A(n9629), .B(n9627), .Z(n9623) );
  IV U13856 ( .A(n9628), .Z(n9629) );
  NAND U13857 ( .A(n9630), .B(n9631), .Z(n9605) );
  NAND U13858 ( .A(n9632), .B(n9633), .Z(n9631) );
  NANDN U13859 ( .A(n9634), .B(n9635), .Z(n9632) );
  NANDN U13860 ( .A(n9635), .B(n9634), .Z(n9630) );
  AND U13861 ( .A(n9636), .B(n9637), .Z(n9607) );
  NAND U13862 ( .A(n9638), .B(n9639), .Z(n9637) );
  OR U13863 ( .A(n9640), .B(n9641), .Z(n9638) );
  NANDN U13864 ( .A(n9642), .B(n9640), .Z(n9636) );
  NAND U13865 ( .A(n9643), .B(n9644), .Z(n9611) );
  NANDN U13866 ( .A(n9645), .B(n9646), .Z(n9644) );
  OR U13867 ( .A(n9647), .B(n9648), .Z(n9646) );
  NANDN U13868 ( .A(n9649), .B(n9647), .Z(n9643) );
  IV U13869 ( .A(n9648), .Z(n9649) );
  XNOR U13870 ( .A(n9619), .B(n9650), .Z(n9614) );
  XNOR U13871 ( .A(n9617), .B(n9620), .Z(n9650) );
  NAND U13872 ( .A(n9651), .B(n9652), .Z(n9620) );
  NAND U13873 ( .A(n9653), .B(n9654), .Z(n9652) );
  OR U13874 ( .A(n9655), .B(n9656), .Z(n9653) );
  NANDN U13875 ( .A(n9657), .B(n9655), .Z(n9651) );
  IV U13876 ( .A(n9656), .Z(n9657) );
  NAND U13877 ( .A(n9658), .B(n9659), .Z(n9617) );
  NAND U13878 ( .A(n9660), .B(n9661), .Z(n9659) );
  NANDN U13879 ( .A(n9662), .B(n9663), .Z(n9660) );
  NANDN U13880 ( .A(n9663), .B(n9662), .Z(n9658) );
  AND U13881 ( .A(n9664), .B(n9665), .Z(n9619) );
  NAND U13882 ( .A(n9666), .B(n9667), .Z(n9665) );
  OR U13883 ( .A(n9668), .B(n9669), .Z(n9666) );
  NANDN U13884 ( .A(n9670), .B(n9668), .Z(n9664) );
  XNOR U13885 ( .A(n9645), .B(n9671), .Z(N29358) );
  XOR U13886 ( .A(n9647), .B(n9648), .Z(n9671) );
  XNOR U13887 ( .A(n9661), .B(n9672), .Z(n9648) );
  XOR U13888 ( .A(n9662), .B(n9663), .Z(n9672) );
  XOR U13889 ( .A(n9668), .B(n9673), .Z(n9663) );
  XOR U13890 ( .A(n9667), .B(n9670), .Z(n9673) );
  IV U13891 ( .A(n9669), .Z(n9670) );
  NAND U13892 ( .A(n9674), .B(n9675), .Z(n9669) );
  OR U13893 ( .A(n9676), .B(n9677), .Z(n9675) );
  OR U13894 ( .A(n9678), .B(n9679), .Z(n9674) );
  NAND U13895 ( .A(n9680), .B(n9681), .Z(n9667) );
  OR U13896 ( .A(n9682), .B(n9683), .Z(n9681) );
  OR U13897 ( .A(n9684), .B(n9685), .Z(n9680) );
  NOR U13898 ( .A(n9686), .B(n9687), .Z(n9668) );
  ANDN U13899 ( .B(n9688), .A(n9689), .Z(n9662) );
  XNOR U13900 ( .A(n9655), .B(n9690), .Z(n9661) );
  XNOR U13901 ( .A(n9654), .B(n9656), .Z(n9690) );
  NAND U13902 ( .A(n9691), .B(n9692), .Z(n9656) );
  OR U13903 ( .A(n9693), .B(n9694), .Z(n9692) );
  OR U13904 ( .A(n9695), .B(n9696), .Z(n9691) );
  NAND U13905 ( .A(n9697), .B(n9698), .Z(n9654) );
  OR U13906 ( .A(n9699), .B(n9700), .Z(n9698) );
  OR U13907 ( .A(n9701), .B(n9702), .Z(n9697) );
  ANDN U13908 ( .B(n9703), .A(n9704), .Z(n9655) );
  IV U13909 ( .A(n9705), .Z(n9703) );
  ANDN U13910 ( .B(n9706), .A(n9707), .Z(n9647) );
  XOR U13911 ( .A(n9633), .B(n9708), .Z(n9645) );
  XOR U13912 ( .A(n9634), .B(n9635), .Z(n9708) );
  XOR U13913 ( .A(n9640), .B(n9709), .Z(n9635) );
  XOR U13914 ( .A(n9639), .B(n9642), .Z(n9709) );
  IV U13915 ( .A(n9641), .Z(n9642) );
  NAND U13916 ( .A(n9710), .B(n9711), .Z(n9641) );
  OR U13917 ( .A(n9712), .B(n9713), .Z(n9711) );
  OR U13918 ( .A(n9714), .B(n9715), .Z(n9710) );
  NAND U13919 ( .A(n9716), .B(n9717), .Z(n9639) );
  OR U13920 ( .A(n9718), .B(n9719), .Z(n9717) );
  OR U13921 ( .A(n9720), .B(n9721), .Z(n9716) );
  NOR U13922 ( .A(n9722), .B(n9723), .Z(n9640) );
  ANDN U13923 ( .B(n9724), .A(n9725), .Z(n9634) );
  IV U13924 ( .A(n9726), .Z(n9724) );
  XNOR U13925 ( .A(n9627), .B(n9727), .Z(n9633) );
  XNOR U13926 ( .A(n9626), .B(n9628), .Z(n9727) );
  NAND U13927 ( .A(n9728), .B(n9729), .Z(n9628) );
  OR U13928 ( .A(n9730), .B(n9731), .Z(n9729) );
  OR U13929 ( .A(n9732), .B(n9733), .Z(n9728) );
  NAND U13930 ( .A(n9734), .B(n9735), .Z(n9626) );
  OR U13931 ( .A(n9736), .B(n9737), .Z(n9735) );
  OR U13932 ( .A(n9738), .B(n9739), .Z(n9734) );
  ANDN U13933 ( .B(n9740), .A(n9741), .Z(n9627) );
  IV U13934 ( .A(n9742), .Z(n9740) );
  XNOR U13935 ( .A(n9707), .B(n9706), .Z(N29357) );
  XOR U13936 ( .A(n9726), .B(n9725), .Z(n9706) );
  XNOR U13937 ( .A(n9741), .B(n9742), .Z(n9725) );
  XNOR U13938 ( .A(n9736), .B(n9737), .Z(n9742) );
  XNOR U13939 ( .A(n9738), .B(n9739), .Z(n9737) );
  XNOR U13940 ( .A(y[2860]), .B(x[2860]), .Z(n9739) );
  XNOR U13941 ( .A(y[2861]), .B(x[2861]), .Z(n9738) );
  XNOR U13942 ( .A(y[2859]), .B(x[2859]), .Z(n9736) );
  XNOR U13943 ( .A(n9730), .B(n9731), .Z(n9741) );
  XNOR U13944 ( .A(y[2856]), .B(x[2856]), .Z(n9731) );
  XNOR U13945 ( .A(n9732), .B(n9733), .Z(n9730) );
  XNOR U13946 ( .A(y[2857]), .B(x[2857]), .Z(n9733) );
  XNOR U13947 ( .A(y[2858]), .B(x[2858]), .Z(n9732) );
  XNOR U13948 ( .A(n9723), .B(n9722), .Z(n9726) );
  XNOR U13949 ( .A(n9718), .B(n9719), .Z(n9722) );
  XNOR U13950 ( .A(y[2853]), .B(x[2853]), .Z(n9719) );
  XNOR U13951 ( .A(n9720), .B(n9721), .Z(n9718) );
  XNOR U13952 ( .A(y[2854]), .B(x[2854]), .Z(n9721) );
  XNOR U13953 ( .A(y[2855]), .B(x[2855]), .Z(n9720) );
  XNOR U13954 ( .A(n9712), .B(n9713), .Z(n9723) );
  XNOR U13955 ( .A(y[2850]), .B(x[2850]), .Z(n9713) );
  XNOR U13956 ( .A(n9714), .B(n9715), .Z(n9712) );
  XNOR U13957 ( .A(y[2851]), .B(x[2851]), .Z(n9715) );
  XNOR U13958 ( .A(y[2852]), .B(x[2852]), .Z(n9714) );
  XOR U13959 ( .A(n9688), .B(n9689), .Z(n9707) );
  XNOR U13960 ( .A(n9704), .B(n9705), .Z(n9689) );
  XNOR U13961 ( .A(n9699), .B(n9700), .Z(n9705) );
  XNOR U13962 ( .A(n9701), .B(n9702), .Z(n9700) );
  XNOR U13963 ( .A(y[2848]), .B(x[2848]), .Z(n9702) );
  XNOR U13964 ( .A(y[2849]), .B(x[2849]), .Z(n9701) );
  XNOR U13965 ( .A(y[2847]), .B(x[2847]), .Z(n9699) );
  XNOR U13966 ( .A(n9693), .B(n9694), .Z(n9704) );
  XNOR U13967 ( .A(y[2844]), .B(x[2844]), .Z(n9694) );
  XNOR U13968 ( .A(n9695), .B(n9696), .Z(n9693) );
  XNOR U13969 ( .A(y[2845]), .B(x[2845]), .Z(n9696) );
  XNOR U13970 ( .A(y[2846]), .B(x[2846]), .Z(n9695) );
  XOR U13971 ( .A(n9687), .B(n9686), .Z(n9688) );
  XNOR U13972 ( .A(n9682), .B(n9683), .Z(n9686) );
  XNOR U13973 ( .A(y[2841]), .B(x[2841]), .Z(n9683) );
  XNOR U13974 ( .A(n9684), .B(n9685), .Z(n9682) );
  XNOR U13975 ( .A(y[2842]), .B(x[2842]), .Z(n9685) );
  XNOR U13976 ( .A(y[2843]), .B(x[2843]), .Z(n9684) );
  XNOR U13977 ( .A(n9676), .B(n9677), .Z(n9687) );
  XNOR U13978 ( .A(y[2838]), .B(x[2838]), .Z(n9677) );
  XNOR U13979 ( .A(n9678), .B(n9679), .Z(n9676) );
  XNOR U13980 ( .A(y[2839]), .B(x[2839]), .Z(n9679) );
  XNOR U13981 ( .A(y[2840]), .B(x[2840]), .Z(n9678) );
  NAND U13982 ( .A(n9743), .B(n9744), .Z(N29349) );
  NANDN U13983 ( .A(n9745), .B(n9746), .Z(n9744) );
  OR U13984 ( .A(n9747), .B(n9748), .Z(n9746) );
  NAND U13985 ( .A(n9747), .B(n9748), .Z(n9743) );
  XOR U13986 ( .A(n9747), .B(n9749), .Z(N29348) );
  XNOR U13987 ( .A(n9745), .B(n9748), .Z(n9749) );
  AND U13988 ( .A(n9750), .B(n9751), .Z(n9748) );
  NANDN U13989 ( .A(n9752), .B(n9753), .Z(n9751) );
  NANDN U13990 ( .A(n9754), .B(n9755), .Z(n9753) );
  NANDN U13991 ( .A(n9755), .B(n9754), .Z(n9750) );
  NAND U13992 ( .A(n9756), .B(n9757), .Z(n9745) );
  NANDN U13993 ( .A(n9758), .B(n9759), .Z(n9757) );
  OR U13994 ( .A(n9760), .B(n9761), .Z(n9759) );
  NAND U13995 ( .A(n9761), .B(n9760), .Z(n9756) );
  AND U13996 ( .A(n9762), .B(n9763), .Z(n9747) );
  NANDN U13997 ( .A(n9764), .B(n9765), .Z(n9763) );
  NANDN U13998 ( .A(n9766), .B(n9767), .Z(n9765) );
  NANDN U13999 ( .A(n9767), .B(n9766), .Z(n9762) );
  XOR U14000 ( .A(n9761), .B(n9768), .Z(N29347) );
  XOR U14001 ( .A(n9758), .B(n9760), .Z(n9768) );
  XNOR U14002 ( .A(n9754), .B(n9769), .Z(n9760) );
  XNOR U14003 ( .A(n9752), .B(n9755), .Z(n9769) );
  NAND U14004 ( .A(n9770), .B(n9771), .Z(n9755) );
  NAND U14005 ( .A(n9772), .B(n9773), .Z(n9771) );
  OR U14006 ( .A(n9774), .B(n9775), .Z(n9772) );
  NANDN U14007 ( .A(n9776), .B(n9774), .Z(n9770) );
  IV U14008 ( .A(n9775), .Z(n9776) );
  NAND U14009 ( .A(n9777), .B(n9778), .Z(n9752) );
  NAND U14010 ( .A(n9779), .B(n9780), .Z(n9778) );
  NANDN U14011 ( .A(n9781), .B(n9782), .Z(n9779) );
  NANDN U14012 ( .A(n9782), .B(n9781), .Z(n9777) );
  AND U14013 ( .A(n9783), .B(n9784), .Z(n9754) );
  NAND U14014 ( .A(n9785), .B(n9786), .Z(n9784) );
  OR U14015 ( .A(n9787), .B(n9788), .Z(n9785) );
  NANDN U14016 ( .A(n9789), .B(n9787), .Z(n9783) );
  NAND U14017 ( .A(n9790), .B(n9791), .Z(n9758) );
  NANDN U14018 ( .A(n9792), .B(n9793), .Z(n9791) );
  OR U14019 ( .A(n9794), .B(n9795), .Z(n9793) );
  NANDN U14020 ( .A(n9796), .B(n9794), .Z(n9790) );
  IV U14021 ( .A(n9795), .Z(n9796) );
  XNOR U14022 ( .A(n9766), .B(n9797), .Z(n9761) );
  XNOR U14023 ( .A(n9764), .B(n9767), .Z(n9797) );
  NAND U14024 ( .A(n9798), .B(n9799), .Z(n9767) );
  NAND U14025 ( .A(n9800), .B(n9801), .Z(n9799) );
  OR U14026 ( .A(n9802), .B(n9803), .Z(n9800) );
  NANDN U14027 ( .A(n9804), .B(n9802), .Z(n9798) );
  IV U14028 ( .A(n9803), .Z(n9804) );
  NAND U14029 ( .A(n9805), .B(n9806), .Z(n9764) );
  NAND U14030 ( .A(n9807), .B(n9808), .Z(n9806) );
  NANDN U14031 ( .A(n9809), .B(n9810), .Z(n9807) );
  NANDN U14032 ( .A(n9810), .B(n9809), .Z(n9805) );
  AND U14033 ( .A(n9811), .B(n9812), .Z(n9766) );
  NAND U14034 ( .A(n9813), .B(n9814), .Z(n9812) );
  OR U14035 ( .A(n9815), .B(n9816), .Z(n9813) );
  NANDN U14036 ( .A(n9817), .B(n9815), .Z(n9811) );
  XNOR U14037 ( .A(n9792), .B(n9818), .Z(N29346) );
  XOR U14038 ( .A(n9794), .B(n9795), .Z(n9818) );
  XNOR U14039 ( .A(n9808), .B(n9819), .Z(n9795) );
  XOR U14040 ( .A(n9809), .B(n9810), .Z(n9819) );
  XOR U14041 ( .A(n9815), .B(n9820), .Z(n9810) );
  XOR U14042 ( .A(n9814), .B(n9817), .Z(n9820) );
  IV U14043 ( .A(n9816), .Z(n9817) );
  NAND U14044 ( .A(n9821), .B(n9822), .Z(n9816) );
  OR U14045 ( .A(n9823), .B(n9824), .Z(n9822) );
  OR U14046 ( .A(n9825), .B(n9826), .Z(n9821) );
  NAND U14047 ( .A(n9827), .B(n9828), .Z(n9814) );
  OR U14048 ( .A(n9829), .B(n9830), .Z(n9828) );
  OR U14049 ( .A(n9831), .B(n9832), .Z(n9827) );
  NOR U14050 ( .A(n9833), .B(n9834), .Z(n9815) );
  ANDN U14051 ( .B(n9835), .A(n9836), .Z(n9809) );
  XNOR U14052 ( .A(n9802), .B(n9837), .Z(n9808) );
  XNOR U14053 ( .A(n9801), .B(n9803), .Z(n9837) );
  NAND U14054 ( .A(n9838), .B(n9839), .Z(n9803) );
  OR U14055 ( .A(n9840), .B(n9841), .Z(n9839) );
  OR U14056 ( .A(n9842), .B(n9843), .Z(n9838) );
  NAND U14057 ( .A(n9844), .B(n9845), .Z(n9801) );
  OR U14058 ( .A(n9846), .B(n9847), .Z(n9845) );
  OR U14059 ( .A(n9848), .B(n9849), .Z(n9844) );
  ANDN U14060 ( .B(n9850), .A(n9851), .Z(n9802) );
  IV U14061 ( .A(n9852), .Z(n9850) );
  ANDN U14062 ( .B(n9853), .A(n9854), .Z(n9794) );
  XOR U14063 ( .A(n9780), .B(n9855), .Z(n9792) );
  XOR U14064 ( .A(n9781), .B(n9782), .Z(n9855) );
  XOR U14065 ( .A(n9787), .B(n9856), .Z(n9782) );
  XOR U14066 ( .A(n9786), .B(n9789), .Z(n9856) );
  IV U14067 ( .A(n9788), .Z(n9789) );
  NAND U14068 ( .A(n9857), .B(n9858), .Z(n9788) );
  OR U14069 ( .A(n9859), .B(n9860), .Z(n9858) );
  OR U14070 ( .A(n9861), .B(n9862), .Z(n9857) );
  NAND U14071 ( .A(n9863), .B(n9864), .Z(n9786) );
  OR U14072 ( .A(n9865), .B(n9866), .Z(n9864) );
  OR U14073 ( .A(n9867), .B(n9868), .Z(n9863) );
  NOR U14074 ( .A(n9869), .B(n9870), .Z(n9787) );
  ANDN U14075 ( .B(n9871), .A(n9872), .Z(n9781) );
  IV U14076 ( .A(n9873), .Z(n9871) );
  XNOR U14077 ( .A(n9774), .B(n9874), .Z(n9780) );
  XNOR U14078 ( .A(n9773), .B(n9775), .Z(n9874) );
  NAND U14079 ( .A(n9875), .B(n9876), .Z(n9775) );
  OR U14080 ( .A(n9877), .B(n9878), .Z(n9876) );
  OR U14081 ( .A(n9879), .B(n9880), .Z(n9875) );
  NAND U14082 ( .A(n9881), .B(n9882), .Z(n9773) );
  OR U14083 ( .A(n9883), .B(n9884), .Z(n9882) );
  OR U14084 ( .A(n9885), .B(n9886), .Z(n9881) );
  ANDN U14085 ( .B(n9887), .A(n9888), .Z(n9774) );
  IV U14086 ( .A(n9889), .Z(n9887) );
  XNOR U14087 ( .A(n9854), .B(n9853), .Z(N29345) );
  XOR U14088 ( .A(n9873), .B(n9872), .Z(n9853) );
  XNOR U14089 ( .A(n9888), .B(n9889), .Z(n9872) );
  XNOR U14090 ( .A(n9883), .B(n9884), .Z(n9889) );
  XNOR U14091 ( .A(n9885), .B(n9886), .Z(n9884) );
  XNOR U14092 ( .A(y[2836]), .B(x[2836]), .Z(n9886) );
  XNOR U14093 ( .A(y[2837]), .B(x[2837]), .Z(n9885) );
  XNOR U14094 ( .A(y[2835]), .B(x[2835]), .Z(n9883) );
  XNOR U14095 ( .A(n9877), .B(n9878), .Z(n9888) );
  XNOR U14096 ( .A(y[2832]), .B(x[2832]), .Z(n9878) );
  XNOR U14097 ( .A(n9879), .B(n9880), .Z(n9877) );
  XNOR U14098 ( .A(y[2833]), .B(x[2833]), .Z(n9880) );
  XNOR U14099 ( .A(y[2834]), .B(x[2834]), .Z(n9879) );
  XNOR U14100 ( .A(n9870), .B(n9869), .Z(n9873) );
  XNOR U14101 ( .A(n9865), .B(n9866), .Z(n9869) );
  XNOR U14102 ( .A(y[2829]), .B(x[2829]), .Z(n9866) );
  XNOR U14103 ( .A(n9867), .B(n9868), .Z(n9865) );
  XNOR U14104 ( .A(y[2830]), .B(x[2830]), .Z(n9868) );
  XNOR U14105 ( .A(y[2831]), .B(x[2831]), .Z(n9867) );
  XNOR U14106 ( .A(n9859), .B(n9860), .Z(n9870) );
  XNOR U14107 ( .A(y[2826]), .B(x[2826]), .Z(n9860) );
  XNOR U14108 ( .A(n9861), .B(n9862), .Z(n9859) );
  XNOR U14109 ( .A(y[2827]), .B(x[2827]), .Z(n9862) );
  XNOR U14110 ( .A(y[2828]), .B(x[2828]), .Z(n9861) );
  XOR U14111 ( .A(n9835), .B(n9836), .Z(n9854) );
  XNOR U14112 ( .A(n9851), .B(n9852), .Z(n9836) );
  XNOR U14113 ( .A(n9846), .B(n9847), .Z(n9852) );
  XNOR U14114 ( .A(n9848), .B(n9849), .Z(n9847) );
  XNOR U14115 ( .A(y[2824]), .B(x[2824]), .Z(n9849) );
  XNOR U14116 ( .A(y[2825]), .B(x[2825]), .Z(n9848) );
  XNOR U14117 ( .A(y[2823]), .B(x[2823]), .Z(n9846) );
  XNOR U14118 ( .A(n9840), .B(n9841), .Z(n9851) );
  XNOR U14119 ( .A(y[2820]), .B(x[2820]), .Z(n9841) );
  XNOR U14120 ( .A(n9842), .B(n9843), .Z(n9840) );
  XNOR U14121 ( .A(y[2821]), .B(x[2821]), .Z(n9843) );
  XNOR U14122 ( .A(y[2822]), .B(x[2822]), .Z(n9842) );
  XOR U14123 ( .A(n9834), .B(n9833), .Z(n9835) );
  XNOR U14124 ( .A(n9829), .B(n9830), .Z(n9833) );
  XNOR U14125 ( .A(y[2817]), .B(x[2817]), .Z(n9830) );
  XNOR U14126 ( .A(n9831), .B(n9832), .Z(n9829) );
  XNOR U14127 ( .A(y[2818]), .B(x[2818]), .Z(n9832) );
  XNOR U14128 ( .A(y[2819]), .B(x[2819]), .Z(n9831) );
  XNOR U14129 ( .A(n9823), .B(n9824), .Z(n9834) );
  XNOR U14130 ( .A(y[2814]), .B(x[2814]), .Z(n9824) );
  XNOR U14131 ( .A(n9825), .B(n9826), .Z(n9823) );
  XNOR U14132 ( .A(y[2815]), .B(x[2815]), .Z(n9826) );
  XNOR U14133 ( .A(y[2816]), .B(x[2816]), .Z(n9825) );
  NAND U14134 ( .A(n9890), .B(n9891), .Z(N29337) );
  NANDN U14135 ( .A(n9892), .B(n9893), .Z(n9891) );
  OR U14136 ( .A(n9894), .B(n9895), .Z(n9893) );
  NAND U14137 ( .A(n9894), .B(n9895), .Z(n9890) );
  XOR U14138 ( .A(n9894), .B(n9896), .Z(N29336) );
  XNOR U14139 ( .A(n9892), .B(n9895), .Z(n9896) );
  AND U14140 ( .A(n9897), .B(n9898), .Z(n9895) );
  NANDN U14141 ( .A(n9899), .B(n9900), .Z(n9898) );
  NANDN U14142 ( .A(n9901), .B(n9902), .Z(n9900) );
  NANDN U14143 ( .A(n9902), .B(n9901), .Z(n9897) );
  NAND U14144 ( .A(n9903), .B(n9904), .Z(n9892) );
  NANDN U14145 ( .A(n9905), .B(n9906), .Z(n9904) );
  OR U14146 ( .A(n9907), .B(n9908), .Z(n9906) );
  NAND U14147 ( .A(n9908), .B(n9907), .Z(n9903) );
  AND U14148 ( .A(n9909), .B(n9910), .Z(n9894) );
  NANDN U14149 ( .A(n9911), .B(n9912), .Z(n9910) );
  NANDN U14150 ( .A(n9913), .B(n9914), .Z(n9912) );
  NANDN U14151 ( .A(n9914), .B(n9913), .Z(n9909) );
  XOR U14152 ( .A(n9908), .B(n9915), .Z(N29335) );
  XOR U14153 ( .A(n9905), .B(n9907), .Z(n9915) );
  XNOR U14154 ( .A(n9901), .B(n9916), .Z(n9907) );
  XNOR U14155 ( .A(n9899), .B(n9902), .Z(n9916) );
  NAND U14156 ( .A(n9917), .B(n9918), .Z(n9902) );
  NAND U14157 ( .A(n9919), .B(n9920), .Z(n9918) );
  OR U14158 ( .A(n9921), .B(n9922), .Z(n9919) );
  NANDN U14159 ( .A(n9923), .B(n9921), .Z(n9917) );
  IV U14160 ( .A(n9922), .Z(n9923) );
  NAND U14161 ( .A(n9924), .B(n9925), .Z(n9899) );
  NAND U14162 ( .A(n9926), .B(n9927), .Z(n9925) );
  NANDN U14163 ( .A(n9928), .B(n9929), .Z(n9926) );
  NANDN U14164 ( .A(n9929), .B(n9928), .Z(n9924) );
  AND U14165 ( .A(n9930), .B(n9931), .Z(n9901) );
  NAND U14166 ( .A(n9932), .B(n9933), .Z(n9931) );
  OR U14167 ( .A(n9934), .B(n9935), .Z(n9932) );
  NANDN U14168 ( .A(n9936), .B(n9934), .Z(n9930) );
  NAND U14169 ( .A(n9937), .B(n9938), .Z(n9905) );
  NANDN U14170 ( .A(n9939), .B(n9940), .Z(n9938) );
  OR U14171 ( .A(n9941), .B(n9942), .Z(n9940) );
  NANDN U14172 ( .A(n9943), .B(n9941), .Z(n9937) );
  IV U14173 ( .A(n9942), .Z(n9943) );
  XNOR U14174 ( .A(n9913), .B(n9944), .Z(n9908) );
  XNOR U14175 ( .A(n9911), .B(n9914), .Z(n9944) );
  NAND U14176 ( .A(n9945), .B(n9946), .Z(n9914) );
  NAND U14177 ( .A(n9947), .B(n9948), .Z(n9946) );
  OR U14178 ( .A(n9949), .B(n9950), .Z(n9947) );
  NANDN U14179 ( .A(n9951), .B(n9949), .Z(n9945) );
  IV U14180 ( .A(n9950), .Z(n9951) );
  NAND U14181 ( .A(n9952), .B(n9953), .Z(n9911) );
  NAND U14182 ( .A(n9954), .B(n9955), .Z(n9953) );
  NANDN U14183 ( .A(n9956), .B(n9957), .Z(n9954) );
  NANDN U14184 ( .A(n9957), .B(n9956), .Z(n9952) );
  AND U14185 ( .A(n9958), .B(n9959), .Z(n9913) );
  NAND U14186 ( .A(n9960), .B(n9961), .Z(n9959) );
  OR U14187 ( .A(n9962), .B(n9963), .Z(n9960) );
  NANDN U14188 ( .A(n9964), .B(n9962), .Z(n9958) );
  XNOR U14189 ( .A(n9939), .B(n9965), .Z(N29334) );
  XOR U14190 ( .A(n9941), .B(n9942), .Z(n9965) );
  XNOR U14191 ( .A(n9955), .B(n9966), .Z(n9942) );
  XOR U14192 ( .A(n9956), .B(n9957), .Z(n9966) );
  XOR U14193 ( .A(n9962), .B(n9967), .Z(n9957) );
  XOR U14194 ( .A(n9961), .B(n9964), .Z(n9967) );
  IV U14195 ( .A(n9963), .Z(n9964) );
  NAND U14196 ( .A(n9968), .B(n9969), .Z(n9963) );
  OR U14197 ( .A(n9970), .B(n9971), .Z(n9969) );
  OR U14198 ( .A(n9972), .B(n9973), .Z(n9968) );
  NAND U14199 ( .A(n9974), .B(n9975), .Z(n9961) );
  OR U14200 ( .A(n9976), .B(n9977), .Z(n9975) );
  OR U14201 ( .A(n9978), .B(n9979), .Z(n9974) );
  NOR U14202 ( .A(n9980), .B(n9981), .Z(n9962) );
  ANDN U14203 ( .B(n9982), .A(n9983), .Z(n9956) );
  XNOR U14204 ( .A(n9949), .B(n9984), .Z(n9955) );
  XNOR U14205 ( .A(n9948), .B(n9950), .Z(n9984) );
  NAND U14206 ( .A(n9985), .B(n9986), .Z(n9950) );
  OR U14207 ( .A(n9987), .B(n9988), .Z(n9986) );
  OR U14208 ( .A(n9989), .B(n9990), .Z(n9985) );
  NAND U14209 ( .A(n9991), .B(n9992), .Z(n9948) );
  OR U14210 ( .A(n9993), .B(n9994), .Z(n9992) );
  OR U14211 ( .A(n9995), .B(n9996), .Z(n9991) );
  ANDN U14212 ( .B(n9997), .A(n9998), .Z(n9949) );
  IV U14213 ( .A(n9999), .Z(n9997) );
  ANDN U14214 ( .B(n10000), .A(n10001), .Z(n9941) );
  XOR U14215 ( .A(n9927), .B(n10002), .Z(n9939) );
  XOR U14216 ( .A(n9928), .B(n9929), .Z(n10002) );
  XOR U14217 ( .A(n9934), .B(n10003), .Z(n9929) );
  XOR U14218 ( .A(n9933), .B(n9936), .Z(n10003) );
  IV U14219 ( .A(n9935), .Z(n9936) );
  NAND U14220 ( .A(n10004), .B(n10005), .Z(n9935) );
  OR U14221 ( .A(n10006), .B(n10007), .Z(n10005) );
  OR U14222 ( .A(n10008), .B(n10009), .Z(n10004) );
  NAND U14223 ( .A(n10010), .B(n10011), .Z(n9933) );
  OR U14224 ( .A(n10012), .B(n10013), .Z(n10011) );
  OR U14225 ( .A(n10014), .B(n10015), .Z(n10010) );
  NOR U14226 ( .A(n10016), .B(n10017), .Z(n9934) );
  ANDN U14227 ( .B(n10018), .A(n10019), .Z(n9928) );
  IV U14228 ( .A(n10020), .Z(n10018) );
  XNOR U14229 ( .A(n9921), .B(n10021), .Z(n9927) );
  XNOR U14230 ( .A(n9920), .B(n9922), .Z(n10021) );
  NAND U14231 ( .A(n10022), .B(n10023), .Z(n9922) );
  OR U14232 ( .A(n10024), .B(n10025), .Z(n10023) );
  OR U14233 ( .A(n10026), .B(n10027), .Z(n10022) );
  NAND U14234 ( .A(n10028), .B(n10029), .Z(n9920) );
  OR U14235 ( .A(n10030), .B(n10031), .Z(n10029) );
  OR U14236 ( .A(n10032), .B(n10033), .Z(n10028) );
  ANDN U14237 ( .B(n10034), .A(n10035), .Z(n9921) );
  IV U14238 ( .A(n10036), .Z(n10034) );
  XNOR U14239 ( .A(n10001), .B(n10000), .Z(N29333) );
  XOR U14240 ( .A(n10020), .B(n10019), .Z(n10000) );
  XNOR U14241 ( .A(n10035), .B(n10036), .Z(n10019) );
  XNOR U14242 ( .A(n10030), .B(n10031), .Z(n10036) );
  XNOR U14243 ( .A(n10032), .B(n10033), .Z(n10031) );
  XNOR U14244 ( .A(y[2812]), .B(x[2812]), .Z(n10033) );
  XNOR U14245 ( .A(y[2813]), .B(x[2813]), .Z(n10032) );
  XNOR U14246 ( .A(y[2811]), .B(x[2811]), .Z(n10030) );
  XNOR U14247 ( .A(n10024), .B(n10025), .Z(n10035) );
  XNOR U14248 ( .A(y[2808]), .B(x[2808]), .Z(n10025) );
  XNOR U14249 ( .A(n10026), .B(n10027), .Z(n10024) );
  XNOR U14250 ( .A(y[2809]), .B(x[2809]), .Z(n10027) );
  XNOR U14251 ( .A(y[2810]), .B(x[2810]), .Z(n10026) );
  XNOR U14252 ( .A(n10017), .B(n10016), .Z(n10020) );
  XNOR U14253 ( .A(n10012), .B(n10013), .Z(n10016) );
  XNOR U14254 ( .A(y[2805]), .B(x[2805]), .Z(n10013) );
  XNOR U14255 ( .A(n10014), .B(n10015), .Z(n10012) );
  XNOR U14256 ( .A(y[2806]), .B(x[2806]), .Z(n10015) );
  XNOR U14257 ( .A(y[2807]), .B(x[2807]), .Z(n10014) );
  XNOR U14258 ( .A(n10006), .B(n10007), .Z(n10017) );
  XNOR U14259 ( .A(y[2802]), .B(x[2802]), .Z(n10007) );
  XNOR U14260 ( .A(n10008), .B(n10009), .Z(n10006) );
  XNOR U14261 ( .A(y[2803]), .B(x[2803]), .Z(n10009) );
  XNOR U14262 ( .A(y[2804]), .B(x[2804]), .Z(n10008) );
  XOR U14263 ( .A(n9982), .B(n9983), .Z(n10001) );
  XNOR U14264 ( .A(n9998), .B(n9999), .Z(n9983) );
  XNOR U14265 ( .A(n9993), .B(n9994), .Z(n9999) );
  XNOR U14266 ( .A(n9995), .B(n9996), .Z(n9994) );
  XNOR U14267 ( .A(y[2800]), .B(x[2800]), .Z(n9996) );
  XNOR U14268 ( .A(y[2801]), .B(x[2801]), .Z(n9995) );
  XNOR U14269 ( .A(y[2799]), .B(x[2799]), .Z(n9993) );
  XNOR U14270 ( .A(n9987), .B(n9988), .Z(n9998) );
  XNOR U14271 ( .A(y[2796]), .B(x[2796]), .Z(n9988) );
  XNOR U14272 ( .A(n9989), .B(n9990), .Z(n9987) );
  XNOR U14273 ( .A(y[2797]), .B(x[2797]), .Z(n9990) );
  XNOR U14274 ( .A(y[2798]), .B(x[2798]), .Z(n9989) );
  XOR U14275 ( .A(n9981), .B(n9980), .Z(n9982) );
  XNOR U14276 ( .A(n9976), .B(n9977), .Z(n9980) );
  XNOR U14277 ( .A(y[2793]), .B(x[2793]), .Z(n9977) );
  XNOR U14278 ( .A(n9978), .B(n9979), .Z(n9976) );
  XNOR U14279 ( .A(y[2794]), .B(x[2794]), .Z(n9979) );
  XNOR U14280 ( .A(y[2795]), .B(x[2795]), .Z(n9978) );
  XNOR U14281 ( .A(n9970), .B(n9971), .Z(n9981) );
  XNOR U14282 ( .A(y[2790]), .B(x[2790]), .Z(n9971) );
  XNOR U14283 ( .A(n9972), .B(n9973), .Z(n9970) );
  XNOR U14284 ( .A(y[2791]), .B(x[2791]), .Z(n9973) );
  XNOR U14285 ( .A(y[2792]), .B(x[2792]), .Z(n9972) );
  NAND U14286 ( .A(n10037), .B(n10038), .Z(N29325) );
  NANDN U14287 ( .A(n10039), .B(n10040), .Z(n10038) );
  OR U14288 ( .A(n10041), .B(n10042), .Z(n10040) );
  NAND U14289 ( .A(n10041), .B(n10042), .Z(n10037) );
  XOR U14290 ( .A(n10041), .B(n10043), .Z(N29324) );
  XNOR U14291 ( .A(n10039), .B(n10042), .Z(n10043) );
  AND U14292 ( .A(n10044), .B(n10045), .Z(n10042) );
  NANDN U14293 ( .A(n10046), .B(n10047), .Z(n10045) );
  NANDN U14294 ( .A(n10048), .B(n10049), .Z(n10047) );
  NANDN U14295 ( .A(n10049), .B(n10048), .Z(n10044) );
  NAND U14296 ( .A(n10050), .B(n10051), .Z(n10039) );
  NANDN U14297 ( .A(n10052), .B(n10053), .Z(n10051) );
  OR U14298 ( .A(n10054), .B(n10055), .Z(n10053) );
  NAND U14299 ( .A(n10055), .B(n10054), .Z(n10050) );
  AND U14300 ( .A(n10056), .B(n10057), .Z(n10041) );
  NANDN U14301 ( .A(n10058), .B(n10059), .Z(n10057) );
  NANDN U14302 ( .A(n10060), .B(n10061), .Z(n10059) );
  NANDN U14303 ( .A(n10061), .B(n10060), .Z(n10056) );
  XOR U14304 ( .A(n10055), .B(n10062), .Z(N29323) );
  XOR U14305 ( .A(n10052), .B(n10054), .Z(n10062) );
  XNOR U14306 ( .A(n10048), .B(n10063), .Z(n10054) );
  XNOR U14307 ( .A(n10046), .B(n10049), .Z(n10063) );
  NAND U14308 ( .A(n10064), .B(n10065), .Z(n10049) );
  NAND U14309 ( .A(n10066), .B(n10067), .Z(n10065) );
  OR U14310 ( .A(n10068), .B(n10069), .Z(n10066) );
  NANDN U14311 ( .A(n10070), .B(n10068), .Z(n10064) );
  IV U14312 ( .A(n10069), .Z(n10070) );
  NAND U14313 ( .A(n10071), .B(n10072), .Z(n10046) );
  NAND U14314 ( .A(n10073), .B(n10074), .Z(n10072) );
  NANDN U14315 ( .A(n10075), .B(n10076), .Z(n10073) );
  NANDN U14316 ( .A(n10076), .B(n10075), .Z(n10071) );
  AND U14317 ( .A(n10077), .B(n10078), .Z(n10048) );
  NAND U14318 ( .A(n10079), .B(n10080), .Z(n10078) );
  OR U14319 ( .A(n10081), .B(n10082), .Z(n10079) );
  NANDN U14320 ( .A(n10083), .B(n10081), .Z(n10077) );
  NAND U14321 ( .A(n10084), .B(n10085), .Z(n10052) );
  NANDN U14322 ( .A(n10086), .B(n10087), .Z(n10085) );
  OR U14323 ( .A(n10088), .B(n10089), .Z(n10087) );
  NANDN U14324 ( .A(n10090), .B(n10088), .Z(n10084) );
  IV U14325 ( .A(n10089), .Z(n10090) );
  XNOR U14326 ( .A(n10060), .B(n10091), .Z(n10055) );
  XNOR U14327 ( .A(n10058), .B(n10061), .Z(n10091) );
  NAND U14328 ( .A(n10092), .B(n10093), .Z(n10061) );
  NAND U14329 ( .A(n10094), .B(n10095), .Z(n10093) );
  OR U14330 ( .A(n10096), .B(n10097), .Z(n10094) );
  NANDN U14331 ( .A(n10098), .B(n10096), .Z(n10092) );
  IV U14332 ( .A(n10097), .Z(n10098) );
  NAND U14333 ( .A(n10099), .B(n10100), .Z(n10058) );
  NAND U14334 ( .A(n10101), .B(n10102), .Z(n10100) );
  NANDN U14335 ( .A(n10103), .B(n10104), .Z(n10101) );
  NANDN U14336 ( .A(n10104), .B(n10103), .Z(n10099) );
  AND U14337 ( .A(n10105), .B(n10106), .Z(n10060) );
  NAND U14338 ( .A(n10107), .B(n10108), .Z(n10106) );
  OR U14339 ( .A(n10109), .B(n10110), .Z(n10107) );
  NANDN U14340 ( .A(n10111), .B(n10109), .Z(n10105) );
  XNOR U14341 ( .A(n10086), .B(n10112), .Z(N29322) );
  XOR U14342 ( .A(n10088), .B(n10089), .Z(n10112) );
  XNOR U14343 ( .A(n10102), .B(n10113), .Z(n10089) );
  XOR U14344 ( .A(n10103), .B(n10104), .Z(n10113) );
  XOR U14345 ( .A(n10109), .B(n10114), .Z(n10104) );
  XOR U14346 ( .A(n10108), .B(n10111), .Z(n10114) );
  IV U14347 ( .A(n10110), .Z(n10111) );
  NAND U14348 ( .A(n10115), .B(n10116), .Z(n10110) );
  OR U14349 ( .A(n10117), .B(n10118), .Z(n10116) );
  OR U14350 ( .A(n10119), .B(n10120), .Z(n10115) );
  NAND U14351 ( .A(n10121), .B(n10122), .Z(n10108) );
  OR U14352 ( .A(n10123), .B(n10124), .Z(n10122) );
  OR U14353 ( .A(n10125), .B(n10126), .Z(n10121) );
  NOR U14354 ( .A(n10127), .B(n10128), .Z(n10109) );
  ANDN U14355 ( .B(n10129), .A(n10130), .Z(n10103) );
  XNOR U14356 ( .A(n10096), .B(n10131), .Z(n10102) );
  XNOR U14357 ( .A(n10095), .B(n10097), .Z(n10131) );
  NAND U14358 ( .A(n10132), .B(n10133), .Z(n10097) );
  OR U14359 ( .A(n10134), .B(n10135), .Z(n10133) );
  OR U14360 ( .A(n10136), .B(n10137), .Z(n10132) );
  NAND U14361 ( .A(n10138), .B(n10139), .Z(n10095) );
  OR U14362 ( .A(n10140), .B(n10141), .Z(n10139) );
  OR U14363 ( .A(n10142), .B(n10143), .Z(n10138) );
  ANDN U14364 ( .B(n10144), .A(n10145), .Z(n10096) );
  IV U14365 ( .A(n10146), .Z(n10144) );
  ANDN U14366 ( .B(n10147), .A(n10148), .Z(n10088) );
  XOR U14367 ( .A(n10074), .B(n10149), .Z(n10086) );
  XOR U14368 ( .A(n10075), .B(n10076), .Z(n10149) );
  XOR U14369 ( .A(n10081), .B(n10150), .Z(n10076) );
  XOR U14370 ( .A(n10080), .B(n10083), .Z(n10150) );
  IV U14371 ( .A(n10082), .Z(n10083) );
  NAND U14372 ( .A(n10151), .B(n10152), .Z(n10082) );
  OR U14373 ( .A(n10153), .B(n10154), .Z(n10152) );
  OR U14374 ( .A(n10155), .B(n10156), .Z(n10151) );
  NAND U14375 ( .A(n10157), .B(n10158), .Z(n10080) );
  OR U14376 ( .A(n10159), .B(n10160), .Z(n10158) );
  OR U14377 ( .A(n10161), .B(n10162), .Z(n10157) );
  NOR U14378 ( .A(n10163), .B(n10164), .Z(n10081) );
  ANDN U14379 ( .B(n10165), .A(n10166), .Z(n10075) );
  IV U14380 ( .A(n10167), .Z(n10165) );
  XNOR U14381 ( .A(n10068), .B(n10168), .Z(n10074) );
  XNOR U14382 ( .A(n10067), .B(n10069), .Z(n10168) );
  NAND U14383 ( .A(n10169), .B(n10170), .Z(n10069) );
  OR U14384 ( .A(n10171), .B(n10172), .Z(n10170) );
  OR U14385 ( .A(n10173), .B(n10174), .Z(n10169) );
  NAND U14386 ( .A(n10175), .B(n10176), .Z(n10067) );
  OR U14387 ( .A(n10177), .B(n10178), .Z(n10176) );
  OR U14388 ( .A(n10179), .B(n10180), .Z(n10175) );
  ANDN U14389 ( .B(n10181), .A(n10182), .Z(n10068) );
  IV U14390 ( .A(n10183), .Z(n10181) );
  XNOR U14391 ( .A(n10148), .B(n10147), .Z(N29321) );
  XOR U14392 ( .A(n10167), .B(n10166), .Z(n10147) );
  XNOR U14393 ( .A(n10182), .B(n10183), .Z(n10166) );
  XNOR U14394 ( .A(n10177), .B(n10178), .Z(n10183) );
  XNOR U14395 ( .A(n10179), .B(n10180), .Z(n10178) );
  XNOR U14396 ( .A(y[2788]), .B(x[2788]), .Z(n10180) );
  XNOR U14397 ( .A(y[2789]), .B(x[2789]), .Z(n10179) );
  XNOR U14398 ( .A(y[2787]), .B(x[2787]), .Z(n10177) );
  XNOR U14399 ( .A(n10171), .B(n10172), .Z(n10182) );
  XNOR U14400 ( .A(y[2784]), .B(x[2784]), .Z(n10172) );
  XNOR U14401 ( .A(n10173), .B(n10174), .Z(n10171) );
  XNOR U14402 ( .A(y[2785]), .B(x[2785]), .Z(n10174) );
  XNOR U14403 ( .A(y[2786]), .B(x[2786]), .Z(n10173) );
  XNOR U14404 ( .A(n10164), .B(n10163), .Z(n10167) );
  XNOR U14405 ( .A(n10159), .B(n10160), .Z(n10163) );
  XNOR U14406 ( .A(y[2781]), .B(x[2781]), .Z(n10160) );
  XNOR U14407 ( .A(n10161), .B(n10162), .Z(n10159) );
  XNOR U14408 ( .A(y[2782]), .B(x[2782]), .Z(n10162) );
  XNOR U14409 ( .A(y[2783]), .B(x[2783]), .Z(n10161) );
  XNOR U14410 ( .A(n10153), .B(n10154), .Z(n10164) );
  XNOR U14411 ( .A(y[2778]), .B(x[2778]), .Z(n10154) );
  XNOR U14412 ( .A(n10155), .B(n10156), .Z(n10153) );
  XNOR U14413 ( .A(y[2779]), .B(x[2779]), .Z(n10156) );
  XNOR U14414 ( .A(y[2780]), .B(x[2780]), .Z(n10155) );
  XOR U14415 ( .A(n10129), .B(n10130), .Z(n10148) );
  XNOR U14416 ( .A(n10145), .B(n10146), .Z(n10130) );
  XNOR U14417 ( .A(n10140), .B(n10141), .Z(n10146) );
  XNOR U14418 ( .A(n10142), .B(n10143), .Z(n10141) );
  XNOR U14419 ( .A(y[2776]), .B(x[2776]), .Z(n10143) );
  XNOR U14420 ( .A(y[2777]), .B(x[2777]), .Z(n10142) );
  XNOR U14421 ( .A(y[2775]), .B(x[2775]), .Z(n10140) );
  XNOR U14422 ( .A(n10134), .B(n10135), .Z(n10145) );
  XNOR U14423 ( .A(y[2772]), .B(x[2772]), .Z(n10135) );
  XNOR U14424 ( .A(n10136), .B(n10137), .Z(n10134) );
  XNOR U14425 ( .A(y[2773]), .B(x[2773]), .Z(n10137) );
  XNOR U14426 ( .A(y[2774]), .B(x[2774]), .Z(n10136) );
  XOR U14427 ( .A(n10128), .B(n10127), .Z(n10129) );
  XNOR U14428 ( .A(n10123), .B(n10124), .Z(n10127) );
  XNOR U14429 ( .A(y[2769]), .B(x[2769]), .Z(n10124) );
  XNOR U14430 ( .A(n10125), .B(n10126), .Z(n10123) );
  XNOR U14431 ( .A(y[2770]), .B(x[2770]), .Z(n10126) );
  XNOR U14432 ( .A(y[2771]), .B(x[2771]), .Z(n10125) );
  XNOR U14433 ( .A(n10117), .B(n10118), .Z(n10128) );
  XNOR U14434 ( .A(y[2766]), .B(x[2766]), .Z(n10118) );
  XNOR U14435 ( .A(n10119), .B(n10120), .Z(n10117) );
  XNOR U14436 ( .A(y[2767]), .B(x[2767]), .Z(n10120) );
  XNOR U14437 ( .A(y[2768]), .B(x[2768]), .Z(n10119) );
  NAND U14438 ( .A(n10184), .B(n10185), .Z(N29313) );
  NANDN U14439 ( .A(n10186), .B(n10187), .Z(n10185) );
  OR U14440 ( .A(n10188), .B(n10189), .Z(n10187) );
  NAND U14441 ( .A(n10188), .B(n10189), .Z(n10184) );
  XOR U14442 ( .A(n10188), .B(n10190), .Z(N29312) );
  XNOR U14443 ( .A(n10186), .B(n10189), .Z(n10190) );
  AND U14444 ( .A(n10191), .B(n10192), .Z(n10189) );
  NANDN U14445 ( .A(n10193), .B(n10194), .Z(n10192) );
  NANDN U14446 ( .A(n10195), .B(n10196), .Z(n10194) );
  NANDN U14447 ( .A(n10196), .B(n10195), .Z(n10191) );
  NAND U14448 ( .A(n10197), .B(n10198), .Z(n10186) );
  NANDN U14449 ( .A(n10199), .B(n10200), .Z(n10198) );
  OR U14450 ( .A(n10201), .B(n10202), .Z(n10200) );
  NAND U14451 ( .A(n10202), .B(n10201), .Z(n10197) );
  AND U14452 ( .A(n10203), .B(n10204), .Z(n10188) );
  NANDN U14453 ( .A(n10205), .B(n10206), .Z(n10204) );
  NANDN U14454 ( .A(n10207), .B(n10208), .Z(n10206) );
  NANDN U14455 ( .A(n10208), .B(n10207), .Z(n10203) );
  XOR U14456 ( .A(n10202), .B(n10209), .Z(N29311) );
  XOR U14457 ( .A(n10199), .B(n10201), .Z(n10209) );
  XNOR U14458 ( .A(n10195), .B(n10210), .Z(n10201) );
  XNOR U14459 ( .A(n10193), .B(n10196), .Z(n10210) );
  NAND U14460 ( .A(n10211), .B(n10212), .Z(n10196) );
  NAND U14461 ( .A(n10213), .B(n10214), .Z(n10212) );
  OR U14462 ( .A(n10215), .B(n10216), .Z(n10213) );
  NANDN U14463 ( .A(n10217), .B(n10215), .Z(n10211) );
  IV U14464 ( .A(n10216), .Z(n10217) );
  NAND U14465 ( .A(n10218), .B(n10219), .Z(n10193) );
  NAND U14466 ( .A(n10220), .B(n10221), .Z(n10219) );
  NANDN U14467 ( .A(n10222), .B(n10223), .Z(n10220) );
  NANDN U14468 ( .A(n10223), .B(n10222), .Z(n10218) );
  AND U14469 ( .A(n10224), .B(n10225), .Z(n10195) );
  NAND U14470 ( .A(n10226), .B(n10227), .Z(n10225) );
  OR U14471 ( .A(n10228), .B(n10229), .Z(n10226) );
  NANDN U14472 ( .A(n10230), .B(n10228), .Z(n10224) );
  NAND U14473 ( .A(n10231), .B(n10232), .Z(n10199) );
  NANDN U14474 ( .A(n10233), .B(n10234), .Z(n10232) );
  OR U14475 ( .A(n10235), .B(n10236), .Z(n10234) );
  NANDN U14476 ( .A(n10237), .B(n10235), .Z(n10231) );
  IV U14477 ( .A(n10236), .Z(n10237) );
  XNOR U14478 ( .A(n10207), .B(n10238), .Z(n10202) );
  XNOR U14479 ( .A(n10205), .B(n10208), .Z(n10238) );
  NAND U14480 ( .A(n10239), .B(n10240), .Z(n10208) );
  NAND U14481 ( .A(n10241), .B(n10242), .Z(n10240) );
  OR U14482 ( .A(n10243), .B(n10244), .Z(n10241) );
  NANDN U14483 ( .A(n10245), .B(n10243), .Z(n10239) );
  IV U14484 ( .A(n10244), .Z(n10245) );
  NAND U14485 ( .A(n10246), .B(n10247), .Z(n10205) );
  NAND U14486 ( .A(n10248), .B(n10249), .Z(n10247) );
  NANDN U14487 ( .A(n10250), .B(n10251), .Z(n10248) );
  NANDN U14488 ( .A(n10251), .B(n10250), .Z(n10246) );
  AND U14489 ( .A(n10252), .B(n10253), .Z(n10207) );
  NAND U14490 ( .A(n10254), .B(n10255), .Z(n10253) );
  OR U14491 ( .A(n10256), .B(n10257), .Z(n10254) );
  NANDN U14492 ( .A(n10258), .B(n10256), .Z(n10252) );
  XNOR U14493 ( .A(n10233), .B(n10259), .Z(N29310) );
  XOR U14494 ( .A(n10235), .B(n10236), .Z(n10259) );
  XNOR U14495 ( .A(n10249), .B(n10260), .Z(n10236) );
  XOR U14496 ( .A(n10250), .B(n10251), .Z(n10260) );
  XOR U14497 ( .A(n10256), .B(n10261), .Z(n10251) );
  XOR U14498 ( .A(n10255), .B(n10258), .Z(n10261) );
  IV U14499 ( .A(n10257), .Z(n10258) );
  NAND U14500 ( .A(n10262), .B(n10263), .Z(n10257) );
  OR U14501 ( .A(n10264), .B(n10265), .Z(n10263) );
  OR U14502 ( .A(n10266), .B(n10267), .Z(n10262) );
  NAND U14503 ( .A(n10268), .B(n10269), .Z(n10255) );
  OR U14504 ( .A(n10270), .B(n10271), .Z(n10269) );
  OR U14505 ( .A(n10272), .B(n10273), .Z(n10268) );
  NOR U14506 ( .A(n10274), .B(n10275), .Z(n10256) );
  ANDN U14507 ( .B(n10276), .A(n10277), .Z(n10250) );
  XNOR U14508 ( .A(n10243), .B(n10278), .Z(n10249) );
  XNOR U14509 ( .A(n10242), .B(n10244), .Z(n10278) );
  NAND U14510 ( .A(n10279), .B(n10280), .Z(n10244) );
  OR U14511 ( .A(n10281), .B(n10282), .Z(n10280) );
  OR U14512 ( .A(n10283), .B(n10284), .Z(n10279) );
  NAND U14513 ( .A(n10285), .B(n10286), .Z(n10242) );
  OR U14514 ( .A(n10287), .B(n10288), .Z(n10286) );
  OR U14515 ( .A(n10289), .B(n10290), .Z(n10285) );
  ANDN U14516 ( .B(n10291), .A(n10292), .Z(n10243) );
  IV U14517 ( .A(n10293), .Z(n10291) );
  ANDN U14518 ( .B(n10294), .A(n10295), .Z(n10235) );
  XOR U14519 ( .A(n10221), .B(n10296), .Z(n10233) );
  XOR U14520 ( .A(n10222), .B(n10223), .Z(n10296) );
  XOR U14521 ( .A(n10228), .B(n10297), .Z(n10223) );
  XOR U14522 ( .A(n10227), .B(n10230), .Z(n10297) );
  IV U14523 ( .A(n10229), .Z(n10230) );
  NAND U14524 ( .A(n10298), .B(n10299), .Z(n10229) );
  OR U14525 ( .A(n10300), .B(n10301), .Z(n10299) );
  OR U14526 ( .A(n10302), .B(n10303), .Z(n10298) );
  NAND U14527 ( .A(n10304), .B(n10305), .Z(n10227) );
  OR U14528 ( .A(n10306), .B(n10307), .Z(n10305) );
  OR U14529 ( .A(n10308), .B(n10309), .Z(n10304) );
  NOR U14530 ( .A(n10310), .B(n10311), .Z(n10228) );
  ANDN U14531 ( .B(n10312), .A(n10313), .Z(n10222) );
  IV U14532 ( .A(n10314), .Z(n10312) );
  XNOR U14533 ( .A(n10215), .B(n10315), .Z(n10221) );
  XNOR U14534 ( .A(n10214), .B(n10216), .Z(n10315) );
  NAND U14535 ( .A(n10316), .B(n10317), .Z(n10216) );
  OR U14536 ( .A(n10318), .B(n10319), .Z(n10317) );
  OR U14537 ( .A(n10320), .B(n10321), .Z(n10316) );
  NAND U14538 ( .A(n10322), .B(n10323), .Z(n10214) );
  OR U14539 ( .A(n10324), .B(n10325), .Z(n10323) );
  OR U14540 ( .A(n10326), .B(n10327), .Z(n10322) );
  ANDN U14541 ( .B(n10328), .A(n10329), .Z(n10215) );
  IV U14542 ( .A(n10330), .Z(n10328) );
  XNOR U14543 ( .A(n10295), .B(n10294), .Z(N29309) );
  XOR U14544 ( .A(n10314), .B(n10313), .Z(n10294) );
  XNOR U14545 ( .A(n10329), .B(n10330), .Z(n10313) );
  XNOR U14546 ( .A(n10324), .B(n10325), .Z(n10330) );
  XNOR U14547 ( .A(n10326), .B(n10327), .Z(n10325) );
  XNOR U14548 ( .A(y[2764]), .B(x[2764]), .Z(n10327) );
  XNOR U14549 ( .A(y[2765]), .B(x[2765]), .Z(n10326) );
  XNOR U14550 ( .A(y[2763]), .B(x[2763]), .Z(n10324) );
  XNOR U14551 ( .A(n10318), .B(n10319), .Z(n10329) );
  XNOR U14552 ( .A(y[2760]), .B(x[2760]), .Z(n10319) );
  XNOR U14553 ( .A(n10320), .B(n10321), .Z(n10318) );
  XNOR U14554 ( .A(y[2761]), .B(x[2761]), .Z(n10321) );
  XNOR U14555 ( .A(y[2762]), .B(x[2762]), .Z(n10320) );
  XNOR U14556 ( .A(n10311), .B(n10310), .Z(n10314) );
  XNOR U14557 ( .A(n10306), .B(n10307), .Z(n10310) );
  XNOR U14558 ( .A(y[2757]), .B(x[2757]), .Z(n10307) );
  XNOR U14559 ( .A(n10308), .B(n10309), .Z(n10306) );
  XNOR U14560 ( .A(y[2758]), .B(x[2758]), .Z(n10309) );
  XNOR U14561 ( .A(y[2759]), .B(x[2759]), .Z(n10308) );
  XNOR U14562 ( .A(n10300), .B(n10301), .Z(n10311) );
  XNOR U14563 ( .A(y[2754]), .B(x[2754]), .Z(n10301) );
  XNOR U14564 ( .A(n10302), .B(n10303), .Z(n10300) );
  XNOR U14565 ( .A(y[2755]), .B(x[2755]), .Z(n10303) );
  XNOR U14566 ( .A(y[2756]), .B(x[2756]), .Z(n10302) );
  XOR U14567 ( .A(n10276), .B(n10277), .Z(n10295) );
  XNOR U14568 ( .A(n10292), .B(n10293), .Z(n10277) );
  XNOR U14569 ( .A(n10287), .B(n10288), .Z(n10293) );
  XNOR U14570 ( .A(n10289), .B(n10290), .Z(n10288) );
  XNOR U14571 ( .A(y[2752]), .B(x[2752]), .Z(n10290) );
  XNOR U14572 ( .A(y[2753]), .B(x[2753]), .Z(n10289) );
  XNOR U14573 ( .A(y[2751]), .B(x[2751]), .Z(n10287) );
  XNOR U14574 ( .A(n10281), .B(n10282), .Z(n10292) );
  XNOR U14575 ( .A(y[2748]), .B(x[2748]), .Z(n10282) );
  XNOR U14576 ( .A(n10283), .B(n10284), .Z(n10281) );
  XNOR U14577 ( .A(y[2749]), .B(x[2749]), .Z(n10284) );
  XNOR U14578 ( .A(y[2750]), .B(x[2750]), .Z(n10283) );
  XOR U14579 ( .A(n10275), .B(n10274), .Z(n10276) );
  XNOR U14580 ( .A(n10270), .B(n10271), .Z(n10274) );
  XNOR U14581 ( .A(y[2745]), .B(x[2745]), .Z(n10271) );
  XNOR U14582 ( .A(n10272), .B(n10273), .Z(n10270) );
  XNOR U14583 ( .A(y[2746]), .B(x[2746]), .Z(n10273) );
  XNOR U14584 ( .A(y[2747]), .B(x[2747]), .Z(n10272) );
  XNOR U14585 ( .A(n10264), .B(n10265), .Z(n10275) );
  XNOR U14586 ( .A(y[2742]), .B(x[2742]), .Z(n10265) );
  XNOR U14587 ( .A(n10266), .B(n10267), .Z(n10264) );
  XNOR U14588 ( .A(y[2743]), .B(x[2743]), .Z(n10267) );
  XNOR U14589 ( .A(y[2744]), .B(x[2744]), .Z(n10266) );
  NAND U14590 ( .A(n10331), .B(n10332), .Z(N29301) );
  NANDN U14591 ( .A(n10333), .B(n10334), .Z(n10332) );
  OR U14592 ( .A(n10335), .B(n10336), .Z(n10334) );
  NAND U14593 ( .A(n10335), .B(n10336), .Z(n10331) );
  XOR U14594 ( .A(n10335), .B(n10337), .Z(N29300) );
  XNOR U14595 ( .A(n10333), .B(n10336), .Z(n10337) );
  AND U14596 ( .A(n10338), .B(n10339), .Z(n10336) );
  NANDN U14597 ( .A(n10340), .B(n10341), .Z(n10339) );
  NANDN U14598 ( .A(n10342), .B(n10343), .Z(n10341) );
  NANDN U14599 ( .A(n10343), .B(n10342), .Z(n10338) );
  NAND U14600 ( .A(n10344), .B(n10345), .Z(n10333) );
  NANDN U14601 ( .A(n10346), .B(n10347), .Z(n10345) );
  OR U14602 ( .A(n10348), .B(n10349), .Z(n10347) );
  NAND U14603 ( .A(n10349), .B(n10348), .Z(n10344) );
  AND U14604 ( .A(n10350), .B(n10351), .Z(n10335) );
  NANDN U14605 ( .A(n10352), .B(n10353), .Z(n10351) );
  NANDN U14606 ( .A(n10354), .B(n10355), .Z(n10353) );
  NANDN U14607 ( .A(n10355), .B(n10354), .Z(n10350) );
  XOR U14608 ( .A(n10349), .B(n10356), .Z(N29299) );
  XOR U14609 ( .A(n10346), .B(n10348), .Z(n10356) );
  XNOR U14610 ( .A(n10342), .B(n10357), .Z(n10348) );
  XNOR U14611 ( .A(n10340), .B(n10343), .Z(n10357) );
  NAND U14612 ( .A(n10358), .B(n10359), .Z(n10343) );
  NAND U14613 ( .A(n10360), .B(n10361), .Z(n10359) );
  OR U14614 ( .A(n10362), .B(n10363), .Z(n10360) );
  NANDN U14615 ( .A(n10364), .B(n10362), .Z(n10358) );
  IV U14616 ( .A(n10363), .Z(n10364) );
  NAND U14617 ( .A(n10365), .B(n10366), .Z(n10340) );
  NAND U14618 ( .A(n10367), .B(n10368), .Z(n10366) );
  NANDN U14619 ( .A(n10369), .B(n10370), .Z(n10367) );
  NANDN U14620 ( .A(n10370), .B(n10369), .Z(n10365) );
  AND U14621 ( .A(n10371), .B(n10372), .Z(n10342) );
  NAND U14622 ( .A(n10373), .B(n10374), .Z(n10372) );
  OR U14623 ( .A(n10375), .B(n10376), .Z(n10373) );
  NANDN U14624 ( .A(n10377), .B(n10375), .Z(n10371) );
  NAND U14625 ( .A(n10378), .B(n10379), .Z(n10346) );
  NANDN U14626 ( .A(n10380), .B(n10381), .Z(n10379) );
  OR U14627 ( .A(n10382), .B(n10383), .Z(n10381) );
  NANDN U14628 ( .A(n10384), .B(n10382), .Z(n10378) );
  IV U14629 ( .A(n10383), .Z(n10384) );
  XNOR U14630 ( .A(n10354), .B(n10385), .Z(n10349) );
  XNOR U14631 ( .A(n10352), .B(n10355), .Z(n10385) );
  NAND U14632 ( .A(n10386), .B(n10387), .Z(n10355) );
  NAND U14633 ( .A(n10388), .B(n10389), .Z(n10387) );
  OR U14634 ( .A(n10390), .B(n10391), .Z(n10388) );
  NANDN U14635 ( .A(n10392), .B(n10390), .Z(n10386) );
  IV U14636 ( .A(n10391), .Z(n10392) );
  NAND U14637 ( .A(n10393), .B(n10394), .Z(n10352) );
  NAND U14638 ( .A(n10395), .B(n10396), .Z(n10394) );
  NANDN U14639 ( .A(n10397), .B(n10398), .Z(n10395) );
  NANDN U14640 ( .A(n10398), .B(n10397), .Z(n10393) );
  AND U14641 ( .A(n10399), .B(n10400), .Z(n10354) );
  NAND U14642 ( .A(n10401), .B(n10402), .Z(n10400) );
  OR U14643 ( .A(n10403), .B(n10404), .Z(n10401) );
  NANDN U14644 ( .A(n10405), .B(n10403), .Z(n10399) );
  XNOR U14645 ( .A(n10380), .B(n10406), .Z(N29298) );
  XOR U14646 ( .A(n10382), .B(n10383), .Z(n10406) );
  XNOR U14647 ( .A(n10396), .B(n10407), .Z(n10383) );
  XOR U14648 ( .A(n10397), .B(n10398), .Z(n10407) );
  XOR U14649 ( .A(n10403), .B(n10408), .Z(n10398) );
  XOR U14650 ( .A(n10402), .B(n10405), .Z(n10408) );
  IV U14651 ( .A(n10404), .Z(n10405) );
  NAND U14652 ( .A(n10409), .B(n10410), .Z(n10404) );
  OR U14653 ( .A(n10411), .B(n10412), .Z(n10410) );
  OR U14654 ( .A(n10413), .B(n10414), .Z(n10409) );
  NAND U14655 ( .A(n10415), .B(n10416), .Z(n10402) );
  OR U14656 ( .A(n10417), .B(n10418), .Z(n10416) );
  OR U14657 ( .A(n10419), .B(n10420), .Z(n10415) );
  NOR U14658 ( .A(n10421), .B(n10422), .Z(n10403) );
  ANDN U14659 ( .B(n10423), .A(n10424), .Z(n10397) );
  XNOR U14660 ( .A(n10390), .B(n10425), .Z(n10396) );
  XNOR U14661 ( .A(n10389), .B(n10391), .Z(n10425) );
  NAND U14662 ( .A(n10426), .B(n10427), .Z(n10391) );
  OR U14663 ( .A(n10428), .B(n10429), .Z(n10427) );
  OR U14664 ( .A(n10430), .B(n10431), .Z(n10426) );
  NAND U14665 ( .A(n10432), .B(n10433), .Z(n10389) );
  OR U14666 ( .A(n10434), .B(n10435), .Z(n10433) );
  OR U14667 ( .A(n10436), .B(n10437), .Z(n10432) );
  ANDN U14668 ( .B(n10438), .A(n10439), .Z(n10390) );
  IV U14669 ( .A(n10440), .Z(n10438) );
  ANDN U14670 ( .B(n10441), .A(n10442), .Z(n10382) );
  XOR U14671 ( .A(n10368), .B(n10443), .Z(n10380) );
  XOR U14672 ( .A(n10369), .B(n10370), .Z(n10443) );
  XOR U14673 ( .A(n10375), .B(n10444), .Z(n10370) );
  XOR U14674 ( .A(n10374), .B(n10377), .Z(n10444) );
  IV U14675 ( .A(n10376), .Z(n10377) );
  NAND U14676 ( .A(n10445), .B(n10446), .Z(n10376) );
  OR U14677 ( .A(n10447), .B(n10448), .Z(n10446) );
  OR U14678 ( .A(n10449), .B(n10450), .Z(n10445) );
  NAND U14679 ( .A(n10451), .B(n10452), .Z(n10374) );
  OR U14680 ( .A(n10453), .B(n10454), .Z(n10452) );
  OR U14681 ( .A(n10455), .B(n10456), .Z(n10451) );
  NOR U14682 ( .A(n10457), .B(n10458), .Z(n10375) );
  ANDN U14683 ( .B(n10459), .A(n10460), .Z(n10369) );
  IV U14684 ( .A(n10461), .Z(n10459) );
  XNOR U14685 ( .A(n10362), .B(n10462), .Z(n10368) );
  XNOR U14686 ( .A(n10361), .B(n10363), .Z(n10462) );
  NAND U14687 ( .A(n10463), .B(n10464), .Z(n10363) );
  OR U14688 ( .A(n10465), .B(n10466), .Z(n10464) );
  OR U14689 ( .A(n10467), .B(n10468), .Z(n10463) );
  NAND U14690 ( .A(n10469), .B(n10470), .Z(n10361) );
  OR U14691 ( .A(n10471), .B(n10472), .Z(n10470) );
  OR U14692 ( .A(n10473), .B(n10474), .Z(n10469) );
  ANDN U14693 ( .B(n10475), .A(n10476), .Z(n10362) );
  IV U14694 ( .A(n10477), .Z(n10475) );
  XNOR U14695 ( .A(n10442), .B(n10441), .Z(N29297) );
  XOR U14696 ( .A(n10461), .B(n10460), .Z(n10441) );
  XNOR U14697 ( .A(n10476), .B(n10477), .Z(n10460) );
  XNOR U14698 ( .A(n10471), .B(n10472), .Z(n10477) );
  XNOR U14699 ( .A(n10473), .B(n10474), .Z(n10472) );
  XNOR U14700 ( .A(y[2740]), .B(x[2740]), .Z(n10474) );
  XNOR U14701 ( .A(y[2741]), .B(x[2741]), .Z(n10473) );
  XNOR U14702 ( .A(y[2739]), .B(x[2739]), .Z(n10471) );
  XNOR U14703 ( .A(n10465), .B(n10466), .Z(n10476) );
  XNOR U14704 ( .A(y[2736]), .B(x[2736]), .Z(n10466) );
  XNOR U14705 ( .A(n10467), .B(n10468), .Z(n10465) );
  XNOR U14706 ( .A(y[2737]), .B(x[2737]), .Z(n10468) );
  XNOR U14707 ( .A(y[2738]), .B(x[2738]), .Z(n10467) );
  XNOR U14708 ( .A(n10458), .B(n10457), .Z(n10461) );
  XNOR U14709 ( .A(n10453), .B(n10454), .Z(n10457) );
  XNOR U14710 ( .A(y[2733]), .B(x[2733]), .Z(n10454) );
  XNOR U14711 ( .A(n10455), .B(n10456), .Z(n10453) );
  XNOR U14712 ( .A(y[2734]), .B(x[2734]), .Z(n10456) );
  XNOR U14713 ( .A(y[2735]), .B(x[2735]), .Z(n10455) );
  XNOR U14714 ( .A(n10447), .B(n10448), .Z(n10458) );
  XNOR U14715 ( .A(y[2730]), .B(x[2730]), .Z(n10448) );
  XNOR U14716 ( .A(n10449), .B(n10450), .Z(n10447) );
  XNOR U14717 ( .A(y[2731]), .B(x[2731]), .Z(n10450) );
  XNOR U14718 ( .A(y[2732]), .B(x[2732]), .Z(n10449) );
  XOR U14719 ( .A(n10423), .B(n10424), .Z(n10442) );
  XNOR U14720 ( .A(n10439), .B(n10440), .Z(n10424) );
  XNOR U14721 ( .A(n10434), .B(n10435), .Z(n10440) );
  XNOR U14722 ( .A(n10436), .B(n10437), .Z(n10435) );
  XNOR U14723 ( .A(y[2728]), .B(x[2728]), .Z(n10437) );
  XNOR U14724 ( .A(y[2729]), .B(x[2729]), .Z(n10436) );
  XNOR U14725 ( .A(y[2727]), .B(x[2727]), .Z(n10434) );
  XNOR U14726 ( .A(n10428), .B(n10429), .Z(n10439) );
  XNOR U14727 ( .A(y[2724]), .B(x[2724]), .Z(n10429) );
  XNOR U14728 ( .A(n10430), .B(n10431), .Z(n10428) );
  XNOR U14729 ( .A(y[2725]), .B(x[2725]), .Z(n10431) );
  XNOR U14730 ( .A(y[2726]), .B(x[2726]), .Z(n10430) );
  XOR U14731 ( .A(n10422), .B(n10421), .Z(n10423) );
  XNOR U14732 ( .A(n10417), .B(n10418), .Z(n10421) );
  XNOR U14733 ( .A(y[2721]), .B(x[2721]), .Z(n10418) );
  XNOR U14734 ( .A(n10419), .B(n10420), .Z(n10417) );
  XNOR U14735 ( .A(y[2722]), .B(x[2722]), .Z(n10420) );
  XNOR U14736 ( .A(y[2723]), .B(x[2723]), .Z(n10419) );
  XNOR U14737 ( .A(n10411), .B(n10412), .Z(n10422) );
  XNOR U14738 ( .A(y[2718]), .B(x[2718]), .Z(n10412) );
  XNOR U14739 ( .A(n10413), .B(n10414), .Z(n10411) );
  XNOR U14740 ( .A(y[2719]), .B(x[2719]), .Z(n10414) );
  XNOR U14741 ( .A(y[2720]), .B(x[2720]), .Z(n10413) );
  NAND U14742 ( .A(n10478), .B(n10479), .Z(N29289) );
  NANDN U14743 ( .A(n10480), .B(n10481), .Z(n10479) );
  OR U14744 ( .A(n10482), .B(n10483), .Z(n10481) );
  NAND U14745 ( .A(n10482), .B(n10483), .Z(n10478) );
  XOR U14746 ( .A(n10482), .B(n10484), .Z(N29288) );
  XNOR U14747 ( .A(n10480), .B(n10483), .Z(n10484) );
  AND U14748 ( .A(n10485), .B(n10486), .Z(n10483) );
  NANDN U14749 ( .A(n10487), .B(n10488), .Z(n10486) );
  NANDN U14750 ( .A(n10489), .B(n10490), .Z(n10488) );
  NANDN U14751 ( .A(n10490), .B(n10489), .Z(n10485) );
  NAND U14752 ( .A(n10491), .B(n10492), .Z(n10480) );
  NANDN U14753 ( .A(n10493), .B(n10494), .Z(n10492) );
  OR U14754 ( .A(n10495), .B(n10496), .Z(n10494) );
  NAND U14755 ( .A(n10496), .B(n10495), .Z(n10491) );
  AND U14756 ( .A(n10497), .B(n10498), .Z(n10482) );
  NANDN U14757 ( .A(n10499), .B(n10500), .Z(n10498) );
  NANDN U14758 ( .A(n10501), .B(n10502), .Z(n10500) );
  NANDN U14759 ( .A(n10502), .B(n10501), .Z(n10497) );
  XOR U14760 ( .A(n10496), .B(n10503), .Z(N29287) );
  XOR U14761 ( .A(n10493), .B(n10495), .Z(n10503) );
  XNOR U14762 ( .A(n10489), .B(n10504), .Z(n10495) );
  XNOR U14763 ( .A(n10487), .B(n10490), .Z(n10504) );
  NAND U14764 ( .A(n10505), .B(n10506), .Z(n10490) );
  NAND U14765 ( .A(n10507), .B(n10508), .Z(n10506) );
  OR U14766 ( .A(n10509), .B(n10510), .Z(n10507) );
  NANDN U14767 ( .A(n10511), .B(n10509), .Z(n10505) );
  IV U14768 ( .A(n10510), .Z(n10511) );
  NAND U14769 ( .A(n10512), .B(n10513), .Z(n10487) );
  NAND U14770 ( .A(n10514), .B(n10515), .Z(n10513) );
  NANDN U14771 ( .A(n10516), .B(n10517), .Z(n10514) );
  NANDN U14772 ( .A(n10517), .B(n10516), .Z(n10512) );
  AND U14773 ( .A(n10518), .B(n10519), .Z(n10489) );
  NAND U14774 ( .A(n10520), .B(n10521), .Z(n10519) );
  OR U14775 ( .A(n10522), .B(n10523), .Z(n10520) );
  NANDN U14776 ( .A(n10524), .B(n10522), .Z(n10518) );
  NAND U14777 ( .A(n10525), .B(n10526), .Z(n10493) );
  NANDN U14778 ( .A(n10527), .B(n10528), .Z(n10526) );
  OR U14779 ( .A(n10529), .B(n10530), .Z(n10528) );
  NANDN U14780 ( .A(n10531), .B(n10529), .Z(n10525) );
  IV U14781 ( .A(n10530), .Z(n10531) );
  XNOR U14782 ( .A(n10501), .B(n10532), .Z(n10496) );
  XNOR U14783 ( .A(n10499), .B(n10502), .Z(n10532) );
  NAND U14784 ( .A(n10533), .B(n10534), .Z(n10502) );
  NAND U14785 ( .A(n10535), .B(n10536), .Z(n10534) );
  OR U14786 ( .A(n10537), .B(n10538), .Z(n10535) );
  NANDN U14787 ( .A(n10539), .B(n10537), .Z(n10533) );
  IV U14788 ( .A(n10538), .Z(n10539) );
  NAND U14789 ( .A(n10540), .B(n10541), .Z(n10499) );
  NAND U14790 ( .A(n10542), .B(n10543), .Z(n10541) );
  NANDN U14791 ( .A(n10544), .B(n10545), .Z(n10542) );
  NANDN U14792 ( .A(n10545), .B(n10544), .Z(n10540) );
  AND U14793 ( .A(n10546), .B(n10547), .Z(n10501) );
  NAND U14794 ( .A(n10548), .B(n10549), .Z(n10547) );
  OR U14795 ( .A(n10550), .B(n10551), .Z(n10548) );
  NANDN U14796 ( .A(n10552), .B(n10550), .Z(n10546) );
  XNOR U14797 ( .A(n10527), .B(n10553), .Z(N29286) );
  XOR U14798 ( .A(n10529), .B(n10530), .Z(n10553) );
  XNOR U14799 ( .A(n10543), .B(n10554), .Z(n10530) );
  XOR U14800 ( .A(n10544), .B(n10545), .Z(n10554) );
  XOR U14801 ( .A(n10550), .B(n10555), .Z(n10545) );
  XOR U14802 ( .A(n10549), .B(n10552), .Z(n10555) );
  IV U14803 ( .A(n10551), .Z(n10552) );
  NAND U14804 ( .A(n10556), .B(n10557), .Z(n10551) );
  OR U14805 ( .A(n10558), .B(n10559), .Z(n10557) );
  OR U14806 ( .A(n10560), .B(n10561), .Z(n10556) );
  NAND U14807 ( .A(n10562), .B(n10563), .Z(n10549) );
  OR U14808 ( .A(n10564), .B(n10565), .Z(n10563) );
  OR U14809 ( .A(n10566), .B(n10567), .Z(n10562) );
  NOR U14810 ( .A(n10568), .B(n10569), .Z(n10550) );
  ANDN U14811 ( .B(n10570), .A(n10571), .Z(n10544) );
  XNOR U14812 ( .A(n10537), .B(n10572), .Z(n10543) );
  XNOR U14813 ( .A(n10536), .B(n10538), .Z(n10572) );
  NAND U14814 ( .A(n10573), .B(n10574), .Z(n10538) );
  OR U14815 ( .A(n10575), .B(n10576), .Z(n10574) );
  OR U14816 ( .A(n10577), .B(n10578), .Z(n10573) );
  NAND U14817 ( .A(n10579), .B(n10580), .Z(n10536) );
  OR U14818 ( .A(n10581), .B(n10582), .Z(n10580) );
  OR U14819 ( .A(n10583), .B(n10584), .Z(n10579) );
  ANDN U14820 ( .B(n10585), .A(n10586), .Z(n10537) );
  IV U14821 ( .A(n10587), .Z(n10585) );
  ANDN U14822 ( .B(n10588), .A(n10589), .Z(n10529) );
  XOR U14823 ( .A(n10515), .B(n10590), .Z(n10527) );
  XOR U14824 ( .A(n10516), .B(n10517), .Z(n10590) );
  XOR U14825 ( .A(n10522), .B(n10591), .Z(n10517) );
  XOR U14826 ( .A(n10521), .B(n10524), .Z(n10591) );
  IV U14827 ( .A(n10523), .Z(n10524) );
  NAND U14828 ( .A(n10592), .B(n10593), .Z(n10523) );
  OR U14829 ( .A(n10594), .B(n10595), .Z(n10593) );
  OR U14830 ( .A(n10596), .B(n10597), .Z(n10592) );
  NAND U14831 ( .A(n10598), .B(n10599), .Z(n10521) );
  OR U14832 ( .A(n10600), .B(n10601), .Z(n10599) );
  OR U14833 ( .A(n10602), .B(n10603), .Z(n10598) );
  NOR U14834 ( .A(n10604), .B(n10605), .Z(n10522) );
  ANDN U14835 ( .B(n10606), .A(n10607), .Z(n10516) );
  IV U14836 ( .A(n10608), .Z(n10606) );
  XNOR U14837 ( .A(n10509), .B(n10609), .Z(n10515) );
  XNOR U14838 ( .A(n10508), .B(n10510), .Z(n10609) );
  NAND U14839 ( .A(n10610), .B(n10611), .Z(n10510) );
  OR U14840 ( .A(n10612), .B(n10613), .Z(n10611) );
  OR U14841 ( .A(n10614), .B(n10615), .Z(n10610) );
  NAND U14842 ( .A(n10616), .B(n10617), .Z(n10508) );
  OR U14843 ( .A(n10618), .B(n10619), .Z(n10617) );
  OR U14844 ( .A(n10620), .B(n10621), .Z(n10616) );
  ANDN U14845 ( .B(n10622), .A(n10623), .Z(n10509) );
  IV U14846 ( .A(n10624), .Z(n10622) );
  XNOR U14847 ( .A(n10589), .B(n10588), .Z(N29285) );
  XOR U14848 ( .A(n10608), .B(n10607), .Z(n10588) );
  XNOR U14849 ( .A(n10623), .B(n10624), .Z(n10607) );
  XNOR U14850 ( .A(n10618), .B(n10619), .Z(n10624) );
  XNOR U14851 ( .A(n10620), .B(n10621), .Z(n10619) );
  XNOR U14852 ( .A(y[2716]), .B(x[2716]), .Z(n10621) );
  XNOR U14853 ( .A(y[2717]), .B(x[2717]), .Z(n10620) );
  XNOR U14854 ( .A(y[2715]), .B(x[2715]), .Z(n10618) );
  XNOR U14855 ( .A(n10612), .B(n10613), .Z(n10623) );
  XNOR U14856 ( .A(y[2712]), .B(x[2712]), .Z(n10613) );
  XNOR U14857 ( .A(n10614), .B(n10615), .Z(n10612) );
  XNOR U14858 ( .A(y[2713]), .B(x[2713]), .Z(n10615) );
  XNOR U14859 ( .A(y[2714]), .B(x[2714]), .Z(n10614) );
  XNOR U14860 ( .A(n10605), .B(n10604), .Z(n10608) );
  XNOR U14861 ( .A(n10600), .B(n10601), .Z(n10604) );
  XNOR U14862 ( .A(y[2709]), .B(x[2709]), .Z(n10601) );
  XNOR U14863 ( .A(n10602), .B(n10603), .Z(n10600) );
  XNOR U14864 ( .A(y[2710]), .B(x[2710]), .Z(n10603) );
  XNOR U14865 ( .A(y[2711]), .B(x[2711]), .Z(n10602) );
  XNOR U14866 ( .A(n10594), .B(n10595), .Z(n10605) );
  XNOR U14867 ( .A(y[2706]), .B(x[2706]), .Z(n10595) );
  XNOR U14868 ( .A(n10596), .B(n10597), .Z(n10594) );
  XNOR U14869 ( .A(y[2707]), .B(x[2707]), .Z(n10597) );
  XNOR U14870 ( .A(y[2708]), .B(x[2708]), .Z(n10596) );
  XOR U14871 ( .A(n10570), .B(n10571), .Z(n10589) );
  XNOR U14872 ( .A(n10586), .B(n10587), .Z(n10571) );
  XNOR U14873 ( .A(n10581), .B(n10582), .Z(n10587) );
  XNOR U14874 ( .A(n10583), .B(n10584), .Z(n10582) );
  XNOR U14875 ( .A(y[2704]), .B(x[2704]), .Z(n10584) );
  XNOR U14876 ( .A(y[2705]), .B(x[2705]), .Z(n10583) );
  XNOR U14877 ( .A(y[2703]), .B(x[2703]), .Z(n10581) );
  XNOR U14878 ( .A(n10575), .B(n10576), .Z(n10586) );
  XNOR U14879 ( .A(y[2700]), .B(x[2700]), .Z(n10576) );
  XNOR U14880 ( .A(n10577), .B(n10578), .Z(n10575) );
  XNOR U14881 ( .A(y[2701]), .B(x[2701]), .Z(n10578) );
  XNOR U14882 ( .A(y[2702]), .B(x[2702]), .Z(n10577) );
  XOR U14883 ( .A(n10569), .B(n10568), .Z(n10570) );
  XNOR U14884 ( .A(n10564), .B(n10565), .Z(n10568) );
  XNOR U14885 ( .A(y[2697]), .B(x[2697]), .Z(n10565) );
  XNOR U14886 ( .A(n10566), .B(n10567), .Z(n10564) );
  XNOR U14887 ( .A(y[2698]), .B(x[2698]), .Z(n10567) );
  XNOR U14888 ( .A(y[2699]), .B(x[2699]), .Z(n10566) );
  XNOR U14889 ( .A(n10558), .B(n10559), .Z(n10569) );
  XNOR U14890 ( .A(y[2694]), .B(x[2694]), .Z(n10559) );
  XNOR U14891 ( .A(n10560), .B(n10561), .Z(n10558) );
  XNOR U14892 ( .A(y[2695]), .B(x[2695]), .Z(n10561) );
  XNOR U14893 ( .A(y[2696]), .B(x[2696]), .Z(n10560) );
  NAND U14894 ( .A(n10625), .B(n10626), .Z(N29277) );
  NANDN U14895 ( .A(n10627), .B(n10628), .Z(n10626) );
  OR U14896 ( .A(n10629), .B(n10630), .Z(n10628) );
  NAND U14897 ( .A(n10629), .B(n10630), .Z(n10625) );
  XOR U14898 ( .A(n10629), .B(n10631), .Z(N29276) );
  XNOR U14899 ( .A(n10627), .B(n10630), .Z(n10631) );
  AND U14900 ( .A(n10632), .B(n10633), .Z(n10630) );
  NANDN U14901 ( .A(n10634), .B(n10635), .Z(n10633) );
  NANDN U14902 ( .A(n10636), .B(n10637), .Z(n10635) );
  NANDN U14903 ( .A(n10637), .B(n10636), .Z(n10632) );
  NAND U14904 ( .A(n10638), .B(n10639), .Z(n10627) );
  NANDN U14905 ( .A(n10640), .B(n10641), .Z(n10639) );
  OR U14906 ( .A(n10642), .B(n10643), .Z(n10641) );
  NAND U14907 ( .A(n10643), .B(n10642), .Z(n10638) );
  AND U14908 ( .A(n10644), .B(n10645), .Z(n10629) );
  NANDN U14909 ( .A(n10646), .B(n10647), .Z(n10645) );
  NANDN U14910 ( .A(n10648), .B(n10649), .Z(n10647) );
  NANDN U14911 ( .A(n10649), .B(n10648), .Z(n10644) );
  XOR U14912 ( .A(n10643), .B(n10650), .Z(N29275) );
  XOR U14913 ( .A(n10640), .B(n10642), .Z(n10650) );
  XNOR U14914 ( .A(n10636), .B(n10651), .Z(n10642) );
  XNOR U14915 ( .A(n10634), .B(n10637), .Z(n10651) );
  NAND U14916 ( .A(n10652), .B(n10653), .Z(n10637) );
  NAND U14917 ( .A(n10654), .B(n10655), .Z(n10653) );
  OR U14918 ( .A(n10656), .B(n10657), .Z(n10654) );
  NANDN U14919 ( .A(n10658), .B(n10656), .Z(n10652) );
  IV U14920 ( .A(n10657), .Z(n10658) );
  NAND U14921 ( .A(n10659), .B(n10660), .Z(n10634) );
  NAND U14922 ( .A(n10661), .B(n10662), .Z(n10660) );
  NANDN U14923 ( .A(n10663), .B(n10664), .Z(n10661) );
  NANDN U14924 ( .A(n10664), .B(n10663), .Z(n10659) );
  AND U14925 ( .A(n10665), .B(n10666), .Z(n10636) );
  NAND U14926 ( .A(n10667), .B(n10668), .Z(n10666) );
  OR U14927 ( .A(n10669), .B(n10670), .Z(n10667) );
  NANDN U14928 ( .A(n10671), .B(n10669), .Z(n10665) );
  NAND U14929 ( .A(n10672), .B(n10673), .Z(n10640) );
  NANDN U14930 ( .A(n10674), .B(n10675), .Z(n10673) );
  OR U14931 ( .A(n10676), .B(n10677), .Z(n10675) );
  NANDN U14932 ( .A(n10678), .B(n10676), .Z(n10672) );
  IV U14933 ( .A(n10677), .Z(n10678) );
  XNOR U14934 ( .A(n10648), .B(n10679), .Z(n10643) );
  XNOR U14935 ( .A(n10646), .B(n10649), .Z(n10679) );
  NAND U14936 ( .A(n10680), .B(n10681), .Z(n10649) );
  NAND U14937 ( .A(n10682), .B(n10683), .Z(n10681) );
  OR U14938 ( .A(n10684), .B(n10685), .Z(n10682) );
  NANDN U14939 ( .A(n10686), .B(n10684), .Z(n10680) );
  IV U14940 ( .A(n10685), .Z(n10686) );
  NAND U14941 ( .A(n10687), .B(n10688), .Z(n10646) );
  NAND U14942 ( .A(n10689), .B(n10690), .Z(n10688) );
  NANDN U14943 ( .A(n10691), .B(n10692), .Z(n10689) );
  NANDN U14944 ( .A(n10692), .B(n10691), .Z(n10687) );
  AND U14945 ( .A(n10693), .B(n10694), .Z(n10648) );
  NAND U14946 ( .A(n10695), .B(n10696), .Z(n10694) );
  OR U14947 ( .A(n10697), .B(n10698), .Z(n10695) );
  NANDN U14948 ( .A(n10699), .B(n10697), .Z(n10693) );
  XNOR U14949 ( .A(n10674), .B(n10700), .Z(N29274) );
  XOR U14950 ( .A(n10676), .B(n10677), .Z(n10700) );
  XNOR U14951 ( .A(n10690), .B(n10701), .Z(n10677) );
  XOR U14952 ( .A(n10691), .B(n10692), .Z(n10701) );
  XOR U14953 ( .A(n10697), .B(n10702), .Z(n10692) );
  XOR U14954 ( .A(n10696), .B(n10699), .Z(n10702) );
  IV U14955 ( .A(n10698), .Z(n10699) );
  NAND U14956 ( .A(n10703), .B(n10704), .Z(n10698) );
  OR U14957 ( .A(n10705), .B(n10706), .Z(n10704) );
  OR U14958 ( .A(n10707), .B(n10708), .Z(n10703) );
  NAND U14959 ( .A(n10709), .B(n10710), .Z(n10696) );
  OR U14960 ( .A(n10711), .B(n10712), .Z(n10710) );
  OR U14961 ( .A(n10713), .B(n10714), .Z(n10709) );
  NOR U14962 ( .A(n10715), .B(n10716), .Z(n10697) );
  ANDN U14963 ( .B(n10717), .A(n10718), .Z(n10691) );
  XNOR U14964 ( .A(n10684), .B(n10719), .Z(n10690) );
  XNOR U14965 ( .A(n10683), .B(n10685), .Z(n10719) );
  NAND U14966 ( .A(n10720), .B(n10721), .Z(n10685) );
  OR U14967 ( .A(n10722), .B(n10723), .Z(n10721) );
  OR U14968 ( .A(n10724), .B(n10725), .Z(n10720) );
  NAND U14969 ( .A(n10726), .B(n10727), .Z(n10683) );
  OR U14970 ( .A(n10728), .B(n10729), .Z(n10727) );
  OR U14971 ( .A(n10730), .B(n10731), .Z(n10726) );
  ANDN U14972 ( .B(n10732), .A(n10733), .Z(n10684) );
  IV U14973 ( .A(n10734), .Z(n10732) );
  ANDN U14974 ( .B(n10735), .A(n10736), .Z(n10676) );
  XOR U14975 ( .A(n10662), .B(n10737), .Z(n10674) );
  XOR U14976 ( .A(n10663), .B(n10664), .Z(n10737) );
  XOR U14977 ( .A(n10669), .B(n10738), .Z(n10664) );
  XOR U14978 ( .A(n10668), .B(n10671), .Z(n10738) );
  IV U14979 ( .A(n10670), .Z(n10671) );
  NAND U14980 ( .A(n10739), .B(n10740), .Z(n10670) );
  OR U14981 ( .A(n10741), .B(n10742), .Z(n10740) );
  OR U14982 ( .A(n10743), .B(n10744), .Z(n10739) );
  NAND U14983 ( .A(n10745), .B(n10746), .Z(n10668) );
  OR U14984 ( .A(n10747), .B(n10748), .Z(n10746) );
  OR U14985 ( .A(n10749), .B(n10750), .Z(n10745) );
  NOR U14986 ( .A(n10751), .B(n10752), .Z(n10669) );
  ANDN U14987 ( .B(n10753), .A(n10754), .Z(n10663) );
  IV U14988 ( .A(n10755), .Z(n10753) );
  XNOR U14989 ( .A(n10656), .B(n10756), .Z(n10662) );
  XNOR U14990 ( .A(n10655), .B(n10657), .Z(n10756) );
  NAND U14991 ( .A(n10757), .B(n10758), .Z(n10657) );
  OR U14992 ( .A(n10759), .B(n10760), .Z(n10758) );
  OR U14993 ( .A(n10761), .B(n10762), .Z(n10757) );
  NAND U14994 ( .A(n10763), .B(n10764), .Z(n10655) );
  OR U14995 ( .A(n10765), .B(n10766), .Z(n10764) );
  OR U14996 ( .A(n10767), .B(n10768), .Z(n10763) );
  ANDN U14997 ( .B(n10769), .A(n10770), .Z(n10656) );
  IV U14998 ( .A(n10771), .Z(n10769) );
  XNOR U14999 ( .A(n10736), .B(n10735), .Z(N29273) );
  XOR U15000 ( .A(n10755), .B(n10754), .Z(n10735) );
  XNOR U15001 ( .A(n10770), .B(n10771), .Z(n10754) );
  XNOR U15002 ( .A(n10765), .B(n10766), .Z(n10771) );
  XNOR U15003 ( .A(n10767), .B(n10768), .Z(n10766) );
  XNOR U15004 ( .A(y[2692]), .B(x[2692]), .Z(n10768) );
  XNOR U15005 ( .A(y[2693]), .B(x[2693]), .Z(n10767) );
  XNOR U15006 ( .A(y[2691]), .B(x[2691]), .Z(n10765) );
  XNOR U15007 ( .A(n10759), .B(n10760), .Z(n10770) );
  XNOR U15008 ( .A(y[2688]), .B(x[2688]), .Z(n10760) );
  XNOR U15009 ( .A(n10761), .B(n10762), .Z(n10759) );
  XNOR U15010 ( .A(y[2689]), .B(x[2689]), .Z(n10762) );
  XNOR U15011 ( .A(y[2690]), .B(x[2690]), .Z(n10761) );
  XNOR U15012 ( .A(n10752), .B(n10751), .Z(n10755) );
  XNOR U15013 ( .A(n10747), .B(n10748), .Z(n10751) );
  XNOR U15014 ( .A(y[2685]), .B(x[2685]), .Z(n10748) );
  XNOR U15015 ( .A(n10749), .B(n10750), .Z(n10747) );
  XNOR U15016 ( .A(y[2686]), .B(x[2686]), .Z(n10750) );
  XNOR U15017 ( .A(y[2687]), .B(x[2687]), .Z(n10749) );
  XNOR U15018 ( .A(n10741), .B(n10742), .Z(n10752) );
  XNOR U15019 ( .A(y[2682]), .B(x[2682]), .Z(n10742) );
  XNOR U15020 ( .A(n10743), .B(n10744), .Z(n10741) );
  XNOR U15021 ( .A(y[2683]), .B(x[2683]), .Z(n10744) );
  XNOR U15022 ( .A(y[2684]), .B(x[2684]), .Z(n10743) );
  XOR U15023 ( .A(n10717), .B(n10718), .Z(n10736) );
  XNOR U15024 ( .A(n10733), .B(n10734), .Z(n10718) );
  XNOR U15025 ( .A(n10728), .B(n10729), .Z(n10734) );
  XNOR U15026 ( .A(n10730), .B(n10731), .Z(n10729) );
  XNOR U15027 ( .A(y[2680]), .B(x[2680]), .Z(n10731) );
  XNOR U15028 ( .A(y[2681]), .B(x[2681]), .Z(n10730) );
  XNOR U15029 ( .A(y[2679]), .B(x[2679]), .Z(n10728) );
  XNOR U15030 ( .A(n10722), .B(n10723), .Z(n10733) );
  XNOR U15031 ( .A(y[2676]), .B(x[2676]), .Z(n10723) );
  XNOR U15032 ( .A(n10724), .B(n10725), .Z(n10722) );
  XNOR U15033 ( .A(y[2677]), .B(x[2677]), .Z(n10725) );
  XNOR U15034 ( .A(y[2678]), .B(x[2678]), .Z(n10724) );
  XOR U15035 ( .A(n10716), .B(n10715), .Z(n10717) );
  XNOR U15036 ( .A(n10711), .B(n10712), .Z(n10715) );
  XNOR U15037 ( .A(y[2673]), .B(x[2673]), .Z(n10712) );
  XNOR U15038 ( .A(n10713), .B(n10714), .Z(n10711) );
  XNOR U15039 ( .A(y[2674]), .B(x[2674]), .Z(n10714) );
  XNOR U15040 ( .A(y[2675]), .B(x[2675]), .Z(n10713) );
  XNOR U15041 ( .A(n10705), .B(n10706), .Z(n10716) );
  XNOR U15042 ( .A(y[2670]), .B(x[2670]), .Z(n10706) );
  XNOR U15043 ( .A(n10707), .B(n10708), .Z(n10705) );
  XNOR U15044 ( .A(y[2671]), .B(x[2671]), .Z(n10708) );
  XNOR U15045 ( .A(y[2672]), .B(x[2672]), .Z(n10707) );
  NAND U15046 ( .A(n10772), .B(n10773), .Z(N29265) );
  NANDN U15047 ( .A(n10774), .B(n10775), .Z(n10773) );
  OR U15048 ( .A(n10776), .B(n10777), .Z(n10775) );
  NAND U15049 ( .A(n10776), .B(n10777), .Z(n10772) );
  XOR U15050 ( .A(n10776), .B(n10778), .Z(N29264) );
  XNOR U15051 ( .A(n10774), .B(n10777), .Z(n10778) );
  AND U15052 ( .A(n10779), .B(n10780), .Z(n10777) );
  NANDN U15053 ( .A(n10781), .B(n10782), .Z(n10780) );
  NANDN U15054 ( .A(n10783), .B(n10784), .Z(n10782) );
  NANDN U15055 ( .A(n10784), .B(n10783), .Z(n10779) );
  NAND U15056 ( .A(n10785), .B(n10786), .Z(n10774) );
  NANDN U15057 ( .A(n10787), .B(n10788), .Z(n10786) );
  OR U15058 ( .A(n10789), .B(n10790), .Z(n10788) );
  NAND U15059 ( .A(n10790), .B(n10789), .Z(n10785) );
  AND U15060 ( .A(n10791), .B(n10792), .Z(n10776) );
  NANDN U15061 ( .A(n10793), .B(n10794), .Z(n10792) );
  NANDN U15062 ( .A(n10795), .B(n10796), .Z(n10794) );
  NANDN U15063 ( .A(n10796), .B(n10795), .Z(n10791) );
  XOR U15064 ( .A(n10790), .B(n10797), .Z(N29263) );
  XOR U15065 ( .A(n10787), .B(n10789), .Z(n10797) );
  XNOR U15066 ( .A(n10783), .B(n10798), .Z(n10789) );
  XNOR U15067 ( .A(n10781), .B(n10784), .Z(n10798) );
  NAND U15068 ( .A(n10799), .B(n10800), .Z(n10784) );
  NAND U15069 ( .A(n10801), .B(n10802), .Z(n10800) );
  OR U15070 ( .A(n10803), .B(n10804), .Z(n10801) );
  NANDN U15071 ( .A(n10805), .B(n10803), .Z(n10799) );
  IV U15072 ( .A(n10804), .Z(n10805) );
  NAND U15073 ( .A(n10806), .B(n10807), .Z(n10781) );
  NAND U15074 ( .A(n10808), .B(n10809), .Z(n10807) );
  NANDN U15075 ( .A(n10810), .B(n10811), .Z(n10808) );
  NANDN U15076 ( .A(n10811), .B(n10810), .Z(n10806) );
  AND U15077 ( .A(n10812), .B(n10813), .Z(n10783) );
  NAND U15078 ( .A(n10814), .B(n10815), .Z(n10813) );
  OR U15079 ( .A(n10816), .B(n10817), .Z(n10814) );
  NANDN U15080 ( .A(n10818), .B(n10816), .Z(n10812) );
  NAND U15081 ( .A(n10819), .B(n10820), .Z(n10787) );
  NANDN U15082 ( .A(n10821), .B(n10822), .Z(n10820) );
  OR U15083 ( .A(n10823), .B(n10824), .Z(n10822) );
  NANDN U15084 ( .A(n10825), .B(n10823), .Z(n10819) );
  IV U15085 ( .A(n10824), .Z(n10825) );
  XNOR U15086 ( .A(n10795), .B(n10826), .Z(n10790) );
  XNOR U15087 ( .A(n10793), .B(n10796), .Z(n10826) );
  NAND U15088 ( .A(n10827), .B(n10828), .Z(n10796) );
  NAND U15089 ( .A(n10829), .B(n10830), .Z(n10828) );
  OR U15090 ( .A(n10831), .B(n10832), .Z(n10829) );
  NANDN U15091 ( .A(n10833), .B(n10831), .Z(n10827) );
  IV U15092 ( .A(n10832), .Z(n10833) );
  NAND U15093 ( .A(n10834), .B(n10835), .Z(n10793) );
  NAND U15094 ( .A(n10836), .B(n10837), .Z(n10835) );
  NANDN U15095 ( .A(n10838), .B(n10839), .Z(n10836) );
  NANDN U15096 ( .A(n10839), .B(n10838), .Z(n10834) );
  AND U15097 ( .A(n10840), .B(n10841), .Z(n10795) );
  NAND U15098 ( .A(n10842), .B(n10843), .Z(n10841) );
  OR U15099 ( .A(n10844), .B(n10845), .Z(n10842) );
  NANDN U15100 ( .A(n10846), .B(n10844), .Z(n10840) );
  XNOR U15101 ( .A(n10821), .B(n10847), .Z(N29262) );
  XOR U15102 ( .A(n10823), .B(n10824), .Z(n10847) );
  XNOR U15103 ( .A(n10837), .B(n10848), .Z(n10824) );
  XOR U15104 ( .A(n10838), .B(n10839), .Z(n10848) );
  XOR U15105 ( .A(n10844), .B(n10849), .Z(n10839) );
  XOR U15106 ( .A(n10843), .B(n10846), .Z(n10849) );
  IV U15107 ( .A(n10845), .Z(n10846) );
  NAND U15108 ( .A(n10850), .B(n10851), .Z(n10845) );
  OR U15109 ( .A(n10852), .B(n10853), .Z(n10851) );
  OR U15110 ( .A(n10854), .B(n10855), .Z(n10850) );
  NAND U15111 ( .A(n10856), .B(n10857), .Z(n10843) );
  OR U15112 ( .A(n10858), .B(n10859), .Z(n10857) );
  OR U15113 ( .A(n10860), .B(n10861), .Z(n10856) );
  NOR U15114 ( .A(n10862), .B(n10863), .Z(n10844) );
  ANDN U15115 ( .B(n10864), .A(n10865), .Z(n10838) );
  XNOR U15116 ( .A(n10831), .B(n10866), .Z(n10837) );
  XNOR U15117 ( .A(n10830), .B(n10832), .Z(n10866) );
  NAND U15118 ( .A(n10867), .B(n10868), .Z(n10832) );
  OR U15119 ( .A(n10869), .B(n10870), .Z(n10868) );
  OR U15120 ( .A(n10871), .B(n10872), .Z(n10867) );
  NAND U15121 ( .A(n10873), .B(n10874), .Z(n10830) );
  OR U15122 ( .A(n10875), .B(n10876), .Z(n10874) );
  OR U15123 ( .A(n10877), .B(n10878), .Z(n10873) );
  ANDN U15124 ( .B(n10879), .A(n10880), .Z(n10831) );
  IV U15125 ( .A(n10881), .Z(n10879) );
  ANDN U15126 ( .B(n10882), .A(n10883), .Z(n10823) );
  XOR U15127 ( .A(n10809), .B(n10884), .Z(n10821) );
  XOR U15128 ( .A(n10810), .B(n10811), .Z(n10884) );
  XOR U15129 ( .A(n10816), .B(n10885), .Z(n10811) );
  XOR U15130 ( .A(n10815), .B(n10818), .Z(n10885) );
  IV U15131 ( .A(n10817), .Z(n10818) );
  NAND U15132 ( .A(n10886), .B(n10887), .Z(n10817) );
  OR U15133 ( .A(n10888), .B(n10889), .Z(n10887) );
  OR U15134 ( .A(n10890), .B(n10891), .Z(n10886) );
  NAND U15135 ( .A(n10892), .B(n10893), .Z(n10815) );
  OR U15136 ( .A(n10894), .B(n10895), .Z(n10893) );
  OR U15137 ( .A(n10896), .B(n10897), .Z(n10892) );
  NOR U15138 ( .A(n10898), .B(n10899), .Z(n10816) );
  ANDN U15139 ( .B(n10900), .A(n10901), .Z(n10810) );
  IV U15140 ( .A(n10902), .Z(n10900) );
  XNOR U15141 ( .A(n10803), .B(n10903), .Z(n10809) );
  XNOR U15142 ( .A(n10802), .B(n10804), .Z(n10903) );
  NAND U15143 ( .A(n10904), .B(n10905), .Z(n10804) );
  OR U15144 ( .A(n10906), .B(n10907), .Z(n10905) );
  OR U15145 ( .A(n10908), .B(n10909), .Z(n10904) );
  NAND U15146 ( .A(n10910), .B(n10911), .Z(n10802) );
  OR U15147 ( .A(n10912), .B(n10913), .Z(n10911) );
  OR U15148 ( .A(n10914), .B(n10915), .Z(n10910) );
  ANDN U15149 ( .B(n10916), .A(n10917), .Z(n10803) );
  IV U15150 ( .A(n10918), .Z(n10916) );
  XNOR U15151 ( .A(n10883), .B(n10882), .Z(N29261) );
  XOR U15152 ( .A(n10902), .B(n10901), .Z(n10882) );
  XNOR U15153 ( .A(n10917), .B(n10918), .Z(n10901) );
  XNOR U15154 ( .A(n10912), .B(n10913), .Z(n10918) );
  XNOR U15155 ( .A(n10914), .B(n10915), .Z(n10913) );
  XNOR U15156 ( .A(y[2668]), .B(x[2668]), .Z(n10915) );
  XNOR U15157 ( .A(y[2669]), .B(x[2669]), .Z(n10914) );
  XNOR U15158 ( .A(y[2667]), .B(x[2667]), .Z(n10912) );
  XNOR U15159 ( .A(n10906), .B(n10907), .Z(n10917) );
  XNOR U15160 ( .A(y[2664]), .B(x[2664]), .Z(n10907) );
  XNOR U15161 ( .A(n10908), .B(n10909), .Z(n10906) );
  XNOR U15162 ( .A(y[2665]), .B(x[2665]), .Z(n10909) );
  XNOR U15163 ( .A(y[2666]), .B(x[2666]), .Z(n10908) );
  XNOR U15164 ( .A(n10899), .B(n10898), .Z(n10902) );
  XNOR U15165 ( .A(n10894), .B(n10895), .Z(n10898) );
  XNOR U15166 ( .A(y[2661]), .B(x[2661]), .Z(n10895) );
  XNOR U15167 ( .A(n10896), .B(n10897), .Z(n10894) );
  XNOR U15168 ( .A(y[2662]), .B(x[2662]), .Z(n10897) );
  XNOR U15169 ( .A(y[2663]), .B(x[2663]), .Z(n10896) );
  XNOR U15170 ( .A(n10888), .B(n10889), .Z(n10899) );
  XNOR U15171 ( .A(y[2658]), .B(x[2658]), .Z(n10889) );
  XNOR U15172 ( .A(n10890), .B(n10891), .Z(n10888) );
  XNOR U15173 ( .A(y[2659]), .B(x[2659]), .Z(n10891) );
  XNOR U15174 ( .A(y[2660]), .B(x[2660]), .Z(n10890) );
  XOR U15175 ( .A(n10864), .B(n10865), .Z(n10883) );
  XNOR U15176 ( .A(n10880), .B(n10881), .Z(n10865) );
  XNOR U15177 ( .A(n10875), .B(n10876), .Z(n10881) );
  XNOR U15178 ( .A(n10877), .B(n10878), .Z(n10876) );
  XNOR U15179 ( .A(y[2656]), .B(x[2656]), .Z(n10878) );
  XNOR U15180 ( .A(y[2657]), .B(x[2657]), .Z(n10877) );
  XNOR U15181 ( .A(y[2655]), .B(x[2655]), .Z(n10875) );
  XNOR U15182 ( .A(n10869), .B(n10870), .Z(n10880) );
  XNOR U15183 ( .A(y[2652]), .B(x[2652]), .Z(n10870) );
  XNOR U15184 ( .A(n10871), .B(n10872), .Z(n10869) );
  XNOR U15185 ( .A(y[2653]), .B(x[2653]), .Z(n10872) );
  XNOR U15186 ( .A(y[2654]), .B(x[2654]), .Z(n10871) );
  XOR U15187 ( .A(n10863), .B(n10862), .Z(n10864) );
  XNOR U15188 ( .A(n10858), .B(n10859), .Z(n10862) );
  XNOR U15189 ( .A(y[2649]), .B(x[2649]), .Z(n10859) );
  XNOR U15190 ( .A(n10860), .B(n10861), .Z(n10858) );
  XNOR U15191 ( .A(y[2650]), .B(x[2650]), .Z(n10861) );
  XNOR U15192 ( .A(y[2651]), .B(x[2651]), .Z(n10860) );
  XNOR U15193 ( .A(n10852), .B(n10853), .Z(n10863) );
  XNOR U15194 ( .A(y[2646]), .B(x[2646]), .Z(n10853) );
  XNOR U15195 ( .A(n10854), .B(n10855), .Z(n10852) );
  XNOR U15196 ( .A(y[2647]), .B(x[2647]), .Z(n10855) );
  XNOR U15197 ( .A(y[2648]), .B(x[2648]), .Z(n10854) );
  NAND U15198 ( .A(n10919), .B(n10920), .Z(N29253) );
  NANDN U15199 ( .A(n10921), .B(n10922), .Z(n10920) );
  OR U15200 ( .A(n10923), .B(n10924), .Z(n10922) );
  NAND U15201 ( .A(n10923), .B(n10924), .Z(n10919) );
  XOR U15202 ( .A(n10923), .B(n10925), .Z(N29252) );
  XNOR U15203 ( .A(n10921), .B(n10924), .Z(n10925) );
  AND U15204 ( .A(n10926), .B(n10927), .Z(n10924) );
  NANDN U15205 ( .A(n10928), .B(n10929), .Z(n10927) );
  NANDN U15206 ( .A(n10930), .B(n10931), .Z(n10929) );
  NANDN U15207 ( .A(n10931), .B(n10930), .Z(n10926) );
  NAND U15208 ( .A(n10932), .B(n10933), .Z(n10921) );
  NANDN U15209 ( .A(n10934), .B(n10935), .Z(n10933) );
  OR U15210 ( .A(n10936), .B(n10937), .Z(n10935) );
  NAND U15211 ( .A(n10937), .B(n10936), .Z(n10932) );
  AND U15212 ( .A(n10938), .B(n10939), .Z(n10923) );
  NANDN U15213 ( .A(n10940), .B(n10941), .Z(n10939) );
  NANDN U15214 ( .A(n10942), .B(n10943), .Z(n10941) );
  NANDN U15215 ( .A(n10943), .B(n10942), .Z(n10938) );
  XOR U15216 ( .A(n10937), .B(n10944), .Z(N29251) );
  XOR U15217 ( .A(n10934), .B(n10936), .Z(n10944) );
  XNOR U15218 ( .A(n10930), .B(n10945), .Z(n10936) );
  XNOR U15219 ( .A(n10928), .B(n10931), .Z(n10945) );
  NAND U15220 ( .A(n10946), .B(n10947), .Z(n10931) );
  NAND U15221 ( .A(n10948), .B(n10949), .Z(n10947) );
  OR U15222 ( .A(n10950), .B(n10951), .Z(n10948) );
  NANDN U15223 ( .A(n10952), .B(n10950), .Z(n10946) );
  IV U15224 ( .A(n10951), .Z(n10952) );
  NAND U15225 ( .A(n10953), .B(n10954), .Z(n10928) );
  NAND U15226 ( .A(n10955), .B(n10956), .Z(n10954) );
  NANDN U15227 ( .A(n10957), .B(n10958), .Z(n10955) );
  NANDN U15228 ( .A(n10958), .B(n10957), .Z(n10953) );
  AND U15229 ( .A(n10959), .B(n10960), .Z(n10930) );
  NAND U15230 ( .A(n10961), .B(n10962), .Z(n10960) );
  OR U15231 ( .A(n10963), .B(n10964), .Z(n10961) );
  NANDN U15232 ( .A(n10965), .B(n10963), .Z(n10959) );
  NAND U15233 ( .A(n10966), .B(n10967), .Z(n10934) );
  NANDN U15234 ( .A(n10968), .B(n10969), .Z(n10967) );
  OR U15235 ( .A(n10970), .B(n10971), .Z(n10969) );
  NANDN U15236 ( .A(n10972), .B(n10970), .Z(n10966) );
  IV U15237 ( .A(n10971), .Z(n10972) );
  XNOR U15238 ( .A(n10942), .B(n10973), .Z(n10937) );
  XNOR U15239 ( .A(n10940), .B(n10943), .Z(n10973) );
  NAND U15240 ( .A(n10974), .B(n10975), .Z(n10943) );
  NAND U15241 ( .A(n10976), .B(n10977), .Z(n10975) );
  OR U15242 ( .A(n10978), .B(n10979), .Z(n10976) );
  NANDN U15243 ( .A(n10980), .B(n10978), .Z(n10974) );
  IV U15244 ( .A(n10979), .Z(n10980) );
  NAND U15245 ( .A(n10981), .B(n10982), .Z(n10940) );
  NAND U15246 ( .A(n10983), .B(n10984), .Z(n10982) );
  NANDN U15247 ( .A(n10985), .B(n10986), .Z(n10983) );
  NANDN U15248 ( .A(n10986), .B(n10985), .Z(n10981) );
  AND U15249 ( .A(n10987), .B(n10988), .Z(n10942) );
  NAND U15250 ( .A(n10989), .B(n10990), .Z(n10988) );
  OR U15251 ( .A(n10991), .B(n10992), .Z(n10989) );
  NANDN U15252 ( .A(n10993), .B(n10991), .Z(n10987) );
  XNOR U15253 ( .A(n10968), .B(n10994), .Z(N29250) );
  XOR U15254 ( .A(n10970), .B(n10971), .Z(n10994) );
  XNOR U15255 ( .A(n10984), .B(n10995), .Z(n10971) );
  XOR U15256 ( .A(n10985), .B(n10986), .Z(n10995) );
  XOR U15257 ( .A(n10991), .B(n10996), .Z(n10986) );
  XOR U15258 ( .A(n10990), .B(n10993), .Z(n10996) );
  IV U15259 ( .A(n10992), .Z(n10993) );
  NAND U15260 ( .A(n10997), .B(n10998), .Z(n10992) );
  OR U15261 ( .A(n10999), .B(n11000), .Z(n10998) );
  OR U15262 ( .A(n11001), .B(n11002), .Z(n10997) );
  NAND U15263 ( .A(n11003), .B(n11004), .Z(n10990) );
  OR U15264 ( .A(n11005), .B(n11006), .Z(n11004) );
  OR U15265 ( .A(n11007), .B(n11008), .Z(n11003) );
  NOR U15266 ( .A(n11009), .B(n11010), .Z(n10991) );
  ANDN U15267 ( .B(n11011), .A(n11012), .Z(n10985) );
  XNOR U15268 ( .A(n10978), .B(n11013), .Z(n10984) );
  XNOR U15269 ( .A(n10977), .B(n10979), .Z(n11013) );
  NAND U15270 ( .A(n11014), .B(n11015), .Z(n10979) );
  OR U15271 ( .A(n11016), .B(n11017), .Z(n11015) );
  OR U15272 ( .A(n11018), .B(n11019), .Z(n11014) );
  NAND U15273 ( .A(n11020), .B(n11021), .Z(n10977) );
  OR U15274 ( .A(n11022), .B(n11023), .Z(n11021) );
  OR U15275 ( .A(n11024), .B(n11025), .Z(n11020) );
  ANDN U15276 ( .B(n11026), .A(n11027), .Z(n10978) );
  IV U15277 ( .A(n11028), .Z(n11026) );
  ANDN U15278 ( .B(n11029), .A(n11030), .Z(n10970) );
  XOR U15279 ( .A(n10956), .B(n11031), .Z(n10968) );
  XOR U15280 ( .A(n10957), .B(n10958), .Z(n11031) );
  XOR U15281 ( .A(n10963), .B(n11032), .Z(n10958) );
  XOR U15282 ( .A(n10962), .B(n10965), .Z(n11032) );
  IV U15283 ( .A(n10964), .Z(n10965) );
  NAND U15284 ( .A(n11033), .B(n11034), .Z(n10964) );
  OR U15285 ( .A(n11035), .B(n11036), .Z(n11034) );
  OR U15286 ( .A(n11037), .B(n11038), .Z(n11033) );
  NAND U15287 ( .A(n11039), .B(n11040), .Z(n10962) );
  OR U15288 ( .A(n11041), .B(n11042), .Z(n11040) );
  OR U15289 ( .A(n11043), .B(n11044), .Z(n11039) );
  NOR U15290 ( .A(n11045), .B(n11046), .Z(n10963) );
  ANDN U15291 ( .B(n11047), .A(n11048), .Z(n10957) );
  IV U15292 ( .A(n11049), .Z(n11047) );
  XNOR U15293 ( .A(n10950), .B(n11050), .Z(n10956) );
  XNOR U15294 ( .A(n10949), .B(n10951), .Z(n11050) );
  NAND U15295 ( .A(n11051), .B(n11052), .Z(n10951) );
  OR U15296 ( .A(n11053), .B(n11054), .Z(n11052) );
  OR U15297 ( .A(n11055), .B(n11056), .Z(n11051) );
  NAND U15298 ( .A(n11057), .B(n11058), .Z(n10949) );
  OR U15299 ( .A(n11059), .B(n11060), .Z(n11058) );
  OR U15300 ( .A(n11061), .B(n11062), .Z(n11057) );
  ANDN U15301 ( .B(n11063), .A(n11064), .Z(n10950) );
  IV U15302 ( .A(n11065), .Z(n11063) );
  XNOR U15303 ( .A(n11030), .B(n11029), .Z(N29249) );
  XOR U15304 ( .A(n11049), .B(n11048), .Z(n11029) );
  XNOR U15305 ( .A(n11064), .B(n11065), .Z(n11048) );
  XNOR U15306 ( .A(n11059), .B(n11060), .Z(n11065) );
  XNOR U15307 ( .A(n11061), .B(n11062), .Z(n11060) );
  XNOR U15308 ( .A(y[2644]), .B(x[2644]), .Z(n11062) );
  XNOR U15309 ( .A(y[2645]), .B(x[2645]), .Z(n11061) );
  XNOR U15310 ( .A(y[2643]), .B(x[2643]), .Z(n11059) );
  XNOR U15311 ( .A(n11053), .B(n11054), .Z(n11064) );
  XNOR U15312 ( .A(y[2640]), .B(x[2640]), .Z(n11054) );
  XNOR U15313 ( .A(n11055), .B(n11056), .Z(n11053) );
  XNOR U15314 ( .A(y[2641]), .B(x[2641]), .Z(n11056) );
  XNOR U15315 ( .A(y[2642]), .B(x[2642]), .Z(n11055) );
  XNOR U15316 ( .A(n11046), .B(n11045), .Z(n11049) );
  XNOR U15317 ( .A(n11041), .B(n11042), .Z(n11045) );
  XNOR U15318 ( .A(y[2637]), .B(x[2637]), .Z(n11042) );
  XNOR U15319 ( .A(n11043), .B(n11044), .Z(n11041) );
  XNOR U15320 ( .A(y[2638]), .B(x[2638]), .Z(n11044) );
  XNOR U15321 ( .A(y[2639]), .B(x[2639]), .Z(n11043) );
  XNOR U15322 ( .A(n11035), .B(n11036), .Z(n11046) );
  XNOR U15323 ( .A(y[2634]), .B(x[2634]), .Z(n11036) );
  XNOR U15324 ( .A(n11037), .B(n11038), .Z(n11035) );
  XNOR U15325 ( .A(y[2635]), .B(x[2635]), .Z(n11038) );
  XNOR U15326 ( .A(y[2636]), .B(x[2636]), .Z(n11037) );
  XOR U15327 ( .A(n11011), .B(n11012), .Z(n11030) );
  XNOR U15328 ( .A(n11027), .B(n11028), .Z(n11012) );
  XNOR U15329 ( .A(n11022), .B(n11023), .Z(n11028) );
  XNOR U15330 ( .A(n11024), .B(n11025), .Z(n11023) );
  XNOR U15331 ( .A(y[2632]), .B(x[2632]), .Z(n11025) );
  XNOR U15332 ( .A(y[2633]), .B(x[2633]), .Z(n11024) );
  XNOR U15333 ( .A(y[2631]), .B(x[2631]), .Z(n11022) );
  XNOR U15334 ( .A(n11016), .B(n11017), .Z(n11027) );
  XNOR U15335 ( .A(y[2628]), .B(x[2628]), .Z(n11017) );
  XNOR U15336 ( .A(n11018), .B(n11019), .Z(n11016) );
  XNOR U15337 ( .A(y[2629]), .B(x[2629]), .Z(n11019) );
  XNOR U15338 ( .A(y[2630]), .B(x[2630]), .Z(n11018) );
  XOR U15339 ( .A(n11010), .B(n11009), .Z(n11011) );
  XNOR U15340 ( .A(n11005), .B(n11006), .Z(n11009) );
  XNOR U15341 ( .A(y[2625]), .B(x[2625]), .Z(n11006) );
  XNOR U15342 ( .A(n11007), .B(n11008), .Z(n11005) );
  XNOR U15343 ( .A(y[2626]), .B(x[2626]), .Z(n11008) );
  XNOR U15344 ( .A(y[2627]), .B(x[2627]), .Z(n11007) );
  XNOR U15345 ( .A(n10999), .B(n11000), .Z(n11010) );
  XNOR U15346 ( .A(y[2622]), .B(x[2622]), .Z(n11000) );
  XNOR U15347 ( .A(n11001), .B(n11002), .Z(n10999) );
  XNOR U15348 ( .A(y[2623]), .B(x[2623]), .Z(n11002) );
  XNOR U15349 ( .A(y[2624]), .B(x[2624]), .Z(n11001) );
  NAND U15350 ( .A(n11066), .B(n11067), .Z(N29241) );
  NANDN U15351 ( .A(n11068), .B(n11069), .Z(n11067) );
  OR U15352 ( .A(n11070), .B(n11071), .Z(n11069) );
  NAND U15353 ( .A(n11070), .B(n11071), .Z(n11066) );
  XOR U15354 ( .A(n11070), .B(n11072), .Z(N29240) );
  XNOR U15355 ( .A(n11068), .B(n11071), .Z(n11072) );
  AND U15356 ( .A(n11073), .B(n11074), .Z(n11071) );
  NANDN U15357 ( .A(n11075), .B(n11076), .Z(n11074) );
  NANDN U15358 ( .A(n11077), .B(n11078), .Z(n11076) );
  NANDN U15359 ( .A(n11078), .B(n11077), .Z(n11073) );
  NAND U15360 ( .A(n11079), .B(n11080), .Z(n11068) );
  NANDN U15361 ( .A(n11081), .B(n11082), .Z(n11080) );
  OR U15362 ( .A(n11083), .B(n11084), .Z(n11082) );
  NAND U15363 ( .A(n11084), .B(n11083), .Z(n11079) );
  AND U15364 ( .A(n11085), .B(n11086), .Z(n11070) );
  NANDN U15365 ( .A(n11087), .B(n11088), .Z(n11086) );
  NANDN U15366 ( .A(n11089), .B(n11090), .Z(n11088) );
  NANDN U15367 ( .A(n11090), .B(n11089), .Z(n11085) );
  XOR U15368 ( .A(n11084), .B(n11091), .Z(N29239) );
  XOR U15369 ( .A(n11081), .B(n11083), .Z(n11091) );
  XNOR U15370 ( .A(n11077), .B(n11092), .Z(n11083) );
  XNOR U15371 ( .A(n11075), .B(n11078), .Z(n11092) );
  NAND U15372 ( .A(n11093), .B(n11094), .Z(n11078) );
  NAND U15373 ( .A(n11095), .B(n11096), .Z(n11094) );
  OR U15374 ( .A(n11097), .B(n11098), .Z(n11095) );
  NANDN U15375 ( .A(n11099), .B(n11097), .Z(n11093) );
  IV U15376 ( .A(n11098), .Z(n11099) );
  NAND U15377 ( .A(n11100), .B(n11101), .Z(n11075) );
  NAND U15378 ( .A(n11102), .B(n11103), .Z(n11101) );
  NANDN U15379 ( .A(n11104), .B(n11105), .Z(n11102) );
  NANDN U15380 ( .A(n11105), .B(n11104), .Z(n11100) );
  AND U15381 ( .A(n11106), .B(n11107), .Z(n11077) );
  NAND U15382 ( .A(n11108), .B(n11109), .Z(n11107) );
  OR U15383 ( .A(n11110), .B(n11111), .Z(n11108) );
  NANDN U15384 ( .A(n11112), .B(n11110), .Z(n11106) );
  NAND U15385 ( .A(n11113), .B(n11114), .Z(n11081) );
  NANDN U15386 ( .A(n11115), .B(n11116), .Z(n11114) );
  OR U15387 ( .A(n11117), .B(n11118), .Z(n11116) );
  NANDN U15388 ( .A(n11119), .B(n11117), .Z(n11113) );
  IV U15389 ( .A(n11118), .Z(n11119) );
  XNOR U15390 ( .A(n11089), .B(n11120), .Z(n11084) );
  XNOR U15391 ( .A(n11087), .B(n11090), .Z(n11120) );
  NAND U15392 ( .A(n11121), .B(n11122), .Z(n11090) );
  NAND U15393 ( .A(n11123), .B(n11124), .Z(n11122) );
  OR U15394 ( .A(n11125), .B(n11126), .Z(n11123) );
  NANDN U15395 ( .A(n11127), .B(n11125), .Z(n11121) );
  IV U15396 ( .A(n11126), .Z(n11127) );
  NAND U15397 ( .A(n11128), .B(n11129), .Z(n11087) );
  NAND U15398 ( .A(n11130), .B(n11131), .Z(n11129) );
  NANDN U15399 ( .A(n11132), .B(n11133), .Z(n11130) );
  NANDN U15400 ( .A(n11133), .B(n11132), .Z(n11128) );
  AND U15401 ( .A(n11134), .B(n11135), .Z(n11089) );
  NAND U15402 ( .A(n11136), .B(n11137), .Z(n11135) );
  OR U15403 ( .A(n11138), .B(n11139), .Z(n11136) );
  NANDN U15404 ( .A(n11140), .B(n11138), .Z(n11134) );
  XNOR U15405 ( .A(n11115), .B(n11141), .Z(N29238) );
  XOR U15406 ( .A(n11117), .B(n11118), .Z(n11141) );
  XNOR U15407 ( .A(n11131), .B(n11142), .Z(n11118) );
  XOR U15408 ( .A(n11132), .B(n11133), .Z(n11142) );
  XOR U15409 ( .A(n11138), .B(n11143), .Z(n11133) );
  XOR U15410 ( .A(n11137), .B(n11140), .Z(n11143) );
  IV U15411 ( .A(n11139), .Z(n11140) );
  NAND U15412 ( .A(n11144), .B(n11145), .Z(n11139) );
  OR U15413 ( .A(n11146), .B(n11147), .Z(n11145) );
  OR U15414 ( .A(n11148), .B(n11149), .Z(n11144) );
  NAND U15415 ( .A(n11150), .B(n11151), .Z(n11137) );
  OR U15416 ( .A(n11152), .B(n11153), .Z(n11151) );
  OR U15417 ( .A(n11154), .B(n11155), .Z(n11150) );
  NOR U15418 ( .A(n11156), .B(n11157), .Z(n11138) );
  ANDN U15419 ( .B(n11158), .A(n11159), .Z(n11132) );
  XNOR U15420 ( .A(n11125), .B(n11160), .Z(n11131) );
  XNOR U15421 ( .A(n11124), .B(n11126), .Z(n11160) );
  NAND U15422 ( .A(n11161), .B(n11162), .Z(n11126) );
  OR U15423 ( .A(n11163), .B(n11164), .Z(n11162) );
  OR U15424 ( .A(n11165), .B(n11166), .Z(n11161) );
  NAND U15425 ( .A(n11167), .B(n11168), .Z(n11124) );
  OR U15426 ( .A(n11169), .B(n11170), .Z(n11168) );
  OR U15427 ( .A(n11171), .B(n11172), .Z(n11167) );
  ANDN U15428 ( .B(n11173), .A(n11174), .Z(n11125) );
  IV U15429 ( .A(n11175), .Z(n11173) );
  ANDN U15430 ( .B(n11176), .A(n11177), .Z(n11117) );
  XOR U15431 ( .A(n11103), .B(n11178), .Z(n11115) );
  XOR U15432 ( .A(n11104), .B(n11105), .Z(n11178) );
  XOR U15433 ( .A(n11110), .B(n11179), .Z(n11105) );
  XOR U15434 ( .A(n11109), .B(n11112), .Z(n11179) );
  IV U15435 ( .A(n11111), .Z(n11112) );
  NAND U15436 ( .A(n11180), .B(n11181), .Z(n11111) );
  OR U15437 ( .A(n11182), .B(n11183), .Z(n11181) );
  OR U15438 ( .A(n11184), .B(n11185), .Z(n11180) );
  NAND U15439 ( .A(n11186), .B(n11187), .Z(n11109) );
  OR U15440 ( .A(n11188), .B(n11189), .Z(n11187) );
  OR U15441 ( .A(n11190), .B(n11191), .Z(n11186) );
  NOR U15442 ( .A(n11192), .B(n11193), .Z(n11110) );
  ANDN U15443 ( .B(n11194), .A(n11195), .Z(n11104) );
  IV U15444 ( .A(n11196), .Z(n11194) );
  XNOR U15445 ( .A(n11097), .B(n11197), .Z(n11103) );
  XNOR U15446 ( .A(n11096), .B(n11098), .Z(n11197) );
  NAND U15447 ( .A(n11198), .B(n11199), .Z(n11098) );
  OR U15448 ( .A(n11200), .B(n11201), .Z(n11199) );
  OR U15449 ( .A(n11202), .B(n11203), .Z(n11198) );
  NAND U15450 ( .A(n11204), .B(n11205), .Z(n11096) );
  OR U15451 ( .A(n11206), .B(n11207), .Z(n11205) );
  OR U15452 ( .A(n11208), .B(n11209), .Z(n11204) );
  ANDN U15453 ( .B(n11210), .A(n11211), .Z(n11097) );
  IV U15454 ( .A(n11212), .Z(n11210) );
  XNOR U15455 ( .A(n11177), .B(n11176), .Z(N29237) );
  XOR U15456 ( .A(n11196), .B(n11195), .Z(n11176) );
  XNOR U15457 ( .A(n11211), .B(n11212), .Z(n11195) );
  XNOR U15458 ( .A(n11206), .B(n11207), .Z(n11212) );
  XNOR U15459 ( .A(n11208), .B(n11209), .Z(n11207) );
  XNOR U15460 ( .A(y[2620]), .B(x[2620]), .Z(n11209) );
  XNOR U15461 ( .A(y[2621]), .B(x[2621]), .Z(n11208) );
  XNOR U15462 ( .A(y[2619]), .B(x[2619]), .Z(n11206) );
  XNOR U15463 ( .A(n11200), .B(n11201), .Z(n11211) );
  XNOR U15464 ( .A(y[2616]), .B(x[2616]), .Z(n11201) );
  XNOR U15465 ( .A(n11202), .B(n11203), .Z(n11200) );
  XNOR U15466 ( .A(y[2617]), .B(x[2617]), .Z(n11203) );
  XNOR U15467 ( .A(y[2618]), .B(x[2618]), .Z(n11202) );
  XNOR U15468 ( .A(n11193), .B(n11192), .Z(n11196) );
  XNOR U15469 ( .A(n11188), .B(n11189), .Z(n11192) );
  XNOR U15470 ( .A(y[2613]), .B(x[2613]), .Z(n11189) );
  XNOR U15471 ( .A(n11190), .B(n11191), .Z(n11188) );
  XNOR U15472 ( .A(y[2614]), .B(x[2614]), .Z(n11191) );
  XNOR U15473 ( .A(y[2615]), .B(x[2615]), .Z(n11190) );
  XNOR U15474 ( .A(n11182), .B(n11183), .Z(n11193) );
  XNOR U15475 ( .A(y[2610]), .B(x[2610]), .Z(n11183) );
  XNOR U15476 ( .A(n11184), .B(n11185), .Z(n11182) );
  XNOR U15477 ( .A(y[2611]), .B(x[2611]), .Z(n11185) );
  XNOR U15478 ( .A(y[2612]), .B(x[2612]), .Z(n11184) );
  XOR U15479 ( .A(n11158), .B(n11159), .Z(n11177) );
  XNOR U15480 ( .A(n11174), .B(n11175), .Z(n11159) );
  XNOR U15481 ( .A(n11169), .B(n11170), .Z(n11175) );
  XNOR U15482 ( .A(n11171), .B(n11172), .Z(n11170) );
  XNOR U15483 ( .A(y[2608]), .B(x[2608]), .Z(n11172) );
  XNOR U15484 ( .A(y[2609]), .B(x[2609]), .Z(n11171) );
  XNOR U15485 ( .A(y[2607]), .B(x[2607]), .Z(n11169) );
  XNOR U15486 ( .A(n11163), .B(n11164), .Z(n11174) );
  XNOR U15487 ( .A(y[2604]), .B(x[2604]), .Z(n11164) );
  XNOR U15488 ( .A(n11165), .B(n11166), .Z(n11163) );
  XNOR U15489 ( .A(y[2605]), .B(x[2605]), .Z(n11166) );
  XNOR U15490 ( .A(y[2606]), .B(x[2606]), .Z(n11165) );
  XOR U15491 ( .A(n11157), .B(n11156), .Z(n11158) );
  XNOR U15492 ( .A(n11152), .B(n11153), .Z(n11156) );
  XNOR U15493 ( .A(y[2601]), .B(x[2601]), .Z(n11153) );
  XNOR U15494 ( .A(n11154), .B(n11155), .Z(n11152) );
  XNOR U15495 ( .A(y[2602]), .B(x[2602]), .Z(n11155) );
  XNOR U15496 ( .A(y[2603]), .B(x[2603]), .Z(n11154) );
  XNOR U15497 ( .A(n11146), .B(n11147), .Z(n11157) );
  XNOR U15498 ( .A(y[2598]), .B(x[2598]), .Z(n11147) );
  XNOR U15499 ( .A(n11148), .B(n11149), .Z(n11146) );
  XNOR U15500 ( .A(y[2599]), .B(x[2599]), .Z(n11149) );
  XNOR U15501 ( .A(y[2600]), .B(x[2600]), .Z(n11148) );
  NAND U15502 ( .A(n11213), .B(n11214), .Z(N29229) );
  NANDN U15503 ( .A(n11215), .B(n11216), .Z(n11214) );
  OR U15504 ( .A(n11217), .B(n11218), .Z(n11216) );
  NAND U15505 ( .A(n11217), .B(n11218), .Z(n11213) );
  XOR U15506 ( .A(n11217), .B(n11219), .Z(N29228) );
  XNOR U15507 ( .A(n11215), .B(n11218), .Z(n11219) );
  AND U15508 ( .A(n11220), .B(n11221), .Z(n11218) );
  NANDN U15509 ( .A(n11222), .B(n11223), .Z(n11221) );
  NANDN U15510 ( .A(n11224), .B(n11225), .Z(n11223) );
  NANDN U15511 ( .A(n11225), .B(n11224), .Z(n11220) );
  NAND U15512 ( .A(n11226), .B(n11227), .Z(n11215) );
  NANDN U15513 ( .A(n11228), .B(n11229), .Z(n11227) );
  OR U15514 ( .A(n11230), .B(n11231), .Z(n11229) );
  NAND U15515 ( .A(n11231), .B(n11230), .Z(n11226) );
  AND U15516 ( .A(n11232), .B(n11233), .Z(n11217) );
  NANDN U15517 ( .A(n11234), .B(n11235), .Z(n11233) );
  NANDN U15518 ( .A(n11236), .B(n11237), .Z(n11235) );
  NANDN U15519 ( .A(n11237), .B(n11236), .Z(n11232) );
  XOR U15520 ( .A(n11231), .B(n11238), .Z(N29227) );
  XOR U15521 ( .A(n11228), .B(n11230), .Z(n11238) );
  XNOR U15522 ( .A(n11224), .B(n11239), .Z(n11230) );
  XNOR U15523 ( .A(n11222), .B(n11225), .Z(n11239) );
  NAND U15524 ( .A(n11240), .B(n11241), .Z(n11225) );
  NAND U15525 ( .A(n11242), .B(n11243), .Z(n11241) );
  OR U15526 ( .A(n11244), .B(n11245), .Z(n11242) );
  NANDN U15527 ( .A(n11246), .B(n11244), .Z(n11240) );
  IV U15528 ( .A(n11245), .Z(n11246) );
  NAND U15529 ( .A(n11247), .B(n11248), .Z(n11222) );
  NAND U15530 ( .A(n11249), .B(n11250), .Z(n11248) );
  NANDN U15531 ( .A(n11251), .B(n11252), .Z(n11249) );
  NANDN U15532 ( .A(n11252), .B(n11251), .Z(n11247) );
  AND U15533 ( .A(n11253), .B(n11254), .Z(n11224) );
  NAND U15534 ( .A(n11255), .B(n11256), .Z(n11254) );
  OR U15535 ( .A(n11257), .B(n11258), .Z(n11255) );
  NANDN U15536 ( .A(n11259), .B(n11257), .Z(n11253) );
  NAND U15537 ( .A(n11260), .B(n11261), .Z(n11228) );
  NANDN U15538 ( .A(n11262), .B(n11263), .Z(n11261) );
  OR U15539 ( .A(n11264), .B(n11265), .Z(n11263) );
  NANDN U15540 ( .A(n11266), .B(n11264), .Z(n11260) );
  IV U15541 ( .A(n11265), .Z(n11266) );
  XNOR U15542 ( .A(n11236), .B(n11267), .Z(n11231) );
  XNOR U15543 ( .A(n11234), .B(n11237), .Z(n11267) );
  NAND U15544 ( .A(n11268), .B(n11269), .Z(n11237) );
  NAND U15545 ( .A(n11270), .B(n11271), .Z(n11269) );
  OR U15546 ( .A(n11272), .B(n11273), .Z(n11270) );
  NANDN U15547 ( .A(n11274), .B(n11272), .Z(n11268) );
  IV U15548 ( .A(n11273), .Z(n11274) );
  NAND U15549 ( .A(n11275), .B(n11276), .Z(n11234) );
  NAND U15550 ( .A(n11277), .B(n11278), .Z(n11276) );
  NANDN U15551 ( .A(n11279), .B(n11280), .Z(n11277) );
  NANDN U15552 ( .A(n11280), .B(n11279), .Z(n11275) );
  AND U15553 ( .A(n11281), .B(n11282), .Z(n11236) );
  NAND U15554 ( .A(n11283), .B(n11284), .Z(n11282) );
  OR U15555 ( .A(n11285), .B(n11286), .Z(n11283) );
  NANDN U15556 ( .A(n11287), .B(n11285), .Z(n11281) );
  XNOR U15557 ( .A(n11262), .B(n11288), .Z(N29226) );
  XOR U15558 ( .A(n11264), .B(n11265), .Z(n11288) );
  XNOR U15559 ( .A(n11278), .B(n11289), .Z(n11265) );
  XOR U15560 ( .A(n11279), .B(n11280), .Z(n11289) );
  XOR U15561 ( .A(n11285), .B(n11290), .Z(n11280) );
  XOR U15562 ( .A(n11284), .B(n11287), .Z(n11290) );
  IV U15563 ( .A(n11286), .Z(n11287) );
  NAND U15564 ( .A(n11291), .B(n11292), .Z(n11286) );
  OR U15565 ( .A(n11293), .B(n11294), .Z(n11292) );
  OR U15566 ( .A(n11295), .B(n11296), .Z(n11291) );
  NAND U15567 ( .A(n11297), .B(n11298), .Z(n11284) );
  OR U15568 ( .A(n11299), .B(n11300), .Z(n11298) );
  OR U15569 ( .A(n11301), .B(n11302), .Z(n11297) );
  NOR U15570 ( .A(n11303), .B(n11304), .Z(n11285) );
  ANDN U15571 ( .B(n11305), .A(n11306), .Z(n11279) );
  XNOR U15572 ( .A(n11272), .B(n11307), .Z(n11278) );
  XNOR U15573 ( .A(n11271), .B(n11273), .Z(n11307) );
  NAND U15574 ( .A(n11308), .B(n11309), .Z(n11273) );
  OR U15575 ( .A(n11310), .B(n11311), .Z(n11309) );
  OR U15576 ( .A(n11312), .B(n11313), .Z(n11308) );
  NAND U15577 ( .A(n11314), .B(n11315), .Z(n11271) );
  OR U15578 ( .A(n11316), .B(n11317), .Z(n11315) );
  OR U15579 ( .A(n11318), .B(n11319), .Z(n11314) );
  ANDN U15580 ( .B(n11320), .A(n11321), .Z(n11272) );
  IV U15581 ( .A(n11322), .Z(n11320) );
  ANDN U15582 ( .B(n11323), .A(n11324), .Z(n11264) );
  XOR U15583 ( .A(n11250), .B(n11325), .Z(n11262) );
  XOR U15584 ( .A(n11251), .B(n11252), .Z(n11325) );
  XOR U15585 ( .A(n11257), .B(n11326), .Z(n11252) );
  XOR U15586 ( .A(n11256), .B(n11259), .Z(n11326) );
  IV U15587 ( .A(n11258), .Z(n11259) );
  NAND U15588 ( .A(n11327), .B(n11328), .Z(n11258) );
  OR U15589 ( .A(n11329), .B(n11330), .Z(n11328) );
  OR U15590 ( .A(n11331), .B(n11332), .Z(n11327) );
  NAND U15591 ( .A(n11333), .B(n11334), .Z(n11256) );
  OR U15592 ( .A(n11335), .B(n11336), .Z(n11334) );
  OR U15593 ( .A(n11337), .B(n11338), .Z(n11333) );
  NOR U15594 ( .A(n11339), .B(n11340), .Z(n11257) );
  ANDN U15595 ( .B(n11341), .A(n11342), .Z(n11251) );
  IV U15596 ( .A(n11343), .Z(n11341) );
  XNOR U15597 ( .A(n11244), .B(n11344), .Z(n11250) );
  XNOR U15598 ( .A(n11243), .B(n11245), .Z(n11344) );
  NAND U15599 ( .A(n11345), .B(n11346), .Z(n11245) );
  OR U15600 ( .A(n11347), .B(n11348), .Z(n11346) );
  OR U15601 ( .A(n11349), .B(n11350), .Z(n11345) );
  NAND U15602 ( .A(n11351), .B(n11352), .Z(n11243) );
  OR U15603 ( .A(n11353), .B(n11354), .Z(n11352) );
  OR U15604 ( .A(n11355), .B(n11356), .Z(n11351) );
  ANDN U15605 ( .B(n11357), .A(n11358), .Z(n11244) );
  IV U15606 ( .A(n11359), .Z(n11357) );
  XNOR U15607 ( .A(n11324), .B(n11323), .Z(N29225) );
  XOR U15608 ( .A(n11343), .B(n11342), .Z(n11323) );
  XNOR U15609 ( .A(n11358), .B(n11359), .Z(n11342) );
  XNOR U15610 ( .A(n11353), .B(n11354), .Z(n11359) );
  XNOR U15611 ( .A(n11355), .B(n11356), .Z(n11354) );
  XNOR U15612 ( .A(y[2596]), .B(x[2596]), .Z(n11356) );
  XNOR U15613 ( .A(y[2597]), .B(x[2597]), .Z(n11355) );
  XNOR U15614 ( .A(y[2595]), .B(x[2595]), .Z(n11353) );
  XNOR U15615 ( .A(n11347), .B(n11348), .Z(n11358) );
  XNOR U15616 ( .A(y[2592]), .B(x[2592]), .Z(n11348) );
  XNOR U15617 ( .A(n11349), .B(n11350), .Z(n11347) );
  XNOR U15618 ( .A(y[2593]), .B(x[2593]), .Z(n11350) );
  XNOR U15619 ( .A(y[2594]), .B(x[2594]), .Z(n11349) );
  XNOR U15620 ( .A(n11340), .B(n11339), .Z(n11343) );
  XNOR U15621 ( .A(n11335), .B(n11336), .Z(n11339) );
  XNOR U15622 ( .A(y[2589]), .B(x[2589]), .Z(n11336) );
  XNOR U15623 ( .A(n11337), .B(n11338), .Z(n11335) );
  XNOR U15624 ( .A(y[2590]), .B(x[2590]), .Z(n11338) );
  XNOR U15625 ( .A(y[2591]), .B(x[2591]), .Z(n11337) );
  XNOR U15626 ( .A(n11329), .B(n11330), .Z(n11340) );
  XNOR U15627 ( .A(y[2586]), .B(x[2586]), .Z(n11330) );
  XNOR U15628 ( .A(n11331), .B(n11332), .Z(n11329) );
  XNOR U15629 ( .A(y[2587]), .B(x[2587]), .Z(n11332) );
  XNOR U15630 ( .A(y[2588]), .B(x[2588]), .Z(n11331) );
  XOR U15631 ( .A(n11305), .B(n11306), .Z(n11324) );
  XNOR U15632 ( .A(n11321), .B(n11322), .Z(n11306) );
  XNOR U15633 ( .A(n11316), .B(n11317), .Z(n11322) );
  XNOR U15634 ( .A(n11318), .B(n11319), .Z(n11317) );
  XNOR U15635 ( .A(y[2584]), .B(x[2584]), .Z(n11319) );
  XNOR U15636 ( .A(y[2585]), .B(x[2585]), .Z(n11318) );
  XNOR U15637 ( .A(y[2583]), .B(x[2583]), .Z(n11316) );
  XNOR U15638 ( .A(n11310), .B(n11311), .Z(n11321) );
  XNOR U15639 ( .A(y[2580]), .B(x[2580]), .Z(n11311) );
  XNOR U15640 ( .A(n11312), .B(n11313), .Z(n11310) );
  XNOR U15641 ( .A(y[2581]), .B(x[2581]), .Z(n11313) );
  XNOR U15642 ( .A(y[2582]), .B(x[2582]), .Z(n11312) );
  XOR U15643 ( .A(n11304), .B(n11303), .Z(n11305) );
  XNOR U15644 ( .A(n11299), .B(n11300), .Z(n11303) );
  XNOR U15645 ( .A(y[2577]), .B(x[2577]), .Z(n11300) );
  XNOR U15646 ( .A(n11301), .B(n11302), .Z(n11299) );
  XNOR U15647 ( .A(y[2578]), .B(x[2578]), .Z(n11302) );
  XNOR U15648 ( .A(y[2579]), .B(x[2579]), .Z(n11301) );
  XNOR U15649 ( .A(n11293), .B(n11294), .Z(n11304) );
  XNOR U15650 ( .A(y[2574]), .B(x[2574]), .Z(n11294) );
  XNOR U15651 ( .A(n11295), .B(n11296), .Z(n11293) );
  XNOR U15652 ( .A(y[2575]), .B(x[2575]), .Z(n11296) );
  XNOR U15653 ( .A(y[2576]), .B(x[2576]), .Z(n11295) );
  NAND U15654 ( .A(n11360), .B(n11361), .Z(N29217) );
  NANDN U15655 ( .A(n11362), .B(n11363), .Z(n11361) );
  OR U15656 ( .A(n11364), .B(n11365), .Z(n11363) );
  NAND U15657 ( .A(n11364), .B(n11365), .Z(n11360) );
  XOR U15658 ( .A(n11364), .B(n11366), .Z(N29216) );
  XNOR U15659 ( .A(n11362), .B(n11365), .Z(n11366) );
  AND U15660 ( .A(n11367), .B(n11368), .Z(n11365) );
  NANDN U15661 ( .A(n11369), .B(n11370), .Z(n11368) );
  NANDN U15662 ( .A(n11371), .B(n11372), .Z(n11370) );
  NANDN U15663 ( .A(n11372), .B(n11371), .Z(n11367) );
  NAND U15664 ( .A(n11373), .B(n11374), .Z(n11362) );
  NANDN U15665 ( .A(n11375), .B(n11376), .Z(n11374) );
  OR U15666 ( .A(n11377), .B(n11378), .Z(n11376) );
  NAND U15667 ( .A(n11378), .B(n11377), .Z(n11373) );
  AND U15668 ( .A(n11379), .B(n11380), .Z(n11364) );
  NANDN U15669 ( .A(n11381), .B(n11382), .Z(n11380) );
  NANDN U15670 ( .A(n11383), .B(n11384), .Z(n11382) );
  NANDN U15671 ( .A(n11384), .B(n11383), .Z(n11379) );
  XOR U15672 ( .A(n11378), .B(n11385), .Z(N29215) );
  XOR U15673 ( .A(n11375), .B(n11377), .Z(n11385) );
  XNOR U15674 ( .A(n11371), .B(n11386), .Z(n11377) );
  XNOR U15675 ( .A(n11369), .B(n11372), .Z(n11386) );
  NAND U15676 ( .A(n11387), .B(n11388), .Z(n11372) );
  NAND U15677 ( .A(n11389), .B(n11390), .Z(n11388) );
  OR U15678 ( .A(n11391), .B(n11392), .Z(n11389) );
  NANDN U15679 ( .A(n11393), .B(n11391), .Z(n11387) );
  IV U15680 ( .A(n11392), .Z(n11393) );
  NAND U15681 ( .A(n11394), .B(n11395), .Z(n11369) );
  NAND U15682 ( .A(n11396), .B(n11397), .Z(n11395) );
  NANDN U15683 ( .A(n11398), .B(n11399), .Z(n11396) );
  NANDN U15684 ( .A(n11399), .B(n11398), .Z(n11394) );
  AND U15685 ( .A(n11400), .B(n11401), .Z(n11371) );
  NAND U15686 ( .A(n11402), .B(n11403), .Z(n11401) );
  OR U15687 ( .A(n11404), .B(n11405), .Z(n11402) );
  NANDN U15688 ( .A(n11406), .B(n11404), .Z(n11400) );
  NAND U15689 ( .A(n11407), .B(n11408), .Z(n11375) );
  NANDN U15690 ( .A(n11409), .B(n11410), .Z(n11408) );
  OR U15691 ( .A(n11411), .B(n11412), .Z(n11410) );
  NANDN U15692 ( .A(n11413), .B(n11411), .Z(n11407) );
  IV U15693 ( .A(n11412), .Z(n11413) );
  XNOR U15694 ( .A(n11383), .B(n11414), .Z(n11378) );
  XNOR U15695 ( .A(n11381), .B(n11384), .Z(n11414) );
  NAND U15696 ( .A(n11415), .B(n11416), .Z(n11384) );
  NAND U15697 ( .A(n11417), .B(n11418), .Z(n11416) );
  OR U15698 ( .A(n11419), .B(n11420), .Z(n11417) );
  NANDN U15699 ( .A(n11421), .B(n11419), .Z(n11415) );
  IV U15700 ( .A(n11420), .Z(n11421) );
  NAND U15701 ( .A(n11422), .B(n11423), .Z(n11381) );
  NAND U15702 ( .A(n11424), .B(n11425), .Z(n11423) );
  NANDN U15703 ( .A(n11426), .B(n11427), .Z(n11424) );
  NANDN U15704 ( .A(n11427), .B(n11426), .Z(n11422) );
  AND U15705 ( .A(n11428), .B(n11429), .Z(n11383) );
  NAND U15706 ( .A(n11430), .B(n11431), .Z(n11429) );
  OR U15707 ( .A(n11432), .B(n11433), .Z(n11430) );
  NANDN U15708 ( .A(n11434), .B(n11432), .Z(n11428) );
  XNOR U15709 ( .A(n11409), .B(n11435), .Z(N29214) );
  XOR U15710 ( .A(n11411), .B(n11412), .Z(n11435) );
  XNOR U15711 ( .A(n11425), .B(n11436), .Z(n11412) );
  XOR U15712 ( .A(n11426), .B(n11427), .Z(n11436) );
  XOR U15713 ( .A(n11432), .B(n11437), .Z(n11427) );
  XOR U15714 ( .A(n11431), .B(n11434), .Z(n11437) );
  IV U15715 ( .A(n11433), .Z(n11434) );
  NAND U15716 ( .A(n11438), .B(n11439), .Z(n11433) );
  OR U15717 ( .A(n11440), .B(n11441), .Z(n11439) );
  OR U15718 ( .A(n11442), .B(n11443), .Z(n11438) );
  NAND U15719 ( .A(n11444), .B(n11445), .Z(n11431) );
  OR U15720 ( .A(n11446), .B(n11447), .Z(n11445) );
  OR U15721 ( .A(n11448), .B(n11449), .Z(n11444) );
  NOR U15722 ( .A(n11450), .B(n11451), .Z(n11432) );
  ANDN U15723 ( .B(n11452), .A(n11453), .Z(n11426) );
  XNOR U15724 ( .A(n11419), .B(n11454), .Z(n11425) );
  XNOR U15725 ( .A(n11418), .B(n11420), .Z(n11454) );
  NAND U15726 ( .A(n11455), .B(n11456), .Z(n11420) );
  OR U15727 ( .A(n11457), .B(n11458), .Z(n11456) );
  OR U15728 ( .A(n11459), .B(n11460), .Z(n11455) );
  NAND U15729 ( .A(n11461), .B(n11462), .Z(n11418) );
  OR U15730 ( .A(n11463), .B(n11464), .Z(n11462) );
  OR U15731 ( .A(n11465), .B(n11466), .Z(n11461) );
  ANDN U15732 ( .B(n11467), .A(n11468), .Z(n11419) );
  IV U15733 ( .A(n11469), .Z(n11467) );
  ANDN U15734 ( .B(n11470), .A(n11471), .Z(n11411) );
  XOR U15735 ( .A(n11397), .B(n11472), .Z(n11409) );
  XOR U15736 ( .A(n11398), .B(n11399), .Z(n11472) );
  XOR U15737 ( .A(n11404), .B(n11473), .Z(n11399) );
  XOR U15738 ( .A(n11403), .B(n11406), .Z(n11473) );
  IV U15739 ( .A(n11405), .Z(n11406) );
  NAND U15740 ( .A(n11474), .B(n11475), .Z(n11405) );
  OR U15741 ( .A(n11476), .B(n11477), .Z(n11475) );
  OR U15742 ( .A(n11478), .B(n11479), .Z(n11474) );
  NAND U15743 ( .A(n11480), .B(n11481), .Z(n11403) );
  OR U15744 ( .A(n11482), .B(n11483), .Z(n11481) );
  OR U15745 ( .A(n11484), .B(n11485), .Z(n11480) );
  NOR U15746 ( .A(n11486), .B(n11487), .Z(n11404) );
  ANDN U15747 ( .B(n11488), .A(n11489), .Z(n11398) );
  IV U15748 ( .A(n11490), .Z(n11488) );
  XNOR U15749 ( .A(n11391), .B(n11491), .Z(n11397) );
  XNOR U15750 ( .A(n11390), .B(n11392), .Z(n11491) );
  NAND U15751 ( .A(n11492), .B(n11493), .Z(n11392) );
  OR U15752 ( .A(n11494), .B(n11495), .Z(n11493) );
  OR U15753 ( .A(n11496), .B(n11497), .Z(n11492) );
  NAND U15754 ( .A(n11498), .B(n11499), .Z(n11390) );
  OR U15755 ( .A(n11500), .B(n11501), .Z(n11499) );
  OR U15756 ( .A(n11502), .B(n11503), .Z(n11498) );
  ANDN U15757 ( .B(n11504), .A(n11505), .Z(n11391) );
  IV U15758 ( .A(n11506), .Z(n11504) );
  XNOR U15759 ( .A(n11471), .B(n11470), .Z(N29213) );
  XOR U15760 ( .A(n11490), .B(n11489), .Z(n11470) );
  XNOR U15761 ( .A(n11505), .B(n11506), .Z(n11489) );
  XNOR U15762 ( .A(n11500), .B(n11501), .Z(n11506) );
  XNOR U15763 ( .A(n11502), .B(n11503), .Z(n11501) );
  XNOR U15764 ( .A(y[2572]), .B(x[2572]), .Z(n11503) );
  XNOR U15765 ( .A(y[2573]), .B(x[2573]), .Z(n11502) );
  XNOR U15766 ( .A(y[2571]), .B(x[2571]), .Z(n11500) );
  XNOR U15767 ( .A(n11494), .B(n11495), .Z(n11505) );
  XNOR U15768 ( .A(y[2568]), .B(x[2568]), .Z(n11495) );
  XNOR U15769 ( .A(n11496), .B(n11497), .Z(n11494) );
  XNOR U15770 ( .A(y[2569]), .B(x[2569]), .Z(n11497) );
  XNOR U15771 ( .A(y[2570]), .B(x[2570]), .Z(n11496) );
  XNOR U15772 ( .A(n11487), .B(n11486), .Z(n11490) );
  XNOR U15773 ( .A(n11482), .B(n11483), .Z(n11486) );
  XNOR U15774 ( .A(y[2565]), .B(x[2565]), .Z(n11483) );
  XNOR U15775 ( .A(n11484), .B(n11485), .Z(n11482) );
  XNOR U15776 ( .A(y[2566]), .B(x[2566]), .Z(n11485) );
  XNOR U15777 ( .A(y[2567]), .B(x[2567]), .Z(n11484) );
  XNOR U15778 ( .A(n11476), .B(n11477), .Z(n11487) );
  XNOR U15779 ( .A(y[2562]), .B(x[2562]), .Z(n11477) );
  XNOR U15780 ( .A(n11478), .B(n11479), .Z(n11476) );
  XNOR U15781 ( .A(y[2563]), .B(x[2563]), .Z(n11479) );
  XNOR U15782 ( .A(y[2564]), .B(x[2564]), .Z(n11478) );
  XOR U15783 ( .A(n11452), .B(n11453), .Z(n11471) );
  XNOR U15784 ( .A(n11468), .B(n11469), .Z(n11453) );
  XNOR U15785 ( .A(n11463), .B(n11464), .Z(n11469) );
  XNOR U15786 ( .A(n11465), .B(n11466), .Z(n11464) );
  XNOR U15787 ( .A(y[2560]), .B(x[2560]), .Z(n11466) );
  XNOR U15788 ( .A(y[2561]), .B(x[2561]), .Z(n11465) );
  XNOR U15789 ( .A(y[2559]), .B(x[2559]), .Z(n11463) );
  XNOR U15790 ( .A(n11457), .B(n11458), .Z(n11468) );
  XNOR U15791 ( .A(y[2556]), .B(x[2556]), .Z(n11458) );
  XNOR U15792 ( .A(n11459), .B(n11460), .Z(n11457) );
  XNOR U15793 ( .A(y[2557]), .B(x[2557]), .Z(n11460) );
  XNOR U15794 ( .A(y[2558]), .B(x[2558]), .Z(n11459) );
  XOR U15795 ( .A(n11451), .B(n11450), .Z(n11452) );
  XNOR U15796 ( .A(n11446), .B(n11447), .Z(n11450) );
  XNOR U15797 ( .A(y[2553]), .B(x[2553]), .Z(n11447) );
  XNOR U15798 ( .A(n11448), .B(n11449), .Z(n11446) );
  XNOR U15799 ( .A(y[2554]), .B(x[2554]), .Z(n11449) );
  XNOR U15800 ( .A(y[2555]), .B(x[2555]), .Z(n11448) );
  XNOR U15801 ( .A(n11440), .B(n11441), .Z(n11451) );
  XNOR U15802 ( .A(y[2550]), .B(x[2550]), .Z(n11441) );
  XNOR U15803 ( .A(n11442), .B(n11443), .Z(n11440) );
  XNOR U15804 ( .A(y[2551]), .B(x[2551]), .Z(n11443) );
  XNOR U15805 ( .A(y[2552]), .B(x[2552]), .Z(n11442) );
  NAND U15806 ( .A(n11507), .B(n11508), .Z(N29205) );
  NANDN U15807 ( .A(n11509), .B(n11510), .Z(n11508) );
  OR U15808 ( .A(n11511), .B(n11512), .Z(n11510) );
  NAND U15809 ( .A(n11511), .B(n11512), .Z(n11507) );
  XOR U15810 ( .A(n11511), .B(n11513), .Z(N29204) );
  XNOR U15811 ( .A(n11509), .B(n11512), .Z(n11513) );
  AND U15812 ( .A(n11514), .B(n11515), .Z(n11512) );
  NANDN U15813 ( .A(n11516), .B(n11517), .Z(n11515) );
  NANDN U15814 ( .A(n11518), .B(n11519), .Z(n11517) );
  NANDN U15815 ( .A(n11519), .B(n11518), .Z(n11514) );
  NAND U15816 ( .A(n11520), .B(n11521), .Z(n11509) );
  NANDN U15817 ( .A(n11522), .B(n11523), .Z(n11521) );
  OR U15818 ( .A(n11524), .B(n11525), .Z(n11523) );
  NAND U15819 ( .A(n11525), .B(n11524), .Z(n11520) );
  AND U15820 ( .A(n11526), .B(n11527), .Z(n11511) );
  NANDN U15821 ( .A(n11528), .B(n11529), .Z(n11527) );
  NANDN U15822 ( .A(n11530), .B(n11531), .Z(n11529) );
  NANDN U15823 ( .A(n11531), .B(n11530), .Z(n11526) );
  XOR U15824 ( .A(n11525), .B(n11532), .Z(N29203) );
  XOR U15825 ( .A(n11522), .B(n11524), .Z(n11532) );
  XNOR U15826 ( .A(n11518), .B(n11533), .Z(n11524) );
  XNOR U15827 ( .A(n11516), .B(n11519), .Z(n11533) );
  NAND U15828 ( .A(n11534), .B(n11535), .Z(n11519) );
  NAND U15829 ( .A(n11536), .B(n11537), .Z(n11535) );
  OR U15830 ( .A(n11538), .B(n11539), .Z(n11536) );
  NANDN U15831 ( .A(n11540), .B(n11538), .Z(n11534) );
  IV U15832 ( .A(n11539), .Z(n11540) );
  NAND U15833 ( .A(n11541), .B(n11542), .Z(n11516) );
  NAND U15834 ( .A(n11543), .B(n11544), .Z(n11542) );
  NANDN U15835 ( .A(n11545), .B(n11546), .Z(n11543) );
  NANDN U15836 ( .A(n11546), .B(n11545), .Z(n11541) );
  AND U15837 ( .A(n11547), .B(n11548), .Z(n11518) );
  NAND U15838 ( .A(n11549), .B(n11550), .Z(n11548) );
  OR U15839 ( .A(n11551), .B(n11552), .Z(n11549) );
  NANDN U15840 ( .A(n11553), .B(n11551), .Z(n11547) );
  NAND U15841 ( .A(n11554), .B(n11555), .Z(n11522) );
  NANDN U15842 ( .A(n11556), .B(n11557), .Z(n11555) );
  OR U15843 ( .A(n11558), .B(n11559), .Z(n11557) );
  NANDN U15844 ( .A(n11560), .B(n11558), .Z(n11554) );
  IV U15845 ( .A(n11559), .Z(n11560) );
  XNOR U15846 ( .A(n11530), .B(n11561), .Z(n11525) );
  XNOR U15847 ( .A(n11528), .B(n11531), .Z(n11561) );
  NAND U15848 ( .A(n11562), .B(n11563), .Z(n11531) );
  NAND U15849 ( .A(n11564), .B(n11565), .Z(n11563) );
  OR U15850 ( .A(n11566), .B(n11567), .Z(n11564) );
  NANDN U15851 ( .A(n11568), .B(n11566), .Z(n11562) );
  IV U15852 ( .A(n11567), .Z(n11568) );
  NAND U15853 ( .A(n11569), .B(n11570), .Z(n11528) );
  NAND U15854 ( .A(n11571), .B(n11572), .Z(n11570) );
  NANDN U15855 ( .A(n11573), .B(n11574), .Z(n11571) );
  NANDN U15856 ( .A(n11574), .B(n11573), .Z(n11569) );
  AND U15857 ( .A(n11575), .B(n11576), .Z(n11530) );
  NAND U15858 ( .A(n11577), .B(n11578), .Z(n11576) );
  OR U15859 ( .A(n11579), .B(n11580), .Z(n11577) );
  NANDN U15860 ( .A(n11581), .B(n11579), .Z(n11575) );
  XNOR U15861 ( .A(n11556), .B(n11582), .Z(N29202) );
  XOR U15862 ( .A(n11558), .B(n11559), .Z(n11582) );
  XNOR U15863 ( .A(n11572), .B(n11583), .Z(n11559) );
  XOR U15864 ( .A(n11573), .B(n11574), .Z(n11583) );
  XOR U15865 ( .A(n11579), .B(n11584), .Z(n11574) );
  XOR U15866 ( .A(n11578), .B(n11581), .Z(n11584) );
  IV U15867 ( .A(n11580), .Z(n11581) );
  NAND U15868 ( .A(n11585), .B(n11586), .Z(n11580) );
  OR U15869 ( .A(n11587), .B(n11588), .Z(n11586) );
  OR U15870 ( .A(n11589), .B(n11590), .Z(n11585) );
  NAND U15871 ( .A(n11591), .B(n11592), .Z(n11578) );
  OR U15872 ( .A(n11593), .B(n11594), .Z(n11592) );
  OR U15873 ( .A(n11595), .B(n11596), .Z(n11591) );
  NOR U15874 ( .A(n11597), .B(n11598), .Z(n11579) );
  ANDN U15875 ( .B(n11599), .A(n11600), .Z(n11573) );
  XNOR U15876 ( .A(n11566), .B(n11601), .Z(n11572) );
  XNOR U15877 ( .A(n11565), .B(n11567), .Z(n11601) );
  NAND U15878 ( .A(n11602), .B(n11603), .Z(n11567) );
  OR U15879 ( .A(n11604), .B(n11605), .Z(n11603) );
  OR U15880 ( .A(n11606), .B(n11607), .Z(n11602) );
  NAND U15881 ( .A(n11608), .B(n11609), .Z(n11565) );
  OR U15882 ( .A(n11610), .B(n11611), .Z(n11609) );
  OR U15883 ( .A(n11612), .B(n11613), .Z(n11608) );
  ANDN U15884 ( .B(n11614), .A(n11615), .Z(n11566) );
  IV U15885 ( .A(n11616), .Z(n11614) );
  ANDN U15886 ( .B(n11617), .A(n11618), .Z(n11558) );
  XOR U15887 ( .A(n11544), .B(n11619), .Z(n11556) );
  XOR U15888 ( .A(n11545), .B(n11546), .Z(n11619) );
  XOR U15889 ( .A(n11551), .B(n11620), .Z(n11546) );
  XOR U15890 ( .A(n11550), .B(n11553), .Z(n11620) );
  IV U15891 ( .A(n11552), .Z(n11553) );
  NAND U15892 ( .A(n11621), .B(n11622), .Z(n11552) );
  OR U15893 ( .A(n11623), .B(n11624), .Z(n11622) );
  OR U15894 ( .A(n11625), .B(n11626), .Z(n11621) );
  NAND U15895 ( .A(n11627), .B(n11628), .Z(n11550) );
  OR U15896 ( .A(n11629), .B(n11630), .Z(n11628) );
  OR U15897 ( .A(n11631), .B(n11632), .Z(n11627) );
  NOR U15898 ( .A(n11633), .B(n11634), .Z(n11551) );
  ANDN U15899 ( .B(n11635), .A(n11636), .Z(n11545) );
  IV U15900 ( .A(n11637), .Z(n11635) );
  XNOR U15901 ( .A(n11538), .B(n11638), .Z(n11544) );
  XNOR U15902 ( .A(n11537), .B(n11539), .Z(n11638) );
  NAND U15903 ( .A(n11639), .B(n11640), .Z(n11539) );
  OR U15904 ( .A(n11641), .B(n11642), .Z(n11640) );
  OR U15905 ( .A(n11643), .B(n11644), .Z(n11639) );
  NAND U15906 ( .A(n11645), .B(n11646), .Z(n11537) );
  OR U15907 ( .A(n11647), .B(n11648), .Z(n11646) );
  OR U15908 ( .A(n11649), .B(n11650), .Z(n11645) );
  ANDN U15909 ( .B(n11651), .A(n11652), .Z(n11538) );
  IV U15910 ( .A(n11653), .Z(n11651) );
  XNOR U15911 ( .A(n11618), .B(n11617), .Z(N29201) );
  XOR U15912 ( .A(n11637), .B(n11636), .Z(n11617) );
  XNOR U15913 ( .A(n11652), .B(n11653), .Z(n11636) );
  XNOR U15914 ( .A(n11647), .B(n11648), .Z(n11653) );
  XNOR U15915 ( .A(n11649), .B(n11650), .Z(n11648) );
  XNOR U15916 ( .A(y[2548]), .B(x[2548]), .Z(n11650) );
  XNOR U15917 ( .A(y[2549]), .B(x[2549]), .Z(n11649) );
  XNOR U15918 ( .A(y[2547]), .B(x[2547]), .Z(n11647) );
  XNOR U15919 ( .A(n11641), .B(n11642), .Z(n11652) );
  XNOR U15920 ( .A(y[2544]), .B(x[2544]), .Z(n11642) );
  XNOR U15921 ( .A(n11643), .B(n11644), .Z(n11641) );
  XNOR U15922 ( .A(y[2545]), .B(x[2545]), .Z(n11644) );
  XNOR U15923 ( .A(y[2546]), .B(x[2546]), .Z(n11643) );
  XNOR U15924 ( .A(n11634), .B(n11633), .Z(n11637) );
  XNOR U15925 ( .A(n11629), .B(n11630), .Z(n11633) );
  XNOR U15926 ( .A(y[2541]), .B(x[2541]), .Z(n11630) );
  XNOR U15927 ( .A(n11631), .B(n11632), .Z(n11629) );
  XNOR U15928 ( .A(y[2542]), .B(x[2542]), .Z(n11632) );
  XNOR U15929 ( .A(y[2543]), .B(x[2543]), .Z(n11631) );
  XNOR U15930 ( .A(n11623), .B(n11624), .Z(n11634) );
  XNOR U15931 ( .A(y[2538]), .B(x[2538]), .Z(n11624) );
  XNOR U15932 ( .A(n11625), .B(n11626), .Z(n11623) );
  XNOR U15933 ( .A(y[2539]), .B(x[2539]), .Z(n11626) );
  XNOR U15934 ( .A(y[2540]), .B(x[2540]), .Z(n11625) );
  XOR U15935 ( .A(n11599), .B(n11600), .Z(n11618) );
  XNOR U15936 ( .A(n11615), .B(n11616), .Z(n11600) );
  XNOR U15937 ( .A(n11610), .B(n11611), .Z(n11616) );
  XNOR U15938 ( .A(n11612), .B(n11613), .Z(n11611) );
  XNOR U15939 ( .A(y[2536]), .B(x[2536]), .Z(n11613) );
  XNOR U15940 ( .A(y[2537]), .B(x[2537]), .Z(n11612) );
  XNOR U15941 ( .A(y[2535]), .B(x[2535]), .Z(n11610) );
  XNOR U15942 ( .A(n11604), .B(n11605), .Z(n11615) );
  XNOR U15943 ( .A(y[2532]), .B(x[2532]), .Z(n11605) );
  XNOR U15944 ( .A(n11606), .B(n11607), .Z(n11604) );
  XNOR U15945 ( .A(y[2533]), .B(x[2533]), .Z(n11607) );
  XNOR U15946 ( .A(y[2534]), .B(x[2534]), .Z(n11606) );
  XOR U15947 ( .A(n11598), .B(n11597), .Z(n11599) );
  XNOR U15948 ( .A(n11593), .B(n11594), .Z(n11597) );
  XNOR U15949 ( .A(y[2529]), .B(x[2529]), .Z(n11594) );
  XNOR U15950 ( .A(n11595), .B(n11596), .Z(n11593) );
  XNOR U15951 ( .A(y[2530]), .B(x[2530]), .Z(n11596) );
  XNOR U15952 ( .A(y[2531]), .B(x[2531]), .Z(n11595) );
  XNOR U15953 ( .A(n11587), .B(n11588), .Z(n11598) );
  XNOR U15954 ( .A(y[2526]), .B(x[2526]), .Z(n11588) );
  XNOR U15955 ( .A(n11589), .B(n11590), .Z(n11587) );
  XNOR U15956 ( .A(y[2527]), .B(x[2527]), .Z(n11590) );
  XNOR U15957 ( .A(y[2528]), .B(x[2528]), .Z(n11589) );
  NAND U15958 ( .A(n11654), .B(n11655), .Z(N29193) );
  NANDN U15959 ( .A(n11656), .B(n11657), .Z(n11655) );
  OR U15960 ( .A(n11658), .B(n11659), .Z(n11657) );
  NAND U15961 ( .A(n11658), .B(n11659), .Z(n11654) );
  XOR U15962 ( .A(n11658), .B(n11660), .Z(N29192) );
  XNOR U15963 ( .A(n11656), .B(n11659), .Z(n11660) );
  AND U15964 ( .A(n11661), .B(n11662), .Z(n11659) );
  NANDN U15965 ( .A(n11663), .B(n11664), .Z(n11662) );
  NANDN U15966 ( .A(n11665), .B(n11666), .Z(n11664) );
  NANDN U15967 ( .A(n11666), .B(n11665), .Z(n11661) );
  NAND U15968 ( .A(n11667), .B(n11668), .Z(n11656) );
  NANDN U15969 ( .A(n11669), .B(n11670), .Z(n11668) );
  OR U15970 ( .A(n11671), .B(n11672), .Z(n11670) );
  NAND U15971 ( .A(n11672), .B(n11671), .Z(n11667) );
  AND U15972 ( .A(n11673), .B(n11674), .Z(n11658) );
  NANDN U15973 ( .A(n11675), .B(n11676), .Z(n11674) );
  NANDN U15974 ( .A(n11677), .B(n11678), .Z(n11676) );
  NANDN U15975 ( .A(n11678), .B(n11677), .Z(n11673) );
  XOR U15976 ( .A(n11672), .B(n11679), .Z(N29191) );
  XOR U15977 ( .A(n11669), .B(n11671), .Z(n11679) );
  XNOR U15978 ( .A(n11665), .B(n11680), .Z(n11671) );
  XNOR U15979 ( .A(n11663), .B(n11666), .Z(n11680) );
  NAND U15980 ( .A(n11681), .B(n11682), .Z(n11666) );
  NAND U15981 ( .A(n11683), .B(n11684), .Z(n11682) );
  OR U15982 ( .A(n11685), .B(n11686), .Z(n11683) );
  NANDN U15983 ( .A(n11687), .B(n11685), .Z(n11681) );
  IV U15984 ( .A(n11686), .Z(n11687) );
  NAND U15985 ( .A(n11688), .B(n11689), .Z(n11663) );
  NAND U15986 ( .A(n11690), .B(n11691), .Z(n11689) );
  NANDN U15987 ( .A(n11692), .B(n11693), .Z(n11690) );
  NANDN U15988 ( .A(n11693), .B(n11692), .Z(n11688) );
  AND U15989 ( .A(n11694), .B(n11695), .Z(n11665) );
  NAND U15990 ( .A(n11696), .B(n11697), .Z(n11695) );
  OR U15991 ( .A(n11698), .B(n11699), .Z(n11696) );
  NANDN U15992 ( .A(n11700), .B(n11698), .Z(n11694) );
  NAND U15993 ( .A(n11701), .B(n11702), .Z(n11669) );
  NANDN U15994 ( .A(n11703), .B(n11704), .Z(n11702) );
  OR U15995 ( .A(n11705), .B(n11706), .Z(n11704) );
  NANDN U15996 ( .A(n11707), .B(n11705), .Z(n11701) );
  IV U15997 ( .A(n11706), .Z(n11707) );
  XNOR U15998 ( .A(n11677), .B(n11708), .Z(n11672) );
  XNOR U15999 ( .A(n11675), .B(n11678), .Z(n11708) );
  NAND U16000 ( .A(n11709), .B(n11710), .Z(n11678) );
  NAND U16001 ( .A(n11711), .B(n11712), .Z(n11710) );
  OR U16002 ( .A(n11713), .B(n11714), .Z(n11711) );
  NANDN U16003 ( .A(n11715), .B(n11713), .Z(n11709) );
  IV U16004 ( .A(n11714), .Z(n11715) );
  NAND U16005 ( .A(n11716), .B(n11717), .Z(n11675) );
  NAND U16006 ( .A(n11718), .B(n11719), .Z(n11717) );
  NANDN U16007 ( .A(n11720), .B(n11721), .Z(n11718) );
  NANDN U16008 ( .A(n11721), .B(n11720), .Z(n11716) );
  AND U16009 ( .A(n11722), .B(n11723), .Z(n11677) );
  NAND U16010 ( .A(n11724), .B(n11725), .Z(n11723) );
  OR U16011 ( .A(n11726), .B(n11727), .Z(n11724) );
  NANDN U16012 ( .A(n11728), .B(n11726), .Z(n11722) );
  XNOR U16013 ( .A(n11703), .B(n11729), .Z(N29190) );
  XOR U16014 ( .A(n11705), .B(n11706), .Z(n11729) );
  XNOR U16015 ( .A(n11719), .B(n11730), .Z(n11706) );
  XOR U16016 ( .A(n11720), .B(n11721), .Z(n11730) );
  XOR U16017 ( .A(n11726), .B(n11731), .Z(n11721) );
  XOR U16018 ( .A(n11725), .B(n11728), .Z(n11731) );
  IV U16019 ( .A(n11727), .Z(n11728) );
  NAND U16020 ( .A(n11732), .B(n11733), .Z(n11727) );
  OR U16021 ( .A(n11734), .B(n11735), .Z(n11733) );
  OR U16022 ( .A(n11736), .B(n11737), .Z(n11732) );
  NAND U16023 ( .A(n11738), .B(n11739), .Z(n11725) );
  OR U16024 ( .A(n11740), .B(n11741), .Z(n11739) );
  OR U16025 ( .A(n11742), .B(n11743), .Z(n11738) );
  NOR U16026 ( .A(n11744), .B(n11745), .Z(n11726) );
  ANDN U16027 ( .B(n11746), .A(n11747), .Z(n11720) );
  XNOR U16028 ( .A(n11713), .B(n11748), .Z(n11719) );
  XNOR U16029 ( .A(n11712), .B(n11714), .Z(n11748) );
  NAND U16030 ( .A(n11749), .B(n11750), .Z(n11714) );
  OR U16031 ( .A(n11751), .B(n11752), .Z(n11750) );
  OR U16032 ( .A(n11753), .B(n11754), .Z(n11749) );
  NAND U16033 ( .A(n11755), .B(n11756), .Z(n11712) );
  OR U16034 ( .A(n11757), .B(n11758), .Z(n11756) );
  OR U16035 ( .A(n11759), .B(n11760), .Z(n11755) );
  ANDN U16036 ( .B(n11761), .A(n11762), .Z(n11713) );
  IV U16037 ( .A(n11763), .Z(n11761) );
  ANDN U16038 ( .B(n11764), .A(n11765), .Z(n11705) );
  XOR U16039 ( .A(n11691), .B(n11766), .Z(n11703) );
  XOR U16040 ( .A(n11692), .B(n11693), .Z(n11766) );
  XOR U16041 ( .A(n11698), .B(n11767), .Z(n11693) );
  XOR U16042 ( .A(n11697), .B(n11700), .Z(n11767) );
  IV U16043 ( .A(n11699), .Z(n11700) );
  NAND U16044 ( .A(n11768), .B(n11769), .Z(n11699) );
  OR U16045 ( .A(n11770), .B(n11771), .Z(n11769) );
  OR U16046 ( .A(n11772), .B(n11773), .Z(n11768) );
  NAND U16047 ( .A(n11774), .B(n11775), .Z(n11697) );
  OR U16048 ( .A(n11776), .B(n11777), .Z(n11775) );
  OR U16049 ( .A(n11778), .B(n11779), .Z(n11774) );
  NOR U16050 ( .A(n11780), .B(n11781), .Z(n11698) );
  ANDN U16051 ( .B(n11782), .A(n11783), .Z(n11692) );
  IV U16052 ( .A(n11784), .Z(n11782) );
  XNOR U16053 ( .A(n11685), .B(n11785), .Z(n11691) );
  XNOR U16054 ( .A(n11684), .B(n11686), .Z(n11785) );
  NAND U16055 ( .A(n11786), .B(n11787), .Z(n11686) );
  OR U16056 ( .A(n11788), .B(n11789), .Z(n11787) );
  OR U16057 ( .A(n11790), .B(n11791), .Z(n11786) );
  NAND U16058 ( .A(n11792), .B(n11793), .Z(n11684) );
  OR U16059 ( .A(n11794), .B(n11795), .Z(n11793) );
  OR U16060 ( .A(n11796), .B(n11797), .Z(n11792) );
  ANDN U16061 ( .B(n11798), .A(n11799), .Z(n11685) );
  IV U16062 ( .A(n11800), .Z(n11798) );
  XNOR U16063 ( .A(n11765), .B(n11764), .Z(N29189) );
  XOR U16064 ( .A(n11784), .B(n11783), .Z(n11764) );
  XNOR U16065 ( .A(n11799), .B(n11800), .Z(n11783) );
  XNOR U16066 ( .A(n11794), .B(n11795), .Z(n11800) );
  XNOR U16067 ( .A(n11796), .B(n11797), .Z(n11795) );
  XNOR U16068 ( .A(y[2524]), .B(x[2524]), .Z(n11797) );
  XNOR U16069 ( .A(y[2525]), .B(x[2525]), .Z(n11796) );
  XNOR U16070 ( .A(y[2523]), .B(x[2523]), .Z(n11794) );
  XNOR U16071 ( .A(n11788), .B(n11789), .Z(n11799) );
  XNOR U16072 ( .A(y[2520]), .B(x[2520]), .Z(n11789) );
  XNOR U16073 ( .A(n11790), .B(n11791), .Z(n11788) );
  XNOR U16074 ( .A(y[2521]), .B(x[2521]), .Z(n11791) );
  XNOR U16075 ( .A(y[2522]), .B(x[2522]), .Z(n11790) );
  XNOR U16076 ( .A(n11781), .B(n11780), .Z(n11784) );
  XNOR U16077 ( .A(n11776), .B(n11777), .Z(n11780) );
  XNOR U16078 ( .A(y[2517]), .B(x[2517]), .Z(n11777) );
  XNOR U16079 ( .A(n11778), .B(n11779), .Z(n11776) );
  XNOR U16080 ( .A(y[2518]), .B(x[2518]), .Z(n11779) );
  XNOR U16081 ( .A(y[2519]), .B(x[2519]), .Z(n11778) );
  XNOR U16082 ( .A(n11770), .B(n11771), .Z(n11781) );
  XNOR U16083 ( .A(y[2514]), .B(x[2514]), .Z(n11771) );
  XNOR U16084 ( .A(n11772), .B(n11773), .Z(n11770) );
  XNOR U16085 ( .A(y[2515]), .B(x[2515]), .Z(n11773) );
  XNOR U16086 ( .A(y[2516]), .B(x[2516]), .Z(n11772) );
  XOR U16087 ( .A(n11746), .B(n11747), .Z(n11765) );
  XNOR U16088 ( .A(n11762), .B(n11763), .Z(n11747) );
  XNOR U16089 ( .A(n11757), .B(n11758), .Z(n11763) );
  XNOR U16090 ( .A(n11759), .B(n11760), .Z(n11758) );
  XNOR U16091 ( .A(y[2512]), .B(x[2512]), .Z(n11760) );
  XNOR U16092 ( .A(y[2513]), .B(x[2513]), .Z(n11759) );
  XNOR U16093 ( .A(y[2511]), .B(x[2511]), .Z(n11757) );
  XNOR U16094 ( .A(n11751), .B(n11752), .Z(n11762) );
  XNOR U16095 ( .A(y[2508]), .B(x[2508]), .Z(n11752) );
  XNOR U16096 ( .A(n11753), .B(n11754), .Z(n11751) );
  XNOR U16097 ( .A(y[2509]), .B(x[2509]), .Z(n11754) );
  XNOR U16098 ( .A(y[2510]), .B(x[2510]), .Z(n11753) );
  XOR U16099 ( .A(n11745), .B(n11744), .Z(n11746) );
  XNOR U16100 ( .A(n11740), .B(n11741), .Z(n11744) );
  XNOR U16101 ( .A(y[2505]), .B(x[2505]), .Z(n11741) );
  XNOR U16102 ( .A(n11742), .B(n11743), .Z(n11740) );
  XNOR U16103 ( .A(y[2506]), .B(x[2506]), .Z(n11743) );
  XNOR U16104 ( .A(y[2507]), .B(x[2507]), .Z(n11742) );
  XNOR U16105 ( .A(n11734), .B(n11735), .Z(n11745) );
  XNOR U16106 ( .A(y[2502]), .B(x[2502]), .Z(n11735) );
  XNOR U16107 ( .A(n11736), .B(n11737), .Z(n11734) );
  XNOR U16108 ( .A(y[2503]), .B(x[2503]), .Z(n11737) );
  XNOR U16109 ( .A(y[2504]), .B(x[2504]), .Z(n11736) );
  NAND U16110 ( .A(n11801), .B(n11802), .Z(N29181) );
  NANDN U16111 ( .A(n11803), .B(n11804), .Z(n11802) );
  OR U16112 ( .A(n11805), .B(n11806), .Z(n11804) );
  NAND U16113 ( .A(n11805), .B(n11806), .Z(n11801) );
  XOR U16114 ( .A(n11805), .B(n11807), .Z(N29180) );
  XNOR U16115 ( .A(n11803), .B(n11806), .Z(n11807) );
  AND U16116 ( .A(n11808), .B(n11809), .Z(n11806) );
  NANDN U16117 ( .A(n11810), .B(n11811), .Z(n11809) );
  NANDN U16118 ( .A(n11812), .B(n11813), .Z(n11811) );
  NANDN U16119 ( .A(n11813), .B(n11812), .Z(n11808) );
  NAND U16120 ( .A(n11814), .B(n11815), .Z(n11803) );
  NANDN U16121 ( .A(n11816), .B(n11817), .Z(n11815) );
  OR U16122 ( .A(n11818), .B(n11819), .Z(n11817) );
  NAND U16123 ( .A(n11819), .B(n11818), .Z(n11814) );
  AND U16124 ( .A(n11820), .B(n11821), .Z(n11805) );
  NANDN U16125 ( .A(n11822), .B(n11823), .Z(n11821) );
  NANDN U16126 ( .A(n11824), .B(n11825), .Z(n11823) );
  NANDN U16127 ( .A(n11825), .B(n11824), .Z(n11820) );
  XOR U16128 ( .A(n11819), .B(n11826), .Z(N29179) );
  XOR U16129 ( .A(n11816), .B(n11818), .Z(n11826) );
  XNOR U16130 ( .A(n11812), .B(n11827), .Z(n11818) );
  XNOR U16131 ( .A(n11810), .B(n11813), .Z(n11827) );
  NAND U16132 ( .A(n11828), .B(n11829), .Z(n11813) );
  NAND U16133 ( .A(n11830), .B(n11831), .Z(n11829) );
  OR U16134 ( .A(n11832), .B(n11833), .Z(n11830) );
  NANDN U16135 ( .A(n11834), .B(n11832), .Z(n11828) );
  IV U16136 ( .A(n11833), .Z(n11834) );
  NAND U16137 ( .A(n11835), .B(n11836), .Z(n11810) );
  NAND U16138 ( .A(n11837), .B(n11838), .Z(n11836) );
  NANDN U16139 ( .A(n11839), .B(n11840), .Z(n11837) );
  NANDN U16140 ( .A(n11840), .B(n11839), .Z(n11835) );
  AND U16141 ( .A(n11841), .B(n11842), .Z(n11812) );
  NAND U16142 ( .A(n11843), .B(n11844), .Z(n11842) );
  OR U16143 ( .A(n11845), .B(n11846), .Z(n11843) );
  NANDN U16144 ( .A(n11847), .B(n11845), .Z(n11841) );
  NAND U16145 ( .A(n11848), .B(n11849), .Z(n11816) );
  NANDN U16146 ( .A(n11850), .B(n11851), .Z(n11849) );
  OR U16147 ( .A(n11852), .B(n11853), .Z(n11851) );
  NANDN U16148 ( .A(n11854), .B(n11852), .Z(n11848) );
  IV U16149 ( .A(n11853), .Z(n11854) );
  XNOR U16150 ( .A(n11824), .B(n11855), .Z(n11819) );
  XNOR U16151 ( .A(n11822), .B(n11825), .Z(n11855) );
  NAND U16152 ( .A(n11856), .B(n11857), .Z(n11825) );
  NAND U16153 ( .A(n11858), .B(n11859), .Z(n11857) );
  OR U16154 ( .A(n11860), .B(n11861), .Z(n11858) );
  NANDN U16155 ( .A(n11862), .B(n11860), .Z(n11856) );
  IV U16156 ( .A(n11861), .Z(n11862) );
  NAND U16157 ( .A(n11863), .B(n11864), .Z(n11822) );
  NAND U16158 ( .A(n11865), .B(n11866), .Z(n11864) );
  NANDN U16159 ( .A(n11867), .B(n11868), .Z(n11865) );
  NANDN U16160 ( .A(n11868), .B(n11867), .Z(n11863) );
  AND U16161 ( .A(n11869), .B(n11870), .Z(n11824) );
  NAND U16162 ( .A(n11871), .B(n11872), .Z(n11870) );
  OR U16163 ( .A(n11873), .B(n11874), .Z(n11871) );
  NANDN U16164 ( .A(n11875), .B(n11873), .Z(n11869) );
  XNOR U16165 ( .A(n11850), .B(n11876), .Z(N29178) );
  XOR U16166 ( .A(n11852), .B(n11853), .Z(n11876) );
  XNOR U16167 ( .A(n11866), .B(n11877), .Z(n11853) );
  XOR U16168 ( .A(n11867), .B(n11868), .Z(n11877) );
  XOR U16169 ( .A(n11873), .B(n11878), .Z(n11868) );
  XOR U16170 ( .A(n11872), .B(n11875), .Z(n11878) );
  IV U16171 ( .A(n11874), .Z(n11875) );
  NAND U16172 ( .A(n11879), .B(n11880), .Z(n11874) );
  OR U16173 ( .A(n11881), .B(n11882), .Z(n11880) );
  OR U16174 ( .A(n11883), .B(n11884), .Z(n11879) );
  NAND U16175 ( .A(n11885), .B(n11886), .Z(n11872) );
  OR U16176 ( .A(n11887), .B(n11888), .Z(n11886) );
  OR U16177 ( .A(n11889), .B(n11890), .Z(n11885) );
  NOR U16178 ( .A(n11891), .B(n11892), .Z(n11873) );
  ANDN U16179 ( .B(n11893), .A(n11894), .Z(n11867) );
  XNOR U16180 ( .A(n11860), .B(n11895), .Z(n11866) );
  XNOR U16181 ( .A(n11859), .B(n11861), .Z(n11895) );
  NAND U16182 ( .A(n11896), .B(n11897), .Z(n11861) );
  OR U16183 ( .A(n11898), .B(n11899), .Z(n11897) );
  OR U16184 ( .A(n11900), .B(n11901), .Z(n11896) );
  NAND U16185 ( .A(n11902), .B(n11903), .Z(n11859) );
  OR U16186 ( .A(n11904), .B(n11905), .Z(n11903) );
  OR U16187 ( .A(n11906), .B(n11907), .Z(n11902) );
  ANDN U16188 ( .B(n11908), .A(n11909), .Z(n11860) );
  IV U16189 ( .A(n11910), .Z(n11908) );
  ANDN U16190 ( .B(n11911), .A(n11912), .Z(n11852) );
  XOR U16191 ( .A(n11838), .B(n11913), .Z(n11850) );
  XOR U16192 ( .A(n11839), .B(n11840), .Z(n11913) );
  XOR U16193 ( .A(n11845), .B(n11914), .Z(n11840) );
  XOR U16194 ( .A(n11844), .B(n11847), .Z(n11914) );
  IV U16195 ( .A(n11846), .Z(n11847) );
  NAND U16196 ( .A(n11915), .B(n11916), .Z(n11846) );
  OR U16197 ( .A(n11917), .B(n11918), .Z(n11916) );
  OR U16198 ( .A(n11919), .B(n11920), .Z(n11915) );
  NAND U16199 ( .A(n11921), .B(n11922), .Z(n11844) );
  OR U16200 ( .A(n11923), .B(n11924), .Z(n11922) );
  OR U16201 ( .A(n11925), .B(n11926), .Z(n11921) );
  NOR U16202 ( .A(n11927), .B(n11928), .Z(n11845) );
  ANDN U16203 ( .B(n11929), .A(n11930), .Z(n11839) );
  IV U16204 ( .A(n11931), .Z(n11929) );
  XNOR U16205 ( .A(n11832), .B(n11932), .Z(n11838) );
  XNOR U16206 ( .A(n11831), .B(n11833), .Z(n11932) );
  NAND U16207 ( .A(n11933), .B(n11934), .Z(n11833) );
  OR U16208 ( .A(n11935), .B(n11936), .Z(n11934) );
  OR U16209 ( .A(n11937), .B(n11938), .Z(n11933) );
  NAND U16210 ( .A(n11939), .B(n11940), .Z(n11831) );
  OR U16211 ( .A(n11941), .B(n11942), .Z(n11940) );
  OR U16212 ( .A(n11943), .B(n11944), .Z(n11939) );
  ANDN U16213 ( .B(n11945), .A(n11946), .Z(n11832) );
  IV U16214 ( .A(n11947), .Z(n11945) );
  XNOR U16215 ( .A(n11912), .B(n11911), .Z(N29177) );
  XOR U16216 ( .A(n11931), .B(n11930), .Z(n11911) );
  XNOR U16217 ( .A(n11946), .B(n11947), .Z(n11930) );
  XNOR U16218 ( .A(n11941), .B(n11942), .Z(n11947) );
  XNOR U16219 ( .A(n11943), .B(n11944), .Z(n11942) );
  XNOR U16220 ( .A(y[2500]), .B(x[2500]), .Z(n11944) );
  XNOR U16221 ( .A(y[2501]), .B(x[2501]), .Z(n11943) );
  XNOR U16222 ( .A(y[2499]), .B(x[2499]), .Z(n11941) );
  XNOR U16223 ( .A(n11935), .B(n11936), .Z(n11946) );
  XNOR U16224 ( .A(y[2496]), .B(x[2496]), .Z(n11936) );
  XNOR U16225 ( .A(n11937), .B(n11938), .Z(n11935) );
  XNOR U16226 ( .A(y[2497]), .B(x[2497]), .Z(n11938) );
  XNOR U16227 ( .A(y[2498]), .B(x[2498]), .Z(n11937) );
  XNOR U16228 ( .A(n11928), .B(n11927), .Z(n11931) );
  XNOR U16229 ( .A(n11923), .B(n11924), .Z(n11927) );
  XNOR U16230 ( .A(y[2493]), .B(x[2493]), .Z(n11924) );
  XNOR U16231 ( .A(n11925), .B(n11926), .Z(n11923) );
  XNOR U16232 ( .A(y[2494]), .B(x[2494]), .Z(n11926) );
  XNOR U16233 ( .A(y[2495]), .B(x[2495]), .Z(n11925) );
  XNOR U16234 ( .A(n11917), .B(n11918), .Z(n11928) );
  XNOR U16235 ( .A(y[2490]), .B(x[2490]), .Z(n11918) );
  XNOR U16236 ( .A(n11919), .B(n11920), .Z(n11917) );
  XNOR U16237 ( .A(y[2491]), .B(x[2491]), .Z(n11920) );
  XNOR U16238 ( .A(y[2492]), .B(x[2492]), .Z(n11919) );
  XOR U16239 ( .A(n11893), .B(n11894), .Z(n11912) );
  XNOR U16240 ( .A(n11909), .B(n11910), .Z(n11894) );
  XNOR U16241 ( .A(n11904), .B(n11905), .Z(n11910) );
  XNOR U16242 ( .A(n11906), .B(n11907), .Z(n11905) );
  XNOR U16243 ( .A(y[2488]), .B(x[2488]), .Z(n11907) );
  XNOR U16244 ( .A(y[2489]), .B(x[2489]), .Z(n11906) );
  XNOR U16245 ( .A(y[2487]), .B(x[2487]), .Z(n11904) );
  XNOR U16246 ( .A(n11898), .B(n11899), .Z(n11909) );
  XNOR U16247 ( .A(y[2484]), .B(x[2484]), .Z(n11899) );
  XNOR U16248 ( .A(n11900), .B(n11901), .Z(n11898) );
  XNOR U16249 ( .A(y[2485]), .B(x[2485]), .Z(n11901) );
  XNOR U16250 ( .A(y[2486]), .B(x[2486]), .Z(n11900) );
  XOR U16251 ( .A(n11892), .B(n11891), .Z(n11893) );
  XNOR U16252 ( .A(n11887), .B(n11888), .Z(n11891) );
  XNOR U16253 ( .A(y[2481]), .B(x[2481]), .Z(n11888) );
  XNOR U16254 ( .A(n11889), .B(n11890), .Z(n11887) );
  XNOR U16255 ( .A(y[2482]), .B(x[2482]), .Z(n11890) );
  XNOR U16256 ( .A(y[2483]), .B(x[2483]), .Z(n11889) );
  XNOR U16257 ( .A(n11881), .B(n11882), .Z(n11892) );
  XNOR U16258 ( .A(y[2478]), .B(x[2478]), .Z(n11882) );
  XNOR U16259 ( .A(n11883), .B(n11884), .Z(n11881) );
  XNOR U16260 ( .A(y[2479]), .B(x[2479]), .Z(n11884) );
  XNOR U16261 ( .A(y[2480]), .B(x[2480]), .Z(n11883) );
  NAND U16262 ( .A(n11948), .B(n11949), .Z(N29169) );
  NANDN U16263 ( .A(n11950), .B(n11951), .Z(n11949) );
  OR U16264 ( .A(n11952), .B(n11953), .Z(n11951) );
  NAND U16265 ( .A(n11952), .B(n11953), .Z(n11948) );
  XOR U16266 ( .A(n11952), .B(n11954), .Z(N29168) );
  XNOR U16267 ( .A(n11950), .B(n11953), .Z(n11954) );
  AND U16268 ( .A(n11955), .B(n11956), .Z(n11953) );
  NANDN U16269 ( .A(n11957), .B(n11958), .Z(n11956) );
  NANDN U16270 ( .A(n11959), .B(n11960), .Z(n11958) );
  NANDN U16271 ( .A(n11960), .B(n11959), .Z(n11955) );
  NAND U16272 ( .A(n11961), .B(n11962), .Z(n11950) );
  NANDN U16273 ( .A(n11963), .B(n11964), .Z(n11962) );
  OR U16274 ( .A(n11965), .B(n11966), .Z(n11964) );
  NAND U16275 ( .A(n11966), .B(n11965), .Z(n11961) );
  AND U16276 ( .A(n11967), .B(n11968), .Z(n11952) );
  NANDN U16277 ( .A(n11969), .B(n11970), .Z(n11968) );
  NANDN U16278 ( .A(n11971), .B(n11972), .Z(n11970) );
  NANDN U16279 ( .A(n11972), .B(n11971), .Z(n11967) );
  XOR U16280 ( .A(n11966), .B(n11973), .Z(N29167) );
  XOR U16281 ( .A(n11963), .B(n11965), .Z(n11973) );
  XNOR U16282 ( .A(n11959), .B(n11974), .Z(n11965) );
  XNOR U16283 ( .A(n11957), .B(n11960), .Z(n11974) );
  NAND U16284 ( .A(n11975), .B(n11976), .Z(n11960) );
  NAND U16285 ( .A(n11977), .B(n11978), .Z(n11976) );
  OR U16286 ( .A(n11979), .B(n11980), .Z(n11977) );
  NANDN U16287 ( .A(n11981), .B(n11979), .Z(n11975) );
  IV U16288 ( .A(n11980), .Z(n11981) );
  NAND U16289 ( .A(n11982), .B(n11983), .Z(n11957) );
  NAND U16290 ( .A(n11984), .B(n11985), .Z(n11983) );
  NANDN U16291 ( .A(n11986), .B(n11987), .Z(n11984) );
  NANDN U16292 ( .A(n11987), .B(n11986), .Z(n11982) );
  AND U16293 ( .A(n11988), .B(n11989), .Z(n11959) );
  NAND U16294 ( .A(n11990), .B(n11991), .Z(n11989) );
  OR U16295 ( .A(n11992), .B(n11993), .Z(n11990) );
  NANDN U16296 ( .A(n11994), .B(n11992), .Z(n11988) );
  NAND U16297 ( .A(n11995), .B(n11996), .Z(n11963) );
  NANDN U16298 ( .A(n11997), .B(n11998), .Z(n11996) );
  OR U16299 ( .A(n11999), .B(n12000), .Z(n11998) );
  NANDN U16300 ( .A(n12001), .B(n11999), .Z(n11995) );
  IV U16301 ( .A(n12000), .Z(n12001) );
  XNOR U16302 ( .A(n11971), .B(n12002), .Z(n11966) );
  XNOR U16303 ( .A(n11969), .B(n11972), .Z(n12002) );
  NAND U16304 ( .A(n12003), .B(n12004), .Z(n11972) );
  NAND U16305 ( .A(n12005), .B(n12006), .Z(n12004) );
  OR U16306 ( .A(n12007), .B(n12008), .Z(n12005) );
  NANDN U16307 ( .A(n12009), .B(n12007), .Z(n12003) );
  IV U16308 ( .A(n12008), .Z(n12009) );
  NAND U16309 ( .A(n12010), .B(n12011), .Z(n11969) );
  NAND U16310 ( .A(n12012), .B(n12013), .Z(n12011) );
  NANDN U16311 ( .A(n12014), .B(n12015), .Z(n12012) );
  NANDN U16312 ( .A(n12015), .B(n12014), .Z(n12010) );
  AND U16313 ( .A(n12016), .B(n12017), .Z(n11971) );
  NAND U16314 ( .A(n12018), .B(n12019), .Z(n12017) );
  OR U16315 ( .A(n12020), .B(n12021), .Z(n12018) );
  NANDN U16316 ( .A(n12022), .B(n12020), .Z(n12016) );
  XNOR U16317 ( .A(n11997), .B(n12023), .Z(N29166) );
  XOR U16318 ( .A(n11999), .B(n12000), .Z(n12023) );
  XNOR U16319 ( .A(n12013), .B(n12024), .Z(n12000) );
  XOR U16320 ( .A(n12014), .B(n12015), .Z(n12024) );
  XOR U16321 ( .A(n12020), .B(n12025), .Z(n12015) );
  XOR U16322 ( .A(n12019), .B(n12022), .Z(n12025) );
  IV U16323 ( .A(n12021), .Z(n12022) );
  NAND U16324 ( .A(n12026), .B(n12027), .Z(n12021) );
  OR U16325 ( .A(n12028), .B(n12029), .Z(n12027) );
  OR U16326 ( .A(n12030), .B(n12031), .Z(n12026) );
  NAND U16327 ( .A(n12032), .B(n12033), .Z(n12019) );
  OR U16328 ( .A(n12034), .B(n12035), .Z(n12033) );
  OR U16329 ( .A(n12036), .B(n12037), .Z(n12032) );
  NOR U16330 ( .A(n12038), .B(n12039), .Z(n12020) );
  ANDN U16331 ( .B(n12040), .A(n12041), .Z(n12014) );
  XNOR U16332 ( .A(n12007), .B(n12042), .Z(n12013) );
  XNOR U16333 ( .A(n12006), .B(n12008), .Z(n12042) );
  NAND U16334 ( .A(n12043), .B(n12044), .Z(n12008) );
  OR U16335 ( .A(n12045), .B(n12046), .Z(n12044) );
  OR U16336 ( .A(n12047), .B(n12048), .Z(n12043) );
  NAND U16337 ( .A(n12049), .B(n12050), .Z(n12006) );
  OR U16338 ( .A(n12051), .B(n12052), .Z(n12050) );
  OR U16339 ( .A(n12053), .B(n12054), .Z(n12049) );
  ANDN U16340 ( .B(n12055), .A(n12056), .Z(n12007) );
  IV U16341 ( .A(n12057), .Z(n12055) );
  ANDN U16342 ( .B(n12058), .A(n12059), .Z(n11999) );
  XOR U16343 ( .A(n11985), .B(n12060), .Z(n11997) );
  XOR U16344 ( .A(n11986), .B(n11987), .Z(n12060) );
  XOR U16345 ( .A(n11992), .B(n12061), .Z(n11987) );
  XOR U16346 ( .A(n11991), .B(n11994), .Z(n12061) );
  IV U16347 ( .A(n11993), .Z(n11994) );
  NAND U16348 ( .A(n12062), .B(n12063), .Z(n11993) );
  OR U16349 ( .A(n12064), .B(n12065), .Z(n12063) );
  OR U16350 ( .A(n12066), .B(n12067), .Z(n12062) );
  NAND U16351 ( .A(n12068), .B(n12069), .Z(n11991) );
  OR U16352 ( .A(n12070), .B(n12071), .Z(n12069) );
  OR U16353 ( .A(n12072), .B(n12073), .Z(n12068) );
  NOR U16354 ( .A(n12074), .B(n12075), .Z(n11992) );
  ANDN U16355 ( .B(n12076), .A(n12077), .Z(n11986) );
  IV U16356 ( .A(n12078), .Z(n12076) );
  XNOR U16357 ( .A(n11979), .B(n12079), .Z(n11985) );
  XNOR U16358 ( .A(n11978), .B(n11980), .Z(n12079) );
  NAND U16359 ( .A(n12080), .B(n12081), .Z(n11980) );
  OR U16360 ( .A(n12082), .B(n12083), .Z(n12081) );
  OR U16361 ( .A(n12084), .B(n12085), .Z(n12080) );
  NAND U16362 ( .A(n12086), .B(n12087), .Z(n11978) );
  OR U16363 ( .A(n12088), .B(n12089), .Z(n12087) );
  OR U16364 ( .A(n12090), .B(n12091), .Z(n12086) );
  ANDN U16365 ( .B(n12092), .A(n12093), .Z(n11979) );
  IV U16366 ( .A(n12094), .Z(n12092) );
  XNOR U16367 ( .A(n12059), .B(n12058), .Z(N29165) );
  XOR U16368 ( .A(n12078), .B(n12077), .Z(n12058) );
  XNOR U16369 ( .A(n12093), .B(n12094), .Z(n12077) );
  XNOR U16370 ( .A(n12088), .B(n12089), .Z(n12094) );
  XNOR U16371 ( .A(n12090), .B(n12091), .Z(n12089) );
  XNOR U16372 ( .A(y[2476]), .B(x[2476]), .Z(n12091) );
  XNOR U16373 ( .A(y[2477]), .B(x[2477]), .Z(n12090) );
  XNOR U16374 ( .A(y[2475]), .B(x[2475]), .Z(n12088) );
  XNOR U16375 ( .A(n12082), .B(n12083), .Z(n12093) );
  XNOR U16376 ( .A(y[2472]), .B(x[2472]), .Z(n12083) );
  XNOR U16377 ( .A(n12084), .B(n12085), .Z(n12082) );
  XNOR U16378 ( .A(y[2473]), .B(x[2473]), .Z(n12085) );
  XNOR U16379 ( .A(y[2474]), .B(x[2474]), .Z(n12084) );
  XNOR U16380 ( .A(n12075), .B(n12074), .Z(n12078) );
  XNOR U16381 ( .A(n12070), .B(n12071), .Z(n12074) );
  XNOR U16382 ( .A(y[2469]), .B(x[2469]), .Z(n12071) );
  XNOR U16383 ( .A(n12072), .B(n12073), .Z(n12070) );
  XNOR U16384 ( .A(y[2470]), .B(x[2470]), .Z(n12073) );
  XNOR U16385 ( .A(y[2471]), .B(x[2471]), .Z(n12072) );
  XNOR U16386 ( .A(n12064), .B(n12065), .Z(n12075) );
  XNOR U16387 ( .A(y[2466]), .B(x[2466]), .Z(n12065) );
  XNOR U16388 ( .A(n12066), .B(n12067), .Z(n12064) );
  XNOR U16389 ( .A(y[2467]), .B(x[2467]), .Z(n12067) );
  XNOR U16390 ( .A(y[2468]), .B(x[2468]), .Z(n12066) );
  XOR U16391 ( .A(n12040), .B(n12041), .Z(n12059) );
  XNOR U16392 ( .A(n12056), .B(n12057), .Z(n12041) );
  XNOR U16393 ( .A(n12051), .B(n12052), .Z(n12057) );
  XNOR U16394 ( .A(n12053), .B(n12054), .Z(n12052) );
  XNOR U16395 ( .A(y[2464]), .B(x[2464]), .Z(n12054) );
  XNOR U16396 ( .A(y[2465]), .B(x[2465]), .Z(n12053) );
  XNOR U16397 ( .A(y[2463]), .B(x[2463]), .Z(n12051) );
  XNOR U16398 ( .A(n12045), .B(n12046), .Z(n12056) );
  XNOR U16399 ( .A(y[2460]), .B(x[2460]), .Z(n12046) );
  XNOR U16400 ( .A(n12047), .B(n12048), .Z(n12045) );
  XNOR U16401 ( .A(y[2461]), .B(x[2461]), .Z(n12048) );
  XNOR U16402 ( .A(y[2462]), .B(x[2462]), .Z(n12047) );
  XOR U16403 ( .A(n12039), .B(n12038), .Z(n12040) );
  XNOR U16404 ( .A(n12034), .B(n12035), .Z(n12038) );
  XNOR U16405 ( .A(y[2457]), .B(x[2457]), .Z(n12035) );
  XNOR U16406 ( .A(n12036), .B(n12037), .Z(n12034) );
  XNOR U16407 ( .A(y[2458]), .B(x[2458]), .Z(n12037) );
  XNOR U16408 ( .A(y[2459]), .B(x[2459]), .Z(n12036) );
  XNOR U16409 ( .A(n12028), .B(n12029), .Z(n12039) );
  XNOR U16410 ( .A(y[2454]), .B(x[2454]), .Z(n12029) );
  XNOR U16411 ( .A(n12030), .B(n12031), .Z(n12028) );
  XNOR U16412 ( .A(y[2455]), .B(x[2455]), .Z(n12031) );
  XNOR U16413 ( .A(y[2456]), .B(x[2456]), .Z(n12030) );
  NAND U16414 ( .A(n12095), .B(n12096), .Z(N29157) );
  NANDN U16415 ( .A(n12097), .B(n12098), .Z(n12096) );
  OR U16416 ( .A(n12099), .B(n12100), .Z(n12098) );
  NAND U16417 ( .A(n12099), .B(n12100), .Z(n12095) );
  XOR U16418 ( .A(n12099), .B(n12101), .Z(N29156) );
  XNOR U16419 ( .A(n12097), .B(n12100), .Z(n12101) );
  AND U16420 ( .A(n12102), .B(n12103), .Z(n12100) );
  NANDN U16421 ( .A(n12104), .B(n12105), .Z(n12103) );
  NANDN U16422 ( .A(n12106), .B(n12107), .Z(n12105) );
  NANDN U16423 ( .A(n12107), .B(n12106), .Z(n12102) );
  NAND U16424 ( .A(n12108), .B(n12109), .Z(n12097) );
  NANDN U16425 ( .A(n12110), .B(n12111), .Z(n12109) );
  OR U16426 ( .A(n12112), .B(n12113), .Z(n12111) );
  NAND U16427 ( .A(n12113), .B(n12112), .Z(n12108) );
  AND U16428 ( .A(n12114), .B(n12115), .Z(n12099) );
  NANDN U16429 ( .A(n12116), .B(n12117), .Z(n12115) );
  NANDN U16430 ( .A(n12118), .B(n12119), .Z(n12117) );
  NANDN U16431 ( .A(n12119), .B(n12118), .Z(n12114) );
  XOR U16432 ( .A(n12113), .B(n12120), .Z(N29155) );
  XOR U16433 ( .A(n12110), .B(n12112), .Z(n12120) );
  XNOR U16434 ( .A(n12106), .B(n12121), .Z(n12112) );
  XNOR U16435 ( .A(n12104), .B(n12107), .Z(n12121) );
  NAND U16436 ( .A(n12122), .B(n12123), .Z(n12107) );
  NAND U16437 ( .A(n12124), .B(n12125), .Z(n12123) );
  OR U16438 ( .A(n12126), .B(n12127), .Z(n12124) );
  NANDN U16439 ( .A(n12128), .B(n12126), .Z(n12122) );
  IV U16440 ( .A(n12127), .Z(n12128) );
  NAND U16441 ( .A(n12129), .B(n12130), .Z(n12104) );
  NAND U16442 ( .A(n12131), .B(n12132), .Z(n12130) );
  NANDN U16443 ( .A(n12133), .B(n12134), .Z(n12131) );
  NANDN U16444 ( .A(n12134), .B(n12133), .Z(n12129) );
  AND U16445 ( .A(n12135), .B(n12136), .Z(n12106) );
  NAND U16446 ( .A(n12137), .B(n12138), .Z(n12136) );
  OR U16447 ( .A(n12139), .B(n12140), .Z(n12137) );
  NANDN U16448 ( .A(n12141), .B(n12139), .Z(n12135) );
  NAND U16449 ( .A(n12142), .B(n12143), .Z(n12110) );
  NANDN U16450 ( .A(n12144), .B(n12145), .Z(n12143) );
  OR U16451 ( .A(n12146), .B(n12147), .Z(n12145) );
  NANDN U16452 ( .A(n12148), .B(n12146), .Z(n12142) );
  IV U16453 ( .A(n12147), .Z(n12148) );
  XNOR U16454 ( .A(n12118), .B(n12149), .Z(n12113) );
  XNOR U16455 ( .A(n12116), .B(n12119), .Z(n12149) );
  NAND U16456 ( .A(n12150), .B(n12151), .Z(n12119) );
  NAND U16457 ( .A(n12152), .B(n12153), .Z(n12151) );
  OR U16458 ( .A(n12154), .B(n12155), .Z(n12152) );
  NANDN U16459 ( .A(n12156), .B(n12154), .Z(n12150) );
  IV U16460 ( .A(n12155), .Z(n12156) );
  NAND U16461 ( .A(n12157), .B(n12158), .Z(n12116) );
  NAND U16462 ( .A(n12159), .B(n12160), .Z(n12158) );
  NANDN U16463 ( .A(n12161), .B(n12162), .Z(n12159) );
  NANDN U16464 ( .A(n12162), .B(n12161), .Z(n12157) );
  AND U16465 ( .A(n12163), .B(n12164), .Z(n12118) );
  NAND U16466 ( .A(n12165), .B(n12166), .Z(n12164) );
  OR U16467 ( .A(n12167), .B(n12168), .Z(n12165) );
  NANDN U16468 ( .A(n12169), .B(n12167), .Z(n12163) );
  XNOR U16469 ( .A(n12144), .B(n12170), .Z(N29154) );
  XOR U16470 ( .A(n12146), .B(n12147), .Z(n12170) );
  XNOR U16471 ( .A(n12160), .B(n12171), .Z(n12147) );
  XOR U16472 ( .A(n12161), .B(n12162), .Z(n12171) );
  XOR U16473 ( .A(n12167), .B(n12172), .Z(n12162) );
  XOR U16474 ( .A(n12166), .B(n12169), .Z(n12172) );
  IV U16475 ( .A(n12168), .Z(n12169) );
  NAND U16476 ( .A(n12173), .B(n12174), .Z(n12168) );
  OR U16477 ( .A(n12175), .B(n12176), .Z(n12174) );
  OR U16478 ( .A(n12177), .B(n12178), .Z(n12173) );
  NAND U16479 ( .A(n12179), .B(n12180), .Z(n12166) );
  OR U16480 ( .A(n12181), .B(n12182), .Z(n12180) );
  OR U16481 ( .A(n12183), .B(n12184), .Z(n12179) );
  NOR U16482 ( .A(n12185), .B(n12186), .Z(n12167) );
  ANDN U16483 ( .B(n12187), .A(n12188), .Z(n12161) );
  XNOR U16484 ( .A(n12154), .B(n12189), .Z(n12160) );
  XNOR U16485 ( .A(n12153), .B(n12155), .Z(n12189) );
  NAND U16486 ( .A(n12190), .B(n12191), .Z(n12155) );
  OR U16487 ( .A(n12192), .B(n12193), .Z(n12191) );
  OR U16488 ( .A(n12194), .B(n12195), .Z(n12190) );
  NAND U16489 ( .A(n12196), .B(n12197), .Z(n12153) );
  OR U16490 ( .A(n12198), .B(n12199), .Z(n12197) );
  OR U16491 ( .A(n12200), .B(n12201), .Z(n12196) );
  ANDN U16492 ( .B(n12202), .A(n12203), .Z(n12154) );
  IV U16493 ( .A(n12204), .Z(n12202) );
  ANDN U16494 ( .B(n12205), .A(n12206), .Z(n12146) );
  XOR U16495 ( .A(n12132), .B(n12207), .Z(n12144) );
  XOR U16496 ( .A(n12133), .B(n12134), .Z(n12207) );
  XOR U16497 ( .A(n12139), .B(n12208), .Z(n12134) );
  XOR U16498 ( .A(n12138), .B(n12141), .Z(n12208) );
  IV U16499 ( .A(n12140), .Z(n12141) );
  NAND U16500 ( .A(n12209), .B(n12210), .Z(n12140) );
  OR U16501 ( .A(n12211), .B(n12212), .Z(n12210) );
  OR U16502 ( .A(n12213), .B(n12214), .Z(n12209) );
  NAND U16503 ( .A(n12215), .B(n12216), .Z(n12138) );
  OR U16504 ( .A(n12217), .B(n12218), .Z(n12216) );
  OR U16505 ( .A(n12219), .B(n12220), .Z(n12215) );
  NOR U16506 ( .A(n12221), .B(n12222), .Z(n12139) );
  ANDN U16507 ( .B(n12223), .A(n12224), .Z(n12133) );
  IV U16508 ( .A(n12225), .Z(n12223) );
  XNOR U16509 ( .A(n12126), .B(n12226), .Z(n12132) );
  XNOR U16510 ( .A(n12125), .B(n12127), .Z(n12226) );
  NAND U16511 ( .A(n12227), .B(n12228), .Z(n12127) );
  OR U16512 ( .A(n12229), .B(n12230), .Z(n12228) );
  OR U16513 ( .A(n12231), .B(n12232), .Z(n12227) );
  NAND U16514 ( .A(n12233), .B(n12234), .Z(n12125) );
  OR U16515 ( .A(n12235), .B(n12236), .Z(n12234) );
  OR U16516 ( .A(n12237), .B(n12238), .Z(n12233) );
  ANDN U16517 ( .B(n12239), .A(n12240), .Z(n12126) );
  IV U16518 ( .A(n12241), .Z(n12239) );
  XNOR U16519 ( .A(n12206), .B(n12205), .Z(N29153) );
  XOR U16520 ( .A(n12225), .B(n12224), .Z(n12205) );
  XNOR U16521 ( .A(n12240), .B(n12241), .Z(n12224) );
  XNOR U16522 ( .A(n12235), .B(n12236), .Z(n12241) );
  XNOR U16523 ( .A(n12237), .B(n12238), .Z(n12236) );
  XNOR U16524 ( .A(y[2452]), .B(x[2452]), .Z(n12238) );
  XNOR U16525 ( .A(y[2453]), .B(x[2453]), .Z(n12237) );
  XNOR U16526 ( .A(y[2451]), .B(x[2451]), .Z(n12235) );
  XNOR U16527 ( .A(n12229), .B(n12230), .Z(n12240) );
  XNOR U16528 ( .A(y[2448]), .B(x[2448]), .Z(n12230) );
  XNOR U16529 ( .A(n12231), .B(n12232), .Z(n12229) );
  XNOR U16530 ( .A(y[2449]), .B(x[2449]), .Z(n12232) );
  XNOR U16531 ( .A(y[2450]), .B(x[2450]), .Z(n12231) );
  XNOR U16532 ( .A(n12222), .B(n12221), .Z(n12225) );
  XNOR U16533 ( .A(n12217), .B(n12218), .Z(n12221) );
  XNOR U16534 ( .A(y[2445]), .B(x[2445]), .Z(n12218) );
  XNOR U16535 ( .A(n12219), .B(n12220), .Z(n12217) );
  XNOR U16536 ( .A(y[2446]), .B(x[2446]), .Z(n12220) );
  XNOR U16537 ( .A(y[2447]), .B(x[2447]), .Z(n12219) );
  XNOR U16538 ( .A(n12211), .B(n12212), .Z(n12222) );
  XNOR U16539 ( .A(y[2442]), .B(x[2442]), .Z(n12212) );
  XNOR U16540 ( .A(n12213), .B(n12214), .Z(n12211) );
  XNOR U16541 ( .A(y[2443]), .B(x[2443]), .Z(n12214) );
  XNOR U16542 ( .A(y[2444]), .B(x[2444]), .Z(n12213) );
  XOR U16543 ( .A(n12187), .B(n12188), .Z(n12206) );
  XNOR U16544 ( .A(n12203), .B(n12204), .Z(n12188) );
  XNOR U16545 ( .A(n12198), .B(n12199), .Z(n12204) );
  XNOR U16546 ( .A(n12200), .B(n12201), .Z(n12199) );
  XNOR U16547 ( .A(y[2440]), .B(x[2440]), .Z(n12201) );
  XNOR U16548 ( .A(y[2441]), .B(x[2441]), .Z(n12200) );
  XNOR U16549 ( .A(y[2439]), .B(x[2439]), .Z(n12198) );
  XNOR U16550 ( .A(n12192), .B(n12193), .Z(n12203) );
  XNOR U16551 ( .A(y[2436]), .B(x[2436]), .Z(n12193) );
  XNOR U16552 ( .A(n12194), .B(n12195), .Z(n12192) );
  XNOR U16553 ( .A(y[2437]), .B(x[2437]), .Z(n12195) );
  XNOR U16554 ( .A(y[2438]), .B(x[2438]), .Z(n12194) );
  XOR U16555 ( .A(n12186), .B(n12185), .Z(n12187) );
  XNOR U16556 ( .A(n12181), .B(n12182), .Z(n12185) );
  XNOR U16557 ( .A(y[2433]), .B(x[2433]), .Z(n12182) );
  XNOR U16558 ( .A(n12183), .B(n12184), .Z(n12181) );
  XNOR U16559 ( .A(y[2434]), .B(x[2434]), .Z(n12184) );
  XNOR U16560 ( .A(y[2435]), .B(x[2435]), .Z(n12183) );
  XNOR U16561 ( .A(n12175), .B(n12176), .Z(n12186) );
  XNOR U16562 ( .A(y[2430]), .B(x[2430]), .Z(n12176) );
  XNOR U16563 ( .A(n12177), .B(n12178), .Z(n12175) );
  XNOR U16564 ( .A(y[2431]), .B(x[2431]), .Z(n12178) );
  XNOR U16565 ( .A(y[2432]), .B(x[2432]), .Z(n12177) );
  NAND U16566 ( .A(n12242), .B(n12243), .Z(N29145) );
  NANDN U16567 ( .A(n12244), .B(n12245), .Z(n12243) );
  OR U16568 ( .A(n12246), .B(n12247), .Z(n12245) );
  NAND U16569 ( .A(n12246), .B(n12247), .Z(n12242) );
  XOR U16570 ( .A(n12246), .B(n12248), .Z(N29144) );
  XNOR U16571 ( .A(n12244), .B(n12247), .Z(n12248) );
  AND U16572 ( .A(n12249), .B(n12250), .Z(n12247) );
  NANDN U16573 ( .A(n12251), .B(n12252), .Z(n12250) );
  NANDN U16574 ( .A(n12253), .B(n12254), .Z(n12252) );
  NANDN U16575 ( .A(n12254), .B(n12253), .Z(n12249) );
  NAND U16576 ( .A(n12255), .B(n12256), .Z(n12244) );
  NANDN U16577 ( .A(n12257), .B(n12258), .Z(n12256) );
  OR U16578 ( .A(n12259), .B(n12260), .Z(n12258) );
  NAND U16579 ( .A(n12260), .B(n12259), .Z(n12255) );
  AND U16580 ( .A(n12261), .B(n12262), .Z(n12246) );
  NANDN U16581 ( .A(n12263), .B(n12264), .Z(n12262) );
  NANDN U16582 ( .A(n12265), .B(n12266), .Z(n12264) );
  NANDN U16583 ( .A(n12266), .B(n12265), .Z(n12261) );
  XOR U16584 ( .A(n12260), .B(n12267), .Z(N29143) );
  XOR U16585 ( .A(n12257), .B(n12259), .Z(n12267) );
  XNOR U16586 ( .A(n12253), .B(n12268), .Z(n12259) );
  XNOR U16587 ( .A(n12251), .B(n12254), .Z(n12268) );
  NAND U16588 ( .A(n12269), .B(n12270), .Z(n12254) );
  NAND U16589 ( .A(n12271), .B(n12272), .Z(n12270) );
  OR U16590 ( .A(n12273), .B(n12274), .Z(n12271) );
  NANDN U16591 ( .A(n12275), .B(n12273), .Z(n12269) );
  IV U16592 ( .A(n12274), .Z(n12275) );
  NAND U16593 ( .A(n12276), .B(n12277), .Z(n12251) );
  NAND U16594 ( .A(n12278), .B(n12279), .Z(n12277) );
  NANDN U16595 ( .A(n12280), .B(n12281), .Z(n12278) );
  NANDN U16596 ( .A(n12281), .B(n12280), .Z(n12276) );
  AND U16597 ( .A(n12282), .B(n12283), .Z(n12253) );
  NAND U16598 ( .A(n12284), .B(n12285), .Z(n12283) );
  OR U16599 ( .A(n12286), .B(n12287), .Z(n12284) );
  NANDN U16600 ( .A(n12288), .B(n12286), .Z(n12282) );
  NAND U16601 ( .A(n12289), .B(n12290), .Z(n12257) );
  NANDN U16602 ( .A(n12291), .B(n12292), .Z(n12290) );
  OR U16603 ( .A(n12293), .B(n12294), .Z(n12292) );
  NANDN U16604 ( .A(n12295), .B(n12293), .Z(n12289) );
  IV U16605 ( .A(n12294), .Z(n12295) );
  XNOR U16606 ( .A(n12265), .B(n12296), .Z(n12260) );
  XNOR U16607 ( .A(n12263), .B(n12266), .Z(n12296) );
  NAND U16608 ( .A(n12297), .B(n12298), .Z(n12266) );
  NAND U16609 ( .A(n12299), .B(n12300), .Z(n12298) );
  OR U16610 ( .A(n12301), .B(n12302), .Z(n12299) );
  NANDN U16611 ( .A(n12303), .B(n12301), .Z(n12297) );
  IV U16612 ( .A(n12302), .Z(n12303) );
  NAND U16613 ( .A(n12304), .B(n12305), .Z(n12263) );
  NAND U16614 ( .A(n12306), .B(n12307), .Z(n12305) );
  NANDN U16615 ( .A(n12308), .B(n12309), .Z(n12306) );
  NANDN U16616 ( .A(n12309), .B(n12308), .Z(n12304) );
  AND U16617 ( .A(n12310), .B(n12311), .Z(n12265) );
  NAND U16618 ( .A(n12312), .B(n12313), .Z(n12311) );
  OR U16619 ( .A(n12314), .B(n12315), .Z(n12312) );
  NANDN U16620 ( .A(n12316), .B(n12314), .Z(n12310) );
  XNOR U16621 ( .A(n12291), .B(n12317), .Z(N29142) );
  XOR U16622 ( .A(n12293), .B(n12294), .Z(n12317) );
  XNOR U16623 ( .A(n12307), .B(n12318), .Z(n12294) );
  XOR U16624 ( .A(n12308), .B(n12309), .Z(n12318) );
  XOR U16625 ( .A(n12314), .B(n12319), .Z(n12309) );
  XOR U16626 ( .A(n12313), .B(n12316), .Z(n12319) );
  IV U16627 ( .A(n12315), .Z(n12316) );
  NAND U16628 ( .A(n12320), .B(n12321), .Z(n12315) );
  OR U16629 ( .A(n12322), .B(n12323), .Z(n12321) );
  OR U16630 ( .A(n12324), .B(n12325), .Z(n12320) );
  NAND U16631 ( .A(n12326), .B(n12327), .Z(n12313) );
  OR U16632 ( .A(n12328), .B(n12329), .Z(n12327) );
  OR U16633 ( .A(n12330), .B(n12331), .Z(n12326) );
  NOR U16634 ( .A(n12332), .B(n12333), .Z(n12314) );
  ANDN U16635 ( .B(n12334), .A(n12335), .Z(n12308) );
  XNOR U16636 ( .A(n12301), .B(n12336), .Z(n12307) );
  XNOR U16637 ( .A(n12300), .B(n12302), .Z(n12336) );
  NAND U16638 ( .A(n12337), .B(n12338), .Z(n12302) );
  OR U16639 ( .A(n12339), .B(n12340), .Z(n12338) );
  OR U16640 ( .A(n12341), .B(n12342), .Z(n12337) );
  NAND U16641 ( .A(n12343), .B(n12344), .Z(n12300) );
  OR U16642 ( .A(n12345), .B(n12346), .Z(n12344) );
  OR U16643 ( .A(n12347), .B(n12348), .Z(n12343) );
  ANDN U16644 ( .B(n12349), .A(n12350), .Z(n12301) );
  IV U16645 ( .A(n12351), .Z(n12349) );
  ANDN U16646 ( .B(n12352), .A(n12353), .Z(n12293) );
  XOR U16647 ( .A(n12279), .B(n12354), .Z(n12291) );
  XOR U16648 ( .A(n12280), .B(n12281), .Z(n12354) );
  XOR U16649 ( .A(n12286), .B(n12355), .Z(n12281) );
  XOR U16650 ( .A(n12285), .B(n12288), .Z(n12355) );
  IV U16651 ( .A(n12287), .Z(n12288) );
  NAND U16652 ( .A(n12356), .B(n12357), .Z(n12287) );
  OR U16653 ( .A(n12358), .B(n12359), .Z(n12357) );
  OR U16654 ( .A(n12360), .B(n12361), .Z(n12356) );
  NAND U16655 ( .A(n12362), .B(n12363), .Z(n12285) );
  OR U16656 ( .A(n12364), .B(n12365), .Z(n12363) );
  OR U16657 ( .A(n12366), .B(n12367), .Z(n12362) );
  NOR U16658 ( .A(n12368), .B(n12369), .Z(n12286) );
  ANDN U16659 ( .B(n12370), .A(n12371), .Z(n12280) );
  IV U16660 ( .A(n12372), .Z(n12370) );
  XNOR U16661 ( .A(n12273), .B(n12373), .Z(n12279) );
  XNOR U16662 ( .A(n12272), .B(n12274), .Z(n12373) );
  NAND U16663 ( .A(n12374), .B(n12375), .Z(n12274) );
  OR U16664 ( .A(n12376), .B(n12377), .Z(n12375) );
  OR U16665 ( .A(n12378), .B(n12379), .Z(n12374) );
  NAND U16666 ( .A(n12380), .B(n12381), .Z(n12272) );
  OR U16667 ( .A(n12382), .B(n12383), .Z(n12381) );
  OR U16668 ( .A(n12384), .B(n12385), .Z(n12380) );
  ANDN U16669 ( .B(n12386), .A(n12387), .Z(n12273) );
  IV U16670 ( .A(n12388), .Z(n12386) );
  XNOR U16671 ( .A(n12353), .B(n12352), .Z(N29141) );
  XOR U16672 ( .A(n12372), .B(n12371), .Z(n12352) );
  XNOR U16673 ( .A(n12387), .B(n12388), .Z(n12371) );
  XNOR U16674 ( .A(n12382), .B(n12383), .Z(n12388) );
  XNOR U16675 ( .A(n12384), .B(n12385), .Z(n12383) );
  XNOR U16676 ( .A(y[2428]), .B(x[2428]), .Z(n12385) );
  XNOR U16677 ( .A(y[2429]), .B(x[2429]), .Z(n12384) );
  XNOR U16678 ( .A(y[2427]), .B(x[2427]), .Z(n12382) );
  XNOR U16679 ( .A(n12376), .B(n12377), .Z(n12387) );
  XNOR U16680 ( .A(y[2424]), .B(x[2424]), .Z(n12377) );
  XNOR U16681 ( .A(n12378), .B(n12379), .Z(n12376) );
  XNOR U16682 ( .A(y[2425]), .B(x[2425]), .Z(n12379) );
  XNOR U16683 ( .A(y[2426]), .B(x[2426]), .Z(n12378) );
  XNOR U16684 ( .A(n12369), .B(n12368), .Z(n12372) );
  XNOR U16685 ( .A(n12364), .B(n12365), .Z(n12368) );
  XNOR U16686 ( .A(y[2421]), .B(x[2421]), .Z(n12365) );
  XNOR U16687 ( .A(n12366), .B(n12367), .Z(n12364) );
  XNOR U16688 ( .A(y[2422]), .B(x[2422]), .Z(n12367) );
  XNOR U16689 ( .A(y[2423]), .B(x[2423]), .Z(n12366) );
  XNOR U16690 ( .A(n12358), .B(n12359), .Z(n12369) );
  XNOR U16691 ( .A(y[2418]), .B(x[2418]), .Z(n12359) );
  XNOR U16692 ( .A(n12360), .B(n12361), .Z(n12358) );
  XNOR U16693 ( .A(y[2419]), .B(x[2419]), .Z(n12361) );
  XNOR U16694 ( .A(y[2420]), .B(x[2420]), .Z(n12360) );
  XOR U16695 ( .A(n12334), .B(n12335), .Z(n12353) );
  XNOR U16696 ( .A(n12350), .B(n12351), .Z(n12335) );
  XNOR U16697 ( .A(n12345), .B(n12346), .Z(n12351) );
  XNOR U16698 ( .A(n12347), .B(n12348), .Z(n12346) );
  XNOR U16699 ( .A(y[2416]), .B(x[2416]), .Z(n12348) );
  XNOR U16700 ( .A(y[2417]), .B(x[2417]), .Z(n12347) );
  XNOR U16701 ( .A(y[2415]), .B(x[2415]), .Z(n12345) );
  XNOR U16702 ( .A(n12339), .B(n12340), .Z(n12350) );
  XNOR U16703 ( .A(y[2412]), .B(x[2412]), .Z(n12340) );
  XNOR U16704 ( .A(n12341), .B(n12342), .Z(n12339) );
  XNOR U16705 ( .A(y[2413]), .B(x[2413]), .Z(n12342) );
  XNOR U16706 ( .A(y[2414]), .B(x[2414]), .Z(n12341) );
  XOR U16707 ( .A(n12333), .B(n12332), .Z(n12334) );
  XNOR U16708 ( .A(n12328), .B(n12329), .Z(n12332) );
  XNOR U16709 ( .A(y[2409]), .B(x[2409]), .Z(n12329) );
  XNOR U16710 ( .A(n12330), .B(n12331), .Z(n12328) );
  XNOR U16711 ( .A(y[2410]), .B(x[2410]), .Z(n12331) );
  XNOR U16712 ( .A(y[2411]), .B(x[2411]), .Z(n12330) );
  XNOR U16713 ( .A(n12322), .B(n12323), .Z(n12333) );
  XNOR U16714 ( .A(y[2406]), .B(x[2406]), .Z(n12323) );
  XNOR U16715 ( .A(n12324), .B(n12325), .Z(n12322) );
  XNOR U16716 ( .A(y[2407]), .B(x[2407]), .Z(n12325) );
  XNOR U16717 ( .A(y[2408]), .B(x[2408]), .Z(n12324) );
  NAND U16718 ( .A(n12389), .B(n12390), .Z(N29133) );
  NANDN U16719 ( .A(n12391), .B(n12392), .Z(n12390) );
  OR U16720 ( .A(n12393), .B(n12394), .Z(n12392) );
  NAND U16721 ( .A(n12393), .B(n12394), .Z(n12389) );
  XOR U16722 ( .A(n12393), .B(n12395), .Z(N29132) );
  XNOR U16723 ( .A(n12391), .B(n12394), .Z(n12395) );
  AND U16724 ( .A(n12396), .B(n12397), .Z(n12394) );
  NANDN U16725 ( .A(n12398), .B(n12399), .Z(n12397) );
  NANDN U16726 ( .A(n12400), .B(n12401), .Z(n12399) );
  NANDN U16727 ( .A(n12401), .B(n12400), .Z(n12396) );
  NAND U16728 ( .A(n12402), .B(n12403), .Z(n12391) );
  NANDN U16729 ( .A(n12404), .B(n12405), .Z(n12403) );
  OR U16730 ( .A(n12406), .B(n12407), .Z(n12405) );
  NAND U16731 ( .A(n12407), .B(n12406), .Z(n12402) );
  AND U16732 ( .A(n12408), .B(n12409), .Z(n12393) );
  NANDN U16733 ( .A(n12410), .B(n12411), .Z(n12409) );
  NANDN U16734 ( .A(n12412), .B(n12413), .Z(n12411) );
  NANDN U16735 ( .A(n12413), .B(n12412), .Z(n12408) );
  XOR U16736 ( .A(n12407), .B(n12414), .Z(N29131) );
  XOR U16737 ( .A(n12404), .B(n12406), .Z(n12414) );
  XNOR U16738 ( .A(n12400), .B(n12415), .Z(n12406) );
  XNOR U16739 ( .A(n12398), .B(n12401), .Z(n12415) );
  NAND U16740 ( .A(n12416), .B(n12417), .Z(n12401) );
  NAND U16741 ( .A(n12418), .B(n12419), .Z(n12417) );
  OR U16742 ( .A(n12420), .B(n12421), .Z(n12418) );
  NANDN U16743 ( .A(n12422), .B(n12420), .Z(n12416) );
  IV U16744 ( .A(n12421), .Z(n12422) );
  NAND U16745 ( .A(n12423), .B(n12424), .Z(n12398) );
  NAND U16746 ( .A(n12425), .B(n12426), .Z(n12424) );
  NANDN U16747 ( .A(n12427), .B(n12428), .Z(n12425) );
  NANDN U16748 ( .A(n12428), .B(n12427), .Z(n12423) );
  AND U16749 ( .A(n12429), .B(n12430), .Z(n12400) );
  NAND U16750 ( .A(n12431), .B(n12432), .Z(n12430) );
  OR U16751 ( .A(n12433), .B(n12434), .Z(n12431) );
  NANDN U16752 ( .A(n12435), .B(n12433), .Z(n12429) );
  NAND U16753 ( .A(n12436), .B(n12437), .Z(n12404) );
  NANDN U16754 ( .A(n12438), .B(n12439), .Z(n12437) );
  OR U16755 ( .A(n12440), .B(n12441), .Z(n12439) );
  NANDN U16756 ( .A(n12442), .B(n12440), .Z(n12436) );
  IV U16757 ( .A(n12441), .Z(n12442) );
  XNOR U16758 ( .A(n12412), .B(n12443), .Z(n12407) );
  XNOR U16759 ( .A(n12410), .B(n12413), .Z(n12443) );
  NAND U16760 ( .A(n12444), .B(n12445), .Z(n12413) );
  NAND U16761 ( .A(n12446), .B(n12447), .Z(n12445) );
  OR U16762 ( .A(n12448), .B(n12449), .Z(n12446) );
  NANDN U16763 ( .A(n12450), .B(n12448), .Z(n12444) );
  IV U16764 ( .A(n12449), .Z(n12450) );
  NAND U16765 ( .A(n12451), .B(n12452), .Z(n12410) );
  NAND U16766 ( .A(n12453), .B(n12454), .Z(n12452) );
  NANDN U16767 ( .A(n12455), .B(n12456), .Z(n12453) );
  NANDN U16768 ( .A(n12456), .B(n12455), .Z(n12451) );
  AND U16769 ( .A(n12457), .B(n12458), .Z(n12412) );
  NAND U16770 ( .A(n12459), .B(n12460), .Z(n12458) );
  OR U16771 ( .A(n12461), .B(n12462), .Z(n12459) );
  NANDN U16772 ( .A(n12463), .B(n12461), .Z(n12457) );
  XNOR U16773 ( .A(n12438), .B(n12464), .Z(N29130) );
  XOR U16774 ( .A(n12440), .B(n12441), .Z(n12464) );
  XNOR U16775 ( .A(n12454), .B(n12465), .Z(n12441) );
  XOR U16776 ( .A(n12455), .B(n12456), .Z(n12465) );
  XOR U16777 ( .A(n12461), .B(n12466), .Z(n12456) );
  XOR U16778 ( .A(n12460), .B(n12463), .Z(n12466) );
  IV U16779 ( .A(n12462), .Z(n12463) );
  NAND U16780 ( .A(n12467), .B(n12468), .Z(n12462) );
  OR U16781 ( .A(n12469), .B(n12470), .Z(n12468) );
  OR U16782 ( .A(n12471), .B(n12472), .Z(n12467) );
  NAND U16783 ( .A(n12473), .B(n12474), .Z(n12460) );
  OR U16784 ( .A(n12475), .B(n12476), .Z(n12474) );
  OR U16785 ( .A(n12477), .B(n12478), .Z(n12473) );
  NOR U16786 ( .A(n12479), .B(n12480), .Z(n12461) );
  ANDN U16787 ( .B(n12481), .A(n12482), .Z(n12455) );
  XNOR U16788 ( .A(n12448), .B(n12483), .Z(n12454) );
  XNOR U16789 ( .A(n12447), .B(n12449), .Z(n12483) );
  NAND U16790 ( .A(n12484), .B(n12485), .Z(n12449) );
  OR U16791 ( .A(n12486), .B(n12487), .Z(n12485) );
  OR U16792 ( .A(n12488), .B(n12489), .Z(n12484) );
  NAND U16793 ( .A(n12490), .B(n12491), .Z(n12447) );
  OR U16794 ( .A(n12492), .B(n12493), .Z(n12491) );
  OR U16795 ( .A(n12494), .B(n12495), .Z(n12490) );
  ANDN U16796 ( .B(n12496), .A(n12497), .Z(n12448) );
  IV U16797 ( .A(n12498), .Z(n12496) );
  ANDN U16798 ( .B(n12499), .A(n12500), .Z(n12440) );
  XOR U16799 ( .A(n12426), .B(n12501), .Z(n12438) );
  XOR U16800 ( .A(n12427), .B(n12428), .Z(n12501) );
  XOR U16801 ( .A(n12433), .B(n12502), .Z(n12428) );
  XOR U16802 ( .A(n12432), .B(n12435), .Z(n12502) );
  IV U16803 ( .A(n12434), .Z(n12435) );
  NAND U16804 ( .A(n12503), .B(n12504), .Z(n12434) );
  OR U16805 ( .A(n12505), .B(n12506), .Z(n12504) );
  OR U16806 ( .A(n12507), .B(n12508), .Z(n12503) );
  NAND U16807 ( .A(n12509), .B(n12510), .Z(n12432) );
  OR U16808 ( .A(n12511), .B(n12512), .Z(n12510) );
  OR U16809 ( .A(n12513), .B(n12514), .Z(n12509) );
  NOR U16810 ( .A(n12515), .B(n12516), .Z(n12433) );
  ANDN U16811 ( .B(n12517), .A(n12518), .Z(n12427) );
  IV U16812 ( .A(n12519), .Z(n12517) );
  XNOR U16813 ( .A(n12420), .B(n12520), .Z(n12426) );
  XNOR U16814 ( .A(n12419), .B(n12421), .Z(n12520) );
  NAND U16815 ( .A(n12521), .B(n12522), .Z(n12421) );
  OR U16816 ( .A(n12523), .B(n12524), .Z(n12522) );
  OR U16817 ( .A(n12525), .B(n12526), .Z(n12521) );
  NAND U16818 ( .A(n12527), .B(n12528), .Z(n12419) );
  OR U16819 ( .A(n12529), .B(n12530), .Z(n12528) );
  OR U16820 ( .A(n12531), .B(n12532), .Z(n12527) );
  ANDN U16821 ( .B(n12533), .A(n12534), .Z(n12420) );
  IV U16822 ( .A(n12535), .Z(n12533) );
  XNOR U16823 ( .A(n12500), .B(n12499), .Z(N29129) );
  XOR U16824 ( .A(n12519), .B(n12518), .Z(n12499) );
  XNOR U16825 ( .A(n12534), .B(n12535), .Z(n12518) );
  XNOR U16826 ( .A(n12529), .B(n12530), .Z(n12535) );
  XNOR U16827 ( .A(n12531), .B(n12532), .Z(n12530) );
  XNOR U16828 ( .A(y[2404]), .B(x[2404]), .Z(n12532) );
  XNOR U16829 ( .A(y[2405]), .B(x[2405]), .Z(n12531) );
  XNOR U16830 ( .A(y[2403]), .B(x[2403]), .Z(n12529) );
  XNOR U16831 ( .A(n12523), .B(n12524), .Z(n12534) );
  XNOR U16832 ( .A(y[2400]), .B(x[2400]), .Z(n12524) );
  XNOR U16833 ( .A(n12525), .B(n12526), .Z(n12523) );
  XNOR U16834 ( .A(y[2401]), .B(x[2401]), .Z(n12526) );
  XNOR U16835 ( .A(y[2402]), .B(x[2402]), .Z(n12525) );
  XNOR U16836 ( .A(n12516), .B(n12515), .Z(n12519) );
  XNOR U16837 ( .A(n12511), .B(n12512), .Z(n12515) );
  XNOR U16838 ( .A(y[2397]), .B(x[2397]), .Z(n12512) );
  XNOR U16839 ( .A(n12513), .B(n12514), .Z(n12511) );
  XNOR U16840 ( .A(y[2398]), .B(x[2398]), .Z(n12514) );
  XNOR U16841 ( .A(y[2399]), .B(x[2399]), .Z(n12513) );
  XNOR U16842 ( .A(n12505), .B(n12506), .Z(n12516) );
  XNOR U16843 ( .A(y[2394]), .B(x[2394]), .Z(n12506) );
  XNOR U16844 ( .A(n12507), .B(n12508), .Z(n12505) );
  XNOR U16845 ( .A(y[2395]), .B(x[2395]), .Z(n12508) );
  XNOR U16846 ( .A(y[2396]), .B(x[2396]), .Z(n12507) );
  XOR U16847 ( .A(n12481), .B(n12482), .Z(n12500) );
  XNOR U16848 ( .A(n12497), .B(n12498), .Z(n12482) );
  XNOR U16849 ( .A(n12492), .B(n12493), .Z(n12498) );
  XNOR U16850 ( .A(n12494), .B(n12495), .Z(n12493) );
  XNOR U16851 ( .A(y[2392]), .B(x[2392]), .Z(n12495) );
  XNOR U16852 ( .A(y[2393]), .B(x[2393]), .Z(n12494) );
  XNOR U16853 ( .A(y[2391]), .B(x[2391]), .Z(n12492) );
  XNOR U16854 ( .A(n12486), .B(n12487), .Z(n12497) );
  XNOR U16855 ( .A(y[2388]), .B(x[2388]), .Z(n12487) );
  XNOR U16856 ( .A(n12488), .B(n12489), .Z(n12486) );
  XNOR U16857 ( .A(y[2389]), .B(x[2389]), .Z(n12489) );
  XNOR U16858 ( .A(y[2390]), .B(x[2390]), .Z(n12488) );
  XOR U16859 ( .A(n12480), .B(n12479), .Z(n12481) );
  XNOR U16860 ( .A(n12475), .B(n12476), .Z(n12479) );
  XNOR U16861 ( .A(y[2385]), .B(x[2385]), .Z(n12476) );
  XNOR U16862 ( .A(n12477), .B(n12478), .Z(n12475) );
  XNOR U16863 ( .A(y[2386]), .B(x[2386]), .Z(n12478) );
  XNOR U16864 ( .A(y[2387]), .B(x[2387]), .Z(n12477) );
  XNOR U16865 ( .A(n12469), .B(n12470), .Z(n12480) );
  XNOR U16866 ( .A(y[2382]), .B(x[2382]), .Z(n12470) );
  XNOR U16867 ( .A(n12471), .B(n12472), .Z(n12469) );
  XNOR U16868 ( .A(y[2383]), .B(x[2383]), .Z(n12472) );
  XNOR U16869 ( .A(y[2384]), .B(x[2384]), .Z(n12471) );
  NAND U16870 ( .A(n12536), .B(n12537), .Z(N29121) );
  NANDN U16871 ( .A(n12538), .B(n12539), .Z(n12537) );
  OR U16872 ( .A(n12540), .B(n12541), .Z(n12539) );
  NAND U16873 ( .A(n12540), .B(n12541), .Z(n12536) );
  XOR U16874 ( .A(n12540), .B(n12542), .Z(N29120) );
  XNOR U16875 ( .A(n12538), .B(n12541), .Z(n12542) );
  AND U16876 ( .A(n12543), .B(n12544), .Z(n12541) );
  NANDN U16877 ( .A(n12545), .B(n12546), .Z(n12544) );
  NANDN U16878 ( .A(n12547), .B(n12548), .Z(n12546) );
  NANDN U16879 ( .A(n12548), .B(n12547), .Z(n12543) );
  NAND U16880 ( .A(n12549), .B(n12550), .Z(n12538) );
  NANDN U16881 ( .A(n12551), .B(n12552), .Z(n12550) );
  OR U16882 ( .A(n12553), .B(n12554), .Z(n12552) );
  NAND U16883 ( .A(n12554), .B(n12553), .Z(n12549) );
  AND U16884 ( .A(n12555), .B(n12556), .Z(n12540) );
  NANDN U16885 ( .A(n12557), .B(n12558), .Z(n12556) );
  NANDN U16886 ( .A(n12559), .B(n12560), .Z(n12558) );
  NANDN U16887 ( .A(n12560), .B(n12559), .Z(n12555) );
  XOR U16888 ( .A(n12554), .B(n12561), .Z(N29119) );
  XOR U16889 ( .A(n12551), .B(n12553), .Z(n12561) );
  XNOR U16890 ( .A(n12547), .B(n12562), .Z(n12553) );
  XNOR U16891 ( .A(n12545), .B(n12548), .Z(n12562) );
  NAND U16892 ( .A(n12563), .B(n12564), .Z(n12548) );
  NAND U16893 ( .A(n12565), .B(n12566), .Z(n12564) );
  OR U16894 ( .A(n12567), .B(n12568), .Z(n12565) );
  NANDN U16895 ( .A(n12569), .B(n12567), .Z(n12563) );
  IV U16896 ( .A(n12568), .Z(n12569) );
  NAND U16897 ( .A(n12570), .B(n12571), .Z(n12545) );
  NAND U16898 ( .A(n12572), .B(n12573), .Z(n12571) );
  NANDN U16899 ( .A(n12574), .B(n12575), .Z(n12572) );
  NANDN U16900 ( .A(n12575), .B(n12574), .Z(n12570) );
  AND U16901 ( .A(n12576), .B(n12577), .Z(n12547) );
  NAND U16902 ( .A(n12578), .B(n12579), .Z(n12577) );
  OR U16903 ( .A(n12580), .B(n12581), .Z(n12578) );
  NANDN U16904 ( .A(n12582), .B(n12580), .Z(n12576) );
  NAND U16905 ( .A(n12583), .B(n12584), .Z(n12551) );
  NANDN U16906 ( .A(n12585), .B(n12586), .Z(n12584) );
  OR U16907 ( .A(n12587), .B(n12588), .Z(n12586) );
  NANDN U16908 ( .A(n12589), .B(n12587), .Z(n12583) );
  IV U16909 ( .A(n12588), .Z(n12589) );
  XNOR U16910 ( .A(n12559), .B(n12590), .Z(n12554) );
  XNOR U16911 ( .A(n12557), .B(n12560), .Z(n12590) );
  NAND U16912 ( .A(n12591), .B(n12592), .Z(n12560) );
  NAND U16913 ( .A(n12593), .B(n12594), .Z(n12592) );
  OR U16914 ( .A(n12595), .B(n12596), .Z(n12593) );
  NANDN U16915 ( .A(n12597), .B(n12595), .Z(n12591) );
  IV U16916 ( .A(n12596), .Z(n12597) );
  NAND U16917 ( .A(n12598), .B(n12599), .Z(n12557) );
  NAND U16918 ( .A(n12600), .B(n12601), .Z(n12599) );
  NANDN U16919 ( .A(n12602), .B(n12603), .Z(n12600) );
  NANDN U16920 ( .A(n12603), .B(n12602), .Z(n12598) );
  AND U16921 ( .A(n12604), .B(n12605), .Z(n12559) );
  NAND U16922 ( .A(n12606), .B(n12607), .Z(n12605) );
  OR U16923 ( .A(n12608), .B(n12609), .Z(n12606) );
  NANDN U16924 ( .A(n12610), .B(n12608), .Z(n12604) );
  XNOR U16925 ( .A(n12585), .B(n12611), .Z(N29118) );
  XOR U16926 ( .A(n12587), .B(n12588), .Z(n12611) );
  XNOR U16927 ( .A(n12601), .B(n12612), .Z(n12588) );
  XOR U16928 ( .A(n12602), .B(n12603), .Z(n12612) );
  XOR U16929 ( .A(n12608), .B(n12613), .Z(n12603) );
  XOR U16930 ( .A(n12607), .B(n12610), .Z(n12613) );
  IV U16931 ( .A(n12609), .Z(n12610) );
  NAND U16932 ( .A(n12614), .B(n12615), .Z(n12609) );
  OR U16933 ( .A(n12616), .B(n12617), .Z(n12615) );
  OR U16934 ( .A(n12618), .B(n12619), .Z(n12614) );
  NAND U16935 ( .A(n12620), .B(n12621), .Z(n12607) );
  OR U16936 ( .A(n12622), .B(n12623), .Z(n12621) );
  OR U16937 ( .A(n12624), .B(n12625), .Z(n12620) );
  NOR U16938 ( .A(n12626), .B(n12627), .Z(n12608) );
  ANDN U16939 ( .B(n12628), .A(n12629), .Z(n12602) );
  XNOR U16940 ( .A(n12595), .B(n12630), .Z(n12601) );
  XNOR U16941 ( .A(n12594), .B(n12596), .Z(n12630) );
  NAND U16942 ( .A(n12631), .B(n12632), .Z(n12596) );
  OR U16943 ( .A(n12633), .B(n12634), .Z(n12632) );
  OR U16944 ( .A(n12635), .B(n12636), .Z(n12631) );
  NAND U16945 ( .A(n12637), .B(n12638), .Z(n12594) );
  OR U16946 ( .A(n12639), .B(n12640), .Z(n12638) );
  OR U16947 ( .A(n12641), .B(n12642), .Z(n12637) );
  ANDN U16948 ( .B(n12643), .A(n12644), .Z(n12595) );
  IV U16949 ( .A(n12645), .Z(n12643) );
  ANDN U16950 ( .B(n12646), .A(n12647), .Z(n12587) );
  XOR U16951 ( .A(n12573), .B(n12648), .Z(n12585) );
  XOR U16952 ( .A(n12574), .B(n12575), .Z(n12648) );
  XOR U16953 ( .A(n12580), .B(n12649), .Z(n12575) );
  XOR U16954 ( .A(n12579), .B(n12582), .Z(n12649) );
  IV U16955 ( .A(n12581), .Z(n12582) );
  NAND U16956 ( .A(n12650), .B(n12651), .Z(n12581) );
  OR U16957 ( .A(n12652), .B(n12653), .Z(n12651) );
  OR U16958 ( .A(n12654), .B(n12655), .Z(n12650) );
  NAND U16959 ( .A(n12656), .B(n12657), .Z(n12579) );
  OR U16960 ( .A(n12658), .B(n12659), .Z(n12657) );
  OR U16961 ( .A(n12660), .B(n12661), .Z(n12656) );
  NOR U16962 ( .A(n12662), .B(n12663), .Z(n12580) );
  ANDN U16963 ( .B(n12664), .A(n12665), .Z(n12574) );
  IV U16964 ( .A(n12666), .Z(n12664) );
  XNOR U16965 ( .A(n12567), .B(n12667), .Z(n12573) );
  XNOR U16966 ( .A(n12566), .B(n12568), .Z(n12667) );
  NAND U16967 ( .A(n12668), .B(n12669), .Z(n12568) );
  OR U16968 ( .A(n12670), .B(n12671), .Z(n12669) );
  OR U16969 ( .A(n12672), .B(n12673), .Z(n12668) );
  NAND U16970 ( .A(n12674), .B(n12675), .Z(n12566) );
  OR U16971 ( .A(n12676), .B(n12677), .Z(n12675) );
  OR U16972 ( .A(n12678), .B(n12679), .Z(n12674) );
  ANDN U16973 ( .B(n12680), .A(n12681), .Z(n12567) );
  IV U16974 ( .A(n12682), .Z(n12680) );
  XNOR U16975 ( .A(n12647), .B(n12646), .Z(N29117) );
  XOR U16976 ( .A(n12666), .B(n12665), .Z(n12646) );
  XNOR U16977 ( .A(n12681), .B(n12682), .Z(n12665) );
  XNOR U16978 ( .A(n12676), .B(n12677), .Z(n12682) );
  XNOR U16979 ( .A(n12678), .B(n12679), .Z(n12677) );
  XNOR U16980 ( .A(y[2380]), .B(x[2380]), .Z(n12679) );
  XNOR U16981 ( .A(y[2381]), .B(x[2381]), .Z(n12678) );
  XNOR U16982 ( .A(y[2379]), .B(x[2379]), .Z(n12676) );
  XNOR U16983 ( .A(n12670), .B(n12671), .Z(n12681) );
  XNOR U16984 ( .A(y[2376]), .B(x[2376]), .Z(n12671) );
  XNOR U16985 ( .A(n12672), .B(n12673), .Z(n12670) );
  XNOR U16986 ( .A(y[2377]), .B(x[2377]), .Z(n12673) );
  XNOR U16987 ( .A(y[2378]), .B(x[2378]), .Z(n12672) );
  XNOR U16988 ( .A(n12663), .B(n12662), .Z(n12666) );
  XNOR U16989 ( .A(n12658), .B(n12659), .Z(n12662) );
  XNOR U16990 ( .A(y[2373]), .B(x[2373]), .Z(n12659) );
  XNOR U16991 ( .A(n12660), .B(n12661), .Z(n12658) );
  XNOR U16992 ( .A(y[2374]), .B(x[2374]), .Z(n12661) );
  XNOR U16993 ( .A(y[2375]), .B(x[2375]), .Z(n12660) );
  XNOR U16994 ( .A(n12652), .B(n12653), .Z(n12663) );
  XNOR U16995 ( .A(y[2370]), .B(x[2370]), .Z(n12653) );
  XNOR U16996 ( .A(n12654), .B(n12655), .Z(n12652) );
  XNOR U16997 ( .A(y[2371]), .B(x[2371]), .Z(n12655) );
  XNOR U16998 ( .A(y[2372]), .B(x[2372]), .Z(n12654) );
  XOR U16999 ( .A(n12628), .B(n12629), .Z(n12647) );
  XNOR U17000 ( .A(n12644), .B(n12645), .Z(n12629) );
  XNOR U17001 ( .A(n12639), .B(n12640), .Z(n12645) );
  XNOR U17002 ( .A(n12641), .B(n12642), .Z(n12640) );
  XNOR U17003 ( .A(y[2368]), .B(x[2368]), .Z(n12642) );
  XNOR U17004 ( .A(y[2369]), .B(x[2369]), .Z(n12641) );
  XNOR U17005 ( .A(y[2367]), .B(x[2367]), .Z(n12639) );
  XNOR U17006 ( .A(n12633), .B(n12634), .Z(n12644) );
  XNOR U17007 ( .A(y[2364]), .B(x[2364]), .Z(n12634) );
  XNOR U17008 ( .A(n12635), .B(n12636), .Z(n12633) );
  XNOR U17009 ( .A(y[2365]), .B(x[2365]), .Z(n12636) );
  XNOR U17010 ( .A(y[2366]), .B(x[2366]), .Z(n12635) );
  XOR U17011 ( .A(n12627), .B(n12626), .Z(n12628) );
  XNOR U17012 ( .A(n12622), .B(n12623), .Z(n12626) );
  XNOR U17013 ( .A(y[2361]), .B(x[2361]), .Z(n12623) );
  XNOR U17014 ( .A(n12624), .B(n12625), .Z(n12622) );
  XNOR U17015 ( .A(y[2362]), .B(x[2362]), .Z(n12625) );
  XNOR U17016 ( .A(y[2363]), .B(x[2363]), .Z(n12624) );
  XNOR U17017 ( .A(n12616), .B(n12617), .Z(n12627) );
  XNOR U17018 ( .A(y[2358]), .B(x[2358]), .Z(n12617) );
  XNOR U17019 ( .A(n12618), .B(n12619), .Z(n12616) );
  XNOR U17020 ( .A(y[2359]), .B(x[2359]), .Z(n12619) );
  XNOR U17021 ( .A(y[2360]), .B(x[2360]), .Z(n12618) );
  NAND U17022 ( .A(n12683), .B(n12684), .Z(N29109) );
  NANDN U17023 ( .A(n12685), .B(n12686), .Z(n12684) );
  OR U17024 ( .A(n12687), .B(n12688), .Z(n12686) );
  NAND U17025 ( .A(n12687), .B(n12688), .Z(n12683) );
  XOR U17026 ( .A(n12687), .B(n12689), .Z(N29108) );
  XNOR U17027 ( .A(n12685), .B(n12688), .Z(n12689) );
  AND U17028 ( .A(n12690), .B(n12691), .Z(n12688) );
  NANDN U17029 ( .A(n12692), .B(n12693), .Z(n12691) );
  NANDN U17030 ( .A(n12694), .B(n12695), .Z(n12693) );
  NANDN U17031 ( .A(n12695), .B(n12694), .Z(n12690) );
  NAND U17032 ( .A(n12696), .B(n12697), .Z(n12685) );
  NANDN U17033 ( .A(n12698), .B(n12699), .Z(n12697) );
  OR U17034 ( .A(n12700), .B(n12701), .Z(n12699) );
  NAND U17035 ( .A(n12701), .B(n12700), .Z(n12696) );
  AND U17036 ( .A(n12702), .B(n12703), .Z(n12687) );
  NANDN U17037 ( .A(n12704), .B(n12705), .Z(n12703) );
  NANDN U17038 ( .A(n12706), .B(n12707), .Z(n12705) );
  NANDN U17039 ( .A(n12707), .B(n12706), .Z(n12702) );
  XOR U17040 ( .A(n12701), .B(n12708), .Z(N29107) );
  XOR U17041 ( .A(n12698), .B(n12700), .Z(n12708) );
  XNOR U17042 ( .A(n12694), .B(n12709), .Z(n12700) );
  XNOR U17043 ( .A(n12692), .B(n12695), .Z(n12709) );
  NAND U17044 ( .A(n12710), .B(n12711), .Z(n12695) );
  NAND U17045 ( .A(n12712), .B(n12713), .Z(n12711) );
  OR U17046 ( .A(n12714), .B(n12715), .Z(n12712) );
  NANDN U17047 ( .A(n12716), .B(n12714), .Z(n12710) );
  IV U17048 ( .A(n12715), .Z(n12716) );
  NAND U17049 ( .A(n12717), .B(n12718), .Z(n12692) );
  NAND U17050 ( .A(n12719), .B(n12720), .Z(n12718) );
  NANDN U17051 ( .A(n12721), .B(n12722), .Z(n12719) );
  NANDN U17052 ( .A(n12722), .B(n12721), .Z(n12717) );
  AND U17053 ( .A(n12723), .B(n12724), .Z(n12694) );
  NAND U17054 ( .A(n12725), .B(n12726), .Z(n12724) );
  OR U17055 ( .A(n12727), .B(n12728), .Z(n12725) );
  NANDN U17056 ( .A(n12729), .B(n12727), .Z(n12723) );
  NAND U17057 ( .A(n12730), .B(n12731), .Z(n12698) );
  NANDN U17058 ( .A(n12732), .B(n12733), .Z(n12731) );
  OR U17059 ( .A(n12734), .B(n12735), .Z(n12733) );
  NANDN U17060 ( .A(n12736), .B(n12734), .Z(n12730) );
  IV U17061 ( .A(n12735), .Z(n12736) );
  XNOR U17062 ( .A(n12706), .B(n12737), .Z(n12701) );
  XNOR U17063 ( .A(n12704), .B(n12707), .Z(n12737) );
  NAND U17064 ( .A(n12738), .B(n12739), .Z(n12707) );
  NAND U17065 ( .A(n12740), .B(n12741), .Z(n12739) );
  OR U17066 ( .A(n12742), .B(n12743), .Z(n12740) );
  NANDN U17067 ( .A(n12744), .B(n12742), .Z(n12738) );
  IV U17068 ( .A(n12743), .Z(n12744) );
  NAND U17069 ( .A(n12745), .B(n12746), .Z(n12704) );
  NAND U17070 ( .A(n12747), .B(n12748), .Z(n12746) );
  NANDN U17071 ( .A(n12749), .B(n12750), .Z(n12747) );
  NANDN U17072 ( .A(n12750), .B(n12749), .Z(n12745) );
  AND U17073 ( .A(n12751), .B(n12752), .Z(n12706) );
  NAND U17074 ( .A(n12753), .B(n12754), .Z(n12752) );
  OR U17075 ( .A(n12755), .B(n12756), .Z(n12753) );
  NANDN U17076 ( .A(n12757), .B(n12755), .Z(n12751) );
  XNOR U17077 ( .A(n12732), .B(n12758), .Z(N29106) );
  XOR U17078 ( .A(n12734), .B(n12735), .Z(n12758) );
  XNOR U17079 ( .A(n12748), .B(n12759), .Z(n12735) );
  XOR U17080 ( .A(n12749), .B(n12750), .Z(n12759) );
  XOR U17081 ( .A(n12755), .B(n12760), .Z(n12750) );
  XOR U17082 ( .A(n12754), .B(n12757), .Z(n12760) );
  IV U17083 ( .A(n12756), .Z(n12757) );
  NAND U17084 ( .A(n12761), .B(n12762), .Z(n12756) );
  OR U17085 ( .A(n12763), .B(n12764), .Z(n12762) );
  OR U17086 ( .A(n12765), .B(n12766), .Z(n12761) );
  NAND U17087 ( .A(n12767), .B(n12768), .Z(n12754) );
  OR U17088 ( .A(n12769), .B(n12770), .Z(n12768) );
  OR U17089 ( .A(n12771), .B(n12772), .Z(n12767) );
  NOR U17090 ( .A(n12773), .B(n12774), .Z(n12755) );
  ANDN U17091 ( .B(n12775), .A(n12776), .Z(n12749) );
  XNOR U17092 ( .A(n12742), .B(n12777), .Z(n12748) );
  XNOR U17093 ( .A(n12741), .B(n12743), .Z(n12777) );
  NAND U17094 ( .A(n12778), .B(n12779), .Z(n12743) );
  OR U17095 ( .A(n12780), .B(n12781), .Z(n12779) );
  OR U17096 ( .A(n12782), .B(n12783), .Z(n12778) );
  NAND U17097 ( .A(n12784), .B(n12785), .Z(n12741) );
  OR U17098 ( .A(n12786), .B(n12787), .Z(n12785) );
  OR U17099 ( .A(n12788), .B(n12789), .Z(n12784) );
  ANDN U17100 ( .B(n12790), .A(n12791), .Z(n12742) );
  IV U17101 ( .A(n12792), .Z(n12790) );
  ANDN U17102 ( .B(n12793), .A(n12794), .Z(n12734) );
  XOR U17103 ( .A(n12720), .B(n12795), .Z(n12732) );
  XOR U17104 ( .A(n12721), .B(n12722), .Z(n12795) );
  XOR U17105 ( .A(n12727), .B(n12796), .Z(n12722) );
  XOR U17106 ( .A(n12726), .B(n12729), .Z(n12796) );
  IV U17107 ( .A(n12728), .Z(n12729) );
  NAND U17108 ( .A(n12797), .B(n12798), .Z(n12728) );
  OR U17109 ( .A(n12799), .B(n12800), .Z(n12798) );
  OR U17110 ( .A(n12801), .B(n12802), .Z(n12797) );
  NAND U17111 ( .A(n12803), .B(n12804), .Z(n12726) );
  OR U17112 ( .A(n12805), .B(n12806), .Z(n12804) );
  OR U17113 ( .A(n12807), .B(n12808), .Z(n12803) );
  NOR U17114 ( .A(n12809), .B(n12810), .Z(n12727) );
  ANDN U17115 ( .B(n12811), .A(n12812), .Z(n12721) );
  IV U17116 ( .A(n12813), .Z(n12811) );
  XNOR U17117 ( .A(n12714), .B(n12814), .Z(n12720) );
  XNOR U17118 ( .A(n12713), .B(n12715), .Z(n12814) );
  NAND U17119 ( .A(n12815), .B(n12816), .Z(n12715) );
  OR U17120 ( .A(n12817), .B(n12818), .Z(n12816) );
  OR U17121 ( .A(n12819), .B(n12820), .Z(n12815) );
  NAND U17122 ( .A(n12821), .B(n12822), .Z(n12713) );
  OR U17123 ( .A(n12823), .B(n12824), .Z(n12822) );
  OR U17124 ( .A(n12825), .B(n12826), .Z(n12821) );
  ANDN U17125 ( .B(n12827), .A(n12828), .Z(n12714) );
  IV U17126 ( .A(n12829), .Z(n12827) );
  XNOR U17127 ( .A(n12794), .B(n12793), .Z(N29105) );
  XOR U17128 ( .A(n12813), .B(n12812), .Z(n12793) );
  XNOR U17129 ( .A(n12828), .B(n12829), .Z(n12812) );
  XNOR U17130 ( .A(n12823), .B(n12824), .Z(n12829) );
  XNOR U17131 ( .A(n12825), .B(n12826), .Z(n12824) );
  XNOR U17132 ( .A(y[2356]), .B(x[2356]), .Z(n12826) );
  XNOR U17133 ( .A(y[2357]), .B(x[2357]), .Z(n12825) );
  XNOR U17134 ( .A(y[2355]), .B(x[2355]), .Z(n12823) );
  XNOR U17135 ( .A(n12817), .B(n12818), .Z(n12828) );
  XNOR U17136 ( .A(y[2352]), .B(x[2352]), .Z(n12818) );
  XNOR U17137 ( .A(n12819), .B(n12820), .Z(n12817) );
  XNOR U17138 ( .A(y[2353]), .B(x[2353]), .Z(n12820) );
  XNOR U17139 ( .A(y[2354]), .B(x[2354]), .Z(n12819) );
  XNOR U17140 ( .A(n12810), .B(n12809), .Z(n12813) );
  XNOR U17141 ( .A(n12805), .B(n12806), .Z(n12809) );
  XNOR U17142 ( .A(y[2349]), .B(x[2349]), .Z(n12806) );
  XNOR U17143 ( .A(n12807), .B(n12808), .Z(n12805) );
  XNOR U17144 ( .A(y[2350]), .B(x[2350]), .Z(n12808) );
  XNOR U17145 ( .A(y[2351]), .B(x[2351]), .Z(n12807) );
  XNOR U17146 ( .A(n12799), .B(n12800), .Z(n12810) );
  XNOR U17147 ( .A(y[2346]), .B(x[2346]), .Z(n12800) );
  XNOR U17148 ( .A(n12801), .B(n12802), .Z(n12799) );
  XNOR U17149 ( .A(y[2347]), .B(x[2347]), .Z(n12802) );
  XNOR U17150 ( .A(y[2348]), .B(x[2348]), .Z(n12801) );
  XOR U17151 ( .A(n12775), .B(n12776), .Z(n12794) );
  XNOR U17152 ( .A(n12791), .B(n12792), .Z(n12776) );
  XNOR U17153 ( .A(n12786), .B(n12787), .Z(n12792) );
  XNOR U17154 ( .A(n12788), .B(n12789), .Z(n12787) );
  XNOR U17155 ( .A(y[2344]), .B(x[2344]), .Z(n12789) );
  XNOR U17156 ( .A(y[2345]), .B(x[2345]), .Z(n12788) );
  XNOR U17157 ( .A(y[2343]), .B(x[2343]), .Z(n12786) );
  XNOR U17158 ( .A(n12780), .B(n12781), .Z(n12791) );
  XNOR U17159 ( .A(y[2340]), .B(x[2340]), .Z(n12781) );
  XNOR U17160 ( .A(n12782), .B(n12783), .Z(n12780) );
  XNOR U17161 ( .A(y[2341]), .B(x[2341]), .Z(n12783) );
  XNOR U17162 ( .A(y[2342]), .B(x[2342]), .Z(n12782) );
  XOR U17163 ( .A(n12774), .B(n12773), .Z(n12775) );
  XNOR U17164 ( .A(n12769), .B(n12770), .Z(n12773) );
  XNOR U17165 ( .A(y[2337]), .B(x[2337]), .Z(n12770) );
  XNOR U17166 ( .A(n12771), .B(n12772), .Z(n12769) );
  XNOR U17167 ( .A(y[2338]), .B(x[2338]), .Z(n12772) );
  XNOR U17168 ( .A(y[2339]), .B(x[2339]), .Z(n12771) );
  XNOR U17169 ( .A(n12763), .B(n12764), .Z(n12774) );
  XNOR U17170 ( .A(y[2334]), .B(x[2334]), .Z(n12764) );
  XNOR U17171 ( .A(n12765), .B(n12766), .Z(n12763) );
  XNOR U17172 ( .A(y[2335]), .B(x[2335]), .Z(n12766) );
  XNOR U17173 ( .A(y[2336]), .B(x[2336]), .Z(n12765) );
  NAND U17174 ( .A(n12830), .B(n12831), .Z(N29097) );
  NANDN U17175 ( .A(n12832), .B(n12833), .Z(n12831) );
  OR U17176 ( .A(n12834), .B(n12835), .Z(n12833) );
  NAND U17177 ( .A(n12834), .B(n12835), .Z(n12830) );
  XOR U17178 ( .A(n12834), .B(n12836), .Z(N29096) );
  XNOR U17179 ( .A(n12832), .B(n12835), .Z(n12836) );
  AND U17180 ( .A(n12837), .B(n12838), .Z(n12835) );
  NANDN U17181 ( .A(n12839), .B(n12840), .Z(n12838) );
  NANDN U17182 ( .A(n12841), .B(n12842), .Z(n12840) );
  NANDN U17183 ( .A(n12842), .B(n12841), .Z(n12837) );
  NAND U17184 ( .A(n12843), .B(n12844), .Z(n12832) );
  NANDN U17185 ( .A(n12845), .B(n12846), .Z(n12844) );
  OR U17186 ( .A(n12847), .B(n12848), .Z(n12846) );
  NAND U17187 ( .A(n12848), .B(n12847), .Z(n12843) );
  AND U17188 ( .A(n12849), .B(n12850), .Z(n12834) );
  NANDN U17189 ( .A(n12851), .B(n12852), .Z(n12850) );
  NANDN U17190 ( .A(n12853), .B(n12854), .Z(n12852) );
  NANDN U17191 ( .A(n12854), .B(n12853), .Z(n12849) );
  XOR U17192 ( .A(n12848), .B(n12855), .Z(N29095) );
  XOR U17193 ( .A(n12845), .B(n12847), .Z(n12855) );
  XNOR U17194 ( .A(n12841), .B(n12856), .Z(n12847) );
  XNOR U17195 ( .A(n12839), .B(n12842), .Z(n12856) );
  NAND U17196 ( .A(n12857), .B(n12858), .Z(n12842) );
  NAND U17197 ( .A(n12859), .B(n12860), .Z(n12858) );
  OR U17198 ( .A(n12861), .B(n12862), .Z(n12859) );
  NANDN U17199 ( .A(n12863), .B(n12861), .Z(n12857) );
  IV U17200 ( .A(n12862), .Z(n12863) );
  NAND U17201 ( .A(n12864), .B(n12865), .Z(n12839) );
  NAND U17202 ( .A(n12866), .B(n12867), .Z(n12865) );
  NANDN U17203 ( .A(n12868), .B(n12869), .Z(n12866) );
  NANDN U17204 ( .A(n12869), .B(n12868), .Z(n12864) );
  AND U17205 ( .A(n12870), .B(n12871), .Z(n12841) );
  NAND U17206 ( .A(n12872), .B(n12873), .Z(n12871) );
  OR U17207 ( .A(n12874), .B(n12875), .Z(n12872) );
  NANDN U17208 ( .A(n12876), .B(n12874), .Z(n12870) );
  NAND U17209 ( .A(n12877), .B(n12878), .Z(n12845) );
  NANDN U17210 ( .A(n12879), .B(n12880), .Z(n12878) );
  OR U17211 ( .A(n12881), .B(n12882), .Z(n12880) );
  NANDN U17212 ( .A(n12883), .B(n12881), .Z(n12877) );
  IV U17213 ( .A(n12882), .Z(n12883) );
  XNOR U17214 ( .A(n12853), .B(n12884), .Z(n12848) );
  XNOR U17215 ( .A(n12851), .B(n12854), .Z(n12884) );
  NAND U17216 ( .A(n12885), .B(n12886), .Z(n12854) );
  NAND U17217 ( .A(n12887), .B(n12888), .Z(n12886) );
  OR U17218 ( .A(n12889), .B(n12890), .Z(n12887) );
  NANDN U17219 ( .A(n12891), .B(n12889), .Z(n12885) );
  IV U17220 ( .A(n12890), .Z(n12891) );
  NAND U17221 ( .A(n12892), .B(n12893), .Z(n12851) );
  NAND U17222 ( .A(n12894), .B(n12895), .Z(n12893) );
  NANDN U17223 ( .A(n12896), .B(n12897), .Z(n12894) );
  NANDN U17224 ( .A(n12897), .B(n12896), .Z(n12892) );
  AND U17225 ( .A(n12898), .B(n12899), .Z(n12853) );
  NAND U17226 ( .A(n12900), .B(n12901), .Z(n12899) );
  OR U17227 ( .A(n12902), .B(n12903), .Z(n12900) );
  NANDN U17228 ( .A(n12904), .B(n12902), .Z(n12898) );
  XNOR U17229 ( .A(n12879), .B(n12905), .Z(N29094) );
  XOR U17230 ( .A(n12881), .B(n12882), .Z(n12905) );
  XNOR U17231 ( .A(n12895), .B(n12906), .Z(n12882) );
  XOR U17232 ( .A(n12896), .B(n12897), .Z(n12906) );
  XOR U17233 ( .A(n12902), .B(n12907), .Z(n12897) );
  XOR U17234 ( .A(n12901), .B(n12904), .Z(n12907) );
  IV U17235 ( .A(n12903), .Z(n12904) );
  NAND U17236 ( .A(n12908), .B(n12909), .Z(n12903) );
  OR U17237 ( .A(n12910), .B(n12911), .Z(n12909) );
  OR U17238 ( .A(n12912), .B(n12913), .Z(n12908) );
  NAND U17239 ( .A(n12914), .B(n12915), .Z(n12901) );
  OR U17240 ( .A(n12916), .B(n12917), .Z(n12915) );
  OR U17241 ( .A(n12918), .B(n12919), .Z(n12914) );
  NOR U17242 ( .A(n12920), .B(n12921), .Z(n12902) );
  ANDN U17243 ( .B(n12922), .A(n12923), .Z(n12896) );
  XNOR U17244 ( .A(n12889), .B(n12924), .Z(n12895) );
  XNOR U17245 ( .A(n12888), .B(n12890), .Z(n12924) );
  NAND U17246 ( .A(n12925), .B(n12926), .Z(n12890) );
  OR U17247 ( .A(n12927), .B(n12928), .Z(n12926) );
  OR U17248 ( .A(n12929), .B(n12930), .Z(n12925) );
  NAND U17249 ( .A(n12931), .B(n12932), .Z(n12888) );
  OR U17250 ( .A(n12933), .B(n12934), .Z(n12932) );
  OR U17251 ( .A(n12935), .B(n12936), .Z(n12931) );
  ANDN U17252 ( .B(n12937), .A(n12938), .Z(n12889) );
  IV U17253 ( .A(n12939), .Z(n12937) );
  ANDN U17254 ( .B(n12940), .A(n12941), .Z(n12881) );
  XOR U17255 ( .A(n12867), .B(n12942), .Z(n12879) );
  XOR U17256 ( .A(n12868), .B(n12869), .Z(n12942) );
  XOR U17257 ( .A(n12874), .B(n12943), .Z(n12869) );
  XOR U17258 ( .A(n12873), .B(n12876), .Z(n12943) );
  IV U17259 ( .A(n12875), .Z(n12876) );
  NAND U17260 ( .A(n12944), .B(n12945), .Z(n12875) );
  OR U17261 ( .A(n12946), .B(n12947), .Z(n12945) );
  OR U17262 ( .A(n12948), .B(n12949), .Z(n12944) );
  NAND U17263 ( .A(n12950), .B(n12951), .Z(n12873) );
  OR U17264 ( .A(n12952), .B(n12953), .Z(n12951) );
  OR U17265 ( .A(n12954), .B(n12955), .Z(n12950) );
  NOR U17266 ( .A(n12956), .B(n12957), .Z(n12874) );
  ANDN U17267 ( .B(n12958), .A(n12959), .Z(n12868) );
  IV U17268 ( .A(n12960), .Z(n12958) );
  XNOR U17269 ( .A(n12861), .B(n12961), .Z(n12867) );
  XNOR U17270 ( .A(n12860), .B(n12862), .Z(n12961) );
  NAND U17271 ( .A(n12962), .B(n12963), .Z(n12862) );
  OR U17272 ( .A(n12964), .B(n12965), .Z(n12963) );
  OR U17273 ( .A(n12966), .B(n12967), .Z(n12962) );
  NAND U17274 ( .A(n12968), .B(n12969), .Z(n12860) );
  OR U17275 ( .A(n12970), .B(n12971), .Z(n12969) );
  OR U17276 ( .A(n12972), .B(n12973), .Z(n12968) );
  ANDN U17277 ( .B(n12974), .A(n12975), .Z(n12861) );
  IV U17278 ( .A(n12976), .Z(n12974) );
  XNOR U17279 ( .A(n12941), .B(n12940), .Z(N29093) );
  XOR U17280 ( .A(n12960), .B(n12959), .Z(n12940) );
  XNOR U17281 ( .A(n12975), .B(n12976), .Z(n12959) );
  XNOR U17282 ( .A(n12970), .B(n12971), .Z(n12976) );
  XNOR U17283 ( .A(n12972), .B(n12973), .Z(n12971) );
  XNOR U17284 ( .A(y[2332]), .B(x[2332]), .Z(n12973) );
  XNOR U17285 ( .A(y[2333]), .B(x[2333]), .Z(n12972) );
  XNOR U17286 ( .A(y[2331]), .B(x[2331]), .Z(n12970) );
  XNOR U17287 ( .A(n12964), .B(n12965), .Z(n12975) );
  XNOR U17288 ( .A(y[2328]), .B(x[2328]), .Z(n12965) );
  XNOR U17289 ( .A(n12966), .B(n12967), .Z(n12964) );
  XNOR U17290 ( .A(y[2329]), .B(x[2329]), .Z(n12967) );
  XNOR U17291 ( .A(y[2330]), .B(x[2330]), .Z(n12966) );
  XNOR U17292 ( .A(n12957), .B(n12956), .Z(n12960) );
  XNOR U17293 ( .A(n12952), .B(n12953), .Z(n12956) );
  XNOR U17294 ( .A(y[2325]), .B(x[2325]), .Z(n12953) );
  XNOR U17295 ( .A(n12954), .B(n12955), .Z(n12952) );
  XNOR U17296 ( .A(y[2326]), .B(x[2326]), .Z(n12955) );
  XNOR U17297 ( .A(y[2327]), .B(x[2327]), .Z(n12954) );
  XNOR U17298 ( .A(n12946), .B(n12947), .Z(n12957) );
  XNOR U17299 ( .A(y[2322]), .B(x[2322]), .Z(n12947) );
  XNOR U17300 ( .A(n12948), .B(n12949), .Z(n12946) );
  XNOR U17301 ( .A(y[2323]), .B(x[2323]), .Z(n12949) );
  XNOR U17302 ( .A(y[2324]), .B(x[2324]), .Z(n12948) );
  XOR U17303 ( .A(n12922), .B(n12923), .Z(n12941) );
  XNOR U17304 ( .A(n12938), .B(n12939), .Z(n12923) );
  XNOR U17305 ( .A(n12933), .B(n12934), .Z(n12939) );
  XNOR U17306 ( .A(n12935), .B(n12936), .Z(n12934) );
  XNOR U17307 ( .A(y[2320]), .B(x[2320]), .Z(n12936) );
  XNOR U17308 ( .A(y[2321]), .B(x[2321]), .Z(n12935) );
  XNOR U17309 ( .A(y[2319]), .B(x[2319]), .Z(n12933) );
  XNOR U17310 ( .A(n12927), .B(n12928), .Z(n12938) );
  XNOR U17311 ( .A(y[2316]), .B(x[2316]), .Z(n12928) );
  XNOR U17312 ( .A(n12929), .B(n12930), .Z(n12927) );
  XNOR U17313 ( .A(y[2317]), .B(x[2317]), .Z(n12930) );
  XNOR U17314 ( .A(y[2318]), .B(x[2318]), .Z(n12929) );
  XOR U17315 ( .A(n12921), .B(n12920), .Z(n12922) );
  XNOR U17316 ( .A(n12916), .B(n12917), .Z(n12920) );
  XNOR U17317 ( .A(y[2313]), .B(x[2313]), .Z(n12917) );
  XNOR U17318 ( .A(n12918), .B(n12919), .Z(n12916) );
  XNOR U17319 ( .A(y[2314]), .B(x[2314]), .Z(n12919) );
  XNOR U17320 ( .A(y[2315]), .B(x[2315]), .Z(n12918) );
  XNOR U17321 ( .A(n12910), .B(n12911), .Z(n12921) );
  XNOR U17322 ( .A(y[2310]), .B(x[2310]), .Z(n12911) );
  XNOR U17323 ( .A(n12912), .B(n12913), .Z(n12910) );
  XNOR U17324 ( .A(y[2311]), .B(x[2311]), .Z(n12913) );
  XNOR U17325 ( .A(y[2312]), .B(x[2312]), .Z(n12912) );
  NAND U17326 ( .A(n12977), .B(n12978), .Z(N29085) );
  NANDN U17327 ( .A(n12979), .B(n12980), .Z(n12978) );
  OR U17328 ( .A(n12981), .B(n12982), .Z(n12980) );
  NAND U17329 ( .A(n12981), .B(n12982), .Z(n12977) );
  XOR U17330 ( .A(n12981), .B(n12983), .Z(N29084) );
  XNOR U17331 ( .A(n12979), .B(n12982), .Z(n12983) );
  AND U17332 ( .A(n12984), .B(n12985), .Z(n12982) );
  NANDN U17333 ( .A(n12986), .B(n12987), .Z(n12985) );
  NANDN U17334 ( .A(n12988), .B(n12989), .Z(n12987) );
  NANDN U17335 ( .A(n12989), .B(n12988), .Z(n12984) );
  NAND U17336 ( .A(n12990), .B(n12991), .Z(n12979) );
  NANDN U17337 ( .A(n12992), .B(n12993), .Z(n12991) );
  OR U17338 ( .A(n12994), .B(n12995), .Z(n12993) );
  NAND U17339 ( .A(n12995), .B(n12994), .Z(n12990) );
  AND U17340 ( .A(n12996), .B(n12997), .Z(n12981) );
  NANDN U17341 ( .A(n12998), .B(n12999), .Z(n12997) );
  NANDN U17342 ( .A(n13000), .B(n13001), .Z(n12999) );
  NANDN U17343 ( .A(n13001), .B(n13000), .Z(n12996) );
  XOR U17344 ( .A(n12995), .B(n13002), .Z(N29083) );
  XOR U17345 ( .A(n12992), .B(n12994), .Z(n13002) );
  XNOR U17346 ( .A(n12988), .B(n13003), .Z(n12994) );
  XNOR U17347 ( .A(n12986), .B(n12989), .Z(n13003) );
  NAND U17348 ( .A(n13004), .B(n13005), .Z(n12989) );
  NAND U17349 ( .A(n13006), .B(n13007), .Z(n13005) );
  OR U17350 ( .A(n13008), .B(n13009), .Z(n13006) );
  NANDN U17351 ( .A(n13010), .B(n13008), .Z(n13004) );
  IV U17352 ( .A(n13009), .Z(n13010) );
  NAND U17353 ( .A(n13011), .B(n13012), .Z(n12986) );
  NAND U17354 ( .A(n13013), .B(n13014), .Z(n13012) );
  NANDN U17355 ( .A(n13015), .B(n13016), .Z(n13013) );
  NANDN U17356 ( .A(n13016), .B(n13015), .Z(n13011) );
  AND U17357 ( .A(n13017), .B(n13018), .Z(n12988) );
  NAND U17358 ( .A(n13019), .B(n13020), .Z(n13018) );
  OR U17359 ( .A(n13021), .B(n13022), .Z(n13019) );
  NANDN U17360 ( .A(n13023), .B(n13021), .Z(n13017) );
  NAND U17361 ( .A(n13024), .B(n13025), .Z(n12992) );
  NANDN U17362 ( .A(n13026), .B(n13027), .Z(n13025) );
  OR U17363 ( .A(n13028), .B(n13029), .Z(n13027) );
  NANDN U17364 ( .A(n13030), .B(n13028), .Z(n13024) );
  IV U17365 ( .A(n13029), .Z(n13030) );
  XNOR U17366 ( .A(n13000), .B(n13031), .Z(n12995) );
  XNOR U17367 ( .A(n12998), .B(n13001), .Z(n13031) );
  NAND U17368 ( .A(n13032), .B(n13033), .Z(n13001) );
  NAND U17369 ( .A(n13034), .B(n13035), .Z(n13033) );
  OR U17370 ( .A(n13036), .B(n13037), .Z(n13034) );
  NANDN U17371 ( .A(n13038), .B(n13036), .Z(n13032) );
  IV U17372 ( .A(n13037), .Z(n13038) );
  NAND U17373 ( .A(n13039), .B(n13040), .Z(n12998) );
  NAND U17374 ( .A(n13041), .B(n13042), .Z(n13040) );
  NANDN U17375 ( .A(n13043), .B(n13044), .Z(n13041) );
  NANDN U17376 ( .A(n13044), .B(n13043), .Z(n13039) );
  AND U17377 ( .A(n13045), .B(n13046), .Z(n13000) );
  NAND U17378 ( .A(n13047), .B(n13048), .Z(n13046) );
  OR U17379 ( .A(n13049), .B(n13050), .Z(n13047) );
  NANDN U17380 ( .A(n13051), .B(n13049), .Z(n13045) );
  XNOR U17381 ( .A(n13026), .B(n13052), .Z(N29082) );
  XOR U17382 ( .A(n13028), .B(n13029), .Z(n13052) );
  XNOR U17383 ( .A(n13042), .B(n13053), .Z(n13029) );
  XOR U17384 ( .A(n13043), .B(n13044), .Z(n13053) );
  XOR U17385 ( .A(n13049), .B(n13054), .Z(n13044) );
  XOR U17386 ( .A(n13048), .B(n13051), .Z(n13054) );
  IV U17387 ( .A(n13050), .Z(n13051) );
  NAND U17388 ( .A(n13055), .B(n13056), .Z(n13050) );
  OR U17389 ( .A(n13057), .B(n13058), .Z(n13056) );
  OR U17390 ( .A(n13059), .B(n13060), .Z(n13055) );
  NAND U17391 ( .A(n13061), .B(n13062), .Z(n13048) );
  OR U17392 ( .A(n13063), .B(n13064), .Z(n13062) );
  OR U17393 ( .A(n13065), .B(n13066), .Z(n13061) );
  NOR U17394 ( .A(n13067), .B(n13068), .Z(n13049) );
  ANDN U17395 ( .B(n13069), .A(n13070), .Z(n13043) );
  XNOR U17396 ( .A(n13036), .B(n13071), .Z(n13042) );
  XNOR U17397 ( .A(n13035), .B(n13037), .Z(n13071) );
  NAND U17398 ( .A(n13072), .B(n13073), .Z(n13037) );
  OR U17399 ( .A(n13074), .B(n13075), .Z(n13073) );
  OR U17400 ( .A(n13076), .B(n13077), .Z(n13072) );
  NAND U17401 ( .A(n13078), .B(n13079), .Z(n13035) );
  OR U17402 ( .A(n13080), .B(n13081), .Z(n13079) );
  OR U17403 ( .A(n13082), .B(n13083), .Z(n13078) );
  ANDN U17404 ( .B(n13084), .A(n13085), .Z(n13036) );
  IV U17405 ( .A(n13086), .Z(n13084) );
  ANDN U17406 ( .B(n13087), .A(n13088), .Z(n13028) );
  XOR U17407 ( .A(n13014), .B(n13089), .Z(n13026) );
  XOR U17408 ( .A(n13015), .B(n13016), .Z(n13089) );
  XOR U17409 ( .A(n13021), .B(n13090), .Z(n13016) );
  XOR U17410 ( .A(n13020), .B(n13023), .Z(n13090) );
  IV U17411 ( .A(n13022), .Z(n13023) );
  NAND U17412 ( .A(n13091), .B(n13092), .Z(n13022) );
  OR U17413 ( .A(n13093), .B(n13094), .Z(n13092) );
  OR U17414 ( .A(n13095), .B(n13096), .Z(n13091) );
  NAND U17415 ( .A(n13097), .B(n13098), .Z(n13020) );
  OR U17416 ( .A(n13099), .B(n13100), .Z(n13098) );
  OR U17417 ( .A(n13101), .B(n13102), .Z(n13097) );
  NOR U17418 ( .A(n13103), .B(n13104), .Z(n13021) );
  ANDN U17419 ( .B(n13105), .A(n13106), .Z(n13015) );
  IV U17420 ( .A(n13107), .Z(n13105) );
  XNOR U17421 ( .A(n13008), .B(n13108), .Z(n13014) );
  XNOR U17422 ( .A(n13007), .B(n13009), .Z(n13108) );
  NAND U17423 ( .A(n13109), .B(n13110), .Z(n13009) );
  OR U17424 ( .A(n13111), .B(n13112), .Z(n13110) );
  OR U17425 ( .A(n13113), .B(n13114), .Z(n13109) );
  NAND U17426 ( .A(n13115), .B(n13116), .Z(n13007) );
  OR U17427 ( .A(n13117), .B(n13118), .Z(n13116) );
  OR U17428 ( .A(n13119), .B(n13120), .Z(n13115) );
  ANDN U17429 ( .B(n13121), .A(n13122), .Z(n13008) );
  IV U17430 ( .A(n13123), .Z(n13121) );
  XNOR U17431 ( .A(n13088), .B(n13087), .Z(N29081) );
  XOR U17432 ( .A(n13107), .B(n13106), .Z(n13087) );
  XNOR U17433 ( .A(n13122), .B(n13123), .Z(n13106) );
  XNOR U17434 ( .A(n13117), .B(n13118), .Z(n13123) );
  XNOR U17435 ( .A(n13119), .B(n13120), .Z(n13118) );
  XNOR U17436 ( .A(y[2308]), .B(x[2308]), .Z(n13120) );
  XNOR U17437 ( .A(y[2309]), .B(x[2309]), .Z(n13119) );
  XNOR U17438 ( .A(y[2307]), .B(x[2307]), .Z(n13117) );
  XNOR U17439 ( .A(n13111), .B(n13112), .Z(n13122) );
  XNOR U17440 ( .A(y[2304]), .B(x[2304]), .Z(n13112) );
  XNOR U17441 ( .A(n13113), .B(n13114), .Z(n13111) );
  XNOR U17442 ( .A(y[2305]), .B(x[2305]), .Z(n13114) );
  XNOR U17443 ( .A(y[2306]), .B(x[2306]), .Z(n13113) );
  XNOR U17444 ( .A(n13104), .B(n13103), .Z(n13107) );
  XNOR U17445 ( .A(n13099), .B(n13100), .Z(n13103) );
  XNOR U17446 ( .A(y[2301]), .B(x[2301]), .Z(n13100) );
  XNOR U17447 ( .A(n13101), .B(n13102), .Z(n13099) );
  XNOR U17448 ( .A(y[2302]), .B(x[2302]), .Z(n13102) );
  XNOR U17449 ( .A(y[2303]), .B(x[2303]), .Z(n13101) );
  XNOR U17450 ( .A(n13093), .B(n13094), .Z(n13104) );
  XNOR U17451 ( .A(y[2298]), .B(x[2298]), .Z(n13094) );
  XNOR U17452 ( .A(n13095), .B(n13096), .Z(n13093) );
  XNOR U17453 ( .A(y[2299]), .B(x[2299]), .Z(n13096) );
  XNOR U17454 ( .A(y[2300]), .B(x[2300]), .Z(n13095) );
  XOR U17455 ( .A(n13069), .B(n13070), .Z(n13088) );
  XNOR U17456 ( .A(n13085), .B(n13086), .Z(n13070) );
  XNOR U17457 ( .A(n13080), .B(n13081), .Z(n13086) );
  XNOR U17458 ( .A(n13082), .B(n13083), .Z(n13081) );
  XNOR U17459 ( .A(y[2296]), .B(x[2296]), .Z(n13083) );
  XNOR U17460 ( .A(y[2297]), .B(x[2297]), .Z(n13082) );
  XNOR U17461 ( .A(y[2295]), .B(x[2295]), .Z(n13080) );
  XNOR U17462 ( .A(n13074), .B(n13075), .Z(n13085) );
  XNOR U17463 ( .A(y[2292]), .B(x[2292]), .Z(n13075) );
  XNOR U17464 ( .A(n13076), .B(n13077), .Z(n13074) );
  XNOR U17465 ( .A(y[2293]), .B(x[2293]), .Z(n13077) );
  XNOR U17466 ( .A(y[2294]), .B(x[2294]), .Z(n13076) );
  XOR U17467 ( .A(n13068), .B(n13067), .Z(n13069) );
  XNOR U17468 ( .A(n13063), .B(n13064), .Z(n13067) );
  XNOR U17469 ( .A(y[2289]), .B(x[2289]), .Z(n13064) );
  XNOR U17470 ( .A(n13065), .B(n13066), .Z(n13063) );
  XNOR U17471 ( .A(y[2290]), .B(x[2290]), .Z(n13066) );
  XNOR U17472 ( .A(y[2291]), .B(x[2291]), .Z(n13065) );
  XNOR U17473 ( .A(n13057), .B(n13058), .Z(n13068) );
  XNOR U17474 ( .A(y[2286]), .B(x[2286]), .Z(n13058) );
  XNOR U17475 ( .A(n13059), .B(n13060), .Z(n13057) );
  XNOR U17476 ( .A(y[2287]), .B(x[2287]), .Z(n13060) );
  XNOR U17477 ( .A(y[2288]), .B(x[2288]), .Z(n13059) );
  NAND U17478 ( .A(n13124), .B(n13125), .Z(N29073) );
  NANDN U17479 ( .A(n13126), .B(n13127), .Z(n13125) );
  OR U17480 ( .A(n13128), .B(n13129), .Z(n13127) );
  NAND U17481 ( .A(n13128), .B(n13129), .Z(n13124) );
  XOR U17482 ( .A(n13128), .B(n13130), .Z(N29072) );
  XNOR U17483 ( .A(n13126), .B(n13129), .Z(n13130) );
  AND U17484 ( .A(n13131), .B(n13132), .Z(n13129) );
  NANDN U17485 ( .A(n13133), .B(n13134), .Z(n13132) );
  NANDN U17486 ( .A(n13135), .B(n13136), .Z(n13134) );
  NANDN U17487 ( .A(n13136), .B(n13135), .Z(n13131) );
  NAND U17488 ( .A(n13137), .B(n13138), .Z(n13126) );
  NANDN U17489 ( .A(n13139), .B(n13140), .Z(n13138) );
  OR U17490 ( .A(n13141), .B(n13142), .Z(n13140) );
  NAND U17491 ( .A(n13142), .B(n13141), .Z(n13137) );
  AND U17492 ( .A(n13143), .B(n13144), .Z(n13128) );
  NANDN U17493 ( .A(n13145), .B(n13146), .Z(n13144) );
  NANDN U17494 ( .A(n13147), .B(n13148), .Z(n13146) );
  NANDN U17495 ( .A(n13148), .B(n13147), .Z(n13143) );
  XOR U17496 ( .A(n13142), .B(n13149), .Z(N29071) );
  XOR U17497 ( .A(n13139), .B(n13141), .Z(n13149) );
  XNOR U17498 ( .A(n13135), .B(n13150), .Z(n13141) );
  XNOR U17499 ( .A(n13133), .B(n13136), .Z(n13150) );
  NAND U17500 ( .A(n13151), .B(n13152), .Z(n13136) );
  NAND U17501 ( .A(n13153), .B(n13154), .Z(n13152) );
  OR U17502 ( .A(n13155), .B(n13156), .Z(n13153) );
  NANDN U17503 ( .A(n13157), .B(n13155), .Z(n13151) );
  IV U17504 ( .A(n13156), .Z(n13157) );
  NAND U17505 ( .A(n13158), .B(n13159), .Z(n13133) );
  NAND U17506 ( .A(n13160), .B(n13161), .Z(n13159) );
  NANDN U17507 ( .A(n13162), .B(n13163), .Z(n13160) );
  NANDN U17508 ( .A(n13163), .B(n13162), .Z(n13158) );
  AND U17509 ( .A(n13164), .B(n13165), .Z(n13135) );
  NAND U17510 ( .A(n13166), .B(n13167), .Z(n13165) );
  OR U17511 ( .A(n13168), .B(n13169), .Z(n13166) );
  NANDN U17512 ( .A(n13170), .B(n13168), .Z(n13164) );
  NAND U17513 ( .A(n13171), .B(n13172), .Z(n13139) );
  NANDN U17514 ( .A(n13173), .B(n13174), .Z(n13172) );
  OR U17515 ( .A(n13175), .B(n13176), .Z(n13174) );
  NANDN U17516 ( .A(n13177), .B(n13175), .Z(n13171) );
  IV U17517 ( .A(n13176), .Z(n13177) );
  XNOR U17518 ( .A(n13147), .B(n13178), .Z(n13142) );
  XNOR U17519 ( .A(n13145), .B(n13148), .Z(n13178) );
  NAND U17520 ( .A(n13179), .B(n13180), .Z(n13148) );
  NAND U17521 ( .A(n13181), .B(n13182), .Z(n13180) );
  OR U17522 ( .A(n13183), .B(n13184), .Z(n13181) );
  NANDN U17523 ( .A(n13185), .B(n13183), .Z(n13179) );
  IV U17524 ( .A(n13184), .Z(n13185) );
  NAND U17525 ( .A(n13186), .B(n13187), .Z(n13145) );
  NAND U17526 ( .A(n13188), .B(n13189), .Z(n13187) );
  NANDN U17527 ( .A(n13190), .B(n13191), .Z(n13188) );
  NANDN U17528 ( .A(n13191), .B(n13190), .Z(n13186) );
  AND U17529 ( .A(n13192), .B(n13193), .Z(n13147) );
  NAND U17530 ( .A(n13194), .B(n13195), .Z(n13193) );
  OR U17531 ( .A(n13196), .B(n13197), .Z(n13194) );
  NANDN U17532 ( .A(n13198), .B(n13196), .Z(n13192) );
  XNOR U17533 ( .A(n13173), .B(n13199), .Z(N29070) );
  XOR U17534 ( .A(n13175), .B(n13176), .Z(n13199) );
  XNOR U17535 ( .A(n13189), .B(n13200), .Z(n13176) );
  XOR U17536 ( .A(n13190), .B(n13191), .Z(n13200) );
  XOR U17537 ( .A(n13196), .B(n13201), .Z(n13191) );
  XOR U17538 ( .A(n13195), .B(n13198), .Z(n13201) );
  IV U17539 ( .A(n13197), .Z(n13198) );
  NAND U17540 ( .A(n13202), .B(n13203), .Z(n13197) );
  OR U17541 ( .A(n13204), .B(n13205), .Z(n13203) );
  OR U17542 ( .A(n13206), .B(n13207), .Z(n13202) );
  NAND U17543 ( .A(n13208), .B(n13209), .Z(n13195) );
  OR U17544 ( .A(n13210), .B(n13211), .Z(n13209) );
  OR U17545 ( .A(n13212), .B(n13213), .Z(n13208) );
  NOR U17546 ( .A(n13214), .B(n13215), .Z(n13196) );
  ANDN U17547 ( .B(n13216), .A(n13217), .Z(n13190) );
  XNOR U17548 ( .A(n13183), .B(n13218), .Z(n13189) );
  XNOR U17549 ( .A(n13182), .B(n13184), .Z(n13218) );
  NAND U17550 ( .A(n13219), .B(n13220), .Z(n13184) );
  OR U17551 ( .A(n13221), .B(n13222), .Z(n13220) );
  OR U17552 ( .A(n13223), .B(n13224), .Z(n13219) );
  NAND U17553 ( .A(n13225), .B(n13226), .Z(n13182) );
  OR U17554 ( .A(n13227), .B(n13228), .Z(n13226) );
  OR U17555 ( .A(n13229), .B(n13230), .Z(n13225) );
  ANDN U17556 ( .B(n13231), .A(n13232), .Z(n13183) );
  IV U17557 ( .A(n13233), .Z(n13231) );
  ANDN U17558 ( .B(n13234), .A(n13235), .Z(n13175) );
  XOR U17559 ( .A(n13161), .B(n13236), .Z(n13173) );
  XOR U17560 ( .A(n13162), .B(n13163), .Z(n13236) );
  XOR U17561 ( .A(n13168), .B(n13237), .Z(n13163) );
  XOR U17562 ( .A(n13167), .B(n13170), .Z(n13237) );
  IV U17563 ( .A(n13169), .Z(n13170) );
  NAND U17564 ( .A(n13238), .B(n13239), .Z(n13169) );
  OR U17565 ( .A(n13240), .B(n13241), .Z(n13239) );
  OR U17566 ( .A(n13242), .B(n13243), .Z(n13238) );
  NAND U17567 ( .A(n13244), .B(n13245), .Z(n13167) );
  OR U17568 ( .A(n13246), .B(n13247), .Z(n13245) );
  OR U17569 ( .A(n13248), .B(n13249), .Z(n13244) );
  NOR U17570 ( .A(n13250), .B(n13251), .Z(n13168) );
  ANDN U17571 ( .B(n13252), .A(n13253), .Z(n13162) );
  IV U17572 ( .A(n13254), .Z(n13252) );
  XNOR U17573 ( .A(n13155), .B(n13255), .Z(n13161) );
  XNOR U17574 ( .A(n13154), .B(n13156), .Z(n13255) );
  NAND U17575 ( .A(n13256), .B(n13257), .Z(n13156) );
  OR U17576 ( .A(n13258), .B(n13259), .Z(n13257) );
  OR U17577 ( .A(n13260), .B(n13261), .Z(n13256) );
  NAND U17578 ( .A(n13262), .B(n13263), .Z(n13154) );
  OR U17579 ( .A(n13264), .B(n13265), .Z(n13263) );
  OR U17580 ( .A(n13266), .B(n13267), .Z(n13262) );
  ANDN U17581 ( .B(n13268), .A(n13269), .Z(n13155) );
  IV U17582 ( .A(n13270), .Z(n13268) );
  XNOR U17583 ( .A(n13235), .B(n13234), .Z(N29069) );
  XOR U17584 ( .A(n13254), .B(n13253), .Z(n13234) );
  XNOR U17585 ( .A(n13269), .B(n13270), .Z(n13253) );
  XNOR U17586 ( .A(n13264), .B(n13265), .Z(n13270) );
  XNOR U17587 ( .A(n13266), .B(n13267), .Z(n13265) );
  XNOR U17588 ( .A(y[2284]), .B(x[2284]), .Z(n13267) );
  XNOR U17589 ( .A(y[2285]), .B(x[2285]), .Z(n13266) );
  XNOR U17590 ( .A(y[2283]), .B(x[2283]), .Z(n13264) );
  XNOR U17591 ( .A(n13258), .B(n13259), .Z(n13269) );
  XNOR U17592 ( .A(y[2280]), .B(x[2280]), .Z(n13259) );
  XNOR U17593 ( .A(n13260), .B(n13261), .Z(n13258) );
  XNOR U17594 ( .A(y[2281]), .B(x[2281]), .Z(n13261) );
  XNOR U17595 ( .A(y[2282]), .B(x[2282]), .Z(n13260) );
  XNOR U17596 ( .A(n13251), .B(n13250), .Z(n13254) );
  XNOR U17597 ( .A(n13246), .B(n13247), .Z(n13250) );
  XNOR U17598 ( .A(y[2277]), .B(x[2277]), .Z(n13247) );
  XNOR U17599 ( .A(n13248), .B(n13249), .Z(n13246) );
  XNOR U17600 ( .A(y[2278]), .B(x[2278]), .Z(n13249) );
  XNOR U17601 ( .A(y[2279]), .B(x[2279]), .Z(n13248) );
  XNOR U17602 ( .A(n13240), .B(n13241), .Z(n13251) );
  XNOR U17603 ( .A(y[2274]), .B(x[2274]), .Z(n13241) );
  XNOR U17604 ( .A(n13242), .B(n13243), .Z(n13240) );
  XNOR U17605 ( .A(y[2275]), .B(x[2275]), .Z(n13243) );
  XNOR U17606 ( .A(y[2276]), .B(x[2276]), .Z(n13242) );
  XOR U17607 ( .A(n13216), .B(n13217), .Z(n13235) );
  XNOR U17608 ( .A(n13232), .B(n13233), .Z(n13217) );
  XNOR U17609 ( .A(n13227), .B(n13228), .Z(n13233) );
  XNOR U17610 ( .A(n13229), .B(n13230), .Z(n13228) );
  XNOR U17611 ( .A(y[2272]), .B(x[2272]), .Z(n13230) );
  XNOR U17612 ( .A(y[2273]), .B(x[2273]), .Z(n13229) );
  XNOR U17613 ( .A(y[2271]), .B(x[2271]), .Z(n13227) );
  XNOR U17614 ( .A(n13221), .B(n13222), .Z(n13232) );
  XNOR U17615 ( .A(y[2268]), .B(x[2268]), .Z(n13222) );
  XNOR U17616 ( .A(n13223), .B(n13224), .Z(n13221) );
  XNOR U17617 ( .A(y[2269]), .B(x[2269]), .Z(n13224) );
  XNOR U17618 ( .A(y[2270]), .B(x[2270]), .Z(n13223) );
  XOR U17619 ( .A(n13215), .B(n13214), .Z(n13216) );
  XNOR U17620 ( .A(n13210), .B(n13211), .Z(n13214) );
  XNOR U17621 ( .A(y[2265]), .B(x[2265]), .Z(n13211) );
  XNOR U17622 ( .A(n13212), .B(n13213), .Z(n13210) );
  XNOR U17623 ( .A(y[2266]), .B(x[2266]), .Z(n13213) );
  XNOR U17624 ( .A(y[2267]), .B(x[2267]), .Z(n13212) );
  XNOR U17625 ( .A(n13204), .B(n13205), .Z(n13215) );
  XNOR U17626 ( .A(y[2262]), .B(x[2262]), .Z(n13205) );
  XNOR U17627 ( .A(n13206), .B(n13207), .Z(n13204) );
  XNOR U17628 ( .A(y[2263]), .B(x[2263]), .Z(n13207) );
  XNOR U17629 ( .A(y[2264]), .B(x[2264]), .Z(n13206) );
  NAND U17630 ( .A(n13271), .B(n13272), .Z(N29061) );
  NANDN U17631 ( .A(n13273), .B(n13274), .Z(n13272) );
  OR U17632 ( .A(n13275), .B(n13276), .Z(n13274) );
  NAND U17633 ( .A(n13275), .B(n13276), .Z(n13271) );
  XOR U17634 ( .A(n13275), .B(n13277), .Z(N29060) );
  XNOR U17635 ( .A(n13273), .B(n13276), .Z(n13277) );
  AND U17636 ( .A(n13278), .B(n13279), .Z(n13276) );
  NANDN U17637 ( .A(n13280), .B(n13281), .Z(n13279) );
  NANDN U17638 ( .A(n13282), .B(n13283), .Z(n13281) );
  NANDN U17639 ( .A(n13283), .B(n13282), .Z(n13278) );
  NAND U17640 ( .A(n13284), .B(n13285), .Z(n13273) );
  NANDN U17641 ( .A(n13286), .B(n13287), .Z(n13285) );
  OR U17642 ( .A(n13288), .B(n13289), .Z(n13287) );
  NAND U17643 ( .A(n13289), .B(n13288), .Z(n13284) );
  AND U17644 ( .A(n13290), .B(n13291), .Z(n13275) );
  NANDN U17645 ( .A(n13292), .B(n13293), .Z(n13291) );
  NANDN U17646 ( .A(n13294), .B(n13295), .Z(n13293) );
  NANDN U17647 ( .A(n13295), .B(n13294), .Z(n13290) );
  XOR U17648 ( .A(n13289), .B(n13296), .Z(N29059) );
  XOR U17649 ( .A(n13286), .B(n13288), .Z(n13296) );
  XNOR U17650 ( .A(n13282), .B(n13297), .Z(n13288) );
  XNOR U17651 ( .A(n13280), .B(n13283), .Z(n13297) );
  NAND U17652 ( .A(n13298), .B(n13299), .Z(n13283) );
  NAND U17653 ( .A(n13300), .B(n13301), .Z(n13299) );
  OR U17654 ( .A(n13302), .B(n13303), .Z(n13300) );
  NANDN U17655 ( .A(n13304), .B(n13302), .Z(n13298) );
  IV U17656 ( .A(n13303), .Z(n13304) );
  NAND U17657 ( .A(n13305), .B(n13306), .Z(n13280) );
  NAND U17658 ( .A(n13307), .B(n13308), .Z(n13306) );
  NANDN U17659 ( .A(n13309), .B(n13310), .Z(n13307) );
  NANDN U17660 ( .A(n13310), .B(n13309), .Z(n13305) );
  AND U17661 ( .A(n13311), .B(n13312), .Z(n13282) );
  NAND U17662 ( .A(n13313), .B(n13314), .Z(n13312) );
  OR U17663 ( .A(n13315), .B(n13316), .Z(n13313) );
  NANDN U17664 ( .A(n13317), .B(n13315), .Z(n13311) );
  NAND U17665 ( .A(n13318), .B(n13319), .Z(n13286) );
  NANDN U17666 ( .A(n13320), .B(n13321), .Z(n13319) );
  OR U17667 ( .A(n13322), .B(n13323), .Z(n13321) );
  NANDN U17668 ( .A(n13324), .B(n13322), .Z(n13318) );
  IV U17669 ( .A(n13323), .Z(n13324) );
  XNOR U17670 ( .A(n13294), .B(n13325), .Z(n13289) );
  XNOR U17671 ( .A(n13292), .B(n13295), .Z(n13325) );
  NAND U17672 ( .A(n13326), .B(n13327), .Z(n13295) );
  NAND U17673 ( .A(n13328), .B(n13329), .Z(n13327) );
  OR U17674 ( .A(n13330), .B(n13331), .Z(n13328) );
  NANDN U17675 ( .A(n13332), .B(n13330), .Z(n13326) );
  IV U17676 ( .A(n13331), .Z(n13332) );
  NAND U17677 ( .A(n13333), .B(n13334), .Z(n13292) );
  NAND U17678 ( .A(n13335), .B(n13336), .Z(n13334) );
  NANDN U17679 ( .A(n13337), .B(n13338), .Z(n13335) );
  NANDN U17680 ( .A(n13338), .B(n13337), .Z(n13333) );
  AND U17681 ( .A(n13339), .B(n13340), .Z(n13294) );
  NAND U17682 ( .A(n13341), .B(n13342), .Z(n13340) );
  OR U17683 ( .A(n13343), .B(n13344), .Z(n13341) );
  NANDN U17684 ( .A(n13345), .B(n13343), .Z(n13339) );
  XNOR U17685 ( .A(n13320), .B(n13346), .Z(N29058) );
  XOR U17686 ( .A(n13322), .B(n13323), .Z(n13346) );
  XNOR U17687 ( .A(n13336), .B(n13347), .Z(n13323) );
  XOR U17688 ( .A(n13337), .B(n13338), .Z(n13347) );
  XOR U17689 ( .A(n13343), .B(n13348), .Z(n13338) );
  XOR U17690 ( .A(n13342), .B(n13345), .Z(n13348) );
  IV U17691 ( .A(n13344), .Z(n13345) );
  NAND U17692 ( .A(n13349), .B(n13350), .Z(n13344) );
  OR U17693 ( .A(n13351), .B(n13352), .Z(n13350) );
  OR U17694 ( .A(n13353), .B(n13354), .Z(n13349) );
  NAND U17695 ( .A(n13355), .B(n13356), .Z(n13342) );
  OR U17696 ( .A(n13357), .B(n13358), .Z(n13356) );
  OR U17697 ( .A(n13359), .B(n13360), .Z(n13355) );
  NOR U17698 ( .A(n13361), .B(n13362), .Z(n13343) );
  ANDN U17699 ( .B(n13363), .A(n13364), .Z(n13337) );
  XNOR U17700 ( .A(n13330), .B(n13365), .Z(n13336) );
  XNOR U17701 ( .A(n13329), .B(n13331), .Z(n13365) );
  NAND U17702 ( .A(n13366), .B(n13367), .Z(n13331) );
  OR U17703 ( .A(n13368), .B(n13369), .Z(n13367) );
  OR U17704 ( .A(n13370), .B(n13371), .Z(n13366) );
  NAND U17705 ( .A(n13372), .B(n13373), .Z(n13329) );
  OR U17706 ( .A(n13374), .B(n13375), .Z(n13373) );
  OR U17707 ( .A(n13376), .B(n13377), .Z(n13372) );
  ANDN U17708 ( .B(n13378), .A(n13379), .Z(n13330) );
  IV U17709 ( .A(n13380), .Z(n13378) );
  ANDN U17710 ( .B(n13381), .A(n13382), .Z(n13322) );
  XOR U17711 ( .A(n13308), .B(n13383), .Z(n13320) );
  XOR U17712 ( .A(n13309), .B(n13310), .Z(n13383) );
  XOR U17713 ( .A(n13315), .B(n13384), .Z(n13310) );
  XOR U17714 ( .A(n13314), .B(n13317), .Z(n13384) );
  IV U17715 ( .A(n13316), .Z(n13317) );
  NAND U17716 ( .A(n13385), .B(n13386), .Z(n13316) );
  OR U17717 ( .A(n13387), .B(n13388), .Z(n13386) );
  OR U17718 ( .A(n13389), .B(n13390), .Z(n13385) );
  NAND U17719 ( .A(n13391), .B(n13392), .Z(n13314) );
  OR U17720 ( .A(n13393), .B(n13394), .Z(n13392) );
  OR U17721 ( .A(n13395), .B(n13396), .Z(n13391) );
  NOR U17722 ( .A(n13397), .B(n13398), .Z(n13315) );
  ANDN U17723 ( .B(n13399), .A(n13400), .Z(n13309) );
  IV U17724 ( .A(n13401), .Z(n13399) );
  XNOR U17725 ( .A(n13302), .B(n13402), .Z(n13308) );
  XNOR U17726 ( .A(n13301), .B(n13303), .Z(n13402) );
  NAND U17727 ( .A(n13403), .B(n13404), .Z(n13303) );
  OR U17728 ( .A(n13405), .B(n13406), .Z(n13404) );
  OR U17729 ( .A(n13407), .B(n13408), .Z(n13403) );
  NAND U17730 ( .A(n13409), .B(n13410), .Z(n13301) );
  OR U17731 ( .A(n13411), .B(n13412), .Z(n13410) );
  OR U17732 ( .A(n13413), .B(n13414), .Z(n13409) );
  ANDN U17733 ( .B(n13415), .A(n13416), .Z(n13302) );
  IV U17734 ( .A(n13417), .Z(n13415) );
  XNOR U17735 ( .A(n13382), .B(n13381), .Z(N29057) );
  XOR U17736 ( .A(n13401), .B(n13400), .Z(n13381) );
  XNOR U17737 ( .A(n13416), .B(n13417), .Z(n13400) );
  XNOR U17738 ( .A(n13411), .B(n13412), .Z(n13417) );
  XNOR U17739 ( .A(n13413), .B(n13414), .Z(n13412) );
  XNOR U17740 ( .A(y[2260]), .B(x[2260]), .Z(n13414) );
  XNOR U17741 ( .A(y[2261]), .B(x[2261]), .Z(n13413) );
  XNOR U17742 ( .A(y[2259]), .B(x[2259]), .Z(n13411) );
  XNOR U17743 ( .A(n13405), .B(n13406), .Z(n13416) );
  XNOR U17744 ( .A(y[2256]), .B(x[2256]), .Z(n13406) );
  XNOR U17745 ( .A(n13407), .B(n13408), .Z(n13405) );
  XNOR U17746 ( .A(y[2257]), .B(x[2257]), .Z(n13408) );
  XNOR U17747 ( .A(y[2258]), .B(x[2258]), .Z(n13407) );
  XNOR U17748 ( .A(n13398), .B(n13397), .Z(n13401) );
  XNOR U17749 ( .A(n13393), .B(n13394), .Z(n13397) );
  XNOR U17750 ( .A(y[2253]), .B(x[2253]), .Z(n13394) );
  XNOR U17751 ( .A(n13395), .B(n13396), .Z(n13393) );
  XNOR U17752 ( .A(y[2254]), .B(x[2254]), .Z(n13396) );
  XNOR U17753 ( .A(y[2255]), .B(x[2255]), .Z(n13395) );
  XNOR U17754 ( .A(n13387), .B(n13388), .Z(n13398) );
  XNOR U17755 ( .A(y[2250]), .B(x[2250]), .Z(n13388) );
  XNOR U17756 ( .A(n13389), .B(n13390), .Z(n13387) );
  XNOR U17757 ( .A(y[2251]), .B(x[2251]), .Z(n13390) );
  XNOR U17758 ( .A(y[2252]), .B(x[2252]), .Z(n13389) );
  XOR U17759 ( .A(n13363), .B(n13364), .Z(n13382) );
  XNOR U17760 ( .A(n13379), .B(n13380), .Z(n13364) );
  XNOR U17761 ( .A(n13374), .B(n13375), .Z(n13380) );
  XNOR U17762 ( .A(n13376), .B(n13377), .Z(n13375) );
  XNOR U17763 ( .A(y[2248]), .B(x[2248]), .Z(n13377) );
  XNOR U17764 ( .A(y[2249]), .B(x[2249]), .Z(n13376) );
  XNOR U17765 ( .A(y[2247]), .B(x[2247]), .Z(n13374) );
  XNOR U17766 ( .A(n13368), .B(n13369), .Z(n13379) );
  XNOR U17767 ( .A(y[2244]), .B(x[2244]), .Z(n13369) );
  XNOR U17768 ( .A(n13370), .B(n13371), .Z(n13368) );
  XNOR U17769 ( .A(y[2245]), .B(x[2245]), .Z(n13371) );
  XNOR U17770 ( .A(y[2246]), .B(x[2246]), .Z(n13370) );
  XOR U17771 ( .A(n13362), .B(n13361), .Z(n13363) );
  XNOR U17772 ( .A(n13357), .B(n13358), .Z(n13361) );
  XNOR U17773 ( .A(y[2241]), .B(x[2241]), .Z(n13358) );
  XNOR U17774 ( .A(n13359), .B(n13360), .Z(n13357) );
  XNOR U17775 ( .A(y[2242]), .B(x[2242]), .Z(n13360) );
  XNOR U17776 ( .A(y[2243]), .B(x[2243]), .Z(n13359) );
  XNOR U17777 ( .A(n13351), .B(n13352), .Z(n13362) );
  XNOR U17778 ( .A(y[2238]), .B(x[2238]), .Z(n13352) );
  XNOR U17779 ( .A(n13353), .B(n13354), .Z(n13351) );
  XNOR U17780 ( .A(y[2239]), .B(x[2239]), .Z(n13354) );
  XNOR U17781 ( .A(y[2240]), .B(x[2240]), .Z(n13353) );
  NAND U17782 ( .A(n13418), .B(n13419), .Z(N29049) );
  NANDN U17783 ( .A(n13420), .B(n13421), .Z(n13419) );
  OR U17784 ( .A(n13422), .B(n13423), .Z(n13421) );
  NAND U17785 ( .A(n13422), .B(n13423), .Z(n13418) );
  XOR U17786 ( .A(n13422), .B(n13424), .Z(N29048) );
  XNOR U17787 ( .A(n13420), .B(n13423), .Z(n13424) );
  AND U17788 ( .A(n13425), .B(n13426), .Z(n13423) );
  NANDN U17789 ( .A(n13427), .B(n13428), .Z(n13426) );
  NANDN U17790 ( .A(n13429), .B(n13430), .Z(n13428) );
  NANDN U17791 ( .A(n13430), .B(n13429), .Z(n13425) );
  NAND U17792 ( .A(n13431), .B(n13432), .Z(n13420) );
  NANDN U17793 ( .A(n13433), .B(n13434), .Z(n13432) );
  OR U17794 ( .A(n13435), .B(n13436), .Z(n13434) );
  NAND U17795 ( .A(n13436), .B(n13435), .Z(n13431) );
  AND U17796 ( .A(n13437), .B(n13438), .Z(n13422) );
  NANDN U17797 ( .A(n13439), .B(n13440), .Z(n13438) );
  NANDN U17798 ( .A(n13441), .B(n13442), .Z(n13440) );
  NANDN U17799 ( .A(n13442), .B(n13441), .Z(n13437) );
  XOR U17800 ( .A(n13436), .B(n13443), .Z(N29047) );
  XOR U17801 ( .A(n13433), .B(n13435), .Z(n13443) );
  XNOR U17802 ( .A(n13429), .B(n13444), .Z(n13435) );
  XNOR U17803 ( .A(n13427), .B(n13430), .Z(n13444) );
  NAND U17804 ( .A(n13445), .B(n13446), .Z(n13430) );
  NAND U17805 ( .A(n13447), .B(n13448), .Z(n13446) );
  OR U17806 ( .A(n13449), .B(n13450), .Z(n13447) );
  NANDN U17807 ( .A(n13451), .B(n13449), .Z(n13445) );
  IV U17808 ( .A(n13450), .Z(n13451) );
  NAND U17809 ( .A(n13452), .B(n13453), .Z(n13427) );
  NAND U17810 ( .A(n13454), .B(n13455), .Z(n13453) );
  NANDN U17811 ( .A(n13456), .B(n13457), .Z(n13454) );
  NANDN U17812 ( .A(n13457), .B(n13456), .Z(n13452) );
  AND U17813 ( .A(n13458), .B(n13459), .Z(n13429) );
  NAND U17814 ( .A(n13460), .B(n13461), .Z(n13459) );
  OR U17815 ( .A(n13462), .B(n13463), .Z(n13460) );
  NANDN U17816 ( .A(n13464), .B(n13462), .Z(n13458) );
  NAND U17817 ( .A(n13465), .B(n13466), .Z(n13433) );
  NANDN U17818 ( .A(n13467), .B(n13468), .Z(n13466) );
  OR U17819 ( .A(n13469), .B(n13470), .Z(n13468) );
  NANDN U17820 ( .A(n13471), .B(n13469), .Z(n13465) );
  IV U17821 ( .A(n13470), .Z(n13471) );
  XNOR U17822 ( .A(n13441), .B(n13472), .Z(n13436) );
  XNOR U17823 ( .A(n13439), .B(n13442), .Z(n13472) );
  NAND U17824 ( .A(n13473), .B(n13474), .Z(n13442) );
  NAND U17825 ( .A(n13475), .B(n13476), .Z(n13474) );
  OR U17826 ( .A(n13477), .B(n13478), .Z(n13475) );
  NANDN U17827 ( .A(n13479), .B(n13477), .Z(n13473) );
  IV U17828 ( .A(n13478), .Z(n13479) );
  NAND U17829 ( .A(n13480), .B(n13481), .Z(n13439) );
  NAND U17830 ( .A(n13482), .B(n13483), .Z(n13481) );
  NANDN U17831 ( .A(n13484), .B(n13485), .Z(n13482) );
  NANDN U17832 ( .A(n13485), .B(n13484), .Z(n13480) );
  AND U17833 ( .A(n13486), .B(n13487), .Z(n13441) );
  NAND U17834 ( .A(n13488), .B(n13489), .Z(n13487) );
  OR U17835 ( .A(n13490), .B(n13491), .Z(n13488) );
  NANDN U17836 ( .A(n13492), .B(n13490), .Z(n13486) );
  XNOR U17837 ( .A(n13467), .B(n13493), .Z(N29046) );
  XOR U17838 ( .A(n13469), .B(n13470), .Z(n13493) );
  XNOR U17839 ( .A(n13483), .B(n13494), .Z(n13470) );
  XOR U17840 ( .A(n13484), .B(n13485), .Z(n13494) );
  XOR U17841 ( .A(n13490), .B(n13495), .Z(n13485) );
  XOR U17842 ( .A(n13489), .B(n13492), .Z(n13495) );
  IV U17843 ( .A(n13491), .Z(n13492) );
  NAND U17844 ( .A(n13496), .B(n13497), .Z(n13491) );
  OR U17845 ( .A(n13498), .B(n13499), .Z(n13497) );
  OR U17846 ( .A(n13500), .B(n13501), .Z(n13496) );
  NAND U17847 ( .A(n13502), .B(n13503), .Z(n13489) );
  OR U17848 ( .A(n13504), .B(n13505), .Z(n13503) );
  OR U17849 ( .A(n13506), .B(n13507), .Z(n13502) );
  NOR U17850 ( .A(n13508), .B(n13509), .Z(n13490) );
  ANDN U17851 ( .B(n13510), .A(n13511), .Z(n13484) );
  XNOR U17852 ( .A(n13477), .B(n13512), .Z(n13483) );
  XNOR U17853 ( .A(n13476), .B(n13478), .Z(n13512) );
  NAND U17854 ( .A(n13513), .B(n13514), .Z(n13478) );
  OR U17855 ( .A(n13515), .B(n13516), .Z(n13514) );
  OR U17856 ( .A(n13517), .B(n13518), .Z(n13513) );
  NAND U17857 ( .A(n13519), .B(n13520), .Z(n13476) );
  OR U17858 ( .A(n13521), .B(n13522), .Z(n13520) );
  OR U17859 ( .A(n13523), .B(n13524), .Z(n13519) );
  ANDN U17860 ( .B(n13525), .A(n13526), .Z(n13477) );
  IV U17861 ( .A(n13527), .Z(n13525) );
  ANDN U17862 ( .B(n13528), .A(n13529), .Z(n13469) );
  XOR U17863 ( .A(n13455), .B(n13530), .Z(n13467) );
  XOR U17864 ( .A(n13456), .B(n13457), .Z(n13530) );
  XOR U17865 ( .A(n13462), .B(n13531), .Z(n13457) );
  XOR U17866 ( .A(n13461), .B(n13464), .Z(n13531) );
  IV U17867 ( .A(n13463), .Z(n13464) );
  NAND U17868 ( .A(n13532), .B(n13533), .Z(n13463) );
  OR U17869 ( .A(n13534), .B(n13535), .Z(n13533) );
  OR U17870 ( .A(n13536), .B(n13537), .Z(n13532) );
  NAND U17871 ( .A(n13538), .B(n13539), .Z(n13461) );
  OR U17872 ( .A(n13540), .B(n13541), .Z(n13539) );
  OR U17873 ( .A(n13542), .B(n13543), .Z(n13538) );
  NOR U17874 ( .A(n13544), .B(n13545), .Z(n13462) );
  ANDN U17875 ( .B(n13546), .A(n13547), .Z(n13456) );
  IV U17876 ( .A(n13548), .Z(n13546) );
  XNOR U17877 ( .A(n13449), .B(n13549), .Z(n13455) );
  XNOR U17878 ( .A(n13448), .B(n13450), .Z(n13549) );
  NAND U17879 ( .A(n13550), .B(n13551), .Z(n13450) );
  OR U17880 ( .A(n13552), .B(n13553), .Z(n13551) );
  OR U17881 ( .A(n13554), .B(n13555), .Z(n13550) );
  NAND U17882 ( .A(n13556), .B(n13557), .Z(n13448) );
  OR U17883 ( .A(n13558), .B(n13559), .Z(n13557) );
  OR U17884 ( .A(n13560), .B(n13561), .Z(n13556) );
  ANDN U17885 ( .B(n13562), .A(n13563), .Z(n13449) );
  IV U17886 ( .A(n13564), .Z(n13562) );
  XNOR U17887 ( .A(n13529), .B(n13528), .Z(N29045) );
  XOR U17888 ( .A(n13548), .B(n13547), .Z(n13528) );
  XNOR U17889 ( .A(n13563), .B(n13564), .Z(n13547) );
  XNOR U17890 ( .A(n13558), .B(n13559), .Z(n13564) );
  XNOR U17891 ( .A(n13560), .B(n13561), .Z(n13559) );
  XNOR U17892 ( .A(y[2236]), .B(x[2236]), .Z(n13561) );
  XNOR U17893 ( .A(y[2237]), .B(x[2237]), .Z(n13560) );
  XNOR U17894 ( .A(y[2235]), .B(x[2235]), .Z(n13558) );
  XNOR U17895 ( .A(n13552), .B(n13553), .Z(n13563) );
  XNOR U17896 ( .A(y[2232]), .B(x[2232]), .Z(n13553) );
  XNOR U17897 ( .A(n13554), .B(n13555), .Z(n13552) );
  XNOR U17898 ( .A(y[2233]), .B(x[2233]), .Z(n13555) );
  XNOR U17899 ( .A(y[2234]), .B(x[2234]), .Z(n13554) );
  XNOR U17900 ( .A(n13545), .B(n13544), .Z(n13548) );
  XNOR U17901 ( .A(n13540), .B(n13541), .Z(n13544) );
  XNOR U17902 ( .A(y[2229]), .B(x[2229]), .Z(n13541) );
  XNOR U17903 ( .A(n13542), .B(n13543), .Z(n13540) );
  XNOR U17904 ( .A(y[2230]), .B(x[2230]), .Z(n13543) );
  XNOR U17905 ( .A(y[2231]), .B(x[2231]), .Z(n13542) );
  XNOR U17906 ( .A(n13534), .B(n13535), .Z(n13545) );
  XNOR U17907 ( .A(y[2226]), .B(x[2226]), .Z(n13535) );
  XNOR U17908 ( .A(n13536), .B(n13537), .Z(n13534) );
  XNOR U17909 ( .A(y[2227]), .B(x[2227]), .Z(n13537) );
  XNOR U17910 ( .A(y[2228]), .B(x[2228]), .Z(n13536) );
  XOR U17911 ( .A(n13510), .B(n13511), .Z(n13529) );
  XNOR U17912 ( .A(n13526), .B(n13527), .Z(n13511) );
  XNOR U17913 ( .A(n13521), .B(n13522), .Z(n13527) );
  XNOR U17914 ( .A(n13523), .B(n13524), .Z(n13522) );
  XNOR U17915 ( .A(y[2224]), .B(x[2224]), .Z(n13524) );
  XNOR U17916 ( .A(y[2225]), .B(x[2225]), .Z(n13523) );
  XNOR U17917 ( .A(y[2223]), .B(x[2223]), .Z(n13521) );
  XNOR U17918 ( .A(n13515), .B(n13516), .Z(n13526) );
  XNOR U17919 ( .A(y[2220]), .B(x[2220]), .Z(n13516) );
  XNOR U17920 ( .A(n13517), .B(n13518), .Z(n13515) );
  XNOR U17921 ( .A(y[2221]), .B(x[2221]), .Z(n13518) );
  XNOR U17922 ( .A(y[2222]), .B(x[2222]), .Z(n13517) );
  XOR U17923 ( .A(n13509), .B(n13508), .Z(n13510) );
  XNOR U17924 ( .A(n13504), .B(n13505), .Z(n13508) );
  XNOR U17925 ( .A(y[2217]), .B(x[2217]), .Z(n13505) );
  XNOR U17926 ( .A(n13506), .B(n13507), .Z(n13504) );
  XNOR U17927 ( .A(y[2218]), .B(x[2218]), .Z(n13507) );
  XNOR U17928 ( .A(y[2219]), .B(x[2219]), .Z(n13506) );
  XNOR U17929 ( .A(n13498), .B(n13499), .Z(n13509) );
  XNOR U17930 ( .A(y[2214]), .B(x[2214]), .Z(n13499) );
  XNOR U17931 ( .A(n13500), .B(n13501), .Z(n13498) );
  XNOR U17932 ( .A(y[2215]), .B(x[2215]), .Z(n13501) );
  XNOR U17933 ( .A(y[2216]), .B(x[2216]), .Z(n13500) );
  NAND U17934 ( .A(n13565), .B(n13566), .Z(N29037) );
  NANDN U17935 ( .A(n13567), .B(n13568), .Z(n13566) );
  OR U17936 ( .A(n13569), .B(n13570), .Z(n13568) );
  NAND U17937 ( .A(n13569), .B(n13570), .Z(n13565) );
  XOR U17938 ( .A(n13569), .B(n13571), .Z(N29036) );
  XNOR U17939 ( .A(n13567), .B(n13570), .Z(n13571) );
  AND U17940 ( .A(n13572), .B(n13573), .Z(n13570) );
  NANDN U17941 ( .A(n13574), .B(n13575), .Z(n13573) );
  NANDN U17942 ( .A(n13576), .B(n13577), .Z(n13575) );
  NANDN U17943 ( .A(n13577), .B(n13576), .Z(n13572) );
  NAND U17944 ( .A(n13578), .B(n13579), .Z(n13567) );
  NANDN U17945 ( .A(n13580), .B(n13581), .Z(n13579) );
  OR U17946 ( .A(n13582), .B(n13583), .Z(n13581) );
  NAND U17947 ( .A(n13583), .B(n13582), .Z(n13578) );
  AND U17948 ( .A(n13584), .B(n13585), .Z(n13569) );
  NANDN U17949 ( .A(n13586), .B(n13587), .Z(n13585) );
  NANDN U17950 ( .A(n13588), .B(n13589), .Z(n13587) );
  NANDN U17951 ( .A(n13589), .B(n13588), .Z(n13584) );
  XOR U17952 ( .A(n13583), .B(n13590), .Z(N29035) );
  XOR U17953 ( .A(n13580), .B(n13582), .Z(n13590) );
  XNOR U17954 ( .A(n13576), .B(n13591), .Z(n13582) );
  XNOR U17955 ( .A(n13574), .B(n13577), .Z(n13591) );
  NAND U17956 ( .A(n13592), .B(n13593), .Z(n13577) );
  NAND U17957 ( .A(n13594), .B(n13595), .Z(n13593) );
  OR U17958 ( .A(n13596), .B(n13597), .Z(n13594) );
  NANDN U17959 ( .A(n13598), .B(n13596), .Z(n13592) );
  IV U17960 ( .A(n13597), .Z(n13598) );
  NAND U17961 ( .A(n13599), .B(n13600), .Z(n13574) );
  NAND U17962 ( .A(n13601), .B(n13602), .Z(n13600) );
  NANDN U17963 ( .A(n13603), .B(n13604), .Z(n13601) );
  NANDN U17964 ( .A(n13604), .B(n13603), .Z(n13599) );
  AND U17965 ( .A(n13605), .B(n13606), .Z(n13576) );
  NAND U17966 ( .A(n13607), .B(n13608), .Z(n13606) );
  OR U17967 ( .A(n13609), .B(n13610), .Z(n13607) );
  NANDN U17968 ( .A(n13611), .B(n13609), .Z(n13605) );
  NAND U17969 ( .A(n13612), .B(n13613), .Z(n13580) );
  NANDN U17970 ( .A(n13614), .B(n13615), .Z(n13613) );
  OR U17971 ( .A(n13616), .B(n13617), .Z(n13615) );
  NANDN U17972 ( .A(n13618), .B(n13616), .Z(n13612) );
  IV U17973 ( .A(n13617), .Z(n13618) );
  XNOR U17974 ( .A(n13588), .B(n13619), .Z(n13583) );
  XNOR U17975 ( .A(n13586), .B(n13589), .Z(n13619) );
  NAND U17976 ( .A(n13620), .B(n13621), .Z(n13589) );
  NAND U17977 ( .A(n13622), .B(n13623), .Z(n13621) );
  OR U17978 ( .A(n13624), .B(n13625), .Z(n13622) );
  NANDN U17979 ( .A(n13626), .B(n13624), .Z(n13620) );
  IV U17980 ( .A(n13625), .Z(n13626) );
  NAND U17981 ( .A(n13627), .B(n13628), .Z(n13586) );
  NAND U17982 ( .A(n13629), .B(n13630), .Z(n13628) );
  NANDN U17983 ( .A(n13631), .B(n13632), .Z(n13629) );
  NANDN U17984 ( .A(n13632), .B(n13631), .Z(n13627) );
  AND U17985 ( .A(n13633), .B(n13634), .Z(n13588) );
  NAND U17986 ( .A(n13635), .B(n13636), .Z(n13634) );
  OR U17987 ( .A(n13637), .B(n13638), .Z(n13635) );
  NANDN U17988 ( .A(n13639), .B(n13637), .Z(n13633) );
  XNOR U17989 ( .A(n13614), .B(n13640), .Z(N29034) );
  XOR U17990 ( .A(n13616), .B(n13617), .Z(n13640) );
  XNOR U17991 ( .A(n13630), .B(n13641), .Z(n13617) );
  XOR U17992 ( .A(n13631), .B(n13632), .Z(n13641) );
  XOR U17993 ( .A(n13637), .B(n13642), .Z(n13632) );
  XOR U17994 ( .A(n13636), .B(n13639), .Z(n13642) );
  IV U17995 ( .A(n13638), .Z(n13639) );
  NAND U17996 ( .A(n13643), .B(n13644), .Z(n13638) );
  OR U17997 ( .A(n13645), .B(n13646), .Z(n13644) );
  OR U17998 ( .A(n13647), .B(n13648), .Z(n13643) );
  NAND U17999 ( .A(n13649), .B(n13650), .Z(n13636) );
  OR U18000 ( .A(n13651), .B(n13652), .Z(n13650) );
  OR U18001 ( .A(n13653), .B(n13654), .Z(n13649) );
  NOR U18002 ( .A(n13655), .B(n13656), .Z(n13637) );
  ANDN U18003 ( .B(n13657), .A(n13658), .Z(n13631) );
  XNOR U18004 ( .A(n13624), .B(n13659), .Z(n13630) );
  XNOR U18005 ( .A(n13623), .B(n13625), .Z(n13659) );
  NAND U18006 ( .A(n13660), .B(n13661), .Z(n13625) );
  OR U18007 ( .A(n13662), .B(n13663), .Z(n13661) );
  OR U18008 ( .A(n13664), .B(n13665), .Z(n13660) );
  NAND U18009 ( .A(n13666), .B(n13667), .Z(n13623) );
  OR U18010 ( .A(n13668), .B(n13669), .Z(n13667) );
  OR U18011 ( .A(n13670), .B(n13671), .Z(n13666) );
  ANDN U18012 ( .B(n13672), .A(n13673), .Z(n13624) );
  IV U18013 ( .A(n13674), .Z(n13672) );
  ANDN U18014 ( .B(n13675), .A(n13676), .Z(n13616) );
  XOR U18015 ( .A(n13602), .B(n13677), .Z(n13614) );
  XOR U18016 ( .A(n13603), .B(n13604), .Z(n13677) );
  XOR U18017 ( .A(n13609), .B(n13678), .Z(n13604) );
  XOR U18018 ( .A(n13608), .B(n13611), .Z(n13678) );
  IV U18019 ( .A(n13610), .Z(n13611) );
  NAND U18020 ( .A(n13679), .B(n13680), .Z(n13610) );
  OR U18021 ( .A(n13681), .B(n13682), .Z(n13680) );
  OR U18022 ( .A(n13683), .B(n13684), .Z(n13679) );
  NAND U18023 ( .A(n13685), .B(n13686), .Z(n13608) );
  OR U18024 ( .A(n13687), .B(n13688), .Z(n13686) );
  OR U18025 ( .A(n13689), .B(n13690), .Z(n13685) );
  NOR U18026 ( .A(n13691), .B(n13692), .Z(n13609) );
  ANDN U18027 ( .B(n13693), .A(n13694), .Z(n13603) );
  IV U18028 ( .A(n13695), .Z(n13693) );
  XNOR U18029 ( .A(n13596), .B(n13696), .Z(n13602) );
  XNOR U18030 ( .A(n13595), .B(n13597), .Z(n13696) );
  NAND U18031 ( .A(n13697), .B(n13698), .Z(n13597) );
  OR U18032 ( .A(n13699), .B(n13700), .Z(n13698) );
  OR U18033 ( .A(n13701), .B(n13702), .Z(n13697) );
  NAND U18034 ( .A(n13703), .B(n13704), .Z(n13595) );
  OR U18035 ( .A(n13705), .B(n13706), .Z(n13704) );
  OR U18036 ( .A(n13707), .B(n13708), .Z(n13703) );
  ANDN U18037 ( .B(n13709), .A(n13710), .Z(n13596) );
  IV U18038 ( .A(n13711), .Z(n13709) );
  XNOR U18039 ( .A(n13676), .B(n13675), .Z(N29033) );
  XOR U18040 ( .A(n13695), .B(n13694), .Z(n13675) );
  XNOR U18041 ( .A(n13710), .B(n13711), .Z(n13694) );
  XNOR U18042 ( .A(n13705), .B(n13706), .Z(n13711) );
  XNOR U18043 ( .A(n13707), .B(n13708), .Z(n13706) );
  XNOR U18044 ( .A(y[2212]), .B(x[2212]), .Z(n13708) );
  XNOR U18045 ( .A(y[2213]), .B(x[2213]), .Z(n13707) );
  XNOR U18046 ( .A(y[2211]), .B(x[2211]), .Z(n13705) );
  XNOR U18047 ( .A(n13699), .B(n13700), .Z(n13710) );
  XNOR U18048 ( .A(y[2208]), .B(x[2208]), .Z(n13700) );
  XNOR U18049 ( .A(n13701), .B(n13702), .Z(n13699) );
  XNOR U18050 ( .A(y[2209]), .B(x[2209]), .Z(n13702) );
  XNOR U18051 ( .A(y[2210]), .B(x[2210]), .Z(n13701) );
  XNOR U18052 ( .A(n13692), .B(n13691), .Z(n13695) );
  XNOR U18053 ( .A(n13687), .B(n13688), .Z(n13691) );
  XNOR U18054 ( .A(y[2205]), .B(x[2205]), .Z(n13688) );
  XNOR U18055 ( .A(n13689), .B(n13690), .Z(n13687) );
  XNOR U18056 ( .A(y[2206]), .B(x[2206]), .Z(n13690) );
  XNOR U18057 ( .A(y[2207]), .B(x[2207]), .Z(n13689) );
  XNOR U18058 ( .A(n13681), .B(n13682), .Z(n13692) );
  XNOR U18059 ( .A(y[2202]), .B(x[2202]), .Z(n13682) );
  XNOR U18060 ( .A(n13683), .B(n13684), .Z(n13681) );
  XNOR U18061 ( .A(y[2203]), .B(x[2203]), .Z(n13684) );
  XNOR U18062 ( .A(y[2204]), .B(x[2204]), .Z(n13683) );
  XOR U18063 ( .A(n13657), .B(n13658), .Z(n13676) );
  XNOR U18064 ( .A(n13673), .B(n13674), .Z(n13658) );
  XNOR U18065 ( .A(n13668), .B(n13669), .Z(n13674) );
  XNOR U18066 ( .A(n13670), .B(n13671), .Z(n13669) );
  XNOR U18067 ( .A(y[2200]), .B(x[2200]), .Z(n13671) );
  XNOR U18068 ( .A(y[2201]), .B(x[2201]), .Z(n13670) );
  XNOR U18069 ( .A(y[2199]), .B(x[2199]), .Z(n13668) );
  XNOR U18070 ( .A(n13662), .B(n13663), .Z(n13673) );
  XNOR U18071 ( .A(y[2196]), .B(x[2196]), .Z(n13663) );
  XNOR U18072 ( .A(n13664), .B(n13665), .Z(n13662) );
  XNOR U18073 ( .A(y[2197]), .B(x[2197]), .Z(n13665) );
  XNOR U18074 ( .A(y[2198]), .B(x[2198]), .Z(n13664) );
  XOR U18075 ( .A(n13656), .B(n13655), .Z(n13657) );
  XNOR U18076 ( .A(n13651), .B(n13652), .Z(n13655) );
  XNOR U18077 ( .A(y[2193]), .B(x[2193]), .Z(n13652) );
  XNOR U18078 ( .A(n13653), .B(n13654), .Z(n13651) );
  XNOR U18079 ( .A(y[2194]), .B(x[2194]), .Z(n13654) );
  XNOR U18080 ( .A(y[2195]), .B(x[2195]), .Z(n13653) );
  XNOR U18081 ( .A(n13645), .B(n13646), .Z(n13656) );
  XNOR U18082 ( .A(y[2190]), .B(x[2190]), .Z(n13646) );
  XNOR U18083 ( .A(n13647), .B(n13648), .Z(n13645) );
  XNOR U18084 ( .A(y[2191]), .B(x[2191]), .Z(n13648) );
  XNOR U18085 ( .A(y[2192]), .B(x[2192]), .Z(n13647) );
  NAND U18086 ( .A(n13712), .B(n13713), .Z(N29025) );
  NANDN U18087 ( .A(n13714), .B(n13715), .Z(n13713) );
  OR U18088 ( .A(n13716), .B(n13717), .Z(n13715) );
  NAND U18089 ( .A(n13716), .B(n13717), .Z(n13712) );
  XOR U18090 ( .A(n13716), .B(n13718), .Z(N29024) );
  XNOR U18091 ( .A(n13714), .B(n13717), .Z(n13718) );
  AND U18092 ( .A(n13719), .B(n13720), .Z(n13717) );
  NANDN U18093 ( .A(n13721), .B(n13722), .Z(n13720) );
  NANDN U18094 ( .A(n13723), .B(n13724), .Z(n13722) );
  NANDN U18095 ( .A(n13724), .B(n13723), .Z(n13719) );
  NAND U18096 ( .A(n13725), .B(n13726), .Z(n13714) );
  NANDN U18097 ( .A(n13727), .B(n13728), .Z(n13726) );
  OR U18098 ( .A(n13729), .B(n13730), .Z(n13728) );
  NAND U18099 ( .A(n13730), .B(n13729), .Z(n13725) );
  AND U18100 ( .A(n13731), .B(n13732), .Z(n13716) );
  NANDN U18101 ( .A(n13733), .B(n13734), .Z(n13732) );
  NANDN U18102 ( .A(n13735), .B(n13736), .Z(n13734) );
  NANDN U18103 ( .A(n13736), .B(n13735), .Z(n13731) );
  XOR U18104 ( .A(n13730), .B(n13737), .Z(N29023) );
  XOR U18105 ( .A(n13727), .B(n13729), .Z(n13737) );
  XNOR U18106 ( .A(n13723), .B(n13738), .Z(n13729) );
  XNOR U18107 ( .A(n13721), .B(n13724), .Z(n13738) );
  NAND U18108 ( .A(n13739), .B(n13740), .Z(n13724) );
  NAND U18109 ( .A(n13741), .B(n13742), .Z(n13740) );
  OR U18110 ( .A(n13743), .B(n13744), .Z(n13741) );
  NANDN U18111 ( .A(n13745), .B(n13743), .Z(n13739) );
  IV U18112 ( .A(n13744), .Z(n13745) );
  NAND U18113 ( .A(n13746), .B(n13747), .Z(n13721) );
  NAND U18114 ( .A(n13748), .B(n13749), .Z(n13747) );
  NANDN U18115 ( .A(n13750), .B(n13751), .Z(n13748) );
  NANDN U18116 ( .A(n13751), .B(n13750), .Z(n13746) );
  AND U18117 ( .A(n13752), .B(n13753), .Z(n13723) );
  NAND U18118 ( .A(n13754), .B(n13755), .Z(n13753) );
  OR U18119 ( .A(n13756), .B(n13757), .Z(n13754) );
  NANDN U18120 ( .A(n13758), .B(n13756), .Z(n13752) );
  NAND U18121 ( .A(n13759), .B(n13760), .Z(n13727) );
  NANDN U18122 ( .A(n13761), .B(n13762), .Z(n13760) );
  OR U18123 ( .A(n13763), .B(n13764), .Z(n13762) );
  NANDN U18124 ( .A(n13765), .B(n13763), .Z(n13759) );
  IV U18125 ( .A(n13764), .Z(n13765) );
  XNOR U18126 ( .A(n13735), .B(n13766), .Z(n13730) );
  XNOR U18127 ( .A(n13733), .B(n13736), .Z(n13766) );
  NAND U18128 ( .A(n13767), .B(n13768), .Z(n13736) );
  NAND U18129 ( .A(n13769), .B(n13770), .Z(n13768) );
  OR U18130 ( .A(n13771), .B(n13772), .Z(n13769) );
  NANDN U18131 ( .A(n13773), .B(n13771), .Z(n13767) );
  IV U18132 ( .A(n13772), .Z(n13773) );
  NAND U18133 ( .A(n13774), .B(n13775), .Z(n13733) );
  NAND U18134 ( .A(n13776), .B(n13777), .Z(n13775) );
  NANDN U18135 ( .A(n13778), .B(n13779), .Z(n13776) );
  NANDN U18136 ( .A(n13779), .B(n13778), .Z(n13774) );
  AND U18137 ( .A(n13780), .B(n13781), .Z(n13735) );
  NAND U18138 ( .A(n13782), .B(n13783), .Z(n13781) );
  OR U18139 ( .A(n13784), .B(n13785), .Z(n13782) );
  NANDN U18140 ( .A(n13786), .B(n13784), .Z(n13780) );
  XNOR U18141 ( .A(n13761), .B(n13787), .Z(N29022) );
  XOR U18142 ( .A(n13763), .B(n13764), .Z(n13787) );
  XNOR U18143 ( .A(n13777), .B(n13788), .Z(n13764) );
  XOR U18144 ( .A(n13778), .B(n13779), .Z(n13788) );
  XOR U18145 ( .A(n13784), .B(n13789), .Z(n13779) );
  XOR U18146 ( .A(n13783), .B(n13786), .Z(n13789) );
  IV U18147 ( .A(n13785), .Z(n13786) );
  NAND U18148 ( .A(n13790), .B(n13791), .Z(n13785) );
  OR U18149 ( .A(n13792), .B(n13793), .Z(n13791) );
  OR U18150 ( .A(n13794), .B(n13795), .Z(n13790) );
  NAND U18151 ( .A(n13796), .B(n13797), .Z(n13783) );
  OR U18152 ( .A(n13798), .B(n13799), .Z(n13797) );
  OR U18153 ( .A(n13800), .B(n13801), .Z(n13796) );
  NOR U18154 ( .A(n13802), .B(n13803), .Z(n13784) );
  ANDN U18155 ( .B(n13804), .A(n13805), .Z(n13778) );
  XNOR U18156 ( .A(n13771), .B(n13806), .Z(n13777) );
  XNOR U18157 ( .A(n13770), .B(n13772), .Z(n13806) );
  NAND U18158 ( .A(n13807), .B(n13808), .Z(n13772) );
  OR U18159 ( .A(n13809), .B(n13810), .Z(n13808) );
  OR U18160 ( .A(n13811), .B(n13812), .Z(n13807) );
  NAND U18161 ( .A(n13813), .B(n13814), .Z(n13770) );
  OR U18162 ( .A(n13815), .B(n13816), .Z(n13814) );
  OR U18163 ( .A(n13817), .B(n13818), .Z(n13813) );
  ANDN U18164 ( .B(n13819), .A(n13820), .Z(n13771) );
  IV U18165 ( .A(n13821), .Z(n13819) );
  ANDN U18166 ( .B(n13822), .A(n13823), .Z(n13763) );
  XOR U18167 ( .A(n13749), .B(n13824), .Z(n13761) );
  XOR U18168 ( .A(n13750), .B(n13751), .Z(n13824) );
  XOR U18169 ( .A(n13756), .B(n13825), .Z(n13751) );
  XOR U18170 ( .A(n13755), .B(n13758), .Z(n13825) );
  IV U18171 ( .A(n13757), .Z(n13758) );
  NAND U18172 ( .A(n13826), .B(n13827), .Z(n13757) );
  OR U18173 ( .A(n13828), .B(n13829), .Z(n13827) );
  OR U18174 ( .A(n13830), .B(n13831), .Z(n13826) );
  NAND U18175 ( .A(n13832), .B(n13833), .Z(n13755) );
  OR U18176 ( .A(n13834), .B(n13835), .Z(n13833) );
  OR U18177 ( .A(n13836), .B(n13837), .Z(n13832) );
  NOR U18178 ( .A(n13838), .B(n13839), .Z(n13756) );
  ANDN U18179 ( .B(n13840), .A(n13841), .Z(n13750) );
  IV U18180 ( .A(n13842), .Z(n13840) );
  XNOR U18181 ( .A(n13743), .B(n13843), .Z(n13749) );
  XNOR U18182 ( .A(n13742), .B(n13744), .Z(n13843) );
  NAND U18183 ( .A(n13844), .B(n13845), .Z(n13744) );
  OR U18184 ( .A(n13846), .B(n13847), .Z(n13845) );
  OR U18185 ( .A(n13848), .B(n13849), .Z(n13844) );
  NAND U18186 ( .A(n13850), .B(n13851), .Z(n13742) );
  OR U18187 ( .A(n13852), .B(n13853), .Z(n13851) );
  OR U18188 ( .A(n13854), .B(n13855), .Z(n13850) );
  ANDN U18189 ( .B(n13856), .A(n13857), .Z(n13743) );
  IV U18190 ( .A(n13858), .Z(n13856) );
  XNOR U18191 ( .A(n13823), .B(n13822), .Z(N29021) );
  XOR U18192 ( .A(n13842), .B(n13841), .Z(n13822) );
  XNOR U18193 ( .A(n13857), .B(n13858), .Z(n13841) );
  XNOR U18194 ( .A(n13852), .B(n13853), .Z(n13858) );
  XNOR U18195 ( .A(n13854), .B(n13855), .Z(n13853) );
  XNOR U18196 ( .A(y[2188]), .B(x[2188]), .Z(n13855) );
  XNOR U18197 ( .A(y[2189]), .B(x[2189]), .Z(n13854) );
  XNOR U18198 ( .A(y[2187]), .B(x[2187]), .Z(n13852) );
  XNOR U18199 ( .A(n13846), .B(n13847), .Z(n13857) );
  XNOR U18200 ( .A(y[2184]), .B(x[2184]), .Z(n13847) );
  XNOR U18201 ( .A(n13848), .B(n13849), .Z(n13846) );
  XNOR U18202 ( .A(y[2185]), .B(x[2185]), .Z(n13849) );
  XNOR U18203 ( .A(y[2186]), .B(x[2186]), .Z(n13848) );
  XNOR U18204 ( .A(n13839), .B(n13838), .Z(n13842) );
  XNOR U18205 ( .A(n13834), .B(n13835), .Z(n13838) );
  XNOR U18206 ( .A(y[2181]), .B(x[2181]), .Z(n13835) );
  XNOR U18207 ( .A(n13836), .B(n13837), .Z(n13834) );
  XNOR U18208 ( .A(y[2182]), .B(x[2182]), .Z(n13837) );
  XNOR U18209 ( .A(y[2183]), .B(x[2183]), .Z(n13836) );
  XNOR U18210 ( .A(n13828), .B(n13829), .Z(n13839) );
  XNOR U18211 ( .A(y[2178]), .B(x[2178]), .Z(n13829) );
  XNOR U18212 ( .A(n13830), .B(n13831), .Z(n13828) );
  XNOR U18213 ( .A(y[2179]), .B(x[2179]), .Z(n13831) );
  XNOR U18214 ( .A(y[2180]), .B(x[2180]), .Z(n13830) );
  XOR U18215 ( .A(n13804), .B(n13805), .Z(n13823) );
  XNOR U18216 ( .A(n13820), .B(n13821), .Z(n13805) );
  XNOR U18217 ( .A(n13815), .B(n13816), .Z(n13821) );
  XNOR U18218 ( .A(n13817), .B(n13818), .Z(n13816) );
  XNOR U18219 ( .A(y[2176]), .B(x[2176]), .Z(n13818) );
  XNOR U18220 ( .A(y[2177]), .B(x[2177]), .Z(n13817) );
  XNOR U18221 ( .A(y[2175]), .B(x[2175]), .Z(n13815) );
  XNOR U18222 ( .A(n13809), .B(n13810), .Z(n13820) );
  XNOR U18223 ( .A(y[2172]), .B(x[2172]), .Z(n13810) );
  XNOR U18224 ( .A(n13811), .B(n13812), .Z(n13809) );
  XNOR U18225 ( .A(y[2173]), .B(x[2173]), .Z(n13812) );
  XNOR U18226 ( .A(y[2174]), .B(x[2174]), .Z(n13811) );
  XOR U18227 ( .A(n13803), .B(n13802), .Z(n13804) );
  XNOR U18228 ( .A(n13798), .B(n13799), .Z(n13802) );
  XNOR U18229 ( .A(y[2169]), .B(x[2169]), .Z(n13799) );
  XNOR U18230 ( .A(n13800), .B(n13801), .Z(n13798) );
  XNOR U18231 ( .A(y[2170]), .B(x[2170]), .Z(n13801) );
  XNOR U18232 ( .A(y[2171]), .B(x[2171]), .Z(n13800) );
  XNOR U18233 ( .A(n13792), .B(n13793), .Z(n13803) );
  XNOR U18234 ( .A(y[2166]), .B(x[2166]), .Z(n13793) );
  XNOR U18235 ( .A(n13794), .B(n13795), .Z(n13792) );
  XNOR U18236 ( .A(y[2167]), .B(x[2167]), .Z(n13795) );
  XNOR U18237 ( .A(y[2168]), .B(x[2168]), .Z(n13794) );
  NAND U18238 ( .A(n13859), .B(n13860), .Z(N29013) );
  NANDN U18239 ( .A(n13861), .B(n13862), .Z(n13860) );
  OR U18240 ( .A(n13863), .B(n13864), .Z(n13862) );
  NAND U18241 ( .A(n13863), .B(n13864), .Z(n13859) );
  XOR U18242 ( .A(n13863), .B(n13865), .Z(N29012) );
  XNOR U18243 ( .A(n13861), .B(n13864), .Z(n13865) );
  AND U18244 ( .A(n13866), .B(n13867), .Z(n13864) );
  NANDN U18245 ( .A(n13868), .B(n13869), .Z(n13867) );
  NANDN U18246 ( .A(n13870), .B(n13871), .Z(n13869) );
  NANDN U18247 ( .A(n13871), .B(n13870), .Z(n13866) );
  NAND U18248 ( .A(n13872), .B(n13873), .Z(n13861) );
  NANDN U18249 ( .A(n13874), .B(n13875), .Z(n13873) );
  OR U18250 ( .A(n13876), .B(n13877), .Z(n13875) );
  NAND U18251 ( .A(n13877), .B(n13876), .Z(n13872) );
  AND U18252 ( .A(n13878), .B(n13879), .Z(n13863) );
  NANDN U18253 ( .A(n13880), .B(n13881), .Z(n13879) );
  NANDN U18254 ( .A(n13882), .B(n13883), .Z(n13881) );
  NANDN U18255 ( .A(n13883), .B(n13882), .Z(n13878) );
  XOR U18256 ( .A(n13877), .B(n13884), .Z(N29011) );
  XOR U18257 ( .A(n13874), .B(n13876), .Z(n13884) );
  XNOR U18258 ( .A(n13870), .B(n13885), .Z(n13876) );
  XNOR U18259 ( .A(n13868), .B(n13871), .Z(n13885) );
  NAND U18260 ( .A(n13886), .B(n13887), .Z(n13871) );
  NAND U18261 ( .A(n13888), .B(n13889), .Z(n13887) );
  OR U18262 ( .A(n13890), .B(n13891), .Z(n13888) );
  NANDN U18263 ( .A(n13892), .B(n13890), .Z(n13886) );
  IV U18264 ( .A(n13891), .Z(n13892) );
  NAND U18265 ( .A(n13893), .B(n13894), .Z(n13868) );
  NAND U18266 ( .A(n13895), .B(n13896), .Z(n13894) );
  NANDN U18267 ( .A(n13897), .B(n13898), .Z(n13895) );
  NANDN U18268 ( .A(n13898), .B(n13897), .Z(n13893) );
  AND U18269 ( .A(n13899), .B(n13900), .Z(n13870) );
  NAND U18270 ( .A(n13901), .B(n13902), .Z(n13900) );
  OR U18271 ( .A(n13903), .B(n13904), .Z(n13901) );
  NANDN U18272 ( .A(n13905), .B(n13903), .Z(n13899) );
  NAND U18273 ( .A(n13906), .B(n13907), .Z(n13874) );
  NANDN U18274 ( .A(n13908), .B(n13909), .Z(n13907) );
  OR U18275 ( .A(n13910), .B(n13911), .Z(n13909) );
  NANDN U18276 ( .A(n13912), .B(n13910), .Z(n13906) );
  IV U18277 ( .A(n13911), .Z(n13912) );
  XNOR U18278 ( .A(n13882), .B(n13913), .Z(n13877) );
  XNOR U18279 ( .A(n13880), .B(n13883), .Z(n13913) );
  NAND U18280 ( .A(n13914), .B(n13915), .Z(n13883) );
  NAND U18281 ( .A(n13916), .B(n13917), .Z(n13915) );
  OR U18282 ( .A(n13918), .B(n13919), .Z(n13916) );
  NANDN U18283 ( .A(n13920), .B(n13918), .Z(n13914) );
  IV U18284 ( .A(n13919), .Z(n13920) );
  NAND U18285 ( .A(n13921), .B(n13922), .Z(n13880) );
  NAND U18286 ( .A(n13923), .B(n13924), .Z(n13922) );
  NANDN U18287 ( .A(n13925), .B(n13926), .Z(n13923) );
  NANDN U18288 ( .A(n13926), .B(n13925), .Z(n13921) );
  AND U18289 ( .A(n13927), .B(n13928), .Z(n13882) );
  NAND U18290 ( .A(n13929), .B(n13930), .Z(n13928) );
  OR U18291 ( .A(n13931), .B(n13932), .Z(n13929) );
  NANDN U18292 ( .A(n13933), .B(n13931), .Z(n13927) );
  XNOR U18293 ( .A(n13908), .B(n13934), .Z(N29010) );
  XOR U18294 ( .A(n13910), .B(n13911), .Z(n13934) );
  XNOR U18295 ( .A(n13924), .B(n13935), .Z(n13911) );
  XOR U18296 ( .A(n13925), .B(n13926), .Z(n13935) );
  XOR U18297 ( .A(n13931), .B(n13936), .Z(n13926) );
  XOR U18298 ( .A(n13930), .B(n13933), .Z(n13936) );
  IV U18299 ( .A(n13932), .Z(n13933) );
  NAND U18300 ( .A(n13937), .B(n13938), .Z(n13932) );
  OR U18301 ( .A(n13939), .B(n13940), .Z(n13938) );
  OR U18302 ( .A(n13941), .B(n13942), .Z(n13937) );
  NAND U18303 ( .A(n13943), .B(n13944), .Z(n13930) );
  OR U18304 ( .A(n13945), .B(n13946), .Z(n13944) );
  OR U18305 ( .A(n13947), .B(n13948), .Z(n13943) );
  NOR U18306 ( .A(n13949), .B(n13950), .Z(n13931) );
  ANDN U18307 ( .B(n13951), .A(n13952), .Z(n13925) );
  XNOR U18308 ( .A(n13918), .B(n13953), .Z(n13924) );
  XNOR U18309 ( .A(n13917), .B(n13919), .Z(n13953) );
  NAND U18310 ( .A(n13954), .B(n13955), .Z(n13919) );
  OR U18311 ( .A(n13956), .B(n13957), .Z(n13955) );
  OR U18312 ( .A(n13958), .B(n13959), .Z(n13954) );
  NAND U18313 ( .A(n13960), .B(n13961), .Z(n13917) );
  OR U18314 ( .A(n13962), .B(n13963), .Z(n13961) );
  OR U18315 ( .A(n13964), .B(n13965), .Z(n13960) );
  ANDN U18316 ( .B(n13966), .A(n13967), .Z(n13918) );
  IV U18317 ( .A(n13968), .Z(n13966) );
  ANDN U18318 ( .B(n13969), .A(n13970), .Z(n13910) );
  XOR U18319 ( .A(n13896), .B(n13971), .Z(n13908) );
  XOR U18320 ( .A(n13897), .B(n13898), .Z(n13971) );
  XOR U18321 ( .A(n13903), .B(n13972), .Z(n13898) );
  XOR U18322 ( .A(n13902), .B(n13905), .Z(n13972) );
  IV U18323 ( .A(n13904), .Z(n13905) );
  NAND U18324 ( .A(n13973), .B(n13974), .Z(n13904) );
  OR U18325 ( .A(n13975), .B(n13976), .Z(n13974) );
  OR U18326 ( .A(n13977), .B(n13978), .Z(n13973) );
  NAND U18327 ( .A(n13979), .B(n13980), .Z(n13902) );
  OR U18328 ( .A(n13981), .B(n13982), .Z(n13980) );
  OR U18329 ( .A(n13983), .B(n13984), .Z(n13979) );
  NOR U18330 ( .A(n13985), .B(n13986), .Z(n13903) );
  ANDN U18331 ( .B(n13987), .A(n13988), .Z(n13897) );
  IV U18332 ( .A(n13989), .Z(n13987) );
  XNOR U18333 ( .A(n13890), .B(n13990), .Z(n13896) );
  XNOR U18334 ( .A(n13889), .B(n13891), .Z(n13990) );
  NAND U18335 ( .A(n13991), .B(n13992), .Z(n13891) );
  OR U18336 ( .A(n13993), .B(n13994), .Z(n13992) );
  OR U18337 ( .A(n13995), .B(n13996), .Z(n13991) );
  NAND U18338 ( .A(n13997), .B(n13998), .Z(n13889) );
  OR U18339 ( .A(n13999), .B(n14000), .Z(n13998) );
  OR U18340 ( .A(n14001), .B(n14002), .Z(n13997) );
  ANDN U18341 ( .B(n14003), .A(n14004), .Z(n13890) );
  IV U18342 ( .A(n14005), .Z(n14003) );
  XNOR U18343 ( .A(n13970), .B(n13969), .Z(N29009) );
  XOR U18344 ( .A(n13989), .B(n13988), .Z(n13969) );
  XNOR U18345 ( .A(n14004), .B(n14005), .Z(n13988) );
  XNOR U18346 ( .A(n13999), .B(n14000), .Z(n14005) );
  XNOR U18347 ( .A(n14001), .B(n14002), .Z(n14000) );
  XNOR U18348 ( .A(y[2164]), .B(x[2164]), .Z(n14002) );
  XNOR U18349 ( .A(y[2165]), .B(x[2165]), .Z(n14001) );
  XNOR U18350 ( .A(y[2163]), .B(x[2163]), .Z(n13999) );
  XNOR U18351 ( .A(n13993), .B(n13994), .Z(n14004) );
  XNOR U18352 ( .A(y[2160]), .B(x[2160]), .Z(n13994) );
  XNOR U18353 ( .A(n13995), .B(n13996), .Z(n13993) );
  XNOR U18354 ( .A(y[2161]), .B(x[2161]), .Z(n13996) );
  XNOR U18355 ( .A(y[2162]), .B(x[2162]), .Z(n13995) );
  XNOR U18356 ( .A(n13986), .B(n13985), .Z(n13989) );
  XNOR U18357 ( .A(n13981), .B(n13982), .Z(n13985) );
  XNOR U18358 ( .A(y[2157]), .B(x[2157]), .Z(n13982) );
  XNOR U18359 ( .A(n13983), .B(n13984), .Z(n13981) );
  XNOR U18360 ( .A(y[2158]), .B(x[2158]), .Z(n13984) );
  XNOR U18361 ( .A(y[2159]), .B(x[2159]), .Z(n13983) );
  XNOR U18362 ( .A(n13975), .B(n13976), .Z(n13986) );
  XNOR U18363 ( .A(y[2154]), .B(x[2154]), .Z(n13976) );
  XNOR U18364 ( .A(n13977), .B(n13978), .Z(n13975) );
  XNOR U18365 ( .A(y[2155]), .B(x[2155]), .Z(n13978) );
  XNOR U18366 ( .A(y[2156]), .B(x[2156]), .Z(n13977) );
  XOR U18367 ( .A(n13951), .B(n13952), .Z(n13970) );
  XNOR U18368 ( .A(n13967), .B(n13968), .Z(n13952) );
  XNOR U18369 ( .A(n13962), .B(n13963), .Z(n13968) );
  XNOR U18370 ( .A(n13964), .B(n13965), .Z(n13963) );
  XNOR U18371 ( .A(y[2152]), .B(x[2152]), .Z(n13965) );
  XNOR U18372 ( .A(y[2153]), .B(x[2153]), .Z(n13964) );
  XNOR U18373 ( .A(y[2151]), .B(x[2151]), .Z(n13962) );
  XNOR U18374 ( .A(n13956), .B(n13957), .Z(n13967) );
  XNOR U18375 ( .A(y[2148]), .B(x[2148]), .Z(n13957) );
  XNOR U18376 ( .A(n13958), .B(n13959), .Z(n13956) );
  XNOR U18377 ( .A(y[2149]), .B(x[2149]), .Z(n13959) );
  XNOR U18378 ( .A(y[2150]), .B(x[2150]), .Z(n13958) );
  XOR U18379 ( .A(n13950), .B(n13949), .Z(n13951) );
  XNOR U18380 ( .A(n13945), .B(n13946), .Z(n13949) );
  XNOR U18381 ( .A(y[2145]), .B(x[2145]), .Z(n13946) );
  XNOR U18382 ( .A(n13947), .B(n13948), .Z(n13945) );
  XNOR U18383 ( .A(y[2146]), .B(x[2146]), .Z(n13948) );
  XNOR U18384 ( .A(y[2147]), .B(x[2147]), .Z(n13947) );
  XNOR U18385 ( .A(n13939), .B(n13940), .Z(n13950) );
  XNOR U18386 ( .A(y[2142]), .B(x[2142]), .Z(n13940) );
  XNOR U18387 ( .A(n13941), .B(n13942), .Z(n13939) );
  XNOR U18388 ( .A(y[2143]), .B(x[2143]), .Z(n13942) );
  XNOR U18389 ( .A(y[2144]), .B(x[2144]), .Z(n13941) );
  NAND U18390 ( .A(n14006), .B(n14007), .Z(N29001) );
  NANDN U18391 ( .A(n14008), .B(n14009), .Z(n14007) );
  OR U18392 ( .A(n14010), .B(n14011), .Z(n14009) );
  NAND U18393 ( .A(n14010), .B(n14011), .Z(n14006) );
  XOR U18394 ( .A(n14010), .B(n14012), .Z(N29000) );
  XNOR U18395 ( .A(n14008), .B(n14011), .Z(n14012) );
  AND U18396 ( .A(n14013), .B(n14014), .Z(n14011) );
  NANDN U18397 ( .A(n14015), .B(n14016), .Z(n14014) );
  NANDN U18398 ( .A(n14017), .B(n14018), .Z(n14016) );
  NANDN U18399 ( .A(n14018), .B(n14017), .Z(n14013) );
  NAND U18400 ( .A(n14019), .B(n14020), .Z(n14008) );
  NANDN U18401 ( .A(n14021), .B(n14022), .Z(n14020) );
  OR U18402 ( .A(n14023), .B(n14024), .Z(n14022) );
  NAND U18403 ( .A(n14024), .B(n14023), .Z(n14019) );
  AND U18404 ( .A(n14025), .B(n14026), .Z(n14010) );
  NANDN U18405 ( .A(n14027), .B(n14028), .Z(n14026) );
  NANDN U18406 ( .A(n14029), .B(n14030), .Z(n14028) );
  NANDN U18407 ( .A(n14030), .B(n14029), .Z(n14025) );
  XOR U18408 ( .A(n14024), .B(n14031), .Z(N28999) );
  XOR U18409 ( .A(n14021), .B(n14023), .Z(n14031) );
  XNOR U18410 ( .A(n14017), .B(n14032), .Z(n14023) );
  XNOR U18411 ( .A(n14015), .B(n14018), .Z(n14032) );
  NAND U18412 ( .A(n14033), .B(n14034), .Z(n14018) );
  NAND U18413 ( .A(n14035), .B(n14036), .Z(n14034) );
  OR U18414 ( .A(n14037), .B(n14038), .Z(n14035) );
  NANDN U18415 ( .A(n14039), .B(n14037), .Z(n14033) );
  IV U18416 ( .A(n14038), .Z(n14039) );
  NAND U18417 ( .A(n14040), .B(n14041), .Z(n14015) );
  NAND U18418 ( .A(n14042), .B(n14043), .Z(n14041) );
  NANDN U18419 ( .A(n14044), .B(n14045), .Z(n14042) );
  NANDN U18420 ( .A(n14045), .B(n14044), .Z(n14040) );
  AND U18421 ( .A(n14046), .B(n14047), .Z(n14017) );
  NAND U18422 ( .A(n14048), .B(n14049), .Z(n14047) );
  OR U18423 ( .A(n14050), .B(n14051), .Z(n14048) );
  NANDN U18424 ( .A(n14052), .B(n14050), .Z(n14046) );
  NAND U18425 ( .A(n14053), .B(n14054), .Z(n14021) );
  NANDN U18426 ( .A(n14055), .B(n14056), .Z(n14054) );
  OR U18427 ( .A(n14057), .B(n14058), .Z(n14056) );
  NANDN U18428 ( .A(n14059), .B(n14057), .Z(n14053) );
  IV U18429 ( .A(n14058), .Z(n14059) );
  XNOR U18430 ( .A(n14029), .B(n14060), .Z(n14024) );
  XNOR U18431 ( .A(n14027), .B(n14030), .Z(n14060) );
  NAND U18432 ( .A(n14061), .B(n14062), .Z(n14030) );
  NAND U18433 ( .A(n14063), .B(n14064), .Z(n14062) );
  OR U18434 ( .A(n14065), .B(n14066), .Z(n14063) );
  NANDN U18435 ( .A(n14067), .B(n14065), .Z(n14061) );
  IV U18436 ( .A(n14066), .Z(n14067) );
  NAND U18437 ( .A(n14068), .B(n14069), .Z(n14027) );
  NAND U18438 ( .A(n14070), .B(n14071), .Z(n14069) );
  NANDN U18439 ( .A(n14072), .B(n14073), .Z(n14070) );
  NANDN U18440 ( .A(n14073), .B(n14072), .Z(n14068) );
  AND U18441 ( .A(n14074), .B(n14075), .Z(n14029) );
  NAND U18442 ( .A(n14076), .B(n14077), .Z(n14075) );
  OR U18443 ( .A(n14078), .B(n14079), .Z(n14076) );
  NANDN U18444 ( .A(n14080), .B(n14078), .Z(n14074) );
  XNOR U18445 ( .A(n14055), .B(n14081), .Z(N28998) );
  XOR U18446 ( .A(n14057), .B(n14058), .Z(n14081) );
  XNOR U18447 ( .A(n14071), .B(n14082), .Z(n14058) );
  XOR U18448 ( .A(n14072), .B(n14073), .Z(n14082) );
  XOR U18449 ( .A(n14078), .B(n14083), .Z(n14073) );
  XOR U18450 ( .A(n14077), .B(n14080), .Z(n14083) );
  IV U18451 ( .A(n14079), .Z(n14080) );
  NAND U18452 ( .A(n14084), .B(n14085), .Z(n14079) );
  OR U18453 ( .A(n14086), .B(n14087), .Z(n14085) );
  OR U18454 ( .A(n14088), .B(n14089), .Z(n14084) );
  NAND U18455 ( .A(n14090), .B(n14091), .Z(n14077) );
  OR U18456 ( .A(n14092), .B(n14093), .Z(n14091) );
  OR U18457 ( .A(n14094), .B(n14095), .Z(n14090) );
  NOR U18458 ( .A(n14096), .B(n14097), .Z(n14078) );
  ANDN U18459 ( .B(n14098), .A(n14099), .Z(n14072) );
  XNOR U18460 ( .A(n14065), .B(n14100), .Z(n14071) );
  XNOR U18461 ( .A(n14064), .B(n14066), .Z(n14100) );
  NAND U18462 ( .A(n14101), .B(n14102), .Z(n14066) );
  OR U18463 ( .A(n14103), .B(n14104), .Z(n14102) );
  OR U18464 ( .A(n14105), .B(n14106), .Z(n14101) );
  NAND U18465 ( .A(n14107), .B(n14108), .Z(n14064) );
  OR U18466 ( .A(n14109), .B(n14110), .Z(n14108) );
  OR U18467 ( .A(n14111), .B(n14112), .Z(n14107) );
  ANDN U18468 ( .B(n14113), .A(n14114), .Z(n14065) );
  IV U18469 ( .A(n14115), .Z(n14113) );
  ANDN U18470 ( .B(n14116), .A(n14117), .Z(n14057) );
  XOR U18471 ( .A(n14043), .B(n14118), .Z(n14055) );
  XOR U18472 ( .A(n14044), .B(n14045), .Z(n14118) );
  XOR U18473 ( .A(n14050), .B(n14119), .Z(n14045) );
  XOR U18474 ( .A(n14049), .B(n14052), .Z(n14119) );
  IV U18475 ( .A(n14051), .Z(n14052) );
  NAND U18476 ( .A(n14120), .B(n14121), .Z(n14051) );
  OR U18477 ( .A(n14122), .B(n14123), .Z(n14121) );
  OR U18478 ( .A(n14124), .B(n14125), .Z(n14120) );
  NAND U18479 ( .A(n14126), .B(n14127), .Z(n14049) );
  OR U18480 ( .A(n14128), .B(n14129), .Z(n14127) );
  OR U18481 ( .A(n14130), .B(n14131), .Z(n14126) );
  NOR U18482 ( .A(n14132), .B(n14133), .Z(n14050) );
  ANDN U18483 ( .B(n14134), .A(n14135), .Z(n14044) );
  IV U18484 ( .A(n14136), .Z(n14134) );
  XNOR U18485 ( .A(n14037), .B(n14137), .Z(n14043) );
  XNOR U18486 ( .A(n14036), .B(n14038), .Z(n14137) );
  NAND U18487 ( .A(n14138), .B(n14139), .Z(n14038) );
  OR U18488 ( .A(n14140), .B(n14141), .Z(n14139) );
  OR U18489 ( .A(n14142), .B(n14143), .Z(n14138) );
  NAND U18490 ( .A(n14144), .B(n14145), .Z(n14036) );
  OR U18491 ( .A(n14146), .B(n14147), .Z(n14145) );
  OR U18492 ( .A(n14148), .B(n14149), .Z(n14144) );
  ANDN U18493 ( .B(n14150), .A(n14151), .Z(n14037) );
  IV U18494 ( .A(n14152), .Z(n14150) );
  XNOR U18495 ( .A(n14117), .B(n14116), .Z(N28997) );
  XOR U18496 ( .A(n14136), .B(n14135), .Z(n14116) );
  XNOR U18497 ( .A(n14151), .B(n14152), .Z(n14135) );
  XNOR U18498 ( .A(n14146), .B(n14147), .Z(n14152) );
  XNOR U18499 ( .A(n14148), .B(n14149), .Z(n14147) );
  XNOR U18500 ( .A(y[2140]), .B(x[2140]), .Z(n14149) );
  XNOR U18501 ( .A(y[2141]), .B(x[2141]), .Z(n14148) );
  XNOR U18502 ( .A(y[2139]), .B(x[2139]), .Z(n14146) );
  XNOR U18503 ( .A(n14140), .B(n14141), .Z(n14151) );
  XNOR U18504 ( .A(y[2136]), .B(x[2136]), .Z(n14141) );
  XNOR U18505 ( .A(n14142), .B(n14143), .Z(n14140) );
  XNOR U18506 ( .A(y[2137]), .B(x[2137]), .Z(n14143) );
  XNOR U18507 ( .A(y[2138]), .B(x[2138]), .Z(n14142) );
  XNOR U18508 ( .A(n14133), .B(n14132), .Z(n14136) );
  XNOR U18509 ( .A(n14128), .B(n14129), .Z(n14132) );
  XNOR U18510 ( .A(y[2133]), .B(x[2133]), .Z(n14129) );
  XNOR U18511 ( .A(n14130), .B(n14131), .Z(n14128) );
  XNOR U18512 ( .A(y[2134]), .B(x[2134]), .Z(n14131) );
  XNOR U18513 ( .A(y[2135]), .B(x[2135]), .Z(n14130) );
  XNOR U18514 ( .A(n14122), .B(n14123), .Z(n14133) );
  XNOR U18515 ( .A(y[2130]), .B(x[2130]), .Z(n14123) );
  XNOR U18516 ( .A(n14124), .B(n14125), .Z(n14122) );
  XNOR U18517 ( .A(y[2131]), .B(x[2131]), .Z(n14125) );
  XNOR U18518 ( .A(y[2132]), .B(x[2132]), .Z(n14124) );
  XOR U18519 ( .A(n14098), .B(n14099), .Z(n14117) );
  XNOR U18520 ( .A(n14114), .B(n14115), .Z(n14099) );
  XNOR U18521 ( .A(n14109), .B(n14110), .Z(n14115) );
  XNOR U18522 ( .A(n14111), .B(n14112), .Z(n14110) );
  XNOR U18523 ( .A(y[2128]), .B(x[2128]), .Z(n14112) );
  XNOR U18524 ( .A(y[2129]), .B(x[2129]), .Z(n14111) );
  XNOR U18525 ( .A(y[2127]), .B(x[2127]), .Z(n14109) );
  XNOR U18526 ( .A(n14103), .B(n14104), .Z(n14114) );
  XNOR U18527 ( .A(y[2124]), .B(x[2124]), .Z(n14104) );
  XNOR U18528 ( .A(n14105), .B(n14106), .Z(n14103) );
  XNOR U18529 ( .A(y[2125]), .B(x[2125]), .Z(n14106) );
  XNOR U18530 ( .A(y[2126]), .B(x[2126]), .Z(n14105) );
  XOR U18531 ( .A(n14097), .B(n14096), .Z(n14098) );
  XNOR U18532 ( .A(n14092), .B(n14093), .Z(n14096) );
  XNOR U18533 ( .A(y[2121]), .B(x[2121]), .Z(n14093) );
  XNOR U18534 ( .A(n14094), .B(n14095), .Z(n14092) );
  XNOR U18535 ( .A(y[2122]), .B(x[2122]), .Z(n14095) );
  XNOR U18536 ( .A(y[2123]), .B(x[2123]), .Z(n14094) );
  XNOR U18537 ( .A(n14086), .B(n14087), .Z(n14097) );
  XNOR U18538 ( .A(y[2118]), .B(x[2118]), .Z(n14087) );
  XNOR U18539 ( .A(n14088), .B(n14089), .Z(n14086) );
  XNOR U18540 ( .A(y[2119]), .B(x[2119]), .Z(n14089) );
  XNOR U18541 ( .A(y[2120]), .B(x[2120]), .Z(n14088) );
  NAND U18542 ( .A(n14153), .B(n14154), .Z(N28989) );
  NANDN U18543 ( .A(n14155), .B(n14156), .Z(n14154) );
  OR U18544 ( .A(n14157), .B(n14158), .Z(n14156) );
  NAND U18545 ( .A(n14157), .B(n14158), .Z(n14153) );
  XOR U18546 ( .A(n14157), .B(n14159), .Z(N28988) );
  XNOR U18547 ( .A(n14155), .B(n14158), .Z(n14159) );
  AND U18548 ( .A(n14160), .B(n14161), .Z(n14158) );
  NANDN U18549 ( .A(n14162), .B(n14163), .Z(n14161) );
  NANDN U18550 ( .A(n14164), .B(n14165), .Z(n14163) );
  NANDN U18551 ( .A(n14165), .B(n14164), .Z(n14160) );
  NAND U18552 ( .A(n14166), .B(n14167), .Z(n14155) );
  NANDN U18553 ( .A(n14168), .B(n14169), .Z(n14167) );
  OR U18554 ( .A(n14170), .B(n14171), .Z(n14169) );
  NAND U18555 ( .A(n14171), .B(n14170), .Z(n14166) );
  AND U18556 ( .A(n14172), .B(n14173), .Z(n14157) );
  NANDN U18557 ( .A(n14174), .B(n14175), .Z(n14173) );
  NANDN U18558 ( .A(n14176), .B(n14177), .Z(n14175) );
  NANDN U18559 ( .A(n14177), .B(n14176), .Z(n14172) );
  XOR U18560 ( .A(n14171), .B(n14178), .Z(N28987) );
  XOR U18561 ( .A(n14168), .B(n14170), .Z(n14178) );
  XNOR U18562 ( .A(n14164), .B(n14179), .Z(n14170) );
  XNOR U18563 ( .A(n14162), .B(n14165), .Z(n14179) );
  NAND U18564 ( .A(n14180), .B(n14181), .Z(n14165) );
  NAND U18565 ( .A(n14182), .B(n14183), .Z(n14181) );
  OR U18566 ( .A(n14184), .B(n14185), .Z(n14182) );
  NANDN U18567 ( .A(n14186), .B(n14184), .Z(n14180) );
  IV U18568 ( .A(n14185), .Z(n14186) );
  NAND U18569 ( .A(n14187), .B(n14188), .Z(n14162) );
  NAND U18570 ( .A(n14189), .B(n14190), .Z(n14188) );
  NANDN U18571 ( .A(n14191), .B(n14192), .Z(n14189) );
  NANDN U18572 ( .A(n14192), .B(n14191), .Z(n14187) );
  AND U18573 ( .A(n14193), .B(n14194), .Z(n14164) );
  NAND U18574 ( .A(n14195), .B(n14196), .Z(n14194) );
  OR U18575 ( .A(n14197), .B(n14198), .Z(n14195) );
  NANDN U18576 ( .A(n14199), .B(n14197), .Z(n14193) );
  NAND U18577 ( .A(n14200), .B(n14201), .Z(n14168) );
  NANDN U18578 ( .A(n14202), .B(n14203), .Z(n14201) );
  OR U18579 ( .A(n14204), .B(n14205), .Z(n14203) );
  NANDN U18580 ( .A(n14206), .B(n14204), .Z(n14200) );
  IV U18581 ( .A(n14205), .Z(n14206) );
  XNOR U18582 ( .A(n14176), .B(n14207), .Z(n14171) );
  XNOR U18583 ( .A(n14174), .B(n14177), .Z(n14207) );
  NAND U18584 ( .A(n14208), .B(n14209), .Z(n14177) );
  NAND U18585 ( .A(n14210), .B(n14211), .Z(n14209) );
  OR U18586 ( .A(n14212), .B(n14213), .Z(n14210) );
  NANDN U18587 ( .A(n14214), .B(n14212), .Z(n14208) );
  IV U18588 ( .A(n14213), .Z(n14214) );
  NAND U18589 ( .A(n14215), .B(n14216), .Z(n14174) );
  NAND U18590 ( .A(n14217), .B(n14218), .Z(n14216) );
  NANDN U18591 ( .A(n14219), .B(n14220), .Z(n14217) );
  NANDN U18592 ( .A(n14220), .B(n14219), .Z(n14215) );
  AND U18593 ( .A(n14221), .B(n14222), .Z(n14176) );
  NAND U18594 ( .A(n14223), .B(n14224), .Z(n14222) );
  OR U18595 ( .A(n14225), .B(n14226), .Z(n14223) );
  NANDN U18596 ( .A(n14227), .B(n14225), .Z(n14221) );
  XNOR U18597 ( .A(n14202), .B(n14228), .Z(N28986) );
  XOR U18598 ( .A(n14204), .B(n14205), .Z(n14228) );
  XNOR U18599 ( .A(n14218), .B(n14229), .Z(n14205) );
  XOR U18600 ( .A(n14219), .B(n14220), .Z(n14229) );
  XOR U18601 ( .A(n14225), .B(n14230), .Z(n14220) );
  XOR U18602 ( .A(n14224), .B(n14227), .Z(n14230) );
  IV U18603 ( .A(n14226), .Z(n14227) );
  NAND U18604 ( .A(n14231), .B(n14232), .Z(n14226) );
  OR U18605 ( .A(n14233), .B(n14234), .Z(n14232) );
  OR U18606 ( .A(n14235), .B(n14236), .Z(n14231) );
  NAND U18607 ( .A(n14237), .B(n14238), .Z(n14224) );
  OR U18608 ( .A(n14239), .B(n14240), .Z(n14238) );
  OR U18609 ( .A(n14241), .B(n14242), .Z(n14237) );
  NOR U18610 ( .A(n14243), .B(n14244), .Z(n14225) );
  ANDN U18611 ( .B(n14245), .A(n14246), .Z(n14219) );
  XNOR U18612 ( .A(n14212), .B(n14247), .Z(n14218) );
  XNOR U18613 ( .A(n14211), .B(n14213), .Z(n14247) );
  NAND U18614 ( .A(n14248), .B(n14249), .Z(n14213) );
  OR U18615 ( .A(n14250), .B(n14251), .Z(n14249) );
  OR U18616 ( .A(n14252), .B(n14253), .Z(n14248) );
  NAND U18617 ( .A(n14254), .B(n14255), .Z(n14211) );
  OR U18618 ( .A(n14256), .B(n14257), .Z(n14255) );
  OR U18619 ( .A(n14258), .B(n14259), .Z(n14254) );
  ANDN U18620 ( .B(n14260), .A(n14261), .Z(n14212) );
  IV U18621 ( .A(n14262), .Z(n14260) );
  ANDN U18622 ( .B(n14263), .A(n14264), .Z(n14204) );
  XOR U18623 ( .A(n14190), .B(n14265), .Z(n14202) );
  XOR U18624 ( .A(n14191), .B(n14192), .Z(n14265) );
  XOR U18625 ( .A(n14197), .B(n14266), .Z(n14192) );
  XOR U18626 ( .A(n14196), .B(n14199), .Z(n14266) );
  IV U18627 ( .A(n14198), .Z(n14199) );
  NAND U18628 ( .A(n14267), .B(n14268), .Z(n14198) );
  OR U18629 ( .A(n14269), .B(n14270), .Z(n14268) );
  OR U18630 ( .A(n14271), .B(n14272), .Z(n14267) );
  NAND U18631 ( .A(n14273), .B(n14274), .Z(n14196) );
  OR U18632 ( .A(n14275), .B(n14276), .Z(n14274) );
  OR U18633 ( .A(n14277), .B(n14278), .Z(n14273) );
  NOR U18634 ( .A(n14279), .B(n14280), .Z(n14197) );
  ANDN U18635 ( .B(n14281), .A(n14282), .Z(n14191) );
  IV U18636 ( .A(n14283), .Z(n14281) );
  XNOR U18637 ( .A(n14184), .B(n14284), .Z(n14190) );
  XNOR U18638 ( .A(n14183), .B(n14185), .Z(n14284) );
  NAND U18639 ( .A(n14285), .B(n14286), .Z(n14185) );
  OR U18640 ( .A(n14287), .B(n14288), .Z(n14286) );
  OR U18641 ( .A(n14289), .B(n14290), .Z(n14285) );
  NAND U18642 ( .A(n14291), .B(n14292), .Z(n14183) );
  OR U18643 ( .A(n14293), .B(n14294), .Z(n14292) );
  OR U18644 ( .A(n14295), .B(n14296), .Z(n14291) );
  ANDN U18645 ( .B(n14297), .A(n14298), .Z(n14184) );
  IV U18646 ( .A(n14299), .Z(n14297) );
  XNOR U18647 ( .A(n14264), .B(n14263), .Z(N28985) );
  XOR U18648 ( .A(n14283), .B(n14282), .Z(n14263) );
  XNOR U18649 ( .A(n14298), .B(n14299), .Z(n14282) );
  XNOR U18650 ( .A(n14293), .B(n14294), .Z(n14299) );
  XNOR U18651 ( .A(n14295), .B(n14296), .Z(n14294) );
  XNOR U18652 ( .A(y[2116]), .B(x[2116]), .Z(n14296) );
  XNOR U18653 ( .A(y[2117]), .B(x[2117]), .Z(n14295) );
  XNOR U18654 ( .A(y[2115]), .B(x[2115]), .Z(n14293) );
  XNOR U18655 ( .A(n14287), .B(n14288), .Z(n14298) );
  XNOR U18656 ( .A(y[2112]), .B(x[2112]), .Z(n14288) );
  XNOR U18657 ( .A(n14289), .B(n14290), .Z(n14287) );
  XNOR U18658 ( .A(y[2113]), .B(x[2113]), .Z(n14290) );
  XNOR U18659 ( .A(y[2114]), .B(x[2114]), .Z(n14289) );
  XNOR U18660 ( .A(n14280), .B(n14279), .Z(n14283) );
  XNOR U18661 ( .A(n14275), .B(n14276), .Z(n14279) );
  XNOR U18662 ( .A(y[2109]), .B(x[2109]), .Z(n14276) );
  XNOR U18663 ( .A(n14277), .B(n14278), .Z(n14275) );
  XNOR U18664 ( .A(y[2110]), .B(x[2110]), .Z(n14278) );
  XNOR U18665 ( .A(y[2111]), .B(x[2111]), .Z(n14277) );
  XNOR U18666 ( .A(n14269), .B(n14270), .Z(n14280) );
  XNOR U18667 ( .A(y[2106]), .B(x[2106]), .Z(n14270) );
  XNOR U18668 ( .A(n14271), .B(n14272), .Z(n14269) );
  XNOR U18669 ( .A(y[2107]), .B(x[2107]), .Z(n14272) );
  XNOR U18670 ( .A(y[2108]), .B(x[2108]), .Z(n14271) );
  XOR U18671 ( .A(n14245), .B(n14246), .Z(n14264) );
  XNOR U18672 ( .A(n14261), .B(n14262), .Z(n14246) );
  XNOR U18673 ( .A(n14256), .B(n14257), .Z(n14262) );
  XNOR U18674 ( .A(n14258), .B(n14259), .Z(n14257) );
  XNOR U18675 ( .A(y[2104]), .B(x[2104]), .Z(n14259) );
  XNOR U18676 ( .A(y[2105]), .B(x[2105]), .Z(n14258) );
  XNOR U18677 ( .A(y[2103]), .B(x[2103]), .Z(n14256) );
  XNOR U18678 ( .A(n14250), .B(n14251), .Z(n14261) );
  XNOR U18679 ( .A(y[2100]), .B(x[2100]), .Z(n14251) );
  XNOR U18680 ( .A(n14252), .B(n14253), .Z(n14250) );
  XNOR U18681 ( .A(y[2101]), .B(x[2101]), .Z(n14253) );
  XNOR U18682 ( .A(y[2102]), .B(x[2102]), .Z(n14252) );
  XOR U18683 ( .A(n14244), .B(n14243), .Z(n14245) );
  XNOR U18684 ( .A(n14239), .B(n14240), .Z(n14243) );
  XNOR U18685 ( .A(y[2097]), .B(x[2097]), .Z(n14240) );
  XNOR U18686 ( .A(n14241), .B(n14242), .Z(n14239) );
  XNOR U18687 ( .A(y[2098]), .B(x[2098]), .Z(n14242) );
  XNOR U18688 ( .A(y[2099]), .B(x[2099]), .Z(n14241) );
  XNOR U18689 ( .A(n14233), .B(n14234), .Z(n14244) );
  XNOR U18690 ( .A(y[2094]), .B(x[2094]), .Z(n14234) );
  XNOR U18691 ( .A(n14235), .B(n14236), .Z(n14233) );
  XNOR U18692 ( .A(y[2095]), .B(x[2095]), .Z(n14236) );
  XNOR U18693 ( .A(y[2096]), .B(x[2096]), .Z(n14235) );
  NAND U18694 ( .A(n14300), .B(n14301), .Z(N28977) );
  NANDN U18695 ( .A(n14302), .B(n14303), .Z(n14301) );
  OR U18696 ( .A(n14304), .B(n14305), .Z(n14303) );
  NAND U18697 ( .A(n14304), .B(n14305), .Z(n14300) );
  XOR U18698 ( .A(n14304), .B(n14306), .Z(N28976) );
  XNOR U18699 ( .A(n14302), .B(n14305), .Z(n14306) );
  AND U18700 ( .A(n14307), .B(n14308), .Z(n14305) );
  NANDN U18701 ( .A(n14309), .B(n14310), .Z(n14308) );
  NANDN U18702 ( .A(n14311), .B(n14312), .Z(n14310) );
  NANDN U18703 ( .A(n14312), .B(n14311), .Z(n14307) );
  NAND U18704 ( .A(n14313), .B(n14314), .Z(n14302) );
  NANDN U18705 ( .A(n14315), .B(n14316), .Z(n14314) );
  OR U18706 ( .A(n14317), .B(n14318), .Z(n14316) );
  NAND U18707 ( .A(n14318), .B(n14317), .Z(n14313) );
  AND U18708 ( .A(n14319), .B(n14320), .Z(n14304) );
  NANDN U18709 ( .A(n14321), .B(n14322), .Z(n14320) );
  NANDN U18710 ( .A(n14323), .B(n14324), .Z(n14322) );
  NANDN U18711 ( .A(n14324), .B(n14323), .Z(n14319) );
  XOR U18712 ( .A(n14318), .B(n14325), .Z(N28975) );
  XOR U18713 ( .A(n14315), .B(n14317), .Z(n14325) );
  XNOR U18714 ( .A(n14311), .B(n14326), .Z(n14317) );
  XNOR U18715 ( .A(n14309), .B(n14312), .Z(n14326) );
  NAND U18716 ( .A(n14327), .B(n14328), .Z(n14312) );
  NAND U18717 ( .A(n14329), .B(n14330), .Z(n14328) );
  OR U18718 ( .A(n14331), .B(n14332), .Z(n14329) );
  NANDN U18719 ( .A(n14333), .B(n14331), .Z(n14327) );
  IV U18720 ( .A(n14332), .Z(n14333) );
  NAND U18721 ( .A(n14334), .B(n14335), .Z(n14309) );
  NAND U18722 ( .A(n14336), .B(n14337), .Z(n14335) );
  NANDN U18723 ( .A(n14338), .B(n14339), .Z(n14336) );
  NANDN U18724 ( .A(n14339), .B(n14338), .Z(n14334) );
  AND U18725 ( .A(n14340), .B(n14341), .Z(n14311) );
  NAND U18726 ( .A(n14342), .B(n14343), .Z(n14341) );
  OR U18727 ( .A(n14344), .B(n14345), .Z(n14342) );
  NANDN U18728 ( .A(n14346), .B(n14344), .Z(n14340) );
  NAND U18729 ( .A(n14347), .B(n14348), .Z(n14315) );
  NANDN U18730 ( .A(n14349), .B(n14350), .Z(n14348) );
  OR U18731 ( .A(n14351), .B(n14352), .Z(n14350) );
  NANDN U18732 ( .A(n14353), .B(n14351), .Z(n14347) );
  IV U18733 ( .A(n14352), .Z(n14353) );
  XNOR U18734 ( .A(n14323), .B(n14354), .Z(n14318) );
  XNOR U18735 ( .A(n14321), .B(n14324), .Z(n14354) );
  NAND U18736 ( .A(n14355), .B(n14356), .Z(n14324) );
  NAND U18737 ( .A(n14357), .B(n14358), .Z(n14356) );
  OR U18738 ( .A(n14359), .B(n14360), .Z(n14357) );
  NANDN U18739 ( .A(n14361), .B(n14359), .Z(n14355) );
  IV U18740 ( .A(n14360), .Z(n14361) );
  NAND U18741 ( .A(n14362), .B(n14363), .Z(n14321) );
  NAND U18742 ( .A(n14364), .B(n14365), .Z(n14363) );
  NANDN U18743 ( .A(n14366), .B(n14367), .Z(n14364) );
  NANDN U18744 ( .A(n14367), .B(n14366), .Z(n14362) );
  AND U18745 ( .A(n14368), .B(n14369), .Z(n14323) );
  NAND U18746 ( .A(n14370), .B(n14371), .Z(n14369) );
  OR U18747 ( .A(n14372), .B(n14373), .Z(n14370) );
  NANDN U18748 ( .A(n14374), .B(n14372), .Z(n14368) );
  XNOR U18749 ( .A(n14349), .B(n14375), .Z(N28974) );
  XOR U18750 ( .A(n14351), .B(n14352), .Z(n14375) );
  XNOR U18751 ( .A(n14365), .B(n14376), .Z(n14352) );
  XOR U18752 ( .A(n14366), .B(n14367), .Z(n14376) );
  XOR U18753 ( .A(n14372), .B(n14377), .Z(n14367) );
  XOR U18754 ( .A(n14371), .B(n14374), .Z(n14377) );
  IV U18755 ( .A(n14373), .Z(n14374) );
  NAND U18756 ( .A(n14378), .B(n14379), .Z(n14373) );
  OR U18757 ( .A(n14380), .B(n14381), .Z(n14379) );
  OR U18758 ( .A(n14382), .B(n14383), .Z(n14378) );
  NAND U18759 ( .A(n14384), .B(n14385), .Z(n14371) );
  OR U18760 ( .A(n14386), .B(n14387), .Z(n14385) );
  OR U18761 ( .A(n14388), .B(n14389), .Z(n14384) );
  NOR U18762 ( .A(n14390), .B(n14391), .Z(n14372) );
  ANDN U18763 ( .B(n14392), .A(n14393), .Z(n14366) );
  XNOR U18764 ( .A(n14359), .B(n14394), .Z(n14365) );
  XNOR U18765 ( .A(n14358), .B(n14360), .Z(n14394) );
  NAND U18766 ( .A(n14395), .B(n14396), .Z(n14360) );
  OR U18767 ( .A(n14397), .B(n14398), .Z(n14396) );
  OR U18768 ( .A(n14399), .B(n14400), .Z(n14395) );
  NAND U18769 ( .A(n14401), .B(n14402), .Z(n14358) );
  OR U18770 ( .A(n14403), .B(n14404), .Z(n14402) );
  OR U18771 ( .A(n14405), .B(n14406), .Z(n14401) );
  ANDN U18772 ( .B(n14407), .A(n14408), .Z(n14359) );
  IV U18773 ( .A(n14409), .Z(n14407) );
  ANDN U18774 ( .B(n14410), .A(n14411), .Z(n14351) );
  XOR U18775 ( .A(n14337), .B(n14412), .Z(n14349) );
  XOR U18776 ( .A(n14338), .B(n14339), .Z(n14412) );
  XOR U18777 ( .A(n14344), .B(n14413), .Z(n14339) );
  XOR U18778 ( .A(n14343), .B(n14346), .Z(n14413) );
  IV U18779 ( .A(n14345), .Z(n14346) );
  NAND U18780 ( .A(n14414), .B(n14415), .Z(n14345) );
  OR U18781 ( .A(n14416), .B(n14417), .Z(n14415) );
  OR U18782 ( .A(n14418), .B(n14419), .Z(n14414) );
  NAND U18783 ( .A(n14420), .B(n14421), .Z(n14343) );
  OR U18784 ( .A(n14422), .B(n14423), .Z(n14421) );
  OR U18785 ( .A(n14424), .B(n14425), .Z(n14420) );
  NOR U18786 ( .A(n14426), .B(n14427), .Z(n14344) );
  ANDN U18787 ( .B(n14428), .A(n14429), .Z(n14338) );
  IV U18788 ( .A(n14430), .Z(n14428) );
  XNOR U18789 ( .A(n14331), .B(n14431), .Z(n14337) );
  XNOR U18790 ( .A(n14330), .B(n14332), .Z(n14431) );
  NAND U18791 ( .A(n14432), .B(n14433), .Z(n14332) );
  OR U18792 ( .A(n14434), .B(n14435), .Z(n14433) );
  OR U18793 ( .A(n14436), .B(n14437), .Z(n14432) );
  NAND U18794 ( .A(n14438), .B(n14439), .Z(n14330) );
  OR U18795 ( .A(n14440), .B(n14441), .Z(n14439) );
  OR U18796 ( .A(n14442), .B(n14443), .Z(n14438) );
  ANDN U18797 ( .B(n14444), .A(n14445), .Z(n14331) );
  IV U18798 ( .A(n14446), .Z(n14444) );
  XNOR U18799 ( .A(n14411), .B(n14410), .Z(N28973) );
  XOR U18800 ( .A(n14430), .B(n14429), .Z(n14410) );
  XNOR U18801 ( .A(n14445), .B(n14446), .Z(n14429) );
  XNOR U18802 ( .A(n14440), .B(n14441), .Z(n14446) );
  XNOR U18803 ( .A(n14442), .B(n14443), .Z(n14441) );
  XNOR U18804 ( .A(y[2092]), .B(x[2092]), .Z(n14443) );
  XNOR U18805 ( .A(y[2093]), .B(x[2093]), .Z(n14442) );
  XNOR U18806 ( .A(y[2091]), .B(x[2091]), .Z(n14440) );
  XNOR U18807 ( .A(n14434), .B(n14435), .Z(n14445) );
  XNOR U18808 ( .A(y[2088]), .B(x[2088]), .Z(n14435) );
  XNOR U18809 ( .A(n14436), .B(n14437), .Z(n14434) );
  XNOR U18810 ( .A(y[2089]), .B(x[2089]), .Z(n14437) );
  XNOR U18811 ( .A(y[2090]), .B(x[2090]), .Z(n14436) );
  XNOR U18812 ( .A(n14427), .B(n14426), .Z(n14430) );
  XNOR U18813 ( .A(n14422), .B(n14423), .Z(n14426) );
  XNOR U18814 ( .A(y[2085]), .B(x[2085]), .Z(n14423) );
  XNOR U18815 ( .A(n14424), .B(n14425), .Z(n14422) );
  XNOR U18816 ( .A(y[2086]), .B(x[2086]), .Z(n14425) );
  XNOR U18817 ( .A(y[2087]), .B(x[2087]), .Z(n14424) );
  XNOR U18818 ( .A(n14416), .B(n14417), .Z(n14427) );
  XNOR U18819 ( .A(y[2082]), .B(x[2082]), .Z(n14417) );
  XNOR U18820 ( .A(n14418), .B(n14419), .Z(n14416) );
  XNOR U18821 ( .A(y[2083]), .B(x[2083]), .Z(n14419) );
  XNOR U18822 ( .A(y[2084]), .B(x[2084]), .Z(n14418) );
  XOR U18823 ( .A(n14392), .B(n14393), .Z(n14411) );
  XNOR U18824 ( .A(n14408), .B(n14409), .Z(n14393) );
  XNOR U18825 ( .A(n14403), .B(n14404), .Z(n14409) );
  XNOR U18826 ( .A(n14405), .B(n14406), .Z(n14404) );
  XNOR U18827 ( .A(y[2080]), .B(x[2080]), .Z(n14406) );
  XNOR U18828 ( .A(y[2081]), .B(x[2081]), .Z(n14405) );
  XNOR U18829 ( .A(y[2079]), .B(x[2079]), .Z(n14403) );
  XNOR U18830 ( .A(n14397), .B(n14398), .Z(n14408) );
  XNOR U18831 ( .A(y[2076]), .B(x[2076]), .Z(n14398) );
  XNOR U18832 ( .A(n14399), .B(n14400), .Z(n14397) );
  XNOR U18833 ( .A(y[2077]), .B(x[2077]), .Z(n14400) );
  XNOR U18834 ( .A(y[2078]), .B(x[2078]), .Z(n14399) );
  XOR U18835 ( .A(n14391), .B(n14390), .Z(n14392) );
  XNOR U18836 ( .A(n14386), .B(n14387), .Z(n14390) );
  XNOR U18837 ( .A(y[2073]), .B(x[2073]), .Z(n14387) );
  XNOR U18838 ( .A(n14388), .B(n14389), .Z(n14386) );
  XNOR U18839 ( .A(y[2074]), .B(x[2074]), .Z(n14389) );
  XNOR U18840 ( .A(y[2075]), .B(x[2075]), .Z(n14388) );
  XNOR U18841 ( .A(n14380), .B(n14381), .Z(n14391) );
  XNOR U18842 ( .A(y[2070]), .B(x[2070]), .Z(n14381) );
  XNOR U18843 ( .A(n14382), .B(n14383), .Z(n14380) );
  XNOR U18844 ( .A(y[2071]), .B(x[2071]), .Z(n14383) );
  XNOR U18845 ( .A(y[2072]), .B(x[2072]), .Z(n14382) );
  NAND U18846 ( .A(n14447), .B(n14448), .Z(N28965) );
  NANDN U18847 ( .A(n14449), .B(n14450), .Z(n14448) );
  OR U18848 ( .A(n14451), .B(n14452), .Z(n14450) );
  NAND U18849 ( .A(n14451), .B(n14452), .Z(n14447) );
  XOR U18850 ( .A(n14451), .B(n14453), .Z(N28964) );
  XNOR U18851 ( .A(n14449), .B(n14452), .Z(n14453) );
  AND U18852 ( .A(n14454), .B(n14455), .Z(n14452) );
  NANDN U18853 ( .A(n14456), .B(n14457), .Z(n14455) );
  NANDN U18854 ( .A(n14458), .B(n14459), .Z(n14457) );
  NANDN U18855 ( .A(n14459), .B(n14458), .Z(n14454) );
  NAND U18856 ( .A(n14460), .B(n14461), .Z(n14449) );
  NANDN U18857 ( .A(n14462), .B(n14463), .Z(n14461) );
  OR U18858 ( .A(n14464), .B(n14465), .Z(n14463) );
  NAND U18859 ( .A(n14465), .B(n14464), .Z(n14460) );
  AND U18860 ( .A(n14466), .B(n14467), .Z(n14451) );
  NANDN U18861 ( .A(n14468), .B(n14469), .Z(n14467) );
  NANDN U18862 ( .A(n14470), .B(n14471), .Z(n14469) );
  NANDN U18863 ( .A(n14471), .B(n14470), .Z(n14466) );
  XOR U18864 ( .A(n14465), .B(n14472), .Z(N28963) );
  XOR U18865 ( .A(n14462), .B(n14464), .Z(n14472) );
  XNOR U18866 ( .A(n14458), .B(n14473), .Z(n14464) );
  XNOR U18867 ( .A(n14456), .B(n14459), .Z(n14473) );
  NAND U18868 ( .A(n14474), .B(n14475), .Z(n14459) );
  NAND U18869 ( .A(n14476), .B(n14477), .Z(n14475) );
  OR U18870 ( .A(n14478), .B(n14479), .Z(n14476) );
  NANDN U18871 ( .A(n14480), .B(n14478), .Z(n14474) );
  IV U18872 ( .A(n14479), .Z(n14480) );
  NAND U18873 ( .A(n14481), .B(n14482), .Z(n14456) );
  NAND U18874 ( .A(n14483), .B(n14484), .Z(n14482) );
  NANDN U18875 ( .A(n14485), .B(n14486), .Z(n14483) );
  NANDN U18876 ( .A(n14486), .B(n14485), .Z(n14481) );
  AND U18877 ( .A(n14487), .B(n14488), .Z(n14458) );
  NAND U18878 ( .A(n14489), .B(n14490), .Z(n14488) );
  OR U18879 ( .A(n14491), .B(n14492), .Z(n14489) );
  NANDN U18880 ( .A(n14493), .B(n14491), .Z(n14487) );
  NAND U18881 ( .A(n14494), .B(n14495), .Z(n14462) );
  NANDN U18882 ( .A(n14496), .B(n14497), .Z(n14495) );
  OR U18883 ( .A(n14498), .B(n14499), .Z(n14497) );
  NANDN U18884 ( .A(n14500), .B(n14498), .Z(n14494) );
  IV U18885 ( .A(n14499), .Z(n14500) );
  XNOR U18886 ( .A(n14470), .B(n14501), .Z(n14465) );
  XNOR U18887 ( .A(n14468), .B(n14471), .Z(n14501) );
  NAND U18888 ( .A(n14502), .B(n14503), .Z(n14471) );
  NAND U18889 ( .A(n14504), .B(n14505), .Z(n14503) );
  OR U18890 ( .A(n14506), .B(n14507), .Z(n14504) );
  NANDN U18891 ( .A(n14508), .B(n14506), .Z(n14502) );
  IV U18892 ( .A(n14507), .Z(n14508) );
  NAND U18893 ( .A(n14509), .B(n14510), .Z(n14468) );
  NAND U18894 ( .A(n14511), .B(n14512), .Z(n14510) );
  NANDN U18895 ( .A(n14513), .B(n14514), .Z(n14511) );
  NANDN U18896 ( .A(n14514), .B(n14513), .Z(n14509) );
  AND U18897 ( .A(n14515), .B(n14516), .Z(n14470) );
  NAND U18898 ( .A(n14517), .B(n14518), .Z(n14516) );
  OR U18899 ( .A(n14519), .B(n14520), .Z(n14517) );
  NANDN U18900 ( .A(n14521), .B(n14519), .Z(n14515) );
  XNOR U18901 ( .A(n14496), .B(n14522), .Z(N28962) );
  XOR U18902 ( .A(n14498), .B(n14499), .Z(n14522) );
  XNOR U18903 ( .A(n14512), .B(n14523), .Z(n14499) );
  XOR U18904 ( .A(n14513), .B(n14514), .Z(n14523) );
  XOR U18905 ( .A(n14519), .B(n14524), .Z(n14514) );
  XOR U18906 ( .A(n14518), .B(n14521), .Z(n14524) );
  IV U18907 ( .A(n14520), .Z(n14521) );
  NAND U18908 ( .A(n14525), .B(n14526), .Z(n14520) );
  OR U18909 ( .A(n14527), .B(n14528), .Z(n14526) );
  OR U18910 ( .A(n14529), .B(n14530), .Z(n14525) );
  NAND U18911 ( .A(n14531), .B(n14532), .Z(n14518) );
  OR U18912 ( .A(n14533), .B(n14534), .Z(n14532) );
  OR U18913 ( .A(n14535), .B(n14536), .Z(n14531) );
  NOR U18914 ( .A(n14537), .B(n14538), .Z(n14519) );
  ANDN U18915 ( .B(n14539), .A(n14540), .Z(n14513) );
  XNOR U18916 ( .A(n14506), .B(n14541), .Z(n14512) );
  XNOR U18917 ( .A(n14505), .B(n14507), .Z(n14541) );
  NAND U18918 ( .A(n14542), .B(n14543), .Z(n14507) );
  OR U18919 ( .A(n14544), .B(n14545), .Z(n14543) );
  OR U18920 ( .A(n14546), .B(n14547), .Z(n14542) );
  NAND U18921 ( .A(n14548), .B(n14549), .Z(n14505) );
  OR U18922 ( .A(n14550), .B(n14551), .Z(n14549) );
  OR U18923 ( .A(n14552), .B(n14553), .Z(n14548) );
  ANDN U18924 ( .B(n14554), .A(n14555), .Z(n14506) );
  IV U18925 ( .A(n14556), .Z(n14554) );
  ANDN U18926 ( .B(n14557), .A(n14558), .Z(n14498) );
  XOR U18927 ( .A(n14484), .B(n14559), .Z(n14496) );
  XOR U18928 ( .A(n14485), .B(n14486), .Z(n14559) );
  XOR U18929 ( .A(n14491), .B(n14560), .Z(n14486) );
  XOR U18930 ( .A(n14490), .B(n14493), .Z(n14560) );
  IV U18931 ( .A(n14492), .Z(n14493) );
  NAND U18932 ( .A(n14561), .B(n14562), .Z(n14492) );
  OR U18933 ( .A(n14563), .B(n14564), .Z(n14562) );
  OR U18934 ( .A(n14565), .B(n14566), .Z(n14561) );
  NAND U18935 ( .A(n14567), .B(n14568), .Z(n14490) );
  OR U18936 ( .A(n14569), .B(n14570), .Z(n14568) );
  OR U18937 ( .A(n14571), .B(n14572), .Z(n14567) );
  NOR U18938 ( .A(n14573), .B(n14574), .Z(n14491) );
  ANDN U18939 ( .B(n14575), .A(n14576), .Z(n14485) );
  IV U18940 ( .A(n14577), .Z(n14575) );
  XNOR U18941 ( .A(n14478), .B(n14578), .Z(n14484) );
  XNOR U18942 ( .A(n14477), .B(n14479), .Z(n14578) );
  NAND U18943 ( .A(n14579), .B(n14580), .Z(n14479) );
  OR U18944 ( .A(n14581), .B(n14582), .Z(n14580) );
  OR U18945 ( .A(n14583), .B(n14584), .Z(n14579) );
  NAND U18946 ( .A(n14585), .B(n14586), .Z(n14477) );
  OR U18947 ( .A(n14587), .B(n14588), .Z(n14586) );
  OR U18948 ( .A(n14589), .B(n14590), .Z(n14585) );
  ANDN U18949 ( .B(n14591), .A(n14592), .Z(n14478) );
  IV U18950 ( .A(n14593), .Z(n14591) );
  XNOR U18951 ( .A(n14558), .B(n14557), .Z(N28961) );
  XOR U18952 ( .A(n14577), .B(n14576), .Z(n14557) );
  XNOR U18953 ( .A(n14592), .B(n14593), .Z(n14576) );
  XNOR U18954 ( .A(n14587), .B(n14588), .Z(n14593) );
  XNOR U18955 ( .A(n14589), .B(n14590), .Z(n14588) );
  XNOR U18956 ( .A(y[2068]), .B(x[2068]), .Z(n14590) );
  XNOR U18957 ( .A(y[2069]), .B(x[2069]), .Z(n14589) );
  XNOR U18958 ( .A(y[2067]), .B(x[2067]), .Z(n14587) );
  XNOR U18959 ( .A(n14581), .B(n14582), .Z(n14592) );
  XNOR U18960 ( .A(y[2064]), .B(x[2064]), .Z(n14582) );
  XNOR U18961 ( .A(n14583), .B(n14584), .Z(n14581) );
  XNOR U18962 ( .A(y[2065]), .B(x[2065]), .Z(n14584) );
  XNOR U18963 ( .A(y[2066]), .B(x[2066]), .Z(n14583) );
  XNOR U18964 ( .A(n14574), .B(n14573), .Z(n14577) );
  XNOR U18965 ( .A(n14569), .B(n14570), .Z(n14573) );
  XNOR U18966 ( .A(y[2061]), .B(x[2061]), .Z(n14570) );
  XNOR U18967 ( .A(n14571), .B(n14572), .Z(n14569) );
  XNOR U18968 ( .A(y[2062]), .B(x[2062]), .Z(n14572) );
  XNOR U18969 ( .A(y[2063]), .B(x[2063]), .Z(n14571) );
  XNOR U18970 ( .A(n14563), .B(n14564), .Z(n14574) );
  XNOR U18971 ( .A(y[2058]), .B(x[2058]), .Z(n14564) );
  XNOR U18972 ( .A(n14565), .B(n14566), .Z(n14563) );
  XNOR U18973 ( .A(y[2059]), .B(x[2059]), .Z(n14566) );
  XNOR U18974 ( .A(y[2060]), .B(x[2060]), .Z(n14565) );
  XOR U18975 ( .A(n14539), .B(n14540), .Z(n14558) );
  XNOR U18976 ( .A(n14555), .B(n14556), .Z(n14540) );
  XNOR U18977 ( .A(n14550), .B(n14551), .Z(n14556) );
  XNOR U18978 ( .A(n14552), .B(n14553), .Z(n14551) );
  XNOR U18979 ( .A(y[2056]), .B(x[2056]), .Z(n14553) );
  XNOR U18980 ( .A(y[2057]), .B(x[2057]), .Z(n14552) );
  XNOR U18981 ( .A(y[2055]), .B(x[2055]), .Z(n14550) );
  XNOR U18982 ( .A(n14544), .B(n14545), .Z(n14555) );
  XNOR U18983 ( .A(y[2052]), .B(x[2052]), .Z(n14545) );
  XNOR U18984 ( .A(n14546), .B(n14547), .Z(n14544) );
  XNOR U18985 ( .A(y[2053]), .B(x[2053]), .Z(n14547) );
  XNOR U18986 ( .A(y[2054]), .B(x[2054]), .Z(n14546) );
  XOR U18987 ( .A(n14538), .B(n14537), .Z(n14539) );
  XNOR U18988 ( .A(n14533), .B(n14534), .Z(n14537) );
  XNOR U18989 ( .A(y[2049]), .B(x[2049]), .Z(n14534) );
  XNOR U18990 ( .A(n14535), .B(n14536), .Z(n14533) );
  XNOR U18991 ( .A(y[2050]), .B(x[2050]), .Z(n14536) );
  XNOR U18992 ( .A(y[2051]), .B(x[2051]), .Z(n14535) );
  XNOR U18993 ( .A(n14527), .B(n14528), .Z(n14538) );
  XNOR U18994 ( .A(y[2046]), .B(x[2046]), .Z(n14528) );
  XNOR U18995 ( .A(n14529), .B(n14530), .Z(n14527) );
  XNOR U18996 ( .A(y[2047]), .B(x[2047]), .Z(n14530) );
  XNOR U18997 ( .A(y[2048]), .B(x[2048]), .Z(n14529) );
  NAND U18998 ( .A(n14594), .B(n14595), .Z(N28953) );
  NANDN U18999 ( .A(n14596), .B(n14597), .Z(n14595) );
  OR U19000 ( .A(n14598), .B(n14599), .Z(n14597) );
  NAND U19001 ( .A(n14598), .B(n14599), .Z(n14594) );
  XOR U19002 ( .A(n14598), .B(n14600), .Z(N28952) );
  XNOR U19003 ( .A(n14596), .B(n14599), .Z(n14600) );
  AND U19004 ( .A(n14601), .B(n14602), .Z(n14599) );
  NANDN U19005 ( .A(n14603), .B(n14604), .Z(n14602) );
  NANDN U19006 ( .A(n14605), .B(n14606), .Z(n14604) );
  NANDN U19007 ( .A(n14606), .B(n14605), .Z(n14601) );
  NAND U19008 ( .A(n14607), .B(n14608), .Z(n14596) );
  NANDN U19009 ( .A(n14609), .B(n14610), .Z(n14608) );
  OR U19010 ( .A(n14611), .B(n14612), .Z(n14610) );
  NAND U19011 ( .A(n14612), .B(n14611), .Z(n14607) );
  AND U19012 ( .A(n14613), .B(n14614), .Z(n14598) );
  NANDN U19013 ( .A(n14615), .B(n14616), .Z(n14614) );
  NANDN U19014 ( .A(n14617), .B(n14618), .Z(n14616) );
  NANDN U19015 ( .A(n14618), .B(n14617), .Z(n14613) );
  XOR U19016 ( .A(n14612), .B(n14619), .Z(N28951) );
  XOR U19017 ( .A(n14609), .B(n14611), .Z(n14619) );
  XNOR U19018 ( .A(n14605), .B(n14620), .Z(n14611) );
  XNOR U19019 ( .A(n14603), .B(n14606), .Z(n14620) );
  NAND U19020 ( .A(n14621), .B(n14622), .Z(n14606) );
  NAND U19021 ( .A(n14623), .B(n14624), .Z(n14622) );
  OR U19022 ( .A(n14625), .B(n14626), .Z(n14623) );
  NANDN U19023 ( .A(n14627), .B(n14625), .Z(n14621) );
  IV U19024 ( .A(n14626), .Z(n14627) );
  NAND U19025 ( .A(n14628), .B(n14629), .Z(n14603) );
  NAND U19026 ( .A(n14630), .B(n14631), .Z(n14629) );
  NANDN U19027 ( .A(n14632), .B(n14633), .Z(n14630) );
  NANDN U19028 ( .A(n14633), .B(n14632), .Z(n14628) );
  AND U19029 ( .A(n14634), .B(n14635), .Z(n14605) );
  NAND U19030 ( .A(n14636), .B(n14637), .Z(n14635) );
  OR U19031 ( .A(n14638), .B(n14639), .Z(n14636) );
  NANDN U19032 ( .A(n14640), .B(n14638), .Z(n14634) );
  NAND U19033 ( .A(n14641), .B(n14642), .Z(n14609) );
  NANDN U19034 ( .A(n14643), .B(n14644), .Z(n14642) );
  OR U19035 ( .A(n14645), .B(n14646), .Z(n14644) );
  NANDN U19036 ( .A(n14647), .B(n14645), .Z(n14641) );
  IV U19037 ( .A(n14646), .Z(n14647) );
  XNOR U19038 ( .A(n14617), .B(n14648), .Z(n14612) );
  XNOR U19039 ( .A(n14615), .B(n14618), .Z(n14648) );
  NAND U19040 ( .A(n14649), .B(n14650), .Z(n14618) );
  NAND U19041 ( .A(n14651), .B(n14652), .Z(n14650) );
  OR U19042 ( .A(n14653), .B(n14654), .Z(n14651) );
  NANDN U19043 ( .A(n14655), .B(n14653), .Z(n14649) );
  IV U19044 ( .A(n14654), .Z(n14655) );
  NAND U19045 ( .A(n14656), .B(n14657), .Z(n14615) );
  NAND U19046 ( .A(n14658), .B(n14659), .Z(n14657) );
  NANDN U19047 ( .A(n14660), .B(n14661), .Z(n14658) );
  NANDN U19048 ( .A(n14661), .B(n14660), .Z(n14656) );
  AND U19049 ( .A(n14662), .B(n14663), .Z(n14617) );
  NAND U19050 ( .A(n14664), .B(n14665), .Z(n14663) );
  OR U19051 ( .A(n14666), .B(n14667), .Z(n14664) );
  NANDN U19052 ( .A(n14668), .B(n14666), .Z(n14662) );
  XNOR U19053 ( .A(n14643), .B(n14669), .Z(N28950) );
  XOR U19054 ( .A(n14645), .B(n14646), .Z(n14669) );
  XNOR U19055 ( .A(n14659), .B(n14670), .Z(n14646) );
  XOR U19056 ( .A(n14660), .B(n14661), .Z(n14670) );
  XOR U19057 ( .A(n14666), .B(n14671), .Z(n14661) );
  XOR U19058 ( .A(n14665), .B(n14668), .Z(n14671) );
  IV U19059 ( .A(n14667), .Z(n14668) );
  NAND U19060 ( .A(n14672), .B(n14673), .Z(n14667) );
  OR U19061 ( .A(n14674), .B(n14675), .Z(n14673) );
  OR U19062 ( .A(n14676), .B(n14677), .Z(n14672) );
  NAND U19063 ( .A(n14678), .B(n14679), .Z(n14665) );
  OR U19064 ( .A(n14680), .B(n14681), .Z(n14679) );
  OR U19065 ( .A(n14682), .B(n14683), .Z(n14678) );
  NOR U19066 ( .A(n14684), .B(n14685), .Z(n14666) );
  ANDN U19067 ( .B(n14686), .A(n14687), .Z(n14660) );
  XNOR U19068 ( .A(n14653), .B(n14688), .Z(n14659) );
  XNOR U19069 ( .A(n14652), .B(n14654), .Z(n14688) );
  NAND U19070 ( .A(n14689), .B(n14690), .Z(n14654) );
  OR U19071 ( .A(n14691), .B(n14692), .Z(n14690) );
  OR U19072 ( .A(n14693), .B(n14694), .Z(n14689) );
  NAND U19073 ( .A(n14695), .B(n14696), .Z(n14652) );
  OR U19074 ( .A(n14697), .B(n14698), .Z(n14696) );
  OR U19075 ( .A(n14699), .B(n14700), .Z(n14695) );
  ANDN U19076 ( .B(n14701), .A(n14702), .Z(n14653) );
  IV U19077 ( .A(n14703), .Z(n14701) );
  ANDN U19078 ( .B(n14704), .A(n14705), .Z(n14645) );
  XOR U19079 ( .A(n14631), .B(n14706), .Z(n14643) );
  XOR U19080 ( .A(n14632), .B(n14633), .Z(n14706) );
  XOR U19081 ( .A(n14638), .B(n14707), .Z(n14633) );
  XOR U19082 ( .A(n14637), .B(n14640), .Z(n14707) );
  IV U19083 ( .A(n14639), .Z(n14640) );
  NAND U19084 ( .A(n14708), .B(n14709), .Z(n14639) );
  OR U19085 ( .A(n14710), .B(n14711), .Z(n14709) );
  OR U19086 ( .A(n14712), .B(n14713), .Z(n14708) );
  NAND U19087 ( .A(n14714), .B(n14715), .Z(n14637) );
  OR U19088 ( .A(n14716), .B(n14717), .Z(n14715) );
  OR U19089 ( .A(n14718), .B(n14719), .Z(n14714) );
  NOR U19090 ( .A(n14720), .B(n14721), .Z(n14638) );
  ANDN U19091 ( .B(n14722), .A(n14723), .Z(n14632) );
  IV U19092 ( .A(n14724), .Z(n14722) );
  XNOR U19093 ( .A(n14625), .B(n14725), .Z(n14631) );
  XNOR U19094 ( .A(n14624), .B(n14626), .Z(n14725) );
  NAND U19095 ( .A(n14726), .B(n14727), .Z(n14626) );
  OR U19096 ( .A(n14728), .B(n14729), .Z(n14727) );
  OR U19097 ( .A(n14730), .B(n14731), .Z(n14726) );
  NAND U19098 ( .A(n14732), .B(n14733), .Z(n14624) );
  OR U19099 ( .A(n14734), .B(n14735), .Z(n14733) );
  OR U19100 ( .A(n14736), .B(n14737), .Z(n14732) );
  ANDN U19101 ( .B(n14738), .A(n14739), .Z(n14625) );
  IV U19102 ( .A(n14740), .Z(n14738) );
  XNOR U19103 ( .A(n14705), .B(n14704), .Z(N28949) );
  XOR U19104 ( .A(n14724), .B(n14723), .Z(n14704) );
  XNOR U19105 ( .A(n14739), .B(n14740), .Z(n14723) );
  XNOR U19106 ( .A(n14734), .B(n14735), .Z(n14740) );
  XNOR U19107 ( .A(n14736), .B(n14737), .Z(n14735) );
  XNOR U19108 ( .A(y[2044]), .B(x[2044]), .Z(n14737) );
  XNOR U19109 ( .A(y[2045]), .B(x[2045]), .Z(n14736) );
  XNOR U19110 ( .A(y[2043]), .B(x[2043]), .Z(n14734) );
  XNOR U19111 ( .A(n14728), .B(n14729), .Z(n14739) );
  XNOR U19112 ( .A(y[2040]), .B(x[2040]), .Z(n14729) );
  XNOR U19113 ( .A(n14730), .B(n14731), .Z(n14728) );
  XNOR U19114 ( .A(y[2041]), .B(x[2041]), .Z(n14731) );
  XNOR U19115 ( .A(y[2042]), .B(x[2042]), .Z(n14730) );
  XNOR U19116 ( .A(n14721), .B(n14720), .Z(n14724) );
  XNOR U19117 ( .A(n14716), .B(n14717), .Z(n14720) );
  XNOR U19118 ( .A(y[2037]), .B(x[2037]), .Z(n14717) );
  XNOR U19119 ( .A(n14718), .B(n14719), .Z(n14716) );
  XNOR U19120 ( .A(y[2038]), .B(x[2038]), .Z(n14719) );
  XNOR U19121 ( .A(y[2039]), .B(x[2039]), .Z(n14718) );
  XNOR U19122 ( .A(n14710), .B(n14711), .Z(n14721) );
  XNOR U19123 ( .A(y[2034]), .B(x[2034]), .Z(n14711) );
  XNOR U19124 ( .A(n14712), .B(n14713), .Z(n14710) );
  XNOR U19125 ( .A(y[2035]), .B(x[2035]), .Z(n14713) );
  XNOR U19126 ( .A(y[2036]), .B(x[2036]), .Z(n14712) );
  XOR U19127 ( .A(n14686), .B(n14687), .Z(n14705) );
  XNOR U19128 ( .A(n14702), .B(n14703), .Z(n14687) );
  XNOR U19129 ( .A(n14697), .B(n14698), .Z(n14703) );
  XNOR U19130 ( .A(n14699), .B(n14700), .Z(n14698) );
  XNOR U19131 ( .A(y[2032]), .B(x[2032]), .Z(n14700) );
  XNOR U19132 ( .A(y[2033]), .B(x[2033]), .Z(n14699) );
  XNOR U19133 ( .A(y[2031]), .B(x[2031]), .Z(n14697) );
  XNOR U19134 ( .A(n14691), .B(n14692), .Z(n14702) );
  XNOR U19135 ( .A(y[2028]), .B(x[2028]), .Z(n14692) );
  XNOR U19136 ( .A(n14693), .B(n14694), .Z(n14691) );
  XNOR U19137 ( .A(y[2029]), .B(x[2029]), .Z(n14694) );
  XNOR U19138 ( .A(y[2030]), .B(x[2030]), .Z(n14693) );
  XOR U19139 ( .A(n14685), .B(n14684), .Z(n14686) );
  XNOR U19140 ( .A(n14680), .B(n14681), .Z(n14684) );
  XNOR U19141 ( .A(y[2025]), .B(x[2025]), .Z(n14681) );
  XNOR U19142 ( .A(n14682), .B(n14683), .Z(n14680) );
  XNOR U19143 ( .A(y[2026]), .B(x[2026]), .Z(n14683) );
  XNOR U19144 ( .A(y[2027]), .B(x[2027]), .Z(n14682) );
  XNOR U19145 ( .A(n14674), .B(n14675), .Z(n14685) );
  XNOR U19146 ( .A(y[2022]), .B(x[2022]), .Z(n14675) );
  XNOR U19147 ( .A(n14676), .B(n14677), .Z(n14674) );
  XNOR U19148 ( .A(y[2023]), .B(x[2023]), .Z(n14677) );
  XNOR U19149 ( .A(y[2024]), .B(x[2024]), .Z(n14676) );
  NAND U19150 ( .A(n14741), .B(n14742), .Z(N28941) );
  NANDN U19151 ( .A(n14743), .B(n14744), .Z(n14742) );
  OR U19152 ( .A(n14745), .B(n14746), .Z(n14744) );
  NAND U19153 ( .A(n14745), .B(n14746), .Z(n14741) );
  XOR U19154 ( .A(n14745), .B(n14747), .Z(N28940) );
  XNOR U19155 ( .A(n14743), .B(n14746), .Z(n14747) );
  AND U19156 ( .A(n14748), .B(n14749), .Z(n14746) );
  NANDN U19157 ( .A(n14750), .B(n14751), .Z(n14749) );
  NANDN U19158 ( .A(n14752), .B(n14753), .Z(n14751) );
  NANDN U19159 ( .A(n14753), .B(n14752), .Z(n14748) );
  NAND U19160 ( .A(n14754), .B(n14755), .Z(n14743) );
  NANDN U19161 ( .A(n14756), .B(n14757), .Z(n14755) );
  OR U19162 ( .A(n14758), .B(n14759), .Z(n14757) );
  NAND U19163 ( .A(n14759), .B(n14758), .Z(n14754) );
  AND U19164 ( .A(n14760), .B(n14761), .Z(n14745) );
  NANDN U19165 ( .A(n14762), .B(n14763), .Z(n14761) );
  NANDN U19166 ( .A(n14764), .B(n14765), .Z(n14763) );
  NANDN U19167 ( .A(n14765), .B(n14764), .Z(n14760) );
  XOR U19168 ( .A(n14759), .B(n14766), .Z(N28939) );
  XOR U19169 ( .A(n14756), .B(n14758), .Z(n14766) );
  XNOR U19170 ( .A(n14752), .B(n14767), .Z(n14758) );
  XNOR U19171 ( .A(n14750), .B(n14753), .Z(n14767) );
  NAND U19172 ( .A(n14768), .B(n14769), .Z(n14753) );
  NAND U19173 ( .A(n14770), .B(n14771), .Z(n14769) );
  OR U19174 ( .A(n14772), .B(n14773), .Z(n14770) );
  NANDN U19175 ( .A(n14774), .B(n14772), .Z(n14768) );
  IV U19176 ( .A(n14773), .Z(n14774) );
  NAND U19177 ( .A(n14775), .B(n14776), .Z(n14750) );
  NAND U19178 ( .A(n14777), .B(n14778), .Z(n14776) );
  NANDN U19179 ( .A(n14779), .B(n14780), .Z(n14777) );
  NANDN U19180 ( .A(n14780), .B(n14779), .Z(n14775) );
  AND U19181 ( .A(n14781), .B(n14782), .Z(n14752) );
  NAND U19182 ( .A(n14783), .B(n14784), .Z(n14782) );
  OR U19183 ( .A(n14785), .B(n14786), .Z(n14783) );
  NANDN U19184 ( .A(n14787), .B(n14785), .Z(n14781) );
  NAND U19185 ( .A(n14788), .B(n14789), .Z(n14756) );
  NANDN U19186 ( .A(n14790), .B(n14791), .Z(n14789) );
  OR U19187 ( .A(n14792), .B(n14793), .Z(n14791) );
  NANDN U19188 ( .A(n14794), .B(n14792), .Z(n14788) );
  IV U19189 ( .A(n14793), .Z(n14794) );
  XNOR U19190 ( .A(n14764), .B(n14795), .Z(n14759) );
  XNOR U19191 ( .A(n14762), .B(n14765), .Z(n14795) );
  NAND U19192 ( .A(n14796), .B(n14797), .Z(n14765) );
  NAND U19193 ( .A(n14798), .B(n14799), .Z(n14797) );
  OR U19194 ( .A(n14800), .B(n14801), .Z(n14798) );
  NANDN U19195 ( .A(n14802), .B(n14800), .Z(n14796) );
  IV U19196 ( .A(n14801), .Z(n14802) );
  NAND U19197 ( .A(n14803), .B(n14804), .Z(n14762) );
  NAND U19198 ( .A(n14805), .B(n14806), .Z(n14804) );
  NANDN U19199 ( .A(n14807), .B(n14808), .Z(n14805) );
  NANDN U19200 ( .A(n14808), .B(n14807), .Z(n14803) );
  AND U19201 ( .A(n14809), .B(n14810), .Z(n14764) );
  NAND U19202 ( .A(n14811), .B(n14812), .Z(n14810) );
  OR U19203 ( .A(n14813), .B(n14814), .Z(n14811) );
  NANDN U19204 ( .A(n14815), .B(n14813), .Z(n14809) );
  XNOR U19205 ( .A(n14790), .B(n14816), .Z(N28938) );
  XOR U19206 ( .A(n14792), .B(n14793), .Z(n14816) );
  XNOR U19207 ( .A(n14806), .B(n14817), .Z(n14793) );
  XOR U19208 ( .A(n14807), .B(n14808), .Z(n14817) );
  XOR U19209 ( .A(n14813), .B(n14818), .Z(n14808) );
  XOR U19210 ( .A(n14812), .B(n14815), .Z(n14818) );
  IV U19211 ( .A(n14814), .Z(n14815) );
  NAND U19212 ( .A(n14819), .B(n14820), .Z(n14814) );
  OR U19213 ( .A(n14821), .B(n14822), .Z(n14820) );
  OR U19214 ( .A(n14823), .B(n14824), .Z(n14819) );
  NAND U19215 ( .A(n14825), .B(n14826), .Z(n14812) );
  OR U19216 ( .A(n14827), .B(n14828), .Z(n14826) );
  OR U19217 ( .A(n14829), .B(n14830), .Z(n14825) );
  NOR U19218 ( .A(n14831), .B(n14832), .Z(n14813) );
  ANDN U19219 ( .B(n14833), .A(n14834), .Z(n14807) );
  XNOR U19220 ( .A(n14800), .B(n14835), .Z(n14806) );
  XNOR U19221 ( .A(n14799), .B(n14801), .Z(n14835) );
  NAND U19222 ( .A(n14836), .B(n14837), .Z(n14801) );
  OR U19223 ( .A(n14838), .B(n14839), .Z(n14837) );
  OR U19224 ( .A(n14840), .B(n14841), .Z(n14836) );
  NAND U19225 ( .A(n14842), .B(n14843), .Z(n14799) );
  OR U19226 ( .A(n14844), .B(n14845), .Z(n14843) );
  OR U19227 ( .A(n14846), .B(n14847), .Z(n14842) );
  ANDN U19228 ( .B(n14848), .A(n14849), .Z(n14800) );
  IV U19229 ( .A(n14850), .Z(n14848) );
  ANDN U19230 ( .B(n14851), .A(n14852), .Z(n14792) );
  XOR U19231 ( .A(n14778), .B(n14853), .Z(n14790) );
  XOR U19232 ( .A(n14779), .B(n14780), .Z(n14853) );
  XOR U19233 ( .A(n14785), .B(n14854), .Z(n14780) );
  XOR U19234 ( .A(n14784), .B(n14787), .Z(n14854) );
  IV U19235 ( .A(n14786), .Z(n14787) );
  NAND U19236 ( .A(n14855), .B(n14856), .Z(n14786) );
  OR U19237 ( .A(n14857), .B(n14858), .Z(n14856) );
  OR U19238 ( .A(n14859), .B(n14860), .Z(n14855) );
  NAND U19239 ( .A(n14861), .B(n14862), .Z(n14784) );
  OR U19240 ( .A(n14863), .B(n14864), .Z(n14862) );
  OR U19241 ( .A(n14865), .B(n14866), .Z(n14861) );
  NOR U19242 ( .A(n14867), .B(n14868), .Z(n14785) );
  ANDN U19243 ( .B(n14869), .A(n14870), .Z(n14779) );
  IV U19244 ( .A(n14871), .Z(n14869) );
  XNOR U19245 ( .A(n14772), .B(n14872), .Z(n14778) );
  XNOR U19246 ( .A(n14771), .B(n14773), .Z(n14872) );
  NAND U19247 ( .A(n14873), .B(n14874), .Z(n14773) );
  OR U19248 ( .A(n14875), .B(n14876), .Z(n14874) );
  OR U19249 ( .A(n14877), .B(n14878), .Z(n14873) );
  NAND U19250 ( .A(n14879), .B(n14880), .Z(n14771) );
  OR U19251 ( .A(n14881), .B(n14882), .Z(n14880) );
  OR U19252 ( .A(n14883), .B(n14884), .Z(n14879) );
  ANDN U19253 ( .B(n14885), .A(n14886), .Z(n14772) );
  IV U19254 ( .A(n14887), .Z(n14885) );
  XNOR U19255 ( .A(n14852), .B(n14851), .Z(N28937) );
  XOR U19256 ( .A(n14871), .B(n14870), .Z(n14851) );
  XNOR U19257 ( .A(n14886), .B(n14887), .Z(n14870) );
  XNOR U19258 ( .A(n14881), .B(n14882), .Z(n14887) );
  XNOR U19259 ( .A(n14883), .B(n14884), .Z(n14882) );
  XNOR U19260 ( .A(y[2020]), .B(x[2020]), .Z(n14884) );
  XNOR U19261 ( .A(y[2021]), .B(x[2021]), .Z(n14883) );
  XNOR U19262 ( .A(y[2019]), .B(x[2019]), .Z(n14881) );
  XNOR U19263 ( .A(n14875), .B(n14876), .Z(n14886) );
  XNOR U19264 ( .A(y[2016]), .B(x[2016]), .Z(n14876) );
  XNOR U19265 ( .A(n14877), .B(n14878), .Z(n14875) );
  XNOR U19266 ( .A(y[2017]), .B(x[2017]), .Z(n14878) );
  XNOR U19267 ( .A(y[2018]), .B(x[2018]), .Z(n14877) );
  XNOR U19268 ( .A(n14868), .B(n14867), .Z(n14871) );
  XNOR U19269 ( .A(n14863), .B(n14864), .Z(n14867) );
  XNOR U19270 ( .A(y[2013]), .B(x[2013]), .Z(n14864) );
  XNOR U19271 ( .A(n14865), .B(n14866), .Z(n14863) );
  XNOR U19272 ( .A(y[2014]), .B(x[2014]), .Z(n14866) );
  XNOR U19273 ( .A(y[2015]), .B(x[2015]), .Z(n14865) );
  XNOR U19274 ( .A(n14857), .B(n14858), .Z(n14868) );
  XNOR U19275 ( .A(y[2010]), .B(x[2010]), .Z(n14858) );
  XNOR U19276 ( .A(n14859), .B(n14860), .Z(n14857) );
  XNOR U19277 ( .A(y[2011]), .B(x[2011]), .Z(n14860) );
  XNOR U19278 ( .A(y[2012]), .B(x[2012]), .Z(n14859) );
  XOR U19279 ( .A(n14833), .B(n14834), .Z(n14852) );
  XNOR U19280 ( .A(n14849), .B(n14850), .Z(n14834) );
  XNOR U19281 ( .A(n14844), .B(n14845), .Z(n14850) );
  XNOR U19282 ( .A(n14846), .B(n14847), .Z(n14845) );
  XNOR U19283 ( .A(y[2008]), .B(x[2008]), .Z(n14847) );
  XNOR U19284 ( .A(y[2009]), .B(x[2009]), .Z(n14846) );
  XNOR U19285 ( .A(y[2007]), .B(x[2007]), .Z(n14844) );
  XNOR U19286 ( .A(n14838), .B(n14839), .Z(n14849) );
  XNOR U19287 ( .A(y[2004]), .B(x[2004]), .Z(n14839) );
  XNOR U19288 ( .A(n14840), .B(n14841), .Z(n14838) );
  XNOR U19289 ( .A(y[2005]), .B(x[2005]), .Z(n14841) );
  XNOR U19290 ( .A(y[2006]), .B(x[2006]), .Z(n14840) );
  XOR U19291 ( .A(n14832), .B(n14831), .Z(n14833) );
  XNOR U19292 ( .A(n14827), .B(n14828), .Z(n14831) );
  XNOR U19293 ( .A(y[2001]), .B(x[2001]), .Z(n14828) );
  XNOR U19294 ( .A(n14829), .B(n14830), .Z(n14827) );
  XNOR U19295 ( .A(y[2002]), .B(x[2002]), .Z(n14830) );
  XNOR U19296 ( .A(y[2003]), .B(x[2003]), .Z(n14829) );
  XNOR U19297 ( .A(n14821), .B(n14822), .Z(n14832) );
  XNOR U19298 ( .A(y[1998]), .B(x[1998]), .Z(n14822) );
  XNOR U19299 ( .A(n14823), .B(n14824), .Z(n14821) );
  XNOR U19300 ( .A(y[1999]), .B(x[1999]), .Z(n14824) );
  XNOR U19301 ( .A(y[2000]), .B(x[2000]), .Z(n14823) );
  NAND U19302 ( .A(n14888), .B(n14889), .Z(N28929) );
  NANDN U19303 ( .A(n14890), .B(n14891), .Z(n14889) );
  OR U19304 ( .A(n14892), .B(n14893), .Z(n14891) );
  NAND U19305 ( .A(n14892), .B(n14893), .Z(n14888) );
  XOR U19306 ( .A(n14892), .B(n14894), .Z(N28928) );
  XNOR U19307 ( .A(n14890), .B(n14893), .Z(n14894) );
  AND U19308 ( .A(n14895), .B(n14896), .Z(n14893) );
  NANDN U19309 ( .A(n14897), .B(n14898), .Z(n14896) );
  NANDN U19310 ( .A(n14899), .B(n14900), .Z(n14898) );
  NANDN U19311 ( .A(n14900), .B(n14899), .Z(n14895) );
  NAND U19312 ( .A(n14901), .B(n14902), .Z(n14890) );
  NANDN U19313 ( .A(n14903), .B(n14904), .Z(n14902) );
  OR U19314 ( .A(n14905), .B(n14906), .Z(n14904) );
  NAND U19315 ( .A(n14906), .B(n14905), .Z(n14901) );
  AND U19316 ( .A(n14907), .B(n14908), .Z(n14892) );
  NANDN U19317 ( .A(n14909), .B(n14910), .Z(n14908) );
  NANDN U19318 ( .A(n14911), .B(n14912), .Z(n14910) );
  NANDN U19319 ( .A(n14912), .B(n14911), .Z(n14907) );
  XOR U19320 ( .A(n14906), .B(n14913), .Z(N28927) );
  XOR U19321 ( .A(n14903), .B(n14905), .Z(n14913) );
  XNOR U19322 ( .A(n14899), .B(n14914), .Z(n14905) );
  XNOR U19323 ( .A(n14897), .B(n14900), .Z(n14914) );
  NAND U19324 ( .A(n14915), .B(n14916), .Z(n14900) );
  NAND U19325 ( .A(n14917), .B(n14918), .Z(n14916) );
  OR U19326 ( .A(n14919), .B(n14920), .Z(n14917) );
  NANDN U19327 ( .A(n14921), .B(n14919), .Z(n14915) );
  IV U19328 ( .A(n14920), .Z(n14921) );
  NAND U19329 ( .A(n14922), .B(n14923), .Z(n14897) );
  NAND U19330 ( .A(n14924), .B(n14925), .Z(n14923) );
  NANDN U19331 ( .A(n14926), .B(n14927), .Z(n14924) );
  NANDN U19332 ( .A(n14927), .B(n14926), .Z(n14922) );
  AND U19333 ( .A(n14928), .B(n14929), .Z(n14899) );
  NAND U19334 ( .A(n14930), .B(n14931), .Z(n14929) );
  OR U19335 ( .A(n14932), .B(n14933), .Z(n14930) );
  NANDN U19336 ( .A(n14934), .B(n14932), .Z(n14928) );
  NAND U19337 ( .A(n14935), .B(n14936), .Z(n14903) );
  NANDN U19338 ( .A(n14937), .B(n14938), .Z(n14936) );
  OR U19339 ( .A(n14939), .B(n14940), .Z(n14938) );
  NANDN U19340 ( .A(n14941), .B(n14939), .Z(n14935) );
  IV U19341 ( .A(n14940), .Z(n14941) );
  XNOR U19342 ( .A(n14911), .B(n14942), .Z(n14906) );
  XNOR U19343 ( .A(n14909), .B(n14912), .Z(n14942) );
  NAND U19344 ( .A(n14943), .B(n14944), .Z(n14912) );
  NAND U19345 ( .A(n14945), .B(n14946), .Z(n14944) );
  OR U19346 ( .A(n14947), .B(n14948), .Z(n14945) );
  NANDN U19347 ( .A(n14949), .B(n14947), .Z(n14943) );
  IV U19348 ( .A(n14948), .Z(n14949) );
  NAND U19349 ( .A(n14950), .B(n14951), .Z(n14909) );
  NAND U19350 ( .A(n14952), .B(n14953), .Z(n14951) );
  NANDN U19351 ( .A(n14954), .B(n14955), .Z(n14952) );
  NANDN U19352 ( .A(n14955), .B(n14954), .Z(n14950) );
  AND U19353 ( .A(n14956), .B(n14957), .Z(n14911) );
  NAND U19354 ( .A(n14958), .B(n14959), .Z(n14957) );
  OR U19355 ( .A(n14960), .B(n14961), .Z(n14958) );
  NANDN U19356 ( .A(n14962), .B(n14960), .Z(n14956) );
  XNOR U19357 ( .A(n14937), .B(n14963), .Z(N28926) );
  XOR U19358 ( .A(n14939), .B(n14940), .Z(n14963) );
  XNOR U19359 ( .A(n14953), .B(n14964), .Z(n14940) );
  XOR U19360 ( .A(n14954), .B(n14955), .Z(n14964) );
  XOR U19361 ( .A(n14960), .B(n14965), .Z(n14955) );
  XOR U19362 ( .A(n14959), .B(n14962), .Z(n14965) );
  IV U19363 ( .A(n14961), .Z(n14962) );
  NAND U19364 ( .A(n14966), .B(n14967), .Z(n14961) );
  OR U19365 ( .A(n14968), .B(n14969), .Z(n14967) );
  OR U19366 ( .A(n14970), .B(n14971), .Z(n14966) );
  NAND U19367 ( .A(n14972), .B(n14973), .Z(n14959) );
  OR U19368 ( .A(n14974), .B(n14975), .Z(n14973) );
  OR U19369 ( .A(n14976), .B(n14977), .Z(n14972) );
  NOR U19370 ( .A(n14978), .B(n14979), .Z(n14960) );
  ANDN U19371 ( .B(n14980), .A(n14981), .Z(n14954) );
  XNOR U19372 ( .A(n14947), .B(n14982), .Z(n14953) );
  XNOR U19373 ( .A(n14946), .B(n14948), .Z(n14982) );
  NAND U19374 ( .A(n14983), .B(n14984), .Z(n14948) );
  OR U19375 ( .A(n14985), .B(n14986), .Z(n14984) );
  OR U19376 ( .A(n14987), .B(n14988), .Z(n14983) );
  NAND U19377 ( .A(n14989), .B(n14990), .Z(n14946) );
  OR U19378 ( .A(n14991), .B(n14992), .Z(n14990) );
  OR U19379 ( .A(n14993), .B(n14994), .Z(n14989) );
  ANDN U19380 ( .B(n14995), .A(n14996), .Z(n14947) );
  IV U19381 ( .A(n14997), .Z(n14995) );
  ANDN U19382 ( .B(n14998), .A(n14999), .Z(n14939) );
  XOR U19383 ( .A(n14925), .B(n15000), .Z(n14937) );
  XOR U19384 ( .A(n14926), .B(n14927), .Z(n15000) );
  XOR U19385 ( .A(n14932), .B(n15001), .Z(n14927) );
  XOR U19386 ( .A(n14931), .B(n14934), .Z(n15001) );
  IV U19387 ( .A(n14933), .Z(n14934) );
  NAND U19388 ( .A(n15002), .B(n15003), .Z(n14933) );
  OR U19389 ( .A(n15004), .B(n15005), .Z(n15003) );
  OR U19390 ( .A(n15006), .B(n15007), .Z(n15002) );
  NAND U19391 ( .A(n15008), .B(n15009), .Z(n14931) );
  OR U19392 ( .A(n15010), .B(n15011), .Z(n15009) );
  OR U19393 ( .A(n15012), .B(n15013), .Z(n15008) );
  NOR U19394 ( .A(n15014), .B(n15015), .Z(n14932) );
  ANDN U19395 ( .B(n15016), .A(n15017), .Z(n14926) );
  IV U19396 ( .A(n15018), .Z(n15016) );
  XNOR U19397 ( .A(n14919), .B(n15019), .Z(n14925) );
  XNOR U19398 ( .A(n14918), .B(n14920), .Z(n15019) );
  NAND U19399 ( .A(n15020), .B(n15021), .Z(n14920) );
  OR U19400 ( .A(n15022), .B(n15023), .Z(n15021) );
  OR U19401 ( .A(n15024), .B(n15025), .Z(n15020) );
  NAND U19402 ( .A(n15026), .B(n15027), .Z(n14918) );
  OR U19403 ( .A(n15028), .B(n15029), .Z(n15027) );
  OR U19404 ( .A(n15030), .B(n15031), .Z(n15026) );
  ANDN U19405 ( .B(n15032), .A(n15033), .Z(n14919) );
  IV U19406 ( .A(n15034), .Z(n15032) );
  XNOR U19407 ( .A(n14999), .B(n14998), .Z(N28925) );
  XOR U19408 ( .A(n15018), .B(n15017), .Z(n14998) );
  XNOR U19409 ( .A(n15033), .B(n15034), .Z(n15017) );
  XNOR U19410 ( .A(n15028), .B(n15029), .Z(n15034) );
  XNOR U19411 ( .A(n15030), .B(n15031), .Z(n15029) );
  XNOR U19412 ( .A(y[1996]), .B(x[1996]), .Z(n15031) );
  XNOR U19413 ( .A(y[1997]), .B(x[1997]), .Z(n15030) );
  XNOR U19414 ( .A(y[1995]), .B(x[1995]), .Z(n15028) );
  XNOR U19415 ( .A(n15022), .B(n15023), .Z(n15033) );
  XNOR U19416 ( .A(y[1992]), .B(x[1992]), .Z(n15023) );
  XNOR U19417 ( .A(n15024), .B(n15025), .Z(n15022) );
  XNOR U19418 ( .A(y[1993]), .B(x[1993]), .Z(n15025) );
  XNOR U19419 ( .A(y[1994]), .B(x[1994]), .Z(n15024) );
  XNOR U19420 ( .A(n15015), .B(n15014), .Z(n15018) );
  XNOR U19421 ( .A(n15010), .B(n15011), .Z(n15014) );
  XNOR U19422 ( .A(y[1989]), .B(x[1989]), .Z(n15011) );
  XNOR U19423 ( .A(n15012), .B(n15013), .Z(n15010) );
  XNOR U19424 ( .A(y[1990]), .B(x[1990]), .Z(n15013) );
  XNOR U19425 ( .A(y[1991]), .B(x[1991]), .Z(n15012) );
  XNOR U19426 ( .A(n15004), .B(n15005), .Z(n15015) );
  XNOR U19427 ( .A(y[1986]), .B(x[1986]), .Z(n15005) );
  XNOR U19428 ( .A(n15006), .B(n15007), .Z(n15004) );
  XNOR U19429 ( .A(y[1987]), .B(x[1987]), .Z(n15007) );
  XNOR U19430 ( .A(y[1988]), .B(x[1988]), .Z(n15006) );
  XOR U19431 ( .A(n14980), .B(n14981), .Z(n14999) );
  XNOR U19432 ( .A(n14996), .B(n14997), .Z(n14981) );
  XNOR U19433 ( .A(n14991), .B(n14992), .Z(n14997) );
  XNOR U19434 ( .A(n14993), .B(n14994), .Z(n14992) );
  XNOR U19435 ( .A(y[1984]), .B(x[1984]), .Z(n14994) );
  XNOR U19436 ( .A(y[1985]), .B(x[1985]), .Z(n14993) );
  XNOR U19437 ( .A(y[1983]), .B(x[1983]), .Z(n14991) );
  XNOR U19438 ( .A(n14985), .B(n14986), .Z(n14996) );
  XNOR U19439 ( .A(y[1980]), .B(x[1980]), .Z(n14986) );
  XNOR U19440 ( .A(n14987), .B(n14988), .Z(n14985) );
  XNOR U19441 ( .A(y[1981]), .B(x[1981]), .Z(n14988) );
  XNOR U19442 ( .A(y[1982]), .B(x[1982]), .Z(n14987) );
  XOR U19443 ( .A(n14979), .B(n14978), .Z(n14980) );
  XNOR U19444 ( .A(n14974), .B(n14975), .Z(n14978) );
  XNOR U19445 ( .A(y[1977]), .B(x[1977]), .Z(n14975) );
  XNOR U19446 ( .A(n14976), .B(n14977), .Z(n14974) );
  XNOR U19447 ( .A(y[1978]), .B(x[1978]), .Z(n14977) );
  XNOR U19448 ( .A(y[1979]), .B(x[1979]), .Z(n14976) );
  XNOR U19449 ( .A(n14968), .B(n14969), .Z(n14979) );
  XNOR U19450 ( .A(y[1974]), .B(x[1974]), .Z(n14969) );
  XNOR U19451 ( .A(n14970), .B(n14971), .Z(n14968) );
  XNOR U19452 ( .A(y[1975]), .B(x[1975]), .Z(n14971) );
  XNOR U19453 ( .A(y[1976]), .B(x[1976]), .Z(n14970) );
  NAND U19454 ( .A(n15035), .B(n15036), .Z(N28917) );
  NANDN U19455 ( .A(n15037), .B(n15038), .Z(n15036) );
  OR U19456 ( .A(n15039), .B(n15040), .Z(n15038) );
  NAND U19457 ( .A(n15039), .B(n15040), .Z(n15035) );
  XOR U19458 ( .A(n15039), .B(n15041), .Z(N28916) );
  XNOR U19459 ( .A(n15037), .B(n15040), .Z(n15041) );
  AND U19460 ( .A(n15042), .B(n15043), .Z(n15040) );
  NANDN U19461 ( .A(n15044), .B(n15045), .Z(n15043) );
  NANDN U19462 ( .A(n15046), .B(n15047), .Z(n15045) );
  NANDN U19463 ( .A(n15047), .B(n15046), .Z(n15042) );
  NAND U19464 ( .A(n15048), .B(n15049), .Z(n15037) );
  NANDN U19465 ( .A(n15050), .B(n15051), .Z(n15049) );
  OR U19466 ( .A(n15052), .B(n15053), .Z(n15051) );
  NAND U19467 ( .A(n15053), .B(n15052), .Z(n15048) );
  AND U19468 ( .A(n15054), .B(n15055), .Z(n15039) );
  NANDN U19469 ( .A(n15056), .B(n15057), .Z(n15055) );
  NANDN U19470 ( .A(n15058), .B(n15059), .Z(n15057) );
  NANDN U19471 ( .A(n15059), .B(n15058), .Z(n15054) );
  XOR U19472 ( .A(n15053), .B(n15060), .Z(N28915) );
  XOR U19473 ( .A(n15050), .B(n15052), .Z(n15060) );
  XNOR U19474 ( .A(n15046), .B(n15061), .Z(n15052) );
  XNOR U19475 ( .A(n15044), .B(n15047), .Z(n15061) );
  NAND U19476 ( .A(n15062), .B(n15063), .Z(n15047) );
  NAND U19477 ( .A(n15064), .B(n15065), .Z(n15063) );
  OR U19478 ( .A(n15066), .B(n15067), .Z(n15064) );
  NANDN U19479 ( .A(n15068), .B(n15066), .Z(n15062) );
  IV U19480 ( .A(n15067), .Z(n15068) );
  NAND U19481 ( .A(n15069), .B(n15070), .Z(n15044) );
  NAND U19482 ( .A(n15071), .B(n15072), .Z(n15070) );
  NANDN U19483 ( .A(n15073), .B(n15074), .Z(n15071) );
  NANDN U19484 ( .A(n15074), .B(n15073), .Z(n15069) );
  AND U19485 ( .A(n15075), .B(n15076), .Z(n15046) );
  NAND U19486 ( .A(n15077), .B(n15078), .Z(n15076) );
  OR U19487 ( .A(n15079), .B(n15080), .Z(n15077) );
  NANDN U19488 ( .A(n15081), .B(n15079), .Z(n15075) );
  NAND U19489 ( .A(n15082), .B(n15083), .Z(n15050) );
  NANDN U19490 ( .A(n15084), .B(n15085), .Z(n15083) );
  OR U19491 ( .A(n15086), .B(n15087), .Z(n15085) );
  NANDN U19492 ( .A(n15088), .B(n15086), .Z(n15082) );
  IV U19493 ( .A(n15087), .Z(n15088) );
  XNOR U19494 ( .A(n15058), .B(n15089), .Z(n15053) );
  XNOR U19495 ( .A(n15056), .B(n15059), .Z(n15089) );
  NAND U19496 ( .A(n15090), .B(n15091), .Z(n15059) );
  NAND U19497 ( .A(n15092), .B(n15093), .Z(n15091) );
  OR U19498 ( .A(n15094), .B(n15095), .Z(n15092) );
  NANDN U19499 ( .A(n15096), .B(n15094), .Z(n15090) );
  IV U19500 ( .A(n15095), .Z(n15096) );
  NAND U19501 ( .A(n15097), .B(n15098), .Z(n15056) );
  NAND U19502 ( .A(n15099), .B(n15100), .Z(n15098) );
  NANDN U19503 ( .A(n15101), .B(n15102), .Z(n15099) );
  NANDN U19504 ( .A(n15102), .B(n15101), .Z(n15097) );
  AND U19505 ( .A(n15103), .B(n15104), .Z(n15058) );
  NAND U19506 ( .A(n15105), .B(n15106), .Z(n15104) );
  OR U19507 ( .A(n15107), .B(n15108), .Z(n15105) );
  NANDN U19508 ( .A(n15109), .B(n15107), .Z(n15103) );
  XNOR U19509 ( .A(n15084), .B(n15110), .Z(N28914) );
  XOR U19510 ( .A(n15086), .B(n15087), .Z(n15110) );
  XNOR U19511 ( .A(n15100), .B(n15111), .Z(n15087) );
  XOR U19512 ( .A(n15101), .B(n15102), .Z(n15111) );
  XOR U19513 ( .A(n15107), .B(n15112), .Z(n15102) );
  XOR U19514 ( .A(n15106), .B(n15109), .Z(n15112) );
  IV U19515 ( .A(n15108), .Z(n15109) );
  NAND U19516 ( .A(n15113), .B(n15114), .Z(n15108) );
  OR U19517 ( .A(n15115), .B(n15116), .Z(n15114) );
  OR U19518 ( .A(n15117), .B(n15118), .Z(n15113) );
  NAND U19519 ( .A(n15119), .B(n15120), .Z(n15106) );
  OR U19520 ( .A(n15121), .B(n15122), .Z(n15120) );
  OR U19521 ( .A(n15123), .B(n15124), .Z(n15119) );
  NOR U19522 ( .A(n15125), .B(n15126), .Z(n15107) );
  ANDN U19523 ( .B(n15127), .A(n15128), .Z(n15101) );
  XNOR U19524 ( .A(n15094), .B(n15129), .Z(n15100) );
  XNOR U19525 ( .A(n15093), .B(n15095), .Z(n15129) );
  NAND U19526 ( .A(n15130), .B(n15131), .Z(n15095) );
  OR U19527 ( .A(n15132), .B(n15133), .Z(n15131) );
  OR U19528 ( .A(n15134), .B(n15135), .Z(n15130) );
  NAND U19529 ( .A(n15136), .B(n15137), .Z(n15093) );
  OR U19530 ( .A(n15138), .B(n15139), .Z(n15137) );
  OR U19531 ( .A(n15140), .B(n15141), .Z(n15136) );
  ANDN U19532 ( .B(n15142), .A(n15143), .Z(n15094) );
  IV U19533 ( .A(n15144), .Z(n15142) );
  ANDN U19534 ( .B(n15145), .A(n15146), .Z(n15086) );
  XOR U19535 ( .A(n15072), .B(n15147), .Z(n15084) );
  XOR U19536 ( .A(n15073), .B(n15074), .Z(n15147) );
  XOR U19537 ( .A(n15079), .B(n15148), .Z(n15074) );
  XOR U19538 ( .A(n15078), .B(n15081), .Z(n15148) );
  IV U19539 ( .A(n15080), .Z(n15081) );
  NAND U19540 ( .A(n15149), .B(n15150), .Z(n15080) );
  OR U19541 ( .A(n15151), .B(n15152), .Z(n15150) );
  OR U19542 ( .A(n15153), .B(n15154), .Z(n15149) );
  NAND U19543 ( .A(n15155), .B(n15156), .Z(n15078) );
  OR U19544 ( .A(n15157), .B(n15158), .Z(n15156) );
  OR U19545 ( .A(n15159), .B(n15160), .Z(n15155) );
  NOR U19546 ( .A(n15161), .B(n15162), .Z(n15079) );
  ANDN U19547 ( .B(n15163), .A(n15164), .Z(n15073) );
  IV U19548 ( .A(n15165), .Z(n15163) );
  XNOR U19549 ( .A(n15066), .B(n15166), .Z(n15072) );
  XNOR U19550 ( .A(n15065), .B(n15067), .Z(n15166) );
  NAND U19551 ( .A(n15167), .B(n15168), .Z(n15067) );
  OR U19552 ( .A(n15169), .B(n15170), .Z(n15168) );
  OR U19553 ( .A(n15171), .B(n15172), .Z(n15167) );
  NAND U19554 ( .A(n15173), .B(n15174), .Z(n15065) );
  OR U19555 ( .A(n15175), .B(n15176), .Z(n15174) );
  OR U19556 ( .A(n15177), .B(n15178), .Z(n15173) );
  ANDN U19557 ( .B(n15179), .A(n15180), .Z(n15066) );
  IV U19558 ( .A(n15181), .Z(n15179) );
  XNOR U19559 ( .A(n15146), .B(n15145), .Z(N28913) );
  XOR U19560 ( .A(n15165), .B(n15164), .Z(n15145) );
  XNOR U19561 ( .A(n15180), .B(n15181), .Z(n15164) );
  XNOR U19562 ( .A(n15175), .B(n15176), .Z(n15181) );
  XNOR U19563 ( .A(n15177), .B(n15178), .Z(n15176) );
  XNOR U19564 ( .A(y[1972]), .B(x[1972]), .Z(n15178) );
  XNOR U19565 ( .A(y[1973]), .B(x[1973]), .Z(n15177) );
  XNOR U19566 ( .A(y[1971]), .B(x[1971]), .Z(n15175) );
  XNOR U19567 ( .A(n15169), .B(n15170), .Z(n15180) );
  XNOR U19568 ( .A(y[1968]), .B(x[1968]), .Z(n15170) );
  XNOR U19569 ( .A(n15171), .B(n15172), .Z(n15169) );
  XNOR U19570 ( .A(y[1969]), .B(x[1969]), .Z(n15172) );
  XNOR U19571 ( .A(y[1970]), .B(x[1970]), .Z(n15171) );
  XNOR U19572 ( .A(n15162), .B(n15161), .Z(n15165) );
  XNOR U19573 ( .A(n15157), .B(n15158), .Z(n15161) );
  XNOR U19574 ( .A(y[1965]), .B(x[1965]), .Z(n15158) );
  XNOR U19575 ( .A(n15159), .B(n15160), .Z(n15157) );
  XNOR U19576 ( .A(y[1966]), .B(x[1966]), .Z(n15160) );
  XNOR U19577 ( .A(y[1967]), .B(x[1967]), .Z(n15159) );
  XNOR U19578 ( .A(n15151), .B(n15152), .Z(n15162) );
  XNOR U19579 ( .A(y[1962]), .B(x[1962]), .Z(n15152) );
  XNOR U19580 ( .A(n15153), .B(n15154), .Z(n15151) );
  XNOR U19581 ( .A(y[1963]), .B(x[1963]), .Z(n15154) );
  XNOR U19582 ( .A(y[1964]), .B(x[1964]), .Z(n15153) );
  XOR U19583 ( .A(n15127), .B(n15128), .Z(n15146) );
  XNOR U19584 ( .A(n15143), .B(n15144), .Z(n15128) );
  XNOR U19585 ( .A(n15138), .B(n15139), .Z(n15144) );
  XNOR U19586 ( .A(n15140), .B(n15141), .Z(n15139) );
  XNOR U19587 ( .A(y[1960]), .B(x[1960]), .Z(n15141) );
  XNOR U19588 ( .A(y[1961]), .B(x[1961]), .Z(n15140) );
  XNOR U19589 ( .A(y[1959]), .B(x[1959]), .Z(n15138) );
  XNOR U19590 ( .A(n15132), .B(n15133), .Z(n15143) );
  XNOR U19591 ( .A(y[1956]), .B(x[1956]), .Z(n15133) );
  XNOR U19592 ( .A(n15134), .B(n15135), .Z(n15132) );
  XNOR U19593 ( .A(y[1957]), .B(x[1957]), .Z(n15135) );
  XNOR U19594 ( .A(y[1958]), .B(x[1958]), .Z(n15134) );
  XOR U19595 ( .A(n15126), .B(n15125), .Z(n15127) );
  XNOR U19596 ( .A(n15121), .B(n15122), .Z(n15125) );
  XNOR U19597 ( .A(y[1953]), .B(x[1953]), .Z(n15122) );
  XNOR U19598 ( .A(n15123), .B(n15124), .Z(n15121) );
  XNOR U19599 ( .A(y[1954]), .B(x[1954]), .Z(n15124) );
  XNOR U19600 ( .A(y[1955]), .B(x[1955]), .Z(n15123) );
  XNOR U19601 ( .A(n15115), .B(n15116), .Z(n15126) );
  XNOR U19602 ( .A(y[1950]), .B(x[1950]), .Z(n15116) );
  XNOR U19603 ( .A(n15117), .B(n15118), .Z(n15115) );
  XNOR U19604 ( .A(y[1951]), .B(x[1951]), .Z(n15118) );
  XNOR U19605 ( .A(y[1952]), .B(x[1952]), .Z(n15117) );
  NAND U19606 ( .A(n15182), .B(n15183), .Z(N28905) );
  NANDN U19607 ( .A(n15184), .B(n15185), .Z(n15183) );
  OR U19608 ( .A(n15186), .B(n15187), .Z(n15185) );
  NAND U19609 ( .A(n15186), .B(n15187), .Z(n15182) );
  XOR U19610 ( .A(n15186), .B(n15188), .Z(N28904) );
  XNOR U19611 ( .A(n15184), .B(n15187), .Z(n15188) );
  AND U19612 ( .A(n15189), .B(n15190), .Z(n15187) );
  NANDN U19613 ( .A(n15191), .B(n15192), .Z(n15190) );
  NANDN U19614 ( .A(n15193), .B(n15194), .Z(n15192) );
  NANDN U19615 ( .A(n15194), .B(n15193), .Z(n15189) );
  NAND U19616 ( .A(n15195), .B(n15196), .Z(n15184) );
  NANDN U19617 ( .A(n15197), .B(n15198), .Z(n15196) );
  OR U19618 ( .A(n15199), .B(n15200), .Z(n15198) );
  NAND U19619 ( .A(n15200), .B(n15199), .Z(n15195) );
  AND U19620 ( .A(n15201), .B(n15202), .Z(n15186) );
  NANDN U19621 ( .A(n15203), .B(n15204), .Z(n15202) );
  NANDN U19622 ( .A(n15205), .B(n15206), .Z(n15204) );
  NANDN U19623 ( .A(n15206), .B(n15205), .Z(n15201) );
  XOR U19624 ( .A(n15200), .B(n15207), .Z(N28903) );
  XOR U19625 ( .A(n15197), .B(n15199), .Z(n15207) );
  XNOR U19626 ( .A(n15193), .B(n15208), .Z(n15199) );
  XNOR U19627 ( .A(n15191), .B(n15194), .Z(n15208) );
  NAND U19628 ( .A(n15209), .B(n15210), .Z(n15194) );
  NAND U19629 ( .A(n15211), .B(n15212), .Z(n15210) );
  OR U19630 ( .A(n15213), .B(n15214), .Z(n15211) );
  NANDN U19631 ( .A(n15215), .B(n15213), .Z(n15209) );
  IV U19632 ( .A(n15214), .Z(n15215) );
  NAND U19633 ( .A(n15216), .B(n15217), .Z(n15191) );
  NAND U19634 ( .A(n15218), .B(n15219), .Z(n15217) );
  NANDN U19635 ( .A(n15220), .B(n15221), .Z(n15218) );
  NANDN U19636 ( .A(n15221), .B(n15220), .Z(n15216) );
  AND U19637 ( .A(n15222), .B(n15223), .Z(n15193) );
  NAND U19638 ( .A(n15224), .B(n15225), .Z(n15223) );
  OR U19639 ( .A(n15226), .B(n15227), .Z(n15224) );
  NANDN U19640 ( .A(n15228), .B(n15226), .Z(n15222) );
  NAND U19641 ( .A(n15229), .B(n15230), .Z(n15197) );
  NANDN U19642 ( .A(n15231), .B(n15232), .Z(n15230) );
  OR U19643 ( .A(n15233), .B(n15234), .Z(n15232) );
  NANDN U19644 ( .A(n15235), .B(n15233), .Z(n15229) );
  IV U19645 ( .A(n15234), .Z(n15235) );
  XNOR U19646 ( .A(n15205), .B(n15236), .Z(n15200) );
  XNOR U19647 ( .A(n15203), .B(n15206), .Z(n15236) );
  NAND U19648 ( .A(n15237), .B(n15238), .Z(n15206) );
  NAND U19649 ( .A(n15239), .B(n15240), .Z(n15238) );
  OR U19650 ( .A(n15241), .B(n15242), .Z(n15239) );
  NANDN U19651 ( .A(n15243), .B(n15241), .Z(n15237) );
  IV U19652 ( .A(n15242), .Z(n15243) );
  NAND U19653 ( .A(n15244), .B(n15245), .Z(n15203) );
  NAND U19654 ( .A(n15246), .B(n15247), .Z(n15245) );
  NANDN U19655 ( .A(n15248), .B(n15249), .Z(n15246) );
  NANDN U19656 ( .A(n15249), .B(n15248), .Z(n15244) );
  AND U19657 ( .A(n15250), .B(n15251), .Z(n15205) );
  NAND U19658 ( .A(n15252), .B(n15253), .Z(n15251) );
  OR U19659 ( .A(n15254), .B(n15255), .Z(n15252) );
  NANDN U19660 ( .A(n15256), .B(n15254), .Z(n15250) );
  XNOR U19661 ( .A(n15231), .B(n15257), .Z(N28902) );
  XOR U19662 ( .A(n15233), .B(n15234), .Z(n15257) );
  XNOR U19663 ( .A(n15247), .B(n15258), .Z(n15234) );
  XOR U19664 ( .A(n15248), .B(n15249), .Z(n15258) );
  XOR U19665 ( .A(n15254), .B(n15259), .Z(n15249) );
  XOR U19666 ( .A(n15253), .B(n15256), .Z(n15259) );
  IV U19667 ( .A(n15255), .Z(n15256) );
  NAND U19668 ( .A(n15260), .B(n15261), .Z(n15255) );
  OR U19669 ( .A(n15262), .B(n15263), .Z(n15261) );
  OR U19670 ( .A(n15264), .B(n15265), .Z(n15260) );
  NAND U19671 ( .A(n15266), .B(n15267), .Z(n15253) );
  OR U19672 ( .A(n15268), .B(n15269), .Z(n15267) );
  OR U19673 ( .A(n15270), .B(n15271), .Z(n15266) );
  NOR U19674 ( .A(n15272), .B(n15273), .Z(n15254) );
  ANDN U19675 ( .B(n15274), .A(n15275), .Z(n15248) );
  XNOR U19676 ( .A(n15241), .B(n15276), .Z(n15247) );
  XNOR U19677 ( .A(n15240), .B(n15242), .Z(n15276) );
  NAND U19678 ( .A(n15277), .B(n15278), .Z(n15242) );
  OR U19679 ( .A(n15279), .B(n15280), .Z(n15278) );
  OR U19680 ( .A(n15281), .B(n15282), .Z(n15277) );
  NAND U19681 ( .A(n15283), .B(n15284), .Z(n15240) );
  OR U19682 ( .A(n15285), .B(n15286), .Z(n15284) );
  OR U19683 ( .A(n15287), .B(n15288), .Z(n15283) );
  ANDN U19684 ( .B(n15289), .A(n15290), .Z(n15241) );
  IV U19685 ( .A(n15291), .Z(n15289) );
  ANDN U19686 ( .B(n15292), .A(n15293), .Z(n15233) );
  XOR U19687 ( .A(n15219), .B(n15294), .Z(n15231) );
  XOR U19688 ( .A(n15220), .B(n15221), .Z(n15294) );
  XOR U19689 ( .A(n15226), .B(n15295), .Z(n15221) );
  XOR U19690 ( .A(n15225), .B(n15228), .Z(n15295) );
  IV U19691 ( .A(n15227), .Z(n15228) );
  NAND U19692 ( .A(n15296), .B(n15297), .Z(n15227) );
  OR U19693 ( .A(n15298), .B(n15299), .Z(n15297) );
  OR U19694 ( .A(n15300), .B(n15301), .Z(n15296) );
  NAND U19695 ( .A(n15302), .B(n15303), .Z(n15225) );
  OR U19696 ( .A(n15304), .B(n15305), .Z(n15303) );
  OR U19697 ( .A(n15306), .B(n15307), .Z(n15302) );
  NOR U19698 ( .A(n15308), .B(n15309), .Z(n15226) );
  ANDN U19699 ( .B(n15310), .A(n15311), .Z(n15220) );
  IV U19700 ( .A(n15312), .Z(n15310) );
  XNOR U19701 ( .A(n15213), .B(n15313), .Z(n15219) );
  XNOR U19702 ( .A(n15212), .B(n15214), .Z(n15313) );
  NAND U19703 ( .A(n15314), .B(n15315), .Z(n15214) );
  OR U19704 ( .A(n15316), .B(n15317), .Z(n15315) );
  OR U19705 ( .A(n15318), .B(n15319), .Z(n15314) );
  NAND U19706 ( .A(n15320), .B(n15321), .Z(n15212) );
  OR U19707 ( .A(n15322), .B(n15323), .Z(n15321) );
  OR U19708 ( .A(n15324), .B(n15325), .Z(n15320) );
  ANDN U19709 ( .B(n15326), .A(n15327), .Z(n15213) );
  IV U19710 ( .A(n15328), .Z(n15326) );
  XNOR U19711 ( .A(n15293), .B(n15292), .Z(N28901) );
  XOR U19712 ( .A(n15312), .B(n15311), .Z(n15292) );
  XNOR U19713 ( .A(n15327), .B(n15328), .Z(n15311) );
  XNOR U19714 ( .A(n15322), .B(n15323), .Z(n15328) );
  XNOR U19715 ( .A(n15324), .B(n15325), .Z(n15323) );
  XNOR U19716 ( .A(y[1948]), .B(x[1948]), .Z(n15325) );
  XNOR U19717 ( .A(y[1949]), .B(x[1949]), .Z(n15324) );
  XNOR U19718 ( .A(y[1947]), .B(x[1947]), .Z(n15322) );
  XNOR U19719 ( .A(n15316), .B(n15317), .Z(n15327) );
  XNOR U19720 ( .A(y[1944]), .B(x[1944]), .Z(n15317) );
  XNOR U19721 ( .A(n15318), .B(n15319), .Z(n15316) );
  XNOR U19722 ( .A(y[1945]), .B(x[1945]), .Z(n15319) );
  XNOR U19723 ( .A(y[1946]), .B(x[1946]), .Z(n15318) );
  XNOR U19724 ( .A(n15309), .B(n15308), .Z(n15312) );
  XNOR U19725 ( .A(n15304), .B(n15305), .Z(n15308) );
  XNOR U19726 ( .A(y[1941]), .B(x[1941]), .Z(n15305) );
  XNOR U19727 ( .A(n15306), .B(n15307), .Z(n15304) );
  XNOR U19728 ( .A(y[1942]), .B(x[1942]), .Z(n15307) );
  XNOR U19729 ( .A(y[1943]), .B(x[1943]), .Z(n15306) );
  XNOR U19730 ( .A(n15298), .B(n15299), .Z(n15309) );
  XNOR U19731 ( .A(y[1938]), .B(x[1938]), .Z(n15299) );
  XNOR U19732 ( .A(n15300), .B(n15301), .Z(n15298) );
  XNOR U19733 ( .A(y[1939]), .B(x[1939]), .Z(n15301) );
  XNOR U19734 ( .A(y[1940]), .B(x[1940]), .Z(n15300) );
  XOR U19735 ( .A(n15274), .B(n15275), .Z(n15293) );
  XNOR U19736 ( .A(n15290), .B(n15291), .Z(n15275) );
  XNOR U19737 ( .A(n15285), .B(n15286), .Z(n15291) );
  XNOR U19738 ( .A(n15287), .B(n15288), .Z(n15286) );
  XNOR U19739 ( .A(y[1936]), .B(x[1936]), .Z(n15288) );
  XNOR U19740 ( .A(y[1937]), .B(x[1937]), .Z(n15287) );
  XNOR U19741 ( .A(y[1935]), .B(x[1935]), .Z(n15285) );
  XNOR U19742 ( .A(n15279), .B(n15280), .Z(n15290) );
  XNOR U19743 ( .A(y[1932]), .B(x[1932]), .Z(n15280) );
  XNOR U19744 ( .A(n15281), .B(n15282), .Z(n15279) );
  XNOR U19745 ( .A(y[1933]), .B(x[1933]), .Z(n15282) );
  XNOR U19746 ( .A(y[1934]), .B(x[1934]), .Z(n15281) );
  XOR U19747 ( .A(n15273), .B(n15272), .Z(n15274) );
  XNOR U19748 ( .A(n15268), .B(n15269), .Z(n15272) );
  XNOR U19749 ( .A(y[1929]), .B(x[1929]), .Z(n15269) );
  XNOR U19750 ( .A(n15270), .B(n15271), .Z(n15268) );
  XNOR U19751 ( .A(y[1930]), .B(x[1930]), .Z(n15271) );
  XNOR U19752 ( .A(y[1931]), .B(x[1931]), .Z(n15270) );
  XNOR U19753 ( .A(n15262), .B(n15263), .Z(n15273) );
  XNOR U19754 ( .A(y[1926]), .B(x[1926]), .Z(n15263) );
  XNOR U19755 ( .A(n15264), .B(n15265), .Z(n15262) );
  XNOR U19756 ( .A(y[1927]), .B(x[1927]), .Z(n15265) );
  XNOR U19757 ( .A(y[1928]), .B(x[1928]), .Z(n15264) );
  NAND U19758 ( .A(n15329), .B(n15330), .Z(N28893) );
  NANDN U19759 ( .A(n15331), .B(n15332), .Z(n15330) );
  OR U19760 ( .A(n15333), .B(n15334), .Z(n15332) );
  NAND U19761 ( .A(n15333), .B(n15334), .Z(n15329) );
  XOR U19762 ( .A(n15333), .B(n15335), .Z(N28892) );
  XNOR U19763 ( .A(n15331), .B(n15334), .Z(n15335) );
  AND U19764 ( .A(n15336), .B(n15337), .Z(n15334) );
  NANDN U19765 ( .A(n15338), .B(n15339), .Z(n15337) );
  NANDN U19766 ( .A(n15340), .B(n15341), .Z(n15339) );
  NANDN U19767 ( .A(n15341), .B(n15340), .Z(n15336) );
  NAND U19768 ( .A(n15342), .B(n15343), .Z(n15331) );
  NANDN U19769 ( .A(n15344), .B(n15345), .Z(n15343) );
  OR U19770 ( .A(n15346), .B(n15347), .Z(n15345) );
  NAND U19771 ( .A(n15347), .B(n15346), .Z(n15342) );
  AND U19772 ( .A(n15348), .B(n15349), .Z(n15333) );
  NANDN U19773 ( .A(n15350), .B(n15351), .Z(n15349) );
  NANDN U19774 ( .A(n15352), .B(n15353), .Z(n15351) );
  NANDN U19775 ( .A(n15353), .B(n15352), .Z(n15348) );
  XOR U19776 ( .A(n15347), .B(n15354), .Z(N28891) );
  XOR U19777 ( .A(n15344), .B(n15346), .Z(n15354) );
  XNOR U19778 ( .A(n15340), .B(n15355), .Z(n15346) );
  XNOR U19779 ( .A(n15338), .B(n15341), .Z(n15355) );
  NAND U19780 ( .A(n15356), .B(n15357), .Z(n15341) );
  NAND U19781 ( .A(n15358), .B(n15359), .Z(n15357) );
  OR U19782 ( .A(n15360), .B(n15361), .Z(n15358) );
  NANDN U19783 ( .A(n15362), .B(n15360), .Z(n15356) );
  IV U19784 ( .A(n15361), .Z(n15362) );
  NAND U19785 ( .A(n15363), .B(n15364), .Z(n15338) );
  NAND U19786 ( .A(n15365), .B(n15366), .Z(n15364) );
  NANDN U19787 ( .A(n15367), .B(n15368), .Z(n15365) );
  NANDN U19788 ( .A(n15368), .B(n15367), .Z(n15363) );
  AND U19789 ( .A(n15369), .B(n15370), .Z(n15340) );
  NAND U19790 ( .A(n15371), .B(n15372), .Z(n15370) );
  OR U19791 ( .A(n15373), .B(n15374), .Z(n15371) );
  NANDN U19792 ( .A(n15375), .B(n15373), .Z(n15369) );
  NAND U19793 ( .A(n15376), .B(n15377), .Z(n15344) );
  NANDN U19794 ( .A(n15378), .B(n15379), .Z(n15377) );
  OR U19795 ( .A(n15380), .B(n15381), .Z(n15379) );
  NANDN U19796 ( .A(n15382), .B(n15380), .Z(n15376) );
  IV U19797 ( .A(n15381), .Z(n15382) );
  XNOR U19798 ( .A(n15352), .B(n15383), .Z(n15347) );
  XNOR U19799 ( .A(n15350), .B(n15353), .Z(n15383) );
  NAND U19800 ( .A(n15384), .B(n15385), .Z(n15353) );
  NAND U19801 ( .A(n15386), .B(n15387), .Z(n15385) );
  OR U19802 ( .A(n15388), .B(n15389), .Z(n15386) );
  NANDN U19803 ( .A(n15390), .B(n15388), .Z(n15384) );
  IV U19804 ( .A(n15389), .Z(n15390) );
  NAND U19805 ( .A(n15391), .B(n15392), .Z(n15350) );
  NAND U19806 ( .A(n15393), .B(n15394), .Z(n15392) );
  NANDN U19807 ( .A(n15395), .B(n15396), .Z(n15393) );
  NANDN U19808 ( .A(n15396), .B(n15395), .Z(n15391) );
  AND U19809 ( .A(n15397), .B(n15398), .Z(n15352) );
  NAND U19810 ( .A(n15399), .B(n15400), .Z(n15398) );
  OR U19811 ( .A(n15401), .B(n15402), .Z(n15399) );
  NANDN U19812 ( .A(n15403), .B(n15401), .Z(n15397) );
  XNOR U19813 ( .A(n15378), .B(n15404), .Z(N28890) );
  XOR U19814 ( .A(n15380), .B(n15381), .Z(n15404) );
  XNOR U19815 ( .A(n15394), .B(n15405), .Z(n15381) );
  XOR U19816 ( .A(n15395), .B(n15396), .Z(n15405) );
  XOR U19817 ( .A(n15401), .B(n15406), .Z(n15396) );
  XOR U19818 ( .A(n15400), .B(n15403), .Z(n15406) );
  IV U19819 ( .A(n15402), .Z(n15403) );
  NAND U19820 ( .A(n15407), .B(n15408), .Z(n15402) );
  OR U19821 ( .A(n15409), .B(n15410), .Z(n15408) );
  OR U19822 ( .A(n15411), .B(n15412), .Z(n15407) );
  NAND U19823 ( .A(n15413), .B(n15414), .Z(n15400) );
  OR U19824 ( .A(n15415), .B(n15416), .Z(n15414) );
  OR U19825 ( .A(n15417), .B(n15418), .Z(n15413) );
  NOR U19826 ( .A(n15419), .B(n15420), .Z(n15401) );
  ANDN U19827 ( .B(n15421), .A(n15422), .Z(n15395) );
  XNOR U19828 ( .A(n15388), .B(n15423), .Z(n15394) );
  XNOR U19829 ( .A(n15387), .B(n15389), .Z(n15423) );
  NAND U19830 ( .A(n15424), .B(n15425), .Z(n15389) );
  OR U19831 ( .A(n15426), .B(n15427), .Z(n15425) );
  OR U19832 ( .A(n15428), .B(n15429), .Z(n15424) );
  NAND U19833 ( .A(n15430), .B(n15431), .Z(n15387) );
  OR U19834 ( .A(n15432), .B(n15433), .Z(n15431) );
  OR U19835 ( .A(n15434), .B(n15435), .Z(n15430) );
  ANDN U19836 ( .B(n15436), .A(n15437), .Z(n15388) );
  IV U19837 ( .A(n15438), .Z(n15436) );
  ANDN U19838 ( .B(n15439), .A(n15440), .Z(n15380) );
  XOR U19839 ( .A(n15366), .B(n15441), .Z(n15378) );
  XOR U19840 ( .A(n15367), .B(n15368), .Z(n15441) );
  XOR U19841 ( .A(n15373), .B(n15442), .Z(n15368) );
  XOR U19842 ( .A(n15372), .B(n15375), .Z(n15442) );
  IV U19843 ( .A(n15374), .Z(n15375) );
  NAND U19844 ( .A(n15443), .B(n15444), .Z(n15374) );
  OR U19845 ( .A(n15445), .B(n15446), .Z(n15444) );
  OR U19846 ( .A(n15447), .B(n15448), .Z(n15443) );
  NAND U19847 ( .A(n15449), .B(n15450), .Z(n15372) );
  OR U19848 ( .A(n15451), .B(n15452), .Z(n15450) );
  OR U19849 ( .A(n15453), .B(n15454), .Z(n15449) );
  NOR U19850 ( .A(n15455), .B(n15456), .Z(n15373) );
  ANDN U19851 ( .B(n15457), .A(n15458), .Z(n15367) );
  IV U19852 ( .A(n15459), .Z(n15457) );
  XNOR U19853 ( .A(n15360), .B(n15460), .Z(n15366) );
  XNOR U19854 ( .A(n15359), .B(n15361), .Z(n15460) );
  NAND U19855 ( .A(n15461), .B(n15462), .Z(n15361) );
  OR U19856 ( .A(n15463), .B(n15464), .Z(n15462) );
  OR U19857 ( .A(n15465), .B(n15466), .Z(n15461) );
  NAND U19858 ( .A(n15467), .B(n15468), .Z(n15359) );
  OR U19859 ( .A(n15469), .B(n15470), .Z(n15468) );
  OR U19860 ( .A(n15471), .B(n15472), .Z(n15467) );
  ANDN U19861 ( .B(n15473), .A(n15474), .Z(n15360) );
  IV U19862 ( .A(n15475), .Z(n15473) );
  XNOR U19863 ( .A(n15440), .B(n15439), .Z(N28889) );
  XOR U19864 ( .A(n15459), .B(n15458), .Z(n15439) );
  XNOR U19865 ( .A(n15474), .B(n15475), .Z(n15458) );
  XNOR U19866 ( .A(n15469), .B(n15470), .Z(n15475) );
  XNOR U19867 ( .A(n15471), .B(n15472), .Z(n15470) );
  XNOR U19868 ( .A(y[1924]), .B(x[1924]), .Z(n15472) );
  XNOR U19869 ( .A(y[1925]), .B(x[1925]), .Z(n15471) );
  XNOR U19870 ( .A(y[1923]), .B(x[1923]), .Z(n15469) );
  XNOR U19871 ( .A(n15463), .B(n15464), .Z(n15474) );
  XNOR U19872 ( .A(y[1920]), .B(x[1920]), .Z(n15464) );
  XNOR U19873 ( .A(n15465), .B(n15466), .Z(n15463) );
  XNOR U19874 ( .A(y[1921]), .B(x[1921]), .Z(n15466) );
  XNOR U19875 ( .A(y[1922]), .B(x[1922]), .Z(n15465) );
  XNOR U19876 ( .A(n15456), .B(n15455), .Z(n15459) );
  XNOR U19877 ( .A(n15451), .B(n15452), .Z(n15455) );
  XNOR U19878 ( .A(y[1917]), .B(x[1917]), .Z(n15452) );
  XNOR U19879 ( .A(n15453), .B(n15454), .Z(n15451) );
  XNOR U19880 ( .A(y[1918]), .B(x[1918]), .Z(n15454) );
  XNOR U19881 ( .A(y[1919]), .B(x[1919]), .Z(n15453) );
  XNOR U19882 ( .A(n15445), .B(n15446), .Z(n15456) );
  XNOR U19883 ( .A(y[1914]), .B(x[1914]), .Z(n15446) );
  XNOR U19884 ( .A(n15447), .B(n15448), .Z(n15445) );
  XNOR U19885 ( .A(y[1915]), .B(x[1915]), .Z(n15448) );
  XNOR U19886 ( .A(y[1916]), .B(x[1916]), .Z(n15447) );
  XOR U19887 ( .A(n15421), .B(n15422), .Z(n15440) );
  XNOR U19888 ( .A(n15437), .B(n15438), .Z(n15422) );
  XNOR U19889 ( .A(n15432), .B(n15433), .Z(n15438) );
  XNOR U19890 ( .A(n15434), .B(n15435), .Z(n15433) );
  XNOR U19891 ( .A(y[1912]), .B(x[1912]), .Z(n15435) );
  XNOR U19892 ( .A(y[1913]), .B(x[1913]), .Z(n15434) );
  XNOR U19893 ( .A(y[1911]), .B(x[1911]), .Z(n15432) );
  XNOR U19894 ( .A(n15426), .B(n15427), .Z(n15437) );
  XNOR U19895 ( .A(y[1908]), .B(x[1908]), .Z(n15427) );
  XNOR U19896 ( .A(n15428), .B(n15429), .Z(n15426) );
  XNOR U19897 ( .A(y[1909]), .B(x[1909]), .Z(n15429) );
  XNOR U19898 ( .A(y[1910]), .B(x[1910]), .Z(n15428) );
  XOR U19899 ( .A(n15420), .B(n15419), .Z(n15421) );
  XNOR U19900 ( .A(n15415), .B(n15416), .Z(n15419) );
  XNOR U19901 ( .A(y[1905]), .B(x[1905]), .Z(n15416) );
  XNOR U19902 ( .A(n15417), .B(n15418), .Z(n15415) );
  XNOR U19903 ( .A(y[1906]), .B(x[1906]), .Z(n15418) );
  XNOR U19904 ( .A(y[1907]), .B(x[1907]), .Z(n15417) );
  XNOR U19905 ( .A(n15409), .B(n15410), .Z(n15420) );
  XNOR U19906 ( .A(y[1902]), .B(x[1902]), .Z(n15410) );
  XNOR U19907 ( .A(n15411), .B(n15412), .Z(n15409) );
  XNOR U19908 ( .A(y[1903]), .B(x[1903]), .Z(n15412) );
  XNOR U19909 ( .A(y[1904]), .B(x[1904]), .Z(n15411) );
  NAND U19910 ( .A(n15476), .B(n15477), .Z(N28881) );
  NANDN U19911 ( .A(n15478), .B(n15479), .Z(n15477) );
  OR U19912 ( .A(n15480), .B(n15481), .Z(n15479) );
  NAND U19913 ( .A(n15480), .B(n15481), .Z(n15476) );
  XOR U19914 ( .A(n15480), .B(n15482), .Z(N28880) );
  XNOR U19915 ( .A(n15478), .B(n15481), .Z(n15482) );
  AND U19916 ( .A(n15483), .B(n15484), .Z(n15481) );
  NANDN U19917 ( .A(n15485), .B(n15486), .Z(n15484) );
  NANDN U19918 ( .A(n15487), .B(n15488), .Z(n15486) );
  NANDN U19919 ( .A(n15488), .B(n15487), .Z(n15483) );
  NAND U19920 ( .A(n15489), .B(n15490), .Z(n15478) );
  NANDN U19921 ( .A(n15491), .B(n15492), .Z(n15490) );
  OR U19922 ( .A(n15493), .B(n15494), .Z(n15492) );
  NAND U19923 ( .A(n15494), .B(n15493), .Z(n15489) );
  AND U19924 ( .A(n15495), .B(n15496), .Z(n15480) );
  NANDN U19925 ( .A(n15497), .B(n15498), .Z(n15496) );
  NANDN U19926 ( .A(n15499), .B(n15500), .Z(n15498) );
  NANDN U19927 ( .A(n15500), .B(n15499), .Z(n15495) );
  XOR U19928 ( .A(n15494), .B(n15501), .Z(N28879) );
  XOR U19929 ( .A(n15491), .B(n15493), .Z(n15501) );
  XNOR U19930 ( .A(n15487), .B(n15502), .Z(n15493) );
  XNOR U19931 ( .A(n15485), .B(n15488), .Z(n15502) );
  NAND U19932 ( .A(n15503), .B(n15504), .Z(n15488) );
  NAND U19933 ( .A(n15505), .B(n15506), .Z(n15504) );
  OR U19934 ( .A(n15507), .B(n15508), .Z(n15505) );
  NANDN U19935 ( .A(n15509), .B(n15507), .Z(n15503) );
  IV U19936 ( .A(n15508), .Z(n15509) );
  NAND U19937 ( .A(n15510), .B(n15511), .Z(n15485) );
  NAND U19938 ( .A(n15512), .B(n15513), .Z(n15511) );
  NANDN U19939 ( .A(n15514), .B(n15515), .Z(n15512) );
  NANDN U19940 ( .A(n15515), .B(n15514), .Z(n15510) );
  AND U19941 ( .A(n15516), .B(n15517), .Z(n15487) );
  NAND U19942 ( .A(n15518), .B(n15519), .Z(n15517) );
  OR U19943 ( .A(n15520), .B(n15521), .Z(n15518) );
  NANDN U19944 ( .A(n15522), .B(n15520), .Z(n15516) );
  NAND U19945 ( .A(n15523), .B(n15524), .Z(n15491) );
  NANDN U19946 ( .A(n15525), .B(n15526), .Z(n15524) );
  OR U19947 ( .A(n15527), .B(n15528), .Z(n15526) );
  NANDN U19948 ( .A(n15529), .B(n15527), .Z(n15523) );
  IV U19949 ( .A(n15528), .Z(n15529) );
  XNOR U19950 ( .A(n15499), .B(n15530), .Z(n15494) );
  XNOR U19951 ( .A(n15497), .B(n15500), .Z(n15530) );
  NAND U19952 ( .A(n15531), .B(n15532), .Z(n15500) );
  NAND U19953 ( .A(n15533), .B(n15534), .Z(n15532) );
  OR U19954 ( .A(n15535), .B(n15536), .Z(n15533) );
  NANDN U19955 ( .A(n15537), .B(n15535), .Z(n15531) );
  IV U19956 ( .A(n15536), .Z(n15537) );
  NAND U19957 ( .A(n15538), .B(n15539), .Z(n15497) );
  NAND U19958 ( .A(n15540), .B(n15541), .Z(n15539) );
  NANDN U19959 ( .A(n15542), .B(n15543), .Z(n15540) );
  NANDN U19960 ( .A(n15543), .B(n15542), .Z(n15538) );
  AND U19961 ( .A(n15544), .B(n15545), .Z(n15499) );
  NAND U19962 ( .A(n15546), .B(n15547), .Z(n15545) );
  OR U19963 ( .A(n15548), .B(n15549), .Z(n15546) );
  NANDN U19964 ( .A(n15550), .B(n15548), .Z(n15544) );
  XNOR U19965 ( .A(n15525), .B(n15551), .Z(N28878) );
  XOR U19966 ( .A(n15527), .B(n15528), .Z(n15551) );
  XNOR U19967 ( .A(n15541), .B(n15552), .Z(n15528) );
  XOR U19968 ( .A(n15542), .B(n15543), .Z(n15552) );
  XOR U19969 ( .A(n15548), .B(n15553), .Z(n15543) );
  XOR U19970 ( .A(n15547), .B(n15550), .Z(n15553) );
  IV U19971 ( .A(n15549), .Z(n15550) );
  NAND U19972 ( .A(n15554), .B(n15555), .Z(n15549) );
  OR U19973 ( .A(n15556), .B(n15557), .Z(n15555) );
  OR U19974 ( .A(n15558), .B(n15559), .Z(n15554) );
  NAND U19975 ( .A(n15560), .B(n15561), .Z(n15547) );
  OR U19976 ( .A(n15562), .B(n15563), .Z(n15561) );
  OR U19977 ( .A(n15564), .B(n15565), .Z(n15560) );
  NOR U19978 ( .A(n15566), .B(n15567), .Z(n15548) );
  ANDN U19979 ( .B(n15568), .A(n15569), .Z(n15542) );
  XNOR U19980 ( .A(n15535), .B(n15570), .Z(n15541) );
  XNOR U19981 ( .A(n15534), .B(n15536), .Z(n15570) );
  NAND U19982 ( .A(n15571), .B(n15572), .Z(n15536) );
  OR U19983 ( .A(n15573), .B(n15574), .Z(n15572) );
  OR U19984 ( .A(n15575), .B(n15576), .Z(n15571) );
  NAND U19985 ( .A(n15577), .B(n15578), .Z(n15534) );
  OR U19986 ( .A(n15579), .B(n15580), .Z(n15578) );
  OR U19987 ( .A(n15581), .B(n15582), .Z(n15577) );
  ANDN U19988 ( .B(n15583), .A(n15584), .Z(n15535) );
  IV U19989 ( .A(n15585), .Z(n15583) );
  ANDN U19990 ( .B(n15586), .A(n15587), .Z(n15527) );
  XOR U19991 ( .A(n15513), .B(n15588), .Z(n15525) );
  XOR U19992 ( .A(n15514), .B(n15515), .Z(n15588) );
  XOR U19993 ( .A(n15520), .B(n15589), .Z(n15515) );
  XOR U19994 ( .A(n15519), .B(n15522), .Z(n15589) );
  IV U19995 ( .A(n15521), .Z(n15522) );
  NAND U19996 ( .A(n15590), .B(n15591), .Z(n15521) );
  OR U19997 ( .A(n15592), .B(n15593), .Z(n15591) );
  OR U19998 ( .A(n15594), .B(n15595), .Z(n15590) );
  NAND U19999 ( .A(n15596), .B(n15597), .Z(n15519) );
  OR U20000 ( .A(n15598), .B(n15599), .Z(n15597) );
  OR U20001 ( .A(n15600), .B(n15601), .Z(n15596) );
  NOR U20002 ( .A(n15602), .B(n15603), .Z(n15520) );
  ANDN U20003 ( .B(n15604), .A(n15605), .Z(n15514) );
  IV U20004 ( .A(n15606), .Z(n15604) );
  XNOR U20005 ( .A(n15507), .B(n15607), .Z(n15513) );
  XNOR U20006 ( .A(n15506), .B(n15508), .Z(n15607) );
  NAND U20007 ( .A(n15608), .B(n15609), .Z(n15508) );
  OR U20008 ( .A(n15610), .B(n15611), .Z(n15609) );
  OR U20009 ( .A(n15612), .B(n15613), .Z(n15608) );
  NAND U20010 ( .A(n15614), .B(n15615), .Z(n15506) );
  OR U20011 ( .A(n15616), .B(n15617), .Z(n15615) );
  OR U20012 ( .A(n15618), .B(n15619), .Z(n15614) );
  ANDN U20013 ( .B(n15620), .A(n15621), .Z(n15507) );
  IV U20014 ( .A(n15622), .Z(n15620) );
  XNOR U20015 ( .A(n15587), .B(n15586), .Z(N28877) );
  XOR U20016 ( .A(n15606), .B(n15605), .Z(n15586) );
  XNOR U20017 ( .A(n15621), .B(n15622), .Z(n15605) );
  XNOR U20018 ( .A(n15616), .B(n15617), .Z(n15622) );
  XNOR U20019 ( .A(n15618), .B(n15619), .Z(n15617) );
  XNOR U20020 ( .A(y[1900]), .B(x[1900]), .Z(n15619) );
  XNOR U20021 ( .A(y[1901]), .B(x[1901]), .Z(n15618) );
  XNOR U20022 ( .A(y[1899]), .B(x[1899]), .Z(n15616) );
  XNOR U20023 ( .A(n15610), .B(n15611), .Z(n15621) );
  XNOR U20024 ( .A(y[1896]), .B(x[1896]), .Z(n15611) );
  XNOR U20025 ( .A(n15612), .B(n15613), .Z(n15610) );
  XNOR U20026 ( .A(y[1897]), .B(x[1897]), .Z(n15613) );
  XNOR U20027 ( .A(y[1898]), .B(x[1898]), .Z(n15612) );
  XNOR U20028 ( .A(n15603), .B(n15602), .Z(n15606) );
  XNOR U20029 ( .A(n15598), .B(n15599), .Z(n15602) );
  XNOR U20030 ( .A(y[1893]), .B(x[1893]), .Z(n15599) );
  XNOR U20031 ( .A(n15600), .B(n15601), .Z(n15598) );
  XNOR U20032 ( .A(y[1894]), .B(x[1894]), .Z(n15601) );
  XNOR U20033 ( .A(y[1895]), .B(x[1895]), .Z(n15600) );
  XNOR U20034 ( .A(n15592), .B(n15593), .Z(n15603) );
  XNOR U20035 ( .A(y[1890]), .B(x[1890]), .Z(n15593) );
  XNOR U20036 ( .A(n15594), .B(n15595), .Z(n15592) );
  XNOR U20037 ( .A(y[1891]), .B(x[1891]), .Z(n15595) );
  XNOR U20038 ( .A(y[1892]), .B(x[1892]), .Z(n15594) );
  XOR U20039 ( .A(n15568), .B(n15569), .Z(n15587) );
  XNOR U20040 ( .A(n15584), .B(n15585), .Z(n15569) );
  XNOR U20041 ( .A(n15579), .B(n15580), .Z(n15585) );
  XNOR U20042 ( .A(n15581), .B(n15582), .Z(n15580) );
  XNOR U20043 ( .A(y[1888]), .B(x[1888]), .Z(n15582) );
  XNOR U20044 ( .A(y[1889]), .B(x[1889]), .Z(n15581) );
  XNOR U20045 ( .A(y[1887]), .B(x[1887]), .Z(n15579) );
  XNOR U20046 ( .A(n15573), .B(n15574), .Z(n15584) );
  XNOR U20047 ( .A(y[1884]), .B(x[1884]), .Z(n15574) );
  XNOR U20048 ( .A(n15575), .B(n15576), .Z(n15573) );
  XNOR U20049 ( .A(y[1885]), .B(x[1885]), .Z(n15576) );
  XNOR U20050 ( .A(y[1886]), .B(x[1886]), .Z(n15575) );
  XOR U20051 ( .A(n15567), .B(n15566), .Z(n15568) );
  XNOR U20052 ( .A(n15562), .B(n15563), .Z(n15566) );
  XNOR U20053 ( .A(y[1881]), .B(x[1881]), .Z(n15563) );
  XNOR U20054 ( .A(n15564), .B(n15565), .Z(n15562) );
  XNOR U20055 ( .A(y[1882]), .B(x[1882]), .Z(n15565) );
  XNOR U20056 ( .A(y[1883]), .B(x[1883]), .Z(n15564) );
  XNOR U20057 ( .A(n15556), .B(n15557), .Z(n15567) );
  XNOR U20058 ( .A(y[1878]), .B(x[1878]), .Z(n15557) );
  XNOR U20059 ( .A(n15558), .B(n15559), .Z(n15556) );
  XNOR U20060 ( .A(y[1879]), .B(x[1879]), .Z(n15559) );
  XNOR U20061 ( .A(y[1880]), .B(x[1880]), .Z(n15558) );
  NAND U20062 ( .A(n15623), .B(n15624), .Z(N28869) );
  NANDN U20063 ( .A(n15625), .B(n15626), .Z(n15624) );
  OR U20064 ( .A(n15627), .B(n15628), .Z(n15626) );
  NAND U20065 ( .A(n15627), .B(n15628), .Z(n15623) );
  XOR U20066 ( .A(n15627), .B(n15629), .Z(N28868) );
  XNOR U20067 ( .A(n15625), .B(n15628), .Z(n15629) );
  AND U20068 ( .A(n15630), .B(n15631), .Z(n15628) );
  NANDN U20069 ( .A(n15632), .B(n15633), .Z(n15631) );
  NANDN U20070 ( .A(n15634), .B(n15635), .Z(n15633) );
  NANDN U20071 ( .A(n15635), .B(n15634), .Z(n15630) );
  NAND U20072 ( .A(n15636), .B(n15637), .Z(n15625) );
  NANDN U20073 ( .A(n15638), .B(n15639), .Z(n15637) );
  OR U20074 ( .A(n15640), .B(n15641), .Z(n15639) );
  NAND U20075 ( .A(n15641), .B(n15640), .Z(n15636) );
  AND U20076 ( .A(n15642), .B(n15643), .Z(n15627) );
  NANDN U20077 ( .A(n15644), .B(n15645), .Z(n15643) );
  NANDN U20078 ( .A(n15646), .B(n15647), .Z(n15645) );
  NANDN U20079 ( .A(n15647), .B(n15646), .Z(n15642) );
  XOR U20080 ( .A(n15641), .B(n15648), .Z(N28867) );
  XOR U20081 ( .A(n15638), .B(n15640), .Z(n15648) );
  XNOR U20082 ( .A(n15634), .B(n15649), .Z(n15640) );
  XNOR U20083 ( .A(n15632), .B(n15635), .Z(n15649) );
  NAND U20084 ( .A(n15650), .B(n15651), .Z(n15635) );
  NAND U20085 ( .A(n15652), .B(n15653), .Z(n15651) );
  OR U20086 ( .A(n15654), .B(n15655), .Z(n15652) );
  NANDN U20087 ( .A(n15656), .B(n15654), .Z(n15650) );
  IV U20088 ( .A(n15655), .Z(n15656) );
  NAND U20089 ( .A(n15657), .B(n15658), .Z(n15632) );
  NAND U20090 ( .A(n15659), .B(n15660), .Z(n15658) );
  NANDN U20091 ( .A(n15661), .B(n15662), .Z(n15659) );
  NANDN U20092 ( .A(n15662), .B(n15661), .Z(n15657) );
  AND U20093 ( .A(n15663), .B(n15664), .Z(n15634) );
  NAND U20094 ( .A(n15665), .B(n15666), .Z(n15664) );
  OR U20095 ( .A(n15667), .B(n15668), .Z(n15665) );
  NANDN U20096 ( .A(n15669), .B(n15667), .Z(n15663) );
  NAND U20097 ( .A(n15670), .B(n15671), .Z(n15638) );
  NANDN U20098 ( .A(n15672), .B(n15673), .Z(n15671) );
  OR U20099 ( .A(n15674), .B(n15675), .Z(n15673) );
  NANDN U20100 ( .A(n15676), .B(n15674), .Z(n15670) );
  IV U20101 ( .A(n15675), .Z(n15676) );
  XNOR U20102 ( .A(n15646), .B(n15677), .Z(n15641) );
  XNOR U20103 ( .A(n15644), .B(n15647), .Z(n15677) );
  NAND U20104 ( .A(n15678), .B(n15679), .Z(n15647) );
  NAND U20105 ( .A(n15680), .B(n15681), .Z(n15679) );
  OR U20106 ( .A(n15682), .B(n15683), .Z(n15680) );
  NANDN U20107 ( .A(n15684), .B(n15682), .Z(n15678) );
  IV U20108 ( .A(n15683), .Z(n15684) );
  NAND U20109 ( .A(n15685), .B(n15686), .Z(n15644) );
  NAND U20110 ( .A(n15687), .B(n15688), .Z(n15686) );
  NANDN U20111 ( .A(n15689), .B(n15690), .Z(n15687) );
  NANDN U20112 ( .A(n15690), .B(n15689), .Z(n15685) );
  AND U20113 ( .A(n15691), .B(n15692), .Z(n15646) );
  NAND U20114 ( .A(n15693), .B(n15694), .Z(n15692) );
  OR U20115 ( .A(n15695), .B(n15696), .Z(n15693) );
  NANDN U20116 ( .A(n15697), .B(n15695), .Z(n15691) );
  XNOR U20117 ( .A(n15672), .B(n15698), .Z(N28866) );
  XOR U20118 ( .A(n15674), .B(n15675), .Z(n15698) );
  XNOR U20119 ( .A(n15688), .B(n15699), .Z(n15675) );
  XOR U20120 ( .A(n15689), .B(n15690), .Z(n15699) );
  XOR U20121 ( .A(n15695), .B(n15700), .Z(n15690) );
  XOR U20122 ( .A(n15694), .B(n15697), .Z(n15700) );
  IV U20123 ( .A(n15696), .Z(n15697) );
  NAND U20124 ( .A(n15701), .B(n15702), .Z(n15696) );
  OR U20125 ( .A(n15703), .B(n15704), .Z(n15702) );
  OR U20126 ( .A(n15705), .B(n15706), .Z(n15701) );
  NAND U20127 ( .A(n15707), .B(n15708), .Z(n15694) );
  OR U20128 ( .A(n15709), .B(n15710), .Z(n15708) );
  OR U20129 ( .A(n15711), .B(n15712), .Z(n15707) );
  NOR U20130 ( .A(n15713), .B(n15714), .Z(n15695) );
  ANDN U20131 ( .B(n15715), .A(n15716), .Z(n15689) );
  XNOR U20132 ( .A(n15682), .B(n15717), .Z(n15688) );
  XNOR U20133 ( .A(n15681), .B(n15683), .Z(n15717) );
  NAND U20134 ( .A(n15718), .B(n15719), .Z(n15683) );
  OR U20135 ( .A(n15720), .B(n15721), .Z(n15719) );
  OR U20136 ( .A(n15722), .B(n15723), .Z(n15718) );
  NAND U20137 ( .A(n15724), .B(n15725), .Z(n15681) );
  OR U20138 ( .A(n15726), .B(n15727), .Z(n15725) );
  OR U20139 ( .A(n15728), .B(n15729), .Z(n15724) );
  ANDN U20140 ( .B(n15730), .A(n15731), .Z(n15682) );
  IV U20141 ( .A(n15732), .Z(n15730) );
  ANDN U20142 ( .B(n15733), .A(n15734), .Z(n15674) );
  XOR U20143 ( .A(n15660), .B(n15735), .Z(n15672) );
  XOR U20144 ( .A(n15661), .B(n15662), .Z(n15735) );
  XOR U20145 ( .A(n15667), .B(n15736), .Z(n15662) );
  XOR U20146 ( .A(n15666), .B(n15669), .Z(n15736) );
  IV U20147 ( .A(n15668), .Z(n15669) );
  NAND U20148 ( .A(n15737), .B(n15738), .Z(n15668) );
  OR U20149 ( .A(n15739), .B(n15740), .Z(n15738) );
  OR U20150 ( .A(n15741), .B(n15742), .Z(n15737) );
  NAND U20151 ( .A(n15743), .B(n15744), .Z(n15666) );
  OR U20152 ( .A(n15745), .B(n15746), .Z(n15744) );
  OR U20153 ( .A(n15747), .B(n15748), .Z(n15743) );
  NOR U20154 ( .A(n15749), .B(n15750), .Z(n15667) );
  ANDN U20155 ( .B(n15751), .A(n15752), .Z(n15661) );
  IV U20156 ( .A(n15753), .Z(n15751) );
  XNOR U20157 ( .A(n15654), .B(n15754), .Z(n15660) );
  XNOR U20158 ( .A(n15653), .B(n15655), .Z(n15754) );
  NAND U20159 ( .A(n15755), .B(n15756), .Z(n15655) );
  OR U20160 ( .A(n15757), .B(n15758), .Z(n15756) );
  OR U20161 ( .A(n15759), .B(n15760), .Z(n15755) );
  NAND U20162 ( .A(n15761), .B(n15762), .Z(n15653) );
  OR U20163 ( .A(n15763), .B(n15764), .Z(n15762) );
  OR U20164 ( .A(n15765), .B(n15766), .Z(n15761) );
  ANDN U20165 ( .B(n15767), .A(n15768), .Z(n15654) );
  IV U20166 ( .A(n15769), .Z(n15767) );
  XNOR U20167 ( .A(n15734), .B(n15733), .Z(N28865) );
  XOR U20168 ( .A(n15753), .B(n15752), .Z(n15733) );
  XNOR U20169 ( .A(n15768), .B(n15769), .Z(n15752) );
  XNOR U20170 ( .A(n15763), .B(n15764), .Z(n15769) );
  XNOR U20171 ( .A(n15765), .B(n15766), .Z(n15764) );
  XNOR U20172 ( .A(y[1876]), .B(x[1876]), .Z(n15766) );
  XNOR U20173 ( .A(y[1877]), .B(x[1877]), .Z(n15765) );
  XNOR U20174 ( .A(y[1875]), .B(x[1875]), .Z(n15763) );
  XNOR U20175 ( .A(n15757), .B(n15758), .Z(n15768) );
  XNOR U20176 ( .A(y[1872]), .B(x[1872]), .Z(n15758) );
  XNOR U20177 ( .A(n15759), .B(n15760), .Z(n15757) );
  XNOR U20178 ( .A(y[1873]), .B(x[1873]), .Z(n15760) );
  XNOR U20179 ( .A(y[1874]), .B(x[1874]), .Z(n15759) );
  XNOR U20180 ( .A(n15750), .B(n15749), .Z(n15753) );
  XNOR U20181 ( .A(n15745), .B(n15746), .Z(n15749) );
  XNOR U20182 ( .A(y[1869]), .B(x[1869]), .Z(n15746) );
  XNOR U20183 ( .A(n15747), .B(n15748), .Z(n15745) );
  XNOR U20184 ( .A(y[1870]), .B(x[1870]), .Z(n15748) );
  XNOR U20185 ( .A(y[1871]), .B(x[1871]), .Z(n15747) );
  XNOR U20186 ( .A(n15739), .B(n15740), .Z(n15750) );
  XNOR U20187 ( .A(y[1866]), .B(x[1866]), .Z(n15740) );
  XNOR U20188 ( .A(n15741), .B(n15742), .Z(n15739) );
  XNOR U20189 ( .A(y[1867]), .B(x[1867]), .Z(n15742) );
  XNOR U20190 ( .A(y[1868]), .B(x[1868]), .Z(n15741) );
  XOR U20191 ( .A(n15715), .B(n15716), .Z(n15734) );
  XNOR U20192 ( .A(n15731), .B(n15732), .Z(n15716) );
  XNOR U20193 ( .A(n15726), .B(n15727), .Z(n15732) );
  XNOR U20194 ( .A(n15728), .B(n15729), .Z(n15727) );
  XNOR U20195 ( .A(y[1864]), .B(x[1864]), .Z(n15729) );
  XNOR U20196 ( .A(y[1865]), .B(x[1865]), .Z(n15728) );
  XNOR U20197 ( .A(y[1863]), .B(x[1863]), .Z(n15726) );
  XNOR U20198 ( .A(n15720), .B(n15721), .Z(n15731) );
  XNOR U20199 ( .A(y[1860]), .B(x[1860]), .Z(n15721) );
  XNOR U20200 ( .A(n15722), .B(n15723), .Z(n15720) );
  XNOR U20201 ( .A(y[1861]), .B(x[1861]), .Z(n15723) );
  XNOR U20202 ( .A(y[1862]), .B(x[1862]), .Z(n15722) );
  XOR U20203 ( .A(n15714), .B(n15713), .Z(n15715) );
  XNOR U20204 ( .A(n15709), .B(n15710), .Z(n15713) );
  XNOR U20205 ( .A(y[1857]), .B(x[1857]), .Z(n15710) );
  XNOR U20206 ( .A(n15711), .B(n15712), .Z(n15709) );
  XNOR U20207 ( .A(y[1858]), .B(x[1858]), .Z(n15712) );
  XNOR U20208 ( .A(y[1859]), .B(x[1859]), .Z(n15711) );
  XNOR U20209 ( .A(n15703), .B(n15704), .Z(n15714) );
  XNOR U20210 ( .A(y[1854]), .B(x[1854]), .Z(n15704) );
  XNOR U20211 ( .A(n15705), .B(n15706), .Z(n15703) );
  XNOR U20212 ( .A(y[1855]), .B(x[1855]), .Z(n15706) );
  XNOR U20213 ( .A(y[1856]), .B(x[1856]), .Z(n15705) );
  NAND U20214 ( .A(n15770), .B(n15771), .Z(N28857) );
  NANDN U20215 ( .A(n15772), .B(n15773), .Z(n15771) );
  OR U20216 ( .A(n15774), .B(n15775), .Z(n15773) );
  NAND U20217 ( .A(n15774), .B(n15775), .Z(n15770) );
  XOR U20218 ( .A(n15774), .B(n15776), .Z(N28856) );
  XNOR U20219 ( .A(n15772), .B(n15775), .Z(n15776) );
  AND U20220 ( .A(n15777), .B(n15778), .Z(n15775) );
  NANDN U20221 ( .A(n15779), .B(n15780), .Z(n15778) );
  NANDN U20222 ( .A(n15781), .B(n15782), .Z(n15780) );
  NANDN U20223 ( .A(n15782), .B(n15781), .Z(n15777) );
  NAND U20224 ( .A(n15783), .B(n15784), .Z(n15772) );
  NANDN U20225 ( .A(n15785), .B(n15786), .Z(n15784) );
  OR U20226 ( .A(n15787), .B(n15788), .Z(n15786) );
  NAND U20227 ( .A(n15788), .B(n15787), .Z(n15783) );
  AND U20228 ( .A(n15789), .B(n15790), .Z(n15774) );
  NANDN U20229 ( .A(n15791), .B(n15792), .Z(n15790) );
  NANDN U20230 ( .A(n15793), .B(n15794), .Z(n15792) );
  NANDN U20231 ( .A(n15794), .B(n15793), .Z(n15789) );
  XOR U20232 ( .A(n15788), .B(n15795), .Z(N28855) );
  XOR U20233 ( .A(n15785), .B(n15787), .Z(n15795) );
  XNOR U20234 ( .A(n15781), .B(n15796), .Z(n15787) );
  XNOR U20235 ( .A(n15779), .B(n15782), .Z(n15796) );
  NAND U20236 ( .A(n15797), .B(n15798), .Z(n15782) );
  NAND U20237 ( .A(n15799), .B(n15800), .Z(n15798) );
  OR U20238 ( .A(n15801), .B(n15802), .Z(n15799) );
  NANDN U20239 ( .A(n15803), .B(n15801), .Z(n15797) );
  IV U20240 ( .A(n15802), .Z(n15803) );
  NAND U20241 ( .A(n15804), .B(n15805), .Z(n15779) );
  NAND U20242 ( .A(n15806), .B(n15807), .Z(n15805) );
  NANDN U20243 ( .A(n15808), .B(n15809), .Z(n15806) );
  NANDN U20244 ( .A(n15809), .B(n15808), .Z(n15804) );
  AND U20245 ( .A(n15810), .B(n15811), .Z(n15781) );
  NAND U20246 ( .A(n15812), .B(n15813), .Z(n15811) );
  OR U20247 ( .A(n15814), .B(n15815), .Z(n15812) );
  NANDN U20248 ( .A(n15816), .B(n15814), .Z(n15810) );
  NAND U20249 ( .A(n15817), .B(n15818), .Z(n15785) );
  NANDN U20250 ( .A(n15819), .B(n15820), .Z(n15818) );
  OR U20251 ( .A(n15821), .B(n15822), .Z(n15820) );
  NANDN U20252 ( .A(n15823), .B(n15821), .Z(n15817) );
  IV U20253 ( .A(n15822), .Z(n15823) );
  XNOR U20254 ( .A(n15793), .B(n15824), .Z(n15788) );
  XNOR U20255 ( .A(n15791), .B(n15794), .Z(n15824) );
  NAND U20256 ( .A(n15825), .B(n15826), .Z(n15794) );
  NAND U20257 ( .A(n15827), .B(n15828), .Z(n15826) );
  OR U20258 ( .A(n15829), .B(n15830), .Z(n15827) );
  NANDN U20259 ( .A(n15831), .B(n15829), .Z(n15825) );
  IV U20260 ( .A(n15830), .Z(n15831) );
  NAND U20261 ( .A(n15832), .B(n15833), .Z(n15791) );
  NAND U20262 ( .A(n15834), .B(n15835), .Z(n15833) );
  NANDN U20263 ( .A(n15836), .B(n15837), .Z(n15834) );
  NANDN U20264 ( .A(n15837), .B(n15836), .Z(n15832) );
  AND U20265 ( .A(n15838), .B(n15839), .Z(n15793) );
  NAND U20266 ( .A(n15840), .B(n15841), .Z(n15839) );
  OR U20267 ( .A(n15842), .B(n15843), .Z(n15840) );
  NANDN U20268 ( .A(n15844), .B(n15842), .Z(n15838) );
  XNOR U20269 ( .A(n15819), .B(n15845), .Z(N28854) );
  XOR U20270 ( .A(n15821), .B(n15822), .Z(n15845) );
  XNOR U20271 ( .A(n15835), .B(n15846), .Z(n15822) );
  XOR U20272 ( .A(n15836), .B(n15837), .Z(n15846) );
  XOR U20273 ( .A(n15842), .B(n15847), .Z(n15837) );
  XOR U20274 ( .A(n15841), .B(n15844), .Z(n15847) );
  IV U20275 ( .A(n15843), .Z(n15844) );
  NAND U20276 ( .A(n15848), .B(n15849), .Z(n15843) );
  OR U20277 ( .A(n15850), .B(n15851), .Z(n15849) );
  OR U20278 ( .A(n15852), .B(n15853), .Z(n15848) );
  NAND U20279 ( .A(n15854), .B(n15855), .Z(n15841) );
  OR U20280 ( .A(n15856), .B(n15857), .Z(n15855) );
  OR U20281 ( .A(n15858), .B(n15859), .Z(n15854) );
  NOR U20282 ( .A(n15860), .B(n15861), .Z(n15842) );
  ANDN U20283 ( .B(n15862), .A(n15863), .Z(n15836) );
  XNOR U20284 ( .A(n15829), .B(n15864), .Z(n15835) );
  XNOR U20285 ( .A(n15828), .B(n15830), .Z(n15864) );
  NAND U20286 ( .A(n15865), .B(n15866), .Z(n15830) );
  OR U20287 ( .A(n15867), .B(n15868), .Z(n15866) );
  OR U20288 ( .A(n15869), .B(n15870), .Z(n15865) );
  NAND U20289 ( .A(n15871), .B(n15872), .Z(n15828) );
  OR U20290 ( .A(n15873), .B(n15874), .Z(n15872) );
  OR U20291 ( .A(n15875), .B(n15876), .Z(n15871) );
  ANDN U20292 ( .B(n15877), .A(n15878), .Z(n15829) );
  IV U20293 ( .A(n15879), .Z(n15877) );
  ANDN U20294 ( .B(n15880), .A(n15881), .Z(n15821) );
  XOR U20295 ( .A(n15807), .B(n15882), .Z(n15819) );
  XOR U20296 ( .A(n15808), .B(n15809), .Z(n15882) );
  XOR U20297 ( .A(n15814), .B(n15883), .Z(n15809) );
  XOR U20298 ( .A(n15813), .B(n15816), .Z(n15883) );
  IV U20299 ( .A(n15815), .Z(n15816) );
  NAND U20300 ( .A(n15884), .B(n15885), .Z(n15815) );
  OR U20301 ( .A(n15886), .B(n15887), .Z(n15885) );
  OR U20302 ( .A(n15888), .B(n15889), .Z(n15884) );
  NAND U20303 ( .A(n15890), .B(n15891), .Z(n15813) );
  OR U20304 ( .A(n15892), .B(n15893), .Z(n15891) );
  OR U20305 ( .A(n15894), .B(n15895), .Z(n15890) );
  NOR U20306 ( .A(n15896), .B(n15897), .Z(n15814) );
  ANDN U20307 ( .B(n15898), .A(n15899), .Z(n15808) );
  IV U20308 ( .A(n15900), .Z(n15898) );
  XNOR U20309 ( .A(n15801), .B(n15901), .Z(n15807) );
  XNOR U20310 ( .A(n15800), .B(n15802), .Z(n15901) );
  NAND U20311 ( .A(n15902), .B(n15903), .Z(n15802) );
  OR U20312 ( .A(n15904), .B(n15905), .Z(n15903) );
  OR U20313 ( .A(n15906), .B(n15907), .Z(n15902) );
  NAND U20314 ( .A(n15908), .B(n15909), .Z(n15800) );
  OR U20315 ( .A(n15910), .B(n15911), .Z(n15909) );
  OR U20316 ( .A(n15912), .B(n15913), .Z(n15908) );
  ANDN U20317 ( .B(n15914), .A(n15915), .Z(n15801) );
  IV U20318 ( .A(n15916), .Z(n15914) );
  XNOR U20319 ( .A(n15881), .B(n15880), .Z(N28853) );
  XOR U20320 ( .A(n15900), .B(n15899), .Z(n15880) );
  XNOR U20321 ( .A(n15915), .B(n15916), .Z(n15899) );
  XNOR U20322 ( .A(n15910), .B(n15911), .Z(n15916) );
  XNOR U20323 ( .A(n15912), .B(n15913), .Z(n15911) );
  XNOR U20324 ( .A(y[1852]), .B(x[1852]), .Z(n15913) );
  XNOR U20325 ( .A(y[1853]), .B(x[1853]), .Z(n15912) );
  XNOR U20326 ( .A(y[1851]), .B(x[1851]), .Z(n15910) );
  XNOR U20327 ( .A(n15904), .B(n15905), .Z(n15915) );
  XNOR U20328 ( .A(y[1848]), .B(x[1848]), .Z(n15905) );
  XNOR U20329 ( .A(n15906), .B(n15907), .Z(n15904) );
  XNOR U20330 ( .A(y[1849]), .B(x[1849]), .Z(n15907) );
  XNOR U20331 ( .A(y[1850]), .B(x[1850]), .Z(n15906) );
  XNOR U20332 ( .A(n15897), .B(n15896), .Z(n15900) );
  XNOR U20333 ( .A(n15892), .B(n15893), .Z(n15896) );
  XNOR U20334 ( .A(y[1845]), .B(x[1845]), .Z(n15893) );
  XNOR U20335 ( .A(n15894), .B(n15895), .Z(n15892) );
  XNOR U20336 ( .A(y[1846]), .B(x[1846]), .Z(n15895) );
  XNOR U20337 ( .A(y[1847]), .B(x[1847]), .Z(n15894) );
  XNOR U20338 ( .A(n15886), .B(n15887), .Z(n15897) );
  XNOR U20339 ( .A(y[1842]), .B(x[1842]), .Z(n15887) );
  XNOR U20340 ( .A(n15888), .B(n15889), .Z(n15886) );
  XNOR U20341 ( .A(y[1843]), .B(x[1843]), .Z(n15889) );
  XNOR U20342 ( .A(y[1844]), .B(x[1844]), .Z(n15888) );
  XOR U20343 ( .A(n15862), .B(n15863), .Z(n15881) );
  XNOR U20344 ( .A(n15878), .B(n15879), .Z(n15863) );
  XNOR U20345 ( .A(n15873), .B(n15874), .Z(n15879) );
  XNOR U20346 ( .A(n15875), .B(n15876), .Z(n15874) );
  XNOR U20347 ( .A(y[1840]), .B(x[1840]), .Z(n15876) );
  XNOR U20348 ( .A(y[1841]), .B(x[1841]), .Z(n15875) );
  XNOR U20349 ( .A(y[1839]), .B(x[1839]), .Z(n15873) );
  XNOR U20350 ( .A(n15867), .B(n15868), .Z(n15878) );
  XNOR U20351 ( .A(y[1836]), .B(x[1836]), .Z(n15868) );
  XNOR U20352 ( .A(n15869), .B(n15870), .Z(n15867) );
  XNOR U20353 ( .A(y[1837]), .B(x[1837]), .Z(n15870) );
  XNOR U20354 ( .A(y[1838]), .B(x[1838]), .Z(n15869) );
  XOR U20355 ( .A(n15861), .B(n15860), .Z(n15862) );
  XNOR U20356 ( .A(n15856), .B(n15857), .Z(n15860) );
  XNOR U20357 ( .A(y[1833]), .B(x[1833]), .Z(n15857) );
  XNOR U20358 ( .A(n15858), .B(n15859), .Z(n15856) );
  XNOR U20359 ( .A(y[1834]), .B(x[1834]), .Z(n15859) );
  XNOR U20360 ( .A(y[1835]), .B(x[1835]), .Z(n15858) );
  XNOR U20361 ( .A(n15850), .B(n15851), .Z(n15861) );
  XNOR U20362 ( .A(y[1830]), .B(x[1830]), .Z(n15851) );
  XNOR U20363 ( .A(n15852), .B(n15853), .Z(n15850) );
  XNOR U20364 ( .A(y[1831]), .B(x[1831]), .Z(n15853) );
  XNOR U20365 ( .A(y[1832]), .B(x[1832]), .Z(n15852) );
  NAND U20366 ( .A(n15917), .B(n15918), .Z(N28845) );
  NANDN U20367 ( .A(n15919), .B(n15920), .Z(n15918) );
  OR U20368 ( .A(n15921), .B(n15922), .Z(n15920) );
  NAND U20369 ( .A(n15921), .B(n15922), .Z(n15917) );
  XOR U20370 ( .A(n15921), .B(n15923), .Z(N28844) );
  XNOR U20371 ( .A(n15919), .B(n15922), .Z(n15923) );
  AND U20372 ( .A(n15924), .B(n15925), .Z(n15922) );
  NANDN U20373 ( .A(n15926), .B(n15927), .Z(n15925) );
  NANDN U20374 ( .A(n15928), .B(n15929), .Z(n15927) );
  NANDN U20375 ( .A(n15929), .B(n15928), .Z(n15924) );
  NAND U20376 ( .A(n15930), .B(n15931), .Z(n15919) );
  NANDN U20377 ( .A(n15932), .B(n15933), .Z(n15931) );
  OR U20378 ( .A(n15934), .B(n15935), .Z(n15933) );
  NAND U20379 ( .A(n15935), .B(n15934), .Z(n15930) );
  AND U20380 ( .A(n15936), .B(n15937), .Z(n15921) );
  NANDN U20381 ( .A(n15938), .B(n15939), .Z(n15937) );
  NANDN U20382 ( .A(n15940), .B(n15941), .Z(n15939) );
  NANDN U20383 ( .A(n15941), .B(n15940), .Z(n15936) );
  XOR U20384 ( .A(n15935), .B(n15942), .Z(N28843) );
  XOR U20385 ( .A(n15932), .B(n15934), .Z(n15942) );
  XNOR U20386 ( .A(n15928), .B(n15943), .Z(n15934) );
  XNOR U20387 ( .A(n15926), .B(n15929), .Z(n15943) );
  NAND U20388 ( .A(n15944), .B(n15945), .Z(n15929) );
  NAND U20389 ( .A(n15946), .B(n15947), .Z(n15945) );
  OR U20390 ( .A(n15948), .B(n15949), .Z(n15946) );
  NANDN U20391 ( .A(n15950), .B(n15948), .Z(n15944) );
  IV U20392 ( .A(n15949), .Z(n15950) );
  NAND U20393 ( .A(n15951), .B(n15952), .Z(n15926) );
  NAND U20394 ( .A(n15953), .B(n15954), .Z(n15952) );
  NANDN U20395 ( .A(n15955), .B(n15956), .Z(n15953) );
  NANDN U20396 ( .A(n15956), .B(n15955), .Z(n15951) );
  AND U20397 ( .A(n15957), .B(n15958), .Z(n15928) );
  NAND U20398 ( .A(n15959), .B(n15960), .Z(n15958) );
  OR U20399 ( .A(n15961), .B(n15962), .Z(n15959) );
  NANDN U20400 ( .A(n15963), .B(n15961), .Z(n15957) );
  NAND U20401 ( .A(n15964), .B(n15965), .Z(n15932) );
  NANDN U20402 ( .A(n15966), .B(n15967), .Z(n15965) );
  OR U20403 ( .A(n15968), .B(n15969), .Z(n15967) );
  NANDN U20404 ( .A(n15970), .B(n15968), .Z(n15964) );
  IV U20405 ( .A(n15969), .Z(n15970) );
  XNOR U20406 ( .A(n15940), .B(n15971), .Z(n15935) );
  XNOR U20407 ( .A(n15938), .B(n15941), .Z(n15971) );
  NAND U20408 ( .A(n15972), .B(n15973), .Z(n15941) );
  NAND U20409 ( .A(n15974), .B(n15975), .Z(n15973) );
  OR U20410 ( .A(n15976), .B(n15977), .Z(n15974) );
  NANDN U20411 ( .A(n15978), .B(n15976), .Z(n15972) );
  IV U20412 ( .A(n15977), .Z(n15978) );
  NAND U20413 ( .A(n15979), .B(n15980), .Z(n15938) );
  NAND U20414 ( .A(n15981), .B(n15982), .Z(n15980) );
  NANDN U20415 ( .A(n15983), .B(n15984), .Z(n15981) );
  NANDN U20416 ( .A(n15984), .B(n15983), .Z(n15979) );
  AND U20417 ( .A(n15985), .B(n15986), .Z(n15940) );
  NAND U20418 ( .A(n15987), .B(n15988), .Z(n15986) );
  OR U20419 ( .A(n15989), .B(n15990), .Z(n15987) );
  NANDN U20420 ( .A(n15991), .B(n15989), .Z(n15985) );
  XNOR U20421 ( .A(n15966), .B(n15992), .Z(N28842) );
  XOR U20422 ( .A(n15968), .B(n15969), .Z(n15992) );
  XNOR U20423 ( .A(n15982), .B(n15993), .Z(n15969) );
  XOR U20424 ( .A(n15983), .B(n15984), .Z(n15993) );
  XOR U20425 ( .A(n15989), .B(n15994), .Z(n15984) );
  XOR U20426 ( .A(n15988), .B(n15991), .Z(n15994) );
  IV U20427 ( .A(n15990), .Z(n15991) );
  NAND U20428 ( .A(n15995), .B(n15996), .Z(n15990) );
  OR U20429 ( .A(n15997), .B(n15998), .Z(n15996) );
  OR U20430 ( .A(n15999), .B(n16000), .Z(n15995) );
  NAND U20431 ( .A(n16001), .B(n16002), .Z(n15988) );
  OR U20432 ( .A(n16003), .B(n16004), .Z(n16002) );
  OR U20433 ( .A(n16005), .B(n16006), .Z(n16001) );
  NOR U20434 ( .A(n16007), .B(n16008), .Z(n15989) );
  ANDN U20435 ( .B(n16009), .A(n16010), .Z(n15983) );
  XNOR U20436 ( .A(n15976), .B(n16011), .Z(n15982) );
  XNOR U20437 ( .A(n15975), .B(n15977), .Z(n16011) );
  NAND U20438 ( .A(n16012), .B(n16013), .Z(n15977) );
  OR U20439 ( .A(n16014), .B(n16015), .Z(n16013) );
  OR U20440 ( .A(n16016), .B(n16017), .Z(n16012) );
  NAND U20441 ( .A(n16018), .B(n16019), .Z(n15975) );
  OR U20442 ( .A(n16020), .B(n16021), .Z(n16019) );
  OR U20443 ( .A(n16022), .B(n16023), .Z(n16018) );
  ANDN U20444 ( .B(n16024), .A(n16025), .Z(n15976) );
  IV U20445 ( .A(n16026), .Z(n16024) );
  ANDN U20446 ( .B(n16027), .A(n16028), .Z(n15968) );
  XOR U20447 ( .A(n15954), .B(n16029), .Z(n15966) );
  XOR U20448 ( .A(n15955), .B(n15956), .Z(n16029) );
  XOR U20449 ( .A(n15961), .B(n16030), .Z(n15956) );
  XOR U20450 ( .A(n15960), .B(n15963), .Z(n16030) );
  IV U20451 ( .A(n15962), .Z(n15963) );
  NAND U20452 ( .A(n16031), .B(n16032), .Z(n15962) );
  OR U20453 ( .A(n16033), .B(n16034), .Z(n16032) );
  OR U20454 ( .A(n16035), .B(n16036), .Z(n16031) );
  NAND U20455 ( .A(n16037), .B(n16038), .Z(n15960) );
  OR U20456 ( .A(n16039), .B(n16040), .Z(n16038) );
  OR U20457 ( .A(n16041), .B(n16042), .Z(n16037) );
  NOR U20458 ( .A(n16043), .B(n16044), .Z(n15961) );
  ANDN U20459 ( .B(n16045), .A(n16046), .Z(n15955) );
  IV U20460 ( .A(n16047), .Z(n16045) );
  XNOR U20461 ( .A(n15948), .B(n16048), .Z(n15954) );
  XNOR U20462 ( .A(n15947), .B(n15949), .Z(n16048) );
  NAND U20463 ( .A(n16049), .B(n16050), .Z(n15949) );
  OR U20464 ( .A(n16051), .B(n16052), .Z(n16050) );
  OR U20465 ( .A(n16053), .B(n16054), .Z(n16049) );
  NAND U20466 ( .A(n16055), .B(n16056), .Z(n15947) );
  OR U20467 ( .A(n16057), .B(n16058), .Z(n16056) );
  OR U20468 ( .A(n16059), .B(n16060), .Z(n16055) );
  ANDN U20469 ( .B(n16061), .A(n16062), .Z(n15948) );
  IV U20470 ( .A(n16063), .Z(n16061) );
  XNOR U20471 ( .A(n16028), .B(n16027), .Z(N28841) );
  XOR U20472 ( .A(n16047), .B(n16046), .Z(n16027) );
  XNOR U20473 ( .A(n16062), .B(n16063), .Z(n16046) );
  XNOR U20474 ( .A(n16057), .B(n16058), .Z(n16063) );
  XNOR U20475 ( .A(n16059), .B(n16060), .Z(n16058) );
  XNOR U20476 ( .A(y[1828]), .B(x[1828]), .Z(n16060) );
  XNOR U20477 ( .A(y[1829]), .B(x[1829]), .Z(n16059) );
  XNOR U20478 ( .A(y[1827]), .B(x[1827]), .Z(n16057) );
  XNOR U20479 ( .A(n16051), .B(n16052), .Z(n16062) );
  XNOR U20480 ( .A(y[1824]), .B(x[1824]), .Z(n16052) );
  XNOR U20481 ( .A(n16053), .B(n16054), .Z(n16051) );
  XNOR U20482 ( .A(y[1825]), .B(x[1825]), .Z(n16054) );
  XNOR U20483 ( .A(y[1826]), .B(x[1826]), .Z(n16053) );
  XNOR U20484 ( .A(n16044), .B(n16043), .Z(n16047) );
  XNOR U20485 ( .A(n16039), .B(n16040), .Z(n16043) );
  XNOR U20486 ( .A(y[1821]), .B(x[1821]), .Z(n16040) );
  XNOR U20487 ( .A(n16041), .B(n16042), .Z(n16039) );
  XNOR U20488 ( .A(y[1822]), .B(x[1822]), .Z(n16042) );
  XNOR U20489 ( .A(y[1823]), .B(x[1823]), .Z(n16041) );
  XNOR U20490 ( .A(n16033), .B(n16034), .Z(n16044) );
  XNOR U20491 ( .A(y[1818]), .B(x[1818]), .Z(n16034) );
  XNOR U20492 ( .A(n16035), .B(n16036), .Z(n16033) );
  XNOR U20493 ( .A(y[1819]), .B(x[1819]), .Z(n16036) );
  XNOR U20494 ( .A(y[1820]), .B(x[1820]), .Z(n16035) );
  XOR U20495 ( .A(n16009), .B(n16010), .Z(n16028) );
  XNOR U20496 ( .A(n16025), .B(n16026), .Z(n16010) );
  XNOR U20497 ( .A(n16020), .B(n16021), .Z(n16026) );
  XNOR U20498 ( .A(n16022), .B(n16023), .Z(n16021) );
  XNOR U20499 ( .A(y[1816]), .B(x[1816]), .Z(n16023) );
  XNOR U20500 ( .A(y[1817]), .B(x[1817]), .Z(n16022) );
  XNOR U20501 ( .A(y[1815]), .B(x[1815]), .Z(n16020) );
  XNOR U20502 ( .A(n16014), .B(n16015), .Z(n16025) );
  XNOR U20503 ( .A(y[1812]), .B(x[1812]), .Z(n16015) );
  XNOR U20504 ( .A(n16016), .B(n16017), .Z(n16014) );
  XNOR U20505 ( .A(y[1813]), .B(x[1813]), .Z(n16017) );
  XNOR U20506 ( .A(y[1814]), .B(x[1814]), .Z(n16016) );
  XOR U20507 ( .A(n16008), .B(n16007), .Z(n16009) );
  XNOR U20508 ( .A(n16003), .B(n16004), .Z(n16007) );
  XNOR U20509 ( .A(y[1809]), .B(x[1809]), .Z(n16004) );
  XNOR U20510 ( .A(n16005), .B(n16006), .Z(n16003) );
  XNOR U20511 ( .A(y[1810]), .B(x[1810]), .Z(n16006) );
  XNOR U20512 ( .A(y[1811]), .B(x[1811]), .Z(n16005) );
  XNOR U20513 ( .A(n15997), .B(n15998), .Z(n16008) );
  XNOR U20514 ( .A(y[1806]), .B(x[1806]), .Z(n15998) );
  XNOR U20515 ( .A(n15999), .B(n16000), .Z(n15997) );
  XNOR U20516 ( .A(y[1807]), .B(x[1807]), .Z(n16000) );
  XNOR U20517 ( .A(y[1808]), .B(x[1808]), .Z(n15999) );
  NAND U20518 ( .A(n16064), .B(n16065), .Z(N28833) );
  NANDN U20519 ( .A(n16066), .B(n16067), .Z(n16065) );
  OR U20520 ( .A(n16068), .B(n16069), .Z(n16067) );
  NAND U20521 ( .A(n16068), .B(n16069), .Z(n16064) );
  XOR U20522 ( .A(n16068), .B(n16070), .Z(N28832) );
  XNOR U20523 ( .A(n16066), .B(n16069), .Z(n16070) );
  AND U20524 ( .A(n16071), .B(n16072), .Z(n16069) );
  NANDN U20525 ( .A(n16073), .B(n16074), .Z(n16072) );
  NANDN U20526 ( .A(n16075), .B(n16076), .Z(n16074) );
  NANDN U20527 ( .A(n16076), .B(n16075), .Z(n16071) );
  NAND U20528 ( .A(n16077), .B(n16078), .Z(n16066) );
  NANDN U20529 ( .A(n16079), .B(n16080), .Z(n16078) );
  OR U20530 ( .A(n16081), .B(n16082), .Z(n16080) );
  NAND U20531 ( .A(n16082), .B(n16081), .Z(n16077) );
  AND U20532 ( .A(n16083), .B(n16084), .Z(n16068) );
  NANDN U20533 ( .A(n16085), .B(n16086), .Z(n16084) );
  NANDN U20534 ( .A(n16087), .B(n16088), .Z(n16086) );
  NANDN U20535 ( .A(n16088), .B(n16087), .Z(n16083) );
  XOR U20536 ( .A(n16082), .B(n16089), .Z(N28831) );
  XOR U20537 ( .A(n16079), .B(n16081), .Z(n16089) );
  XNOR U20538 ( .A(n16075), .B(n16090), .Z(n16081) );
  XNOR U20539 ( .A(n16073), .B(n16076), .Z(n16090) );
  NAND U20540 ( .A(n16091), .B(n16092), .Z(n16076) );
  NAND U20541 ( .A(n16093), .B(n16094), .Z(n16092) );
  OR U20542 ( .A(n16095), .B(n16096), .Z(n16093) );
  NANDN U20543 ( .A(n16097), .B(n16095), .Z(n16091) );
  IV U20544 ( .A(n16096), .Z(n16097) );
  NAND U20545 ( .A(n16098), .B(n16099), .Z(n16073) );
  NAND U20546 ( .A(n16100), .B(n16101), .Z(n16099) );
  NANDN U20547 ( .A(n16102), .B(n16103), .Z(n16100) );
  NANDN U20548 ( .A(n16103), .B(n16102), .Z(n16098) );
  AND U20549 ( .A(n16104), .B(n16105), .Z(n16075) );
  NAND U20550 ( .A(n16106), .B(n16107), .Z(n16105) );
  OR U20551 ( .A(n16108), .B(n16109), .Z(n16106) );
  NANDN U20552 ( .A(n16110), .B(n16108), .Z(n16104) );
  NAND U20553 ( .A(n16111), .B(n16112), .Z(n16079) );
  NANDN U20554 ( .A(n16113), .B(n16114), .Z(n16112) );
  OR U20555 ( .A(n16115), .B(n16116), .Z(n16114) );
  NANDN U20556 ( .A(n16117), .B(n16115), .Z(n16111) );
  IV U20557 ( .A(n16116), .Z(n16117) );
  XNOR U20558 ( .A(n16087), .B(n16118), .Z(n16082) );
  XNOR U20559 ( .A(n16085), .B(n16088), .Z(n16118) );
  NAND U20560 ( .A(n16119), .B(n16120), .Z(n16088) );
  NAND U20561 ( .A(n16121), .B(n16122), .Z(n16120) );
  OR U20562 ( .A(n16123), .B(n16124), .Z(n16121) );
  NANDN U20563 ( .A(n16125), .B(n16123), .Z(n16119) );
  IV U20564 ( .A(n16124), .Z(n16125) );
  NAND U20565 ( .A(n16126), .B(n16127), .Z(n16085) );
  NAND U20566 ( .A(n16128), .B(n16129), .Z(n16127) );
  NANDN U20567 ( .A(n16130), .B(n16131), .Z(n16128) );
  NANDN U20568 ( .A(n16131), .B(n16130), .Z(n16126) );
  AND U20569 ( .A(n16132), .B(n16133), .Z(n16087) );
  NAND U20570 ( .A(n16134), .B(n16135), .Z(n16133) );
  OR U20571 ( .A(n16136), .B(n16137), .Z(n16134) );
  NANDN U20572 ( .A(n16138), .B(n16136), .Z(n16132) );
  XNOR U20573 ( .A(n16113), .B(n16139), .Z(N28830) );
  XOR U20574 ( .A(n16115), .B(n16116), .Z(n16139) );
  XNOR U20575 ( .A(n16129), .B(n16140), .Z(n16116) );
  XOR U20576 ( .A(n16130), .B(n16131), .Z(n16140) );
  XOR U20577 ( .A(n16136), .B(n16141), .Z(n16131) );
  XOR U20578 ( .A(n16135), .B(n16138), .Z(n16141) );
  IV U20579 ( .A(n16137), .Z(n16138) );
  NAND U20580 ( .A(n16142), .B(n16143), .Z(n16137) );
  OR U20581 ( .A(n16144), .B(n16145), .Z(n16143) );
  OR U20582 ( .A(n16146), .B(n16147), .Z(n16142) );
  NAND U20583 ( .A(n16148), .B(n16149), .Z(n16135) );
  OR U20584 ( .A(n16150), .B(n16151), .Z(n16149) );
  OR U20585 ( .A(n16152), .B(n16153), .Z(n16148) );
  NOR U20586 ( .A(n16154), .B(n16155), .Z(n16136) );
  ANDN U20587 ( .B(n16156), .A(n16157), .Z(n16130) );
  XNOR U20588 ( .A(n16123), .B(n16158), .Z(n16129) );
  XNOR U20589 ( .A(n16122), .B(n16124), .Z(n16158) );
  NAND U20590 ( .A(n16159), .B(n16160), .Z(n16124) );
  OR U20591 ( .A(n16161), .B(n16162), .Z(n16160) );
  OR U20592 ( .A(n16163), .B(n16164), .Z(n16159) );
  NAND U20593 ( .A(n16165), .B(n16166), .Z(n16122) );
  OR U20594 ( .A(n16167), .B(n16168), .Z(n16166) );
  OR U20595 ( .A(n16169), .B(n16170), .Z(n16165) );
  ANDN U20596 ( .B(n16171), .A(n16172), .Z(n16123) );
  IV U20597 ( .A(n16173), .Z(n16171) );
  ANDN U20598 ( .B(n16174), .A(n16175), .Z(n16115) );
  XOR U20599 ( .A(n16101), .B(n16176), .Z(n16113) );
  XOR U20600 ( .A(n16102), .B(n16103), .Z(n16176) );
  XOR U20601 ( .A(n16108), .B(n16177), .Z(n16103) );
  XOR U20602 ( .A(n16107), .B(n16110), .Z(n16177) );
  IV U20603 ( .A(n16109), .Z(n16110) );
  NAND U20604 ( .A(n16178), .B(n16179), .Z(n16109) );
  OR U20605 ( .A(n16180), .B(n16181), .Z(n16179) );
  OR U20606 ( .A(n16182), .B(n16183), .Z(n16178) );
  NAND U20607 ( .A(n16184), .B(n16185), .Z(n16107) );
  OR U20608 ( .A(n16186), .B(n16187), .Z(n16185) );
  OR U20609 ( .A(n16188), .B(n16189), .Z(n16184) );
  NOR U20610 ( .A(n16190), .B(n16191), .Z(n16108) );
  ANDN U20611 ( .B(n16192), .A(n16193), .Z(n16102) );
  IV U20612 ( .A(n16194), .Z(n16192) );
  XNOR U20613 ( .A(n16095), .B(n16195), .Z(n16101) );
  XNOR U20614 ( .A(n16094), .B(n16096), .Z(n16195) );
  NAND U20615 ( .A(n16196), .B(n16197), .Z(n16096) );
  OR U20616 ( .A(n16198), .B(n16199), .Z(n16197) );
  OR U20617 ( .A(n16200), .B(n16201), .Z(n16196) );
  NAND U20618 ( .A(n16202), .B(n16203), .Z(n16094) );
  OR U20619 ( .A(n16204), .B(n16205), .Z(n16203) );
  OR U20620 ( .A(n16206), .B(n16207), .Z(n16202) );
  ANDN U20621 ( .B(n16208), .A(n16209), .Z(n16095) );
  IV U20622 ( .A(n16210), .Z(n16208) );
  XNOR U20623 ( .A(n16175), .B(n16174), .Z(N28829) );
  XOR U20624 ( .A(n16194), .B(n16193), .Z(n16174) );
  XNOR U20625 ( .A(n16209), .B(n16210), .Z(n16193) );
  XNOR U20626 ( .A(n16204), .B(n16205), .Z(n16210) );
  XNOR U20627 ( .A(n16206), .B(n16207), .Z(n16205) );
  XNOR U20628 ( .A(y[1804]), .B(x[1804]), .Z(n16207) );
  XNOR U20629 ( .A(y[1805]), .B(x[1805]), .Z(n16206) );
  XNOR U20630 ( .A(y[1803]), .B(x[1803]), .Z(n16204) );
  XNOR U20631 ( .A(n16198), .B(n16199), .Z(n16209) );
  XNOR U20632 ( .A(y[1800]), .B(x[1800]), .Z(n16199) );
  XNOR U20633 ( .A(n16200), .B(n16201), .Z(n16198) );
  XNOR U20634 ( .A(y[1801]), .B(x[1801]), .Z(n16201) );
  XNOR U20635 ( .A(y[1802]), .B(x[1802]), .Z(n16200) );
  XNOR U20636 ( .A(n16191), .B(n16190), .Z(n16194) );
  XNOR U20637 ( .A(n16186), .B(n16187), .Z(n16190) );
  XNOR U20638 ( .A(y[1797]), .B(x[1797]), .Z(n16187) );
  XNOR U20639 ( .A(n16188), .B(n16189), .Z(n16186) );
  XNOR U20640 ( .A(y[1798]), .B(x[1798]), .Z(n16189) );
  XNOR U20641 ( .A(y[1799]), .B(x[1799]), .Z(n16188) );
  XNOR U20642 ( .A(n16180), .B(n16181), .Z(n16191) );
  XNOR U20643 ( .A(y[1794]), .B(x[1794]), .Z(n16181) );
  XNOR U20644 ( .A(n16182), .B(n16183), .Z(n16180) );
  XNOR U20645 ( .A(y[1795]), .B(x[1795]), .Z(n16183) );
  XNOR U20646 ( .A(y[1796]), .B(x[1796]), .Z(n16182) );
  XOR U20647 ( .A(n16156), .B(n16157), .Z(n16175) );
  XNOR U20648 ( .A(n16172), .B(n16173), .Z(n16157) );
  XNOR U20649 ( .A(n16167), .B(n16168), .Z(n16173) );
  XNOR U20650 ( .A(n16169), .B(n16170), .Z(n16168) );
  XNOR U20651 ( .A(y[1792]), .B(x[1792]), .Z(n16170) );
  XNOR U20652 ( .A(y[1793]), .B(x[1793]), .Z(n16169) );
  XNOR U20653 ( .A(y[1791]), .B(x[1791]), .Z(n16167) );
  XNOR U20654 ( .A(n16161), .B(n16162), .Z(n16172) );
  XNOR U20655 ( .A(y[1788]), .B(x[1788]), .Z(n16162) );
  XNOR U20656 ( .A(n16163), .B(n16164), .Z(n16161) );
  XNOR U20657 ( .A(y[1789]), .B(x[1789]), .Z(n16164) );
  XNOR U20658 ( .A(y[1790]), .B(x[1790]), .Z(n16163) );
  XOR U20659 ( .A(n16155), .B(n16154), .Z(n16156) );
  XNOR U20660 ( .A(n16150), .B(n16151), .Z(n16154) );
  XNOR U20661 ( .A(y[1785]), .B(x[1785]), .Z(n16151) );
  XNOR U20662 ( .A(n16152), .B(n16153), .Z(n16150) );
  XNOR U20663 ( .A(y[1786]), .B(x[1786]), .Z(n16153) );
  XNOR U20664 ( .A(y[1787]), .B(x[1787]), .Z(n16152) );
  XNOR U20665 ( .A(n16144), .B(n16145), .Z(n16155) );
  XNOR U20666 ( .A(y[1782]), .B(x[1782]), .Z(n16145) );
  XNOR U20667 ( .A(n16146), .B(n16147), .Z(n16144) );
  XNOR U20668 ( .A(y[1783]), .B(x[1783]), .Z(n16147) );
  XNOR U20669 ( .A(y[1784]), .B(x[1784]), .Z(n16146) );
  NAND U20670 ( .A(n16211), .B(n16212), .Z(N28821) );
  NANDN U20671 ( .A(n16213), .B(n16214), .Z(n16212) );
  OR U20672 ( .A(n16215), .B(n16216), .Z(n16214) );
  NAND U20673 ( .A(n16215), .B(n16216), .Z(n16211) );
  XOR U20674 ( .A(n16215), .B(n16217), .Z(N28820) );
  XNOR U20675 ( .A(n16213), .B(n16216), .Z(n16217) );
  AND U20676 ( .A(n16218), .B(n16219), .Z(n16216) );
  NANDN U20677 ( .A(n16220), .B(n16221), .Z(n16219) );
  NANDN U20678 ( .A(n16222), .B(n16223), .Z(n16221) );
  NANDN U20679 ( .A(n16223), .B(n16222), .Z(n16218) );
  NAND U20680 ( .A(n16224), .B(n16225), .Z(n16213) );
  NANDN U20681 ( .A(n16226), .B(n16227), .Z(n16225) );
  OR U20682 ( .A(n16228), .B(n16229), .Z(n16227) );
  NAND U20683 ( .A(n16229), .B(n16228), .Z(n16224) );
  AND U20684 ( .A(n16230), .B(n16231), .Z(n16215) );
  NANDN U20685 ( .A(n16232), .B(n16233), .Z(n16231) );
  NANDN U20686 ( .A(n16234), .B(n16235), .Z(n16233) );
  NANDN U20687 ( .A(n16235), .B(n16234), .Z(n16230) );
  XOR U20688 ( .A(n16229), .B(n16236), .Z(N28819) );
  XOR U20689 ( .A(n16226), .B(n16228), .Z(n16236) );
  XNOR U20690 ( .A(n16222), .B(n16237), .Z(n16228) );
  XNOR U20691 ( .A(n16220), .B(n16223), .Z(n16237) );
  NAND U20692 ( .A(n16238), .B(n16239), .Z(n16223) );
  NAND U20693 ( .A(n16240), .B(n16241), .Z(n16239) );
  OR U20694 ( .A(n16242), .B(n16243), .Z(n16240) );
  NANDN U20695 ( .A(n16244), .B(n16242), .Z(n16238) );
  IV U20696 ( .A(n16243), .Z(n16244) );
  NAND U20697 ( .A(n16245), .B(n16246), .Z(n16220) );
  NAND U20698 ( .A(n16247), .B(n16248), .Z(n16246) );
  NANDN U20699 ( .A(n16249), .B(n16250), .Z(n16247) );
  NANDN U20700 ( .A(n16250), .B(n16249), .Z(n16245) );
  AND U20701 ( .A(n16251), .B(n16252), .Z(n16222) );
  NAND U20702 ( .A(n16253), .B(n16254), .Z(n16252) );
  OR U20703 ( .A(n16255), .B(n16256), .Z(n16253) );
  NANDN U20704 ( .A(n16257), .B(n16255), .Z(n16251) );
  NAND U20705 ( .A(n16258), .B(n16259), .Z(n16226) );
  NANDN U20706 ( .A(n16260), .B(n16261), .Z(n16259) );
  OR U20707 ( .A(n16262), .B(n16263), .Z(n16261) );
  NANDN U20708 ( .A(n16264), .B(n16262), .Z(n16258) );
  IV U20709 ( .A(n16263), .Z(n16264) );
  XNOR U20710 ( .A(n16234), .B(n16265), .Z(n16229) );
  XNOR U20711 ( .A(n16232), .B(n16235), .Z(n16265) );
  NAND U20712 ( .A(n16266), .B(n16267), .Z(n16235) );
  NAND U20713 ( .A(n16268), .B(n16269), .Z(n16267) );
  OR U20714 ( .A(n16270), .B(n16271), .Z(n16268) );
  NANDN U20715 ( .A(n16272), .B(n16270), .Z(n16266) );
  IV U20716 ( .A(n16271), .Z(n16272) );
  NAND U20717 ( .A(n16273), .B(n16274), .Z(n16232) );
  NAND U20718 ( .A(n16275), .B(n16276), .Z(n16274) );
  NANDN U20719 ( .A(n16277), .B(n16278), .Z(n16275) );
  NANDN U20720 ( .A(n16278), .B(n16277), .Z(n16273) );
  AND U20721 ( .A(n16279), .B(n16280), .Z(n16234) );
  NAND U20722 ( .A(n16281), .B(n16282), .Z(n16280) );
  OR U20723 ( .A(n16283), .B(n16284), .Z(n16281) );
  NANDN U20724 ( .A(n16285), .B(n16283), .Z(n16279) );
  XNOR U20725 ( .A(n16260), .B(n16286), .Z(N28818) );
  XOR U20726 ( .A(n16262), .B(n16263), .Z(n16286) );
  XNOR U20727 ( .A(n16276), .B(n16287), .Z(n16263) );
  XOR U20728 ( .A(n16277), .B(n16278), .Z(n16287) );
  XOR U20729 ( .A(n16283), .B(n16288), .Z(n16278) );
  XOR U20730 ( .A(n16282), .B(n16285), .Z(n16288) );
  IV U20731 ( .A(n16284), .Z(n16285) );
  NAND U20732 ( .A(n16289), .B(n16290), .Z(n16284) );
  OR U20733 ( .A(n16291), .B(n16292), .Z(n16290) );
  OR U20734 ( .A(n16293), .B(n16294), .Z(n16289) );
  NAND U20735 ( .A(n16295), .B(n16296), .Z(n16282) );
  OR U20736 ( .A(n16297), .B(n16298), .Z(n16296) );
  OR U20737 ( .A(n16299), .B(n16300), .Z(n16295) );
  NOR U20738 ( .A(n16301), .B(n16302), .Z(n16283) );
  ANDN U20739 ( .B(n16303), .A(n16304), .Z(n16277) );
  XNOR U20740 ( .A(n16270), .B(n16305), .Z(n16276) );
  XNOR U20741 ( .A(n16269), .B(n16271), .Z(n16305) );
  NAND U20742 ( .A(n16306), .B(n16307), .Z(n16271) );
  OR U20743 ( .A(n16308), .B(n16309), .Z(n16307) );
  OR U20744 ( .A(n16310), .B(n16311), .Z(n16306) );
  NAND U20745 ( .A(n16312), .B(n16313), .Z(n16269) );
  OR U20746 ( .A(n16314), .B(n16315), .Z(n16313) );
  OR U20747 ( .A(n16316), .B(n16317), .Z(n16312) );
  ANDN U20748 ( .B(n16318), .A(n16319), .Z(n16270) );
  IV U20749 ( .A(n16320), .Z(n16318) );
  ANDN U20750 ( .B(n16321), .A(n16322), .Z(n16262) );
  XOR U20751 ( .A(n16248), .B(n16323), .Z(n16260) );
  XOR U20752 ( .A(n16249), .B(n16250), .Z(n16323) );
  XOR U20753 ( .A(n16255), .B(n16324), .Z(n16250) );
  XOR U20754 ( .A(n16254), .B(n16257), .Z(n16324) );
  IV U20755 ( .A(n16256), .Z(n16257) );
  NAND U20756 ( .A(n16325), .B(n16326), .Z(n16256) );
  OR U20757 ( .A(n16327), .B(n16328), .Z(n16326) );
  OR U20758 ( .A(n16329), .B(n16330), .Z(n16325) );
  NAND U20759 ( .A(n16331), .B(n16332), .Z(n16254) );
  OR U20760 ( .A(n16333), .B(n16334), .Z(n16332) );
  OR U20761 ( .A(n16335), .B(n16336), .Z(n16331) );
  NOR U20762 ( .A(n16337), .B(n16338), .Z(n16255) );
  ANDN U20763 ( .B(n16339), .A(n16340), .Z(n16249) );
  IV U20764 ( .A(n16341), .Z(n16339) );
  XNOR U20765 ( .A(n16242), .B(n16342), .Z(n16248) );
  XNOR U20766 ( .A(n16241), .B(n16243), .Z(n16342) );
  NAND U20767 ( .A(n16343), .B(n16344), .Z(n16243) );
  OR U20768 ( .A(n16345), .B(n16346), .Z(n16344) );
  OR U20769 ( .A(n16347), .B(n16348), .Z(n16343) );
  NAND U20770 ( .A(n16349), .B(n16350), .Z(n16241) );
  OR U20771 ( .A(n16351), .B(n16352), .Z(n16350) );
  OR U20772 ( .A(n16353), .B(n16354), .Z(n16349) );
  ANDN U20773 ( .B(n16355), .A(n16356), .Z(n16242) );
  IV U20774 ( .A(n16357), .Z(n16355) );
  XNOR U20775 ( .A(n16322), .B(n16321), .Z(N28817) );
  XOR U20776 ( .A(n16341), .B(n16340), .Z(n16321) );
  XNOR U20777 ( .A(n16356), .B(n16357), .Z(n16340) );
  XNOR U20778 ( .A(n16351), .B(n16352), .Z(n16357) );
  XNOR U20779 ( .A(n16353), .B(n16354), .Z(n16352) );
  XNOR U20780 ( .A(y[1780]), .B(x[1780]), .Z(n16354) );
  XNOR U20781 ( .A(y[1781]), .B(x[1781]), .Z(n16353) );
  XNOR U20782 ( .A(y[1779]), .B(x[1779]), .Z(n16351) );
  XNOR U20783 ( .A(n16345), .B(n16346), .Z(n16356) );
  XNOR U20784 ( .A(y[1776]), .B(x[1776]), .Z(n16346) );
  XNOR U20785 ( .A(n16347), .B(n16348), .Z(n16345) );
  XNOR U20786 ( .A(y[1777]), .B(x[1777]), .Z(n16348) );
  XNOR U20787 ( .A(y[1778]), .B(x[1778]), .Z(n16347) );
  XNOR U20788 ( .A(n16338), .B(n16337), .Z(n16341) );
  XNOR U20789 ( .A(n16333), .B(n16334), .Z(n16337) );
  XNOR U20790 ( .A(y[1773]), .B(x[1773]), .Z(n16334) );
  XNOR U20791 ( .A(n16335), .B(n16336), .Z(n16333) );
  XNOR U20792 ( .A(y[1774]), .B(x[1774]), .Z(n16336) );
  XNOR U20793 ( .A(y[1775]), .B(x[1775]), .Z(n16335) );
  XNOR U20794 ( .A(n16327), .B(n16328), .Z(n16338) );
  XNOR U20795 ( .A(y[1770]), .B(x[1770]), .Z(n16328) );
  XNOR U20796 ( .A(n16329), .B(n16330), .Z(n16327) );
  XNOR U20797 ( .A(y[1771]), .B(x[1771]), .Z(n16330) );
  XNOR U20798 ( .A(y[1772]), .B(x[1772]), .Z(n16329) );
  XOR U20799 ( .A(n16303), .B(n16304), .Z(n16322) );
  XNOR U20800 ( .A(n16319), .B(n16320), .Z(n16304) );
  XNOR U20801 ( .A(n16314), .B(n16315), .Z(n16320) );
  XNOR U20802 ( .A(n16316), .B(n16317), .Z(n16315) );
  XNOR U20803 ( .A(y[1768]), .B(x[1768]), .Z(n16317) );
  XNOR U20804 ( .A(y[1769]), .B(x[1769]), .Z(n16316) );
  XNOR U20805 ( .A(y[1767]), .B(x[1767]), .Z(n16314) );
  XNOR U20806 ( .A(n16308), .B(n16309), .Z(n16319) );
  XNOR U20807 ( .A(y[1764]), .B(x[1764]), .Z(n16309) );
  XNOR U20808 ( .A(n16310), .B(n16311), .Z(n16308) );
  XNOR U20809 ( .A(y[1765]), .B(x[1765]), .Z(n16311) );
  XNOR U20810 ( .A(y[1766]), .B(x[1766]), .Z(n16310) );
  XOR U20811 ( .A(n16302), .B(n16301), .Z(n16303) );
  XNOR U20812 ( .A(n16297), .B(n16298), .Z(n16301) );
  XNOR U20813 ( .A(y[1761]), .B(x[1761]), .Z(n16298) );
  XNOR U20814 ( .A(n16299), .B(n16300), .Z(n16297) );
  XNOR U20815 ( .A(y[1762]), .B(x[1762]), .Z(n16300) );
  XNOR U20816 ( .A(y[1763]), .B(x[1763]), .Z(n16299) );
  XNOR U20817 ( .A(n16291), .B(n16292), .Z(n16302) );
  XNOR U20818 ( .A(y[1758]), .B(x[1758]), .Z(n16292) );
  XNOR U20819 ( .A(n16293), .B(n16294), .Z(n16291) );
  XNOR U20820 ( .A(y[1759]), .B(x[1759]), .Z(n16294) );
  XNOR U20821 ( .A(y[1760]), .B(x[1760]), .Z(n16293) );
  NAND U20822 ( .A(n16358), .B(n16359), .Z(N28809) );
  NANDN U20823 ( .A(n16360), .B(n16361), .Z(n16359) );
  OR U20824 ( .A(n16362), .B(n16363), .Z(n16361) );
  NAND U20825 ( .A(n16362), .B(n16363), .Z(n16358) );
  XOR U20826 ( .A(n16362), .B(n16364), .Z(N28808) );
  XNOR U20827 ( .A(n16360), .B(n16363), .Z(n16364) );
  AND U20828 ( .A(n16365), .B(n16366), .Z(n16363) );
  NANDN U20829 ( .A(n16367), .B(n16368), .Z(n16366) );
  NANDN U20830 ( .A(n16369), .B(n16370), .Z(n16368) );
  NANDN U20831 ( .A(n16370), .B(n16369), .Z(n16365) );
  NAND U20832 ( .A(n16371), .B(n16372), .Z(n16360) );
  NANDN U20833 ( .A(n16373), .B(n16374), .Z(n16372) );
  OR U20834 ( .A(n16375), .B(n16376), .Z(n16374) );
  NAND U20835 ( .A(n16376), .B(n16375), .Z(n16371) );
  AND U20836 ( .A(n16377), .B(n16378), .Z(n16362) );
  NANDN U20837 ( .A(n16379), .B(n16380), .Z(n16378) );
  NANDN U20838 ( .A(n16381), .B(n16382), .Z(n16380) );
  NANDN U20839 ( .A(n16382), .B(n16381), .Z(n16377) );
  XOR U20840 ( .A(n16376), .B(n16383), .Z(N28807) );
  XOR U20841 ( .A(n16373), .B(n16375), .Z(n16383) );
  XNOR U20842 ( .A(n16369), .B(n16384), .Z(n16375) );
  XNOR U20843 ( .A(n16367), .B(n16370), .Z(n16384) );
  NAND U20844 ( .A(n16385), .B(n16386), .Z(n16370) );
  NAND U20845 ( .A(n16387), .B(n16388), .Z(n16386) );
  OR U20846 ( .A(n16389), .B(n16390), .Z(n16387) );
  NANDN U20847 ( .A(n16391), .B(n16389), .Z(n16385) );
  IV U20848 ( .A(n16390), .Z(n16391) );
  NAND U20849 ( .A(n16392), .B(n16393), .Z(n16367) );
  NAND U20850 ( .A(n16394), .B(n16395), .Z(n16393) );
  NANDN U20851 ( .A(n16396), .B(n16397), .Z(n16394) );
  NANDN U20852 ( .A(n16397), .B(n16396), .Z(n16392) );
  AND U20853 ( .A(n16398), .B(n16399), .Z(n16369) );
  NAND U20854 ( .A(n16400), .B(n16401), .Z(n16399) );
  OR U20855 ( .A(n16402), .B(n16403), .Z(n16400) );
  NANDN U20856 ( .A(n16404), .B(n16402), .Z(n16398) );
  NAND U20857 ( .A(n16405), .B(n16406), .Z(n16373) );
  NANDN U20858 ( .A(n16407), .B(n16408), .Z(n16406) );
  OR U20859 ( .A(n16409), .B(n16410), .Z(n16408) );
  NANDN U20860 ( .A(n16411), .B(n16409), .Z(n16405) );
  IV U20861 ( .A(n16410), .Z(n16411) );
  XNOR U20862 ( .A(n16381), .B(n16412), .Z(n16376) );
  XNOR U20863 ( .A(n16379), .B(n16382), .Z(n16412) );
  NAND U20864 ( .A(n16413), .B(n16414), .Z(n16382) );
  NAND U20865 ( .A(n16415), .B(n16416), .Z(n16414) );
  OR U20866 ( .A(n16417), .B(n16418), .Z(n16415) );
  NANDN U20867 ( .A(n16419), .B(n16417), .Z(n16413) );
  IV U20868 ( .A(n16418), .Z(n16419) );
  NAND U20869 ( .A(n16420), .B(n16421), .Z(n16379) );
  NAND U20870 ( .A(n16422), .B(n16423), .Z(n16421) );
  NANDN U20871 ( .A(n16424), .B(n16425), .Z(n16422) );
  NANDN U20872 ( .A(n16425), .B(n16424), .Z(n16420) );
  AND U20873 ( .A(n16426), .B(n16427), .Z(n16381) );
  NAND U20874 ( .A(n16428), .B(n16429), .Z(n16427) );
  OR U20875 ( .A(n16430), .B(n16431), .Z(n16428) );
  NANDN U20876 ( .A(n16432), .B(n16430), .Z(n16426) );
  XNOR U20877 ( .A(n16407), .B(n16433), .Z(N28806) );
  XOR U20878 ( .A(n16409), .B(n16410), .Z(n16433) );
  XNOR U20879 ( .A(n16423), .B(n16434), .Z(n16410) );
  XOR U20880 ( .A(n16424), .B(n16425), .Z(n16434) );
  XOR U20881 ( .A(n16430), .B(n16435), .Z(n16425) );
  XOR U20882 ( .A(n16429), .B(n16432), .Z(n16435) );
  IV U20883 ( .A(n16431), .Z(n16432) );
  NAND U20884 ( .A(n16436), .B(n16437), .Z(n16431) );
  OR U20885 ( .A(n16438), .B(n16439), .Z(n16437) );
  OR U20886 ( .A(n16440), .B(n16441), .Z(n16436) );
  NAND U20887 ( .A(n16442), .B(n16443), .Z(n16429) );
  OR U20888 ( .A(n16444), .B(n16445), .Z(n16443) );
  OR U20889 ( .A(n16446), .B(n16447), .Z(n16442) );
  NOR U20890 ( .A(n16448), .B(n16449), .Z(n16430) );
  ANDN U20891 ( .B(n16450), .A(n16451), .Z(n16424) );
  XNOR U20892 ( .A(n16417), .B(n16452), .Z(n16423) );
  XNOR U20893 ( .A(n16416), .B(n16418), .Z(n16452) );
  NAND U20894 ( .A(n16453), .B(n16454), .Z(n16418) );
  OR U20895 ( .A(n16455), .B(n16456), .Z(n16454) );
  OR U20896 ( .A(n16457), .B(n16458), .Z(n16453) );
  NAND U20897 ( .A(n16459), .B(n16460), .Z(n16416) );
  OR U20898 ( .A(n16461), .B(n16462), .Z(n16460) );
  OR U20899 ( .A(n16463), .B(n16464), .Z(n16459) );
  ANDN U20900 ( .B(n16465), .A(n16466), .Z(n16417) );
  IV U20901 ( .A(n16467), .Z(n16465) );
  ANDN U20902 ( .B(n16468), .A(n16469), .Z(n16409) );
  XOR U20903 ( .A(n16395), .B(n16470), .Z(n16407) );
  XOR U20904 ( .A(n16396), .B(n16397), .Z(n16470) );
  XOR U20905 ( .A(n16402), .B(n16471), .Z(n16397) );
  XOR U20906 ( .A(n16401), .B(n16404), .Z(n16471) );
  IV U20907 ( .A(n16403), .Z(n16404) );
  NAND U20908 ( .A(n16472), .B(n16473), .Z(n16403) );
  OR U20909 ( .A(n16474), .B(n16475), .Z(n16473) );
  OR U20910 ( .A(n16476), .B(n16477), .Z(n16472) );
  NAND U20911 ( .A(n16478), .B(n16479), .Z(n16401) );
  OR U20912 ( .A(n16480), .B(n16481), .Z(n16479) );
  OR U20913 ( .A(n16482), .B(n16483), .Z(n16478) );
  NOR U20914 ( .A(n16484), .B(n16485), .Z(n16402) );
  ANDN U20915 ( .B(n16486), .A(n16487), .Z(n16396) );
  IV U20916 ( .A(n16488), .Z(n16486) );
  XNOR U20917 ( .A(n16389), .B(n16489), .Z(n16395) );
  XNOR U20918 ( .A(n16388), .B(n16390), .Z(n16489) );
  NAND U20919 ( .A(n16490), .B(n16491), .Z(n16390) );
  OR U20920 ( .A(n16492), .B(n16493), .Z(n16491) );
  OR U20921 ( .A(n16494), .B(n16495), .Z(n16490) );
  NAND U20922 ( .A(n16496), .B(n16497), .Z(n16388) );
  OR U20923 ( .A(n16498), .B(n16499), .Z(n16497) );
  OR U20924 ( .A(n16500), .B(n16501), .Z(n16496) );
  ANDN U20925 ( .B(n16502), .A(n16503), .Z(n16389) );
  IV U20926 ( .A(n16504), .Z(n16502) );
  XNOR U20927 ( .A(n16469), .B(n16468), .Z(N28805) );
  XOR U20928 ( .A(n16488), .B(n16487), .Z(n16468) );
  XNOR U20929 ( .A(n16503), .B(n16504), .Z(n16487) );
  XNOR U20930 ( .A(n16498), .B(n16499), .Z(n16504) );
  XNOR U20931 ( .A(n16500), .B(n16501), .Z(n16499) );
  XNOR U20932 ( .A(y[1756]), .B(x[1756]), .Z(n16501) );
  XNOR U20933 ( .A(y[1757]), .B(x[1757]), .Z(n16500) );
  XNOR U20934 ( .A(y[1755]), .B(x[1755]), .Z(n16498) );
  XNOR U20935 ( .A(n16492), .B(n16493), .Z(n16503) );
  XNOR U20936 ( .A(y[1752]), .B(x[1752]), .Z(n16493) );
  XNOR U20937 ( .A(n16494), .B(n16495), .Z(n16492) );
  XNOR U20938 ( .A(y[1753]), .B(x[1753]), .Z(n16495) );
  XNOR U20939 ( .A(y[1754]), .B(x[1754]), .Z(n16494) );
  XNOR U20940 ( .A(n16485), .B(n16484), .Z(n16488) );
  XNOR U20941 ( .A(n16480), .B(n16481), .Z(n16484) );
  XNOR U20942 ( .A(y[1749]), .B(x[1749]), .Z(n16481) );
  XNOR U20943 ( .A(n16482), .B(n16483), .Z(n16480) );
  XNOR U20944 ( .A(y[1750]), .B(x[1750]), .Z(n16483) );
  XNOR U20945 ( .A(y[1751]), .B(x[1751]), .Z(n16482) );
  XNOR U20946 ( .A(n16474), .B(n16475), .Z(n16485) );
  XNOR U20947 ( .A(y[1746]), .B(x[1746]), .Z(n16475) );
  XNOR U20948 ( .A(n16476), .B(n16477), .Z(n16474) );
  XNOR U20949 ( .A(y[1747]), .B(x[1747]), .Z(n16477) );
  XNOR U20950 ( .A(y[1748]), .B(x[1748]), .Z(n16476) );
  XOR U20951 ( .A(n16450), .B(n16451), .Z(n16469) );
  XNOR U20952 ( .A(n16466), .B(n16467), .Z(n16451) );
  XNOR U20953 ( .A(n16461), .B(n16462), .Z(n16467) );
  XNOR U20954 ( .A(n16463), .B(n16464), .Z(n16462) );
  XNOR U20955 ( .A(y[1744]), .B(x[1744]), .Z(n16464) );
  XNOR U20956 ( .A(y[1745]), .B(x[1745]), .Z(n16463) );
  XNOR U20957 ( .A(y[1743]), .B(x[1743]), .Z(n16461) );
  XNOR U20958 ( .A(n16455), .B(n16456), .Z(n16466) );
  XNOR U20959 ( .A(y[1740]), .B(x[1740]), .Z(n16456) );
  XNOR U20960 ( .A(n16457), .B(n16458), .Z(n16455) );
  XNOR U20961 ( .A(y[1741]), .B(x[1741]), .Z(n16458) );
  XNOR U20962 ( .A(y[1742]), .B(x[1742]), .Z(n16457) );
  XOR U20963 ( .A(n16449), .B(n16448), .Z(n16450) );
  XNOR U20964 ( .A(n16444), .B(n16445), .Z(n16448) );
  XNOR U20965 ( .A(y[1737]), .B(x[1737]), .Z(n16445) );
  XNOR U20966 ( .A(n16446), .B(n16447), .Z(n16444) );
  XNOR U20967 ( .A(y[1738]), .B(x[1738]), .Z(n16447) );
  XNOR U20968 ( .A(y[1739]), .B(x[1739]), .Z(n16446) );
  XNOR U20969 ( .A(n16438), .B(n16439), .Z(n16449) );
  XNOR U20970 ( .A(y[1734]), .B(x[1734]), .Z(n16439) );
  XNOR U20971 ( .A(n16440), .B(n16441), .Z(n16438) );
  XNOR U20972 ( .A(y[1735]), .B(x[1735]), .Z(n16441) );
  XNOR U20973 ( .A(y[1736]), .B(x[1736]), .Z(n16440) );
  NAND U20974 ( .A(n16505), .B(n16506), .Z(N28797) );
  NANDN U20975 ( .A(n16507), .B(n16508), .Z(n16506) );
  OR U20976 ( .A(n16509), .B(n16510), .Z(n16508) );
  NAND U20977 ( .A(n16509), .B(n16510), .Z(n16505) );
  XOR U20978 ( .A(n16509), .B(n16511), .Z(N28796) );
  XNOR U20979 ( .A(n16507), .B(n16510), .Z(n16511) );
  AND U20980 ( .A(n16512), .B(n16513), .Z(n16510) );
  NANDN U20981 ( .A(n16514), .B(n16515), .Z(n16513) );
  NANDN U20982 ( .A(n16516), .B(n16517), .Z(n16515) );
  NANDN U20983 ( .A(n16517), .B(n16516), .Z(n16512) );
  NAND U20984 ( .A(n16518), .B(n16519), .Z(n16507) );
  NANDN U20985 ( .A(n16520), .B(n16521), .Z(n16519) );
  OR U20986 ( .A(n16522), .B(n16523), .Z(n16521) );
  NAND U20987 ( .A(n16523), .B(n16522), .Z(n16518) );
  AND U20988 ( .A(n16524), .B(n16525), .Z(n16509) );
  NANDN U20989 ( .A(n16526), .B(n16527), .Z(n16525) );
  NANDN U20990 ( .A(n16528), .B(n16529), .Z(n16527) );
  NANDN U20991 ( .A(n16529), .B(n16528), .Z(n16524) );
  XOR U20992 ( .A(n16523), .B(n16530), .Z(N28795) );
  XOR U20993 ( .A(n16520), .B(n16522), .Z(n16530) );
  XNOR U20994 ( .A(n16516), .B(n16531), .Z(n16522) );
  XNOR U20995 ( .A(n16514), .B(n16517), .Z(n16531) );
  NAND U20996 ( .A(n16532), .B(n16533), .Z(n16517) );
  NAND U20997 ( .A(n16534), .B(n16535), .Z(n16533) );
  OR U20998 ( .A(n16536), .B(n16537), .Z(n16534) );
  NANDN U20999 ( .A(n16538), .B(n16536), .Z(n16532) );
  IV U21000 ( .A(n16537), .Z(n16538) );
  NAND U21001 ( .A(n16539), .B(n16540), .Z(n16514) );
  NAND U21002 ( .A(n16541), .B(n16542), .Z(n16540) );
  NANDN U21003 ( .A(n16543), .B(n16544), .Z(n16541) );
  NANDN U21004 ( .A(n16544), .B(n16543), .Z(n16539) );
  AND U21005 ( .A(n16545), .B(n16546), .Z(n16516) );
  NAND U21006 ( .A(n16547), .B(n16548), .Z(n16546) );
  OR U21007 ( .A(n16549), .B(n16550), .Z(n16547) );
  NANDN U21008 ( .A(n16551), .B(n16549), .Z(n16545) );
  NAND U21009 ( .A(n16552), .B(n16553), .Z(n16520) );
  NANDN U21010 ( .A(n16554), .B(n16555), .Z(n16553) );
  OR U21011 ( .A(n16556), .B(n16557), .Z(n16555) );
  NANDN U21012 ( .A(n16558), .B(n16556), .Z(n16552) );
  IV U21013 ( .A(n16557), .Z(n16558) );
  XNOR U21014 ( .A(n16528), .B(n16559), .Z(n16523) );
  XNOR U21015 ( .A(n16526), .B(n16529), .Z(n16559) );
  NAND U21016 ( .A(n16560), .B(n16561), .Z(n16529) );
  NAND U21017 ( .A(n16562), .B(n16563), .Z(n16561) );
  OR U21018 ( .A(n16564), .B(n16565), .Z(n16562) );
  NANDN U21019 ( .A(n16566), .B(n16564), .Z(n16560) );
  IV U21020 ( .A(n16565), .Z(n16566) );
  NAND U21021 ( .A(n16567), .B(n16568), .Z(n16526) );
  NAND U21022 ( .A(n16569), .B(n16570), .Z(n16568) );
  NANDN U21023 ( .A(n16571), .B(n16572), .Z(n16569) );
  NANDN U21024 ( .A(n16572), .B(n16571), .Z(n16567) );
  AND U21025 ( .A(n16573), .B(n16574), .Z(n16528) );
  NAND U21026 ( .A(n16575), .B(n16576), .Z(n16574) );
  OR U21027 ( .A(n16577), .B(n16578), .Z(n16575) );
  NANDN U21028 ( .A(n16579), .B(n16577), .Z(n16573) );
  XNOR U21029 ( .A(n16554), .B(n16580), .Z(N28794) );
  XOR U21030 ( .A(n16556), .B(n16557), .Z(n16580) );
  XNOR U21031 ( .A(n16570), .B(n16581), .Z(n16557) );
  XOR U21032 ( .A(n16571), .B(n16572), .Z(n16581) );
  XOR U21033 ( .A(n16577), .B(n16582), .Z(n16572) );
  XOR U21034 ( .A(n16576), .B(n16579), .Z(n16582) );
  IV U21035 ( .A(n16578), .Z(n16579) );
  NAND U21036 ( .A(n16583), .B(n16584), .Z(n16578) );
  OR U21037 ( .A(n16585), .B(n16586), .Z(n16584) );
  OR U21038 ( .A(n16587), .B(n16588), .Z(n16583) );
  NAND U21039 ( .A(n16589), .B(n16590), .Z(n16576) );
  OR U21040 ( .A(n16591), .B(n16592), .Z(n16590) );
  OR U21041 ( .A(n16593), .B(n16594), .Z(n16589) );
  NOR U21042 ( .A(n16595), .B(n16596), .Z(n16577) );
  ANDN U21043 ( .B(n16597), .A(n16598), .Z(n16571) );
  XNOR U21044 ( .A(n16564), .B(n16599), .Z(n16570) );
  XNOR U21045 ( .A(n16563), .B(n16565), .Z(n16599) );
  NAND U21046 ( .A(n16600), .B(n16601), .Z(n16565) );
  OR U21047 ( .A(n16602), .B(n16603), .Z(n16601) );
  OR U21048 ( .A(n16604), .B(n16605), .Z(n16600) );
  NAND U21049 ( .A(n16606), .B(n16607), .Z(n16563) );
  OR U21050 ( .A(n16608), .B(n16609), .Z(n16607) );
  OR U21051 ( .A(n16610), .B(n16611), .Z(n16606) );
  ANDN U21052 ( .B(n16612), .A(n16613), .Z(n16564) );
  IV U21053 ( .A(n16614), .Z(n16612) );
  ANDN U21054 ( .B(n16615), .A(n16616), .Z(n16556) );
  XOR U21055 ( .A(n16542), .B(n16617), .Z(n16554) );
  XOR U21056 ( .A(n16543), .B(n16544), .Z(n16617) );
  XOR U21057 ( .A(n16549), .B(n16618), .Z(n16544) );
  XOR U21058 ( .A(n16548), .B(n16551), .Z(n16618) );
  IV U21059 ( .A(n16550), .Z(n16551) );
  NAND U21060 ( .A(n16619), .B(n16620), .Z(n16550) );
  OR U21061 ( .A(n16621), .B(n16622), .Z(n16620) );
  OR U21062 ( .A(n16623), .B(n16624), .Z(n16619) );
  NAND U21063 ( .A(n16625), .B(n16626), .Z(n16548) );
  OR U21064 ( .A(n16627), .B(n16628), .Z(n16626) );
  OR U21065 ( .A(n16629), .B(n16630), .Z(n16625) );
  NOR U21066 ( .A(n16631), .B(n16632), .Z(n16549) );
  ANDN U21067 ( .B(n16633), .A(n16634), .Z(n16543) );
  IV U21068 ( .A(n16635), .Z(n16633) );
  XNOR U21069 ( .A(n16536), .B(n16636), .Z(n16542) );
  XNOR U21070 ( .A(n16535), .B(n16537), .Z(n16636) );
  NAND U21071 ( .A(n16637), .B(n16638), .Z(n16537) );
  OR U21072 ( .A(n16639), .B(n16640), .Z(n16638) );
  OR U21073 ( .A(n16641), .B(n16642), .Z(n16637) );
  NAND U21074 ( .A(n16643), .B(n16644), .Z(n16535) );
  OR U21075 ( .A(n16645), .B(n16646), .Z(n16644) );
  OR U21076 ( .A(n16647), .B(n16648), .Z(n16643) );
  ANDN U21077 ( .B(n16649), .A(n16650), .Z(n16536) );
  IV U21078 ( .A(n16651), .Z(n16649) );
  XNOR U21079 ( .A(n16616), .B(n16615), .Z(N28793) );
  XOR U21080 ( .A(n16635), .B(n16634), .Z(n16615) );
  XNOR U21081 ( .A(n16650), .B(n16651), .Z(n16634) );
  XNOR U21082 ( .A(n16645), .B(n16646), .Z(n16651) );
  XNOR U21083 ( .A(n16647), .B(n16648), .Z(n16646) );
  XNOR U21084 ( .A(y[1732]), .B(x[1732]), .Z(n16648) );
  XNOR U21085 ( .A(y[1733]), .B(x[1733]), .Z(n16647) );
  XNOR U21086 ( .A(y[1731]), .B(x[1731]), .Z(n16645) );
  XNOR U21087 ( .A(n16639), .B(n16640), .Z(n16650) );
  XNOR U21088 ( .A(y[1728]), .B(x[1728]), .Z(n16640) );
  XNOR U21089 ( .A(n16641), .B(n16642), .Z(n16639) );
  XNOR U21090 ( .A(y[1729]), .B(x[1729]), .Z(n16642) );
  XNOR U21091 ( .A(y[1730]), .B(x[1730]), .Z(n16641) );
  XNOR U21092 ( .A(n16632), .B(n16631), .Z(n16635) );
  XNOR U21093 ( .A(n16627), .B(n16628), .Z(n16631) );
  XNOR U21094 ( .A(y[1725]), .B(x[1725]), .Z(n16628) );
  XNOR U21095 ( .A(n16629), .B(n16630), .Z(n16627) );
  XNOR U21096 ( .A(y[1726]), .B(x[1726]), .Z(n16630) );
  XNOR U21097 ( .A(y[1727]), .B(x[1727]), .Z(n16629) );
  XNOR U21098 ( .A(n16621), .B(n16622), .Z(n16632) );
  XNOR U21099 ( .A(y[1722]), .B(x[1722]), .Z(n16622) );
  XNOR U21100 ( .A(n16623), .B(n16624), .Z(n16621) );
  XNOR U21101 ( .A(y[1723]), .B(x[1723]), .Z(n16624) );
  XNOR U21102 ( .A(y[1724]), .B(x[1724]), .Z(n16623) );
  XOR U21103 ( .A(n16597), .B(n16598), .Z(n16616) );
  XNOR U21104 ( .A(n16613), .B(n16614), .Z(n16598) );
  XNOR U21105 ( .A(n16608), .B(n16609), .Z(n16614) );
  XNOR U21106 ( .A(n16610), .B(n16611), .Z(n16609) );
  XNOR U21107 ( .A(y[1720]), .B(x[1720]), .Z(n16611) );
  XNOR U21108 ( .A(y[1721]), .B(x[1721]), .Z(n16610) );
  XNOR U21109 ( .A(y[1719]), .B(x[1719]), .Z(n16608) );
  XNOR U21110 ( .A(n16602), .B(n16603), .Z(n16613) );
  XNOR U21111 ( .A(y[1716]), .B(x[1716]), .Z(n16603) );
  XNOR U21112 ( .A(n16604), .B(n16605), .Z(n16602) );
  XNOR U21113 ( .A(y[1717]), .B(x[1717]), .Z(n16605) );
  XNOR U21114 ( .A(y[1718]), .B(x[1718]), .Z(n16604) );
  XOR U21115 ( .A(n16596), .B(n16595), .Z(n16597) );
  XNOR U21116 ( .A(n16591), .B(n16592), .Z(n16595) );
  XNOR U21117 ( .A(y[1713]), .B(x[1713]), .Z(n16592) );
  XNOR U21118 ( .A(n16593), .B(n16594), .Z(n16591) );
  XNOR U21119 ( .A(y[1714]), .B(x[1714]), .Z(n16594) );
  XNOR U21120 ( .A(y[1715]), .B(x[1715]), .Z(n16593) );
  XNOR U21121 ( .A(n16585), .B(n16586), .Z(n16596) );
  XNOR U21122 ( .A(y[1710]), .B(x[1710]), .Z(n16586) );
  XNOR U21123 ( .A(n16587), .B(n16588), .Z(n16585) );
  XNOR U21124 ( .A(y[1711]), .B(x[1711]), .Z(n16588) );
  XNOR U21125 ( .A(y[1712]), .B(x[1712]), .Z(n16587) );
  NAND U21126 ( .A(n16652), .B(n16653), .Z(N28785) );
  NANDN U21127 ( .A(n16654), .B(n16655), .Z(n16653) );
  OR U21128 ( .A(n16656), .B(n16657), .Z(n16655) );
  NAND U21129 ( .A(n16656), .B(n16657), .Z(n16652) );
  XOR U21130 ( .A(n16656), .B(n16658), .Z(N28784) );
  XNOR U21131 ( .A(n16654), .B(n16657), .Z(n16658) );
  AND U21132 ( .A(n16659), .B(n16660), .Z(n16657) );
  NANDN U21133 ( .A(n16661), .B(n16662), .Z(n16660) );
  NANDN U21134 ( .A(n16663), .B(n16664), .Z(n16662) );
  NANDN U21135 ( .A(n16664), .B(n16663), .Z(n16659) );
  NAND U21136 ( .A(n16665), .B(n16666), .Z(n16654) );
  NANDN U21137 ( .A(n16667), .B(n16668), .Z(n16666) );
  OR U21138 ( .A(n16669), .B(n16670), .Z(n16668) );
  NAND U21139 ( .A(n16670), .B(n16669), .Z(n16665) );
  AND U21140 ( .A(n16671), .B(n16672), .Z(n16656) );
  NANDN U21141 ( .A(n16673), .B(n16674), .Z(n16672) );
  NANDN U21142 ( .A(n16675), .B(n16676), .Z(n16674) );
  NANDN U21143 ( .A(n16676), .B(n16675), .Z(n16671) );
  XOR U21144 ( .A(n16670), .B(n16677), .Z(N28783) );
  XOR U21145 ( .A(n16667), .B(n16669), .Z(n16677) );
  XNOR U21146 ( .A(n16663), .B(n16678), .Z(n16669) );
  XNOR U21147 ( .A(n16661), .B(n16664), .Z(n16678) );
  NAND U21148 ( .A(n16679), .B(n16680), .Z(n16664) );
  NAND U21149 ( .A(n16681), .B(n16682), .Z(n16680) );
  OR U21150 ( .A(n16683), .B(n16684), .Z(n16681) );
  NANDN U21151 ( .A(n16685), .B(n16683), .Z(n16679) );
  IV U21152 ( .A(n16684), .Z(n16685) );
  NAND U21153 ( .A(n16686), .B(n16687), .Z(n16661) );
  NAND U21154 ( .A(n16688), .B(n16689), .Z(n16687) );
  NANDN U21155 ( .A(n16690), .B(n16691), .Z(n16688) );
  NANDN U21156 ( .A(n16691), .B(n16690), .Z(n16686) );
  AND U21157 ( .A(n16692), .B(n16693), .Z(n16663) );
  NAND U21158 ( .A(n16694), .B(n16695), .Z(n16693) );
  OR U21159 ( .A(n16696), .B(n16697), .Z(n16694) );
  NANDN U21160 ( .A(n16698), .B(n16696), .Z(n16692) );
  NAND U21161 ( .A(n16699), .B(n16700), .Z(n16667) );
  NANDN U21162 ( .A(n16701), .B(n16702), .Z(n16700) );
  OR U21163 ( .A(n16703), .B(n16704), .Z(n16702) );
  NANDN U21164 ( .A(n16705), .B(n16703), .Z(n16699) );
  IV U21165 ( .A(n16704), .Z(n16705) );
  XNOR U21166 ( .A(n16675), .B(n16706), .Z(n16670) );
  XNOR U21167 ( .A(n16673), .B(n16676), .Z(n16706) );
  NAND U21168 ( .A(n16707), .B(n16708), .Z(n16676) );
  NAND U21169 ( .A(n16709), .B(n16710), .Z(n16708) );
  OR U21170 ( .A(n16711), .B(n16712), .Z(n16709) );
  NANDN U21171 ( .A(n16713), .B(n16711), .Z(n16707) );
  IV U21172 ( .A(n16712), .Z(n16713) );
  NAND U21173 ( .A(n16714), .B(n16715), .Z(n16673) );
  NAND U21174 ( .A(n16716), .B(n16717), .Z(n16715) );
  NANDN U21175 ( .A(n16718), .B(n16719), .Z(n16716) );
  NANDN U21176 ( .A(n16719), .B(n16718), .Z(n16714) );
  AND U21177 ( .A(n16720), .B(n16721), .Z(n16675) );
  NAND U21178 ( .A(n16722), .B(n16723), .Z(n16721) );
  OR U21179 ( .A(n16724), .B(n16725), .Z(n16722) );
  NANDN U21180 ( .A(n16726), .B(n16724), .Z(n16720) );
  XNOR U21181 ( .A(n16701), .B(n16727), .Z(N28782) );
  XOR U21182 ( .A(n16703), .B(n16704), .Z(n16727) );
  XNOR U21183 ( .A(n16717), .B(n16728), .Z(n16704) );
  XOR U21184 ( .A(n16718), .B(n16719), .Z(n16728) );
  XOR U21185 ( .A(n16724), .B(n16729), .Z(n16719) );
  XOR U21186 ( .A(n16723), .B(n16726), .Z(n16729) );
  IV U21187 ( .A(n16725), .Z(n16726) );
  NAND U21188 ( .A(n16730), .B(n16731), .Z(n16725) );
  OR U21189 ( .A(n16732), .B(n16733), .Z(n16731) );
  OR U21190 ( .A(n16734), .B(n16735), .Z(n16730) );
  NAND U21191 ( .A(n16736), .B(n16737), .Z(n16723) );
  OR U21192 ( .A(n16738), .B(n16739), .Z(n16737) );
  OR U21193 ( .A(n16740), .B(n16741), .Z(n16736) );
  NOR U21194 ( .A(n16742), .B(n16743), .Z(n16724) );
  ANDN U21195 ( .B(n16744), .A(n16745), .Z(n16718) );
  XNOR U21196 ( .A(n16711), .B(n16746), .Z(n16717) );
  XNOR U21197 ( .A(n16710), .B(n16712), .Z(n16746) );
  NAND U21198 ( .A(n16747), .B(n16748), .Z(n16712) );
  OR U21199 ( .A(n16749), .B(n16750), .Z(n16748) );
  OR U21200 ( .A(n16751), .B(n16752), .Z(n16747) );
  NAND U21201 ( .A(n16753), .B(n16754), .Z(n16710) );
  OR U21202 ( .A(n16755), .B(n16756), .Z(n16754) );
  OR U21203 ( .A(n16757), .B(n16758), .Z(n16753) );
  ANDN U21204 ( .B(n16759), .A(n16760), .Z(n16711) );
  IV U21205 ( .A(n16761), .Z(n16759) );
  ANDN U21206 ( .B(n16762), .A(n16763), .Z(n16703) );
  XOR U21207 ( .A(n16689), .B(n16764), .Z(n16701) );
  XOR U21208 ( .A(n16690), .B(n16691), .Z(n16764) );
  XOR U21209 ( .A(n16696), .B(n16765), .Z(n16691) );
  XOR U21210 ( .A(n16695), .B(n16698), .Z(n16765) );
  IV U21211 ( .A(n16697), .Z(n16698) );
  NAND U21212 ( .A(n16766), .B(n16767), .Z(n16697) );
  OR U21213 ( .A(n16768), .B(n16769), .Z(n16767) );
  OR U21214 ( .A(n16770), .B(n16771), .Z(n16766) );
  NAND U21215 ( .A(n16772), .B(n16773), .Z(n16695) );
  OR U21216 ( .A(n16774), .B(n16775), .Z(n16773) );
  OR U21217 ( .A(n16776), .B(n16777), .Z(n16772) );
  NOR U21218 ( .A(n16778), .B(n16779), .Z(n16696) );
  ANDN U21219 ( .B(n16780), .A(n16781), .Z(n16690) );
  IV U21220 ( .A(n16782), .Z(n16780) );
  XNOR U21221 ( .A(n16683), .B(n16783), .Z(n16689) );
  XNOR U21222 ( .A(n16682), .B(n16684), .Z(n16783) );
  NAND U21223 ( .A(n16784), .B(n16785), .Z(n16684) );
  OR U21224 ( .A(n16786), .B(n16787), .Z(n16785) );
  OR U21225 ( .A(n16788), .B(n16789), .Z(n16784) );
  NAND U21226 ( .A(n16790), .B(n16791), .Z(n16682) );
  OR U21227 ( .A(n16792), .B(n16793), .Z(n16791) );
  OR U21228 ( .A(n16794), .B(n16795), .Z(n16790) );
  ANDN U21229 ( .B(n16796), .A(n16797), .Z(n16683) );
  IV U21230 ( .A(n16798), .Z(n16796) );
  XNOR U21231 ( .A(n16763), .B(n16762), .Z(N28781) );
  XOR U21232 ( .A(n16782), .B(n16781), .Z(n16762) );
  XNOR U21233 ( .A(n16797), .B(n16798), .Z(n16781) );
  XNOR U21234 ( .A(n16792), .B(n16793), .Z(n16798) );
  XNOR U21235 ( .A(n16794), .B(n16795), .Z(n16793) );
  XNOR U21236 ( .A(y[1708]), .B(x[1708]), .Z(n16795) );
  XNOR U21237 ( .A(y[1709]), .B(x[1709]), .Z(n16794) );
  XNOR U21238 ( .A(y[1707]), .B(x[1707]), .Z(n16792) );
  XNOR U21239 ( .A(n16786), .B(n16787), .Z(n16797) );
  XNOR U21240 ( .A(y[1704]), .B(x[1704]), .Z(n16787) );
  XNOR U21241 ( .A(n16788), .B(n16789), .Z(n16786) );
  XNOR U21242 ( .A(y[1705]), .B(x[1705]), .Z(n16789) );
  XNOR U21243 ( .A(y[1706]), .B(x[1706]), .Z(n16788) );
  XNOR U21244 ( .A(n16779), .B(n16778), .Z(n16782) );
  XNOR U21245 ( .A(n16774), .B(n16775), .Z(n16778) );
  XNOR U21246 ( .A(y[1701]), .B(x[1701]), .Z(n16775) );
  XNOR U21247 ( .A(n16776), .B(n16777), .Z(n16774) );
  XNOR U21248 ( .A(y[1702]), .B(x[1702]), .Z(n16777) );
  XNOR U21249 ( .A(y[1703]), .B(x[1703]), .Z(n16776) );
  XNOR U21250 ( .A(n16768), .B(n16769), .Z(n16779) );
  XNOR U21251 ( .A(y[1698]), .B(x[1698]), .Z(n16769) );
  XNOR U21252 ( .A(n16770), .B(n16771), .Z(n16768) );
  XNOR U21253 ( .A(y[1699]), .B(x[1699]), .Z(n16771) );
  XNOR U21254 ( .A(y[1700]), .B(x[1700]), .Z(n16770) );
  XOR U21255 ( .A(n16744), .B(n16745), .Z(n16763) );
  XNOR U21256 ( .A(n16760), .B(n16761), .Z(n16745) );
  XNOR U21257 ( .A(n16755), .B(n16756), .Z(n16761) );
  XNOR U21258 ( .A(n16757), .B(n16758), .Z(n16756) );
  XNOR U21259 ( .A(y[1696]), .B(x[1696]), .Z(n16758) );
  XNOR U21260 ( .A(y[1697]), .B(x[1697]), .Z(n16757) );
  XNOR U21261 ( .A(y[1695]), .B(x[1695]), .Z(n16755) );
  XNOR U21262 ( .A(n16749), .B(n16750), .Z(n16760) );
  XNOR U21263 ( .A(y[1692]), .B(x[1692]), .Z(n16750) );
  XNOR U21264 ( .A(n16751), .B(n16752), .Z(n16749) );
  XNOR U21265 ( .A(y[1693]), .B(x[1693]), .Z(n16752) );
  XNOR U21266 ( .A(y[1694]), .B(x[1694]), .Z(n16751) );
  XOR U21267 ( .A(n16743), .B(n16742), .Z(n16744) );
  XNOR U21268 ( .A(n16738), .B(n16739), .Z(n16742) );
  XNOR U21269 ( .A(y[1689]), .B(x[1689]), .Z(n16739) );
  XNOR U21270 ( .A(n16740), .B(n16741), .Z(n16738) );
  XNOR U21271 ( .A(y[1690]), .B(x[1690]), .Z(n16741) );
  XNOR U21272 ( .A(y[1691]), .B(x[1691]), .Z(n16740) );
  XNOR U21273 ( .A(n16732), .B(n16733), .Z(n16743) );
  XNOR U21274 ( .A(y[1686]), .B(x[1686]), .Z(n16733) );
  XNOR U21275 ( .A(n16734), .B(n16735), .Z(n16732) );
  XNOR U21276 ( .A(y[1687]), .B(x[1687]), .Z(n16735) );
  XNOR U21277 ( .A(y[1688]), .B(x[1688]), .Z(n16734) );
  NAND U21278 ( .A(n16799), .B(n16800), .Z(N28773) );
  NANDN U21279 ( .A(n16801), .B(n16802), .Z(n16800) );
  OR U21280 ( .A(n16803), .B(n16804), .Z(n16802) );
  NAND U21281 ( .A(n16803), .B(n16804), .Z(n16799) );
  XOR U21282 ( .A(n16803), .B(n16805), .Z(N28772) );
  XNOR U21283 ( .A(n16801), .B(n16804), .Z(n16805) );
  AND U21284 ( .A(n16806), .B(n16807), .Z(n16804) );
  NANDN U21285 ( .A(n16808), .B(n16809), .Z(n16807) );
  NANDN U21286 ( .A(n16810), .B(n16811), .Z(n16809) );
  NANDN U21287 ( .A(n16811), .B(n16810), .Z(n16806) );
  NAND U21288 ( .A(n16812), .B(n16813), .Z(n16801) );
  NANDN U21289 ( .A(n16814), .B(n16815), .Z(n16813) );
  OR U21290 ( .A(n16816), .B(n16817), .Z(n16815) );
  NAND U21291 ( .A(n16817), .B(n16816), .Z(n16812) );
  AND U21292 ( .A(n16818), .B(n16819), .Z(n16803) );
  NANDN U21293 ( .A(n16820), .B(n16821), .Z(n16819) );
  NANDN U21294 ( .A(n16822), .B(n16823), .Z(n16821) );
  NANDN U21295 ( .A(n16823), .B(n16822), .Z(n16818) );
  XOR U21296 ( .A(n16817), .B(n16824), .Z(N28771) );
  XOR U21297 ( .A(n16814), .B(n16816), .Z(n16824) );
  XNOR U21298 ( .A(n16810), .B(n16825), .Z(n16816) );
  XNOR U21299 ( .A(n16808), .B(n16811), .Z(n16825) );
  NAND U21300 ( .A(n16826), .B(n16827), .Z(n16811) );
  NAND U21301 ( .A(n16828), .B(n16829), .Z(n16827) );
  OR U21302 ( .A(n16830), .B(n16831), .Z(n16828) );
  NANDN U21303 ( .A(n16832), .B(n16830), .Z(n16826) );
  IV U21304 ( .A(n16831), .Z(n16832) );
  NAND U21305 ( .A(n16833), .B(n16834), .Z(n16808) );
  NAND U21306 ( .A(n16835), .B(n16836), .Z(n16834) );
  NANDN U21307 ( .A(n16837), .B(n16838), .Z(n16835) );
  NANDN U21308 ( .A(n16838), .B(n16837), .Z(n16833) );
  AND U21309 ( .A(n16839), .B(n16840), .Z(n16810) );
  NAND U21310 ( .A(n16841), .B(n16842), .Z(n16840) );
  OR U21311 ( .A(n16843), .B(n16844), .Z(n16841) );
  NANDN U21312 ( .A(n16845), .B(n16843), .Z(n16839) );
  NAND U21313 ( .A(n16846), .B(n16847), .Z(n16814) );
  NANDN U21314 ( .A(n16848), .B(n16849), .Z(n16847) );
  OR U21315 ( .A(n16850), .B(n16851), .Z(n16849) );
  NANDN U21316 ( .A(n16852), .B(n16850), .Z(n16846) );
  IV U21317 ( .A(n16851), .Z(n16852) );
  XNOR U21318 ( .A(n16822), .B(n16853), .Z(n16817) );
  XNOR U21319 ( .A(n16820), .B(n16823), .Z(n16853) );
  NAND U21320 ( .A(n16854), .B(n16855), .Z(n16823) );
  NAND U21321 ( .A(n16856), .B(n16857), .Z(n16855) );
  OR U21322 ( .A(n16858), .B(n16859), .Z(n16856) );
  NANDN U21323 ( .A(n16860), .B(n16858), .Z(n16854) );
  IV U21324 ( .A(n16859), .Z(n16860) );
  NAND U21325 ( .A(n16861), .B(n16862), .Z(n16820) );
  NAND U21326 ( .A(n16863), .B(n16864), .Z(n16862) );
  NANDN U21327 ( .A(n16865), .B(n16866), .Z(n16863) );
  NANDN U21328 ( .A(n16866), .B(n16865), .Z(n16861) );
  AND U21329 ( .A(n16867), .B(n16868), .Z(n16822) );
  NAND U21330 ( .A(n16869), .B(n16870), .Z(n16868) );
  OR U21331 ( .A(n16871), .B(n16872), .Z(n16869) );
  NANDN U21332 ( .A(n16873), .B(n16871), .Z(n16867) );
  XNOR U21333 ( .A(n16848), .B(n16874), .Z(N28770) );
  XOR U21334 ( .A(n16850), .B(n16851), .Z(n16874) );
  XNOR U21335 ( .A(n16864), .B(n16875), .Z(n16851) );
  XOR U21336 ( .A(n16865), .B(n16866), .Z(n16875) );
  XOR U21337 ( .A(n16871), .B(n16876), .Z(n16866) );
  XOR U21338 ( .A(n16870), .B(n16873), .Z(n16876) );
  IV U21339 ( .A(n16872), .Z(n16873) );
  NAND U21340 ( .A(n16877), .B(n16878), .Z(n16872) );
  OR U21341 ( .A(n16879), .B(n16880), .Z(n16878) );
  OR U21342 ( .A(n16881), .B(n16882), .Z(n16877) );
  NAND U21343 ( .A(n16883), .B(n16884), .Z(n16870) );
  OR U21344 ( .A(n16885), .B(n16886), .Z(n16884) );
  OR U21345 ( .A(n16887), .B(n16888), .Z(n16883) );
  NOR U21346 ( .A(n16889), .B(n16890), .Z(n16871) );
  ANDN U21347 ( .B(n16891), .A(n16892), .Z(n16865) );
  XNOR U21348 ( .A(n16858), .B(n16893), .Z(n16864) );
  XNOR U21349 ( .A(n16857), .B(n16859), .Z(n16893) );
  NAND U21350 ( .A(n16894), .B(n16895), .Z(n16859) );
  OR U21351 ( .A(n16896), .B(n16897), .Z(n16895) );
  OR U21352 ( .A(n16898), .B(n16899), .Z(n16894) );
  NAND U21353 ( .A(n16900), .B(n16901), .Z(n16857) );
  OR U21354 ( .A(n16902), .B(n16903), .Z(n16901) );
  OR U21355 ( .A(n16904), .B(n16905), .Z(n16900) );
  ANDN U21356 ( .B(n16906), .A(n16907), .Z(n16858) );
  IV U21357 ( .A(n16908), .Z(n16906) );
  ANDN U21358 ( .B(n16909), .A(n16910), .Z(n16850) );
  XOR U21359 ( .A(n16836), .B(n16911), .Z(n16848) );
  XOR U21360 ( .A(n16837), .B(n16838), .Z(n16911) );
  XOR U21361 ( .A(n16843), .B(n16912), .Z(n16838) );
  XOR U21362 ( .A(n16842), .B(n16845), .Z(n16912) );
  IV U21363 ( .A(n16844), .Z(n16845) );
  NAND U21364 ( .A(n16913), .B(n16914), .Z(n16844) );
  OR U21365 ( .A(n16915), .B(n16916), .Z(n16914) );
  OR U21366 ( .A(n16917), .B(n16918), .Z(n16913) );
  NAND U21367 ( .A(n16919), .B(n16920), .Z(n16842) );
  OR U21368 ( .A(n16921), .B(n16922), .Z(n16920) );
  OR U21369 ( .A(n16923), .B(n16924), .Z(n16919) );
  NOR U21370 ( .A(n16925), .B(n16926), .Z(n16843) );
  ANDN U21371 ( .B(n16927), .A(n16928), .Z(n16837) );
  IV U21372 ( .A(n16929), .Z(n16927) );
  XNOR U21373 ( .A(n16830), .B(n16930), .Z(n16836) );
  XNOR U21374 ( .A(n16829), .B(n16831), .Z(n16930) );
  NAND U21375 ( .A(n16931), .B(n16932), .Z(n16831) );
  OR U21376 ( .A(n16933), .B(n16934), .Z(n16932) );
  OR U21377 ( .A(n16935), .B(n16936), .Z(n16931) );
  NAND U21378 ( .A(n16937), .B(n16938), .Z(n16829) );
  OR U21379 ( .A(n16939), .B(n16940), .Z(n16938) );
  OR U21380 ( .A(n16941), .B(n16942), .Z(n16937) );
  ANDN U21381 ( .B(n16943), .A(n16944), .Z(n16830) );
  IV U21382 ( .A(n16945), .Z(n16943) );
  XNOR U21383 ( .A(n16910), .B(n16909), .Z(N28769) );
  XOR U21384 ( .A(n16929), .B(n16928), .Z(n16909) );
  XNOR U21385 ( .A(n16944), .B(n16945), .Z(n16928) );
  XNOR U21386 ( .A(n16939), .B(n16940), .Z(n16945) );
  XNOR U21387 ( .A(n16941), .B(n16942), .Z(n16940) );
  XNOR U21388 ( .A(y[1684]), .B(x[1684]), .Z(n16942) );
  XNOR U21389 ( .A(y[1685]), .B(x[1685]), .Z(n16941) );
  XNOR U21390 ( .A(y[1683]), .B(x[1683]), .Z(n16939) );
  XNOR U21391 ( .A(n16933), .B(n16934), .Z(n16944) );
  XNOR U21392 ( .A(y[1680]), .B(x[1680]), .Z(n16934) );
  XNOR U21393 ( .A(n16935), .B(n16936), .Z(n16933) );
  XNOR U21394 ( .A(y[1681]), .B(x[1681]), .Z(n16936) );
  XNOR U21395 ( .A(y[1682]), .B(x[1682]), .Z(n16935) );
  XNOR U21396 ( .A(n16926), .B(n16925), .Z(n16929) );
  XNOR U21397 ( .A(n16921), .B(n16922), .Z(n16925) );
  XNOR U21398 ( .A(y[1677]), .B(x[1677]), .Z(n16922) );
  XNOR U21399 ( .A(n16923), .B(n16924), .Z(n16921) );
  XNOR U21400 ( .A(y[1678]), .B(x[1678]), .Z(n16924) );
  XNOR U21401 ( .A(y[1679]), .B(x[1679]), .Z(n16923) );
  XNOR U21402 ( .A(n16915), .B(n16916), .Z(n16926) );
  XNOR U21403 ( .A(y[1674]), .B(x[1674]), .Z(n16916) );
  XNOR U21404 ( .A(n16917), .B(n16918), .Z(n16915) );
  XNOR U21405 ( .A(y[1675]), .B(x[1675]), .Z(n16918) );
  XNOR U21406 ( .A(y[1676]), .B(x[1676]), .Z(n16917) );
  XOR U21407 ( .A(n16891), .B(n16892), .Z(n16910) );
  XNOR U21408 ( .A(n16907), .B(n16908), .Z(n16892) );
  XNOR U21409 ( .A(n16902), .B(n16903), .Z(n16908) );
  XNOR U21410 ( .A(n16904), .B(n16905), .Z(n16903) );
  XNOR U21411 ( .A(y[1672]), .B(x[1672]), .Z(n16905) );
  XNOR U21412 ( .A(y[1673]), .B(x[1673]), .Z(n16904) );
  XNOR U21413 ( .A(y[1671]), .B(x[1671]), .Z(n16902) );
  XNOR U21414 ( .A(n16896), .B(n16897), .Z(n16907) );
  XNOR U21415 ( .A(y[1668]), .B(x[1668]), .Z(n16897) );
  XNOR U21416 ( .A(n16898), .B(n16899), .Z(n16896) );
  XNOR U21417 ( .A(y[1669]), .B(x[1669]), .Z(n16899) );
  XNOR U21418 ( .A(y[1670]), .B(x[1670]), .Z(n16898) );
  XOR U21419 ( .A(n16890), .B(n16889), .Z(n16891) );
  XNOR U21420 ( .A(n16885), .B(n16886), .Z(n16889) );
  XNOR U21421 ( .A(y[1665]), .B(x[1665]), .Z(n16886) );
  XNOR U21422 ( .A(n16887), .B(n16888), .Z(n16885) );
  XNOR U21423 ( .A(y[1666]), .B(x[1666]), .Z(n16888) );
  XNOR U21424 ( .A(y[1667]), .B(x[1667]), .Z(n16887) );
  XNOR U21425 ( .A(n16879), .B(n16880), .Z(n16890) );
  XNOR U21426 ( .A(y[1662]), .B(x[1662]), .Z(n16880) );
  XNOR U21427 ( .A(n16881), .B(n16882), .Z(n16879) );
  XNOR U21428 ( .A(y[1663]), .B(x[1663]), .Z(n16882) );
  XNOR U21429 ( .A(y[1664]), .B(x[1664]), .Z(n16881) );
  NAND U21430 ( .A(n16946), .B(n16947), .Z(N28761) );
  NANDN U21431 ( .A(n16948), .B(n16949), .Z(n16947) );
  OR U21432 ( .A(n16950), .B(n16951), .Z(n16949) );
  NAND U21433 ( .A(n16950), .B(n16951), .Z(n16946) );
  XOR U21434 ( .A(n16950), .B(n16952), .Z(N28760) );
  XNOR U21435 ( .A(n16948), .B(n16951), .Z(n16952) );
  AND U21436 ( .A(n16953), .B(n16954), .Z(n16951) );
  NANDN U21437 ( .A(n16955), .B(n16956), .Z(n16954) );
  NANDN U21438 ( .A(n16957), .B(n16958), .Z(n16956) );
  NANDN U21439 ( .A(n16958), .B(n16957), .Z(n16953) );
  NAND U21440 ( .A(n16959), .B(n16960), .Z(n16948) );
  NANDN U21441 ( .A(n16961), .B(n16962), .Z(n16960) );
  OR U21442 ( .A(n16963), .B(n16964), .Z(n16962) );
  NAND U21443 ( .A(n16964), .B(n16963), .Z(n16959) );
  AND U21444 ( .A(n16965), .B(n16966), .Z(n16950) );
  NANDN U21445 ( .A(n16967), .B(n16968), .Z(n16966) );
  NANDN U21446 ( .A(n16969), .B(n16970), .Z(n16968) );
  NANDN U21447 ( .A(n16970), .B(n16969), .Z(n16965) );
  XOR U21448 ( .A(n16964), .B(n16971), .Z(N28759) );
  XOR U21449 ( .A(n16961), .B(n16963), .Z(n16971) );
  XNOR U21450 ( .A(n16957), .B(n16972), .Z(n16963) );
  XNOR U21451 ( .A(n16955), .B(n16958), .Z(n16972) );
  NAND U21452 ( .A(n16973), .B(n16974), .Z(n16958) );
  NAND U21453 ( .A(n16975), .B(n16976), .Z(n16974) );
  OR U21454 ( .A(n16977), .B(n16978), .Z(n16975) );
  NANDN U21455 ( .A(n16979), .B(n16977), .Z(n16973) );
  IV U21456 ( .A(n16978), .Z(n16979) );
  NAND U21457 ( .A(n16980), .B(n16981), .Z(n16955) );
  NAND U21458 ( .A(n16982), .B(n16983), .Z(n16981) );
  NANDN U21459 ( .A(n16984), .B(n16985), .Z(n16982) );
  NANDN U21460 ( .A(n16985), .B(n16984), .Z(n16980) );
  AND U21461 ( .A(n16986), .B(n16987), .Z(n16957) );
  NAND U21462 ( .A(n16988), .B(n16989), .Z(n16987) );
  OR U21463 ( .A(n16990), .B(n16991), .Z(n16988) );
  NANDN U21464 ( .A(n16992), .B(n16990), .Z(n16986) );
  NAND U21465 ( .A(n16993), .B(n16994), .Z(n16961) );
  NANDN U21466 ( .A(n16995), .B(n16996), .Z(n16994) );
  OR U21467 ( .A(n16997), .B(n16998), .Z(n16996) );
  NANDN U21468 ( .A(n16999), .B(n16997), .Z(n16993) );
  IV U21469 ( .A(n16998), .Z(n16999) );
  XNOR U21470 ( .A(n16969), .B(n17000), .Z(n16964) );
  XNOR U21471 ( .A(n16967), .B(n16970), .Z(n17000) );
  NAND U21472 ( .A(n17001), .B(n17002), .Z(n16970) );
  NAND U21473 ( .A(n17003), .B(n17004), .Z(n17002) );
  OR U21474 ( .A(n17005), .B(n17006), .Z(n17003) );
  NANDN U21475 ( .A(n17007), .B(n17005), .Z(n17001) );
  IV U21476 ( .A(n17006), .Z(n17007) );
  NAND U21477 ( .A(n17008), .B(n17009), .Z(n16967) );
  NAND U21478 ( .A(n17010), .B(n17011), .Z(n17009) );
  NANDN U21479 ( .A(n17012), .B(n17013), .Z(n17010) );
  NANDN U21480 ( .A(n17013), .B(n17012), .Z(n17008) );
  AND U21481 ( .A(n17014), .B(n17015), .Z(n16969) );
  NAND U21482 ( .A(n17016), .B(n17017), .Z(n17015) );
  OR U21483 ( .A(n17018), .B(n17019), .Z(n17016) );
  NANDN U21484 ( .A(n17020), .B(n17018), .Z(n17014) );
  XNOR U21485 ( .A(n16995), .B(n17021), .Z(N28758) );
  XOR U21486 ( .A(n16997), .B(n16998), .Z(n17021) );
  XNOR U21487 ( .A(n17011), .B(n17022), .Z(n16998) );
  XOR U21488 ( .A(n17012), .B(n17013), .Z(n17022) );
  XOR U21489 ( .A(n17018), .B(n17023), .Z(n17013) );
  XOR U21490 ( .A(n17017), .B(n17020), .Z(n17023) );
  IV U21491 ( .A(n17019), .Z(n17020) );
  NAND U21492 ( .A(n17024), .B(n17025), .Z(n17019) );
  OR U21493 ( .A(n17026), .B(n17027), .Z(n17025) );
  OR U21494 ( .A(n17028), .B(n17029), .Z(n17024) );
  NAND U21495 ( .A(n17030), .B(n17031), .Z(n17017) );
  OR U21496 ( .A(n17032), .B(n17033), .Z(n17031) );
  OR U21497 ( .A(n17034), .B(n17035), .Z(n17030) );
  NOR U21498 ( .A(n17036), .B(n17037), .Z(n17018) );
  ANDN U21499 ( .B(n17038), .A(n17039), .Z(n17012) );
  XNOR U21500 ( .A(n17005), .B(n17040), .Z(n17011) );
  XNOR U21501 ( .A(n17004), .B(n17006), .Z(n17040) );
  NAND U21502 ( .A(n17041), .B(n17042), .Z(n17006) );
  OR U21503 ( .A(n17043), .B(n17044), .Z(n17042) );
  OR U21504 ( .A(n17045), .B(n17046), .Z(n17041) );
  NAND U21505 ( .A(n17047), .B(n17048), .Z(n17004) );
  OR U21506 ( .A(n17049), .B(n17050), .Z(n17048) );
  OR U21507 ( .A(n17051), .B(n17052), .Z(n17047) );
  ANDN U21508 ( .B(n17053), .A(n17054), .Z(n17005) );
  IV U21509 ( .A(n17055), .Z(n17053) );
  ANDN U21510 ( .B(n17056), .A(n17057), .Z(n16997) );
  XOR U21511 ( .A(n16983), .B(n17058), .Z(n16995) );
  XOR U21512 ( .A(n16984), .B(n16985), .Z(n17058) );
  XOR U21513 ( .A(n16990), .B(n17059), .Z(n16985) );
  XOR U21514 ( .A(n16989), .B(n16992), .Z(n17059) );
  IV U21515 ( .A(n16991), .Z(n16992) );
  NAND U21516 ( .A(n17060), .B(n17061), .Z(n16991) );
  OR U21517 ( .A(n17062), .B(n17063), .Z(n17061) );
  OR U21518 ( .A(n17064), .B(n17065), .Z(n17060) );
  NAND U21519 ( .A(n17066), .B(n17067), .Z(n16989) );
  OR U21520 ( .A(n17068), .B(n17069), .Z(n17067) );
  OR U21521 ( .A(n17070), .B(n17071), .Z(n17066) );
  NOR U21522 ( .A(n17072), .B(n17073), .Z(n16990) );
  ANDN U21523 ( .B(n17074), .A(n17075), .Z(n16984) );
  IV U21524 ( .A(n17076), .Z(n17074) );
  XNOR U21525 ( .A(n16977), .B(n17077), .Z(n16983) );
  XNOR U21526 ( .A(n16976), .B(n16978), .Z(n17077) );
  NAND U21527 ( .A(n17078), .B(n17079), .Z(n16978) );
  OR U21528 ( .A(n17080), .B(n17081), .Z(n17079) );
  OR U21529 ( .A(n17082), .B(n17083), .Z(n17078) );
  NAND U21530 ( .A(n17084), .B(n17085), .Z(n16976) );
  OR U21531 ( .A(n17086), .B(n17087), .Z(n17085) );
  OR U21532 ( .A(n17088), .B(n17089), .Z(n17084) );
  ANDN U21533 ( .B(n17090), .A(n17091), .Z(n16977) );
  IV U21534 ( .A(n17092), .Z(n17090) );
  XNOR U21535 ( .A(n17057), .B(n17056), .Z(N28757) );
  XOR U21536 ( .A(n17076), .B(n17075), .Z(n17056) );
  XNOR U21537 ( .A(n17091), .B(n17092), .Z(n17075) );
  XNOR U21538 ( .A(n17086), .B(n17087), .Z(n17092) );
  XNOR U21539 ( .A(n17088), .B(n17089), .Z(n17087) );
  XNOR U21540 ( .A(y[1660]), .B(x[1660]), .Z(n17089) );
  XNOR U21541 ( .A(y[1661]), .B(x[1661]), .Z(n17088) );
  XNOR U21542 ( .A(y[1659]), .B(x[1659]), .Z(n17086) );
  XNOR U21543 ( .A(n17080), .B(n17081), .Z(n17091) );
  XNOR U21544 ( .A(y[1656]), .B(x[1656]), .Z(n17081) );
  XNOR U21545 ( .A(n17082), .B(n17083), .Z(n17080) );
  XNOR U21546 ( .A(y[1657]), .B(x[1657]), .Z(n17083) );
  XNOR U21547 ( .A(y[1658]), .B(x[1658]), .Z(n17082) );
  XNOR U21548 ( .A(n17073), .B(n17072), .Z(n17076) );
  XNOR U21549 ( .A(n17068), .B(n17069), .Z(n17072) );
  XNOR U21550 ( .A(y[1653]), .B(x[1653]), .Z(n17069) );
  XNOR U21551 ( .A(n17070), .B(n17071), .Z(n17068) );
  XNOR U21552 ( .A(y[1654]), .B(x[1654]), .Z(n17071) );
  XNOR U21553 ( .A(y[1655]), .B(x[1655]), .Z(n17070) );
  XNOR U21554 ( .A(n17062), .B(n17063), .Z(n17073) );
  XNOR U21555 ( .A(y[1650]), .B(x[1650]), .Z(n17063) );
  XNOR U21556 ( .A(n17064), .B(n17065), .Z(n17062) );
  XNOR U21557 ( .A(y[1651]), .B(x[1651]), .Z(n17065) );
  XNOR U21558 ( .A(y[1652]), .B(x[1652]), .Z(n17064) );
  XOR U21559 ( .A(n17038), .B(n17039), .Z(n17057) );
  XNOR U21560 ( .A(n17054), .B(n17055), .Z(n17039) );
  XNOR U21561 ( .A(n17049), .B(n17050), .Z(n17055) );
  XNOR U21562 ( .A(n17051), .B(n17052), .Z(n17050) );
  XNOR U21563 ( .A(y[1648]), .B(x[1648]), .Z(n17052) );
  XNOR U21564 ( .A(y[1649]), .B(x[1649]), .Z(n17051) );
  XNOR U21565 ( .A(y[1647]), .B(x[1647]), .Z(n17049) );
  XNOR U21566 ( .A(n17043), .B(n17044), .Z(n17054) );
  XNOR U21567 ( .A(y[1644]), .B(x[1644]), .Z(n17044) );
  XNOR U21568 ( .A(n17045), .B(n17046), .Z(n17043) );
  XNOR U21569 ( .A(y[1645]), .B(x[1645]), .Z(n17046) );
  XNOR U21570 ( .A(y[1646]), .B(x[1646]), .Z(n17045) );
  XOR U21571 ( .A(n17037), .B(n17036), .Z(n17038) );
  XNOR U21572 ( .A(n17032), .B(n17033), .Z(n17036) );
  XNOR U21573 ( .A(y[1641]), .B(x[1641]), .Z(n17033) );
  XNOR U21574 ( .A(n17034), .B(n17035), .Z(n17032) );
  XNOR U21575 ( .A(y[1642]), .B(x[1642]), .Z(n17035) );
  XNOR U21576 ( .A(y[1643]), .B(x[1643]), .Z(n17034) );
  XNOR U21577 ( .A(n17026), .B(n17027), .Z(n17037) );
  XNOR U21578 ( .A(y[1638]), .B(x[1638]), .Z(n17027) );
  XNOR U21579 ( .A(n17028), .B(n17029), .Z(n17026) );
  XNOR U21580 ( .A(y[1639]), .B(x[1639]), .Z(n17029) );
  XNOR U21581 ( .A(y[1640]), .B(x[1640]), .Z(n17028) );
  NAND U21582 ( .A(n17093), .B(n17094), .Z(N28749) );
  NANDN U21583 ( .A(n17095), .B(n17096), .Z(n17094) );
  OR U21584 ( .A(n17097), .B(n17098), .Z(n17096) );
  NAND U21585 ( .A(n17097), .B(n17098), .Z(n17093) );
  XOR U21586 ( .A(n17097), .B(n17099), .Z(N28748) );
  XNOR U21587 ( .A(n17095), .B(n17098), .Z(n17099) );
  AND U21588 ( .A(n17100), .B(n17101), .Z(n17098) );
  NANDN U21589 ( .A(n17102), .B(n17103), .Z(n17101) );
  NANDN U21590 ( .A(n17104), .B(n17105), .Z(n17103) );
  NANDN U21591 ( .A(n17105), .B(n17104), .Z(n17100) );
  NAND U21592 ( .A(n17106), .B(n17107), .Z(n17095) );
  NANDN U21593 ( .A(n17108), .B(n17109), .Z(n17107) );
  OR U21594 ( .A(n17110), .B(n17111), .Z(n17109) );
  NAND U21595 ( .A(n17111), .B(n17110), .Z(n17106) );
  AND U21596 ( .A(n17112), .B(n17113), .Z(n17097) );
  NANDN U21597 ( .A(n17114), .B(n17115), .Z(n17113) );
  NANDN U21598 ( .A(n17116), .B(n17117), .Z(n17115) );
  NANDN U21599 ( .A(n17117), .B(n17116), .Z(n17112) );
  XOR U21600 ( .A(n17111), .B(n17118), .Z(N28747) );
  XOR U21601 ( .A(n17108), .B(n17110), .Z(n17118) );
  XNOR U21602 ( .A(n17104), .B(n17119), .Z(n17110) );
  XNOR U21603 ( .A(n17102), .B(n17105), .Z(n17119) );
  NAND U21604 ( .A(n17120), .B(n17121), .Z(n17105) );
  NAND U21605 ( .A(n17122), .B(n17123), .Z(n17121) );
  OR U21606 ( .A(n17124), .B(n17125), .Z(n17122) );
  NANDN U21607 ( .A(n17126), .B(n17124), .Z(n17120) );
  IV U21608 ( .A(n17125), .Z(n17126) );
  NAND U21609 ( .A(n17127), .B(n17128), .Z(n17102) );
  NAND U21610 ( .A(n17129), .B(n17130), .Z(n17128) );
  NANDN U21611 ( .A(n17131), .B(n17132), .Z(n17129) );
  NANDN U21612 ( .A(n17132), .B(n17131), .Z(n17127) );
  AND U21613 ( .A(n17133), .B(n17134), .Z(n17104) );
  NAND U21614 ( .A(n17135), .B(n17136), .Z(n17134) );
  OR U21615 ( .A(n17137), .B(n17138), .Z(n17135) );
  NANDN U21616 ( .A(n17139), .B(n17137), .Z(n17133) );
  NAND U21617 ( .A(n17140), .B(n17141), .Z(n17108) );
  NANDN U21618 ( .A(n17142), .B(n17143), .Z(n17141) );
  OR U21619 ( .A(n17144), .B(n17145), .Z(n17143) );
  NANDN U21620 ( .A(n17146), .B(n17144), .Z(n17140) );
  IV U21621 ( .A(n17145), .Z(n17146) );
  XNOR U21622 ( .A(n17116), .B(n17147), .Z(n17111) );
  XNOR U21623 ( .A(n17114), .B(n17117), .Z(n17147) );
  NAND U21624 ( .A(n17148), .B(n17149), .Z(n17117) );
  NAND U21625 ( .A(n17150), .B(n17151), .Z(n17149) );
  OR U21626 ( .A(n17152), .B(n17153), .Z(n17150) );
  NANDN U21627 ( .A(n17154), .B(n17152), .Z(n17148) );
  IV U21628 ( .A(n17153), .Z(n17154) );
  NAND U21629 ( .A(n17155), .B(n17156), .Z(n17114) );
  NAND U21630 ( .A(n17157), .B(n17158), .Z(n17156) );
  NANDN U21631 ( .A(n17159), .B(n17160), .Z(n17157) );
  NANDN U21632 ( .A(n17160), .B(n17159), .Z(n17155) );
  AND U21633 ( .A(n17161), .B(n17162), .Z(n17116) );
  NAND U21634 ( .A(n17163), .B(n17164), .Z(n17162) );
  OR U21635 ( .A(n17165), .B(n17166), .Z(n17163) );
  NANDN U21636 ( .A(n17167), .B(n17165), .Z(n17161) );
  XNOR U21637 ( .A(n17142), .B(n17168), .Z(N28746) );
  XOR U21638 ( .A(n17144), .B(n17145), .Z(n17168) );
  XNOR U21639 ( .A(n17158), .B(n17169), .Z(n17145) );
  XOR U21640 ( .A(n17159), .B(n17160), .Z(n17169) );
  XOR U21641 ( .A(n17165), .B(n17170), .Z(n17160) );
  XOR U21642 ( .A(n17164), .B(n17167), .Z(n17170) );
  IV U21643 ( .A(n17166), .Z(n17167) );
  NAND U21644 ( .A(n17171), .B(n17172), .Z(n17166) );
  OR U21645 ( .A(n17173), .B(n17174), .Z(n17172) );
  OR U21646 ( .A(n17175), .B(n17176), .Z(n17171) );
  NAND U21647 ( .A(n17177), .B(n17178), .Z(n17164) );
  OR U21648 ( .A(n17179), .B(n17180), .Z(n17178) );
  OR U21649 ( .A(n17181), .B(n17182), .Z(n17177) );
  NOR U21650 ( .A(n17183), .B(n17184), .Z(n17165) );
  ANDN U21651 ( .B(n17185), .A(n17186), .Z(n17159) );
  XNOR U21652 ( .A(n17152), .B(n17187), .Z(n17158) );
  XNOR U21653 ( .A(n17151), .B(n17153), .Z(n17187) );
  NAND U21654 ( .A(n17188), .B(n17189), .Z(n17153) );
  OR U21655 ( .A(n17190), .B(n17191), .Z(n17189) );
  OR U21656 ( .A(n17192), .B(n17193), .Z(n17188) );
  NAND U21657 ( .A(n17194), .B(n17195), .Z(n17151) );
  OR U21658 ( .A(n17196), .B(n17197), .Z(n17195) );
  OR U21659 ( .A(n17198), .B(n17199), .Z(n17194) );
  ANDN U21660 ( .B(n17200), .A(n17201), .Z(n17152) );
  IV U21661 ( .A(n17202), .Z(n17200) );
  ANDN U21662 ( .B(n17203), .A(n17204), .Z(n17144) );
  XOR U21663 ( .A(n17130), .B(n17205), .Z(n17142) );
  XOR U21664 ( .A(n17131), .B(n17132), .Z(n17205) );
  XOR U21665 ( .A(n17137), .B(n17206), .Z(n17132) );
  XOR U21666 ( .A(n17136), .B(n17139), .Z(n17206) );
  IV U21667 ( .A(n17138), .Z(n17139) );
  NAND U21668 ( .A(n17207), .B(n17208), .Z(n17138) );
  OR U21669 ( .A(n17209), .B(n17210), .Z(n17208) );
  OR U21670 ( .A(n17211), .B(n17212), .Z(n17207) );
  NAND U21671 ( .A(n17213), .B(n17214), .Z(n17136) );
  OR U21672 ( .A(n17215), .B(n17216), .Z(n17214) );
  OR U21673 ( .A(n17217), .B(n17218), .Z(n17213) );
  NOR U21674 ( .A(n17219), .B(n17220), .Z(n17137) );
  ANDN U21675 ( .B(n17221), .A(n17222), .Z(n17131) );
  IV U21676 ( .A(n17223), .Z(n17221) );
  XNOR U21677 ( .A(n17124), .B(n17224), .Z(n17130) );
  XNOR U21678 ( .A(n17123), .B(n17125), .Z(n17224) );
  NAND U21679 ( .A(n17225), .B(n17226), .Z(n17125) );
  OR U21680 ( .A(n17227), .B(n17228), .Z(n17226) );
  OR U21681 ( .A(n17229), .B(n17230), .Z(n17225) );
  NAND U21682 ( .A(n17231), .B(n17232), .Z(n17123) );
  OR U21683 ( .A(n17233), .B(n17234), .Z(n17232) );
  OR U21684 ( .A(n17235), .B(n17236), .Z(n17231) );
  ANDN U21685 ( .B(n17237), .A(n17238), .Z(n17124) );
  IV U21686 ( .A(n17239), .Z(n17237) );
  XNOR U21687 ( .A(n17204), .B(n17203), .Z(N28745) );
  XOR U21688 ( .A(n17223), .B(n17222), .Z(n17203) );
  XNOR U21689 ( .A(n17238), .B(n17239), .Z(n17222) );
  XNOR U21690 ( .A(n17233), .B(n17234), .Z(n17239) );
  XNOR U21691 ( .A(n17235), .B(n17236), .Z(n17234) );
  XNOR U21692 ( .A(y[1636]), .B(x[1636]), .Z(n17236) );
  XNOR U21693 ( .A(y[1637]), .B(x[1637]), .Z(n17235) );
  XNOR U21694 ( .A(y[1635]), .B(x[1635]), .Z(n17233) );
  XNOR U21695 ( .A(n17227), .B(n17228), .Z(n17238) );
  XNOR U21696 ( .A(y[1632]), .B(x[1632]), .Z(n17228) );
  XNOR U21697 ( .A(n17229), .B(n17230), .Z(n17227) );
  XNOR U21698 ( .A(y[1633]), .B(x[1633]), .Z(n17230) );
  XNOR U21699 ( .A(y[1634]), .B(x[1634]), .Z(n17229) );
  XNOR U21700 ( .A(n17220), .B(n17219), .Z(n17223) );
  XNOR U21701 ( .A(n17215), .B(n17216), .Z(n17219) );
  XNOR U21702 ( .A(y[1629]), .B(x[1629]), .Z(n17216) );
  XNOR U21703 ( .A(n17217), .B(n17218), .Z(n17215) );
  XNOR U21704 ( .A(y[1630]), .B(x[1630]), .Z(n17218) );
  XNOR U21705 ( .A(y[1631]), .B(x[1631]), .Z(n17217) );
  XNOR U21706 ( .A(n17209), .B(n17210), .Z(n17220) );
  XNOR U21707 ( .A(y[1626]), .B(x[1626]), .Z(n17210) );
  XNOR U21708 ( .A(n17211), .B(n17212), .Z(n17209) );
  XNOR U21709 ( .A(y[1627]), .B(x[1627]), .Z(n17212) );
  XNOR U21710 ( .A(y[1628]), .B(x[1628]), .Z(n17211) );
  XOR U21711 ( .A(n17185), .B(n17186), .Z(n17204) );
  XNOR U21712 ( .A(n17201), .B(n17202), .Z(n17186) );
  XNOR U21713 ( .A(n17196), .B(n17197), .Z(n17202) );
  XNOR U21714 ( .A(n17198), .B(n17199), .Z(n17197) );
  XNOR U21715 ( .A(y[1624]), .B(x[1624]), .Z(n17199) );
  XNOR U21716 ( .A(y[1625]), .B(x[1625]), .Z(n17198) );
  XNOR U21717 ( .A(y[1623]), .B(x[1623]), .Z(n17196) );
  XNOR U21718 ( .A(n17190), .B(n17191), .Z(n17201) );
  XNOR U21719 ( .A(y[1620]), .B(x[1620]), .Z(n17191) );
  XNOR U21720 ( .A(n17192), .B(n17193), .Z(n17190) );
  XNOR U21721 ( .A(y[1621]), .B(x[1621]), .Z(n17193) );
  XNOR U21722 ( .A(y[1622]), .B(x[1622]), .Z(n17192) );
  XOR U21723 ( .A(n17184), .B(n17183), .Z(n17185) );
  XNOR U21724 ( .A(n17179), .B(n17180), .Z(n17183) );
  XNOR U21725 ( .A(y[1617]), .B(x[1617]), .Z(n17180) );
  XNOR U21726 ( .A(n17181), .B(n17182), .Z(n17179) );
  XNOR U21727 ( .A(y[1618]), .B(x[1618]), .Z(n17182) );
  XNOR U21728 ( .A(y[1619]), .B(x[1619]), .Z(n17181) );
  XNOR U21729 ( .A(n17173), .B(n17174), .Z(n17184) );
  XNOR U21730 ( .A(y[1614]), .B(x[1614]), .Z(n17174) );
  XNOR U21731 ( .A(n17175), .B(n17176), .Z(n17173) );
  XNOR U21732 ( .A(y[1615]), .B(x[1615]), .Z(n17176) );
  XNOR U21733 ( .A(y[1616]), .B(x[1616]), .Z(n17175) );
  NAND U21734 ( .A(n17240), .B(n17241), .Z(N28737) );
  NANDN U21735 ( .A(n17242), .B(n17243), .Z(n17241) );
  OR U21736 ( .A(n17244), .B(n17245), .Z(n17243) );
  NAND U21737 ( .A(n17244), .B(n17245), .Z(n17240) );
  XOR U21738 ( .A(n17244), .B(n17246), .Z(N28736) );
  XNOR U21739 ( .A(n17242), .B(n17245), .Z(n17246) );
  AND U21740 ( .A(n17247), .B(n17248), .Z(n17245) );
  NANDN U21741 ( .A(n17249), .B(n17250), .Z(n17248) );
  NANDN U21742 ( .A(n17251), .B(n17252), .Z(n17250) );
  NANDN U21743 ( .A(n17252), .B(n17251), .Z(n17247) );
  NAND U21744 ( .A(n17253), .B(n17254), .Z(n17242) );
  NANDN U21745 ( .A(n17255), .B(n17256), .Z(n17254) );
  OR U21746 ( .A(n17257), .B(n17258), .Z(n17256) );
  NAND U21747 ( .A(n17258), .B(n17257), .Z(n17253) );
  AND U21748 ( .A(n17259), .B(n17260), .Z(n17244) );
  NANDN U21749 ( .A(n17261), .B(n17262), .Z(n17260) );
  NANDN U21750 ( .A(n17263), .B(n17264), .Z(n17262) );
  NANDN U21751 ( .A(n17264), .B(n17263), .Z(n17259) );
  XOR U21752 ( .A(n17258), .B(n17265), .Z(N28735) );
  XOR U21753 ( .A(n17255), .B(n17257), .Z(n17265) );
  XNOR U21754 ( .A(n17251), .B(n17266), .Z(n17257) );
  XNOR U21755 ( .A(n17249), .B(n17252), .Z(n17266) );
  NAND U21756 ( .A(n17267), .B(n17268), .Z(n17252) );
  NAND U21757 ( .A(n17269), .B(n17270), .Z(n17268) );
  OR U21758 ( .A(n17271), .B(n17272), .Z(n17269) );
  NANDN U21759 ( .A(n17273), .B(n17271), .Z(n17267) );
  IV U21760 ( .A(n17272), .Z(n17273) );
  NAND U21761 ( .A(n17274), .B(n17275), .Z(n17249) );
  NAND U21762 ( .A(n17276), .B(n17277), .Z(n17275) );
  NANDN U21763 ( .A(n17278), .B(n17279), .Z(n17276) );
  NANDN U21764 ( .A(n17279), .B(n17278), .Z(n17274) );
  AND U21765 ( .A(n17280), .B(n17281), .Z(n17251) );
  NAND U21766 ( .A(n17282), .B(n17283), .Z(n17281) );
  OR U21767 ( .A(n17284), .B(n17285), .Z(n17282) );
  NANDN U21768 ( .A(n17286), .B(n17284), .Z(n17280) );
  NAND U21769 ( .A(n17287), .B(n17288), .Z(n17255) );
  NANDN U21770 ( .A(n17289), .B(n17290), .Z(n17288) );
  OR U21771 ( .A(n17291), .B(n17292), .Z(n17290) );
  NANDN U21772 ( .A(n17293), .B(n17291), .Z(n17287) );
  IV U21773 ( .A(n17292), .Z(n17293) );
  XNOR U21774 ( .A(n17263), .B(n17294), .Z(n17258) );
  XNOR U21775 ( .A(n17261), .B(n17264), .Z(n17294) );
  NAND U21776 ( .A(n17295), .B(n17296), .Z(n17264) );
  NAND U21777 ( .A(n17297), .B(n17298), .Z(n17296) );
  OR U21778 ( .A(n17299), .B(n17300), .Z(n17297) );
  NANDN U21779 ( .A(n17301), .B(n17299), .Z(n17295) );
  IV U21780 ( .A(n17300), .Z(n17301) );
  NAND U21781 ( .A(n17302), .B(n17303), .Z(n17261) );
  NAND U21782 ( .A(n17304), .B(n17305), .Z(n17303) );
  NANDN U21783 ( .A(n17306), .B(n17307), .Z(n17304) );
  NANDN U21784 ( .A(n17307), .B(n17306), .Z(n17302) );
  AND U21785 ( .A(n17308), .B(n17309), .Z(n17263) );
  NAND U21786 ( .A(n17310), .B(n17311), .Z(n17309) );
  OR U21787 ( .A(n17312), .B(n17313), .Z(n17310) );
  NANDN U21788 ( .A(n17314), .B(n17312), .Z(n17308) );
  XNOR U21789 ( .A(n17289), .B(n17315), .Z(N28734) );
  XOR U21790 ( .A(n17291), .B(n17292), .Z(n17315) );
  XNOR U21791 ( .A(n17305), .B(n17316), .Z(n17292) );
  XOR U21792 ( .A(n17306), .B(n17307), .Z(n17316) );
  XOR U21793 ( .A(n17312), .B(n17317), .Z(n17307) );
  XOR U21794 ( .A(n17311), .B(n17314), .Z(n17317) );
  IV U21795 ( .A(n17313), .Z(n17314) );
  NAND U21796 ( .A(n17318), .B(n17319), .Z(n17313) );
  OR U21797 ( .A(n17320), .B(n17321), .Z(n17319) );
  OR U21798 ( .A(n17322), .B(n17323), .Z(n17318) );
  NAND U21799 ( .A(n17324), .B(n17325), .Z(n17311) );
  OR U21800 ( .A(n17326), .B(n17327), .Z(n17325) );
  OR U21801 ( .A(n17328), .B(n17329), .Z(n17324) );
  NOR U21802 ( .A(n17330), .B(n17331), .Z(n17312) );
  ANDN U21803 ( .B(n17332), .A(n17333), .Z(n17306) );
  XNOR U21804 ( .A(n17299), .B(n17334), .Z(n17305) );
  XNOR U21805 ( .A(n17298), .B(n17300), .Z(n17334) );
  NAND U21806 ( .A(n17335), .B(n17336), .Z(n17300) );
  OR U21807 ( .A(n17337), .B(n17338), .Z(n17336) );
  OR U21808 ( .A(n17339), .B(n17340), .Z(n17335) );
  NAND U21809 ( .A(n17341), .B(n17342), .Z(n17298) );
  OR U21810 ( .A(n17343), .B(n17344), .Z(n17342) );
  OR U21811 ( .A(n17345), .B(n17346), .Z(n17341) );
  ANDN U21812 ( .B(n17347), .A(n17348), .Z(n17299) );
  IV U21813 ( .A(n17349), .Z(n17347) );
  ANDN U21814 ( .B(n17350), .A(n17351), .Z(n17291) );
  XOR U21815 ( .A(n17277), .B(n17352), .Z(n17289) );
  XOR U21816 ( .A(n17278), .B(n17279), .Z(n17352) );
  XOR U21817 ( .A(n17284), .B(n17353), .Z(n17279) );
  XOR U21818 ( .A(n17283), .B(n17286), .Z(n17353) );
  IV U21819 ( .A(n17285), .Z(n17286) );
  NAND U21820 ( .A(n17354), .B(n17355), .Z(n17285) );
  OR U21821 ( .A(n17356), .B(n17357), .Z(n17355) );
  OR U21822 ( .A(n17358), .B(n17359), .Z(n17354) );
  NAND U21823 ( .A(n17360), .B(n17361), .Z(n17283) );
  OR U21824 ( .A(n17362), .B(n17363), .Z(n17361) );
  OR U21825 ( .A(n17364), .B(n17365), .Z(n17360) );
  NOR U21826 ( .A(n17366), .B(n17367), .Z(n17284) );
  ANDN U21827 ( .B(n17368), .A(n17369), .Z(n17278) );
  IV U21828 ( .A(n17370), .Z(n17368) );
  XNOR U21829 ( .A(n17271), .B(n17371), .Z(n17277) );
  XNOR U21830 ( .A(n17270), .B(n17272), .Z(n17371) );
  NAND U21831 ( .A(n17372), .B(n17373), .Z(n17272) );
  OR U21832 ( .A(n17374), .B(n17375), .Z(n17373) );
  OR U21833 ( .A(n17376), .B(n17377), .Z(n17372) );
  NAND U21834 ( .A(n17378), .B(n17379), .Z(n17270) );
  OR U21835 ( .A(n17380), .B(n17381), .Z(n17379) );
  OR U21836 ( .A(n17382), .B(n17383), .Z(n17378) );
  ANDN U21837 ( .B(n17384), .A(n17385), .Z(n17271) );
  IV U21838 ( .A(n17386), .Z(n17384) );
  XNOR U21839 ( .A(n17351), .B(n17350), .Z(N28733) );
  XOR U21840 ( .A(n17370), .B(n17369), .Z(n17350) );
  XNOR U21841 ( .A(n17385), .B(n17386), .Z(n17369) );
  XNOR U21842 ( .A(n17380), .B(n17381), .Z(n17386) );
  XNOR U21843 ( .A(n17382), .B(n17383), .Z(n17381) );
  XNOR U21844 ( .A(y[1612]), .B(x[1612]), .Z(n17383) );
  XNOR U21845 ( .A(y[1613]), .B(x[1613]), .Z(n17382) );
  XNOR U21846 ( .A(y[1611]), .B(x[1611]), .Z(n17380) );
  XNOR U21847 ( .A(n17374), .B(n17375), .Z(n17385) );
  XNOR U21848 ( .A(y[1608]), .B(x[1608]), .Z(n17375) );
  XNOR U21849 ( .A(n17376), .B(n17377), .Z(n17374) );
  XNOR U21850 ( .A(y[1609]), .B(x[1609]), .Z(n17377) );
  XNOR U21851 ( .A(y[1610]), .B(x[1610]), .Z(n17376) );
  XNOR U21852 ( .A(n17367), .B(n17366), .Z(n17370) );
  XNOR U21853 ( .A(n17362), .B(n17363), .Z(n17366) );
  XNOR U21854 ( .A(y[1605]), .B(x[1605]), .Z(n17363) );
  XNOR U21855 ( .A(n17364), .B(n17365), .Z(n17362) );
  XNOR U21856 ( .A(y[1606]), .B(x[1606]), .Z(n17365) );
  XNOR U21857 ( .A(y[1607]), .B(x[1607]), .Z(n17364) );
  XNOR U21858 ( .A(n17356), .B(n17357), .Z(n17367) );
  XNOR U21859 ( .A(y[1602]), .B(x[1602]), .Z(n17357) );
  XNOR U21860 ( .A(n17358), .B(n17359), .Z(n17356) );
  XNOR U21861 ( .A(y[1603]), .B(x[1603]), .Z(n17359) );
  XNOR U21862 ( .A(y[1604]), .B(x[1604]), .Z(n17358) );
  XOR U21863 ( .A(n17332), .B(n17333), .Z(n17351) );
  XNOR U21864 ( .A(n17348), .B(n17349), .Z(n17333) );
  XNOR U21865 ( .A(n17343), .B(n17344), .Z(n17349) );
  XNOR U21866 ( .A(n17345), .B(n17346), .Z(n17344) );
  XNOR U21867 ( .A(y[1600]), .B(x[1600]), .Z(n17346) );
  XNOR U21868 ( .A(y[1601]), .B(x[1601]), .Z(n17345) );
  XNOR U21869 ( .A(y[1599]), .B(x[1599]), .Z(n17343) );
  XNOR U21870 ( .A(n17337), .B(n17338), .Z(n17348) );
  XNOR U21871 ( .A(y[1596]), .B(x[1596]), .Z(n17338) );
  XNOR U21872 ( .A(n17339), .B(n17340), .Z(n17337) );
  XNOR U21873 ( .A(y[1597]), .B(x[1597]), .Z(n17340) );
  XNOR U21874 ( .A(y[1598]), .B(x[1598]), .Z(n17339) );
  XOR U21875 ( .A(n17331), .B(n17330), .Z(n17332) );
  XNOR U21876 ( .A(n17326), .B(n17327), .Z(n17330) );
  XNOR U21877 ( .A(y[1593]), .B(x[1593]), .Z(n17327) );
  XNOR U21878 ( .A(n17328), .B(n17329), .Z(n17326) );
  XNOR U21879 ( .A(y[1594]), .B(x[1594]), .Z(n17329) );
  XNOR U21880 ( .A(y[1595]), .B(x[1595]), .Z(n17328) );
  XNOR U21881 ( .A(n17320), .B(n17321), .Z(n17331) );
  XNOR U21882 ( .A(y[1590]), .B(x[1590]), .Z(n17321) );
  XNOR U21883 ( .A(n17322), .B(n17323), .Z(n17320) );
  XNOR U21884 ( .A(y[1591]), .B(x[1591]), .Z(n17323) );
  XNOR U21885 ( .A(y[1592]), .B(x[1592]), .Z(n17322) );
  NAND U21886 ( .A(n17387), .B(n17388), .Z(N28725) );
  NANDN U21887 ( .A(n17389), .B(n17390), .Z(n17388) );
  OR U21888 ( .A(n17391), .B(n17392), .Z(n17390) );
  NAND U21889 ( .A(n17391), .B(n17392), .Z(n17387) );
  XOR U21890 ( .A(n17391), .B(n17393), .Z(N28724) );
  XNOR U21891 ( .A(n17389), .B(n17392), .Z(n17393) );
  AND U21892 ( .A(n17394), .B(n17395), .Z(n17392) );
  NANDN U21893 ( .A(n17396), .B(n17397), .Z(n17395) );
  NANDN U21894 ( .A(n17398), .B(n17399), .Z(n17397) );
  NANDN U21895 ( .A(n17399), .B(n17398), .Z(n17394) );
  NAND U21896 ( .A(n17400), .B(n17401), .Z(n17389) );
  NANDN U21897 ( .A(n17402), .B(n17403), .Z(n17401) );
  OR U21898 ( .A(n17404), .B(n17405), .Z(n17403) );
  NAND U21899 ( .A(n17405), .B(n17404), .Z(n17400) );
  AND U21900 ( .A(n17406), .B(n17407), .Z(n17391) );
  NANDN U21901 ( .A(n17408), .B(n17409), .Z(n17407) );
  NANDN U21902 ( .A(n17410), .B(n17411), .Z(n17409) );
  NANDN U21903 ( .A(n17411), .B(n17410), .Z(n17406) );
  XOR U21904 ( .A(n17405), .B(n17412), .Z(N28723) );
  XOR U21905 ( .A(n17402), .B(n17404), .Z(n17412) );
  XNOR U21906 ( .A(n17398), .B(n17413), .Z(n17404) );
  XNOR U21907 ( .A(n17396), .B(n17399), .Z(n17413) );
  NAND U21908 ( .A(n17414), .B(n17415), .Z(n17399) );
  NAND U21909 ( .A(n17416), .B(n17417), .Z(n17415) );
  OR U21910 ( .A(n17418), .B(n17419), .Z(n17416) );
  NANDN U21911 ( .A(n17420), .B(n17418), .Z(n17414) );
  IV U21912 ( .A(n17419), .Z(n17420) );
  NAND U21913 ( .A(n17421), .B(n17422), .Z(n17396) );
  NAND U21914 ( .A(n17423), .B(n17424), .Z(n17422) );
  NANDN U21915 ( .A(n17425), .B(n17426), .Z(n17423) );
  NANDN U21916 ( .A(n17426), .B(n17425), .Z(n17421) );
  AND U21917 ( .A(n17427), .B(n17428), .Z(n17398) );
  NAND U21918 ( .A(n17429), .B(n17430), .Z(n17428) );
  OR U21919 ( .A(n17431), .B(n17432), .Z(n17429) );
  NANDN U21920 ( .A(n17433), .B(n17431), .Z(n17427) );
  NAND U21921 ( .A(n17434), .B(n17435), .Z(n17402) );
  NANDN U21922 ( .A(n17436), .B(n17437), .Z(n17435) );
  OR U21923 ( .A(n17438), .B(n17439), .Z(n17437) );
  NANDN U21924 ( .A(n17440), .B(n17438), .Z(n17434) );
  IV U21925 ( .A(n17439), .Z(n17440) );
  XNOR U21926 ( .A(n17410), .B(n17441), .Z(n17405) );
  XNOR U21927 ( .A(n17408), .B(n17411), .Z(n17441) );
  NAND U21928 ( .A(n17442), .B(n17443), .Z(n17411) );
  NAND U21929 ( .A(n17444), .B(n17445), .Z(n17443) );
  OR U21930 ( .A(n17446), .B(n17447), .Z(n17444) );
  NANDN U21931 ( .A(n17448), .B(n17446), .Z(n17442) );
  IV U21932 ( .A(n17447), .Z(n17448) );
  NAND U21933 ( .A(n17449), .B(n17450), .Z(n17408) );
  NAND U21934 ( .A(n17451), .B(n17452), .Z(n17450) );
  NANDN U21935 ( .A(n17453), .B(n17454), .Z(n17451) );
  NANDN U21936 ( .A(n17454), .B(n17453), .Z(n17449) );
  AND U21937 ( .A(n17455), .B(n17456), .Z(n17410) );
  NAND U21938 ( .A(n17457), .B(n17458), .Z(n17456) );
  OR U21939 ( .A(n17459), .B(n17460), .Z(n17457) );
  NANDN U21940 ( .A(n17461), .B(n17459), .Z(n17455) );
  XNOR U21941 ( .A(n17436), .B(n17462), .Z(N28722) );
  XOR U21942 ( .A(n17438), .B(n17439), .Z(n17462) );
  XNOR U21943 ( .A(n17452), .B(n17463), .Z(n17439) );
  XOR U21944 ( .A(n17453), .B(n17454), .Z(n17463) );
  XOR U21945 ( .A(n17459), .B(n17464), .Z(n17454) );
  XOR U21946 ( .A(n17458), .B(n17461), .Z(n17464) );
  IV U21947 ( .A(n17460), .Z(n17461) );
  NAND U21948 ( .A(n17465), .B(n17466), .Z(n17460) );
  OR U21949 ( .A(n17467), .B(n17468), .Z(n17466) );
  OR U21950 ( .A(n17469), .B(n17470), .Z(n17465) );
  NAND U21951 ( .A(n17471), .B(n17472), .Z(n17458) );
  OR U21952 ( .A(n17473), .B(n17474), .Z(n17472) );
  OR U21953 ( .A(n17475), .B(n17476), .Z(n17471) );
  NOR U21954 ( .A(n17477), .B(n17478), .Z(n17459) );
  ANDN U21955 ( .B(n17479), .A(n17480), .Z(n17453) );
  XNOR U21956 ( .A(n17446), .B(n17481), .Z(n17452) );
  XNOR U21957 ( .A(n17445), .B(n17447), .Z(n17481) );
  NAND U21958 ( .A(n17482), .B(n17483), .Z(n17447) );
  OR U21959 ( .A(n17484), .B(n17485), .Z(n17483) );
  OR U21960 ( .A(n17486), .B(n17487), .Z(n17482) );
  NAND U21961 ( .A(n17488), .B(n17489), .Z(n17445) );
  OR U21962 ( .A(n17490), .B(n17491), .Z(n17489) );
  OR U21963 ( .A(n17492), .B(n17493), .Z(n17488) );
  ANDN U21964 ( .B(n17494), .A(n17495), .Z(n17446) );
  IV U21965 ( .A(n17496), .Z(n17494) );
  ANDN U21966 ( .B(n17497), .A(n17498), .Z(n17438) );
  XOR U21967 ( .A(n17424), .B(n17499), .Z(n17436) );
  XOR U21968 ( .A(n17425), .B(n17426), .Z(n17499) );
  XOR U21969 ( .A(n17431), .B(n17500), .Z(n17426) );
  XOR U21970 ( .A(n17430), .B(n17433), .Z(n17500) );
  IV U21971 ( .A(n17432), .Z(n17433) );
  NAND U21972 ( .A(n17501), .B(n17502), .Z(n17432) );
  OR U21973 ( .A(n17503), .B(n17504), .Z(n17502) );
  OR U21974 ( .A(n17505), .B(n17506), .Z(n17501) );
  NAND U21975 ( .A(n17507), .B(n17508), .Z(n17430) );
  OR U21976 ( .A(n17509), .B(n17510), .Z(n17508) );
  OR U21977 ( .A(n17511), .B(n17512), .Z(n17507) );
  NOR U21978 ( .A(n17513), .B(n17514), .Z(n17431) );
  ANDN U21979 ( .B(n17515), .A(n17516), .Z(n17425) );
  IV U21980 ( .A(n17517), .Z(n17515) );
  XNOR U21981 ( .A(n17418), .B(n17518), .Z(n17424) );
  XNOR U21982 ( .A(n17417), .B(n17419), .Z(n17518) );
  NAND U21983 ( .A(n17519), .B(n17520), .Z(n17419) );
  OR U21984 ( .A(n17521), .B(n17522), .Z(n17520) );
  OR U21985 ( .A(n17523), .B(n17524), .Z(n17519) );
  NAND U21986 ( .A(n17525), .B(n17526), .Z(n17417) );
  OR U21987 ( .A(n17527), .B(n17528), .Z(n17526) );
  OR U21988 ( .A(n17529), .B(n17530), .Z(n17525) );
  ANDN U21989 ( .B(n17531), .A(n17532), .Z(n17418) );
  IV U21990 ( .A(n17533), .Z(n17531) );
  XNOR U21991 ( .A(n17498), .B(n17497), .Z(N28721) );
  XOR U21992 ( .A(n17517), .B(n17516), .Z(n17497) );
  XNOR U21993 ( .A(n17532), .B(n17533), .Z(n17516) );
  XNOR U21994 ( .A(n17527), .B(n17528), .Z(n17533) );
  XNOR U21995 ( .A(n17529), .B(n17530), .Z(n17528) );
  XNOR U21996 ( .A(y[1588]), .B(x[1588]), .Z(n17530) );
  XNOR U21997 ( .A(y[1589]), .B(x[1589]), .Z(n17529) );
  XNOR U21998 ( .A(y[1587]), .B(x[1587]), .Z(n17527) );
  XNOR U21999 ( .A(n17521), .B(n17522), .Z(n17532) );
  XNOR U22000 ( .A(y[1584]), .B(x[1584]), .Z(n17522) );
  XNOR U22001 ( .A(n17523), .B(n17524), .Z(n17521) );
  XNOR U22002 ( .A(y[1585]), .B(x[1585]), .Z(n17524) );
  XNOR U22003 ( .A(y[1586]), .B(x[1586]), .Z(n17523) );
  XNOR U22004 ( .A(n17514), .B(n17513), .Z(n17517) );
  XNOR U22005 ( .A(n17509), .B(n17510), .Z(n17513) );
  XNOR U22006 ( .A(y[1581]), .B(x[1581]), .Z(n17510) );
  XNOR U22007 ( .A(n17511), .B(n17512), .Z(n17509) );
  XNOR U22008 ( .A(y[1582]), .B(x[1582]), .Z(n17512) );
  XNOR U22009 ( .A(y[1583]), .B(x[1583]), .Z(n17511) );
  XNOR U22010 ( .A(n17503), .B(n17504), .Z(n17514) );
  XNOR U22011 ( .A(y[1578]), .B(x[1578]), .Z(n17504) );
  XNOR U22012 ( .A(n17505), .B(n17506), .Z(n17503) );
  XNOR U22013 ( .A(y[1579]), .B(x[1579]), .Z(n17506) );
  XNOR U22014 ( .A(y[1580]), .B(x[1580]), .Z(n17505) );
  XOR U22015 ( .A(n17479), .B(n17480), .Z(n17498) );
  XNOR U22016 ( .A(n17495), .B(n17496), .Z(n17480) );
  XNOR U22017 ( .A(n17490), .B(n17491), .Z(n17496) );
  XNOR U22018 ( .A(n17492), .B(n17493), .Z(n17491) );
  XNOR U22019 ( .A(y[1576]), .B(x[1576]), .Z(n17493) );
  XNOR U22020 ( .A(y[1577]), .B(x[1577]), .Z(n17492) );
  XNOR U22021 ( .A(y[1575]), .B(x[1575]), .Z(n17490) );
  XNOR U22022 ( .A(n17484), .B(n17485), .Z(n17495) );
  XNOR U22023 ( .A(y[1572]), .B(x[1572]), .Z(n17485) );
  XNOR U22024 ( .A(n17486), .B(n17487), .Z(n17484) );
  XNOR U22025 ( .A(y[1573]), .B(x[1573]), .Z(n17487) );
  XNOR U22026 ( .A(y[1574]), .B(x[1574]), .Z(n17486) );
  XOR U22027 ( .A(n17478), .B(n17477), .Z(n17479) );
  XNOR U22028 ( .A(n17473), .B(n17474), .Z(n17477) );
  XNOR U22029 ( .A(y[1569]), .B(x[1569]), .Z(n17474) );
  XNOR U22030 ( .A(n17475), .B(n17476), .Z(n17473) );
  XNOR U22031 ( .A(y[1570]), .B(x[1570]), .Z(n17476) );
  XNOR U22032 ( .A(y[1571]), .B(x[1571]), .Z(n17475) );
  XNOR U22033 ( .A(n17467), .B(n17468), .Z(n17478) );
  XNOR U22034 ( .A(y[1566]), .B(x[1566]), .Z(n17468) );
  XNOR U22035 ( .A(n17469), .B(n17470), .Z(n17467) );
  XNOR U22036 ( .A(y[1567]), .B(x[1567]), .Z(n17470) );
  XNOR U22037 ( .A(y[1568]), .B(x[1568]), .Z(n17469) );
  NAND U22038 ( .A(n17534), .B(n17535), .Z(N28713) );
  NANDN U22039 ( .A(n17536), .B(n17537), .Z(n17535) );
  OR U22040 ( .A(n17538), .B(n17539), .Z(n17537) );
  NAND U22041 ( .A(n17538), .B(n17539), .Z(n17534) );
  XOR U22042 ( .A(n17538), .B(n17540), .Z(N28712) );
  XNOR U22043 ( .A(n17536), .B(n17539), .Z(n17540) );
  AND U22044 ( .A(n17541), .B(n17542), .Z(n17539) );
  NANDN U22045 ( .A(n17543), .B(n17544), .Z(n17542) );
  NANDN U22046 ( .A(n17545), .B(n17546), .Z(n17544) );
  NANDN U22047 ( .A(n17546), .B(n17545), .Z(n17541) );
  NAND U22048 ( .A(n17547), .B(n17548), .Z(n17536) );
  NANDN U22049 ( .A(n17549), .B(n17550), .Z(n17548) );
  OR U22050 ( .A(n17551), .B(n17552), .Z(n17550) );
  NAND U22051 ( .A(n17552), .B(n17551), .Z(n17547) );
  AND U22052 ( .A(n17553), .B(n17554), .Z(n17538) );
  NANDN U22053 ( .A(n17555), .B(n17556), .Z(n17554) );
  NANDN U22054 ( .A(n17557), .B(n17558), .Z(n17556) );
  NANDN U22055 ( .A(n17558), .B(n17557), .Z(n17553) );
  XOR U22056 ( .A(n17552), .B(n17559), .Z(N28711) );
  XOR U22057 ( .A(n17549), .B(n17551), .Z(n17559) );
  XNOR U22058 ( .A(n17545), .B(n17560), .Z(n17551) );
  XNOR U22059 ( .A(n17543), .B(n17546), .Z(n17560) );
  NAND U22060 ( .A(n17561), .B(n17562), .Z(n17546) );
  NAND U22061 ( .A(n17563), .B(n17564), .Z(n17562) );
  OR U22062 ( .A(n17565), .B(n17566), .Z(n17563) );
  NANDN U22063 ( .A(n17567), .B(n17565), .Z(n17561) );
  IV U22064 ( .A(n17566), .Z(n17567) );
  NAND U22065 ( .A(n17568), .B(n17569), .Z(n17543) );
  NAND U22066 ( .A(n17570), .B(n17571), .Z(n17569) );
  NANDN U22067 ( .A(n17572), .B(n17573), .Z(n17570) );
  NANDN U22068 ( .A(n17573), .B(n17572), .Z(n17568) );
  AND U22069 ( .A(n17574), .B(n17575), .Z(n17545) );
  NAND U22070 ( .A(n17576), .B(n17577), .Z(n17575) );
  OR U22071 ( .A(n17578), .B(n17579), .Z(n17576) );
  NANDN U22072 ( .A(n17580), .B(n17578), .Z(n17574) );
  NAND U22073 ( .A(n17581), .B(n17582), .Z(n17549) );
  NANDN U22074 ( .A(n17583), .B(n17584), .Z(n17582) );
  OR U22075 ( .A(n17585), .B(n17586), .Z(n17584) );
  NANDN U22076 ( .A(n17587), .B(n17585), .Z(n17581) );
  IV U22077 ( .A(n17586), .Z(n17587) );
  XNOR U22078 ( .A(n17557), .B(n17588), .Z(n17552) );
  XNOR U22079 ( .A(n17555), .B(n17558), .Z(n17588) );
  NAND U22080 ( .A(n17589), .B(n17590), .Z(n17558) );
  NAND U22081 ( .A(n17591), .B(n17592), .Z(n17590) );
  OR U22082 ( .A(n17593), .B(n17594), .Z(n17591) );
  NANDN U22083 ( .A(n17595), .B(n17593), .Z(n17589) );
  IV U22084 ( .A(n17594), .Z(n17595) );
  NAND U22085 ( .A(n17596), .B(n17597), .Z(n17555) );
  NAND U22086 ( .A(n17598), .B(n17599), .Z(n17597) );
  NANDN U22087 ( .A(n17600), .B(n17601), .Z(n17598) );
  NANDN U22088 ( .A(n17601), .B(n17600), .Z(n17596) );
  AND U22089 ( .A(n17602), .B(n17603), .Z(n17557) );
  NAND U22090 ( .A(n17604), .B(n17605), .Z(n17603) );
  OR U22091 ( .A(n17606), .B(n17607), .Z(n17604) );
  NANDN U22092 ( .A(n17608), .B(n17606), .Z(n17602) );
  XNOR U22093 ( .A(n17583), .B(n17609), .Z(N28710) );
  XOR U22094 ( .A(n17585), .B(n17586), .Z(n17609) );
  XNOR U22095 ( .A(n17599), .B(n17610), .Z(n17586) );
  XOR U22096 ( .A(n17600), .B(n17601), .Z(n17610) );
  XOR U22097 ( .A(n17606), .B(n17611), .Z(n17601) );
  XOR U22098 ( .A(n17605), .B(n17608), .Z(n17611) );
  IV U22099 ( .A(n17607), .Z(n17608) );
  NAND U22100 ( .A(n17612), .B(n17613), .Z(n17607) );
  OR U22101 ( .A(n17614), .B(n17615), .Z(n17613) );
  OR U22102 ( .A(n17616), .B(n17617), .Z(n17612) );
  NAND U22103 ( .A(n17618), .B(n17619), .Z(n17605) );
  OR U22104 ( .A(n17620), .B(n17621), .Z(n17619) );
  OR U22105 ( .A(n17622), .B(n17623), .Z(n17618) );
  NOR U22106 ( .A(n17624), .B(n17625), .Z(n17606) );
  ANDN U22107 ( .B(n17626), .A(n17627), .Z(n17600) );
  XNOR U22108 ( .A(n17593), .B(n17628), .Z(n17599) );
  XNOR U22109 ( .A(n17592), .B(n17594), .Z(n17628) );
  NAND U22110 ( .A(n17629), .B(n17630), .Z(n17594) );
  OR U22111 ( .A(n17631), .B(n17632), .Z(n17630) );
  OR U22112 ( .A(n17633), .B(n17634), .Z(n17629) );
  NAND U22113 ( .A(n17635), .B(n17636), .Z(n17592) );
  OR U22114 ( .A(n17637), .B(n17638), .Z(n17636) );
  OR U22115 ( .A(n17639), .B(n17640), .Z(n17635) );
  ANDN U22116 ( .B(n17641), .A(n17642), .Z(n17593) );
  IV U22117 ( .A(n17643), .Z(n17641) );
  ANDN U22118 ( .B(n17644), .A(n17645), .Z(n17585) );
  XOR U22119 ( .A(n17571), .B(n17646), .Z(n17583) );
  XOR U22120 ( .A(n17572), .B(n17573), .Z(n17646) );
  XOR U22121 ( .A(n17578), .B(n17647), .Z(n17573) );
  XOR U22122 ( .A(n17577), .B(n17580), .Z(n17647) );
  IV U22123 ( .A(n17579), .Z(n17580) );
  NAND U22124 ( .A(n17648), .B(n17649), .Z(n17579) );
  OR U22125 ( .A(n17650), .B(n17651), .Z(n17649) );
  OR U22126 ( .A(n17652), .B(n17653), .Z(n17648) );
  NAND U22127 ( .A(n17654), .B(n17655), .Z(n17577) );
  OR U22128 ( .A(n17656), .B(n17657), .Z(n17655) );
  OR U22129 ( .A(n17658), .B(n17659), .Z(n17654) );
  NOR U22130 ( .A(n17660), .B(n17661), .Z(n17578) );
  ANDN U22131 ( .B(n17662), .A(n17663), .Z(n17572) );
  IV U22132 ( .A(n17664), .Z(n17662) );
  XNOR U22133 ( .A(n17565), .B(n17665), .Z(n17571) );
  XNOR U22134 ( .A(n17564), .B(n17566), .Z(n17665) );
  NAND U22135 ( .A(n17666), .B(n17667), .Z(n17566) );
  OR U22136 ( .A(n17668), .B(n17669), .Z(n17667) );
  OR U22137 ( .A(n17670), .B(n17671), .Z(n17666) );
  NAND U22138 ( .A(n17672), .B(n17673), .Z(n17564) );
  OR U22139 ( .A(n17674), .B(n17675), .Z(n17673) );
  OR U22140 ( .A(n17676), .B(n17677), .Z(n17672) );
  ANDN U22141 ( .B(n17678), .A(n17679), .Z(n17565) );
  IV U22142 ( .A(n17680), .Z(n17678) );
  XNOR U22143 ( .A(n17645), .B(n17644), .Z(N28709) );
  XOR U22144 ( .A(n17664), .B(n17663), .Z(n17644) );
  XNOR U22145 ( .A(n17679), .B(n17680), .Z(n17663) );
  XNOR U22146 ( .A(n17674), .B(n17675), .Z(n17680) );
  XNOR U22147 ( .A(n17676), .B(n17677), .Z(n17675) );
  XNOR U22148 ( .A(y[1564]), .B(x[1564]), .Z(n17677) );
  XNOR U22149 ( .A(y[1565]), .B(x[1565]), .Z(n17676) );
  XNOR U22150 ( .A(y[1563]), .B(x[1563]), .Z(n17674) );
  XNOR U22151 ( .A(n17668), .B(n17669), .Z(n17679) );
  XNOR U22152 ( .A(y[1560]), .B(x[1560]), .Z(n17669) );
  XNOR U22153 ( .A(n17670), .B(n17671), .Z(n17668) );
  XNOR U22154 ( .A(y[1561]), .B(x[1561]), .Z(n17671) );
  XNOR U22155 ( .A(y[1562]), .B(x[1562]), .Z(n17670) );
  XNOR U22156 ( .A(n17661), .B(n17660), .Z(n17664) );
  XNOR U22157 ( .A(n17656), .B(n17657), .Z(n17660) );
  XNOR U22158 ( .A(y[1557]), .B(x[1557]), .Z(n17657) );
  XNOR U22159 ( .A(n17658), .B(n17659), .Z(n17656) );
  XNOR U22160 ( .A(y[1558]), .B(x[1558]), .Z(n17659) );
  XNOR U22161 ( .A(y[1559]), .B(x[1559]), .Z(n17658) );
  XNOR U22162 ( .A(n17650), .B(n17651), .Z(n17661) );
  XNOR U22163 ( .A(y[1554]), .B(x[1554]), .Z(n17651) );
  XNOR U22164 ( .A(n17652), .B(n17653), .Z(n17650) );
  XNOR U22165 ( .A(y[1555]), .B(x[1555]), .Z(n17653) );
  XNOR U22166 ( .A(y[1556]), .B(x[1556]), .Z(n17652) );
  XOR U22167 ( .A(n17626), .B(n17627), .Z(n17645) );
  XNOR U22168 ( .A(n17642), .B(n17643), .Z(n17627) );
  XNOR U22169 ( .A(n17637), .B(n17638), .Z(n17643) );
  XNOR U22170 ( .A(n17639), .B(n17640), .Z(n17638) );
  XNOR U22171 ( .A(y[1552]), .B(x[1552]), .Z(n17640) );
  XNOR U22172 ( .A(y[1553]), .B(x[1553]), .Z(n17639) );
  XNOR U22173 ( .A(y[1551]), .B(x[1551]), .Z(n17637) );
  XNOR U22174 ( .A(n17631), .B(n17632), .Z(n17642) );
  XNOR U22175 ( .A(y[1548]), .B(x[1548]), .Z(n17632) );
  XNOR U22176 ( .A(n17633), .B(n17634), .Z(n17631) );
  XNOR U22177 ( .A(y[1549]), .B(x[1549]), .Z(n17634) );
  XNOR U22178 ( .A(y[1550]), .B(x[1550]), .Z(n17633) );
  XOR U22179 ( .A(n17625), .B(n17624), .Z(n17626) );
  XNOR U22180 ( .A(n17620), .B(n17621), .Z(n17624) );
  XNOR U22181 ( .A(y[1545]), .B(x[1545]), .Z(n17621) );
  XNOR U22182 ( .A(n17622), .B(n17623), .Z(n17620) );
  XNOR U22183 ( .A(y[1546]), .B(x[1546]), .Z(n17623) );
  XNOR U22184 ( .A(y[1547]), .B(x[1547]), .Z(n17622) );
  XNOR U22185 ( .A(n17614), .B(n17615), .Z(n17625) );
  XNOR U22186 ( .A(y[1542]), .B(x[1542]), .Z(n17615) );
  XNOR U22187 ( .A(n17616), .B(n17617), .Z(n17614) );
  XNOR U22188 ( .A(y[1543]), .B(x[1543]), .Z(n17617) );
  XNOR U22189 ( .A(y[1544]), .B(x[1544]), .Z(n17616) );
  NAND U22190 ( .A(n17681), .B(n17682), .Z(N28701) );
  NANDN U22191 ( .A(n17683), .B(n17684), .Z(n17682) );
  OR U22192 ( .A(n17685), .B(n17686), .Z(n17684) );
  NAND U22193 ( .A(n17685), .B(n17686), .Z(n17681) );
  XOR U22194 ( .A(n17685), .B(n17687), .Z(N28700) );
  XNOR U22195 ( .A(n17683), .B(n17686), .Z(n17687) );
  AND U22196 ( .A(n17688), .B(n17689), .Z(n17686) );
  NANDN U22197 ( .A(n17690), .B(n17691), .Z(n17689) );
  NANDN U22198 ( .A(n17692), .B(n17693), .Z(n17691) );
  NANDN U22199 ( .A(n17693), .B(n17692), .Z(n17688) );
  NAND U22200 ( .A(n17694), .B(n17695), .Z(n17683) );
  NANDN U22201 ( .A(n17696), .B(n17697), .Z(n17695) );
  OR U22202 ( .A(n17698), .B(n17699), .Z(n17697) );
  NAND U22203 ( .A(n17699), .B(n17698), .Z(n17694) );
  AND U22204 ( .A(n17700), .B(n17701), .Z(n17685) );
  NANDN U22205 ( .A(n17702), .B(n17703), .Z(n17701) );
  NANDN U22206 ( .A(n17704), .B(n17705), .Z(n17703) );
  NANDN U22207 ( .A(n17705), .B(n17704), .Z(n17700) );
  XOR U22208 ( .A(n17699), .B(n17706), .Z(N28699) );
  XOR U22209 ( .A(n17696), .B(n17698), .Z(n17706) );
  XNOR U22210 ( .A(n17692), .B(n17707), .Z(n17698) );
  XNOR U22211 ( .A(n17690), .B(n17693), .Z(n17707) );
  NAND U22212 ( .A(n17708), .B(n17709), .Z(n17693) );
  NAND U22213 ( .A(n17710), .B(n17711), .Z(n17709) );
  OR U22214 ( .A(n17712), .B(n17713), .Z(n17710) );
  NANDN U22215 ( .A(n17714), .B(n17712), .Z(n17708) );
  IV U22216 ( .A(n17713), .Z(n17714) );
  NAND U22217 ( .A(n17715), .B(n17716), .Z(n17690) );
  NAND U22218 ( .A(n17717), .B(n17718), .Z(n17716) );
  NANDN U22219 ( .A(n17719), .B(n17720), .Z(n17717) );
  NANDN U22220 ( .A(n17720), .B(n17719), .Z(n17715) );
  AND U22221 ( .A(n17721), .B(n17722), .Z(n17692) );
  NAND U22222 ( .A(n17723), .B(n17724), .Z(n17722) );
  OR U22223 ( .A(n17725), .B(n17726), .Z(n17723) );
  NANDN U22224 ( .A(n17727), .B(n17725), .Z(n17721) );
  NAND U22225 ( .A(n17728), .B(n17729), .Z(n17696) );
  NANDN U22226 ( .A(n17730), .B(n17731), .Z(n17729) );
  OR U22227 ( .A(n17732), .B(n17733), .Z(n17731) );
  NANDN U22228 ( .A(n17734), .B(n17732), .Z(n17728) );
  IV U22229 ( .A(n17733), .Z(n17734) );
  XNOR U22230 ( .A(n17704), .B(n17735), .Z(n17699) );
  XNOR U22231 ( .A(n17702), .B(n17705), .Z(n17735) );
  NAND U22232 ( .A(n17736), .B(n17737), .Z(n17705) );
  NAND U22233 ( .A(n17738), .B(n17739), .Z(n17737) );
  OR U22234 ( .A(n17740), .B(n17741), .Z(n17738) );
  NANDN U22235 ( .A(n17742), .B(n17740), .Z(n17736) );
  IV U22236 ( .A(n17741), .Z(n17742) );
  NAND U22237 ( .A(n17743), .B(n17744), .Z(n17702) );
  NAND U22238 ( .A(n17745), .B(n17746), .Z(n17744) );
  NANDN U22239 ( .A(n17747), .B(n17748), .Z(n17745) );
  NANDN U22240 ( .A(n17748), .B(n17747), .Z(n17743) );
  AND U22241 ( .A(n17749), .B(n17750), .Z(n17704) );
  NAND U22242 ( .A(n17751), .B(n17752), .Z(n17750) );
  OR U22243 ( .A(n17753), .B(n17754), .Z(n17751) );
  NANDN U22244 ( .A(n17755), .B(n17753), .Z(n17749) );
  XNOR U22245 ( .A(n17730), .B(n17756), .Z(N28698) );
  XOR U22246 ( .A(n17732), .B(n17733), .Z(n17756) );
  XNOR U22247 ( .A(n17746), .B(n17757), .Z(n17733) );
  XOR U22248 ( .A(n17747), .B(n17748), .Z(n17757) );
  XOR U22249 ( .A(n17753), .B(n17758), .Z(n17748) );
  XOR U22250 ( .A(n17752), .B(n17755), .Z(n17758) );
  IV U22251 ( .A(n17754), .Z(n17755) );
  NAND U22252 ( .A(n17759), .B(n17760), .Z(n17754) );
  OR U22253 ( .A(n17761), .B(n17762), .Z(n17760) );
  OR U22254 ( .A(n17763), .B(n17764), .Z(n17759) );
  NAND U22255 ( .A(n17765), .B(n17766), .Z(n17752) );
  OR U22256 ( .A(n17767), .B(n17768), .Z(n17766) );
  OR U22257 ( .A(n17769), .B(n17770), .Z(n17765) );
  NOR U22258 ( .A(n17771), .B(n17772), .Z(n17753) );
  ANDN U22259 ( .B(n17773), .A(n17774), .Z(n17747) );
  XNOR U22260 ( .A(n17740), .B(n17775), .Z(n17746) );
  XNOR U22261 ( .A(n17739), .B(n17741), .Z(n17775) );
  NAND U22262 ( .A(n17776), .B(n17777), .Z(n17741) );
  OR U22263 ( .A(n17778), .B(n17779), .Z(n17777) );
  OR U22264 ( .A(n17780), .B(n17781), .Z(n17776) );
  NAND U22265 ( .A(n17782), .B(n17783), .Z(n17739) );
  OR U22266 ( .A(n17784), .B(n17785), .Z(n17783) );
  OR U22267 ( .A(n17786), .B(n17787), .Z(n17782) );
  ANDN U22268 ( .B(n17788), .A(n17789), .Z(n17740) );
  IV U22269 ( .A(n17790), .Z(n17788) );
  ANDN U22270 ( .B(n17791), .A(n17792), .Z(n17732) );
  XOR U22271 ( .A(n17718), .B(n17793), .Z(n17730) );
  XOR U22272 ( .A(n17719), .B(n17720), .Z(n17793) );
  XOR U22273 ( .A(n17725), .B(n17794), .Z(n17720) );
  XOR U22274 ( .A(n17724), .B(n17727), .Z(n17794) );
  IV U22275 ( .A(n17726), .Z(n17727) );
  NAND U22276 ( .A(n17795), .B(n17796), .Z(n17726) );
  OR U22277 ( .A(n17797), .B(n17798), .Z(n17796) );
  OR U22278 ( .A(n17799), .B(n17800), .Z(n17795) );
  NAND U22279 ( .A(n17801), .B(n17802), .Z(n17724) );
  OR U22280 ( .A(n17803), .B(n17804), .Z(n17802) );
  OR U22281 ( .A(n17805), .B(n17806), .Z(n17801) );
  NOR U22282 ( .A(n17807), .B(n17808), .Z(n17725) );
  ANDN U22283 ( .B(n17809), .A(n17810), .Z(n17719) );
  IV U22284 ( .A(n17811), .Z(n17809) );
  XNOR U22285 ( .A(n17712), .B(n17812), .Z(n17718) );
  XNOR U22286 ( .A(n17711), .B(n17713), .Z(n17812) );
  NAND U22287 ( .A(n17813), .B(n17814), .Z(n17713) );
  OR U22288 ( .A(n17815), .B(n17816), .Z(n17814) );
  OR U22289 ( .A(n17817), .B(n17818), .Z(n17813) );
  NAND U22290 ( .A(n17819), .B(n17820), .Z(n17711) );
  OR U22291 ( .A(n17821), .B(n17822), .Z(n17820) );
  OR U22292 ( .A(n17823), .B(n17824), .Z(n17819) );
  ANDN U22293 ( .B(n17825), .A(n17826), .Z(n17712) );
  IV U22294 ( .A(n17827), .Z(n17825) );
  XNOR U22295 ( .A(n17792), .B(n17791), .Z(N28697) );
  XOR U22296 ( .A(n17811), .B(n17810), .Z(n17791) );
  XNOR U22297 ( .A(n17826), .B(n17827), .Z(n17810) );
  XNOR U22298 ( .A(n17821), .B(n17822), .Z(n17827) );
  XNOR U22299 ( .A(n17823), .B(n17824), .Z(n17822) );
  XNOR U22300 ( .A(y[1540]), .B(x[1540]), .Z(n17824) );
  XNOR U22301 ( .A(y[1541]), .B(x[1541]), .Z(n17823) );
  XNOR U22302 ( .A(y[1539]), .B(x[1539]), .Z(n17821) );
  XNOR U22303 ( .A(n17815), .B(n17816), .Z(n17826) );
  XNOR U22304 ( .A(y[1536]), .B(x[1536]), .Z(n17816) );
  XNOR U22305 ( .A(n17817), .B(n17818), .Z(n17815) );
  XNOR U22306 ( .A(y[1537]), .B(x[1537]), .Z(n17818) );
  XNOR U22307 ( .A(y[1538]), .B(x[1538]), .Z(n17817) );
  XNOR U22308 ( .A(n17808), .B(n17807), .Z(n17811) );
  XNOR U22309 ( .A(n17803), .B(n17804), .Z(n17807) );
  XNOR U22310 ( .A(y[1533]), .B(x[1533]), .Z(n17804) );
  XNOR U22311 ( .A(n17805), .B(n17806), .Z(n17803) );
  XNOR U22312 ( .A(y[1534]), .B(x[1534]), .Z(n17806) );
  XNOR U22313 ( .A(y[1535]), .B(x[1535]), .Z(n17805) );
  XNOR U22314 ( .A(n17797), .B(n17798), .Z(n17808) );
  XNOR U22315 ( .A(y[1530]), .B(x[1530]), .Z(n17798) );
  XNOR U22316 ( .A(n17799), .B(n17800), .Z(n17797) );
  XNOR U22317 ( .A(y[1531]), .B(x[1531]), .Z(n17800) );
  XNOR U22318 ( .A(y[1532]), .B(x[1532]), .Z(n17799) );
  XOR U22319 ( .A(n17773), .B(n17774), .Z(n17792) );
  XNOR U22320 ( .A(n17789), .B(n17790), .Z(n17774) );
  XNOR U22321 ( .A(n17784), .B(n17785), .Z(n17790) );
  XNOR U22322 ( .A(n17786), .B(n17787), .Z(n17785) );
  XNOR U22323 ( .A(y[1528]), .B(x[1528]), .Z(n17787) );
  XNOR U22324 ( .A(y[1529]), .B(x[1529]), .Z(n17786) );
  XNOR U22325 ( .A(y[1527]), .B(x[1527]), .Z(n17784) );
  XNOR U22326 ( .A(n17778), .B(n17779), .Z(n17789) );
  XNOR U22327 ( .A(y[1524]), .B(x[1524]), .Z(n17779) );
  XNOR U22328 ( .A(n17780), .B(n17781), .Z(n17778) );
  XNOR U22329 ( .A(y[1525]), .B(x[1525]), .Z(n17781) );
  XNOR U22330 ( .A(y[1526]), .B(x[1526]), .Z(n17780) );
  XOR U22331 ( .A(n17772), .B(n17771), .Z(n17773) );
  XNOR U22332 ( .A(n17767), .B(n17768), .Z(n17771) );
  XNOR U22333 ( .A(y[1521]), .B(x[1521]), .Z(n17768) );
  XNOR U22334 ( .A(n17769), .B(n17770), .Z(n17767) );
  XNOR U22335 ( .A(y[1522]), .B(x[1522]), .Z(n17770) );
  XNOR U22336 ( .A(y[1523]), .B(x[1523]), .Z(n17769) );
  XNOR U22337 ( .A(n17761), .B(n17762), .Z(n17772) );
  XNOR U22338 ( .A(y[1518]), .B(x[1518]), .Z(n17762) );
  XNOR U22339 ( .A(n17763), .B(n17764), .Z(n17761) );
  XNOR U22340 ( .A(y[1519]), .B(x[1519]), .Z(n17764) );
  XNOR U22341 ( .A(y[1520]), .B(x[1520]), .Z(n17763) );
  NAND U22342 ( .A(n17828), .B(n17829), .Z(N28689) );
  NANDN U22343 ( .A(n17830), .B(n17831), .Z(n17829) );
  OR U22344 ( .A(n17832), .B(n17833), .Z(n17831) );
  NAND U22345 ( .A(n17832), .B(n17833), .Z(n17828) );
  XOR U22346 ( .A(n17832), .B(n17834), .Z(N28688) );
  XNOR U22347 ( .A(n17830), .B(n17833), .Z(n17834) );
  AND U22348 ( .A(n17835), .B(n17836), .Z(n17833) );
  NANDN U22349 ( .A(n17837), .B(n17838), .Z(n17836) );
  NANDN U22350 ( .A(n17839), .B(n17840), .Z(n17838) );
  NANDN U22351 ( .A(n17840), .B(n17839), .Z(n17835) );
  NAND U22352 ( .A(n17841), .B(n17842), .Z(n17830) );
  NANDN U22353 ( .A(n17843), .B(n17844), .Z(n17842) );
  OR U22354 ( .A(n17845), .B(n17846), .Z(n17844) );
  NAND U22355 ( .A(n17846), .B(n17845), .Z(n17841) );
  AND U22356 ( .A(n17847), .B(n17848), .Z(n17832) );
  NANDN U22357 ( .A(n17849), .B(n17850), .Z(n17848) );
  NANDN U22358 ( .A(n17851), .B(n17852), .Z(n17850) );
  NANDN U22359 ( .A(n17852), .B(n17851), .Z(n17847) );
  XOR U22360 ( .A(n17846), .B(n17853), .Z(N28687) );
  XOR U22361 ( .A(n17843), .B(n17845), .Z(n17853) );
  XNOR U22362 ( .A(n17839), .B(n17854), .Z(n17845) );
  XNOR U22363 ( .A(n17837), .B(n17840), .Z(n17854) );
  NAND U22364 ( .A(n17855), .B(n17856), .Z(n17840) );
  NAND U22365 ( .A(n17857), .B(n17858), .Z(n17856) );
  OR U22366 ( .A(n17859), .B(n17860), .Z(n17857) );
  NANDN U22367 ( .A(n17861), .B(n17859), .Z(n17855) );
  IV U22368 ( .A(n17860), .Z(n17861) );
  NAND U22369 ( .A(n17862), .B(n17863), .Z(n17837) );
  NAND U22370 ( .A(n17864), .B(n17865), .Z(n17863) );
  NANDN U22371 ( .A(n17866), .B(n17867), .Z(n17864) );
  NANDN U22372 ( .A(n17867), .B(n17866), .Z(n17862) );
  AND U22373 ( .A(n17868), .B(n17869), .Z(n17839) );
  NAND U22374 ( .A(n17870), .B(n17871), .Z(n17869) );
  OR U22375 ( .A(n17872), .B(n17873), .Z(n17870) );
  NANDN U22376 ( .A(n17874), .B(n17872), .Z(n17868) );
  NAND U22377 ( .A(n17875), .B(n17876), .Z(n17843) );
  NANDN U22378 ( .A(n17877), .B(n17878), .Z(n17876) );
  OR U22379 ( .A(n17879), .B(n17880), .Z(n17878) );
  NANDN U22380 ( .A(n17881), .B(n17879), .Z(n17875) );
  IV U22381 ( .A(n17880), .Z(n17881) );
  XNOR U22382 ( .A(n17851), .B(n17882), .Z(n17846) );
  XNOR U22383 ( .A(n17849), .B(n17852), .Z(n17882) );
  NAND U22384 ( .A(n17883), .B(n17884), .Z(n17852) );
  NAND U22385 ( .A(n17885), .B(n17886), .Z(n17884) );
  OR U22386 ( .A(n17887), .B(n17888), .Z(n17885) );
  NANDN U22387 ( .A(n17889), .B(n17887), .Z(n17883) );
  IV U22388 ( .A(n17888), .Z(n17889) );
  NAND U22389 ( .A(n17890), .B(n17891), .Z(n17849) );
  NAND U22390 ( .A(n17892), .B(n17893), .Z(n17891) );
  NANDN U22391 ( .A(n17894), .B(n17895), .Z(n17892) );
  NANDN U22392 ( .A(n17895), .B(n17894), .Z(n17890) );
  AND U22393 ( .A(n17896), .B(n17897), .Z(n17851) );
  NAND U22394 ( .A(n17898), .B(n17899), .Z(n17897) );
  OR U22395 ( .A(n17900), .B(n17901), .Z(n17898) );
  NANDN U22396 ( .A(n17902), .B(n17900), .Z(n17896) );
  XNOR U22397 ( .A(n17877), .B(n17903), .Z(N28686) );
  XOR U22398 ( .A(n17879), .B(n17880), .Z(n17903) );
  XNOR U22399 ( .A(n17893), .B(n17904), .Z(n17880) );
  XOR U22400 ( .A(n17894), .B(n17895), .Z(n17904) );
  XOR U22401 ( .A(n17900), .B(n17905), .Z(n17895) );
  XOR U22402 ( .A(n17899), .B(n17902), .Z(n17905) );
  IV U22403 ( .A(n17901), .Z(n17902) );
  NAND U22404 ( .A(n17906), .B(n17907), .Z(n17901) );
  OR U22405 ( .A(n17908), .B(n17909), .Z(n17907) );
  OR U22406 ( .A(n17910), .B(n17911), .Z(n17906) );
  NAND U22407 ( .A(n17912), .B(n17913), .Z(n17899) );
  OR U22408 ( .A(n17914), .B(n17915), .Z(n17913) );
  OR U22409 ( .A(n17916), .B(n17917), .Z(n17912) );
  NOR U22410 ( .A(n17918), .B(n17919), .Z(n17900) );
  ANDN U22411 ( .B(n17920), .A(n17921), .Z(n17894) );
  XNOR U22412 ( .A(n17887), .B(n17922), .Z(n17893) );
  XNOR U22413 ( .A(n17886), .B(n17888), .Z(n17922) );
  NAND U22414 ( .A(n17923), .B(n17924), .Z(n17888) );
  OR U22415 ( .A(n17925), .B(n17926), .Z(n17924) );
  OR U22416 ( .A(n17927), .B(n17928), .Z(n17923) );
  NAND U22417 ( .A(n17929), .B(n17930), .Z(n17886) );
  OR U22418 ( .A(n17931), .B(n17932), .Z(n17930) );
  OR U22419 ( .A(n17933), .B(n17934), .Z(n17929) );
  ANDN U22420 ( .B(n17935), .A(n17936), .Z(n17887) );
  IV U22421 ( .A(n17937), .Z(n17935) );
  ANDN U22422 ( .B(n17938), .A(n17939), .Z(n17879) );
  XOR U22423 ( .A(n17865), .B(n17940), .Z(n17877) );
  XOR U22424 ( .A(n17866), .B(n17867), .Z(n17940) );
  XOR U22425 ( .A(n17872), .B(n17941), .Z(n17867) );
  XOR U22426 ( .A(n17871), .B(n17874), .Z(n17941) );
  IV U22427 ( .A(n17873), .Z(n17874) );
  NAND U22428 ( .A(n17942), .B(n17943), .Z(n17873) );
  OR U22429 ( .A(n17944), .B(n17945), .Z(n17943) );
  OR U22430 ( .A(n17946), .B(n17947), .Z(n17942) );
  NAND U22431 ( .A(n17948), .B(n17949), .Z(n17871) );
  OR U22432 ( .A(n17950), .B(n17951), .Z(n17949) );
  OR U22433 ( .A(n17952), .B(n17953), .Z(n17948) );
  NOR U22434 ( .A(n17954), .B(n17955), .Z(n17872) );
  ANDN U22435 ( .B(n17956), .A(n17957), .Z(n17866) );
  IV U22436 ( .A(n17958), .Z(n17956) );
  XNOR U22437 ( .A(n17859), .B(n17959), .Z(n17865) );
  XNOR U22438 ( .A(n17858), .B(n17860), .Z(n17959) );
  NAND U22439 ( .A(n17960), .B(n17961), .Z(n17860) );
  OR U22440 ( .A(n17962), .B(n17963), .Z(n17961) );
  OR U22441 ( .A(n17964), .B(n17965), .Z(n17960) );
  NAND U22442 ( .A(n17966), .B(n17967), .Z(n17858) );
  OR U22443 ( .A(n17968), .B(n17969), .Z(n17967) );
  OR U22444 ( .A(n17970), .B(n17971), .Z(n17966) );
  ANDN U22445 ( .B(n17972), .A(n17973), .Z(n17859) );
  IV U22446 ( .A(n17974), .Z(n17972) );
  XNOR U22447 ( .A(n17939), .B(n17938), .Z(N28685) );
  XOR U22448 ( .A(n17958), .B(n17957), .Z(n17938) );
  XNOR U22449 ( .A(n17973), .B(n17974), .Z(n17957) );
  XNOR U22450 ( .A(n17968), .B(n17969), .Z(n17974) );
  XNOR U22451 ( .A(n17970), .B(n17971), .Z(n17969) );
  XNOR U22452 ( .A(y[1516]), .B(x[1516]), .Z(n17971) );
  XNOR U22453 ( .A(y[1517]), .B(x[1517]), .Z(n17970) );
  XNOR U22454 ( .A(y[1515]), .B(x[1515]), .Z(n17968) );
  XNOR U22455 ( .A(n17962), .B(n17963), .Z(n17973) );
  XNOR U22456 ( .A(y[1512]), .B(x[1512]), .Z(n17963) );
  XNOR U22457 ( .A(n17964), .B(n17965), .Z(n17962) );
  XNOR U22458 ( .A(y[1513]), .B(x[1513]), .Z(n17965) );
  XNOR U22459 ( .A(y[1514]), .B(x[1514]), .Z(n17964) );
  XNOR U22460 ( .A(n17955), .B(n17954), .Z(n17958) );
  XNOR U22461 ( .A(n17950), .B(n17951), .Z(n17954) );
  XNOR U22462 ( .A(y[1509]), .B(x[1509]), .Z(n17951) );
  XNOR U22463 ( .A(n17952), .B(n17953), .Z(n17950) );
  XNOR U22464 ( .A(y[1510]), .B(x[1510]), .Z(n17953) );
  XNOR U22465 ( .A(y[1511]), .B(x[1511]), .Z(n17952) );
  XNOR U22466 ( .A(n17944), .B(n17945), .Z(n17955) );
  XNOR U22467 ( .A(y[1506]), .B(x[1506]), .Z(n17945) );
  XNOR U22468 ( .A(n17946), .B(n17947), .Z(n17944) );
  XNOR U22469 ( .A(y[1507]), .B(x[1507]), .Z(n17947) );
  XNOR U22470 ( .A(y[1508]), .B(x[1508]), .Z(n17946) );
  XOR U22471 ( .A(n17920), .B(n17921), .Z(n17939) );
  XNOR U22472 ( .A(n17936), .B(n17937), .Z(n17921) );
  XNOR U22473 ( .A(n17931), .B(n17932), .Z(n17937) );
  XNOR U22474 ( .A(n17933), .B(n17934), .Z(n17932) );
  XNOR U22475 ( .A(y[1504]), .B(x[1504]), .Z(n17934) );
  XNOR U22476 ( .A(y[1505]), .B(x[1505]), .Z(n17933) );
  XNOR U22477 ( .A(y[1503]), .B(x[1503]), .Z(n17931) );
  XNOR U22478 ( .A(n17925), .B(n17926), .Z(n17936) );
  XNOR U22479 ( .A(y[1500]), .B(x[1500]), .Z(n17926) );
  XNOR U22480 ( .A(n17927), .B(n17928), .Z(n17925) );
  XNOR U22481 ( .A(y[1501]), .B(x[1501]), .Z(n17928) );
  XNOR U22482 ( .A(y[1502]), .B(x[1502]), .Z(n17927) );
  XOR U22483 ( .A(n17919), .B(n17918), .Z(n17920) );
  XNOR U22484 ( .A(n17914), .B(n17915), .Z(n17918) );
  XNOR U22485 ( .A(y[1497]), .B(x[1497]), .Z(n17915) );
  XNOR U22486 ( .A(n17916), .B(n17917), .Z(n17914) );
  XNOR U22487 ( .A(y[1498]), .B(x[1498]), .Z(n17917) );
  XNOR U22488 ( .A(y[1499]), .B(x[1499]), .Z(n17916) );
  XNOR U22489 ( .A(n17908), .B(n17909), .Z(n17919) );
  XNOR U22490 ( .A(y[1494]), .B(x[1494]), .Z(n17909) );
  XNOR U22491 ( .A(n17910), .B(n17911), .Z(n17908) );
  XNOR U22492 ( .A(y[1495]), .B(x[1495]), .Z(n17911) );
  XNOR U22493 ( .A(y[1496]), .B(x[1496]), .Z(n17910) );
  NAND U22494 ( .A(n17975), .B(n17976), .Z(N28677) );
  NANDN U22495 ( .A(n17977), .B(n17978), .Z(n17976) );
  OR U22496 ( .A(n17979), .B(n17980), .Z(n17978) );
  NAND U22497 ( .A(n17979), .B(n17980), .Z(n17975) );
  XOR U22498 ( .A(n17979), .B(n17981), .Z(N28676) );
  XNOR U22499 ( .A(n17977), .B(n17980), .Z(n17981) );
  AND U22500 ( .A(n17982), .B(n17983), .Z(n17980) );
  NANDN U22501 ( .A(n17984), .B(n17985), .Z(n17983) );
  NANDN U22502 ( .A(n17986), .B(n17987), .Z(n17985) );
  NANDN U22503 ( .A(n17987), .B(n17986), .Z(n17982) );
  NAND U22504 ( .A(n17988), .B(n17989), .Z(n17977) );
  NANDN U22505 ( .A(n17990), .B(n17991), .Z(n17989) );
  OR U22506 ( .A(n17992), .B(n17993), .Z(n17991) );
  NAND U22507 ( .A(n17993), .B(n17992), .Z(n17988) );
  AND U22508 ( .A(n17994), .B(n17995), .Z(n17979) );
  NANDN U22509 ( .A(n17996), .B(n17997), .Z(n17995) );
  NANDN U22510 ( .A(n17998), .B(n17999), .Z(n17997) );
  NANDN U22511 ( .A(n17999), .B(n17998), .Z(n17994) );
  XOR U22512 ( .A(n17993), .B(n18000), .Z(N28675) );
  XOR U22513 ( .A(n17990), .B(n17992), .Z(n18000) );
  XNOR U22514 ( .A(n17986), .B(n18001), .Z(n17992) );
  XNOR U22515 ( .A(n17984), .B(n17987), .Z(n18001) );
  NAND U22516 ( .A(n18002), .B(n18003), .Z(n17987) );
  NAND U22517 ( .A(n18004), .B(n18005), .Z(n18003) );
  OR U22518 ( .A(n18006), .B(n18007), .Z(n18004) );
  NANDN U22519 ( .A(n18008), .B(n18006), .Z(n18002) );
  IV U22520 ( .A(n18007), .Z(n18008) );
  NAND U22521 ( .A(n18009), .B(n18010), .Z(n17984) );
  NAND U22522 ( .A(n18011), .B(n18012), .Z(n18010) );
  NANDN U22523 ( .A(n18013), .B(n18014), .Z(n18011) );
  NANDN U22524 ( .A(n18014), .B(n18013), .Z(n18009) );
  AND U22525 ( .A(n18015), .B(n18016), .Z(n17986) );
  NAND U22526 ( .A(n18017), .B(n18018), .Z(n18016) );
  OR U22527 ( .A(n18019), .B(n18020), .Z(n18017) );
  NANDN U22528 ( .A(n18021), .B(n18019), .Z(n18015) );
  NAND U22529 ( .A(n18022), .B(n18023), .Z(n17990) );
  NANDN U22530 ( .A(n18024), .B(n18025), .Z(n18023) );
  OR U22531 ( .A(n18026), .B(n18027), .Z(n18025) );
  NANDN U22532 ( .A(n18028), .B(n18026), .Z(n18022) );
  IV U22533 ( .A(n18027), .Z(n18028) );
  XNOR U22534 ( .A(n17998), .B(n18029), .Z(n17993) );
  XNOR U22535 ( .A(n17996), .B(n17999), .Z(n18029) );
  NAND U22536 ( .A(n18030), .B(n18031), .Z(n17999) );
  NAND U22537 ( .A(n18032), .B(n18033), .Z(n18031) );
  OR U22538 ( .A(n18034), .B(n18035), .Z(n18032) );
  NANDN U22539 ( .A(n18036), .B(n18034), .Z(n18030) );
  IV U22540 ( .A(n18035), .Z(n18036) );
  NAND U22541 ( .A(n18037), .B(n18038), .Z(n17996) );
  NAND U22542 ( .A(n18039), .B(n18040), .Z(n18038) );
  NANDN U22543 ( .A(n18041), .B(n18042), .Z(n18039) );
  NANDN U22544 ( .A(n18042), .B(n18041), .Z(n18037) );
  AND U22545 ( .A(n18043), .B(n18044), .Z(n17998) );
  NAND U22546 ( .A(n18045), .B(n18046), .Z(n18044) );
  OR U22547 ( .A(n18047), .B(n18048), .Z(n18045) );
  NANDN U22548 ( .A(n18049), .B(n18047), .Z(n18043) );
  XNOR U22549 ( .A(n18024), .B(n18050), .Z(N28674) );
  XOR U22550 ( .A(n18026), .B(n18027), .Z(n18050) );
  XNOR U22551 ( .A(n18040), .B(n18051), .Z(n18027) );
  XOR U22552 ( .A(n18041), .B(n18042), .Z(n18051) );
  XOR U22553 ( .A(n18047), .B(n18052), .Z(n18042) );
  XOR U22554 ( .A(n18046), .B(n18049), .Z(n18052) );
  IV U22555 ( .A(n18048), .Z(n18049) );
  NAND U22556 ( .A(n18053), .B(n18054), .Z(n18048) );
  OR U22557 ( .A(n18055), .B(n18056), .Z(n18054) );
  OR U22558 ( .A(n18057), .B(n18058), .Z(n18053) );
  NAND U22559 ( .A(n18059), .B(n18060), .Z(n18046) );
  OR U22560 ( .A(n18061), .B(n18062), .Z(n18060) );
  OR U22561 ( .A(n18063), .B(n18064), .Z(n18059) );
  NOR U22562 ( .A(n18065), .B(n18066), .Z(n18047) );
  ANDN U22563 ( .B(n18067), .A(n18068), .Z(n18041) );
  XNOR U22564 ( .A(n18034), .B(n18069), .Z(n18040) );
  XNOR U22565 ( .A(n18033), .B(n18035), .Z(n18069) );
  NAND U22566 ( .A(n18070), .B(n18071), .Z(n18035) );
  OR U22567 ( .A(n18072), .B(n18073), .Z(n18071) );
  OR U22568 ( .A(n18074), .B(n18075), .Z(n18070) );
  NAND U22569 ( .A(n18076), .B(n18077), .Z(n18033) );
  OR U22570 ( .A(n18078), .B(n18079), .Z(n18077) );
  OR U22571 ( .A(n18080), .B(n18081), .Z(n18076) );
  ANDN U22572 ( .B(n18082), .A(n18083), .Z(n18034) );
  IV U22573 ( .A(n18084), .Z(n18082) );
  ANDN U22574 ( .B(n18085), .A(n18086), .Z(n18026) );
  XOR U22575 ( .A(n18012), .B(n18087), .Z(n18024) );
  XOR U22576 ( .A(n18013), .B(n18014), .Z(n18087) );
  XOR U22577 ( .A(n18019), .B(n18088), .Z(n18014) );
  XOR U22578 ( .A(n18018), .B(n18021), .Z(n18088) );
  IV U22579 ( .A(n18020), .Z(n18021) );
  NAND U22580 ( .A(n18089), .B(n18090), .Z(n18020) );
  OR U22581 ( .A(n18091), .B(n18092), .Z(n18090) );
  OR U22582 ( .A(n18093), .B(n18094), .Z(n18089) );
  NAND U22583 ( .A(n18095), .B(n18096), .Z(n18018) );
  OR U22584 ( .A(n18097), .B(n18098), .Z(n18096) );
  OR U22585 ( .A(n18099), .B(n18100), .Z(n18095) );
  NOR U22586 ( .A(n18101), .B(n18102), .Z(n18019) );
  ANDN U22587 ( .B(n18103), .A(n18104), .Z(n18013) );
  IV U22588 ( .A(n18105), .Z(n18103) );
  XNOR U22589 ( .A(n18006), .B(n18106), .Z(n18012) );
  XNOR U22590 ( .A(n18005), .B(n18007), .Z(n18106) );
  NAND U22591 ( .A(n18107), .B(n18108), .Z(n18007) );
  OR U22592 ( .A(n18109), .B(n18110), .Z(n18108) );
  OR U22593 ( .A(n18111), .B(n18112), .Z(n18107) );
  NAND U22594 ( .A(n18113), .B(n18114), .Z(n18005) );
  OR U22595 ( .A(n18115), .B(n18116), .Z(n18114) );
  OR U22596 ( .A(n18117), .B(n18118), .Z(n18113) );
  ANDN U22597 ( .B(n18119), .A(n18120), .Z(n18006) );
  IV U22598 ( .A(n18121), .Z(n18119) );
  XNOR U22599 ( .A(n18086), .B(n18085), .Z(N28673) );
  XOR U22600 ( .A(n18105), .B(n18104), .Z(n18085) );
  XNOR U22601 ( .A(n18120), .B(n18121), .Z(n18104) );
  XNOR U22602 ( .A(n18115), .B(n18116), .Z(n18121) );
  XNOR U22603 ( .A(n18117), .B(n18118), .Z(n18116) );
  XNOR U22604 ( .A(y[1492]), .B(x[1492]), .Z(n18118) );
  XNOR U22605 ( .A(y[1493]), .B(x[1493]), .Z(n18117) );
  XNOR U22606 ( .A(y[1491]), .B(x[1491]), .Z(n18115) );
  XNOR U22607 ( .A(n18109), .B(n18110), .Z(n18120) );
  XNOR U22608 ( .A(y[1488]), .B(x[1488]), .Z(n18110) );
  XNOR U22609 ( .A(n18111), .B(n18112), .Z(n18109) );
  XNOR U22610 ( .A(y[1489]), .B(x[1489]), .Z(n18112) );
  XNOR U22611 ( .A(y[1490]), .B(x[1490]), .Z(n18111) );
  XNOR U22612 ( .A(n18102), .B(n18101), .Z(n18105) );
  XNOR U22613 ( .A(n18097), .B(n18098), .Z(n18101) );
  XNOR U22614 ( .A(y[1485]), .B(x[1485]), .Z(n18098) );
  XNOR U22615 ( .A(n18099), .B(n18100), .Z(n18097) );
  XNOR U22616 ( .A(y[1486]), .B(x[1486]), .Z(n18100) );
  XNOR U22617 ( .A(y[1487]), .B(x[1487]), .Z(n18099) );
  XNOR U22618 ( .A(n18091), .B(n18092), .Z(n18102) );
  XNOR U22619 ( .A(y[1482]), .B(x[1482]), .Z(n18092) );
  XNOR U22620 ( .A(n18093), .B(n18094), .Z(n18091) );
  XNOR U22621 ( .A(y[1483]), .B(x[1483]), .Z(n18094) );
  XNOR U22622 ( .A(y[1484]), .B(x[1484]), .Z(n18093) );
  XOR U22623 ( .A(n18067), .B(n18068), .Z(n18086) );
  XNOR U22624 ( .A(n18083), .B(n18084), .Z(n18068) );
  XNOR U22625 ( .A(n18078), .B(n18079), .Z(n18084) );
  XNOR U22626 ( .A(n18080), .B(n18081), .Z(n18079) );
  XNOR U22627 ( .A(y[1480]), .B(x[1480]), .Z(n18081) );
  XNOR U22628 ( .A(y[1481]), .B(x[1481]), .Z(n18080) );
  XNOR U22629 ( .A(y[1479]), .B(x[1479]), .Z(n18078) );
  XNOR U22630 ( .A(n18072), .B(n18073), .Z(n18083) );
  XNOR U22631 ( .A(y[1476]), .B(x[1476]), .Z(n18073) );
  XNOR U22632 ( .A(n18074), .B(n18075), .Z(n18072) );
  XNOR U22633 ( .A(y[1477]), .B(x[1477]), .Z(n18075) );
  XNOR U22634 ( .A(y[1478]), .B(x[1478]), .Z(n18074) );
  XOR U22635 ( .A(n18066), .B(n18065), .Z(n18067) );
  XNOR U22636 ( .A(n18061), .B(n18062), .Z(n18065) );
  XNOR U22637 ( .A(y[1473]), .B(x[1473]), .Z(n18062) );
  XNOR U22638 ( .A(n18063), .B(n18064), .Z(n18061) );
  XNOR U22639 ( .A(y[1474]), .B(x[1474]), .Z(n18064) );
  XNOR U22640 ( .A(y[1475]), .B(x[1475]), .Z(n18063) );
  XNOR U22641 ( .A(n18055), .B(n18056), .Z(n18066) );
  XNOR U22642 ( .A(y[1470]), .B(x[1470]), .Z(n18056) );
  XNOR U22643 ( .A(n18057), .B(n18058), .Z(n18055) );
  XNOR U22644 ( .A(y[1471]), .B(x[1471]), .Z(n18058) );
  XNOR U22645 ( .A(y[1472]), .B(x[1472]), .Z(n18057) );
  NAND U22646 ( .A(n18122), .B(n18123), .Z(N28665) );
  NANDN U22647 ( .A(n18124), .B(n18125), .Z(n18123) );
  OR U22648 ( .A(n18126), .B(n18127), .Z(n18125) );
  NAND U22649 ( .A(n18126), .B(n18127), .Z(n18122) );
  XOR U22650 ( .A(n18126), .B(n18128), .Z(N28664) );
  XNOR U22651 ( .A(n18124), .B(n18127), .Z(n18128) );
  AND U22652 ( .A(n18129), .B(n18130), .Z(n18127) );
  NANDN U22653 ( .A(n18131), .B(n18132), .Z(n18130) );
  NANDN U22654 ( .A(n18133), .B(n18134), .Z(n18132) );
  NANDN U22655 ( .A(n18134), .B(n18133), .Z(n18129) );
  NAND U22656 ( .A(n18135), .B(n18136), .Z(n18124) );
  NANDN U22657 ( .A(n18137), .B(n18138), .Z(n18136) );
  OR U22658 ( .A(n18139), .B(n18140), .Z(n18138) );
  NAND U22659 ( .A(n18140), .B(n18139), .Z(n18135) );
  AND U22660 ( .A(n18141), .B(n18142), .Z(n18126) );
  NANDN U22661 ( .A(n18143), .B(n18144), .Z(n18142) );
  NANDN U22662 ( .A(n18145), .B(n18146), .Z(n18144) );
  NANDN U22663 ( .A(n18146), .B(n18145), .Z(n18141) );
  XOR U22664 ( .A(n18140), .B(n18147), .Z(N28663) );
  XOR U22665 ( .A(n18137), .B(n18139), .Z(n18147) );
  XNOR U22666 ( .A(n18133), .B(n18148), .Z(n18139) );
  XNOR U22667 ( .A(n18131), .B(n18134), .Z(n18148) );
  NAND U22668 ( .A(n18149), .B(n18150), .Z(n18134) );
  NAND U22669 ( .A(n18151), .B(n18152), .Z(n18150) );
  OR U22670 ( .A(n18153), .B(n18154), .Z(n18151) );
  NANDN U22671 ( .A(n18155), .B(n18153), .Z(n18149) );
  IV U22672 ( .A(n18154), .Z(n18155) );
  NAND U22673 ( .A(n18156), .B(n18157), .Z(n18131) );
  NAND U22674 ( .A(n18158), .B(n18159), .Z(n18157) );
  NANDN U22675 ( .A(n18160), .B(n18161), .Z(n18158) );
  NANDN U22676 ( .A(n18161), .B(n18160), .Z(n18156) );
  AND U22677 ( .A(n18162), .B(n18163), .Z(n18133) );
  NAND U22678 ( .A(n18164), .B(n18165), .Z(n18163) );
  OR U22679 ( .A(n18166), .B(n18167), .Z(n18164) );
  NANDN U22680 ( .A(n18168), .B(n18166), .Z(n18162) );
  NAND U22681 ( .A(n18169), .B(n18170), .Z(n18137) );
  NANDN U22682 ( .A(n18171), .B(n18172), .Z(n18170) );
  OR U22683 ( .A(n18173), .B(n18174), .Z(n18172) );
  NANDN U22684 ( .A(n18175), .B(n18173), .Z(n18169) );
  IV U22685 ( .A(n18174), .Z(n18175) );
  XNOR U22686 ( .A(n18145), .B(n18176), .Z(n18140) );
  XNOR U22687 ( .A(n18143), .B(n18146), .Z(n18176) );
  NAND U22688 ( .A(n18177), .B(n18178), .Z(n18146) );
  NAND U22689 ( .A(n18179), .B(n18180), .Z(n18178) );
  OR U22690 ( .A(n18181), .B(n18182), .Z(n18179) );
  NANDN U22691 ( .A(n18183), .B(n18181), .Z(n18177) );
  IV U22692 ( .A(n18182), .Z(n18183) );
  NAND U22693 ( .A(n18184), .B(n18185), .Z(n18143) );
  NAND U22694 ( .A(n18186), .B(n18187), .Z(n18185) );
  NANDN U22695 ( .A(n18188), .B(n18189), .Z(n18186) );
  NANDN U22696 ( .A(n18189), .B(n18188), .Z(n18184) );
  AND U22697 ( .A(n18190), .B(n18191), .Z(n18145) );
  NAND U22698 ( .A(n18192), .B(n18193), .Z(n18191) );
  OR U22699 ( .A(n18194), .B(n18195), .Z(n18192) );
  NANDN U22700 ( .A(n18196), .B(n18194), .Z(n18190) );
  XNOR U22701 ( .A(n18171), .B(n18197), .Z(N28662) );
  XOR U22702 ( .A(n18173), .B(n18174), .Z(n18197) );
  XNOR U22703 ( .A(n18187), .B(n18198), .Z(n18174) );
  XOR U22704 ( .A(n18188), .B(n18189), .Z(n18198) );
  XOR U22705 ( .A(n18194), .B(n18199), .Z(n18189) );
  XOR U22706 ( .A(n18193), .B(n18196), .Z(n18199) );
  IV U22707 ( .A(n18195), .Z(n18196) );
  NAND U22708 ( .A(n18200), .B(n18201), .Z(n18195) );
  OR U22709 ( .A(n18202), .B(n18203), .Z(n18201) );
  OR U22710 ( .A(n18204), .B(n18205), .Z(n18200) );
  NAND U22711 ( .A(n18206), .B(n18207), .Z(n18193) );
  OR U22712 ( .A(n18208), .B(n18209), .Z(n18207) );
  OR U22713 ( .A(n18210), .B(n18211), .Z(n18206) );
  NOR U22714 ( .A(n18212), .B(n18213), .Z(n18194) );
  ANDN U22715 ( .B(n18214), .A(n18215), .Z(n18188) );
  XNOR U22716 ( .A(n18181), .B(n18216), .Z(n18187) );
  XNOR U22717 ( .A(n18180), .B(n18182), .Z(n18216) );
  NAND U22718 ( .A(n18217), .B(n18218), .Z(n18182) );
  OR U22719 ( .A(n18219), .B(n18220), .Z(n18218) );
  OR U22720 ( .A(n18221), .B(n18222), .Z(n18217) );
  NAND U22721 ( .A(n18223), .B(n18224), .Z(n18180) );
  OR U22722 ( .A(n18225), .B(n18226), .Z(n18224) );
  OR U22723 ( .A(n18227), .B(n18228), .Z(n18223) );
  ANDN U22724 ( .B(n18229), .A(n18230), .Z(n18181) );
  IV U22725 ( .A(n18231), .Z(n18229) );
  ANDN U22726 ( .B(n18232), .A(n18233), .Z(n18173) );
  XOR U22727 ( .A(n18159), .B(n18234), .Z(n18171) );
  XOR U22728 ( .A(n18160), .B(n18161), .Z(n18234) );
  XOR U22729 ( .A(n18166), .B(n18235), .Z(n18161) );
  XOR U22730 ( .A(n18165), .B(n18168), .Z(n18235) );
  IV U22731 ( .A(n18167), .Z(n18168) );
  NAND U22732 ( .A(n18236), .B(n18237), .Z(n18167) );
  OR U22733 ( .A(n18238), .B(n18239), .Z(n18237) );
  OR U22734 ( .A(n18240), .B(n18241), .Z(n18236) );
  NAND U22735 ( .A(n18242), .B(n18243), .Z(n18165) );
  OR U22736 ( .A(n18244), .B(n18245), .Z(n18243) );
  OR U22737 ( .A(n18246), .B(n18247), .Z(n18242) );
  NOR U22738 ( .A(n18248), .B(n18249), .Z(n18166) );
  ANDN U22739 ( .B(n18250), .A(n18251), .Z(n18160) );
  IV U22740 ( .A(n18252), .Z(n18250) );
  XNOR U22741 ( .A(n18153), .B(n18253), .Z(n18159) );
  XNOR U22742 ( .A(n18152), .B(n18154), .Z(n18253) );
  NAND U22743 ( .A(n18254), .B(n18255), .Z(n18154) );
  OR U22744 ( .A(n18256), .B(n18257), .Z(n18255) );
  OR U22745 ( .A(n18258), .B(n18259), .Z(n18254) );
  NAND U22746 ( .A(n18260), .B(n18261), .Z(n18152) );
  OR U22747 ( .A(n18262), .B(n18263), .Z(n18261) );
  OR U22748 ( .A(n18264), .B(n18265), .Z(n18260) );
  ANDN U22749 ( .B(n18266), .A(n18267), .Z(n18153) );
  IV U22750 ( .A(n18268), .Z(n18266) );
  XNOR U22751 ( .A(n18233), .B(n18232), .Z(N28661) );
  XOR U22752 ( .A(n18252), .B(n18251), .Z(n18232) );
  XNOR U22753 ( .A(n18267), .B(n18268), .Z(n18251) );
  XNOR U22754 ( .A(n18262), .B(n18263), .Z(n18268) );
  XNOR U22755 ( .A(n18264), .B(n18265), .Z(n18263) );
  XNOR U22756 ( .A(y[1468]), .B(x[1468]), .Z(n18265) );
  XNOR U22757 ( .A(y[1469]), .B(x[1469]), .Z(n18264) );
  XNOR U22758 ( .A(y[1467]), .B(x[1467]), .Z(n18262) );
  XNOR U22759 ( .A(n18256), .B(n18257), .Z(n18267) );
  XNOR U22760 ( .A(y[1464]), .B(x[1464]), .Z(n18257) );
  XNOR U22761 ( .A(n18258), .B(n18259), .Z(n18256) );
  XNOR U22762 ( .A(y[1465]), .B(x[1465]), .Z(n18259) );
  XNOR U22763 ( .A(y[1466]), .B(x[1466]), .Z(n18258) );
  XNOR U22764 ( .A(n18249), .B(n18248), .Z(n18252) );
  XNOR U22765 ( .A(n18244), .B(n18245), .Z(n18248) );
  XNOR U22766 ( .A(y[1461]), .B(x[1461]), .Z(n18245) );
  XNOR U22767 ( .A(n18246), .B(n18247), .Z(n18244) );
  XNOR U22768 ( .A(y[1462]), .B(x[1462]), .Z(n18247) );
  XNOR U22769 ( .A(y[1463]), .B(x[1463]), .Z(n18246) );
  XNOR U22770 ( .A(n18238), .B(n18239), .Z(n18249) );
  XNOR U22771 ( .A(y[1458]), .B(x[1458]), .Z(n18239) );
  XNOR U22772 ( .A(n18240), .B(n18241), .Z(n18238) );
  XNOR U22773 ( .A(y[1459]), .B(x[1459]), .Z(n18241) );
  XNOR U22774 ( .A(y[1460]), .B(x[1460]), .Z(n18240) );
  XOR U22775 ( .A(n18214), .B(n18215), .Z(n18233) );
  XNOR U22776 ( .A(n18230), .B(n18231), .Z(n18215) );
  XNOR U22777 ( .A(n18225), .B(n18226), .Z(n18231) );
  XNOR U22778 ( .A(n18227), .B(n18228), .Z(n18226) );
  XNOR U22779 ( .A(y[1456]), .B(x[1456]), .Z(n18228) );
  XNOR U22780 ( .A(y[1457]), .B(x[1457]), .Z(n18227) );
  XNOR U22781 ( .A(y[1455]), .B(x[1455]), .Z(n18225) );
  XNOR U22782 ( .A(n18219), .B(n18220), .Z(n18230) );
  XNOR U22783 ( .A(y[1452]), .B(x[1452]), .Z(n18220) );
  XNOR U22784 ( .A(n18221), .B(n18222), .Z(n18219) );
  XNOR U22785 ( .A(y[1453]), .B(x[1453]), .Z(n18222) );
  XNOR U22786 ( .A(y[1454]), .B(x[1454]), .Z(n18221) );
  XOR U22787 ( .A(n18213), .B(n18212), .Z(n18214) );
  XNOR U22788 ( .A(n18208), .B(n18209), .Z(n18212) );
  XNOR U22789 ( .A(y[1449]), .B(x[1449]), .Z(n18209) );
  XNOR U22790 ( .A(n18210), .B(n18211), .Z(n18208) );
  XNOR U22791 ( .A(y[1450]), .B(x[1450]), .Z(n18211) );
  XNOR U22792 ( .A(y[1451]), .B(x[1451]), .Z(n18210) );
  XNOR U22793 ( .A(n18202), .B(n18203), .Z(n18213) );
  XNOR U22794 ( .A(y[1446]), .B(x[1446]), .Z(n18203) );
  XNOR U22795 ( .A(n18204), .B(n18205), .Z(n18202) );
  XNOR U22796 ( .A(y[1447]), .B(x[1447]), .Z(n18205) );
  XNOR U22797 ( .A(y[1448]), .B(x[1448]), .Z(n18204) );
  NAND U22798 ( .A(n18269), .B(n18270), .Z(N28653) );
  NANDN U22799 ( .A(n18271), .B(n18272), .Z(n18270) );
  OR U22800 ( .A(n18273), .B(n18274), .Z(n18272) );
  NAND U22801 ( .A(n18273), .B(n18274), .Z(n18269) );
  XOR U22802 ( .A(n18273), .B(n18275), .Z(N28652) );
  XNOR U22803 ( .A(n18271), .B(n18274), .Z(n18275) );
  AND U22804 ( .A(n18276), .B(n18277), .Z(n18274) );
  NANDN U22805 ( .A(n18278), .B(n18279), .Z(n18277) );
  NANDN U22806 ( .A(n18280), .B(n18281), .Z(n18279) );
  NANDN U22807 ( .A(n18281), .B(n18280), .Z(n18276) );
  NAND U22808 ( .A(n18282), .B(n18283), .Z(n18271) );
  NANDN U22809 ( .A(n18284), .B(n18285), .Z(n18283) );
  OR U22810 ( .A(n18286), .B(n18287), .Z(n18285) );
  NAND U22811 ( .A(n18287), .B(n18286), .Z(n18282) );
  AND U22812 ( .A(n18288), .B(n18289), .Z(n18273) );
  NANDN U22813 ( .A(n18290), .B(n18291), .Z(n18289) );
  NANDN U22814 ( .A(n18292), .B(n18293), .Z(n18291) );
  NANDN U22815 ( .A(n18293), .B(n18292), .Z(n18288) );
  XOR U22816 ( .A(n18287), .B(n18294), .Z(N28651) );
  XOR U22817 ( .A(n18284), .B(n18286), .Z(n18294) );
  XNOR U22818 ( .A(n18280), .B(n18295), .Z(n18286) );
  XNOR U22819 ( .A(n18278), .B(n18281), .Z(n18295) );
  NAND U22820 ( .A(n18296), .B(n18297), .Z(n18281) );
  NAND U22821 ( .A(n18298), .B(n18299), .Z(n18297) );
  OR U22822 ( .A(n18300), .B(n18301), .Z(n18298) );
  NANDN U22823 ( .A(n18302), .B(n18300), .Z(n18296) );
  IV U22824 ( .A(n18301), .Z(n18302) );
  NAND U22825 ( .A(n18303), .B(n18304), .Z(n18278) );
  NAND U22826 ( .A(n18305), .B(n18306), .Z(n18304) );
  NANDN U22827 ( .A(n18307), .B(n18308), .Z(n18305) );
  NANDN U22828 ( .A(n18308), .B(n18307), .Z(n18303) );
  AND U22829 ( .A(n18309), .B(n18310), .Z(n18280) );
  NAND U22830 ( .A(n18311), .B(n18312), .Z(n18310) );
  OR U22831 ( .A(n18313), .B(n18314), .Z(n18311) );
  NANDN U22832 ( .A(n18315), .B(n18313), .Z(n18309) );
  NAND U22833 ( .A(n18316), .B(n18317), .Z(n18284) );
  NANDN U22834 ( .A(n18318), .B(n18319), .Z(n18317) );
  OR U22835 ( .A(n18320), .B(n18321), .Z(n18319) );
  NANDN U22836 ( .A(n18322), .B(n18320), .Z(n18316) );
  IV U22837 ( .A(n18321), .Z(n18322) );
  XNOR U22838 ( .A(n18292), .B(n18323), .Z(n18287) );
  XNOR U22839 ( .A(n18290), .B(n18293), .Z(n18323) );
  NAND U22840 ( .A(n18324), .B(n18325), .Z(n18293) );
  NAND U22841 ( .A(n18326), .B(n18327), .Z(n18325) );
  OR U22842 ( .A(n18328), .B(n18329), .Z(n18326) );
  NANDN U22843 ( .A(n18330), .B(n18328), .Z(n18324) );
  IV U22844 ( .A(n18329), .Z(n18330) );
  NAND U22845 ( .A(n18331), .B(n18332), .Z(n18290) );
  NAND U22846 ( .A(n18333), .B(n18334), .Z(n18332) );
  NANDN U22847 ( .A(n18335), .B(n18336), .Z(n18333) );
  NANDN U22848 ( .A(n18336), .B(n18335), .Z(n18331) );
  AND U22849 ( .A(n18337), .B(n18338), .Z(n18292) );
  NAND U22850 ( .A(n18339), .B(n18340), .Z(n18338) );
  OR U22851 ( .A(n18341), .B(n18342), .Z(n18339) );
  NANDN U22852 ( .A(n18343), .B(n18341), .Z(n18337) );
  XNOR U22853 ( .A(n18318), .B(n18344), .Z(N28650) );
  XOR U22854 ( .A(n18320), .B(n18321), .Z(n18344) );
  XNOR U22855 ( .A(n18334), .B(n18345), .Z(n18321) );
  XOR U22856 ( .A(n18335), .B(n18336), .Z(n18345) );
  XOR U22857 ( .A(n18341), .B(n18346), .Z(n18336) );
  XOR U22858 ( .A(n18340), .B(n18343), .Z(n18346) );
  IV U22859 ( .A(n18342), .Z(n18343) );
  NAND U22860 ( .A(n18347), .B(n18348), .Z(n18342) );
  OR U22861 ( .A(n18349), .B(n18350), .Z(n18348) );
  OR U22862 ( .A(n18351), .B(n18352), .Z(n18347) );
  NAND U22863 ( .A(n18353), .B(n18354), .Z(n18340) );
  OR U22864 ( .A(n18355), .B(n18356), .Z(n18354) );
  OR U22865 ( .A(n18357), .B(n18358), .Z(n18353) );
  NOR U22866 ( .A(n18359), .B(n18360), .Z(n18341) );
  ANDN U22867 ( .B(n18361), .A(n18362), .Z(n18335) );
  XNOR U22868 ( .A(n18328), .B(n18363), .Z(n18334) );
  XNOR U22869 ( .A(n18327), .B(n18329), .Z(n18363) );
  NAND U22870 ( .A(n18364), .B(n18365), .Z(n18329) );
  OR U22871 ( .A(n18366), .B(n18367), .Z(n18365) );
  OR U22872 ( .A(n18368), .B(n18369), .Z(n18364) );
  NAND U22873 ( .A(n18370), .B(n18371), .Z(n18327) );
  OR U22874 ( .A(n18372), .B(n18373), .Z(n18371) );
  OR U22875 ( .A(n18374), .B(n18375), .Z(n18370) );
  ANDN U22876 ( .B(n18376), .A(n18377), .Z(n18328) );
  IV U22877 ( .A(n18378), .Z(n18376) );
  ANDN U22878 ( .B(n18379), .A(n18380), .Z(n18320) );
  XOR U22879 ( .A(n18306), .B(n18381), .Z(n18318) );
  XOR U22880 ( .A(n18307), .B(n18308), .Z(n18381) );
  XOR U22881 ( .A(n18313), .B(n18382), .Z(n18308) );
  XOR U22882 ( .A(n18312), .B(n18315), .Z(n18382) );
  IV U22883 ( .A(n18314), .Z(n18315) );
  NAND U22884 ( .A(n18383), .B(n18384), .Z(n18314) );
  OR U22885 ( .A(n18385), .B(n18386), .Z(n18384) );
  OR U22886 ( .A(n18387), .B(n18388), .Z(n18383) );
  NAND U22887 ( .A(n18389), .B(n18390), .Z(n18312) );
  OR U22888 ( .A(n18391), .B(n18392), .Z(n18390) );
  OR U22889 ( .A(n18393), .B(n18394), .Z(n18389) );
  NOR U22890 ( .A(n18395), .B(n18396), .Z(n18313) );
  ANDN U22891 ( .B(n18397), .A(n18398), .Z(n18307) );
  IV U22892 ( .A(n18399), .Z(n18397) );
  XNOR U22893 ( .A(n18300), .B(n18400), .Z(n18306) );
  XNOR U22894 ( .A(n18299), .B(n18301), .Z(n18400) );
  NAND U22895 ( .A(n18401), .B(n18402), .Z(n18301) );
  OR U22896 ( .A(n18403), .B(n18404), .Z(n18402) );
  OR U22897 ( .A(n18405), .B(n18406), .Z(n18401) );
  NAND U22898 ( .A(n18407), .B(n18408), .Z(n18299) );
  OR U22899 ( .A(n18409), .B(n18410), .Z(n18408) );
  OR U22900 ( .A(n18411), .B(n18412), .Z(n18407) );
  ANDN U22901 ( .B(n18413), .A(n18414), .Z(n18300) );
  IV U22902 ( .A(n18415), .Z(n18413) );
  XNOR U22903 ( .A(n18380), .B(n18379), .Z(N28649) );
  XOR U22904 ( .A(n18399), .B(n18398), .Z(n18379) );
  XNOR U22905 ( .A(n18414), .B(n18415), .Z(n18398) );
  XNOR U22906 ( .A(n18409), .B(n18410), .Z(n18415) );
  XNOR U22907 ( .A(n18411), .B(n18412), .Z(n18410) );
  XNOR U22908 ( .A(y[1444]), .B(x[1444]), .Z(n18412) );
  XNOR U22909 ( .A(y[1445]), .B(x[1445]), .Z(n18411) );
  XNOR U22910 ( .A(y[1443]), .B(x[1443]), .Z(n18409) );
  XNOR U22911 ( .A(n18403), .B(n18404), .Z(n18414) );
  XNOR U22912 ( .A(y[1440]), .B(x[1440]), .Z(n18404) );
  XNOR U22913 ( .A(n18405), .B(n18406), .Z(n18403) );
  XNOR U22914 ( .A(y[1441]), .B(x[1441]), .Z(n18406) );
  XNOR U22915 ( .A(y[1442]), .B(x[1442]), .Z(n18405) );
  XNOR U22916 ( .A(n18396), .B(n18395), .Z(n18399) );
  XNOR U22917 ( .A(n18391), .B(n18392), .Z(n18395) );
  XNOR U22918 ( .A(y[1437]), .B(x[1437]), .Z(n18392) );
  XNOR U22919 ( .A(n18393), .B(n18394), .Z(n18391) );
  XNOR U22920 ( .A(y[1438]), .B(x[1438]), .Z(n18394) );
  XNOR U22921 ( .A(y[1439]), .B(x[1439]), .Z(n18393) );
  XNOR U22922 ( .A(n18385), .B(n18386), .Z(n18396) );
  XNOR U22923 ( .A(y[1434]), .B(x[1434]), .Z(n18386) );
  XNOR U22924 ( .A(n18387), .B(n18388), .Z(n18385) );
  XNOR U22925 ( .A(y[1435]), .B(x[1435]), .Z(n18388) );
  XNOR U22926 ( .A(y[1436]), .B(x[1436]), .Z(n18387) );
  XOR U22927 ( .A(n18361), .B(n18362), .Z(n18380) );
  XNOR U22928 ( .A(n18377), .B(n18378), .Z(n18362) );
  XNOR U22929 ( .A(n18372), .B(n18373), .Z(n18378) );
  XNOR U22930 ( .A(n18374), .B(n18375), .Z(n18373) );
  XNOR U22931 ( .A(y[1432]), .B(x[1432]), .Z(n18375) );
  XNOR U22932 ( .A(y[1433]), .B(x[1433]), .Z(n18374) );
  XNOR U22933 ( .A(y[1431]), .B(x[1431]), .Z(n18372) );
  XNOR U22934 ( .A(n18366), .B(n18367), .Z(n18377) );
  XNOR U22935 ( .A(y[1428]), .B(x[1428]), .Z(n18367) );
  XNOR U22936 ( .A(n18368), .B(n18369), .Z(n18366) );
  XNOR U22937 ( .A(y[1429]), .B(x[1429]), .Z(n18369) );
  XNOR U22938 ( .A(y[1430]), .B(x[1430]), .Z(n18368) );
  XOR U22939 ( .A(n18360), .B(n18359), .Z(n18361) );
  XNOR U22940 ( .A(n18355), .B(n18356), .Z(n18359) );
  XNOR U22941 ( .A(y[1425]), .B(x[1425]), .Z(n18356) );
  XNOR U22942 ( .A(n18357), .B(n18358), .Z(n18355) );
  XNOR U22943 ( .A(y[1426]), .B(x[1426]), .Z(n18358) );
  XNOR U22944 ( .A(y[1427]), .B(x[1427]), .Z(n18357) );
  XNOR U22945 ( .A(n18349), .B(n18350), .Z(n18360) );
  XNOR U22946 ( .A(y[1422]), .B(x[1422]), .Z(n18350) );
  XNOR U22947 ( .A(n18351), .B(n18352), .Z(n18349) );
  XNOR U22948 ( .A(y[1423]), .B(x[1423]), .Z(n18352) );
  XNOR U22949 ( .A(y[1424]), .B(x[1424]), .Z(n18351) );
  NAND U22950 ( .A(n18416), .B(n18417), .Z(N28641) );
  NANDN U22951 ( .A(n18418), .B(n18419), .Z(n18417) );
  OR U22952 ( .A(n18420), .B(n18421), .Z(n18419) );
  NAND U22953 ( .A(n18420), .B(n18421), .Z(n18416) );
  XOR U22954 ( .A(n18420), .B(n18422), .Z(N28640) );
  XNOR U22955 ( .A(n18418), .B(n18421), .Z(n18422) );
  AND U22956 ( .A(n18423), .B(n18424), .Z(n18421) );
  NANDN U22957 ( .A(n18425), .B(n18426), .Z(n18424) );
  NANDN U22958 ( .A(n18427), .B(n18428), .Z(n18426) );
  NANDN U22959 ( .A(n18428), .B(n18427), .Z(n18423) );
  NAND U22960 ( .A(n18429), .B(n18430), .Z(n18418) );
  NANDN U22961 ( .A(n18431), .B(n18432), .Z(n18430) );
  OR U22962 ( .A(n18433), .B(n18434), .Z(n18432) );
  NAND U22963 ( .A(n18434), .B(n18433), .Z(n18429) );
  AND U22964 ( .A(n18435), .B(n18436), .Z(n18420) );
  NANDN U22965 ( .A(n18437), .B(n18438), .Z(n18436) );
  NANDN U22966 ( .A(n18439), .B(n18440), .Z(n18438) );
  NANDN U22967 ( .A(n18440), .B(n18439), .Z(n18435) );
  XOR U22968 ( .A(n18434), .B(n18441), .Z(N28639) );
  XOR U22969 ( .A(n18431), .B(n18433), .Z(n18441) );
  XNOR U22970 ( .A(n18427), .B(n18442), .Z(n18433) );
  XNOR U22971 ( .A(n18425), .B(n18428), .Z(n18442) );
  NAND U22972 ( .A(n18443), .B(n18444), .Z(n18428) );
  NAND U22973 ( .A(n18445), .B(n18446), .Z(n18444) );
  OR U22974 ( .A(n18447), .B(n18448), .Z(n18445) );
  NANDN U22975 ( .A(n18449), .B(n18447), .Z(n18443) );
  IV U22976 ( .A(n18448), .Z(n18449) );
  NAND U22977 ( .A(n18450), .B(n18451), .Z(n18425) );
  NAND U22978 ( .A(n18452), .B(n18453), .Z(n18451) );
  NANDN U22979 ( .A(n18454), .B(n18455), .Z(n18452) );
  NANDN U22980 ( .A(n18455), .B(n18454), .Z(n18450) );
  AND U22981 ( .A(n18456), .B(n18457), .Z(n18427) );
  NAND U22982 ( .A(n18458), .B(n18459), .Z(n18457) );
  OR U22983 ( .A(n18460), .B(n18461), .Z(n18458) );
  NANDN U22984 ( .A(n18462), .B(n18460), .Z(n18456) );
  NAND U22985 ( .A(n18463), .B(n18464), .Z(n18431) );
  NANDN U22986 ( .A(n18465), .B(n18466), .Z(n18464) );
  OR U22987 ( .A(n18467), .B(n18468), .Z(n18466) );
  NANDN U22988 ( .A(n18469), .B(n18467), .Z(n18463) );
  IV U22989 ( .A(n18468), .Z(n18469) );
  XNOR U22990 ( .A(n18439), .B(n18470), .Z(n18434) );
  XNOR U22991 ( .A(n18437), .B(n18440), .Z(n18470) );
  NAND U22992 ( .A(n18471), .B(n18472), .Z(n18440) );
  NAND U22993 ( .A(n18473), .B(n18474), .Z(n18472) );
  OR U22994 ( .A(n18475), .B(n18476), .Z(n18473) );
  NANDN U22995 ( .A(n18477), .B(n18475), .Z(n18471) );
  IV U22996 ( .A(n18476), .Z(n18477) );
  NAND U22997 ( .A(n18478), .B(n18479), .Z(n18437) );
  NAND U22998 ( .A(n18480), .B(n18481), .Z(n18479) );
  NANDN U22999 ( .A(n18482), .B(n18483), .Z(n18480) );
  NANDN U23000 ( .A(n18483), .B(n18482), .Z(n18478) );
  AND U23001 ( .A(n18484), .B(n18485), .Z(n18439) );
  NAND U23002 ( .A(n18486), .B(n18487), .Z(n18485) );
  OR U23003 ( .A(n18488), .B(n18489), .Z(n18486) );
  NANDN U23004 ( .A(n18490), .B(n18488), .Z(n18484) );
  XNOR U23005 ( .A(n18465), .B(n18491), .Z(N28638) );
  XOR U23006 ( .A(n18467), .B(n18468), .Z(n18491) );
  XNOR U23007 ( .A(n18481), .B(n18492), .Z(n18468) );
  XOR U23008 ( .A(n18482), .B(n18483), .Z(n18492) );
  XOR U23009 ( .A(n18488), .B(n18493), .Z(n18483) );
  XOR U23010 ( .A(n18487), .B(n18490), .Z(n18493) );
  IV U23011 ( .A(n18489), .Z(n18490) );
  NAND U23012 ( .A(n18494), .B(n18495), .Z(n18489) );
  OR U23013 ( .A(n18496), .B(n18497), .Z(n18495) );
  OR U23014 ( .A(n18498), .B(n18499), .Z(n18494) );
  NAND U23015 ( .A(n18500), .B(n18501), .Z(n18487) );
  OR U23016 ( .A(n18502), .B(n18503), .Z(n18501) );
  OR U23017 ( .A(n18504), .B(n18505), .Z(n18500) );
  NOR U23018 ( .A(n18506), .B(n18507), .Z(n18488) );
  ANDN U23019 ( .B(n18508), .A(n18509), .Z(n18482) );
  XNOR U23020 ( .A(n18475), .B(n18510), .Z(n18481) );
  XNOR U23021 ( .A(n18474), .B(n18476), .Z(n18510) );
  NAND U23022 ( .A(n18511), .B(n18512), .Z(n18476) );
  OR U23023 ( .A(n18513), .B(n18514), .Z(n18512) );
  OR U23024 ( .A(n18515), .B(n18516), .Z(n18511) );
  NAND U23025 ( .A(n18517), .B(n18518), .Z(n18474) );
  OR U23026 ( .A(n18519), .B(n18520), .Z(n18518) );
  OR U23027 ( .A(n18521), .B(n18522), .Z(n18517) );
  ANDN U23028 ( .B(n18523), .A(n18524), .Z(n18475) );
  IV U23029 ( .A(n18525), .Z(n18523) );
  ANDN U23030 ( .B(n18526), .A(n18527), .Z(n18467) );
  XOR U23031 ( .A(n18453), .B(n18528), .Z(n18465) );
  XOR U23032 ( .A(n18454), .B(n18455), .Z(n18528) );
  XOR U23033 ( .A(n18460), .B(n18529), .Z(n18455) );
  XOR U23034 ( .A(n18459), .B(n18462), .Z(n18529) );
  IV U23035 ( .A(n18461), .Z(n18462) );
  NAND U23036 ( .A(n18530), .B(n18531), .Z(n18461) );
  OR U23037 ( .A(n18532), .B(n18533), .Z(n18531) );
  OR U23038 ( .A(n18534), .B(n18535), .Z(n18530) );
  NAND U23039 ( .A(n18536), .B(n18537), .Z(n18459) );
  OR U23040 ( .A(n18538), .B(n18539), .Z(n18537) );
  OR U23041 ( .A(n18540), .B(n18541), .Z(n18536) );
  NOR U23042 ( .A(n18542), .B(n18543), .Z(n18460) );
  ANDN U23043 ( .B(n18544), .A(n18545), .Z(n18454) );
  IV U23044 ( .A(n18546), .Z(n18544) );
  XNOR U23045 ( .A(n18447), .B(n18547), .Z(n18453) );
  XNOR U23046 ( .A(n18446), .B(n18448), .Z(n18547) );
  NAND U23047 ( .A(n18548), .B(n18549), .Z(n18448) );
  OR U23048 ( .A(n18550), .B(n18551), .Z(n18549) );
  OR U23049 ( .A(n18552), .B(n18553), .Z(n18548) );
  NAND U23050 ( .A(n18554), .B(n18555), .Z(n18446) );
  OR U23051 ( .A(n18556), .B(n18557), .Z(n18555) );
  OR U23052 ( .A(n18558), .B(n18559), .Z(n18554) );
  ANDN U23053 ( .B(n18560), .A(n18561), .Z(n18447) );
  IV U23054 ( .A(n18562), .Z(n18560) );
  XNOR U23055 ( .A(n18527), .B(n18526), .Z(N28637) );
  XOR U23056 ( .A(n18546), .B(n18545), .Z(n18526) );
  XNOR U23057 ( .A(n18561), .B(n18562), .Z(n18545) );
  XNOR U23058 ( .A(n18556), .B(n18557), .Z(n18562) );
  XNOR U23059 ( .A(n18558), .B(n18559), .Z(n18557) );
  XNOR U23060 ( .A(y[1420]), .B(x[1420]), .Z(n18559) );
  XNOR U23061 ( .A(y[1421]), .B(x[1421]), .Z(n18558) );
  XNOR U23062 ( .A(y[1419]), .B(x[1419]), .Z(n18556) );
  XNOR U23063 ( .A(n18550), .B(n18551), .Z(n18561) );
  XNOR U23064 ( .A(y[1416]), .B(x[1416]), .Z(n18551) );
  XNOR U23065 ( .A(n18552), .B(n18553), .Z(n18550) );
  XNOR U23066 ( .A(y[1417]), .B(x[1417]), .Z(n18553) );
  XNOR U23067 ( .A(y[1418]), .B(x[1418]), .Z(n18552) );
  XNOR U23068 ( .A(n18543), .B(n18542), .Z(n18546) );
  XNOR U23069 ( .A(n18538), .B(n18539), .Z(n18542) );
  XNOR U23070 ( .A(y[1413]), .B(x[1413]), .Z(n18539) );
  XNOR U23071 ( .A(n18540), .B(n18541), .Z(n18538) );
  XNOR U23072 ( .A(y[1414]), .B(x[1414]), .Z(n18541) );
  XNOR U23073 ( .A(y[1415]), .B(x[1415]), .Z(n18540) );
  XNOR U23074 ( .A(n18532), .B(n18533), .Z(n18543) );
  XNOR U23075 ( .A(y[1410]), .B(x[1410]), .Z(n18533) );
  XNOR U23076 ( .A(n18534), .B(n18535), .Z(n18532) );
  XNOR U23077 ( .A(y[1411]), .B(x[1411]), .Z(n18535) );
  XNOR U23078 ( .A(y[1412]), .B(x[1412]), .Z(n18534) );
  XOR U23079 ( .A(n18508), .B(n18509), .Z(n18527) );
  XNOR U23080 ( .A(n18524), .B(n18525), .Z(n18509) );
  XNOR U23081 ( .A(n18519), .B(n18520), .Z(n18525) );
  XNOR U23082 ( .A(n18521), .B(n18522), .Z(n18520) );
  XNOR U23083 ( .A(y[1408]), .B(x[1408]), .Z(n18522) );
  XNOR U23084 ( .A(y[1409]), .B(x[1409]), .Z(n18521) );
  XNOR U23085 ( .A(y[1407]), .B(x[1407]), .Z(n18519) );
  XNOR U23086 ( .A(n18513), .B(n18514), .Z(n18524) );
  XNOR U23087 ( .A(y[1404]), .B(x[1404]), .Z(n18514) );
  XNOR U23088 ( .A(n18515), .B(n18516), .Z(n18513) );
  XNOR U23089 ( .A(y[1405]), .B(x[1405]), .Z(n18516) );
  XNOR U23090 ( .A(y[1406]), .B(x[1406]), .Z(n18515) );
  XOR U23091 ( .A(n18507), .B(n18506), .Z(n18508) );
  XNOR U23092 ( .A(n18502), .B(n18503), .Z(n18506) );
  XNOR U23093 ( .A(y[1401]), .B(x[1401]), .Z(n18503) );
  XNOR U23094 ( .A(n18504), .B(n18505), .Z(n18502) );
  XNOR U23095 ( .A(y[1402]), .B(x[1402]), .Z(n18505) );
  XNOR U23096 ( .A(y[1403]), .B(x[1403]), .Z(n18504) );
  XNOR U23097 ( .A(n18496), .B(n18497), .Z(n18507) );
  XNOR U23098 ( .A(y[1398]), .B(x[1398]), .Z(n18497) );
  XNOR U23099 ( .A(n18498), .B(n18499), .Z(n18496) );
  XNOR U23100 ( .A(y[1399]), .B(x[1399]), .Z(n18499) );
  XNOR U23101 ( .A(y[1400]), .B(x[1400]), .Z(n18498) );
  NAND U23102 ( .A(n18563), .B(n18564), .Z(N28629) );
  NANDN U23103 ( .A(n18565), .B(n18566), .Z(n18564) );
  OR U23104 ( .A(n18567), .B(n18568), .Z(n18566) );
  NAND U23105 ( .A(n18567), .B(n18568), .Z(n18563) );
  XOR U23106 ( .A(n18567), .B(n18569), .Z(N28628) );
  XNOR U23107 ( .A(n18565), .B(n18568), .Z(n18569) );
  AND U23108 ( .A(n18570), .B(n18571), .Z(n18568) );
  NANDN U23109 ( .A(n18572), .B(n18573), .Z(n18571) );
  NANDN U23110 ( .A(n18574), .B(n18575), .Z(n18573) );
  NANDN U23111 ( .A(n18575), .B(n18574), .Z(n18570) );
  NAND U23112 ( .A(n18576), .B(n18577), .Z(n18565) );
  NANDN U23113 ( .A(n18578), .B(n18579), .Z(n18577) );
  OR U23114 ( .A(n18580), .B(n18581), .Z(n18579) );
  NAND U23115 ( .A(n18581), .B(n18580), .Z(n18576) );
  AND U23116 ( .A(n18582), .B(n18583), .Z(n18567) );
  NANDN U23117 ( .A(n18584), .B(n18585), .Z(n18583) );
  NANDN U23118 ( .A(n18586), .B(n18587), .Z(n18585) );
  NANDN U23119 ( .A(n18587), .B(n18586), .Z(n18582) );
  XOR U23120 ( .A(n18581), .B(n18588), .Z(N28627) );
  XOR U23121 ( .A(n18578), .B(n18580), .Z(n18588) );
  XNOR U23122 ( .A(n18574), .B(n18589), .Z(n18580) );
  XNOR U23123 ( .A(n18572), .B(n18575), .Z(n18589) );
  NAND U23124 ( .A(n18590), .B(n18591), .Z(n18575) );
  NAND U23125 ( .A(n18592), .B(n18593), .Z(n18591) );
  OR U23126 ( .A(n18594), .B(n18595), .Z(n18592) );
  NANDN U23127 ( .A(n18596), .B(n18594), .Z(n18590) );
  IV U23128 ( .A(n18595), .Z(n18596) );
  NAND U23129 ( .A(n18597), .B(n18598), .Z(n18572) );
  NAND U23130 ( .A(n18599), .B(n18600), .Z(n18598) );
  NANDN U23131 ( .A(n18601), .B(n18602), .Z(n18599) );
  NANDN U23132 ( .A(n18602), .B(n18601), .Z(n18597) );
  AND U23133 ( .A(n18603), .B(n18604), .Z(n18574) );
  NAND U23134 ( .A(n18605), .B(n18606), .Z(n18604) );
  OR U23135 ( .A(n18607), .B(n18608), .Z(n18605) );
  NANDN U23136 ( .A(n18609), .B(n18607), .Z(n18603) );
  NAND U23137 ( .A(n18610), .B(n18611), .Z(n18578) );
  NANDN U23138 ( .A(n18612), .B(n18613), .Z(n18611) );
  OR U23139 ( .A(n18614), .B(n18615), .Z(n18613) );
  NANDN U23140 ( .A(n18616), .B(n18614), .Z(n18610) );
  IV U23141 ( .A(n18615), .Z(n18616) );
  XNOR U23142 ( .A(n18586), .B(n18617), .Z(n18581) );
  XNOR U23143 ( .A(n18584), .B(n18587), .Z(n18617) );
  NAND U23144 ( .A(n18618), .B(n18619), .Z(n18587) );
  NAND U23145 ( .A(n18620), .B(n18621), .Z(n18619) );
  OR U23146 ( .A(n18622), .B(n18623), .Z(n18620) );
  NANDN U23147 ( .A(n18624), .B(n18622), .Z(n18618) );
  IV U23148 ( .A(n18623), .Z(n18624) );
  NAND U23149 ( .A(n18625), .B(n18626), .Z(n18584) );
  NAND U23150 ( .A(n18627), .B(n18628), .Z(n18626) );
  NANDN U23151 ( .A(n18629), .B(n18630), .Z(n18627) );
  NANDN U23152 ( .A(n18630), .B(n18629), .Z(n18625) );
  AND U23153 ( .A(n18631), .B(n18632), .Z(n18586) );
  NAND U23154 ( .A(n18633), .B(n18634), .Z(n18632) );
  OR U23155 ( .A(n18635), .B(n18636), .Z(n18633) );
  NANDN U23156 ( .A(n18637), .B(n18635), .Z(n18631) );
  XNOR U23157 ( .A(n18612), .B(n18638), .Z(N28626) );
  XOR U23158 ( .A(n18614), .B(n18615), .Z(n18638) );
  XNOR U23159 ( .A(n18628), .B(n18639), .Z(n18615) );
  XOR U23160 ( .A(n18629), .B(n18630), .Z(n18639) );
  XOR U23161 ( .A(n18635), .B(n18640), .Z(n18630) );
  XOR U23162 ( .A(n18634), .B(n18637), .Z(n18640) );
  IV U23163 ( .A(n18636), .Z(n18637) );
  NAND U23164 ( .A(n18641), .B(n18642), .Z(n18636) );
  OR U23165 ( .A(n18643), .B(n18644), .Z(n18642) );
  OR U23166 ( .A(n18645), .B(n18646), .Z(n18641) );
  NAND U23167 ( .A(n18647), .B(n18648), .Z(n18634) );
  OR U23168 ( .A(n18649), .B(n18650), .Z(n18648) );
  OR U23169 ( .A(n18651), .B(n18652), .Z(n18647) );
  NOR U23170 ( .A(n18653), .B(n18654), .Z(n18635) );
  ANDN U23171 ( .B(n18655), .A(n18656), .Z(n18629) );
  XNOR U23172 ( .A(n18622), .B(n18657), .Z(n18628) );
  XNOR U23173 ( .A(n18621), .B(n18623), .Z(n18657) );
  NAND U23174 ( .A(n18658), .B(n18659), .Z(n18623) );
  OR U23175 ( .A(n18660), .B(n18661), .Z(n18659) );
  OR U23176 ( .A(n18662), .B(n18663), .Z(n18658) );
  NAND U23177 ( .A(n18664), .B(n18665), .Z(n18621) );
  OR U23178 ( .A(n18666), .B(n18667), .Z(n18665) );
  OR U23179 ( .A(n18668), .B(n18669), .Z(n18664) );
  ANDN U23180 ( .B(n18670), .A(n18671), .Z(n18622) );
  IV U23181 ( .A(n18672), .Z(n18670) );
  ANDN U23182 ( .B(n18673), .A(n18674), .Z(n18614) );
  XOR U23183 ( .A(n18600), .B(n18675), .Z(n18612) );
  XOR U23184 ( .A(n18601), .B(n18602), .Z(n18675) );
  XOR U23185 ( .A(n18607), .B(n18676), .Z(n18602) );
  XOR U23186 ( .A(n18606), .B(n18609), .Z(n18676) );
  IV U23187 ( .A(n18608), .Z(n18609) );
  NAND U23188 ( .A(n18677), .B(n18678), .Z(n18608) );
  OR U23189 ( .A(n18679), .B(n18680), .Z(n18678) );
  OR U23190 ( .A(n18681), .B(n18682), .Z(n18677) );
  NAND U23191 ( .A(n18683), .B(n18684), .Z(n18606) );
  OR U23192 ( .A(n18685), .B(n18686), .Z(n18684) );
  OR U23193 ( .A(n18687), .B(n18688), .Z(n18683) );
  NOR U23194 ( .A(n18689), .B(n18690), .Z(n18607) );
  ANDN U23195 ( .B(n18691), .A(n18692), .Z(n18601) );
  IV U23196 ( .A(n18693), .Z(n18691) );
  XNOR U23197 ( .A(n18594), .B(n18694), .Z(n18600) );
  XNOR U23198 ( .A(n18593), .B(n18595), .Z(n18694) );
  NAND U23199 ( .A(n18695), .B(n18696), .Z(n18595) );
  OR U23200 ( .A(n18697), .B(n18698), .Z(n18696) );
  OR U23201 ( .A(n18699), .B(n18700), .Z(n18695) );
  NAND U23202 ( .A(n18701), .B(n18702), .Z(n18593) );
  OR U23203 ( .A(n18703), .B(n18704), .Z(n18702) );
  OR U23204 ( .A(n18705), .B(n18706), .Z(n18701) );
  ANDN U23205 ( .B(n18707), .A(n18708), .Z(n18594) );
  IV U23206 ( .A(n18709), .Z(n18707) );
  XNOR U23207 ( .A(n18674), .B(n18673), .Z(N28625) );
  XOR U23208 ( .A(n18693), .B(n18692), .Z(n18673) );
  XNOR U23209 ( .A(n18708), .B(n18709), .Z(n18692) );
  XNOR U23210 ( .A(n18703), .B(n18704), .Z(n18709) );
  XNOR U23211 ( .A(n18705), .B(n18706), .Z(n18704) );
  XNOR U23212 ( .A(y[1396]), .B(x[1396]), .Z(n18706) );
  XNOR U23213 ( .A(y[1397]), .B(x[1397]), .Z(n18705) );
  XNOR U23214 ( .A(y[1395]), .B(x[1395]), .Z(n18703) );
  XNOR U23215 ( .A(n18697), .B(n18698), .Z(n18708) );
  XNOR U23216 ( .A(y[1392]), .B(x[1392]), .Z(n18698) );
  XNOR U23217 ( .A(n18699), .B(n18700), .Z(n18697) );
  XNOR U23218 ( .A(y[1393]), .B(x[1393]), .Z(n18700) );
  XNOR U23219 ( .A(y[1394]), .B(x[1394]), .Z(n18699) );
  XNOR U23220 ( .A(n18690), .B(n18689), .Z(n18693) );
  XNOR U23221 ( .A(n18685), .B(n18686), .Z(n18689) );
  XNOR U23222 ( .A(y[1389]), .B(x[1389]), .Z(n18686) );
  XNOR U23223 ( .A(n18687), .B(n18688), .Z(n18685) );
  XNOR U23224 ( .A(y[1390]), .B(x[1390]), .Z(n18688) );
  XNOR U23225 ( .A(y[1391]), .B(x[1391]), .Z(n18687) );
  XNOR U23226 ( .A(n18679), .B(n18680), .Z(n18690) );
  XNOR U23227 ( .A(y[1386]), .B(x[1386]), .Z(n18680) );
  XNOR U23228 ( .A(n18681), .B(n18682), .Z(n18679) );
  XNOR U23229 ( .A(y[1387]), .B(x[1387]), .Z(n18682) );
  XNOR U23230 ( .A(y[1388]), .B(x[1388]), .Z(n18681) );
  XOR U23231 ( .A(n18655), .B(n18656), .Z(n18674) );
  XNOR U23232 ( .A(n18671), .B(n18672), .Z(n18656) );
  XNOR U23233 ( .A(n18666), .B(n18667), .Z(n18672) );
  XNOR U23234 ( .A(n18668), .B(n18669), .Z(n18667) );
  XNOR U23235 ( .A(y[1384]), .B(x[1384]), .Z(n18669) );
  XNOR U23236 ( .A(y[1385]), .B(x[1385]), .Z(n18668) );
  XNOR U23237 ( .A(y[1383]), .B(x[1383]), .Z(n18666) );
  XNOR U23238 ( .A(n18660), .B(n18661), .Z(n18671) );
  XNOR U23239 ( .A(y[1380]), .B(x[1380]), .Z(n18661) );
  XNOR U23240 ( .A(n18662), .B(n18663), .Z(n18660) );
  XNOR U23241 ( .A(y[1381]), .B(x[1381]), .Z(n18663) );
  XNOR U23242 ( .A(y[1382]), .B(x[1382]), .Z(n18662) );
  XOR U23243 ( .A(n18654), .B(n18653), .Z(n18655) );
  XNOR U23244 ( .A(n18649), .B(n18650), .Z(n18653) );
  XNOR U23245 ( .A(y[1377]), .B(x[1377]), .Z(n18650) );
  XNOR U23246 ( .A(n18651), .B(n18652), .Z(n18649) );
  XNOR U23247 ( .A(y[1378]), .B(x[1378]), .Z(n18652) );
  XNOR U23248 ( .A(y[1379]), .B(x[1379]), .Z(n18651) );
  XNOR U23249 ( .A(n18643), .B(n18644), .Z(n18654) );
  XNOR U23250 ( .A(y[1374]), .B(x[1374]), .Z(n18644) );
  XNOR U23251 ( .A(n18645), .B(n18646), .Z(n18643) );
  XNOR U23252 ( .A(y[1375]), .B(x[1375]), .Z(n18646) );
  XNOR U23253 ( .A(y[1376]), .B(x[1376]), .Z(n18645) );
  NAND U23254 ( .A(n18710), .B(n18711), .Z(N28617) );
  NANDN U23255 ( .A(n18712), .B(n18713), .Z(n18711) );
  OR U23256 ( .A(n18714), .B(n18715), .Z(n18713) );
  NAND U23257 ( .A(n18714), .B(n18715), .Z(n18710) );
  XOR U23258 ( .A(n18714), .B(n18716), .Z(N28616) );
  XNOR U23259 ( .A(n18712), .B(n18715), .Z(n18716) );
  AND U23260 ( .A(n18717), .B(n18718), .Z(n18715) );
  NANDN U23261 ( .A(n18719), .B(n18720), .Z(n18718) );
  NANDN U23262 ( .A(n18721), .B(n18722), .Z(n18720) );
  NANDN U23263 ( .A(n18722), .B(n18721), .Z(n18717) );
  NAND U23264 ( .A(n18723), .B(n18724), .Z(n18712) );
  NANDN U23265 ( .A(n18725), .B(n18726), .Z(n18724) );
  OR U23266 ( .A(n18727), .B(n18728), .Z(n18726) );
  NAND U23267 ( .A(n18728), .B(n18727), .Z(n18723) );
  AND U23268 ( .A(n18729), .B(n18730), .Z(n18714) );
  NANDN U23269 ( .A(n18731), .B(n18732), .Z(n18730) );
  NANDN U23270 ( .A(n18733), .B(n18734), .Z(n18732) );
  NANDN U23271 ( .A(n18734), .B(n18733), .Z(n18729) );
  XOR U23272 ( .A(n18728), .B(n18735), .Z(N28615) );
  XOR U23273 ( .A(n18725), .B(n18727), .Z(n18735) );
  XNOR U23274 ( .A(n18721), .B(n18736), .Z(n18727) );
  XNOR U23275 ( .A(n18719), .B(n18722), .Z(n18736) );
  NAND U23276 ( .A(n18737), .B(n18738), .Z(n18722) );
  NAND U23277 ( .A(n18739), .B(n18740), .Z(n18738) );
  OR U23278 ( .A(n18741), .B(n18742), .Z(n18739) );
  NANDN U23279 ( .A(n18743), .B(n18741), .Z(n18737) );
  IV U23280 ( .A(n18742), .Z(n18743) );
  NAND U23281 ( .A(n18744), .B(n18745), .Z(n18719) );
  NAND U23282 ( .A(n18746), .B(n18747), .Z(n18745) );
  NANDN U23283 ( .A(n18748), .B(n18749), .Z(n18746) );
  NANDN U23284 ( .A(n18749), .B(n18748), .Z(n18744) );
  AND U23285 ( .A(n18750), .B(n18751), .Z(n18721) );
  NAND U23286 ( .A(n18752), .B(n18753), .Z(n18751) );
  OR U23287 ( .A(n18754), .B(n18755), .Z(n18752) );
  NANDN U23288 ( .A(n18756), .B(n18754), .Z(n18750) );
  NAND U23289 ( .A(n18757), .B(n18758), .Z(n18725) );
  NANDN U23290 ( .A(n18759), .B(n18760), .Z(n18758) );
  OR U23291 ( .A(n18761), .B(n18762), .Z(n18760) );
  NANDN U23292 ( .A(n18763), .B(n18761), .Z(n18757) );
  IV U23293 ( .A(n18762), .Z(n18763) );
  XNOR U23294 ( .A(n18733), .B(n18764), .Z(n18728) );
  XNOR U23295 ( .A(n18731), .B(n18734), .Z(n18764) );
  NAND U23296 ( .A(n18765), .B(n18766), .Z(n18734) );
  NAND U23297 ( .A(n18767), .B(n18768), .Z(n18766) );
  OR U23298 ( .A(n18769), .B(n18770), .Z(n18767) );
  NANDN U23299 ( .A(n18771), .B(n18769), .Z(n18765) );
  IV U23300 ( .A(n18770), .Z(n18771) );
  NAND U23301 ( .A(n18772), .B(n18773), .Z(n18731) );
  NAND U23302 ( .A(n18774), .B(n18775), .Z(n18773) );
  NANDN U23303 ( .A(n18776), .B(n18777), .Z(n18774) );
  NANDN U23304 ( .A(n18777), .B(n18776), .Z(n18772) );
  AND U23305 ( .A(n18778), .B(n18779), .Z(n18733) );
  NAND U23306 ( .A(n18780), .B(n18781), .Z(n18779) );
  OR U23307 ( .A(n18782), .B(n18783), .Z(n18780) );
  NANDN U23308 ( .A(n18784), .B(n18782), .Z(n18778) );
  XNOR U23309 ( .A(n18759), .B(n18785), .Z(N28614) );
  XOR U23310 ( .A(n18761), .B(n18762), .Z(n18785) );
  XNOR U23311 ( .A(n18775), .B(n18786), .Z(n18762) );
  XOR U23312 ( .A(n18776), .B(n18777), .Z(n18786) );
  XOR U23313 ( .A(n18782), .B(n18787), .Z(n18777) );
  XOR U23314 ( .A(n18781), .B(n18784), .Z(n18787) );
  IV U23315 ( .A(n18783), .Z(n18784) );
  NAND U23316 ( .A(n18788), .B(n18789), .Z(n18783) );
  OR U23317 ( .A(n18790), .B(n18791), .Z(n18789) );
  OR U23318 ( .A(n18792), .B(n18793), .Z(n18788) );
  NAND U23319 ( .A(n18794), .B(n18795), .Z(n18781) );
  OR U23320 ( .A(n18796), .B(n18797), .Z(n18795) );
  OR U23321 ( .A(n18798), .B(n18799), .Z(n18794) );
  NOR U23322 ( .A(n18800), .B(n18801), .Z(n18782) );
  ANDN U23323 ( .B(n18802), .A(n18803), .Z(n18776) );
  XNOR U23324 ( .A(n18769), .B(n18804), .Z(n18775) );
  XNOR U23325 ( .A(n18768), .B(n18770), .Z(n18804) );
  NAND U23326 ( .A(n18805), .B(n18806), .Z(n18770) );
  OR U23327 ( .A(n18807), .B(n18808), .Z(n18806) );
  OR U23328 ( .A(n18809), .B(n18810), .Z(n18805) );
  NAND U23329 ( .A(n18811), .B(n18812), .Z(n18768) );
  OR U23330 ( .A(n18813), .B(n18814), .Z(n18812) );
  OR U23331 ( .A(n18815), .B(n18816), .Z(n18811) );
  ANDN U23332 ( .B(n18817), .A(n18818), .Z(n18769) );
  IV U23333 ( .A(n18819), .Z(n18817) );
  ANDN U23334 ( .B(n18820), .A(n18821), .Z(n18761) );
  XOR U23335 ( .A(n18747), .B(n18822), .Z(n18759) );
  XOR U23336 ( .A(n18748), .B(n18749), .Z(n18822) );
  XOR U23337 ( .A(n18754), .B(n18823), .Z(n18749) );
  XOR U23338 ( .A(n18753), .B(n18756), .Z(n18823) );
  IV U23339 ( .A(n18755), .Z(n18756) );
  NAND U23340 ( .A(n18824), .B(n18825), .Z(n18755) );
  OR U23341 ( .A(n18826), .B(n18827), .Z(n18825) );
  OR U23342 ( .A(n18828), .B(n18829), .Z(n18824) );
  NAND U23343 ( .A(n18830), .B(n18831), .Z(n18753) );
  OR U23344 ( .A(n18832), .B(n18833), .Z(n18831) );
  OR U23345 ( .A(n18834), .B(n18835), .Z(n18830) );
  NOR U23346 ( .A(n18836), .B(n18837), .Z(n18754) );
  ANDN U23347 ( .B(n18838), .A(n18839), .Z(n18748) );
  IV U23348 ( .A(n18840), .Z(n18838) );
  XNOR U23349 ( .A(n18741), .B(n18841), .Z(n18747) );
  XNOR U23350 ( .A(n18740), .B(n18742), .Z(n18841) );
  NAND U23351 ( .A(n18842), .B(n18843), .Z(n18742) );
  OR U23352 ( .A(n18844), .B(n18845), .Z(n18843) );
  OR U23353 ( .A(n18846), .B(n18847), .Z(n18842) );
  NAND U23354 ( .A(n18848), .B(n18849), .Z(n18740) );
  OR U23355 ( .A(n18850), .B(n18851), .Z(n18849) );
  OR U23356 ( .A(n18852), .B(n18853), .Z(n18848) );
  ANDN U23357 ( .B(n18854), .A(n18855), .Z(n18741) );
  IV U23358 ( .A(n18856), .Z(n18854) );
  XNOR U23359 ( .A(n18821), .B(n18820), .Z(N28613) );
  XOR U23360 ( .A(n18840), .B(n18839), .Z(n18820) );
  XNOR U23361 ( .A(n18855), .B(n18856), .Z(n18839) );
  XNOR U23362 ( .A(n18850), .B(n18851), .Z(n18856) );
  XNOR U23363 ( .A(n18852), .B(n18853), .Z(n18851) );
  XNOR U23364 ( .A(y[1372]), .B(x[1372]), .Z(n18853) );
  XNOR U23365 ( .A(y[1373]), .B(x[1373]), .Z(n18852) );
  XNOR U23366 ( .A(y[1371]), .B(x[1371]), .Z(n18850) );
  XNOR U23367 ( .A(n18844), .B(n18845), .Z(n18855) );
  XNOR U23368 ( .A(y[1368]), .B(x[1368]), .Z(n18845) );
  XNOR U23369 ( .A(n18846), .B(n18847), .Z(n18844) );
  XNOR U23370 ( .A(y[1369]), .B(x[1369]), .Z(n18847) );
  XNOR U23371 ( .A(y[1370]), .B(x[1370]), .Z(n18846) );
  XNOR U23372 ( .A(n18837), .B(n18836), .Z(n18840) );
  XNOR U23373 ( .A(n18832), .B(n18833), .Z(n18836) );
  XNOR U23374 ( .A(y[1365]), .B(x[1365]), .Z(n18833) );
  XNOR U23375 ( .A(n18834), .B(n18835), .Z(n18832) );
  XNOR U23376 ( .A(y[1366]), .B(x[1366]), .Z(n18835) );
  XNOR U23377 ( .A(y[1367]), .B(x[1367]), .Z(n18834) );
  XNOR U23378 ( .A(n18826), .B(n18827), .Z(n18837) );
  XNOR U23379 ( .A(y[1362]), .B(x[1362]), .Z(n18827) );
  XNOR U23380 ( .A(n18828), .B(n18829), .Z(n18826) );
  XNOR U23381 ( .A(y[1363]), .B(x[1363]), .Z(n18829) );
  XNOR U23382 ( .A(y[1364]), .B(x[1364]), .Z(n18828) );
  XOR U23383 ( .A(n18802), .B(n18803), .Z(n18821) );
  XNOR U23384 ( .A(n18818), .B(n18819), .Z(n18803) );
  XNOR U23385 ( .A(n18813), .B(n18814), .Z(n18819) );
  XNOR U23386 ( .A(n18815), .B(n18816), .Z(n18814) );
  XNOR U23387 ( .A(y[1360]), .B(x[1360]), .Z(n18816) );
  XNOR U23388 ( .A(y[1361]), .B(x[1361]), .Z(n18815) );
  XNOR U23389 ( .A(y[1359]), .B(x[1359]), .Z(n18813) );
  XNOR U23390 ( .A(n18807), .B(n18808), .Z(n18818) );
  XNOR U23391 ( .A(y[1356]), .B(x[1356]), .Z(n18808) );
  XNOR U23392 ( .A(n18809), .B(n18810), .Z(n18807) );
  XNOR U23393 ( .A(y[1357]), .B(x[1357]), .Z(n18810) );
  XNOR U23394 ( .A(y[1358]), .B(x[1358]), .Z(n18809) );
  XOR U23395 ( .A(n18801), .B(n18800), .Z(n18802) );
  XNOR U23396 ( .A(n18796), .B(n18797), .Z(n18800) );
  XNOR U23397 ( .A(y[1353]), .B(x[1353]), .Z(n18797) );
  XNOR U23398 ( .A(n18798), .B(n18799), .Z(n18796) );
  XNOR U23399 ( .A(y[1354]), .B(x[1354]), .Z(n18799) );
  XNOR U23400 ( .A(y[1355]), .B(x[1355]), .Z(n18798) );
  XNOR U23401 ( .A(n18790), .B(n18791), .Z(n18801) );
  XNOR U23402 ( .A(y[1350]), .B(x[1350]), .Z(n18791) );
  XNOR U23403 ( .A(n18792), .B(n18793), .Z(n18790) );
  XNOR U23404 ( .A(y[1351]), .B(x[1351]), .Z(n18793) );
  XNOR U23405 ( .A(y[1352]), .B(x[1352]), .Z(n18792) );
  NAND U23406 ( .A(n18857), .B(n18858), .Z(N28605) );
  NANDN U23407 ( .A(n18859), .B(n18860), .Z(n18858) );
  OR U23408 ( .A(n18861), .B(n18862), .Z(n18860) );
  NAND U23409 ( .A(n18861), .B(n18862), .Z(n18857) );
  XOR U23410 ( .A(n18861), .B(n18863), .Z(N28604) );
  XNOR U23411 ( .A(n18859), .B(n18862), .Z(n18863) );
  AND U23412 ( .A(n18864), .B(n18865), .Z(n18862) );
  NANDN U23413 ( .A(n18866), .B(n18867), .Z(n18865) );
  NANDN U23414 ( .A(n18868), .B(n18869), .Z(n18867) );
  NANDN U23415 ( .A(n18869), .B(n18868), .Z(n18864) );
  NAND U23416 ( .A(n18870), .B(n18871), .Z(n18859) );
  NANDN U23417 ( .A(n18872), .B(n18873), .Z(n18871) );
  OR U23418 ( .A(n18874), .B(n18875), .Z(n18873) );
  NAND U23419 ( .A(n18875), .B(n18874), .Z(n18870) );
  AND U23420 ( .A(n18876), .B(n18877), .Z(n18861) );
  NANDN U23421 ( .A(n18878), .B(n18879), .Z(n18877) );
  NANDN U23422 ( .A(n18880), .B(n18881), .Z(n18879) );
  NANDN U23423 ( .A(n18881), .B(n18880), .Z(n18876) );
  XOR U23424 ( .A(n18875), .B(n18882), .Z(N28603) );
  XOR U23425 ( .A(n18872), .B(n18874), .Z(n18882) );
  XNOR U23426 ( .A(n18868), .B(n18883), .Z(n18874) );
  XNOR U23427 ( .A(n18866), .B(n18869), .Z(n18883) );
  NAND U23428 ( .A(n18884), .B(n18885), .Z(n18869) );
  NAND U23429 ( .A(n18886), .B(n18887), .Z(n18885) );
  OR U23430 ( .A(n18888), .B(n18889), .Z(n18886) );
  NANDN U23431 ( .A(n18890), .B(n18888), .Z(n18884) );
  IV U23432 ( .A(n18889), .Z(n18890) );
  NAND U23433 ( .A(n18891), .B(n18892), .Z(n18866) );
  NAND U23434 ( .A(n18893), .B(n18894), .Z(n18892) );
  NANDN U23435 ( .A(n18895), .B(n18896), .Z(n18893) );
  NANDN U23436 ( .A(n18896), .B(n18895), .Z(n18891) );
  AND U23437 ( .A(n18897), .B(n18898), .Z(n18868) );
  NAND U23438 ( .A(n18899), .B(n18900), .Z(n18898) );
  OR U23439 ( .A(n18901), .B(n18902), .Z(n18899) );
  NANDN U23440 ( .A(n18903), .B(n18901), .Z(n18897) );
  NAND U23441 ( .A(n18904), .B(n18905), .Z(n18872) );
  NANDN U23442 ( .A(n18906), .B(n18907), .Z(n18905) );
  OR U23443 ( .A(n18908), .B(n18909), .Z(n18907) );
  NANDN U23444 ( .A(n18910), .B(n18908), .Z(n18904) );
  IV U23445 ( .A(n18909), .Z(n18910) );
  XNOR U23446 ( .A(n18880), .B(n18911), .Z(n18875) );
  XNOR U23447 ( .A(n18878), .B(n18881), .Z(n18911) );
  NAND U23448 ( .A(n18912), .B(n18913), .Z(n18881) );
  NAND U23449 ( .A(n18914), .B(n18915), .Z(n18913) );
  OR U23450 ( .A(n18916), .B(n18917), .Z(n18914) );
  NANDN U23451 ( .A(n18918), .B(n18916), .Z(n18912) );
  IV U23452 ( .A(n18917), .Z(n18918) );
  NAND U23453 ( .A(n18919), .B(n18920), .Z(n18878) );
  NAND U23454 ( .A(n18921), .B(n18922), .Z(n18920) );
  NANDN U23455 ( .A(n18923), .B(n18924), .Z(n18921) );
  NANDN U23456 ( .A(n18924), .B(n18923), .Z(n18919) );
  AND U23457 ( .A(n18925), .B(n18926), .Z(n18880) );
  NAND U23458 ( .A(n18927), .B(n18928), .Z(n18926) );
  OR U23459 ( .A(n18929), .B(n18930), .Z(n18927) );
  NANDN U23460 ( .A(n18931), .B(n18929), .Z(n18925) );
  XNOR U23461 ( .A(n18906), .B(n18932), .Z(N28602) );
  XOR U23462 ( .A(n18908), .B(n18909), .Z(n18932) );
  XNOR U23463 ( .A(n18922), .B(n18933), .Z(n18909) );
  XOR U23464 ( .A(n18923), .B(n18924), .Z(n18933) );
  XOR U23465 ( .A(n18929), .B(n18934), .Z(n18924) );
  XOR U23466 ( .A(n18928), .B(n18931), .Z(n18934) );
  IV U23467 ( .A(n18930), .Z(n18931) );
  NAND U23468 ( .A(n18935), .B(n18936), .Z(n18930) );
  OR U23469 ( .A(n18937), .B(n18938), .Z(n18936) );
  OR U23470 ( .A(n18939), .B(n18940), .Z(n18935) );
  NAND U23471 ( .A(n18941), .B(n18942), .Z(n18928) );
  OR U23472 ( .A(n18943), .B(n18944), .Z(n18942) );
  OR U23473 ( .A(n18945), .B(n18946), .Z(n18941) );
  NOR U23474 ( .A(n18947), .B(n18948), .Z(n18929) );
  ANDN U23475 ( .B(n18949), .A(n18950), .Z(n18923) );
  XNOR U23476 ( .A(n18916), .B(n18951), .Z(n18922) );
  XNOR U23477 ( .A(n18915), .B(n18917), .Z(n18951) );
  NAND U23478 ( .A(n18952), .B(n18953), .Z(n18917) );
  OR U23479 ( .A(n18954), .B(n18955), .Z(n18953) );
  OR U23480 ( .A(n18956), .B(n18957), .Z(n18952) );
  NAND U23481 ( .A(n18958), .B(n18959), .Z(n18915) );
  OR U23482 ( .A(n18960), .B(n18961), .Z(n18959) );
  OR U23483 ( .A(n18962), .B(n18963), .Z(n18958) );
  ANDN U23484 ( .B(n18964), .A(n18965), .Z(n18916) );
  IV U23485 ( .A(n18966), .Z(n18964) );
  ANDN U23486 ( .B(n18967), .A(n18968), .Z(n18908) );
  XOR U23487 ( .A(n18894), .B(n18969), .Z(n18906) );
  XOR U23488 ( .A(n18895), .B(n18896), .Z(n18969) );
  XOR U23489 ( .A(n18901), .B(n18970), .Z(n18896) );
  XOR U23490 ( .A(n18900), .B(n18903), .Z(n18970) );
  IV U23491 ( .A(n18902), .Z(n18903) );
  NAND U23492 ( .A(n18971), .B(n18972), .Z(n18902) );
  OR U23493 ( .A(n18973), .B(n18974), .Z(n18972) );
  OR U23494 ( .A(n18975), .B(n18976), .Z(n18971) );
  NAND U23495 ( .A(n18977), .B(n18978), .Z(n18900) );
  OR U23496 ( .A(n18979), .B(n18980), .Z(n18978) );
  OR U23497 ( .A(n18981), .B(n18982), .Z(n18977) );
  NOR U23498 ( .A(n18983), .B(n18984), .Z(n18901) );
  ANDN U23499 ( .B(n18985), .A(n18986), .Z(n18895) );
  IV U23500 ( .A(n18987), .Z(n18985) );
  XNOR U23501 ( .A(n18888), .B(n18988), .Z(n18894) );
  XNOR U23502 ( .A(n18887), .B(n18889), .Z(n18988) );
  NAND U23503 ( .A(n18989), .B(n18990), .Z(n18889) );
  OR U23504 ( .A(n18991), .B(n18992), .Z(n18990) );
  OR U23505 ( .A(n18993), .B(n18994), .Z(n18989) );
  NAND U23506 ( .A(n18995), .B(n18996), .Z(n18887) );
  OR U23507 ( .A(n18997), .B(n18998), .Z(n18996) );
  OR U23508 ( .A(n18999), .B(n19000), .Z(n18995) );
  ANDN U23509 ( .B(n19001), .A(n19002), .Z(n18888) );
  IV U23510 ( .A(n19003), .Z(n19001) );
  XNOR U23511 ( .A(n18968), .B(n18967), .Z(N28601) );
  XOR U23512 ( .A(n18987), .B(n18986), .Z(n18967) );
  XNOR U23513 ( .A(n19002), .B(n19003), .Z(n18986) );
  XNOR U23514 ( .A(n18997), .B(n18998), .Z(n19003) );
  XNOR U23515 ( .A(n18999), .B(n19000), .Z(n18998) );
  XNOR U23516 ( .A(y[1348]), .B(x[1348]), .Z(n19000) );
  XNOR U23517 ( .A(y[1349]), .B(x[1349]), .Z(n18999) );
  XNOR U23518 ( .A(y[1347]), .B(x[1347]), .Z(n18997) );
  XNOR U23519 ( .A(n18991), .B(n18992), .Z(n19002) );
  XNOR U23520 ( .A(y[1344]), .B(x[1344]), .Z(n18992) );
  XNOR U23521 ( .A(n18993), .B(n18994), .Z(n18991) );
  XNOR U23522 ( .A(y[1345]), .B(x[1345]), .Z(n18994) );
  XNOR U23523 ( .A(y[1346]), .B(x[1346]), .Z(n18993) );
  XNOR U23524 ( .A(n18984), .B(n18983), .Z(n18987) );
  XNOR U23525 ( .A(n18979), .B(n18980), .Z(n18983) );
  XNOR U23526 ( .A(y[1341]), .B(x[1341]), .Z(n18980) );
  XNOR U23527 ( .A(n18981), .B(n18982), .Z(n18979) );
  XNOR U23528 ( .A(y[1342]), .B(x[1342]), .Z(n18982) );
  XNOR U23529 ( .A(y[1343]), .B(x[1343]), .Z(n18981) );
  XNOR U23530 ( .A(n18973), .B(n18974), .Z(n18984) );
  XNOR U23531 ( .A(y[1338]), .B(x[1338]), .Z(n18974) );
  XNOR U23532 ( .A(n18975), .B(n18976), .Z(n18973) );
  XNOR U23533 ( .A(y[1339]), .B(x[1339]), .Z(n18976) );
  XNOR U23534 ( .A(y[1340]), .B(x[1340]), .Z(n18975) );
  XOR U23535 ( .A(n18949), .B(n18950), .Z(n18968) );
  XNOR U23536 ( .A(n18965), .B(n18966), .Z(n18950) );
  XNOR U23537 ( .A(n18960), .B(n18961), .Z(n18966) );
  XNOR U23538 ( .A(n18962), .B(n18963), .Z(n18961) );
  XNOR U23539 ( .A(y[1336]), .B(x[1336]), .Z(n18963) );
  XNOR U23540 ( .A(y[1337]), .B(x[1337]), .Z(n18962) );
  XNOR U23541 ( .A(y[1335]), .B(x[1335]), .Z(n18960) );
  XNOR U23542 ( .A(n18954), .B(n18955), .Z(n18965) );
  XNOR U23543 ( .A(y[1332]), .B(x[1332]), .Z(n18955) );
  XNOR U23544 ( .A(n18956), .B(n18957), .Z(n18954) );
  XNOR U23545 ( .A(y[1333]), .B(x[1333]), .Z(n18957) );
  XNOR U23546 ( .A(y[1334]), .B(x[1334]), .Z(n18956) );
  XOR U23547 ( .A(n18948), .B(n18947), .Z(n18949) );
  XNOR U23548 ( .A(n18943), .B(n18944), .Z(n18947) );
  XNOR U23549 ( .A(y[1329]), .B(x[1329]), .Z(n18944) );
  XNOR U23550 ( .A(n18945), .B(n18946), .Z(n18943) );
  XNOR U23551 ( .A(y[1330]), .B(x[1330]), .Z(n18946) );
  XNOR U23552 ( .A(y[1331]), .B(x[1331]), .Z(n18945) );
  XNOR U23553 ( .A(n18937), .B(n18938), .Z(n18948) );
  XNOR U23554 ( .A(y[1326]), .B(x[1326]), .Z(n18938) );
  XNOR U23555 ( .A(n18939), .B(n18940), .Z(n18937) );
  XNOR U23556 ( .A(y[1327]), .B(x[1327]), .Z(n18940) );
  XNOR U23557 ( .A(y[1328]), .B(x[1328]), .Z(n18939) );
  NAND U23558 ( .A(n19004), .B(n19005), .Z(N28593) );
  NANDN U23559 ( .A(n19006), .B(n19007), .Z(n19005) );
  OR U23560 ( .A(n19008), .B(n19009), .Z(n19007) );
  NAND U23561 ( .A(n19008), .B(n19009), .Z(n19004) );
  XOR U23562 ( .A(n19008), .B(n19010), .Z(N28592) );
  XNOR U23563 ( .A(n19006), .B(n19009), .Z(n19010) );
  AND U23564 ( .A(n19011), .B(n19012), .Z(n19009) );
  NANDN U23565 ( .A(n19013), .B(n19014), .Z(n19012) );
  NANDN U23566 ( .A(n19015), .B(n19016), .Z(n19014) );
  NANDN U23567 ( .A(n19016), .B(n19015), .Z(n19011) );
  NAND U23568 ( .A(n19017), .B(n19018), .Z(n19006) );
  NANDN U23569 ( .A(n19019), .B(n19020), .Z(n19018) );
  OR U23570 ( .A(n19021), .B(n19022), .Z(n19020) );
  NAND U23571 ( .A(n19022), .B(n19021), .Z(n19017) );
  AND U23572 ( .A(n19023), .B(n19024), .Z(n19008) );
  NANDN U23573 ( .A(n19025), .B(n19026), .Z(n19024) );
  NANDN U23574 ( .A(n19027), .B(n19028), .Z(n19026) );
  NANDN U23575 ( .A(n19028), .B(n19027), .Z(n19023) );
  XOR U23576 ( .A(n19022), .B(n19029), .Z(N28591) );
  XOR U23577 ( .A(n19019), .B(n19021), .Z(n19029) );
  XNOR U23578 ( .A(n19015), .B(n19030), .Z(n19021) );
  XNOR U23579 ( .A(n19013), .B(n19016), .Z(n19030) );
  NAND U23580 ( .A(n19031), .B(n19032), .Z(n19016) );
  NAND U23581 ( .A(n19033), .B(n19034), .Z(n19032) );
  OR U23582 ( .A(n19035), .B(n19036), .Z(n19033) );
  NANDN U23583 ( .A(n19037), .B(n19035), .Z(n19031) );
  IV U23584 ( .A(n19036), .Z(n19037) );
  NAND U23585 ( .A(n19038), .B(n19039), .Z(n19013) );
  NAND U23586 ( .A(n19040), .B(n19041), .Z(n19039) );
  NANDN U23587 ( .A(n19042), .B(n19043), .Z(n19040) );
  NANDN U23588 ( .A(n19043), .B(n19042), .Z(n19038) );
  AND U23589 ( .A(n19044), .B(n19045), .Z(n19015) );
  NAND U23590 ( .A(n19046), .B(n19047), .Z(n19045) );
  OR U23591 ( .A(n19048), .B(n19049), .Z(n19046) );
  NANDN U23592 ( .A(n19050), .B(n19048), .Z(n19044) );
  NAND U23593 ( .A(n19051), .B(n19052), .Z(n19019) );
  NANDN U23594 ( .A(n19053), .B(n19054), .Z(n19052) );
  OR U23595 ( .A(n19055), .B(n19056), .Z(n19054) );
  NANDN U23596 ( .A(n19057), .B(n19055), .Z(n19051) );
  IV U23597 ( .A(n19056), .Z(n19057) );
  XNOR U23598 ( .A(n19027), .B(n19058), .Z(n19022) );
  XNOR U23599 ( .A(n19025), .B(n19028), .Z(n19058) );
  NAND U23600 ( .A(n19059), .B(n19060), .Z(n19028) );
  NAND U23601 ( .A(n19061), .B(n19062), .Z(n19060) );
  OR U23602 ( .A(n19063), .B(n19064), .Z(n19061) );
  NANDN U23603 ( .A(n19065), .B(n19063), .Z(n19059) );
  IV U23604 ( .A(n19064), .Z(n19065) );
  NAND U23605 ( .A(n19066), .B(n19067), .Z(n19025) );
  NAND U23606 ( .A(n19068), .B(n19069), .Z(n19067) );
  NANDN U23607 ( .A(n19070), .B(n19071), .Z(n19068) );
  NANDN U23608 ( .A(n19071), .B(n19070), .Z(n19066) );
  AND U23609 ( .A(n19072), .B(n19073), .Z(n19027) );
  NAND U23610 ( .A(n19074), .B(n19075), .Z(n19073) );
  OR U23611 ( .A(n19076), .B(n19077), .Z(n19074) );
  NANDN U23612 ( .A(n19078), .B(n19076), .Z(n19072) );
  XNOR U23613 ( .A(n19053), .B(n19079), .Z(N28590) );
  XOR U23614 ( .A(n19055), .B(n19056), .Z(n19079) );
  XNOR U23615 ( .A(n19069), .B(n19080), .Z(n19056) );
  XOR U23616 ( .A(n19070), .B(n19071), .Z(n19080) );
  XOR U23617 ( .A(n19076), .B(n19081), .Z(n19071) );
  XOR U23618 ( .A(n19075), .B(n19078), .Z(n19081) );
  IV U23619 ( .A(n19077), .Z(n19078) );
  NAND U23620 ( .A(n19082), .B(n19083), .Z(n19077) );
  OR U23621 ( .A(n19084), .B(n19085), .Z(n19083) );
  OR U23622 ( .A(n19086), .B(n19087), .Z(n19082) );
  NAND U23623 ( .A(n19088), .B(n19089), .Z(n19075) );
  OR U23624 ( .A(n19090), .B(n19091), .Z(n19089) );
  OR U23625 ( .A(n19092), .B(n19093), .Z(n19088) );
  NOR U23626 ( .A(n19094), .B(n19095), .Z(n19076) );
  ANDN U23627 ( .B(n19096), .A(n19097), .Z(n19070) );
  XNOR U23628 ( .A(n19063), .B(n19098), .Z(n19069) );
  XNOR U23629 ( .A(n19062), .B(n19064), .Z(n19098) );
  NAND U23630 ( .A(n19099), .B(n19100), .Z(n19064) );
  OR U23631 ( .A(n19101), .B(n19102), .Z(n19100) );
  OR U23632 ( .A(n19103), .B(n19104), .Z(n19099) );
  NAND U23633 ( .A(n19105), .B(n19106), .Z(n19062) );
  OR U23634 ( .A(n19107), .B(n19108), .Z(n19106) );
  OR U23635 ( .A(n19109), .B(n19110), .Z(n19105) );
  ANDN U23636 ( .B(n19111), .A(n19112), .Z(n19063) );
  IV U23637 ( .A(n19113), .Z(n19111) );
  ANDN U23638 ( .B(n19114), .A(n19115), .Z(n19055) );
  XOR U23639 ( .A(n19041), .B(n19116), .Z(n19053) );
  XOR U23640 ( .A(n19042), .B(n19043), .Z(n19116) );
  XOR U23641 ( .A(n19048), .B(n19117), .Z(n19043) );
  XOR U23642 ( .A(n19047), .B(n19050), .Z(n19117) );
  IV U23643 ( .A(n19049), .Z(n19050) );
  NAND U23644 ( .A(n19118), .B(n19119), .Z(n19049) );
  OR U23645 ( .A(n19120), .B(n19121), .Z(n19119) );
  OR U23646 ( .A(n19122), .B(n19123), .Z(n19118) );
  NAND U23647 ( .A(n19124), .B(n19125), .Z(n19047) );
  OR U23648 ( .A(n19126), .B(n19127), .Z(n19125) );
  OR U23649 ( .A(n19128), .B(n19129), .Z(n19124) );
  NOR U23650 ( .A(n19130), .B(n19131), .Z(n19048) );
  ANDN U23651 ( .B(n19132), .A(n19133), .Z(n19042) );
  IV U23652 ( .A(n19134), .Z(n19132) );
  XNOR U23653 ( .A(n19035), .B(n19135), .Z(n19041) );
  XNOR U23654 ( .A(n19034), .B(n19036), .Z(n19135) );
  NAND U23655 ( .A(n19136), .B(n19137), .Z(n19036) );
  OR U23656 ( .A(n19138), .B(n19139), .Z(n19137) );
  OR U23657 ( .A(n19140), .B(n19141), .Z(n19136) );
  NAND U23658 ( .A(n19142), .B(n19143), .Z(n19034) );
  OR U23659 ( .A(n19144), .B(n19145), .Z(n19143) );
  OR U23660 ( .A(n19146), .B(n19147), .Z(n19142) );
  ANDN U23661 ( .B(n19148), .A(n19149), .Z(n19035) );
  IV U23662 ( .A(n19150), .Z(n19148) );
  XNOR U23663 ( .A(n19115), .B(n19114), .Z(N28589) );
  XOR U23664 ( .A(n19134), .B(n19133), .Z(n19114) );
  XNOR U23665 ( .A(n19149), .B(n19150), .Z(n19133) );
  XNOR U23666 ( .A(n19144), .B(n19145), .Z(n19150) );
  XNOR U23667 ( .A(n19146), .B(n19147), .Z(n19145) );
  XNOR U23668 ( .A(y[1324]), .B(x[1324]), .Z(n19147) );
  XNOR U23669 ( .A(y[1325]), .B(x[1325]), .Z(n19146) );
  XNOR U23670 ( .A(y[1323]), .B(x[1323]), .Z(n19144) );
  XNOR U23671 ( .A(n19138), .B(n19139), .Z(n19149) );
  XNOR U23672 ( .A(y[1320]), .B(x[1320]), .Z(n19139) );
  XNOR U23673 ( .A(n19140), .B(n19141), .Z(n19138) );
  XNOR U23674 ( .A(y[1321]), .B(x[1321]), .Z(n19141) );
  XNOR U23675 ( .A(y[1322]), .B(x[1322]), .Z(n19140) );
  XNOR U23676 ( .A(n19131), .B(n19130), .Z(n19134) );
  XNOR U23677 ( .A(n19126), .B(n19127), .Z(n19130) );
  XNOR U23678 ( .A(y[1317]), .B(x[1317]), .Z(n19127) );
  XNOR U23679 ( .A(n19128), .B(n19129), .Z(n19126) );
  XNOR U23680 ( .A(y[1318]), .B(x[1318]), .Z(n19129) );
  XNOR U23681 ( .A(y[1319]), .B(x[1319]), .Z(n19128) );
  XNOR U23682 ( .A(n19120), .B(n19121), .Z(n19131) );
  XNOR U23683 ( .A(y[1314]), .B(x[1314]), .Z(n19121) );
  XNOR U23684 ( .A(n19122), .B(n19123), .Z(n19120) );
  XNOR U23685 ( .A(y[1315]), .B(x[1315]), .Z(n19123) );
  XNOR U23686 ( .A(y[1316]), .B(x[1316]), .Z(n19122) );
  XOR U23687 ( .A(n19096), .B(n19097), .Z(n19115) );
  XNOR U23688 ( .A(n19112), .B(n19113), .Z(n19097) );
  XNOR U23689 ( .A(n19107), .B(n19108), .Z(n19113) );
  XNOR U23690 ( .A(n19109), .B(n19110), .Z(n19108) );
  XNOR U23691 ( .A(y[1312]), .B(x[1312]), .Z(n19110) );
  XNOR U23692 ( .A(y[1313]), .B(x[1313]), .Z(n19109) );
  XNOR U23693 ( .A(y[1311]), .B(x[1311]), .Z(n19107) );
  XNOR U23694 ( .A(n19101), .B(n19102), .Z(n19112) );
  XNOR U23695 ( .A(y[1308]), .B(x[1308]), .Z(n19102) );
  XNOR U23696 ( .A(n19103), .B(n19104), .Z(n19101) );
  XNOR U23697 ( .A(y[1309]), .B(x[1309]), .Z(n19104) );
  XNOR U23698 ( .A(y[1310]), .B(x[1310]), .Z(n19103) );
  XOR U23699 ( .A(n19095), .B(n19094), .Z(n19096) );
  XNOR U23700 ( .A(n19090), .B(n19091), .Z(n19094) );
  XNOR U23701 ( .A(y[1305]), .B(x[1305]), .Z(n19091) );
  XNOR U23702 ( .A(n19092), .B(n19093), .Z(n19090) );
  XNOR U23703 ( .A(y[1306]), .B(x[1306]), .Z(n19093) );
  XNOR U23704 ( .A(y[1307]), .B(x[1307]), .Z(n19092) );
  XNOR U23705 ( .A(n19084), .B(n19085), .Z(n19095) );
  XNOR U23706 ( .A(y[1302]), .B(x[1302]), .Z(n19085) );
  XNOR U23707 ( .A(n19086), .B(n19087), .Z(n19084) );
  XNOR U23708 ( .A(y[1303]), .B(x[1303]), .Z(n19087) );
  XNOR U23709 ( .A(y[1304]), .B(x[1304]), .Z(n19086) );
  NAND U23710 ( .A(n19151), .B(n19152), .Z(N28581) );
  NANDN U23711 ( .A(n19153), .B(n19154), .Z(n19152) );
  OR U23712 ( .A(n19155), .B(n19156), .Z(n19154) );
  NAND U23713 ( .A(n19155), .B(n19156), .Z(n19151) );
  XOR U23714 ( .A(n19155), .B(n19157), .Z(N28580) );
  XNOR U23715 ( .A(n19153), .B(n19156), .Z(n19157) );
  AND U23716 ( .A(n19158), .B(n19159), .Z(n19156) );
  NANDN U23717 ( .A(n19160), .B(n19161), .Z(n19159) );
  NANDN U23718 ( .A(n19162), .B(n19163), .Z(n19161) );
  NANDN U23719 ( .A(n19163), .B(n19162), .Z(n19158) );
  NAND U23720 ( .A(n19164), .B(n19165), .Z(n19153) );
  NANDN U23721 ( .A(n19166), .B(n19167), .Z(n19165) );
  OR U23722 ( .A(n19168), .B(n19169), .Z(n19167) );
  NAND U23723 ( .A(n19169), .B(n19168), .Z(n19164) );
  AND U23724 ( .A(n19170), .B(n19171), .Z(n19155) );
  NANDN U23725 ( .A(n19172), .B(n19173), .Z(n19171) );
  NANDN U23726 ( .A(n19174), .B(n19175), .Z(n19173) );
  NANDN U23727 ( .A(n19175), .B(n19174), .Z(n19170) );
  XOR U23728 ( .A(n19169), .B(n19176), .Z(N28579) );
  XOR U23729 ( .A(n19166), .B(n19168), .Z(n19176) );
  XNOR U23730 ( .A(n19162), .B(n19177), .Z(n19168) );
  XNOR U23731 ( .A(n19160), .B(n19163), .Z(n19177) );
  NAND U23732 ( .A(n19178), .B(n19179), .Z(n19163) );
  NAND U23733 ( .A(n19180), .B(n19181), .Z(n19179) );
  OR U23734 ( .A(n19182), .B(n19183), .Z(n19180) );
  NANDN U23735 ( .A(n19184), .B(n19182), .Z(n19178) );
  IV U23736 ( .A(n19183), .Z(n19184) );
  NAND U23737 ( .A(n19185), .B(n19186), .Z(n19160) );
  NAND U23738 ( .A(n19187), .B(n19188), .Z(n19186) );
  NANDN U23739 ( .A(n19189), .B(n19190), .Z(n19187) );
  NANDN U23740 ( .A(n19190), .B(n19189), .Z(n19185) );
  AND U23741 ( .A(n19191), .B(n19192), .Z(n19162) );
  NAND U23742 ( .A(n19193), .B(n19194), .Z(n19192) );
  OR U23743 ( .A(n19195), .B(n19196), .Z(n19193) );
  NANDN U23744 ( .A(n19197), .B(n19195), .Z(n19191) );
  NAND U23745 ( .A(n19198), .B(n19199), .Z(n19166) );
  NANDN U23746 ( .A(n19200), .B(n19201), .Z(n19199) );
  OR U23747 ( .A(n19202), .B(n19203), .Z(n19201) );
  NANDN U23748 ( .A(n19204), .B(n19202), .Z(n19198) );
  IV U23749 ( .A(n19203), .Z(n19204) );
  XNOR U23750 ( .A(n19174), .B(n19205), .Z(n19169) );
  XNOR U23751 ( .A(n19172), .B(n19175), .Z(n19205) );
  NAND U23752 ( .A(n19206), .B(n19207), .Z(n19175) );
  NAND U23753 ( .A(n19208), .B(n19209), .Z(n19207) );
  OR U23754 ( .A(n19210), .B(n19211), .Z(n19208) );
  NANDN U23755 ( .A(n19212), .B(n19210), .Z(n19206) );
  IV U23756 ( .A(n19211), .Z(n19212) );
  NAND U23757 ( .A(n19213), .B(n19214), .Z(n19172) );
  NAND U23758 ( .A(n19215), .B(n19216), .Z(n19214) );
  NANDN U23759 ( .A(n19217), .B(n19218), .Z(n19215) );
  NANDN U23760 ( .A(n19218), .B(n19217), .Z(n19213) );
  AND U23761 ( .A(n19219), .B(n19220), .Z(n19174) );
  NAND U23762 ( .A(n19221), .B(n19222), .Z(n19220) );
  OR U23763 ( .A(n19223), .B(n19224), .Z(n19221) );
  NANDN U23764 ( .A(n19225), .B(n19223), .Z(n19219) );
  XNOR U23765 ( .A(n19200), .B(n19226), .Z(N28578) );
  XOR U23766 ( .A(n19202), .B(n19203), .Z(n19226) );
  XNOR U23767 ( .A(n19216), .B(n19227), .Z(n19203) );
  XOR U23768 ( .A(n19217), .B(n19218), .Z(n19227) );
  XOR U23769 ( .A(n19223), .B(n19228), .Z(n19218) );
  XOR U23770 ( .A(n19222), .B(n19225), .Z(n19228) );
  IV U23771 ( .A(n19224), .Z(n19225) );
  NAND U23772 ( .A(n19229), .B(n19230), .Z(n19224) );
  OR U23773 ( .A(n19231), .B(n19232), .Z(n19230) );
  OR U23774 ( .A(n19233), .B(n19234), .Z(n19229) );
  NAND U23775 ( .A(n19235), .B(n19236), .Z(n19222) );
  OR U23776 ( .A(n19237), .B(n19238), .Z(n19236) );
  OR U23777 ( .A(n19239), .B(n19240), .Z(n19235) );
  NOR U23778 ( .A(n19241), .B(n19242), .Z(n19223) );
  ANDN U23779 ( .B(n19243), .A(n19244), .Z(n19217) );
  XNOR U23780 ( .A(n19210), .B(n19245), .Z(n19216) );
  XNOR U23781 ( .A(n19209), .B(n19211), .Z(n19245) );
  NAND U23782 ( .A(n19246), .B(n19247), .Z(n19211) );
  OR U23783 ( .A(n19248), .B(n19249), .Z(n19247) );
  OR U23784 ( .A(n19250), .B(n19251), .Z(n19246) );
  NAND U23785 ( .A(n19252), .B(n19253), .Z(n19209) );
  OR U23786 ( .A(n19254), .B(n19255), .Z(n19253) );
  OR U23787 ( .A(n19256), .B(n19257), .Z(n19252) );
  ANDN U23788 ( .B(n19258), .A(n19259), .Z(n19210) );
  IV U23789 ( .A(n19260), .Z(n19258) );
  ANDN U23790 ( .B(n19261), .A(n19262), .Z(n19202) );
  XOR U23791 ( .A(n19188), .B(n19263), .Z(n19200) );
  XOR U23792 ( .A(n19189), .B(n19190), .Z(n19263) );
  XOR U23793 ( .A(n19195), .B(n19264), .Z(n19190) );
  XOR U23794 ( .A(n19194), .B(n19197), .Z(n19264) );
  IV U23795 ( .A(n19196), .Z(n19197) );
  NAND U23796 ( .A(n19265), .B(n19266), .Z(n19196) );
  OR U23797 ( .A(n19267), .B(n19268), .Z(n19266) );
  OR U23798 ( .A(n19269), .B(n19270), .Z(n19265) );
  NAND U23799 ( .A(n19271), .B(n19272), .Z(n19194) );
  OR U23800 ( .A(n19273), .B(n19274), .Z(n19272) );
  OR U23801 ( .A(n19275), .B(n19276), .Z(n19271) );
  NOR U23802 ( .A(n19277), .B(n19278), .Z(n19195) );
  ANDN U23803 ( .B(n19279), .A(n19280), .Z(n19189) );
  IV U23804 ( .A(n19281), .Z(n19279) );
  XNOR U23805 ( .A(n19182), .B(n19282), .Z(n19188) );
  XNOR U23806 ( .A(n19181), .B(n19183), .Z(n19282) );
  NAND U23807 ( .A(n19283), .B(n19284), .Z(n19183) );
  OR U23808 ( .A(n19285), .B(n19286), .Z(n19284) );
  OR U23809 ( .A(n19287), .B(n19288), .Z(n19283) );
  NAND U23810 ( .A(n19289), .B(n19290), .Z(n19181) );
  OR U23811 ( .A(n19291), .B(n19292), .Z(n19290) );
  OR U23812 ( .A(n19293), .B(n19294), .Z(n19289) );
  ANDN U23813 ( .B(n19295), .A(n19296), .Z(n19182) );
  IV U23814 ( .A(n19297), .Z(n19295) );
  XNOR U23815 ( .A(n19262), .B(n19261), .Z(N28577) );
  XOR U23816 ( .A(n19281), .B(n19280), .Z(n19261) );
  XNOR U23817 ( .A(n19296), .B(n19297), .Z(n19280) );
  XNOR U23818 ( .A(n19291), .B(n19292), .Z(n19297) );
  XNOR U23819 ( .A(n19293), .B(n19294), .Z(n19292) );
  XNOR U23820 ( .A(y[1300]), .B(x[1300]), .Z(n19294) );
  XNOR U23821 ( .A(y[1301]), .B(x[1301]), .Z(n19293) );
  XNOR U23822 ( .A(y[1299]), .B(x[1299]), .Z(n19291) );
  XNOR U23823 ( .A(n19285), .B(n19286), .Z(n19296) );
  XNOR U23824 ( .A(y[1296]), .B(x[1296]), .Z(n19286) );
  XNOR U23825 ( .A(n19287), .B(n19288), .Z(n19285) );
  XNOR U23826 ( .A(y[1297]), .B(x[1297]), .Z(n19288) );
  XNOR U23827 ( .A(y[1298]), .B(x[1298]), .Z(n19287) );
  XNOR U23828 ( .A(n19278), .B(n19277), .Z(n19281) );
  XNOR U23829 ( .A(n19273), .B(n19274), .Z(n19277) );
  XNOR U23830 ( .A(y[1293]), .B(x[1293]), .Z(n19274) );
  XNOR U23831 ( .A(n19275), .B(n19276), .Z(n19273) );
  XNOR U23832 ( .A(y[1294]), .B(x[1294]), .Z(n19276) );
  XNOR U23833 ( .A(y[1295]), .B(x[1295]), .Z(n19275) );
  XNOR U23834 ( .A(n19267), .B(n19268), .Z(n19278) );
  XNOR U23835 ( .A(y[1290]), .B(x[1290]), .Z(n19268) );
  XNOR U23836 ( .A(n19269), .B(n19270), .Z(n19267) );
  XNOR U23837 ( .A(y[1291]), .B(x[1291]), .Z(n19270) );
  XNOR U23838 ( .A(y[1292]), .B(x[1292]), .Z(n19269) );
  XOR U23839 ( .A(n19243), .B(n19244), .Z(n19262) );
  XNOR U23840 ( .A(n19259), .B(n19260), .Z(n19244) );
  XNOR U23841 ( .A(n19254), .B(n19255), .Z(n19260) );
  XNOR U23842 ( .A(n19256), .B(n19257), .Z(n19255) );
  XNOR U23843 ( .A(y[1288]), .B(x[1288]), .Z(n19257) );
  XNOR U23844 ( .A(y[1289]), .B(x[1289]), .Z(n19256) );
  XNOR U23845 ( .A(y[1287]), .B(x[1287]), .Z(n19254) );
  XNOR U23846 ( .A(n19248), .B(n19249), .Z(n19259) );
  XNOR U23847 ( .A(y[1284]), .B(x[1284]), .Z(n19249) );
  XNOR U23848 ( .A(n19250), .B(n19251), .Z(n19248) );
  XNOR U23849 ( .A(y[1285]), .B(x[1285]), .Z(n19251) );
  XNOR U23850 ( .A(y[1286]), .B(x[1286]), .Z(n19250) );
  XOR U23851 ( .A(n19242), .B(n19241), .Z(n19243) );
  XNOR U23852 ( .A(n19237), .B(n19238), .Z(n19241) );
  XNOR U23853 ( .A(y[1281]), .B(x[1281]), .Z(n19238) );
  XNOR U23854 ( .A(n19239), .B(n19240), .Z(n19237) );
  XNOR U23855 ( .A(y[1282]), .B(x[1282]), .Z(n19240) );
  XNOR U23856 ( .A(y[1283]), .B(x[1283]), .Z(n19239) );
  XNOR U23857 ( .A(n19231), .B(n19232), .Z(n19242) );
  XNOR U23858 ( .A(y[1278]), .B(x[1278]), .Z(n19232) );
  XNOR U23859 ( .A(n19233), .B(n19234), .Z(n19231) );
  XNOR U23860 ( .A(y[1279]), .B(x[1279]), .Z(n19234) );
  XNOR U23861 ( .A(y[1280]), .B(x[1280]), .Z(n19233) );
  NAND U23862 ( .A(n19298), .B(n19299), .Z(N28569) );
  NANDN U23863 ( .A(n19300), .B(n19301), .Z(n19299) );
  OR U23864 ( .A(n19302), .B(n19303), .Z(n19301) );
  NAND U23865 ( .A(n19302), .B(n19303), .Z(n19298) );
  XOR U23866 ( .A(n19302), .B(n19304), .Z(N28568) );
  XNOR U23867 ( .A(n19300), .B(n19303), .Z(n19304) );
  AND U23868 ( .A(n19305), .B(n19306), .Z(n19303) );
  NANDN U23869 ( .A(n19307), .B(n19308), .Z(n19306) );
  NANDN U23870 ( .A(n19309), .B(n19310), .Z(n19308) );
  NANDN U23871 ( .A(n19310), .B(n19309), .Z(n19305) );
  NAND U23872 ( .A(n19311), .B(n19312), .Z(n19300) );
  NANDN U23873 ( .A(n19313), .B(n19314), .Z(n19312) );
  OR U23874 ( .A(n19315), .B(n19316), .Z(n19314) );
  NAND U23875 ( .A(n19316), .B(n19315), .Z(n19311) );
  AND U23876 ( .A(n19317), .B(n19318), .Z(n19302) );
  NANDN U23877 ( .A(n19319), .B(n19320), .Z(n19318) );
  NANDN U23878 ( .A(n19321), .B(n19322), .Z(n19320) );
  NANDN U23879 ( .A(n19322), .B(n19321), .Z(n19317) );
  XOR U23880 ( .A(n19316), .B(n19323), .Z(N28567) );
  XOR U23881 ( .A(n19313), .B(n19315), .Z(n19323) );
  XNOR U23882 ( .A(n19309), .B(n19324), .Z(n19315) );
  XNOR U23883 ( .A(n19307), .B(n19310), .Z(n19324) );
  NAND U23884 ( .A(n19325), .B(n19326), .Z(n19310) );
  NAND U23885 ( .A(n19327), .B(n19328), .Z(n19326) );
  OR U23886 ( .A(n19329), .B(n19330), .Z(n19327) );
  NANDN U23887 ( .A(n19331), .B(n19329), .Z(n19325) );
  IV U23888 ( .A(n19330), .Z(n19331) );
  NAND U23889 ( .A(n19332), .B(n19333), .Z(n19307) );
  NAND U23890 ( .A(n19334), .B(n19335), .Z(n19333) );
  NANDN U23891 ( .A(n19336), .B(n19337), .Z(n19334) );
  NANDN U23892 ( .A(n19337), .B(n19336), .Z(n19332) );
  AND U23893 ( .A(n19338), .B(n19339), .Z(n19309) );
  NAND U23894 ( .A(n19340), .B(n19341), .Z(n19339) );
  OR U23895 ( .A(n19342), .B(n19343), .Z(n19340) );
  NANDN U23896 ( .A(n19344), .B(n19342), .Z(n19338) );
  NAND U23897 ( .A(n19345), .B(n19346), .Z(n19313) );
  NANDN U23898 ( .A(n19347), .B(n19348), .Z(n19346) );
  OR U23899 ( .A(n19349), .B(n19350), .Z(n19348) );
  NANDN U23900 ( .A(n19351), .B(n19349), .Z(n19345) );
  IV U23901 ( .A(n19350), .Z(n19351) );
  XNOR U23902 ( .A(n19321), .B(n19352), .Z(n19316) );
  XNOR U23903 ( .A(n19319), .B(n19322), .Z(n19352) );
  NAND U23904 ( .A(n19353), .B(n19354), .Z(n19322) );
  NAND U23905 ( .A(n19355), .B(n19356), .Z(n19354) );
  OR U23906 ( .A(n19357), .B(n19358), .Z(n19355) );
  NANDN U23907 ( .A(n19359), .B(n19357), .Z(n19353) );
  IV U23908 ( .A(n19358), .Z(n19359) );
  NAND U23909 ( .A(n19360), .B(n19361), .Z(n19319) );
  NAND U23910 ( .A(n19362), .B(n19363), .Z(n19361) );
  NANDN U23911 ( .A(n19364), .B(n19365), .Z(n19362) );
  NANDN U23912 ( .A(n19365), .B(n19364), .Z(n19360) );
  AND U23913 ( .A(n19366), .B(n19367), .Z(n19321) );
  NAND U23914 ( .A(n19368), .B(n19369), .Z(n19367) );
  OR U23915 ( .A(n19370), .B(n19371), .Z(n19368) );
  NANDN U23916 ( .A(n19372), .B(n19370), .Z(n19366) );
  XNOR U23917 ( .A(n19347), .B(n19373), .Z(N28566) );
  XOR U23918 ( .A(n19349), .B(n19350), .Z(n19373) );
  XNOR U23919 ( .A(n19363), .B(n19374), .Z(n19350) );
  XOR U23920 ( .A(n19364), .B(n19365), .Z(n19374) );
  XOR U23921 ( .A(n19370), .B(n19375), .Z(n19365) );
  XOR U23922 ( .A(n19369), .B(n19372), .Z(n19375) );
  IV U23923 ( .A(n19371), .Z(n19372) );
  NAND U23924 ( .A(n19376), .B(n19377), .Z(n19371) );
  OR U23925 ( .A(n19378), .B(n19379), .Z(n19377) );
  OR U23926 ( .A(n19380), .B(n19381), .Z(n19376) );
  NAND U23927 ( .A(n19382), .B(n19383), .Z(n19369) );
  OR U23928 ( .A(n19384), .B(n19385), .Z(n19383) );
  OR U23929 ( .A(n19386), .B(n19387), .Z(n19382) );
  NOR U23930 ( .A(n19388), .B(n19389), .Z(n19370) );
  ANDN U23931 ( .B(n19390), .A(n19391), .Z(n19364) );
  XNOR U23932 ( .A(n19357), .B(n19392), .Z(n19363) );
  XNOR U23933 ( .A(n19356), .B(n19358), .Z(n19392) );
  NAND U23934 ( .A(n19393), .B(n19394), .Z(n19358) );
  OR U23935 ( .A(n19395), .B(n19396), .Z(n19394) );
  OR U23936 ( .A(n19397), .B(n19398), .Z(n19393) );
  NAND U23937 ( .A(n19399), .B(n19400), .Z(n19356) );
  OR U23938 ( .A(n19401), .B(n19402), .Z(n19400) );
  OR U23939 ( .A(n19403), .B(n19404), .Z(n19399) );
  ANDN U23940 ( .B(n19405), .A(n19406), .Z(n19357) );
  IV U23941 ( .A(n19407), .Z(n19405) );
  ANDN U23942 ( .B(n19408), .A(n19409), .Z(n19349) );
  XOR U23943 ( .A(n19335), .B(n19410), .Z(n19347) );
  XOR U23944 ( .A(n19336), .B(n19337), .Z(n19410) );
  XOR U23945 ( .A(n19342), .B(n19411), .Z(n19337) );
  XOR U23946 ( .A(n19341), .B(n19344), .Z(n19411) );
  IV U23947 ( .A(n19343), .Z(n19344) );
  NAND U23948 ( .A(n19412), .B(n19413), .Z(n19343) );
  OR U23949 ( .A(n19414), .B(n19415), .Z(n19413) );
  OR U23950 ( .A(n19416), .B(n19417), .Z(n19412) );
  NAND U23951 ( .A(n19418), .B(n19419), .Z(n19341) );
  OR U23952 ( .A(n19420), .B(n19421), .Z(n19419) );
  OR U23953 ( .A(n19422), .B(n19423), .Z(n19418) );
  NOR U23954 ( .A(n19424), .B(n19425), .Z(n19342) );
  ANDN U23955 ( .B(n19426), .A(n19427), .Z(n19336) );
  IV U23956 ( .A(n19428), .Z(n19426) );
  XNOR U23957 ( .A(n19329), .B(n19429), .Z(n19335) );
  XNOR U23958 ( .A(n19328), .B(n19330), .Z(n19429) );
  NAND U23959 ( .A(n19430), .B(n19431), .Z(n19330) );
  OR U23960 ( .A(n19432), .B(n19433), .Z(n19431) );
  OR U23961 ( .A(n19434), .B(n19435), .Z(n19430) );
  NAND U23962 ( .A(n19436), .B(n19437), .Z(n19328) );
  OR U23963 ( .A(n19438), .B(n19439), .Z(n19437) );
  OR U23964 ( .A(n19440), .B(n19441), .Z(n19436) );
  ANDN U23965 ( .B(n19442), .A(n19443), .Z(n19329) );
  IV U23966 ( .A(n19444), .Z(n19442) );
  XNOR U23967 ( .A(n19409), .B(n19408), .Z(N28565) );
  XOR U23968 ( .A(n19428), .B(n19427), .Z(n19408) );
  XNOR U23969 ( .A(n19443), .B(n19444), .Z(n19427) );
  XNOR U23970 ( .A(n19438), .B(n19439), .Z(n19444) );
  XNOR U23971 ( .A(n19440), .B(n19441), .Z(n19439) );
  XNOR U23972 ( .A(y[1276]), .B(x[1276]), .Z(n19441) );
  XNOR U23973 ( .A(y[1277]), .B(x[1277]), .Z(n19440) );
  XNOR U23974 ( .A(y[1275]), .B(x[1275]), .Z(n19438) );
  XNOR U23975 ( .A(n19432), .B(n19433), .Z(n19443) );
  XNOR U23976 ( .A(y[1272]), .B(x[1272]), .Z(n19433) );
  XNOR U23977 ( .A(n19434), .B(n19435), .Z(n19432) );
  XNOR U23978 ( .A(y[1273]), .B(x[1273]), .Z(n19435) );
  XNOR U23979 ( .A(y[1274]), .B(x[1274]), .Z(n19434) );
  XNOR U23980 ( .A(n19425), .B(n19424), .Z(n19428) );
  XNOR U23981 ( .A(n19420), .B(n19421), .Z(n19424) );
  XNOR U23982 ( .A(y[1269]), .B(x[1269]), .Z(n19421) );
  XNOR U23983 ( .A(n19422), .B(n19423), .Z(n19420) );
  XNOR U23984 ( .A(y[1270]), .B(x[1270]), .Z(n19423) );
  XNOR U23985 ( .A(y[1271]), .B(x[1271]), .Z(n19422) );
  XNOR U23986 ( .A(n19414), .B(n19415), .Z(n19425) );
  XNOR U23987 ( .A(y[1266]), .B(x[1266]), .Z(n19415) );
  XNOR U23988 ( .A(n19416), .B(n19417), .Z(n19414) );
  XNOR U23989 ( .A(y[1267]), .B(x[1267]), .Z(n19417) );
  XNOR U23990 ( .A(y[1268]), .B(x[1268]), .Z(n19416) );
  XOR U23991 ( .A(n19390), .B(n19391), .Z(n19409) );
  XNOR U23992 ( .A(n19406), .B(n19407), .Z(n19391) );
  XNOR U23993 ( .A(n19401), .B(n19402), .Z(n19407) );
  XNOR U23994 ( .A(n19403), .B(n19404), .Z(n19402) );
  XNOR U23995 ( .A(y[1264]), .B(x[1264]), .Z(n19404) );
  XNOR U23996 ( .A(y[1265]), .B(x[1265]), .Z(n19403) );
  XNOR U23997 ( .A(y[1263]), .B(x[1263]), .Z(n19401) );
  XNOR U23998 ( .A(n19395), .B(n19396), .Z(n19406) );
  XNOR U23999 ( .A(y[1260]), .B(x[1260]), .Z(n19396) );
  XNOR U24000 ( .A(n19397), .B(n19398), .Z(n19395) );
  XNOR U24001 ( .A(y[1261]), .B(x[1261]), .Z(n19398) );
  XNOR U24002 ( .A(y[1262]), .B(x[1262]), .Z(n19397) );
  XOR U24003 ( .A(n19389), .B(n19388), .Z(n19390) );
  XNOR U24004 ( .A(n19384), .B(n19385), .Z(n19388) );
  XNOR U24005 ( .A(y[1257]), .B(x[1257]), .Z(n19385) );
  XNOR U24006 ( .A(n19386), .B(n19387), .Z(n19384) );
  XNOR U24007 ( .A(y[1258]), .B(x[1258]), .Z(n19387) );
  XNOR U24008 ( .A(y[1259]), .B(x[1259]), .Z(n19386) );
  XNOR U24009 ( .A(n19378), .B(n19379), .Z(n19389) );
  XNOR U24010 ( .A(y[1254]), .B(x[1254]), .Z(n19379) );
  XNOR U24011 ( .A(n19380), .B(n19381), .Z(n19378) );
  XNOR U24012 ( .A(y[1255]), .B(x[1255]), .Z(n19381) );
  XNOR U24013 ( .A(y[1256]), .B(x[1256]), .Z(n19380) );
  NAND U24014 ( .A(n19445), .B(n19446), .Z(N28557) );
  NANDN U24015 ( .A(n19447), .B(n19448), .Z(n19446) );
  OR U24016 ( .A(n19449), .B(n19450), .Z(n19448) );
  NAND U24017 ( .A(n19449), .B(n19450), .Z(n19445) );
  XOR U24018 ( .A(n19449), .B(n19451), .Z(N28556) );
  XNOR U24019 ( .A(n19447), .B(n19450), .Z(n19451) );
  AND U24020 ( .A(n19452), .B(n19453), .Z(n19450) );
  NANDN U24021 ( .A(n19454), .B(n19455), .Z(n19453) );
  NANDN U24022 ( .A(n19456), .B(n19457), .Z(n19455) );
  NANDN U24023 ( .A(n19457), .B(n19456), .Z(n19452) );
  NAND U24024 ( .A(n19458), .B(n19459), .Z(n19447) );
  NANDN U24025 ( .A(n19460), .B(n19461), .Z(n19459) );
  OR U24026 ( .A(n19462), .B(n19463), .Z(n19461) );
  NAND U24027 ( .A(n19463), .B(n19462), .Z(n19458) );
  AND U24028 ( .A(n19464), .B(n19465), .Z(n19449) );
  NANDN U24029 ( .A(n19466), .B(n19467), .Z(n19465) );
  NANDN U24030 ( .A(n19468), .B(n19469), .Z(n19467) );
  NANDN U24031 ( .A(n19469), .B(n19468), .Z(n19464) );
  XOR U24032 ( .A(n19463), .B(n19470), .Z(N28555) );
  XOR U24033 ( .A(n19460), .B(n19462), .Z(n19470) );
  XNOR U24034 ( .A(n19456), .B(n19471), .Z(n19462) );
  XNOR U24035 ( .A(n19454), .B(n19457), .Z(n19471) );
  NAND U24036 ( .A(n19472), .B(n19473), .Z(n19457) );
  NAND U24037 ( .A(n19474), .B(n19475), .Z(n19473) );
  OR U24038 ( .A(n19476), .B(n19477), .Z(n19474) );
  NANDN U24039 ( .A(n19478), .B(n19476), .Z(n19472) );
  IV U24040 ( .A(n19477), .Z(n19478) );
  NAND U24041 ( .A(n19479), .B(n19480), .Z(n19454) );
  NAND U24042 ( .A(n19481), .B(n19482), .Z(n19480) );
  NANDN U24043 ( .A(n19483), .B(n19484), .Z(n19481) );
  NANDN U24044 ( .A(n19484), .B(n19483), .Z(n19479) );
  AND U24045 ( .A(n19485), .B(n19486), .Z(n19456) );
  NAND U24046 ( .A(n19487), .B(n19488), .Z(n19486) );
  OR U24047 ( .A(n19489), .B(n19490), .Z(n19487) );
  NANDN U24048 ( .A(n19491), .B(n19489), .Z(n19485) );
  NAND U24049 ( .A(n19492), .B(n19493), .Z(n19460) );
  NANDN U24050 ( .A(n19494), .B(n19495), .Z(n19493) );
  OR U24051 ( .A(n19496), .B(n19497), .Z(n19495) );
  NANDN U24052 ( .A(n19498), .B(n19496), .Z(n19492) );
  IV U24053 ( .A(n19497), .Z(n19498) );
  XNOR U24054 ( .A(n19468), .B(n19499), .Z(n19463) );
  XNOR U24055 ( .A(n19466), .B(n19469), .Z(n19499) );
  NAND U24056 ( .A(n19500), .B(n19501), .Z(n19469) );
  NAND U24057 ( .A(n19502), .B(n19503), .Z(n19501) );
  OR U24058 ( .A(n19504), .B(n19505), .Z(n19502) );
  NANDN U24059 ( .A(n19506), .B(n19504), .Z(n19500) );
  IV U24060 ( .A(n19505), .Z(n19506) );
  NAND U24061 ( .A(n19507), .B(n19508), .Z(n19466) );
  NAND U24062 ( .A(n19509), .B(n19510), .Z(n19508) );
  NANDN U24063 ( .A(n19511), .B(n19512), .Z(n19509) );
  NANDN U24064 ( .A(n19512), .B(n19511), .Z(n19507) );
  AND U24065 ( .A(n19513), .B(n19514), .Z(n19468) );
  NAND U24066 ( .A(n19515), .B(n19516), .Z(n19514) );
  OR U24067 ( .A(n19517), .B(n19518), .Z(n19515) );
  NANDN U24068 ( .A(n19519), .B(n19517), .Z(n19513) );
  XNOR U24069 ( .A(n19494), .B(n19520), .Z(N28554) );
  XOR U24070 ( .A(n19496), .B(n19497), .Z(n19520) );
  XNOR U24071 ( .A(n19510), .B(n19521), .Z(n19497) );
  XOR U24072 ( .A(n19511), .B(n19512), .Z(n19521) );
  XOR U24073 ( .A(n19517), .B(n19522), .Z(n19512) );
  XOR U24074 ( .A(n19516), .B(n19519), .Z(n19522) );
  IV U24075 ( .A(n19518), .Z(n19519) );
  NAND U24076 ( .A(n19523), .B(n19524), .Z(n19518) );
  OR U24077 ( .A(n19525), .B(n19526), .Z(n19524) );
  OR U24078 ( .A(n19527), .B(n19528), .Z(n19523) );
  NAND U24079 ( .A(n19529), .B(n19530), .Z(n19516) );
  OR U24080 ( .A(n19531), .B(n19532), .Z(n19530) );
  OR U24081 ( .A(n19533), .B(n19534), .Z(n19529) );
  NOR U24082 ( .A(n19535), .B(n19536), .Z(n19517) );
  ANDN U24083 ( .B(n19537), .A(n19538), .Z(n19511) );
  XNOR U24084 ( .A(n19504), .B(n19539), .Z(n19510) );
  XNOR U24085 ( .A(n19503), .B(n19505), .Z(n19539) );
  NAND U24086 ( .A(n19540), .B(n19541), .Z(n19505) );
  OR U24087 ( .A(n19542), .B(n19543), .Z(n19541) );
  OR U24088 ( .A(n19544), .B(n19545), .Z(n19540) );
  NAND U24089 ( .A(n19546), .B(n19547), .Z(n19503) );
  OR U24090 ( .A(n19548), .B(n19549), .Z(n19547) );
  OR U24091 ( .A(n19550), .B(n19551), .Z(n19546) );
  ANDN U24092 ( .B(n19552), .A(n19553), .Z(n19504) );
  IV U24093 ( .A(n19554), .Z(n19552) );
  ANDN U24094 ( .B(n19555), .A(n19556), .Z(n19496) );
  XOR U24095 ( .A(n19482), .B(n19557), .Z(n19494) );
  XOR U24096 ( .A(n19483), .B(n19484), .Z(n19557) );
  XOR U24097 ( .A(n19489), .B(n19558), .Z(n19484) );
  XOR U24098 ( .A(n19488), .B(n19491), .Z(n19558) );
  IV U24099 ( .A(n19490), .Z(n19491) );
  NAND U24100 ( .A(n19559), .B(n19560), .Z(n19490) );
  OR U24101 ( .A(n19561), .B(n19562), .Z(n19560) );
  OR U24102 ( .A(n19563), .B(n19564), .Z(n19559) );
  NAND U24103 ( .A(n19565), .B(n19566), .Z(n19488) );
  OR U24104 ( .A(n19567), .B(n19568), .Z(n19566) );
  OR U24105 ( .A(n19569), .B(n19570), .Z(n19565) );
  NOR U24106 ( .A(n19571), .B(n19572), .Z(n19489) );
  ANDN U24107 ( .B(n19573), .A(n19574), .Z(n19483) );
  IV U24108 ( .A(n19575), .Z(n19573) );
  XNOR U24109 ( .A(n19476), .B(n19576), .Z(n19482) );
  XNOR U24110 ( .A(n19475), .B(n19477), .Z(n19576) );
  NAND U24111 ( .A(n19577), .B(n19578), .Z(n19477) );
  OR U24112 ( .A(n19579), .B(n19580), .Z(n19578) );
  OR U24113 ( .A(n19581), .B(n19582), .Z(n19577) );
  NAND U24114 ( .A(n19583), .B(n19584), .Z(n19475) );
  OR U24115 ( .A(n19585), .B(n19586), .Z(n19584) );
  OR U24116 ( .A(n19587), .B(n19588), .Z(n19583) );
  ANDN U24117 ( .B(n19589), .A(n19590), .Z(n19476) );
  IV U24118 ( .A(n19591), .Z(n19589) );
  XNOR U24119 ( .A(n19556), .B(n19555), .Z(N28553) );
  XOR U24120 ( .A(n19575), .B(n19574), .Z(n19555) );
  XNOR U24121 ( .A(n19590), .B(n19591), .Z(n19574) );
  XNOR U24122 ( .A(n19585), .B(n19586), .Z(n19591) );
  XNOR U24123 ( .A(n19587), .B(n19588), .Z(n19586) );
  XNOR U24124 ( .A(y[1252]), .B(x[1252]), .Z(n19588) );
  XNOR U24125 ( .A(y[1253]), .B(x[1253]), .Z(n19587) );
  XNOR U24126 ( .A(y[1251]), .B(x[1251]), .Z(n19585) );
  XNOR U24127 ( .A(n19579), .B(n19580), .Z(n19590) );
  XNOR U24128 ( .A(y[1248]), .B(x[1248]), .Z(n19580) );
  XNOR U24129 ( .A(n19581), .B(n19582), .Z(n19579) );
  XNOR U24130 ( .A(y[1249]), .B(x[1249]), .Z(n19582) );
  XNOR U24131 ( .A(y[1250]), .B(x[1250]), .Z(n19581) );
  XNOR U24132 ( .A(n19572), .B(n19571), .Z(n19575) );
  XNOR U24133 ( .A(n19567), .B(n19568), .Z(n19571) );
  XNOR U24134 ( .A(y[1245]), .B(x[1245]), .Z(n19568) );
  XNOR U24135 ( .A(n19569), .B(n19570), .Z(n19567) );
  XNOR U24136 ( .A(y[1246]), .B(x[1246]), .Z(n19570) );
  XNOR U24137 ( .A(y[1247]), .B(x[1247]), .Z(n19569) );
  XNOR U24138 ( .A(n19561), .B(n19562), .Z(n19572) );
  XNOR U24139 ( .A(y[1242]), .B(x[1242]), .Z(n19562) );
  XNOR U24140 ( .A(n19563), .B(n19564), .Z(n19561) );
  XNOR U24141 ( .A(y[1243]), .B(x[1243]), .Z(n19564) );
  XNOR U24142 ( .A(y[1244]), .B(x[1244]), .Z(n19563) );
  XOR U24143 ( .A(n19537), .B(n19538), .Z(n19556) );
  XNOR U24144 ( .A(n19553), .B(n19554), .Z(n19538) );
  XNOR U24145 ( .A(n19548), .B(n19549), .Z(n19554) );
  XNOR U24146 ( .A(n19550), .B(n19551), .Z(n19549) );
  XNOR U24147 ( .A(y[1240]), .B(x[1240]), .Z(n19551) );
  XNOR U24148 ( .A(y[1241]), .B(x[1241]), .Z(n19550) );
  XNOR U24149 ( .A(y[1239]), .B(x[1239]), .Z(n19548) );
  XNOR U24150 ( .A(n19542), .B(n19543), .Z(n19553) );
  XNOR U24151 ( .A(y[1236]), .B(x[1236]), .Z(n19543) );
  XNOR U24152 ( .A(n19544), .B(n19545), .Z(n19542) );
  XNOR U24153 ( .A(y[1237]), .B(x[1237]), .Z(n19545) );
  XNOR U24154 ( .A(y[1238]), .B(x[1238]), .Z(n19544) );
  XOR U24155 ( .A(n19536), .B(n19535), .Z(n19537) );
  XNOR U24156 ( .A(n19531), .B(n19532), .Z(n19535) );
  XNOR U24157 ( .A(y[1233]), .B(x[1233]), .Z(n19532) );
  XNOR U24158 ( .A(n19533), .B(n19534), .Z(n19531) );
  XNOR U24159 ( .A(y[1234]), .B(x[1234]), .Z(n19534) );
  XNOR U24160 ( .A(y[1235]), .B(x[1235]), .Z(n19533) );
  XNOR U24161 ( .A(n19525), .B(n19526), .Z(n19536) );
  XNOR U24162 ( .A(y[1230]), .B(x[1230]), .Z(n19526) );
  XNOR U24163 ( .A(n19527), .B(n19528), .Z(n19525) );
  XNOR U24164 ( .A(y[1231]), .B(x[1231]), .Z(n19528) );
  XNOR U24165 ( .A(y[1232]), .B(x[1232]), .Z(n19527) );
  NAND U24166 ( .A(n19592), .B(n19593), .Z(N28545) );
  NANDN U24167 ( .A(n19594), .B(n19595), .Z(n19593) );
  OR U24168 ( .A(n19596), .B(n19597), .Z(n19595) );
  NAND U24169 ( .A(n19596), .B(n19597), .Z(n19592) );
  XOR U24170 ( .A(n19596), .B(n19598), .Z(N28544) );
  XNOR U24171 ( .A(n19594), .B(n19597), .Z(n19598) );
  AND U24172 ( .A(n19599), .B(n19600), .Z(n19597) );
  NANDN U24173 ( .A(n19601), .B(n19602), .Z(n19600) );
  NANDN U24174 ( .A(n19603), .B(n19604), .Z(n19602) );
  NANDN U24175 ( .A(n19604), .B(n19603), .Z(n19599) );
  NAND U24176 ( .A(n19605), .B(n19606), .Z(n19594) );
  NANDN U24177 ( .A(n19607), .B(n19608), .Z(n19606) );
  OR U24178 ( .A(n19609), .B(n19610), .Z(n19608) );
  NAND U24179 ( .A(n19610), .B(n19609), .Z(n19605) );
  AND U24180 ( .A(n19611), .B(n19612), .Z(n19596) );
  NANDN U24181 ( .A(n19613), .B(n19614), .Z(n19612) );
  NANDN U24182 ( .A(n19615), .B(n19616), .Z(n19614) );
  NANDN U24183 ( .A(n19616), .B(n19615), .Z(n19611) );
  XOR U24184 ( .A(n19610), .B(n19617), .Z(N28543) );
  XOR U24185 ( .A(n19607), .B(n19609), .Z(n19617) );
  XNOR U24186 ( .A(n19603), .B(n19618), .Z(n19609) );
  XNOR U24187 ( .A(n19601), .B(n19604), .Z(n19618) );
  NAND U24188 ( .A(n19619), .B(n19620), .Z(n19604) );
  NAND U24189 ( .A(n19621), .B(n19622), .Z(n19620) );
  OR U24190 ( .A(n19623), .B(n19624), .Z(n19621) );
  NANDN U24191 ( .A(n19625), .B(n19623), .Z(n19619) );
  IV U24192 ( .A(n19624), .Z(n19625) );
  NAND U24193 ( .A(n19626), .B(n19627), .Z(n19601) );
  NAND U24194 ( .A(n19628), .B(n19629), .Z(n19627) );
  NANDN U24195 ( .A(n19630), .B(n19631), .Z(n19628) );
  NANDN U24196 ( .A(n19631), .B(n19630), .Z(n19626) );
  AND U24197 ( .A(n19632), .B(n19633), .Z(n19603) );
  NAND U24198 ( .A(n19634), .B(n19635), .Z(n19633) );
  OR U24199 ( .A(n19636), .B(n19637), .Z(n19634) );
  NANDN U24200 ( .A(n19638), .B(n19636), .Z(n19632) );
  NAND U24201 ( .A(n19639), .B(n19640), .Z(n19607) );
  NANDN U24202 ( .A(n19641), .B(n19642), .Z(n19640) );
  OR U24203 ( .A(n19643), .B(n19644), .Z(n19642) );
  NANDN U24204 ( .A(n19645), .B(n19643), .Z(n19639) );
  IV U24205 ( .A(n19644), .Z(n19645) );
  XNOR U24206 ( .A(n19615), .B(n19646), .Z(n19610) );
  XNOR U24207 ( .A(n19613), .B(n19616), .Z(n19646) );
  NAND U24208 ( .A(n19647), .B(n19648), .Z(n19616) );
  NAND U24209 ( .A(n19649), .B(n19650), .Z(n19648) );
  OR U24210 ( .A(n19651), .B(n19652), .Z(n19649) );
  NANDN U24211 ( .A(n19653), .B(n19651), .Z(n19647) );
  IV U24212 ( .A(n19652), .Z(n19653) );
  NAND U24213 ( .A(n19654), .B(n19655), .Z(n19613) );
  NAND U24214 ( .A(n19656), .B(n19657), .Z(n19655) );
  NANDN U24215 ( .A(n19658), .B(n19659), .Z(n19656) );
  NANDN U24216 ( .A(n19659), .B(n19658), .Z(n19654) );
  AND U24217 ( .A(n19660), .B(n19661), .Z(n19615) );
  NAND U24218 ( .A(n19662), .B(n19663), .Z(n19661) );
  OR U24219 ( .A(n19664), .B(n19665), .Z(n19662) );
  NANDN U24220 ( .A(n19666), .B(n19664), .Z(n19660) );
  XNOR U24221 ( .A(n19641), .B(n19667), .Z(N28542) );
  XOR U24222 ( .A(n19643), .B(n19644), .Z(n19667) );
  XNOR U24223 ( .A(n19657), .B(n19668), .Z(n19644) );
  XOR U24224 ( .A(n19658), .B(n19659), .Z(n19668) );
  XOR U24225 ( .A(n19664), .B(n19669), .Z(n19659) );
  XOR U24226 ( .A(n19663), .B(n19666), .Z(n19669) );
  IV U24227 ( .A(n19665), .Z(n19666) );
  NAND U24228 ( .A(n19670), .B(n19671), .Z(n19665) );
  OR U24229 ( .A(n19672), .B(n19673), .Z(n19671) );
  OR U24230 ( .A(n19674), .B(n19675), .Z(n19670) );
  NAND U24231 ( .A(n19676), .B(n19677), .Z(n19663) );
  OR U24232 ( .A(n19678), .B(n19679), .Z(n19677) );
  OR U24233 ( .A(n19680), .B(n19681), .Z(n19676) );
  NOR U24234 ( .A(n19682), .B(n19683), .Z(n19664) );
  ANDN U24235 ( .B(n19684), .A(n19685), .Z(n19658) );
  XNOR U24236 ( .A(n19651), .B(n19686), .Z(n19657) );
  XNOR U24237 ( .A(n19650), .B(n19652), .Z(n19686) );
  NAND U24238 ( .A(n19687), .B(n19688), .Z(n19652) );
  OR U24239 ( .A(n19689), .B(n19690), .Z(n19688) );
  OR U24240 ( .A(n19691), .B(n19692), .Z(n19687) );
  NAND U24241 ( .A(n19693), .B(n19694), .Z(n19650) );
  OR U24242 ( .A(n19695), .B(n19696), .Z(n19694) );
  OR U24243 ( .A(n19697), .B(n19698), .Z(n19693) );
  ANDN U24244 ( .B(n19699), .A(n19700), .Z(n19651) );
  IV U24245 ( .A(n19701), .Z(n19699) );
  ANDN U24246 ( .B(n19702), .A(n19703), .Z(n19643) );
  XOR U24247 ( .A(n19629), .B(n19704), .Z(n19641) );
  XOR U24248 ( .A(n19630), .B(n19631), .Z(n19704) );
  XOR U24249 ( .A(n19636), .B(n19705), .Z(n19631) );
  XOR U24250 ( .A(n19635), .B(n19638), .Z(n19705) );
  IV U24251 ( .A(n19637), .Z(n19638) );
  NAND U24252 ( .A(n19706), .B(n19707), .Z(n19637) );
  OR U24253 ( .A(n19708), .B(n19709), .Z(n19707) );
  OR U24254 ( .A(n19710), .B(n19711), .Z(n19706) );
  NAND U24255 ( .A(n19712), .B(n19713), .Z(n19635) );
  OR U24256 ( .A(n19714), .B(n19715), .Z(n19713) );
  OR U24257 ( .A(n19716), .B(n19717), .Z(n19712) );
  NOR U24258 ( .A(n19718), .B(n19719), .Z(n19636) );
  ANDN U24259 ( .B(n19720), .A(n19721), .Z(n19630) );
  IV U24260 ( .A(n19722), .Z(n19720) );
  XNOR U24261 ( .A(n19623), .B(n19723), .Z(n19629) );
  XNOR U24262 ( .A(n19622), .B(n19624), .Z(n19723) );
  NAND U24263 ( .A(n19724), .B(n19725), .Z(n19624) );
  OR U24264 ( .A(n19726), .B(n19727), .Z(n19725) );
  OR U24265 ( .A(n19728), .B(n19729), .Z(n19724) );
  NAND U24266 ( .A(n19730), .B(n19731), .Z(n19622) );
  OR U24267 ( .A(n19732), .B(n19733), .Z(n19731) );
  OR U24268 ( .A(n19734), .B(n19735), .Z(n19730) );
  ANDN U24269 ( .B(n19736), .A(n19737), .Z(n19623) );
  IV U24270 ( .A(n19738), .Z(n19736) );
  XNOR U24271 ( .A(n19703), .B(n19702), .Z(N28541) );
  XOR U24272 ( .A(n19722), .B(n19721), .Z(n19702) );
  XNOR U24273 ( .A(n19737), .B(n19738), .Z(n19721) );
  XNOR U24274 ( .A(n19732), .B(n19733), .Z(n19738) );
  XNOR U24275 ( .A(n19734), .B(n19735), .Z(n19733) );
  XNOR U24276 ( .A(y[1228]), .B(x[1228]), .Z(n19735) );
  XNOR U24277 ( .A(y[1229]), .B(x[1229]), .Z(n19734) );
  XNOR U24278 ( .A(y[1227]), .B(x[1227]), .Z(n19732) );
  XNOR U24279 ( .A(n19726), .B(n19727), .Z(n19737) );
  XNOR U24280 ( .A(y[1224]), .B(x[1224]), .Z(n19727) );
  XNOR U24281 ( .A(n19728), .B(n19729), .Z(n19726) );
  XNOR U24282 ( .A(y[1225]), .B(x[1225]), .Z(n19729) );
  XNOR U24283 ( .A(y[1226]), .B(x[1226]), .Z(n19728) );
  XNOR U24284 ( .A(n19719), .B(n19718), .Z(n19722) );
  XNOR U24285 ( .A(n19714), .B(n19715), .Z(n19718) );
  XNOR U24286 ( .A(y[1221]), .B(x[1221]), .Z(n19715) );
  XNOR U24287 ( .A(n19716), .B(n19717), .Z(n19714) );
  XNOR U24288 ( .A(y[1222]), .B(x[1222]), .Z(n19717) );
  XNOR U24289 ( .A(y[1223]), .B(x[1223]), .Z(n19716) );
  XNOR U24290 ( .A(n19708), .B(n19709), .Z(n19719) );
  XNOR U24291 ( .A(y[1218]), .B(x[1218]), .Z(n19709) );
  XNOR U24292 ( .A(n19710), .B(n19711), .Z(n19708) );
  XNOR U24293 ( .A(y[1219]), .B(x[1219]), .Z(n19711) );
  XNOR U24294 ( .A(y[1220]), .B(x[1220]), .Z(n19710) );
  XOR U24295 ( .A(n19684), .B(n19685), .Z(n19703) );
  XNOR U24296 ( .A(n19700), .B(n19701), .Z(n19685) );
  XNOR U24297 ( .A(n19695), .B(n19696), .Z(n19701) );
  XNOR U24298 ( .A(n19697), .B(n19698), .Z(n19696) );
  XNOR U24299 ( .A(y[1216]), .B(x[1216]), .Z(n19698) );
  XNOR U24300 ( .A(y[1217]), .B(x[1217]), .Z(n19697) );
  XNOR U24301 ( .A(y[1215]), .B(x[1215]), .Z(n19695) );
  XNOR U24302 ( .A(n19689), .B(n19690), .Z(n19700) );
  XNOR U24303 ( .A(y[1212]), .B(x[1212]), .Z(n19690) );
  XNOR U24304 ( .A(n19691), .B(n19692), .Z(n19689) );
  XNOR U24305 ( .A(y[1213]), .B(x[1213]), .Z(n19692) );
  XNOR U24306 ( .A(y[1214]), .B(x[1214]), .Z(n19691) );
  XOR U24307 ( .A(n19683), .B(n19682), .Z(n19684) );
  XNOR U24308 ( .A(n19678), .B(n19679), .Z(n19682) );
  XNOR U24309 ( .A(y[1209]), .B(x[1209]), .Z(n19679) );
  XNOR U24310 ( .A(n19680), .B(n19681), .Z(n19678) );
  XNOR U24311 ( .A(y[1210]), .B(x[1210]), .Z(n19681) );
  XNOR U24312 ( .A(y[1211]), .B(x[1211]), .Z(n19680) );
  XNOR U24313 ( .A(n19672), .B(n19673), .Z(n19683) );
  XNOR U24314 ( .A(y[1206]), .B(x[1206]), .Z(n19673) );
  XNOR U24315 ( .A(n19674), .B(n19675), .Z(n19672) );
  XNOR U24316 ( .A(y[1207]), .B(x[1207]), .Z(n19675) );
  XNOR U24317 ( .A(y[1208]), .B(x[1208]), .Z(n19674) );
  NAND U24318 ( .A(n19739), .B(n19740), .Z(N28533) );
  NANDN U24319 ( .A(n19741), .B(n19742), .Z(n19740) );
  OR U24320 ( .A(n19743), .B(n19744), .Z(n19742) );
  NAND U24321 ( .A(n19743), .B(n19744), .Z(n19739) );
  XOR U24322 ( .A(n19743), .B(n19745), .Z(N28532) );
  XNOR U24323 ( .A(n19741), .B(n19744), .Z(n19745) );
  AND U24324 ( .A(n19746), .B(n19747), .Z(n19744) );
  NANDN U24325 ( .A(n19748), .B(n19749), .Z(n19747) );
  NANDN U24326 ( .A(n19750), .B(n19751), .Z(n19749) );
  NANDN U24327 ( .A(n19751), .B(n19750), .Z(n19746) );
  NAND U24328 ( .A(n19752), .B(n19753), .Z(n19741) );
  NANDN U24329 ( .A(n19754), .B(n19755), .Z(n19753) );
  OR U24330 ( .A(n19756), .B(n19757), .Z(n19755) );
  NAND U24331 ( .A(n19757), .B(n19756), .Z(n19752) );
  AND U24332 ( .A(n19758), .B(n19759), .Z(n19743) );
  NANDN U24333 ( .A(n19760), .B(n19761), .Z(n19759) );
  NANDN U24334 ( .A(n19762), .B(n19763), .Z(n19761) );
  NANDN U24335 ( .A(n19763), .B(n19762), .Z(n19758) );
  XOR U24336 ( .A(n19757), .B(n19764), .Z(N28531) );
  XOR U24337 ( .A(n19754), .B(n19756), .Z(n19764) );
  XNOR U24338 ( .A(n19750), .B(n19765), .Z(n19756) );
  XNOR U24339 ( .A(n19748), .B(n19751), .Z(n19765) );
  NAND U24340 ( .A(n19766), .B(n19767), .Z(n19751) );
  NAND U24341 ( .A(n19768), .B(n19769), .Z(n19767) );
  OR U24342 ( .A(n19770), .B(n19771), .Z(n19768) );
  NANDN U24343 ( .A(n19772), .B(n19770), .Z(n19766) );
  IV U24344 ( .A(n19771), .Z(n19772) );
  NAND U24345 ( .A(n19773), .B(n19774), .Z(n19748) );
  NAND U24346 ( .A(n19775), .B(n19776), .Z(n19774) );
  NANDN U24347 ( .A(n19777), .B(n19778), .Z(n19775) );
  NANDN U24348 ( .A(n19778), .B(n19777), .Z(n19773) );
  AND U24349 ( .A(n19779), .B(n19780), .Z(n19750) );
  NAND U24350 ( .A(n19781), .B(n19782), .Z(n19780) );
  OR U24351 ( .A(n19783), .B(n19784), .Z(n19781) );
  NANDN U24352 ( .A(n19785), .B(n19783), .Z(n19779) );
  NAND U24353 ( .A(n19786), .B(n19787), .Z(n19754) );
  NANDN U24354 ( .A(n19788), .B(n19789), .Z(n19787) );
  OR U24355 ( .A(n19790), .B(n19791), .Z(n19789) );
  NANDN U24356 ( .A(n19792), .B(n19790), .Z(n19786) );
  IV U24357 ( .A(n19791), .Z(n19792) );
  XNOR U24358 ( .A(n19762), .B(n19793), .Z(n19757) );
  XNOR U24359 ( .A(n19760), .B(n19763), .Z(n19793) );
  NAND U24360 ( .A(n19794), .B(n19795), .Z(n19763) );
  NAND U24361 ( .A(n19796), .B(n19797), .Z(n19795) );
  OR U24362 ( .A(n19798), .B(n19799), .Z(n19796) );
  NANDN U24363 ( .A(n19800), .B(n19798), .Z(n19794) );
  IV U24364 ( .A(n19799), .Z(n19800) );
  NAND U24365 ( .A(n19801), .B(n19802), .Z(n19760) );
  NAND U24366 ( .A(n19803), .B(n19804), .Z(n19802) );
  NANDN U24367 ( .A(n19805), .B(n19806), .Z(n19803) );
  NANDN U24368 ( .A(n19806), .B(n19805), .Z(n19801) );
  AND U24369 ( .A(n19807), .B(n19808), .Z(n19762) );
  NAND U24370 ( .A(n19809), .B(n19810), .Z(n19808) );
  OR U24371 ( .A(n19811), .B(n19812), .Z(n19809) );
  NANDN U24372 ( .A(n19813), .B(n19811), .Z(n19807) );
  XNOR U24373 ( .A(n19788), .B(n19814), .Z(N28530) );
  XOR U24374 ( .A(n19790), .B(n19791), .Z(n19814) );
  XNOR U24375 ( .A(n19804), .B(n19815), .Z(n19791) );
  XOR U24376 ( .A(n19805), .B(n19806), .Z(n19815) );
  XOR U24377 ( .A(n19811), .B(n19816), .Z(n19806) );
  XOR U24378 ( .A(n19810), .B(n19813), .Z(n19816) );
  IV U24379 ( .A(n19812), .Z(n19813) );
  NAND U24380 ( .A(n19817), .B(n19818), .Z(n19812) );
  OR U24381 ( .A(n19819), .B(n19820), .Z(n19818) );
  OR U24382 ( .A(n19821), .B(n19822), .Z(n19817) );
  NAND U24383 ( .A(n19823), .B(n19824), .Z(n19810) );
  OR U24384 ( .A(n19825), .B(n19826), .Z(n19824) );
  OR U24385 ( .A(n19827), .B(n19828), .Z(n19823) );
  NOR U24386 ( .A(n19829), .B(n19830), .Z(n19811) );
  ANDN U24387 ( .B(n19831), .A(n19832), .Z(n19805) );
  XNOR U24388 ( .A(n19798), .B(n19833), .Z(n19804) );
  XNOR U24389 ( .A(n19797), .B(n19799), .Z(n19833) );
  NAND U24390 ( .A(n19834), .B(n19835), .Z(n19799) );
  OR U24391 ( .A(n19836), .B(n19837), .Z(n19835) );
  OR U24392 ( .A(n19838), .B(n19839), .Z(n19834) );
  NAND U24393 ( .A(n19840), .B(n19841), .Z(n19797) );
  OR U24394 ( .A(n19842), .B(n19843), .Z(n19841) );
  OR U24395 ( .A(n19844), .B(n19845), .Z(n19840) );
  ANDN U24396 ( .B(n19846), .A(n19847), .Z(n19798) );
  IV U24397 ( .A(n19848), .Z(n19846) );
  ANDN U24398 ( .B(n19849), .A(n19850), .Z(n19790) );
  XOR U24399 ( .A(n19776), .B(n19851), .Z(n19788) );
  XOR U24400 ( .A(n19777), .B(n19778), .Z(n19851) );
  XOR U24401 ( .A(n19783), .B(n19852), .Z(n19778) );
  XOR U24402 ( .A(n19782), .B(n19785), .Z(n19852) );
  IV U24403 ( .A(n19784), .Z(n19785) );
  NAND U24404 ( .A(n19853), .B(n19854), .Z(n19784) );
  OR U24405 ( .A(n19855), .B(n19856), .Z(n19854) );
  OR U24406 ( .A(n19857), .B(n19858), .Z(n19853) );
  NAND U24407 ( .A(n19859), .B(n19860), .Z(n19782) );
  OR U24408 ( .A(n19861), .B(n19862), .Z(n19860) );
  OR U24409 ( .A(n19863), .B(n19864), .Z(n19859) );
  NOR U24410 ( .A(n19865), .B(n19866), .Z(n19783) );
  ANDN U24411 ( .B(n19867), .A(n19868), .Z(n19777) );
  IV U24412 ( .A(n19869), .Z(n19867) );
  XNOR U24413 ( .A(n19770), .B(n19870), .Z(n19776) );
  XNOR U24414 ( .A(n19769), .B(n19771), .Z(n19870) );
  NAND U24415 ( .A(n19871), .B(n19872), .Z(n19771) );
  OR U24416 ( .A(n19873), .B(n19874), .Z(n19872) );
  OR U24417 ( .A(n19875), .B(n19876), .Z(n19871) );
  NAND U24418 ( .A(n19877), .B(n19878), .Z(n19769) );
  OR U24419 ( .A(n19879), .B(n19880), .Z(n19878) );
  OR U24420 ( .A(n19881), .B(n19882), .Z(n19877) );
  ANDN U24421 ( .B(n19883), .A(n19884), .Z(n19770) );
  IV U24422 ( .A(n19885), .Z(n19883) );
  XNOR U24423 ( .A(n19850), .B(n19849), .Z(N28529) );
  XOR U24424 ( .A(n19869), .B(n19868), .Z(n19849) );
  XNOR U24425 ( .A(n19884), .B(n19885), .Z(n19868) );
  XNOR U24426 ( .A(n19879), .B(n19880), .Z(n19885) );
  XNOR U24427 ( .A(n19881), .B(n19882), .Z(n19880) );
  XNOR U24428 ( .A(y[1204]), .B(x[1204]), .Z(n19882) );
  XNOR U24429 ( .A(y[1205]), .B(x[1205]), .Z(n19881) );
  XNOR U24430 ( .A(y[1203]), .B(x[1203]), .Z(n19879) );
  XNOR U24431 ( .A(n19873), .B(n19874), .Z(n19884) );
  XNOR U24432 ( .A(y[1200]), .B(x[1200]), .Z(n19874) );
  XNOR U24433 ( .A(n19875), .B(n19876), .Z(n19873) );
  XNOR U24434 ( .A(y[1201]), .B(x[1201]), .Z(n19876) );
  XNOR U24435 ( .A(y[1202]), .B(x[1202]), .Z(n19875) );
  XNOR U24436 ( .A(n19866), .B(n19865), .Z(n19869) );
  XNOR U24437 ( .A(n19861), .B(n19862), .Z(n19865) );
  XNOR U24438 ( .A(y[1197]), .B(x[1197]), .Z(n19862) );
  XNOR U24439 ( .A(n19863), .B(n19864), .Z(n19861) );
  XNOR U24440 ( .A(y[1198]), .B(x[1198]), .Z(n19864) );
  XNOR U24441 ( .A(y[1199]), .B(x[1199]), .Z(n19863) );
  XNOR U24442 ( .A(n19855), .B(n19856), .Z(n19866) );
  XNOR U24443 ( .A(y[1194]), .B(x[1194]), .Z(n19856) );
  XNOR U24444 ( .A(n19857), .B(n19858), .Z(n19855) );
  XNOR U24445 ( .A(y[1195]), .B(x[1195]), .Z(n19858) );
  XNOR U24446 ( .A(y[1196]), .B(x[1196]), .Z(n19857) );
  XOR U24447 ( .A(n19831), .B(n19832), .Z(n19850) );
  XNOR U24448 ( .A(n19847), .B(n19848), .Z(n19832) );
  XNOR U24449 ( .A(n19842), .B(n19843), .Z(n19848) );
  XNOR U24450 ( .A(n19844), .B(n19845), .Z(n19843) );
  XNOR U24451 ( .A(y[1192]), .B(x[1192]), .Z(n19845) );
  XNOR U24452 ( .A(y[1193]), .B(x[1193]), .Z(n19844) );
  XNOR U24453 ( .A(y[1191]), .B(x[1191]), .Z(n19842) );
  XNOR U24454 ( .A(n19836), .B(n19837), .Z(n19847) );
  XNOR U24455 ( .A(y[1188]), .B(x[1188]), .Z(n19837) );
  XNOR U24456 ( .A(n19838), .B(n19839), .Z(n19836) );
  XNOR U24457 ( .A(y[1189]), .B(x[1189]), .Z(n19839) );
  XNOR U24458 ( .A(y[1190]), .B(x[1190]), .Z(n19838) );
  XOR U24459 ( .A(n19830), .B(n19829), .Z(n19831) );
  XNOR U24460 ( .A(n19825), .B(n19826), .Z(n19829) );
  XNOR U24461 ( .A(y[1185]), .B(x[1185]), .Z(n19826) );
  XNOR U24462 ( .A(n19827), .B(n19828), .Z(n19825) );
  XNOR U24463 ( .A(y[1186]), .B(x[1186]), .Z(n19828) );
  XNOR U24464 ( .A(y[1187]), .B(x[1187]), .Z(n19827) );
  XNOR U24465 ( .A(n19819), .B(n19820), .Z(n19830) );
  XNOR U24466 ( .A(y[1182]), .B(x[1182]), .Z(n19820) );
  XNOR U24467 ( .A(n19821), .B(n19822), .Z(n19819) );
  XNOR U24468 ( .A(y[1183]), .B(x[1183]), .Z(n19822) );
  XNOR U24469 ( .A(y[1184]), .B(x[1184]), .Z(n19821) );
  NAND U24470 ( .A(n19886), .B(n19887), .Z(N28521) );
  NANDN U24471 ( .A(n19888), .B(n19889), .Z(n19887) );
  OR U24472 ( .A(n19890), .B(n19891), .Z(n19889) );
  NAND U24473 ( .A(n19890), .B(n19891), .Z(n19886) );
  XOR U24474 ( .A(n19890), .B(n19892), .Z(N28520) );
  XNOR U24475 ( .A(n19888), .B(n19891), .Z(n19892) );
  AND U24476 ( .A(n19893), .B(n19894), .Z(n19891) );
  NANDN U24477 ( .A(n19895), .B(n19896), .Z(n19894) );
  NANDN U24478 ( .A(n19897), .B(n19898), .Z(n19896) );
  NANDN U24479 ( .A(n19898), .B(n19897), .Z(n19893) );
  NAND U24480 ( .A(n19899), .B(n19900), .Z(n19888) );
  NANDN U24481 ( .A(n19901), .B(n19902), .Z(n19900) );
  OR U24482 ( .A(n19903), .B(n19904), .Z(n19902) );
  NAND U24483 ( .A(n19904), .B(n19903), .Z(n19899) );
  AND U24484 ( .A(n19905), .B(n19906), .Z(n19890) );
  NANDN U24485 ( .A(n19907), .B(n19908), .Z(n19906) );
  NANDN U24486 ( .A(n19909), .B(n19910), .Z(n19908) );
  NANDN U24487 ( .A(n19910), .B(n19909), .Z(n19905) );
  XOR U24488 ( .A(n19904), .B(n19911), .Z(N28519) );
  XOR U24489 ( .A(n19901), .B(n19903), .Z(n19911) );
  XNOR U24490 ( .A(n19897), .B(n19912), .Z(n19903) );
  XNOR U24491 ( .A(n19895), .B(n19898), .Z(n19912) );
  NAND U24492 ( .A(n19913), .B(n19914), .Z(n19898) );
  NAND U24493 ( .A(n19915), .B(n19916), .Z(n19914) );
  OR U24494 ( .A(n19917), .B(n19918), .Z(n19915) );
  NANDN U24495 ( .A(n19919), .B(n19917), .Z(n19913) );
  IV U24496 ( .A(n19918), .Z(n19919) );
  NAND U24497 ( .A(n19920), .B(n19921), .Z(n19895) );
  NAND U24498 ( .A(n19922), .B(n19923), .Z(n19921) );
  NANDN U24499 ( .A(n19924), .B(n19925), .Z(n19922) );
  NANDN U24500 ( .A(n19925), .B(n19924), .Z(n19920) );
  AND U24501 ( .A(n19926), .B(n19927), .Z(n19897) );
  NAND U24502 ( .A(n19928), .B(n19929), .Z(n19927) );
  OR U24503 ( .A(n19930), .B(n19931), .Z(n19928) );
  NANDN U24504 ( .A(n19932), .B(n19930), .Z(n19926) );
  NAND U24505 ( .A(n19933), .B(n19934), .Z(n19901) );
  NANDN U24506 ( .A(n19935), .B(n19936), .Z(n19934) );
  OR U24507 ( .A(n19937), .B(n19938), .Z(n19936) );
  NANDN U24508 ( .A(n19939), .B(n19937), .Z(n19933) );
  IV U24509 ( .A(n19938), .Z(n19939) );
  XNOR U24510 ( .A(n19909), .B(n19940), .Z(n19904) );
  XNOR U24511 ( .A(n19907), .B(n19910), .Z(n19940) );
  NAND U24512 ( .A(n19941), .B(n19942), .Z(n19910) );
  NAND U24513 ( .A(n19943), .B(n19944), .Z(n19942) );
  OR U24514 ( .A(n19945), .B(n19946), .Z(n19943) );
  NANDN U24515 ( .A(n19947), .B(n19945), .Z(n19941) );
  IV U24516 ( .A(n19946), .Z(n19947) );
  NAND U24517 ( .A(n19948), .B(n19949), .Z(n19907) );
  NAND U24518 ( .A(n19950), .B(n19951), .Z(n19949) );
  NANDN U24519 ( .A(n19952), .B(n19953), .Z(n19950) );
  NANDN U24520 ( .A(n19953), .B(n19952), .Z(n19948) );
  AND U24521 ( .A(n19954), .B(n19955), .Z(n19909) );
  NAND U24522 ( .A(n19956), .B(n19957), .Z(n19955) );
  OR U24523 ( .A(n19958), .B(n19959), .Z(n19956) );
  NANDN U24524 ( .A(n19960), .B(n19958), .Z(n19954) );
  XNOR U24525 ( .A(n19935), .B(n19961), .Z(N28518) );
  XOR U24526 ( .A(n19937), .B(n19938), .Z(n19961) );
  XNOR U24527 ( .A(n19951), .B(n19962), .Z(n19938) );
  XOR U24528 ( .A(n19952), .B(n19953), .Z(n19962) );
  XOR U24529 ( .A(n19958), .B(n19963), .Z(n19953) );
  XOR U24530 ( .A(n19957), .B(n19960), .Z(n19963) );
  IV U24531 ( .A(n19959), .Z(n19960) );
  NAND U24532 ( .A(n19964), .B(n19965), .Z(n19959) );
  OR U24533 ( .A(n19966), .B(n19967), .Z(n19965) );
  OR U24534 ( .A(n19968), .B(n19969), .Z(n19964) );
  NAND U24535 ( .A(n19970), .B(n19971), .Z(n19957) );
  OR U24536 ( .A(n19972), .B(n19973), .Z(n19971) );
  OR U24537 ( .A(n19974), .B(n19975), .Z(n19970) );
  NOR U24538 ( .A(n19976), .B(n19977), .Z(n19958) );
  ANDN U24539 ( .B(n19978), .A(n19979), .Z(n19952) );
  XNOR U24540 ( .A(n19945), .B(n19980), .Z(n19951) );
  XNOR U24541 ( .A(n19944), .B(n19946), .Z(n19980) );
  NAND U24542 ( .A(n19981), .B(n19982), .Z(n19946) );
  OR U24543 ( .A(n19983), .B(n19984), .Z(n19982) );
  OR U24544 ( .A(n19985), .B(n19986), .Z(n19981) );
  NAND U24545 ( .A(n19987), .B(n19988), .Z(n19944) );
  OR U24546 ( .A(n19989), .B(n19990), .Z(n19988) );
  OR U24547 ( .A(n19991), .B(n19992), .Z(n19987) );
  ANDN U24548 ( .B(n19993), .A(n19994), .Z(n19945) );
  IV U24549 ( .A(n19995), .Z(n19993) );
  ANDN U24550 ( .B(n19996), .A(n19997), .Z(n19937) );
  XOR U24551 ( .A(n19923), .B(n19998), .Z(n19935) );
  XOR U24552 ( .A(n19924), .B(n19925), .Z(n19998) );
  XOR U24553 ( .A(n19930), .B(n19999), .Z(n19925) );
  XOR U24554 ( .A(n19929), .B(n19932), .Z(n19999) );
  IV U24555 ( .A(n19931), .Z(n19932) );
  NAND U24556 ( .A(n20000), .B(n20001), .Z(n19931) );
  OR U24557 ( .A(n20002), .B(n20003), .Z(n20001) );
  OR U24558 ( .A(n20004), .B(n20005), .Z(n20000) );
  NAND U24559 ( .A(n20006), .B(n20007), .Z(n19929) );
  OR U24560 ( .A(n20008), .B(n20009), .Z(n20007) );
  OR U24561 ( .A(n20010), .B(n20011), .Z(n20006) );
  NOR U24562 ( .A(n20012), .B(n20013), .Z(n19930) );
  ANDN U24563 ( .B(n20014), .A(n20015), .Z(n19924) );
  IV U24564 ( .A(n20016), .Z(n20014) );
  XNOR U24565 ( .A(n19917), .B(n20017), .Z(n19923) );
  XNOR U24566 ( .A(n19916), .B(n19918), .Z(n20017) );
  NAND U24567 ( .A(n20018), .B(n20019), .Z(n19918) );
  OR U24568 ( .A(n20020), .B(n20021), .Z(n20019) );
  OR U24569 ( .A(n20022), .B(n20023), .Z(n20018) );
  NAND U24570 ( .A(n20024), .B(n20025), .Z(n19916) );
  OR U24571 ( .A(n20026), .B(n20027), .Z(n20025) );
  OR U24572 ( .A(n20028), .B(n20029), .Z(n20024) );
  ANDN U24573 ( .B(n20030), .A(n20031), .Z(n19917) );
  IV U24574 ( .A(n20032), .Z(n20030) );
  XNOR U24575 ( .A(n19997), .B(n19996), .Z(N28517) );
  XOR U24576 ( .A(n20016), .B(n20015), .Z(n19996) );
  XNOR U24577 ( .A(n20031), .B(n20032), .Z(n20015) );
  XNOR U24578 ( .A(n20026), .B(n20027), .Z(n20032) );
  XNOR U24579 ( .A(n20028), .B(n20029), .Z(n20027) );
  XNOR U24580 ( .A(y[1180]), .B(x[1180]), .Z(n20029) );
  XNOR U24581 ( .A(y[1181]), .B(x[1181]), .Z(n20028) );
  XNOR U24582 ( .A(y[1179]), .B(x[1179]), .Z(n20026) );
  XNOR U24583 ( .A(n20020), .B(n20021), .Z(n20031) );
  XNOR U24584 ( .A(y[1176]), .B(x[1176]), .Z(n20021) );
  XNOR U24585 ( .A(n20022), .B(n20023), .Z(n20020) );
  XNOR U24586 ( .A(y[1177]), .B(x[1177]), .Z(n20023) );
  XNOR U24587 ( .A(y[1178]), .B(x[1178]), .Z(n20022) );
  XNOR U24588 ( .A(n20013), .B(n20012), .Z(n20016) );
  XNOR U24589 ( .A(n20008), .B(n20009), .Z(n20012) );
  XNOR U24590 ( .A(y[1173]), .B(x[1173]), .Z(n20009) );
  XNOR U24591 ( .A(n20010), .B(n20011), .Z(n20008) );
  XNOR U24592 ( .A(y[1174]), .B(x[1174]), .Z(n20011) );
  XNOR U24593 ( .A(y[1175]), .B(x[1175]), .Z(n20010) );
  XNOR U24594 ( .A(n20002), .B(n20003), .Z(n20013) );
  XNOR U24595 ( .A(y[1170]), .B(x[1170]), .Z(n20003) );
  XNOR U24596 ( .A(n20004), .B(n20005), .Z(n20002) );
  XNOR U24597 ( .A(y[1171]), .B(x[1171]), .Z(n20005) );
  XNOR U24598 ( .A(y[1172]), .B(x[1172]), .Z(n20004) );
  XOR U24599 ( .A(n19978), .B(n19979), .Z(n19997) );
  XNOR U24600 ( .A(n19994), .B(n19995), .Z(n19979) );
  XNOR U24601 ( .A(n19989), .B(n19990), .Z(n19995) );
  XNOR U24602 ( .A(n19991), .B(n19992), .Z(n19990) );
  XNOR U24603 ( .A(y[1168]), .B(x[1168]), .Z(n19992) );
  XNOR U24604 ( .A(y[1169]), .B(x[1169]), .Z(n19991) );
  XNOR U24605 ( .A(y[1167]), .B(x[1167]), .Z(n19989) );
  XNOR U24606 ( .A(n19983), .B(n19984), .Z(n19994) );
  XNOR U24607 ( .A(y[1164]), .B(x[1164]), .Z(n19984) );
  XNOR U24608 ( .A(n19985), .B(n19986), .Z(n19983) );
  XNOR U24609 ( .A(y[1165]), .B(x[1165]), .Z(n19986) );
  XNOR U24610 ( .A(y[1166]), .B(x[1166]), .Z(n19985) );
  XOR U24611 ( .A(n19977), .B(n19976), .Z(n19978) );
  XNOR U24612 ( .A(n19972), .B(n19973), .Z(n19976) );
  XNOR U24613 ( .A(y[1161]), .B(x[1161]), .Z(n19973) );
  XNOR U24614 ( .A(n19974), .B(n19975), .Z(n19972) );
  XNOR U24615 ( .A(y[1162]), .B(x[1162]), .Z(n19975) );
  XNOR U24616 ( .A(y[1163]), .B(x[1163]), .Z(n19974) );
  XNOR U24617 ( .A(n19966), .B(n19967), .Z(n19977) );
  XNOR U24618 ( .A(y[1158]), .B(x[1158]), .Z(n19967) );
  XNOR U24619 ( .A(n19968), .B(n19969), .Z(n19966) );
  XNOR U24620 ( .A(y[1159]), .B(x[1159]), .Z(n19969) );
  XNOR U24621 ( .A(y[1160]), .B(x[1160]), .Z(n19968) );
  NAND U24622 ( .A(n20033), .B(n20034), .Z(N28509) );
  NANDN U24623 ( .A(n20035), .B(n20036), .Z(n20034) );
  OR U24624 ( .A(n20037), .B(n20038), .Z(n20036) );
  NAND U24625 ( .A(n20037), .B(n20038), .Z(n20033) );
  XOR U24626 ( .A(n20037), .B(n20039), .Z(N28508) );
  XNOR U24627 ( .A(n20035), .B(n20038), .Z(n20039) );
  AND U24628 ( .A(n20040), .B(n20041), .Z(n20038) );
  NANDN U24629 ( .A(n20042), .B(n20043), .Z(n20041) );
  NANDN U24630 ( .A(n20044), .B(n20045), .Z(n20043) );
  NANDN U24631 ( .A(n20045), .B(n20044), .Z(n20040) );
  NAND U24632 ( .A(n20046), .B(n20047), .Z(n20035) );
  NANDN U24633 ( .A(n20048), .B(n20049), .Z(n20047) );
  OR U24634 ( .A(n20050), .B(n20051), .Z(n20049) );
  NAND U24635 ( .A(n20051), .B(n20050), .Z(n20046) );
  AND U24636 ( .A(n20052), .B(n20053), .Z(n20037) );
  NANDN U24637 ( .A(n20054), .B(n20055), .Z(n20053) );
  NANDN U24638 ( .A(n20056), .B(n20057), .Z(n20055) );
  NANDN U24639 ( .A(n20057), .B(n20056), .Z(n20052) );
  XOR U24640 ( .A(n20051), .B(n20058), .Z(N28507) );
  XOR U24641 ( .A(n20048), .B(n20050), .Z(n20058) );
  XNOR U24642 ( .A(n20044), .B(n20059), .Z(n20050) );
  XNOR U24643 ( .A(n20042), .B(n20045), .Z(n20059) );
  NAND U24644 ( .A(n20060), .B(n20061), .Z(n20045) );
  NAND U24645 ( .A(n20062), .B(n20063), .Z(n20061) );
  OR U24646 ( .A(n20064), .B(n20065), .Z(n20062) );
  NANDN U24647 ( .A(n20066), .B(n20064), .Z(n20060) );
  IV U24648 ( .A(n20065), .Z(n20066) );
  NAND U24649 ( .A(n20067), .B(n20068), .Z(n20042) );
  NAND U24650 ( .A(n20069), .B(n20070), .Z(n20068) );
  NANDN U24651 ( .A(n20071), .B(n20072), .Z(n20069) );
  NANDN U24652 ( .A(n20072), .B(n20071), .Z(n20067) );
  AND U24653 ( .A(n20073), .B(n20074), .Z(n20044) );
  NAND U24654 ( .A(n20075), .B(n20076), .Z(n20074) );
  OR U24655 ( .A(n20077), .B(n20078), .Z(n20075) );
  NANDN U24656 ( .A(n20079), .B(n20077), .Z(n20073) );
  NAND U24657 ( .A(n20080), .B(n20081), .Z(n20048) );
  NANDN U24658 ( .A(n20082), .B(n20083), .Z(n20081) );
  OR U24659 ( .A(n20084), .B(n20085), .Z(n20083) );
  NANDN U24660 ( .A(n20086), .B(n20084), .Z(n20080) );
  IV U24661 ( .A(n20085), .Z(n20086) );
  XNOR U24662 ( .A(n20056), .B(n20087), .Z(n20051) );
  XNOR U24663 ( .A(n20054), .B(n20057), .Z(n20087) );
  NAND U24664 ( .A(n20088), .B(n20089), .Z(n20057) );
  NAND U24665 ( .A(n20090), .B(n20091), .Z(n20089) );
  OR U24666 ( .A(n20092), .B(n20093), .Z(n20090) );
  NANDN U24667 ( .A(n20094), .B(n20092), .Z(n20088) );
  IV U24668 ( .A(n20093), .Z(n20094) );
  NAND U24669 ( .A(n20095), .B(n20096), .Z(n20054) );
  NAND U24670 ( .A(n20097), .B(n20098), .Z(n20096) );
  NANDN U24671 ( .A(n20099), .B(n20100), .Z(n20097) );
  NANDN U24672 ( .A(n20100), .B(n20099), .Z(n20095) );
  AND U24673 ( .A(n20101), .B(n20102), .Z(n20056) );
  NAND U24674 ( .A(n20103), .B(n20104), .Z(n20102) );
  OR U24675 ( .A(n20105), .B(n20106), .Z(n20103) );
  NANDN U24676 ( .A(n20107), .B(n20105), .Z(n20101) );
  XNOR U24677 ( .A(n20082), .B(n20108), .Z(N28506) );
  XOR U24678 ( .A(n20084), .B(n20085), .Z(n20108) );
  XNOR U24679 ( .A(n20098), .B(n20109), .Z(n20085) );
  XOR U24680 ( .A(n20099), .B(n20100), .Z(n20109) );
  XOR U24681 ( .A(n20105), .B(n20110), .Z(n20100) );
  XOR U24682 ( .A(n20104), .B(n20107), .Z(n20110) );
  IV U24683 ( .A(n20106), .Z(n20107) );
  NAND U24684 ( .A(n20111), .B(n20112), .Z(n20106) );
  OR U24685 ( .A(n20113), .B(n20114), .Z(n20112) );
  OR U24686 ( .A(n20115), .B(n20116), .Z(n20111) );
  NAND U24687 ( .A(n20117), .B(n20118), .Z(n20104) );
  OR U24688 ( .A(n20119), .B(n20120), .Z(n20118) );
  OR U24689 ( .A(n20121), .B(n20122), .Z(n20117) );
  NOR U24690 ( .A(n20123), .B(n20124), .Z(n20105) );
  ANDN U24691 ( .B(n20125), .A(n20126), .Z(n20099) );
  XNOR U24692 ( .A(n20092), .B(n20127), .Z(n20098) );
  XNOR U24693 ( .A(n20091), .B(n20093), .Z(n20127) );
  NAND U24694 ( .A(n20128), .B(n20129), .Z(n20093) );
  OR U24695 ( .A(n20130), .B(n20131), .Z(n20129) );
  OR U24696 ( .A(n20132), .B(n20133), .Z(n20128) );
  NAND U24697 ( .A(n20134), .B(n20135), .Z(n20091) );
  OR U24698 ( .A(n20136), .B(n20137), .Z(n20135) );
  OR U24699 ( .A(n20138), .B(n20139), .Z(n20134) );
  ANDN U24700 ( .B(n20140), .A(n20141), .Z(n20092) );
  IV U24701 ( .A(n20142), .Z(n20140) );
  ANDN U24702 ( .B(n20143), .A(n20144), .Z(n20084) );
  XOR U24703 ( .A(n20070), .B(n20145), .Z(n20082) );
  XOR U24704 ( .A(n20071), .B(n20072), .Z(n20145) );
  XOR U24705 ( .A(n20077), .B(n20146), .Z(n20072) );
  XOR U24706 ( .A(n20076), .B(n20079), .Z(n20146) );
  IV U24707 ( .A(n20078), .Z(n20079) );
  NAND U24708 ( .A(n20147), .B(n20148), .Z(n20078) );
  OR U24709 ( .A(n20149), .B(n20150), .Z(n20148) );
  OR U24710 ( .A(n20151), .B(n20152), .Z(n20147) );
  NAND U24711 ( .A(n20153), .B(n20154), .Z(n20076) );
  OR U24712 ( .A(n20155), .B(n20156), .Z(n20154) );
  OR U24713 ( .A(n20157), .B(n20158), .Z(n20153) );
  NOR U24714 ( .A(n20159), .B(n20160), .Z(n20077) );
  ANDN U24715 ( .B(n20161), .A(n20162), .Z(n20071) );
  IV U24716 ( .A(n20163), .Z(n20161) );
  XNOR U24717 ( .A(n20064), .B(n20164), .Z(n20070) );
  XNOR U24718 ( .A(n20063), .B(n20065), .Z(n20164) );
  NAND U24719 ( .A(n20165), .B(n20166), .Z(n20065) );
  OR U24720 ( .A(n20167), .B(n20168), .Z(n20166) );
  OR U24721 ( .A(n20169), .B(n20170), .Z(n20165) );
  NAND U24722 ( .A(n20171), .B(n20172), .Z(n20063) );
  OR U24723 ( .A(n20173), .B(n20174), .Z(n20172) );
  OR U24724 ( .A(n20175), .B(n20176), .Z(n20171) );
  ANDN U24725 ( .B(n20177), .A(n20178), .Z(n20064) );
  IV U24726 ( .A(n20179), .Z(n20177) );
  XNOR U24727 ( .A(n20144), .B(n20143), .Z(N28505) );
  XOR U24728 ( .A(n20163), .B(n20162), .Z(n20143) );
  XNOR U24729 ( .A(n20178), .B(n20179), .Z(n20162) );
  XNOR U24730 ( .A(n20173), .B(n20174), .Z(n20179) );
  XNOR U24731 ( .A(n20175), .B(n20176), .Z(n20174) );
  XNOR U24732 ( .A(y[1156]), .B(x[1156]), .Z(n20176) );
  XNOR U24733 ( .A(y[1157]), .B(x[1157]), .Z(n20175) );
  XNOR U24734 ( .A(y[1155]), .B(x[1155]), .Z(n20173) );
  XNOR U24735 ( .A(n20167), .B(n20168), .Z(n20178) );
  XNOR U24736 ( .A(y[1152]), .B(x[1152]), .Z(n20168) );
  XNOR U24737 ( .A(n20169), .B(n20170), .Z(n20167) );
  XNOR U24738 ( .A(y[1153]), .B(x[1153]), .Z(n20170) );
  XNOR U24739 ( .A(y[1154]), .B(x[1154]), .Z(n20169) );
  XNOR U24740 ( .A(n20160), .B(n20159), .Z(n20163) );
  XNOR U24741 ( .A(n20155), .B(n20156), .Z(n20159) );
  XNOR U24742 ( .A(y[1149]), .B(x[1149]), .Z(n20156) );
  XNOR U24743 ( .A(n20157), .B(n20158), .Z(n20155) );
  XNOR U24744 ( .A(y[1150]), .B(x[1150]), .Z(n20158) );
  XNOR U24745 ( .A(y[1151]), .B(x[1151]), .Z(n20157) );
  XNOR U24746 ( .A(n20149), .B(n20150), .Z(n20160) );
  XNOR U24747 ( .A(y[1146]), .B(x[1146]), .Z(n20150) );
  XNOR U24748 ( .A(n20151), .B(n20152), .Z(n20149) );
  XNOR U24749 ( .A(y[1147]), .B(x[1147]), .Z(n20152) );
  XNOR U24750 ( .A(y[1148]), .B(x[1148]), .Z(n20151) );
  XOR U24751 ( .A(n20125), .B(n20126), .Z(n20144) );
  XNOR U24752 ( .A(n20141), .B(n20142), .Z(n20126) );
  XNOR U24753 ( .A(n20136), .B(n20137), .Z(n20142) );
  XNOR U24754 ( .A(n20138), .B(n20139), .Z(n20137) );
  XNOR U24755 ( .A(y[1144]), .B(x[1144]), .Z(n20139) );
  XNOR U24756 ( .A(y[1145]), .B(x[1145]), .Z(n20138) );
  XNOR U24757 ( .A(y[1143]), .B(x[1143]), .Z(n20136) );
  XNOR U24758 ( .A(n20130), .B(n20131), .Z(n20141) );
  XNOR U24759 ( .A(y[1140]), .B(x[1140]), .Z(n20131) );
  XNOR U24760 ( .A(n20132), .B(n20133), .Z(n20130) );
  XNOR U24761 ( .A(y[1141]), .B(x[1141]), .Z(n20133) );
  XNOR U24762 ( .A(y[1142]), .B(x[1142]), .Z(n20132) );
  XOR U24763 ( .A(n20124), .B(n20123), .Z(n20125) );
  XNOR U24764 ( .A(n20119), .B(n20120), .Z(n20123) );
  XNOR U24765 ( .A(y[1137]), .B(x[1137]), .Z(n20120) );
  XNOR U24766 ( .A(n20121), .B(n20122), .Z(n20119) );
  XNOR U24767 ( .A(y[1138]), .B(x[1138]), .Z(n20122) );
  XNOR U24768 ( .A(y[1139]), .B(x[1139]), .Z(n20121) );
  XNOR U24769 ( .A(n20113), .B(n20114), .Z(n20124) );
  XNOR U24770 ( .A(y[1134]), .B(x[1134]), .Z(n20114) );
  XNOR U24771 ( .A(n20115), .B(n20116), .Z(n20113) );
  XNOR U24772 ( .A(y[1135]), .B(x[1135]), .Z(n20116) );
  XNOR U24773 ( .A(y[1136]), .B(x[1136]), .Z(n20115) );
  NAND U24774 ( .A(n20180), .B(n20181), .Z(N28497) );
  NANDN U24775 ( .A(n20182), .B(n20183), .Z(n20181) );
  OR U24776 ( .A(n20184), .B(n20185), .Z(n20183) );
  NAND U24777 ( .A(n20184), .B(n20185), .Z(n20180) );
  XOR U24778 ( .A(n20184), .B(n20186), .Z(N28496) );
  XNOR U24779 ( .A(n20182), .B(n20185), .Z(n20186) );
  AND U24780 ( .A(n20187), .B(n20188), .Z(n20185) );
  NANDN U24781 ( .A(n20189), .B(n20190), .Z(n20188) );
  NANDN U24782 ( .A(n20191), .B(n20192), .Z(n20190) );
  NANDN U24783 ( .A(n20192), .B(n20191), .Z(n20187) );
  NAND U24784 ( .A(n20193), .B(n20194), .Z(n20182) );
  NANDN U24785 ( .A(n20195), .B(n20196), .Z(n20194) );
  OR U24786 ( .A(n20197), .B(n20198), .Z(n20196) );
  NAND U24787 ( .A(n20198), .B(n20197), .Z(n20193) );
  AND U24788 ( .A(n20199), .B(n20200), .Z(n20184) );
  NANDN U24789 ( .A(n20201), .B(n20202), .Z(n20200) );
  NANDN U24790 ( .A(n20203), .B(n20204), .Z(n20202) );
  NANDN U24791 ( .A(n20204), .B(n20203), .Z(n20199) );
  XOR U24792 ( .A(n20198), .B(n20205), .Z(N28495) );
  XOR U24793 ( .A(n20195), .B(n20197), .Z(n20205) );
  XNOR U24794 ( .A(n20191), .B(n20206), .Z(n20197) );
  XNOR U24795 ( .A(n20189), .B(n20192), .Z(n20206) );
  NAND U24796 ( .A(n20207), .B(n20208), .Z(n20192) );
  NAND U24797 ( .A(n20209), .B(n20210), .Z(n20208) );
  OR U24798 ( .A(n20211), .B(n20212), .Z(n20209) );
  NANDN U24799 ( .A(n20213), .B(n20211), .Z(n20207) );
  IV U24800 ( .A(n20212), .Z(n20213) );
  NAND U24801 ( .A(n20214), .B(n20215), .Z(n20189) );
  NAND U24802 ( .A(n20216), .B(n20217), .Z(n20215) );
  NANDN U24803 ( .A(n20218), .B(n20219), .Z(n20216) );
  NANDN U24804 ( .A(n20219), .B(n20218), .Z(n20214) );
  AND U24805 ( .A(n20220), .B(n20221), .Z(n20191) );
  NAND U24806 ( .A(n20222), .B(n20223), .Z(n20221) );
  OR U24807 ( .A(n20224), .B(n20225), .Z(n20222) );
  NANDN U24808 ( .A(n20226), .B(n20224), .Z(n20220) );
  NAND U24809 ( .A(n20227), .B(n20228), .Z(n20195) );
  NANDN U24810 ( .A(n20229), .B(n20230), .Z(n20228) );
  OR U24811 ( .A(n20231), .B(n20232), .Z(n20230) );
  NANDN U24812 ( .A(n20233), .B(n20231), .Z(n20227) );
  IV U24813 ( .A(n20232), .Z(n20233) );
  XNOR U24814 ( .A(n20203), .B(n20234), .Z(n20198) );
  XNOR U24815 ( .A(n20201), .B(n20204), .Z(n20234) );
  NAND U24816 ( .A(n20235), .B(n20236), .Z(n20204) );
  NAND U24817 ( .A(n20237), .B(n20238), .Z(n20236) );
  OR U24818 ( .A(n20239), .B(n20240), .Z(n20237) );
  NANDN U24819 ( .A(n20241), .B(n20239), .Z(n20235) );
  IV U24820 ( .A(n20240), .Z(n20241) );
  NAND U24821 ( .A(n20242), .B(n20243), .Z(n20201) );
  NAND U24822 ( .A(n20244), .B(n20245), .Z(n20243) );
  NANDN U24823 ( .A(n20246), .B(n20247), .Z(n20244) );
  NANDN U24824 ( .A(n20247), .B(n20246), .Z(n20242) );
  AND U24825 ( .A(n20248), .B(n20249), .Z(n20203) );
  NAND U24826 ( .A(n20250), .B(n20251), .Z(n20249) );
  OR U24827 ( .A(n20252), .B(n20253), .Z(n20250) );
  NANDN U24828 ( .A(n20254), .B(n20252), .Z(n20248) );
  XNOR U24829 ( .A(n20229), .B(n20255), .Z(N28494) );
  XOR U24830 ( .A(n20231), .B(n20232), .Z(n20255) );
  XNOR U24831 ( .A(n20245), .B(n20256), .Z(n20232) );
  XOR U24832 ( .A(n20246), .B(n20247), .Z(n20256) );
  XOR U24833 ( .A(n20252), .B(n20257), .Z(n20247) );
  XOR U24834 ( .A(n20251), .B(n20254), .Z(n20257) );
  IV U24835 ( .A(n20253), .Z(n20254) );
  NAND U24836 ( .A(n20258), .B(n20259), .Z(n20253) );
  OR U24837 ( .A(n20260), .B(n20261), .Z(n20259) );
  OR U24838 ( .A(n20262), .B(n20263), .Z(n20258) );
  NAND U24839 ( .A(n20264), .B(n20265), .Z(n20251) );
  OR U24840 ( .A(n20266), .B(n20267), .Z(n20265) );
  OR U24841 ( .A(n20268), .B(n20269), .Z(n20264) );
  NOR U24842 ( .A(n20270), .B(n20271), .Z(n20252) );
  ANDN U24843 ( .B(n20272), .A(n20273), .Z(n20246) );
  XNOR U24844 ( .A(n20239), .B(n20274), .Z(n20245) );
  XNOR U24845 ( .A(n20238), .B(n20240), .Z(n20274) );
  NAND U24846 ( .A(n20275), .B(n20276), .Z(n20240) );
  OR U24847 ( .A(n20277), .B(n20278), .Z(n20276) );
  OR U24848 ( .A(n20279), .B(n20280), .Z(n20275) );
  NAND U24849 ( .A(n20281), .B(n20282), .Z(n20238) );
  OR U24850 ( .A(n20283), .B(n20284), .Z(n20282) );
  OR U24851 ( .A(n20285), .B(n20286), .Z(n20281) );
  ANDN U24852 ( .B(n20287), .A(n20288), .Z(n20239) );
  IV U24853 ( .A(n20289), .Z(n20287) );
  ANDN U24854 ( .B(n20290), .A(n20291), .Z(n20231) );
  XOR U24855 ( .A(n20217), .B(n20292), .Z(n20229) );
  XOR U24856 ( .A(n20218), .B(n20219), .Z(n20292) );
  XOR U24857 ( .A(n20224), .B(n20293), .Z(n20219) );
  XOR U24858 ( .A(n20223), .B(n20226), .Z(n20293) );
  IV U24859 ( .A(n20225), .Z(n20226) );
  NAND U24860 ( .A(n20294), .B(n20295), .Z(n20225) );
  OR U24861 ( .A(n20296), .B(n20297), .Z(n20295) );
  OR U24862 ( .A(n20298), .B(n20299), .Z(n20294) );
  NAND U24863 ( .A(n20300), .B(n20301), .Z(n20223) );
  OR U24864 ( .A(n20302), .B(n20303), .Z(n20301) );
  OR U24865 ( .A(n20304), .B(n20305), .Z(n20300) );
  NOR U24866 ( .A(n20306), .B(n20307), .Z(n20224) );
  ANDN U24867 ( .B(n20308), .A(n20309), .Z(n20218) );
  IV U24868 ( .A(n20310), .Z(n20308) );
  XNOR U24869 ( .A(n20211), .B(n20311), .Z(n20217) );
  XNOR U24870 ( .A(n20210), .B(n20212), .Z(n20311) );
  NAND U24871 ( .A(n20312), .B(n20313), .Z(n20212) );
  OR U24872 ( .A(n20314), .B(n20315), .Z(n20313) );
  OR U24873 ( .A(n20316), .B(n20317), .Z(n20312) );
  NAND U24874 ( .A(n20318), .B(n20319), .Z(n20210) );
  OR U24875 ( .A(n20320), .B(n20321), .Z(n20319) );
  OR U24876 ( .A(n20322), .B(n20323), .Z(n20318) );
  ANDN U24877 ( .B(n20324), .A(n20325), .Z(n20211) );
  IV U24878 ( .A(n20326), .Z(n20324) );
  XNOR U24879 ( .A(n20291), .B(n20290), .Z(N28493) );
  XOR U24880 ( .A(n20310), .B(n20309), .Z(n20290) );
  XNOR U24881 ( .A(n20325), .B(n20326), .Z(n20309) );
  XNOR U24882 ( .A(n20320), .B(n20321), .Z(n20326) );
  XNOR U24883 ( .A(n20322), .B(n20323), .Z(n20321) );
  XNOR U24884 ( .A(y[1132]), .B(x[1132]), .Z(n20323) );
  XNOR U24885 ( .A(y[1133]), .B(x[1133]), .Z(n20322) );
  XNOR U24886 ( .A(y[1131]), .B(x[1131]), .Z(n20320) );
  XNOR U24887 ( .A(n20314), .B(n20315), .Z(n20325) );
  XNOR U24888 ( .A(y[1128]), .B(x[1128]), .Z(n20315) );
  XNOR U24889 ( .A(n20316), .B(n20317), .Z(n20314) );
  XNOR U24890 ( .A(y[1129]), .B(x[1129]), .Z(n20317) );
  XNOR U24891 ( .A(y[1130]), .B(x[1130]), .Z(n20316) );
  XNOR U24892 ( .A(n20307), .B(n20306), .Z(n20310) );
  XNOR U24893 ( .A(n20302), .B(n20303), .Z(n20306) );
  XNOR U24894 ( .A(y[1125]), .B(x[1125]), .Z(n20303) );
  XNOR U24895 ( .A(n20304), .B(n20305), .Z(n20302) );
  XNOR U24896 ( .A(y[1126]), .B(x[1126]), .Z(n20305) );
  XNOR U24897 ( .A(y[1127]), .B(x[1127]), .Z(n20304) );
  XNOR U24898 ( .A(n20296), .B(n20297), .Z(n20307) );
  XNOR U24899 ( .A(y[1122]), .B(x[1122]), .Z(n20297) );
  XNOR U24900 ( .A(n20298), .B(n20299), .Z(n20296) );
  XNOR U24901 ( .A(y[1123]), .B(x[1123]), .Z(n20299) );
  XNOR U24902 ( .A(y[1124]), .B(x[1124]), .Z(n20298) );
  XOR U24903 ( .A(n20272), .B(n20273), .Z(n20291) );
  XNOR U24904 ( .A(n20288), .B(n20289), .Z(n20273) );
  XNOR U24905 ( .A(n20283), .B(n20284), .Z(n20289) );
  XNOR U24906 ( .A(n20285), .B(n20286), .Z(n20284) );
  XNOR U24907 ( .A(y[1120]), .B(x[1120]), .Z(n20286) );
  XNOR U24908 ( .A(y[1121]), .B(x[1121]), .Z(n20285) );
  XNOR U24909 ( .A(y[1119]), .B(x[1119]), .Z(n20283) );
  XNOR U24910 ( .A(n20277), .B(n20278), .Z(n20288) );
  XNOR U24911 ( .A(y[1116]), .B(x[1116]), .Z(n20278) );
  XNOR U24912 ( .A(n20279), .B(n20280), .Z(n20277) );
  XNOR U24913 ( .A(y[1117]), .B(x[1117]), .Z(n20280) );
  XNOR U24914 ( .A(y[1118]), .B(x[1118]), .Z(n20279) );
  XOR U24915 ( .A(n20271), .B(n20270), .Z(n20272) );
  XNOR U24916 ( .A(n20266), .B(n20267), .Z(n20270) );
  XNOR U24917 ( .A(y[1113]), .B(x[1113]), .Z(n20267) );
  XNOR U24918 ( .A(n20268), .B(n20269), .Z(n20266) );
  XNOR U24919 ( .A(y[1114]), .B(x[1114]), .Z(n20269) );
  XNOR U24920 ( .A(y[1115]), .B(x[1115]), .Z(n20268) );
  XNOR U24921 ( .A(n20260), .B(n20261), .Z(n20271) );
  XNOR U24922 ( .A(y[1110]), .B(x[1110]), .Z(n20261) );
  XNOR U24923 ( .A(n20262), .B(n20263), .Z(n20260) );
  XNOR U24924 ( .A(y[1111]), .B(x[1111]), .Z(n20263) );
  XNOR U24925 ( .A(y[1112]), .B(x[1112]), .Z(n20262) );
  NAND U24926 ( .A(n20327), .B(n20328), .Z(N28485) );
  NANDN U24927 ( .A(n20329), .B(n20330), .Z(n20328) );
  OR U24928 ( .A(n20331), .B(n20332), .Z(n20330) );
  NAND U24929 ( .A(n20331), .B(n20332), .Z(n20327) );
  XOR U24930 ( .A(n20331), .B(n20333), .Z(N28484) );
  XNOR U24931 ( .A(n20329), .B(n20332), .Z(n20333) );
  AND U24932 ( .A(n20334), .B(n20335), .Z(n20332) );
  NANDN U24933 ( .A(n20336), .B(n20337), .Z(n20335) );
  NANDN U24934 ( .A(n20338), .B(n20339), .Z(n20337) );
  NANDN U24935 ( .A(n20339), .B(n20338), .Z(n20334) );
  NAND U24936 ( .A(n20340), .B(n20341), .Z(n20329) );
  NANDN U24937 ( .A(n20342), .B(n20343), .Z(n20341) );
  OR U24938 ( .A(n20344), .B(n20345), .Z(n20343) );
  NAND U24939 ( .A(n20345), .B(n20344), .Z(n20340) );
  AND U24940 ( .A(n20346), .B(n20347), .Z(n20331) );
  NANDN U24941 ( .A(n20348), .B(n20349), .Z(n20347) );
  NANDN U24942 ( .A(n20350), .B(n20351), .Z(n20349) );
  NANDN U24943 ( .A(n20351), .B(n20350), .Z(n20346) );
  XOR U24944 ( .A(n20345), .B(n20352), .Z(N28483) );
  XOR U24945 ( .A(n20342), .B(n20344), .Z(n20352) );
  XNOR U24946 ( .A(n20338), .B(n20353), .Z(n20344) );
  XNOR U24947 ( .A(n20336), .B(n20339), .Z(n20353) );
  NAND U24948 ( .A(n20354), .B(n20355), .Z(n20339) );
  NAND U24949 ( .A(n20356), .B(n20357), .Z(n20355) );
  OR U24950 ( .A(n20358), .B(n20359), .Z(n20356) );
  NANDN U24951 ( .A(n20360), .B(n20358), .Z(n20354) );
  IV U24952 ( .A(n20359), .Z(n20360) );
  NAND U24953 ( .A(n20361), .B(n20362), .Z(n20336) );
  NAND U24954 ( .A(n20363), .B(n20364), .Z(n20362) );
  NANDN U24955 ( .A(n20365), .B(n20366), .Z(n20363) );
  NANDN U24956 ( .A(n20366), .B(n20365), .Z(n20361) );
  AND U24957 ( .A(n20367), .B(n20368), .Z(n20338) );
  NAND U24958 ( .A(n20369), .B(n20370), .Z(n20368) );
  OR U24959 ( .A(n20371), .B(n20372), .Z(n20369) );
  NANDN U24960 ( .A(n20373), .B(n20371), .Z(n20367) );
  NAND U24961 ( .A(n20374), .B(n20375), .Z(n20342) );
  NANDN U24962 ( .A(n20376), .B(n20377), .Z(n20375) );
  OR U24963 ( .A(n20378), .B(n20379), .Z(n20377) );
  NANDN U24964 ( .A(n20380), .B(n20378), .Z(n20374) );
  IV U24965 ( .A(n20379), .Z(n20380) );
  XNOR U24966 ( .A(n20350), .B(n20381), .Z(n20345) );
  XNOR U24967 ( .A(n20348), .B(n20351), .Z(n20381) );
  NAND U24968 ( .A(n20382), .B(n20383), .Z(n20351) );
  NAND U24969 ( .A(n20384), .B(n20385), .Z(n20383) );
  OR U24970 ( .A(n20386), .B(n20387), .Z(n20384) );
  NANDN U24971 ( .A(n20388), .B(n20386), .Z(n20382) );
  IV U24972 ( .A(n20387), .Z(n20388) );
  NAND U24973 ( .A(n20389), .B(n20390), .Z(n20348) );
  NAND U24974 ( .A(n20391), .B(n20392), .Z(n20390) );
  NANDN U24975 ( .A(n20393), .B(n20394), .Z(n20391) );
  NANDN U24976 ( .A(n20394), .B(n20393), .Z(n20389) );
  AND U24977 ( .A(n20395), .B(n20396), .Z(n20350) );
  NAND U24978 ( .A(n20397), .B(n20398), .Z(n20396) );
  OR U24979 ( .A(n20399), .B(n20400), .Z(n20397) );
  NANDN U24980 ( .A(n20401), .B(n20399), .Z(n20395) );
  XNOR U24981 ( .A(n20376), .B(n20402), .Z(N28482) );
  XOR U24982 ( .A(n20378), .B(n20379), .Z(n20402) );
  XNOR U24983 ( .A(n20392), .B(n20403), .Z(n20379) );
  XOR U24984 ( .A(n20393), .B(n20394), .Z(n20403) );
  XOR U24985 ( .A(n20399), .B(n20404), .Z(n20394) );
  XOR U24986 ( .A(n20398), .B(n20401), .Z(n20404) );
  IV U24987 ( .A(n20400), .Z(n20401) );
  NAND U24988 ( .A(n20405), .B(n20406), .Z(n20400) );
  OR U24989 ( .A(n20407), .B(n20408), .Z(n20406) );
  OR U24990 ( .A(n20409), .B(n20410), .Z(n20405) );
  NAND U24991 ( .A(n20411), .B(n20412), .Z(n20398) );
  OR U24992 ( .A(n20413), .B(n20414), .Z(n20412) );
  OR U24993 ( .A(n20415), .B(n20416), .Z(n20411) );
  NOR U24994 ( .A(n20417), .B(n20418), .Z(n20399) );
  ANDN U24995 ( .B(n20419), .A(n20420), .Z(n20393) );
  XNOR U24996 ( .A(n20386), .B(n20421), .Z(n20392) );
  XNOR U24997 ( .A(n20385), .B(n20387), .Z(n20421) );
  NAND U24998 ( .A(n20422), .B(n20423), .Z(n20387) );
  OR U24999 ( .A(n20424), .B(n20425), .Z(n20423) );
  OR U25000 ( .A(n20426), .B(n20427), .Z(n20422) );
  NAND U25001 ( .A(n20428), .B(n20429), .Z(n20385) );
  OR U25002 ( .A(n20430), .B(n20431), .Z(n20429) );
  OR U25003 ( .A(n20432), .B(n20433), .Z(n20428) );
  ANDN U25004 ( .B(n20434), .A(n20435), .Z(n20386) );
  IV U25005 ( .A(n20436), .Z(n20434) );
  ANDN U25006 ( .B(n20437), .A(n20438), .Z(n20378) );
  XOR U25007 ( .A(n20364), .B(n20439), .Z(n20376) );
  XOR U25008 ( .A(n20365), .B(n20366), .Z(n20439) );
  XOR U25009 ( .A(n20371), .B(n20440), .Z(n20366) );
  XOR U25010 ( .A(n20370), .B(n20373), .Z(n20440) );
  IV U25011 ( .A(n20372), .Z(n20373) );
  NAND U25012 ( .A(n20441), .B(n20442), .Z(n20372) );
  OR U25013 ( .A(n20443), .B(n20444), .Z(n20442) );
  OR U25014 ( .A(n20445), .B(n20446), .Z(n20441) );
  NAND U25015 ( .A(n20447), .B(n20448), .Z(n20370) );
  OR U25016 ( .A(n20449), .B(n20450), .Z(n20448) );
  OR U25017 ( .A(n20451), .B(n20452), .Z(n20447) );
  NOR U25018 ( .A(n20453), .B(n20454), .Z(n20371) );
  ANDN U25019 ( .B(n20455), .A(n20456), .Z(n20365) );
  IV U25020 ( .A(n20457), .Z(n20455) );
  XNOR U25021 ( .A(n20358), .B(n20458), .Z(n20364) );
  XNOR U25022 ( .A(n20357), .B(n20359), .Z(n20458) );
  NAND U25023 ( .A(n20459), .B(n20460), .Z(n20359) );
  OR U25024 ( .A(n20461), .B(n20462), .Z(n20460) );
  OR U25025 ( .A(n20463), .B(n20464), .Z(n20459) );
  NAND U25026 ( .A(n20465), .B(n20466), .Z(n20357) );
  OR U25027 ( .A(n20467), .B(n20468), .Z(n20466) );
  OR U25028 ( .A(n20469), .B(n20470), .Z(n20465) );
  ANDN U25029 ( .B(n20471), .A(n20472), .Z(n20358) );
  IV U25030 ( .A(n20473), .Z(n20471) );
  XNOR U25031 ( .A(n20438), .B(n20437), .Z(N28481) );
  XOR U25032 ( .A(n20457), .B(n20456), .Z(n20437) );
  XNOR U25033 ( .A(n20472), .B(n20473), .Z(n20456) );
  XNOR U25034 ( .A(n20467), .B(n20468), .Z(n20473) );
  XNOR U25035 ( .A(n20469), .B(n20470), .Z(n20468) );
  XNOR U25036 ( .A(y[1108]), .B(x[1108]), .Z(n20470) );
  XNOR U25037 ( .A(y[1109]), .B(x[1109]), .Z(n20469) );
  XNOR U25038 ( .A(y[1107]), .B(x[1107]), .Z(n20467) );
  XNOR U25039 ( .A(n20461), .B(n20462), .Z(n20472) );
  XNOR U25040 ( .A(y[1104]), .B(x[1104]), .Z(n20462) );
  XNOR U25041 ( .A(n20463), .B(n20464), .Z(n20461) );
  XNOR U25042 ( .A(y[1105]), .B(x[1105]), .Z(n20464) );
  XNOR U25043 ( .A(y[1106]), .B(x[1106]), .Z(n20463) );
  XNOR U25044 ( .A(n20454), .B(n20453), .Z(n20457) );
  XNOR U25045 ( .A(n20449), .B(n20450), .Z(n20453) );
  XNOR U25046 ( .A(y[1101]), .B(x[1101]), .Z(n20450) );
  XNOR U25047 ( .A(n20451), .B(n20452), .Z(n20449) );
  XNOR U25048 ( .A(y[1102]), .B(x[1102]), .Z(n20452) );
  XNOR U25049 ( .A(y[1103]), .B(x[1103]), .Z(n20451) );
  XNOR U25050 ( .A(n20443), .B(n20444), .Z(n20454) );
  XNOR U25051 ( .A(y[1098]), .B(x[1098]), .Z(n20444) );
  XNOR U25052 ( .A(n20445), .B(n20446), .Z(n20443) );
  XNOR U25053 ( .A(y[1099]), .B(x[1099]), .Z(n20446) );
  XNOR U25054 ( .A(y[1100]), .B(x[1100]), .Z(n20445) );
  XOR U25055 ( .A(n20419), .B(n20420), .Z(n20438) );
  XNOR U25056 ( .A(n20435), .B(n20436), .Z(n20420) );
  XNOR U25057 ( .A(n20430), .B(n20431), .Z(n20436) );
  XNOR U25058 ( .A(n20432), .B(n20433), .Z(n20431) );
  XNOR U25059 ( .A(y[1096]), .B(x[1096]), .Z(n20433) );
  XNOR U25060 ( .A(y[1097]), .B(x[1097]), .Z(n20432) );
  XNOR U25061 ( .A(y[1095]), .B(x[1095]), .Z(n20430) );
  XNOR U25062 ( .A(n20424), .B(n20425), .Z(n20435) );
  XNOR U25063 ( .A(y[1092]), .B(x[1092]), .Z(n20425) );
  XNOR U25064 ( .A(n20426), .B(n20427), .Z(n20424) );
  XNOR U25065 ( .A(y[1093]), .B(x[1093]), .Z(n20427) );
  XNOR U25066 ( .A(y[1094]), .B(x[1094]), .Z(n20426) );
  XOR U25067 ( .A(n20418), .B(n20417), .Z(n20419) );
  XNOR U25068 ( .A(n20413), .B(n20414), .Z(n20417) );
  XNOR U25069 ( .A(y[1089]), .B(x[1089]), .Z(n20414) );
  XNOR U25070 ( .A(n20415), .B(n20416), .Z(n20413) );
  XNOR U25071 ( .A(y[1090]), .B(x[1090]), .Z(n20416) );
  XNOR U25072 ( .A(y[1091]), .B(x[1091]), .Z(n20415) );
  XNOR U25073 ( .A(n20407), .B(n20408), .Z(n20418) );
  XNOR U25074 ( .A(y[1086]), .B(x[1086]), .Z(n20408) );
  XNOR U25075 ( .A(n20409), .B(n20410), .Z(n20407) );
  XNOR U25076 ( .A(y[1087]), .B(x[1087]), .Z(n20410) );
  XNOR U25077 ( .A(y[1088]), .B(x[1088]), .Z(n20409) );
  NAND U25078 ( .A(n20474), .B(n20475), .Z(N28473) );
  NANDN U25079 ( .A(n20476), .B(n20477), .Z(n20475) );
  OR U25080 ( .A(n20478), .B(n20479), .Z(n20477) );
  NAND U25081 ( .A(n20478), .B(n20479), .Z(n20474) );
  XOR U25082 ( .A(n20478), .B(n20480), .Z(N28472) );
  XNOR U25083 ( .A(n20476), .B(n20479), .Z(n20480) );
  AND U25084 ( .A(n20481), .B(n20482), .Z(n20479) );
  NANDN U25085 ( .A(n20483), .B(n20484), .Z(n20482) );
  NANDN U25086 ( .A(n20485), .B(n20486), .Z(n20484) );
  NANDN U25087 ( .A(n20486), .B(n20485), .Z(n20481) );
  NAND U25088 ( .A(n20487), .B(n20488), .Z(n20476) );
  NANDN U25089 ( .A(n20489), .B(n20490), .Z(n20488) );
  OR U25090 ( .A(n20491), .B(n20492), .Z(n20490) );
  NAND U25091 ( .A(n20492), .B(n20491), .Z(n20487) );
  AND U25092 ( .A(n20493), .B(n20494), .Z(n20478) );
  NANDN U25093 ( .A(n20495), .B(n20496), .Z(n20494) );
  NANDN U25094 ( .A(n20497), .B(n20498), .Z(n20496) );
  NANDN U25095 ( .A(n20498), .B(n20497), .Z(n20493) );
  XOR U25096 ( .A(n20492), .B(n20499), .Z(N28471) );
  XOR U25097 ( .A(n20489), .B(n20491), .Z(n20499) );
  XNOR U25098 ( .A(n20485), .B(n20500), .Z(n20491) );
  XNOR U25099 ( .A(n20483), .B(n20486), .Z(n20500) );
  NAND U25100 ( .A(n20501), .B(n20502), .Z(n20486) );
  NAND U25101 ( .A(n20503), .B(n20504), .Z(n20502) );
  OR U25102 ( .A(n20505), .B(n20506), .Z(n20503) );
  NANDN U25103 ( .A(n20507), .B(n20505), .Z(n20501) );
  IV U25104 ( .A(n20506), .Z(n20507) );
  NAND U25105 ( .A(n20508), .B(n20509), .Z(n20483) );
  NAND U25106 ( .A(n20510), .B(n20511), .Z(n20509) );
  NANDN U25107 ( .A(n20512), .B(n20513), .Z(n20510) );
  NANDN U25108 ( .A(n20513), .B(n20512), .Z(n20508) );
  AND U25109 ( .A(n20514), .B(n20515), .Z(n20485) );
  NAND U25110 ( .A(n20516), .B(n20517), .Z(n20515) );
  OR U25111 ( .A(n20518), .B(n20519), .Z(n20516) );
  NANDN U25112 ( .A(n20520), .B(n20518), .Z(n20514) );
  NAND U25113 ( .A(n20521), .B(n20522), .Z(n20489) );
  NANDN U25114 ( .A(n20523), .B(n20524), .Z(n20522) );
  OR U25115 ( .A(n20525), .B(n20526), .Z(n20524) );
  NANDN U25116 ( .A(n20527), .B(n20525), .Z(n20521) );
  IV U25117 ( .A(n20526), .Z(n20527) );
  XNOR U25118 ( .A(n20497), .B(n20528), .Z(n20492) );
  XNOR U25119 ( .A(n20495), .B(n20498), .Z(n20528) );
  NAND U25120 ( .A(n20529), .B(n20530), .Z(n20498) );
  NAND U25121 ( .A(n20531), .B(n20532), .Z(n20530) );
  OR U25122 ( .A(n20533), .B(n20534), .Z(n20531) );
  NANDN U25123 ( .A(n20535), .B(n20533), .Z(n20529) );
  IV U25124 ( .A(n20534), .Z(n20535) );
  NAND U25125 ( .A(n20536), .B(n20537), .Z(n20495) );
  NAND U25126 ( .A(n20538), .B(n20539), .Z(n20537) );
  NANDN U25127 ( .A(n20540), .B(n20541), .Z(n20538) );
  NANDN U25128 ( .A(n20541), .B(n20540), .Z(n20536) );
  AND U25129 ( .A(n20542), .B(n20543), .Z(n20497) );
  NAND U25130 ( .A(n20544), .B(n20545), .Z(n20543) );
  OR U25131 ( .A(n20546), .B(n20547), .Z(n20544) );
  NANDN U25132 ( .A(n20548), .B(n20546), .Z(n20542) );
  XNOR U25133 ( .A(n20523), .B(n20549), .Z(N28470) );
  XOR U25134 ( .A(n20525), .B(n20526), .Z(n20549) );
  XNOR U25135 ( .A(n20539), .B(n20550), .Z(n20526) );
  XOR U25136 ( .A(n20540), .B(n20541), .Z(n20550) );
  XOR U25137 ( .A(n20546), .B(n20551), .Z(n20541) );
  XOR U25138 ( .A(n20545), .B(n20548), .Z(n20551) );
  IV U25139 ( .A(n20547), .Z(n20548) );
  NAND U25140 ( .A(n20552), .B(n20553), .Z(n20547) );
  OR U25141 ( .A(n20554), .B(n20555), .Z(n20553) );
  OR U25142 ( .A(n20556), .B(n20557), .Z(n20552) );
  NAND U25143 ( .A(n20558), .B(n20559), .Z(n20545) );
  OR U25144 ( .A(n20560), .B(n20561), .Z(n20559) );
  OR U25145 ( .A(n20562), .B(n20563), .Z(n20558) );
  NOR U25146 ( .A(n20564), .B(n20565), .Z(n20546) );
  ANDN U25147 ( .B(n20566), .A(n20567), .Z(n20540) );
  XNOR U25148 ( .A(n20533), .B(n20568), .Z(n20539) );
  XNOR U25149 ( .A(n20532), .B(n20534), .Z(n20568) );
  NAND U25150 ( .A(n20569), .B(n20570), .Z(n20534) );
  OR U25151 ( .A(n20571), .B(n20572), .Z(n20570) );
  OR U25152 ( .A(n20573), .B(n20574), .Z(n20569) );
  NAND U25153 ( .A(n20575), .B(n20576), .Z(n20532) );
  OR U25154 ( .A(n20577), .B(n20578), .Z(n20576) );
  OR U25155 ( .A(n20579), .B(n20580), .Z(n20575) );
  ANDN U25156 ( .B(n20581), .A(n20582), .Z(n20533) );
  IV U25157 ( .A(n20583), .Z(n20581) );
  ANDN U25158 ( .B(n20584), .A(n20585), .Z(n20525) );
  XOR U25159 ( .A(n20511), .B(n20586), .Z(n20523) );
  XOR U25160 ( .A(n20512), .B(n20513), .Z(n20586) );
  XOR U25161 ( .A(n20518), .B(n20587), .Z(n20513) );
  XOR U25162 ( .A(n20517), .B(n20520), .Z(n20587) );
  IV U25163 ( .A(n20519), .Z(n20520) );
  NAND U25164 ( .A(n20588), .B(n20589), .Z(n20519) );
  OR U25165 ( .A(n20590), .B(n20591), .Z(n20589) );
  OR U25166 ( .A(n20592), .B(n20593), .Z(n20588) );
  NAND U25167 ( .A(n20594), .B(n20595), .Z(n20517) );
  OR U25168 ( .A(n20596), .B(n20597), .Z(n20595) );
  OR U25169 ( .A(n20598), .B(n20599), .Z(n20594) );
  NOR U25170 ( .A(n20600), .B(n20601), .Z(n20518) );
  ANDN U25171 ( .B(n20602), .A(n20603), .Z(n20512) );
  IV U25172 ( .A(n20604), .Z(n20602) );
  XNOR U25173 ( .A(n20505), .B(n20605), .Z(n20511) );
  XNOR U25174 ( .A(n20504), .B(n20506), .Z(n20605) );
  NAND U25175 ( .A(n20606), .B(n20607), .Z(n20506) );
  OR U25176 ( .A(n20608), .B(n20609), .Z(n20607) );
  OR U25177 ( .A(n20610), .B(n20611), .Z(n20606) );
  NAND U25178 ( .A(n20612), .B(n20613), .Z(n20504) );
  OR U25179 ( .A(n20614), .B(n20615), .Z(n20613) );
  OR U25180 ( .A(n20616), .B(n20617), .Z(n20612) );
  ANDN U25181 ( .B(n20618), .A(n20619), .Z(n20505) );
  IV U25182 ( .A(n20620), .Z(n20618) );
  XNOR U25183 ( .A(n20585), .B(n20584), .Z(N28469) );
  XOR U25184 ( .A(n20604), .B(n20603), .Z(n20584) );
  XNOR U25185 ( .A(n20619), .B(n20620), .Z(n20603) );
  XNOR U25186 ( .A(n20614), .B(n20615), .Z(n20620) );
  XNOR U25187 ( .A(n20616), .B(n20617), .Z(n20615) );
  XNOR U25188 ( .A(y[1084]), .B(x[1084]), .Z(n20617) );
  XNOR U25189 ( .A(y[1085]), .B(x[1085]), .Z(n20616) );
  XNOR U25190 ( .A(y[1083]), .B(x[1083]), .Z(n20614) );
  XNOR U25191 ( .A(n20608), .B(n20609), .Z(n20619) );
  XNOR U25192 ( .A(y[1080]), .B(x[1080]), .Z(n20609) );
  XNOR U25193 ( .A(n20610), .B(n20611), .Z(n20608) );
  XNOR U25194 ( .A(y[1081]), .B(x[1081]), .Z(n20611) );
  XNOR U25195 ( .A(y[1082]), .B(x[1082]), .Z(n20610) );
  XNOR U25196 ( .A(n20601), .B(n20600), .Z(n20604) );
  XNOR U25197 ( .A(n20596), .B(n20597), .Z(n20600) );
  XNOR U25198 ( .A(y[1077]), .B(x[1077]), .Z(n20597) );
  XNOR U25199 ( .A(n20598), .B(n20599), .Z(n20596) );
  XNOR U25200 ( .A(y[1078]), .B(x[1078]), .Z(n20599) );
  XNOR U25201 ( .A(y[1079]), .B(x[1079]), .Z(n20598) );
  XNOR U25202 ( .A(n20590), .B(n20591), .Z(n20601) );
  XNOR U25203 ( .A(y[1074]), .B(x[1074]), .Z(n20591) );
  XNOR U25204 ( .A(n20592), .B(n20593), .Z(n20590) );
  XNOR U25205 ( .A(y[1075]), .B(x[1075]), .Z(n20593) );
  XNOR U25206 ( .A(y[1076]), .B(x[1076]), .Z(n20592) );
  XOR U25207 ( .A(n20566), .B(n20567), .Z(n20585) );
  XNOR U25208 ( .A(n20582), .B(n20583), .Z(n20567) );
  XNOR U25209 ( .A(n20577), .B(n20578), .Z(n20583) );
  XNOR U25210 ( .A(n20579), .B(n20580), .Z(n20578) );
  XNOR U25211 ( .A(y[1072]), .B(x[1072]), .Z(n20580) );
  XNOR U25212 ( .A(y[1073]), .B(x[1073]), .Z(n20579) );
  XNOR U25213 ( .A(y[1071]), .B(x[1071]), .Z(n20577) );
  XNOR U25214 ( .A(n20571), .B(n20572), .Z(n20582) );
  XNOR U25215 ( .A(y[1068]), .B(x[1068]), .Z(n20572) );
  XNOR U25216 ( .A(n20573), .B(n20574), .Z(n20571) );
  XNOR U25217 ( .A(y[1069]), .B(x[1069]), .Z(n20574) );
  XNOR U25218 ( .A(y[1070]), .B(x[1070]), .Z(n20573) );
  XOR U25219 ( .A(n20565), .B(n20564), .Z(n20566) );
  XNOR U25220 ( .A(n20560), .B(n20561), .Z(n20564) );
  XNOR U25221 ( .A(y[1065]), .B(x[1065]), .Z(n20561) );
  XNOR U25222 ( .A(n20562), .B(n20563), .Z(n20560) );
  XNOR U25223 ( .A(y[1066]), .B(x[1066]), .Z(n20563) );
  XNOR U25224 ( .A(y[1067]), .B(x[1067]), .Z(n20562) );
  XNOR U25225 ( .A(n20554), .B(n20555), .Z(n20565) );
  XNOR U25226 ( .A(y[1062]), .B(x[1062]), .Z(n20555) );
  XNOR U25227 ( .A(n20556), .B(n20557), .Z(n20554) );
  XNOR U25228 ( .A(y[1063]), .B(x[1063]), .Z(n20557) );
  XNOR U25229 ( .A(y[1064]), .B(x[1064]), .Z(n20556) );
  NAND U25230 ( .A(n20621), .B(n20622), .Z(N28461) );
  NANDN U25231 ( .A(n20623), .B(n20624), .Z(n20622) );
  OR U25232 ( .A(n20625), .B(n20626), .Z(n20624) );
  NAND U25233 ( .A(n20625), .B(n20626), .Z(n20621) );
  XOR U25234 ( .A(n20625), .B(n20627), .Z(N28460) );
  XNOR U25235 ( .A(n20623), .B(n20626), .Z(n20627) );
  AND U25236 ( .A(n20628), .B(n20629), .Z(n20626) );
  NANDN U25237 ( .A(n20630), .B(n20631), .Z(n20629) );
  NANDN U25238 ( .A(n20632), .B(n20633), .Z(n20631) );
  NANDN U25239 ( .A(n20633), .B(n20632), .Z(n20628) );
  NAND U25240 ( .A(n20634), .B(n20635), .Z(n20623) );
  NANDN U25241 ( .A(n20636), .B(n20637), .Z(n20635) );
  OR U25242 ( .A(n20638), .B(n20639), .Z(n20637) );
  NAND U25243 ( .A(n20639), .B(n20638), .Z(n20634) );
  AND U25244 ( .A(n20640), .B(n20641), .Z(n20625) );
  NANDN U25245 ( .A(n20642), .B(n20643), .Z(n20641) );
  NANDN U25246 ( .A(n20644), .B(n20645), .Z(n20643) );
  NANDN U25247 ( .A(n20645), .B(n20644), .Z(n20640) );
  XOR U25248 ( .A(n20639), .B(n20646), .Z(N28459) );
  XOR U25249 ( .A(n20636), .B(n20638), .Z(n20646) );
  XNOR U25250 ( .A(n20632), .B(n20647), .Z(n20638) );
  XNOR U25251 ( .A(n20630), .B(n20633), .Z(n20647) );
  NAND U25252 ( .A(n20648), .B(n20649), .Z(n20633) );
  NAND U25253 ( .A(n20650), .B(n20651), .Z(n20649) );
  OR U25254 ( .A(n20652), .B(n20653), .Z(n20650) );
  NANDN U25255 ( .A(n20654), .B(n20652), .Z(n20648) );
  IV U25256 ( .A(n20653), .Z(n20654) );
  NAND U25257 ( .A(n20655), .B(n20656), .Z(n20630) );
  NAND U25258 ( .A(n20657), .B(n20658), .Z(n20656) );
  NANDN U25259 ( .A(n20659), .B(n20660), .Z(n20657) );
  NANDN U25260 ( .A(n20660), .B(n20659), .Z(n20655) );
  AND U25261 ( .A(n20661), .B(n20662), .Z(n20632) );
  NAND U25262 ( .A(n20663), .B(n20664), .Z(n20662) );
  OR U25263 ( .A(n20665), .B(n20666), .Z(n20663) );
  NANDN U25264 ( .A(n20667), .B(n20665), .Z(n20661) );
  NAND U25265 ( .A(n20668), .B(n20669), .Z(n20636) );
  NANDN U25266 ( .A(n20670), .B(n20671), .Z(n20669) );
  OR U25267 ( .A(n20672), .B(n20673), .Z(n20671) );
  NANDN U25268 ( .A(n20674), .B(n20672), .Z(n20668) );
  IV U25269 ( .A(n20673), .Z(n20674) );
  XNOR U25270 ( .A(n20644), .B(n20675), .Z(n20639) );
  XNOR U25271 ( .A(n20642), .B(n20645), .Z(n20675) );
  NAND U25272 ( .A(n20676), .B(n20677), .Z(n20645) );
  NAND U25273 ( .A(n20678), .B(n20679), .Z(n20677) );
  OR U25274 ( .A(n20680), .B(n20681), .Z(n20678) );
  NANDN U25275 ( .A(n20682), .B(n20680), .Z(n20676) );
  IV U25276 ( .A(n20681), .Z(n20682) );
  NAND U25277 ( .A(n20683), .B(n20684), .Z(n20642) );
  NAND U25278 ( .A(n20685), .B(n20686), .Z(n20684) );
  NANDN U25279 ( .A(n20687), .B(n20688), .Z(n20685) );
  NANDN U25280 ( .A(n20688), .B(n20687), .Z(n20683) );
  AND U25281 ( .A(n20689), .B(n20690), .Z(n20644) );
  NAND U25282 ( .A(n20691), .B(n20692), .Z(n20690) );
  OR U25283 ( .A(n20693), .B(n20694), .Z(n20691) );
  NANDN U25284 ( .A(n20695), .B(n20693), .Z(n20689) );
  XNOR U25285 ( .A(n20670), .B(n20696), .Z(N28458) );
  XOR U25286 ( .A(n20672), .B(n20673), .Z(n20696) );
  XNOR U25287 ( .A(n20686), .B(n20697), .Z(n20673) );
  XOR U25288 ( .A(n20687), .B(n20688), .Z(n20697) );
  XOR U25289 ( .A(n20693), .B(n20698), .Z(n20688) );
  XOR U25290 ( .A(n20692), .B(n20695), .Z(n20698) );
  IV U25291 ( .A(n20694), .Z(n20695) );
  NAND U25292 ( .A(n20699), .B(n20700), .Z(n20694) );
  OR U25293 ( .A(n20701), .B(n20702), .Z(n20700) );
  OR U25294 ( .A(n20703), .B(n20704), .Z(n20699) );
  NAND U25295 ( .A(n20705), .B(n20706), .Z(n20692) );
  OR U25296 ( .A(n20707), .B(n20708), .Z(n20706) );
  OR U25297 ( .A(n20709), .B(n20710), .Z(n20705) );
  NOR U25298 ( .A(n20711), .B(n20712), .Z(n20693) );
  ANDN U25299 ( .B(n20713), .A(n20714), .Z(n20687) );
  XNOR U25300 ( .A(n20680), .B(n20715), .Z(n20686) );
  XNOR U25301 ( .A(n20679), .B(n20681), .Z(n20715) );
  NAND U25302 ( .A(n20716), .B(n20717), .Z(n20681) );
  OR U25303 ( .A(n20718), .B(n20719), .Z(n20717) );
  OR U25304 ( .A(n20720), .B(n20721), .Z(n20716) );
  NAND U25305 ( .A(n20722), .B(n20723), .Z(n20679) );
  OR U25306 ( .A(n20724), .B(n20725), .Z(n20723) );
  OR U25307 ( .A(n20726), .B(n20727), .Z(n20722) );
  ANDN U25308 ( .B(n20728), .A(n20729), .Z(n20680) );
  IV U25309 ( .A(n20730), .Z(n20728) );
  ANDN U25310 ( .B(n20731), .A(n20732), .Z(n20672) );
  XOR U25311 ( .A(n20658), .B(n20733), .Z(n20670) );
  XOR U25312 ( .A(n20659), .B(n20660), .Z(n20733) );
  XOR U25313 ( .A(n20665), .B(n20734), .Z(n20660) );
  XOR U25314 ( .A(n20664), .B(n20667), .Z(n20734) );
  IV U25315 ( .A(n20666), .Z(n20667) );
  NAND U25316 ( .A(n20735), .B(n20736), .Z(n20666) );
  OR U25317 ( .A(n20737), .B(n20738), .Z(n20736) );
  OR U25318 ( .A(n20739), .B(n20740), .Z(n20735) );
  NAND U25319 ( .A(n20741), .B(n20742), .Z(n20664) );
  OR U25320 ( .A(n20743), .B(n20744), .Z(n20742) );
  OR U25321 ( .A(n20745), .B(n20746), .Z(n20741) );
  NOR U25322 ( .A(n20747), .B(n20748), .Z(n20665) );
  ANDN U25323 ( .B(n20749), .A(n20750), .Z(n20659) );
  IV U25324 ( .A(n20751), .Z(n20749) );
  XNOR U25325 ( .A(n20652), .B(n20752), .Z(n20658) );
  XNOR U25326 ( .A(n20651), .B(n20653), .Z(n20752) );
  NAND U25327 ( .A(n20753), .B(n20754), .Z(n20653) );
  OR U25328 ( .A(n20755), .B(n20756), .Z(n20754) );
  OR U25329 ( .A(n20757), .B(n20758), .Z(n20753) );
  NAND U25330 ( .A(n20759), .B(n20760), .Z(n20651) );
  OR U25331 ( .A(n20761), .B(n20762), .Z(n20760) );
  OR U25332 ( .A(n20763), .B(n20764), .Z(n20759) );
  ANDN U25333 ( .B(n20765), .A(n20766), .Z(n20652) );
  IV U25334 ( .A(n20767), .Z(n20765) );
  XNOR U25335 ( .A(n20732), .B(n20731), .Z(N28457) );
  XOR U25336 ( .A(n20751), .B(n20750), .Z(n20731) );
  XNOR U25337 ( .A(n20766), .B(n20767), .Z(n20750) );
  XNOR U25338 ( .A(n20761), .B(n20762), .Z(n20767) );
  XNOR U25339 ( .A(n20763), .B(n20764), .Z(n20762) );
  XNOR U25340 ( .A(y[1060]), .B(x[1060]), .Z(n20764) );
  XNOR U25341 ( .A(y[1061]), .B(x[1061]), .Z(n20763) );
  XNOR U25342 ( .A(y[1059]), .B(x[1059]), .Z(n20761) );
  XNOR U25343 ( .A(n20755), .B(n20756), .Z(n20766) );
  XNOR U25344 ( .A(y[1056]), .B(x[1056]), .Z(n20756) );
  XNOR U25345 ( .A(n20757), .B(n20758), .Z(n20755) );
  XNOR U25346 ( .A(y[1057]), .B(x[1057]), .Z(n20758) );
  XNOR U25347 ( .A(y[1058]), .B(x[1058]), .Z(n20757) );
  XNOR U25348 ( .A(n20748), .B(n20747), .Z(n20751) );
  XNOR U25349 ( .A(n20743), .B(n20744), .Z(n20747) );
  XNOR U25350 ( .A(y[1053]), .B(x[1053]), .Z(n20744) );
  XNOR U25351 ( .A(n20745), .B(n20746), .Z(n20743) );
  XNOR U25352 ( .A(y[1054]), .B(x[1054]), .Z(n20746) );
  XNOR U25353 ( .A(y[1055]), .B(x[1055]), .Z(n20745) );
  XNOR U25354 ( .A(n20737), .B(n20738), .Z(n20748) );
  XNOR U25355 ( .A(y[1050]), .B(x[1050]), .Z(n20738) );
  XNOR U25356 ( .A(n20739), .B(n20740), .Z(n20737) );
  XNOR U25357 ( .A(y[1051]), .B(x[1051]), .Z(n20740) );
  XNOR U25358 ( .A(y[1052]), .B(x[1052]), .Z(n20739) );
  XOR U25359 ( .A(n20713), .B(n20714), .Z(n20732) );
  XNOR U25360 ( .A(n20729), .B(n20730), .Z(n20714) );
  XNOR U25361 ( .A(n20724), .B(n20725), .Z(n20730) );
  XNOR U25362 ( .A(n20726), .B(n20727), .Z(n20725) );
  XNOR U25363 ( .A(y[1048]), .B(x[1048]), .Z(n20727) );
  XNOR U25364 ( .A(y[1049]), .B(x[1049]), .Z(n20726) );
  XNOR U25365 ( .A(y[1047]), .B(x[1047]), .Z(n20724) );
  XNOR U25366 ( .A(n20718), .B(n20719), .Z(n20729) );
  XNOR U25367 ( .A(y[1044]), .B(x[1044]), .Z(n20719) );
  XNOR U25368 ( .A(n20720), .B(n20721), .Z(n20718) );
  XNOR U25369 ( .A(y[1045]), .B(x[1045]), .Z(n20721) );
  XNOR U25370 ( .A(y[1046]), .B(x[1046]), .Z(n20720) );
  XOR U25371 ( .A(n20712), .B(n20711), .Z(n20713) );
  XNOR U25372 ( .A(n20707), .B(n20708), .Z(n20711) );
  XNOR U25373 ( .A(y[1041]), .B(x[1041]), .Z(n20708) );
  XNOR U25374 ( .A(n20709), .B(n20710), .Z(n20707) );
  XNOR U25375 ( .A(y[1042]), .B(x[1042]), .Z(n20710) );
  XNOR U25376 ( .A(y[1043]), .B(x[1043]), .Z(n20709) );
  XNOR U25377 ( .A(n20701), .B(n20702), .Z(n20712) );
  XNOR U25378 ( .A(y[1038]), .B(x[1038]), .Z(n20702) );
  XNOR U25379 ( .A(n20703), .B(n20704), .Z(n20701) );
  XNOR U25380 ( .A(y[1039]), .B(x[1039]), .Z(n20704) );
  XNOR U25381 ( .A(y[1040]), .B(x[1040]), .Z(n20703) );
  NAND U25382 ( .A(n20768), .B(n20769), .Z(N28449) );
  NANDN U25383 ( .A(n20770), .B(n20771), .Z(n20769) );
  OR U25384 ( .A(n20772), .B(n20773), .Z(n20771) );
  NAND U25385 ( .A(n20772), .B(n20773), .Z(n20768) );
  XOR U25386 ( .A(n20772), .B(n20774), .Z(N28448) );
  XNOR U25387 ( .A(n20770), .B(n20773), .Z(n20774) );
  AND U25388 ( .A(n20775), .B(n20776), .Z(n20773) );
  NANDN U25389 ( .A(n20777), .B(n20778), .Z(n20776) );
  NANDN U25390 ( .A(n20779), .B(n20780), .Z(n20778) );
  NANDN U25391 ( .A(n20780), .B(n20779), .Z(n20775) );
  NAND U25392 ( .A(n20781), .B(n20782), .Z(n20770) );
  NANDN U25393 ( .A(n20783), .B(n20784), .Z(n20782) );
  OR U25394 ( .A(n20785), .B(n20786), .Z(n20784) );
  NAND U25395 ( .A(n20786), .B(n20785), .Z(n20781) );
  AND U25396 ( .A(n20787), .B(n20788), .Z(n20772) );
  NANDN U25397 ( .A(n20789), .B(n20790), .Z(n20788) );
  NANDN U25398 ( .A(n20791), .B(n20792), .Z(n20790) );
  NANDN U25399 ( .A(n20792), .B(n20791), .Z(n20787) );
  XOR U25400 ( .A(n20786), .B(n20793), .Z(N28447) );
  XOR U25401 ( .A(n20783), .B(n20785), .Z(n20793) );
  XNOR U25402 ( .A(n20779), .B(n20794), .Z(n20785) );
  XNOR U25403 ( .A(n20777), .B(n20780), .Z(n20794) );
  NAND U25404 ( .A(n20795), .B(n20796), .Z(n20780) );
  NAND U25405 ( .A(n20797), .B(n20798), .Z(n20796) );
  OR U25406 ( .A(n20799), .B(n20800), .Z(n20797) );
  NANDN U25407 ( .A(n20801), .B(n20799), .Z(n20795) );
  IV U25408 ( .A(n20800), .Z(n20801) );
  NAND U25409 ( .A(n20802), .B(n20803), .Z(n20777) );
  NAND U25410 ( .A(n20804), .B(n20805), .Z(n20803) );
  NANDN U25411 ( .A(n20806), .B(n20807), .Z(n20804) );
  NANDN U25412 ( .A(n20807), .B(n20806), .Z(n20802) );
  AND U25413 ( .A(n20808), .B(n20809), .Z(n20779) );
  NAND U25414 ( .A(n20810), .B(n20811), .Z(n20809) );
  OR U25415 ( .A(n20812), .B(n20813), .Z(n20810) );
  NANDN U25416 ( .A(n20814), .B(n20812), .Z(n20808) );
  NAND U25417 ( .A(n20815), .B(n20816), .Z(n20783) );
  NANDN U25418 ( .A(n20817), .B(n20818), .Z(n20816) );
  OR U25419 ( .A(n20819), .B(n20820), .Z(n20818) );
  NANDN U25420 ( .A(n20821), .B(n20819), .Z(n20815) );
  IV U25421 ( .A(n20820), .Z(n20821) );
  XNOR U25422 ( .A(n20791), .B(n20822), .Z(n20786) );
  XNOR U25423 ( .A(n20789), .B(n20792), .Z(n20822) );
  NAND U25424 ( .A(n20823), .B(n20824), .Z(n20792) );
  NAND U25425 ( .A(n20825), .B(n20826), .Z(n20824) );
  OR U25426 ( .A(n20827), .B(n20828), .Z(n20825) );
  NANDN U25427 ( .A(n20829), .B(n20827), .Z(n20823) );
  IV U25428 ( .A(n20828), .Z(n20829) );
  NAND U25429 ( .A(n20830), .B(n20831), .Z(n20789) );
  NAND U25430 ( .A(n20832), .B(n20833), .Z(n20831) );
  NANDN U25431 ( .A(n20834), .B(n20835), .Z(n20832) );
  NANDN U25432 ( .A(n20835), .B(n20834), .Z(n20830) );
  AND U25433 ( .A(n20836), .B(n20837), .Z(n20791) );
  NAND U25434 ( .A(n20838), .B(n20839), .Z(n20837) );
  OR U25435 ( .A(n20840), .B(n20841), .Z(n20838) );
  NANDN U25436 ( .A(n20842), .B(n20840), .Z(n20836) );
  XNOR U25437 ( .A(n20817), .B(n20843), .Z(N28446) );
  XOR U25438 ( .A(n20819), .B(n20820), .Z(n20843) );
  XNOR U25439 ( .A(n20833), .B(n20844), .Z(n20820) );
  XOR U25440 ( .A(n20834), .B(n20835), .Z(n20844) );
  XOR U25441 ( .A(n20840), .B(n20845), .Z(n20835) );
  XOR U25442 ( .A(n20839), .B(n20842), .Z(n20845) );
  IV U25443 ( .A(n20841), .Z(n20842) );
  NAND U25444 ( .A(n20846), .B(n20847), .Z(n20841) );
  OR U25445 ( .A(n20848), .B(n20849), .Z(n20847) );
  OR U25446 ( .A(n20850), .B(n20851), .Z(n20846) );
  NAND U25447 ( .A(n20852), .B(n20853), .Z(n20839) );
  OR U25448 ( .A(n20854), .B(n20855), .Z(n20853) );
  OR U25449 ( .A(n20856), .B(n20857), .Z(n20852) );
  NOR U25450 ( .A(n20858), .B(n20859), .Z(n20840) );
  ANDN U25451 ( .B(n20860), .A(n20861), .Z(n20834) );
  XNOR U25452 ( .A(n20827), .B(n20862), .Z(n20833) );
  XNOR U25453 ( .A(n20826), .B(n20828), .Z(n20862) );
  NAND U25454 ( .A(n20863), .B(n20864), .Z(n20828) );
  OR U25455 ( .A(n20865), .B(n20866), .Z(n20864) );
  OR U25456 ( .A(n20867), .B(n20868), .Z(n20863) );
  NAND U25457 ( .A(n20869), .B(n20870), .Z(n20826) );
  OR U25458 ( .A(n20871), .B(n20872), .Z(n20870) );
  OR U25459 ( .A(n20873), .B(n20874), .Z(n20869) );
  ANDN U25460 ( .B(n20875), .A(n20876), .Z(n20827) );
  IV U25461 ( .A(n20877), .Z(n20875) );
  ANDN U25462 ( .B(n20878), .A(n20879), .Z(n20819) );
  XOR U25463 ( .A(n20805), .B(n20880), .Z(n20817) );
  XOR U25464 ( .A(n20806), .B(n20807), .Z(n20880) );
  XOR U25465 ( .A(n20812), .B(n20881), .Z(n20807) );
  XOR U25466 ( .A(n20811), .B(n20814), .Z(n20881) );
  IV U25467 ( .A(n20813), .Z(n20814) );
  NAND U25468 ( .A(n20882), .B(n20883), .Z(n20813) );
  OR U25469 ( .A(n20884), .B(n20885), .Z(n20883) );
  OR U25470 ( .A(n20886), .B(n20887), .Z(n20882) );
  NAND U25471 ( .A(n20888), .B(n20889), .Z(n20811) );
  OR U25472 ( .A(n20890), .B(n20891), .Z(n20889) );
  OR U25473 ( .A(n20892), .B(n20893), .Z(n20888) );
  NOR U25474 ( .A(n20894), .B(n20895), .Z(n20812) );
  ANDN U25475 ( .B(n20896), .A(n20897), .Z(n20806) );
  IV U25476 ( .A(n20898), .Z(n20896) );
  XNOR U25477 ( .A(n20799), .B(n20899), .Z(n20805) );
  XNOR U25478 ( .A(n20798), .B(n20800), .Z(n20899) );
  NAND U25479 ( .A(n20900), .B(n20901), .Z(n20800) );
  OR U25480 ( .A(n20902), .B(n20903), .Z(n20901) );
  OR U25481 ( .A(n20904), .B(n20905), .Z(n20900) );
  NAND U25482 ( .A(n20906), .B(n20907), .Z(n20798) );
  OR U25483 ( .A(n20908), .B(n20909), .Z(n20907) );
  OR U25484 ( .A(n20910), .B(n20911), .Z(n20906) );
  ANDN U25485 ( .B(n20912), .A(n20913), .Z(n20799) );
  IV U25486 ( .A(n20914), .Z(n20912) );
  XNOR U25487 ( .A(n20879), .B(n20878), .Z(N28445) );
  XOR U25488 ( .A(n20898), .B(n20897), .Z(n20878) );
  XNOR U25489 ( .A(n20913), .B(n20914), .Z(n20897) );
  XNOR U25490 ( .A(n20908), .B(n20909), .Z(n20914) );
  XNOR U25491 ( .A(n20910), .B(n20911), .Z(n20909) );
  XNOR U25492 ( .A(y[1036]), .B(x[1036]), .Z(n20911) );
  XNOR U25493 ( .A(y[1037]), .B(x[1037]), .Z(n20910) );
  XNOR U25494 ( .A(y[1035]), .B(x[1035]), .Z(n20908) );
  XNOR U25495 ( .A(n20902), .B(n20903), .Z(n20913) );
  XNOR U25496 ( .A(y[1032]), .B(x[1032]), .Z(n20903) );
  XNOR U25497 ( .A(n20904), .B(n20905), .Z(n20902) );
  XNOR U25498 ( .A(y[1033]), .B(x[1033]), .Z(n20905) );
  XNOR U25499 ( .A(y[1034]), .B(x[1034]), .Z(n20904) );
  XNOR U25500 ( .A(n20895), .B(n20894), .Z(n20898) );
  XNOR U25501 ( .A(n20890), .B(n20891), .Z(n20894) );
  XNOR U25502 ( .A(y[1029]), .B(x[1029]), .Z(n20891) );
  XNOR U25503 ( .A(n20892), .B(n20893), .Z(n20890) );
  XNOR U25504 ( .A(y[1030]), .B(x[1030]), .Z(n20893) );
  XNOR U25505 ( .A(y[1031]), .B(x[1031]), .Z(n20892) );
  XNOR U25506 ( .A(n20884), .B(n20885), .Z(n20895) );
  XNOR U25507 ( .A(y[1026]), .B(x[1026]), .Z(n20885) );
  XNOR U25508 ( .A(n20886), .B(n20887), .Z(n20884) );
  XNOR U25509 ( .A(y[1027]), .B(x[1027]), .Z(n20887) );
  XNOR U25510 ( .A(y[1028]), .B(x[1028]), .Z(n20886) );
  XOR U25511 ( .A(n20860), .B(n20861), .Z(n20879) );
  XNOR U25512 ( .A(n20876), .B(n20877), .Z(n20861) );
  XNOR U25513 ( .A(n20871), .B(n20872), .Z(n20877) );
  XNOR U25514 ( .A(n20873), .B(n20874), .Z(n20872) );
  XNOR U25515 ( .A(y[1024]), .B(x[1024]), .Z(n20874) );
  XNOR U25516 ( .A(y[1025]), .B(x[1025]), .Z(n20873) );
  XNOR U25517 ( .A(y[1023]), .B(x[1023]), .Z(n20871) );
  XNOR U25518 ( .A(n20865), .B(n20866), .Z(n20876) );
  XNOR U25519 ( .A(y[1020]), .B(x[1020]), .Z(n20866) );
  XNOR U25520 ( .A(n20867), .B(n20868), .Z(n20865) );
  XNOR U25521 ( .A(y[1021]), .B(x[1021]), .Z(n20868) );
  XNOR U25522 ( .A(y[1022]), .B(x[1022]), .Z(n20867) );
  XOR U25523 ( .A(n20859), .B(n20858), .Z(n20860) );
  XNOR U25524 ( .A(n20854), .B(n20855), .Z(n20858) );
  XNOR U25525 ( .A(y[1017]), .B(x[1017]), .Z(n20855) );
  XNOR U25526 ( .A(n20856), .B(n20857), .Z(n20854) );
  XNOR U25527 ( .A(y[1018]), .B(x[1018]), .Z(n20857) );
  XNOR U25528 ( .A(y[1019]), .B(x[1019]), .Z(n20856) );
  XNOR U25529 ( .A(n20848), .B(n20849), .Z(n20859) );
  XNOR U25530 ( .A(y[1014]), .B(x[1014]), .Z(n20849) );
  XNOR U25531 ( .A(n20850), .B(n20851), .Z(n20848) );
  XNOR U25532 ( .A(y[1015]), .B(x[1015]), .Z(n20851) );
  XNOR U25533 ( .A(y[1016]), .B(x[1016]), .Z(n20850) );
  NAND U25534 ( .A(n20915), .B(n20916), .Z(N28437) );
  NANDN U25535 ( .A(n20917), .B(n20918), .Z(n20916) );
  OR U25536 ( .A(n20919), .B(n20920), .Z(n20918) );
  NAND U25537 ( .A(n20919), .B(n20920), .Z(n20915) );
  XOR U25538 ( .A(n20919), .B(n20921), .Z(N28436) );
  XNOR U25539 ( .A(n20917), .B(n20920), .Z(n20921) );
  AND U25540 ( .A(n20922), .B(n20923), .Z(n20920) );
  NANDN U25541 ( .A(n20924), .B(n20925), .Z(n20923) );
  NANDN U25542 ( .A(n20926), .B(n20927), .Z(n20925) );
  NANDN U25543 ( .A(n20927), .B(n20926), .Z(n20922) );
  NAND U25544 ( .A(n20928), .B(n20929), .Z(n20917) );
  NANDN U25545 ( .A(n20930), .B(n20931), .Z(n20929) );
  OR U25546 ( .A(n20932), .B(n20933), .Z(n20931) );
  NAND U25547 ( .A(n20933), .B(n20932), .Z(n20928) );
  AND U25548 ( .A(n20934), .B(n20935), .Z(n20919) );
  NANDN U25549 ( .A(n20936), .B(n20937), .Z(n20935) );
  NANDN U25550 ( .A(n20938), .B(n20939), .Z(n20937) );
  NANDN U25551 ( .A(n20939), .B(n20938), .Z(n20934) );
  XOR U25552 ( .A(n20933), .B(n20940), .Z(N28435) );
  XOR U25553 ( .A(n20930), .B(n20932), .Z(n20940) );
  XNOR U25554 ( .A(n20926), .B(n20941), .Z(n20932) );
  XNOR U25555 ( .A(n20924), .B(n20927), .Z(n20941) );
  NAND U25556 ( .A(n20942), .B(n20943), .Z(n20927) );
  NAND U25557 ( .A(n20944), .B(n20945), .Z(n20943) );
  OR U25558 ( .A(n20946), .B(n20947), .Z(n20944) );
  NANDN U25559 ( .A(n20948), .B(n20946), .Z(n20942) );
  IV U25560 ( .A(n20947), .Z(n20948) );
  NAND U25561 ( .A(n20949), .B(n20950), .Z(n20924) );
  NAND U25562 ( .A(n20951), .B(n20952), .Z(n20950) );
  NANDN U25563 ( .A(n20953), .B(n20954), .Z(n20951) );
  NANDN U25564 ( .A(n20954), .B(n20953), .Z(n20949) );
  AND U25565 ( .A(n20955), .B(n20956), .Z(n20926) );
  NAND U25566 ( .A(n20957), .B(n20958), .Z(n20956) );
  OR U25567 ( .A(n20959), .B(n20960), .Z(n20957) );
  NANDN U25568 ( .A(n20961), .B(n20959), .Z(n20955) );
  NAND U25569 ( .A(n20962), .B(n20963), .Z(n20930) );
  NANDN U25570 ( .A(n20964), .B(n20965), .Z(n20963) );
  OR U25571 ( .A(n20966), .B(n20967), .Z(n20965) );
  NANDN U25572 ( .A(n20968), .B(n20966), .Z(n20962) );
  IV U25573 ( .A(n20967), .Z(n20968) );
  XNOR U25574 ( .A(n20938), .B(n20969), .Z(n20933) );
  XNOR U25575 ( .A(n20936), .B(n20939), .Z(n20969) );
  NAND U25576 ( .A(n20970), .B(n20971), .Z(n20939) );
  NAND U25577 ( .A(n20972), .B(n20973), .Z(n20971) );
  OR U25578 ( .A(n20974), .B(n20975), .Z(n20972) );
  NANDN U25579 ( .A(n20976), .B(n20974), .Z(n20970) );
  IV U25580 ( .A(n20975), .Z(n20976) );
  NAND U25581 ( .A(n20977), .B(n20978), .Z(n20936) );
  NAND U25582 ( .A(n20979), .B(n20980), .Z(n20978) );
  NANDN U25583 ( .A(n20981), .B(n20982), .Z(n20979) );
  NANDN U25584 ( .A(n20982), .B(n20981), .Z(n20977) );
  AND U25585 ( .A(n20983), .B(n20984), .Z(n20938) );
  NAND U25586 ( .A(n20985), .B(n20986), .Z(n20984) );
  OR U25587 ( .A(n20987), .B(n20988), .Z(n20985) );
  NANDN U25588 ( .A(n20989), .B(n20987), .Z(n20983) );
  XNOR U25589 ( .A(n20964), .B(n20990), .Z(N28434) );
  XOR U25590 ( .A(n20966), .B(n20967), .Z(n20990) );
  XNOR U25591 ( .A(n20980), .B(n20991), .Z(n20967) );
  XOR U25592 ( .A(n20981), .B(n20982), .Z(n20991) );
  XOR U25593 ( .A(n20987), .B(n20992), .Z(n20982) );
  XOR U25594 ( .A(n20986), .B(n20989), .Z(n20992) );
  IV U25595 ( .A(n20988), .Z(n20989) );
  NAND U25596 ( .A(n20993), .B(n20994), .Z(n20988) );
  OR U25597 ( .A(n20995), .B(n20996), .Z(n20994) );
  OR U25598 ( .A(n20997), .B(n20998), .Z(n20993) );
  NAND U25599 ( .A(n20999), .B(n21000), .Z(n20986) );
  OR U25600 ( .A(n21001), .B(n21002), .Z(n21000) );
  OR U25601 ( .A(n21003), .B(n21004), .Z(n20999) );
  NOR U25602 ( .A(n21005), .B(n21006), .Z(n20987) );
  ANDN U25603 ( .B(n21007), .A(n21008), .Z(n20981) );
  XNOR U25604 ( .A(n20974), .B(n21009), .Z(n20980) );
  XNOR U25605 ( .A(n20973), .B(n20975), .Z(n21009) );
  NAND U25606 ( .A(n21010), .B(n21011), .Z(n20975) );
  OR U25607 ( .A(n21012), .B(n21013), .Z(n21011) );
  OR U25608 ( .A(n21014), .B(n21015), .Z(n21010) );
  NAND U25609 ( .A(n21016), .B(n21017), .Z(n20973) );
  OR U25610 ( .A(n21018), .B(n21019), .Z(n21017) );
  OR U25611 ( .A(n21020), .B(n21021), .Z(n21016) );
  ANDN U25612 ( .B(n21022), .A(n21023), .Z(n20974) );
  IV U25613 ( .A(n21024), .Z(n21022) );
  ANDN U25614 ( .B(n21025), .A(n21026), .Z(n20966) );
  XOR U25615 ( .A(n20952), .B(n21027), .Z(n20964) );
  XOR U25616 ( .A(n20953), .B(n20954), .Z(n21027) );
  XOR U25617 ( .A(n20959), .B(n21028), .Z(n20954) );
  XOR U25618 ( .A(n20958), .B(n20961), .Z(n21028) );
  IV U25619 ( .A(n20960), .Z(n20961) );
  NAND U25620 ( .A(n21029), .B(n21030), .Z(n20960) );
  OR U25621 ( .A(n21031), .B(n21032), .Z(n21030) );
  OR U25622 ( .A(n21033), .B(n21034), .Z(n21029) );
  NAND U25623 ( .A(n21035), .B(n21036), .Z(n20958) );
  OR U25624 ( .A(n21037), .B(n21038), .Z(n21036) );
  OR U25625 ( .A(n21039), .B(n21040), .Z(n21035) );
  NOR U25626 ( .A(n21041), .B(n21042), .Z(n20959) );
  ANDN U25627 ( .B(n21043), .A(n21044), .Z(n20953) );
  IV U25628 ( .A(n21045), .Z(n21043) );
  XNOR U25629 ( .A(n20946), .B(n21046), .Z(n20952) );
  XNOR U25630 ( .A(n20945), .B(n20947), .Z(n21046) );
  NAND U25631 ( .A(n21047), .B(n21048), .Z(n20947) );
  OR U25632 ( .A(n21049), .B(n21050), .Z(n21048) );
  OR U25633 ( .A(n21051), .B(n21052), .Z(n21047) );
  NAND U25634 ( .A(n21053), .B(n21054), .Z(n20945) );
  OR U25635 ( .A(n21055), .B(n21056), .Z(n21054) );
  OR U25636 ( .A(n21057), .B(n21058), .Z(n21053) );
  ANDN U25637 ( .B(n21059), .A(n21060), .Z(n20946) );
  IV U25638 ( .A(n21061), .Z(n21059) );
  XNOR U25639 ( .A(n21026), .B(n21025), .Z(N28433) );
  XOR U25640 ( .A(n21045), .B(n21044), .Z(n21025) );
  XNOR U25641 ( .A(n21060), .B(n21061), .Z(n21044) );
  XNOR U25642 ( .A(n21055), .B(n21056), .Z(n21061) );
  XNOR U25643 ( .A(n21057), .B(n21058), .Z(n21056) );
  XNOR U25644 ( .A(y[1012]), .B(x[1012]), .Z(n21058) );
  XNOR U25645 ( .A(y[1013]), .B(x[1013]), .Z(n21057) );
  XNOR U25646 ( .A(y[1011]), .B(x[1011]), .Z(n21055) );
  XNOR U25647 ( .A(n21049), .B(n21050), .Z(n21060) );
  XNOR U25648 ( .A(y[1008]), .B(x[1008]), .Z(n21050) );
  XNOR U25649 ( .A(n21051), .B(n21052), .Z(n21049) );
  XNOR U25650 ( .A(y[1009]), .B(x[1009]), .Z(n21052) );
  XNOR U25651 ( .A(y[1010]), .B(x[1010]), .Z(n21051) );
  XNOR U25652 ( .A(n21042), .B(n21041), .Z(n21045) );
  XNOR U25653 ( .A(n21037), .B(n21038), .Z(n21041) );
  XNOR U25654 ( .A(y[1005]), .B(x[1005]), .Z(n21038) );
  XNOR U25655 ( .A(n21039), .B(n21040), .Z(n21037) );
  XNOR U25656 ( .A(y[1006]), .B(x[1006]), .Z(n21040) );
  XNOR U25657 ( .A(y[1007]), .B(x[1007]), .Z(n21039) );
  XNOR U25658 ( .A(n21031), .B(n21032), .Z(n21042) );
  XNOR U25659 ( .A(y[1002]), .B(x[1002]), .Z(n21032) );
  XNOR U25660 ( .A(n21033), .B(n21034), .Z(n21031) );
  XNOR U25661 ( .A(y[1003]), .B(x[1003]), .Z(n21034) );
  XNOR U25662 ( .A(y[1004]), .B(x[1004]), .Z(n21033) );
  XOR U25663 ( .A(n21007), .B(n21008), .Z(n21026) );
  XNOR U25664 ( .A(n21023), .B(n21024), .Z(n21008) );
  XNOR U25665 ( .A(n21018), .B(n21019), .Z(n21024) );
  XNOR U25666 ( .A(n21020), .B(n21021), .Z(n21019) );
  XNOR U25667 ( .A(y[1000]), .B(x[1000]), .Z(n21021) );
  XNOR U25668 ( .A(y[1001]), .B(x[1001]), .Z(n21020) );
  XNOR U25669 ( .A(y[999]), .B(x[999]), .Z(n21018) );
  XNOR U25670 ( .A(n21012), .B(n21013), .Z(n21023) );
  XNOR U25671 ( .A(y[996]), .B(x[996]), .Z(n21013) );
  XNOR U25672 ( .A(n21014), .B(n21015), .Z(n21012) );
  XNOR U25673 ( .A(y[997]), .B(x[997]), .Z(n21015) );
  XNOR U25674 ( .A(y[998]), .B(x[998]), .Z(n21014) );
  XOR U25675 ( .A(n21006), .B(n21005), .Z(n21007) );
  XNOR U25676 ( .A(n21001), .B(n21002), .Z(n21005) );
  XNOR U25677 ( .A(y[993]), .B(x[993]), .Z(n21002) );
  XNOR U25678 ( .A(n21003), .B(n21004), .Z(n21001) );
  XNOR U25679 ( .A(y[994]), .B(x[994]), .Z(n21004) );
  XNOR U25680 ( .A(y[995]), .B(x[995]), .Z(n21003) );
  XNOR U25681 ( .A(n20995), .B(n20996), .Z(n21006) );
  XNOR U25682 ( .A(y[990]), .B(x[990]), .Z(n20996) );
  XNOR U25683 ( .A(n20997), .B(n20998), .Z(n20995) );
  XNOR U25684 ( .A(y[991]), .B(x[991]), .Z(n20998) );
  XNOR U25685 ( .A(y[992]), .B(x[992]), .Z(n20997) );
  NAND U25686 ( .A(n21062), .B(n21063), .Z(N28425) );
  NANDN U25687 ( .A(n21064), .B(n21065), .Z(n21063) );
  OR U25688 ( .A(n21066), .B(n21067), .Z(n21065) );
  NAND U25689 ( .A(n21066), .B(n21067), .Z(n21062) );
  XOR U25690 ( .A(n21066), .B(n21068), .Z(N28424) );
  XNOR U25691 ( .A(n21064), .B(n21067), .Z(n21068) );
  AND U25692 ( .A(n21069), .B(n21070), .Z(n21067) );
  NANDN U25693 ( .A(n21071), .B(n21072), .Z(n21070) );
  NANDN U25694 ( .A(n21073), .B(n21074), .Z(n21072) );
  NANDN U25695 ( .A(n21074), .B(n21073), .Z(n21069) );
  NAND U25696 ( .A(n21075), .B(n21076), .Z(n21064) );
  NANDN U25697 ( .A(n21077), .B(n21078), .Z(n21076) );
  OR U25698 ( .A(n21079), .B(n21080), .Z(n21078) );
  NAND U25699 ( .A(n21080), .B(n21079), .Z(n21075) );
  AND U25700 ( .A(n21081), .B(n21082), .Z(n21066) );
  NANDN U25701 ( .A(n21083), .B(n21084), .Z(n21082) );
  NANDN U25702 ( .A(n21085), .B(n21086), .Z(n21084) );
  NANDN U25703 ( .A(n21086), .B(n21085), .Z(n21081) );
  XOR U25704 ( .A(n21080), .B(n21087), .Z(N28423) );
  XOR U25705 ( .A(n21077), .B(n21079), .Z(n21087) );
  XNOR U25706 ( .A(n21073), .B(n21088), .Z(n21079) );
  XNOR U25707 ( .A(n21071), .B(n21074), .Z(n21088) );
  NAND U25708 ( .A(n21089), .B(n21090), .Z(n21074) );
  NAND U25709 ( .A(n21091), .B(n21092), .Z(n21090) );
  OR U25710 ( .A(n21093), .B(n21094), .Z(n21091) );
  NANDN U25711 ( .A(n21095), .B(n21093), .Z(n21089) );
  IV U25712 ( .A(n21094), .Z(n21095) );
  NAND U25713 ( .A(n21096), .B(n21097), .Z(n21071) );
  NAND U25714 ( .A(n21098), .B(n21099), .Z(n21097) );
  NANDN U25715 ( .A(n21100), .B(n21101), .Z(n21098) );
  NANDN U25716 ( .A(n21101), .B(n21100), .Z(n21096) );
  AND U25717 ( .A(n21102), .B(n21103), .Z(n21073) );
  NAND U25718 ( .A(n21104), .B(n21105), .Z(n21103) );
  OR U25719 ( .A(n21106), .B(n21107), .Z(n21104) );
  NANDN U25720 ( .A(n21108), .B(n21106), .Z(n21102) );
  NAND U25721 ( .A(n21109), .B(n21110), .Z(n21077) );
  NANDN U25722 ( .A(n21111), .B(n21112), .Z(n21110) );
  OR U25723 ( .A(n21113), .B(n21114), .Z(n21112) );
  NANDN U25724 ( .A(n21115), .B(n21113), .Z(n21109) );
  IV U25725 ( .A(n21114), .Z(n21115) );
  XNOR U25726 ( .A(n21085), .B(n21116), .Z(n21080) );
  XNOR U25727 ( .A(n21083), .B(n21086), .Z(n21116) );
  NAND U25728 ( .A(n21117), .B(n21118), .Z(n21086) );
  NAND U25729 ( .A(n21119), .B(n21120), .Z(n21118) );
  OR U25730 ( .A(n21121), .B(n21122), .Z(n21119) );
  NANDN U25731 ( .A(n21123), .B(n21121), .Z(n21117) );
  IV U25732 ( .A(n21122), .Z(n21123) );
  NAND U25733 ( .A(n21124), .B(n21125), .Z(n21083) );
  NAND U25734 ( .A(n21126), .B(n21127), .Z(n21125) );
  NANDN U25735 ( .A(n21128), .B(n21129), .Z(n21126) );
  NANDN U25736 ( .A(n21129), .B(n21128), .Z(n21124) );
  AND U25737 ( .A(n21130), .B(n21131), .Z(n21085) );
  NAND U25738 ( .A(n21132), .B(n21133), .Z(n21131) );
  OR U25739 ( .A(n21134), .B(n21135), .Z(n21132) );
  NANDN U25740 ( .A(n21136), .B(n21134), .Z(n21130) );
  XNOR U25741 ( .A(n21111), .B(n21137), .Z(N28422) );
  XOR U25742 ( .A(n21113), .B(n21114), .Z(n21137) );
  XNOR U25743 ( .A(n21127), .B(n21138), .Z(n21114) );
  XOR U25744 ( .A(n21128), .B(n21129), .Z(n21138) );
  XOR U25745 ( .A(n21134), .B(n21139), .Z(n21129) );
  XOR U25746 ( .A(n21133), .B(n21136), .Z(n21139) );
  IV U25747 ( .A(n21135), .Z(n21136) );
  NAND U25748 ( .A(n21140), .B(n21141), .Z(n21135) );
  OR U25749 ( .A(n21142), .B(n21143), .Z(n21141) );
  OR U25750 ( .A(n21144), .B(n21145), .Z(n21140) );
  NAND U25751 ( .A(n21146), .B(n21147), .Z(n21133) );
  OR U25752 ( .A(n21148), .B(n21149), .Z(n21147) );
  OR U25753 ( .A(n21150), .B(n21151), .Z(n21146) );
  NOR U25754 ( .A(n21152), .B(n21153), .Z(n21134) );
  ANDN U25755 ( .B(n21154), .A(n21155), .Z(n21128) );
  XNOR U25756 ( .A(n21121), .B(n21156), .Z(n21127) );
  XNOR U25757 ( .A(n21120), .B(n21122), .Z(n21156) );
  NAND U25758 ( .A(n21157), .B(n21158), .Z(n21122) );
  OR U25759 ( .A(n21159), .B(n21160), .Z(n21158) );
  OR U25760 ( .A(n21161), .B(n21162), .Z(n21157) );
  NAND U25761 ( .A(n21163), .B(n21164), .Z(n21120) );
  OR U25762 ( .A(n21165), .B(n21166), .Z(n21164) );
  OR U25763 ( .A(n21167), .B(n21168), .Z(n21163) );
  ANDN U25764 ( .B(n21169), .A(n21170), .Z(n21121) );
  IV U25765 ( .A(n21171), .Z(n21169) );
  ANDN U25766 ( .B(n21172), .A(n21173), .Z(n21113) );
  XOR U25767 ( .A(n21099), .B(n21174), .Z(n21111) );
  XOR U25768 ( .A(n21100), .B(n21101), .Z(n21174) );
  XOR U25769 ( .A(n21106), .B(n21175), .Z(n21101) );
  XOR U25770 ( .A(n21105), .B(n21108), .Z(n21175) );
  IV U25771 ( .A(n21107), .Z(n21108) );
  NAND U25772 ( .A(n21176), .B(n21177), .Z(n21107) );
  OR U25773 ( .A(n21178), .B(n21179), .Z(n21177) );
  OR U25774 ( .A(n21180), .B(n21181), .Z(n21176) );
  NAND U25775 ( .A(n21182), .B(n21183), .Z(n21105) );
  OR U25776 ( .A(n21184), .B(n21185), .Z(n21183) );
  OR U25777 ( .A(n21186), .B(n21187), .Z(n21182) );
  NOR U25778 ( .A(n21188), .B(n21189), .Z(n21106) );
  ANDN U25779 ( .B(n21190), .A(n21191), .Z(n21100) );
  IV U25780 ( .A(n21192), .Z(n21190) );
  XNOR U25781 ( .A(n21093), .B(n21193), .Z(n21099) );
  XNOR U25782 ( .A(n21092), .B(n21094), .Z(n21193) );
  NAND U25783 ( .A(n21194), .B(n21195), .Z(n21094) );
  OR U25784 ( .A(n21196), .B(n21197), .Z(n21195) );
  OR U25785 ( .A(n21198), .B(n21199), .Z(n21194) );
  NAND U25786 ( .A(n21200), .B(n21201), .Z(n21092) );
  OR U25787 ( .A(n21202), .B(n21203), .Z(n21201) );
  OR U25788 ( .A(n21204), .B(n21205), .Z(n21200) );
  ANDN U25789 ( .B(n21206), .A(n21207), .Z(n21093) );
  IV U25790 ( .A(n21208), .Z(n21206) );
  XNOR U25791 ( .A(n21173), .B(n21172), .Z(N28421) );
  XOR U25792 ( .A(n21192), .B(n21191), .Z(n21172) );
  XNOR U25793 ( .A(n21207), .B(n21208), .Z(n21191) );
  XNOR U25794 ( .A(n21202), .B(n21203), .Z(n21208) );
  XNOR U25795 ( .A(n21204), .B(n21205), .Z(n21203) );
  XNOR U25796 ( .A(y[988]), .B(x[988]), .Z(n21205) );
  XNOR U25797 ( .A(y[989]), .B(x[989]), .Z(n21204) );
  XNOR U25798 ( .A(y[987]), .B(x[987]), .Z(n21202) );
  XNOR U25799 ( .A(n21196), .B(n21197), .Z(n21207) );
  XNOR U25800 ( .A(y[984]), .B(x[984]), .Z(n21197) );
  XNOR U25801 ( .A(n21198), .B(n21199), .Z(n21196) );
  XNOR U25802 ( .A(y[985]), .B(x[985]), .Z(n21199) );
  XNOR U25803 ( .A(y[986]), .B(x[986]), .Z(n21198) );
  XNOR U25804 ( .A(n21189), .B(n21188), .Z(n21192) );
  XNOR U25805 ( .A(n21184), .B(n21185), .Z(n21188) );
  XNOR U25806 ( .A(y[981]), .B(x[981]), .Z(n21185) );
  XNOR U25807 ( .A(n21186), .B(n21187), .Z(n21184) );
  XNOR U25808 ( .A(y[982]), .B(x[982]), .Z(n21187) );
  XNOR U25809 ( .A(y[983]), .B(x[983]), .Z(n21186) );
  XNOR U25810 ( .A(n21178), .B(n21179), .Z(n21189) );
  XNOR U25811 ( .A(y[978]), .B(x[978]), .Z(n21179) );
  XNOR U25812 ( .A(n21180), .B(n21181), .Z(n21178) );
  XNOR U25813 ( .A(y[979]), .B(x[979]), .Z(n21181) );
  XNOR U25814 ( .A(y[980]), .B(x[980]), .Z(n21180) );
  XOR U25815 ( .A(n21154), .B(n21155), .Z(n21173) );
  XNOR U25816 ( .A(n21170), .B(n21171), .Z(n21155) );
  XNOR U25817 ( .A(n21165), .B(n21166), .Z(n21171) );
  XNOR U25818 ( .A(n21167), .B(n21168), .Z(n21166) );
  XNOR U25819 ( .A(y[976]), .B(x[976]), .Z(n21168) );
  XNOR U25820 ( .A(y[977]), .B(x[977]), .Z(n21167) );
  XNOR U25821 ( .A(y[975]), .B(x[975]), .Z(n21165) );
  XNOR U25822 ( .A(n21159), .B(n21160), .Z(n21170) );
  XNOR U25823 ( .A(y[972]), .B(x[972]), .Z(n21160) );
  XNOR U25824 ( .A(n21161), .B(n21162), .Z(n21159) );
  XNOR U25825 ( .A(y[973]), .B(x[973]), .Z(n21162) );
  XNOR U25826 ( .A(y[974]), .B(x[974]), .Z(n21161) );
  XOR U25827 ( .A(n21153), .B(n21152), .Z(n21154) );
  XNOR U25828 ( .A(n21148), .B(n21149), .Z(n21152) );
  XNOR U25829 ( .A(y[969]), .B(x[969]), .Z(n21149) );
  XNOR U25830 ( .A(n21150), .B(n21151), .Z(n21148) );
  XNOR U25831 ( .A(y[970]), .B(x[970]), .Z(n21151) );
  XNOR U25832 ( .A(y[971]), .B(x[971]), .Z(n21150) );
  XNOR U25833 ( .A(n21142), .B(n21143), .Z(n21153) );
  XNOR U25834 ( .A(y[966]), .B(x[966]), .Z(n21143) );
  XNOR U25835 ( .A(n21144), .B(n21145), .Z(n21142) );
  XNOR U25836 ( .A(y[967]), .B(x[967]), .Z(n21145) );
  XNOR U25837 ( .A(y[968]), .B(x[968]), .Z(n21144) );
  NAND U25838 ( .A(n21209), .B(n21210), .Z(N28413) );
  NANDN U25839 ( .A(n21211), .B(n21212), .Z(n21210) );
  OR U25840 ( .A(n21213), .B(n21214), .Z(n21212) );
  NAND U25841 ( .A(n21213), .B(n21214), .Z(n21209) );
  XOR U25842 ( .A(n21213), .B(n21215), .Z(N28412) );
  XNOR U25843 ( .A(n21211), .B(n21214), .Z(n21215) );
  AND U25844 ( .A(n21216), .B(n21217), .Z(n21214) );
  NANDN U25845 ( .A(n21218), .B(n21219), .Z(n21217) );
  NANDN U25846 ( .A(n21220), .B(n21221), .Z(n21219) );
  NANDN U25847 ( .A(n21221), .B(n21220), .Z(n21216) );
  NAND U25848 ( .A(n21222), .B(n21223), .Z(n21211) );
  NANDN U25849 ( .A(n21224), .B(n21225), .Z(n21223) );
  OR U25850 ( .A(n21226), .B(n21227), .Z(n21225) );
  NAND U25851 ( .A(n21227), .B(n21226), .Z(n21222) );
  AND U25852 ( .A(n21228), .B(n21229), .Z(n21213) );
  NANDN U25853 ( .A(n21230), .B(n21231), .Z(n21229) );
  NANDN U25854 ( .A(n21232), .B(n21233), .Z(n21231) );
  NANDN U25855 ( .A(n21233), .B(n21232), .Z(n21228) );
  XOR U25856 ( .A(n21227), .B(n21234), .Z(N28411) );
  XOR U25857 ( .A(n21224), .B(n21226), .Z(n21234) );
  XNOR U25858 ( .A(n21220), .B(n21235), .Z(n21226) );
  XNOR U25859 ( .A(n21218), .B(n21221), .Z(n21235) );
  NAND U25860 ( .A(n21236), .B(n21237), .Z(n21221) );
  NAND U25861 ( .A(n21238), .B(n21239), .Z(n21237) );
  OR U25862 ( .A(n21240), .B(n21241), .Z(n21238) );
  NANDN U25863 ( .A(n21242), .B(n21240), .Z(n21236) );
  IV U25864 ( .A(n21241), .Z(n21242) );
  NAND U25865 ( .A(n21243), .B(n21244), .Z(n21218) );
  NAND U25866 ( .A(n21245), .B(n21246), .Z(n21244) );
  NANDN U25867 ( .A(n21247), .B(n21248), .Z(n21245) );
  NANDN U25868 ( .A(n21248), .B(n21247), .Z(n21243) );
  AND U25869 ( .A(n21249), .B(n21250), .Z(n21220) );
  NAND U25870 ( .A(n21251), .B(n21252), .Z(n21250) );
  OR U25871 ( .A(n21253), .B(n21254), .Z(n21251) );
  NANDN U25872 ( .A(n21255), .B(n21253), .Z(n21249) );
  NAND U25873 ( .A(n21256), .B(n21257), .Z(n21224) );
  NANDN U25874 ( .A(n21258), .B(n21259), .Z(n21257) );
  OR U25875 ( .A(n21260), .B(n21261), .Z(n21259) );
  NANDN U25876 ( .A(n21262), .B(n21260), .Z(n21256) );
  IV U25877 ( .A(n21261), .Z(n21262) );
  XNOR U25878 ( .A(n21232), .B(n21263), .Z(n21227) );
  XNOR U25879 ( .A(n21230), .B(n21233), .Z(n21263) );
  NAND U25880 ( .A(n21264), .B(n21265), .Z(n21233) );
  NAND U25881 ( .A(n21266), .B(n21267), .Z(n21265) );
  OR U25882 ( .A(n21268), .B(n21269), .Z(n21266) );
  NANDN U25883 ( .A(n21270), .B(n21268), .Z(n21264) );
  IV U25884 ( .A(n21269), .Z(n21270) );
  NAND U25885 ( .A(n21271), .B(n21272), .Z(n21230) );
  NAND U25886 ( .A(n21273), .B(n21274), .Z(n21272) );
  NANDN U25887 ( .A(n21275), .B(n21276), .Z(n21273) );
  NANDN U25888 ( .A(n21276), .B(n21275), .Z(n21271) );
  AND U25889 ( .A(n21277), .B(n21278), .Z(n21232) );
  NAND U25890 ( .A(n21279), .B(n21280), .Z(n21278) );
  OR U25891 ( .A(n21281), .B(n21282), .Z(n21279) );
  NANDN U25892 ( .A(n21283), .B(n21281), .Z(n21277) );
  XNOR U25893 ( .A(n21258), .B(n21284), .Z(N28410) );
  XOR U25894 ( .A(n21260), .B(n21261), .Z(n21284) );
  XNOR U25895 ( .A(n21274), .B(n21285), .Z(n21261) );
  XOR U25896 ( .A(n21275), .B(n21276), .Z(n21285) );
  XOR U25897 ( .A(n21281), .B(n21286), .Z(n21276) );
  XOR U25898 ( .A(n21280), .B(n21283), .Z(n21286) );
  IV U25899 ( .A(n21282), .Z(n21283) );
  NAND U25900 ( .A(n21287), .B(n21288), .Z(n21282) );
  OR U25901 ( .A(n21289), .B(n21290), .Z(n21288) );
  OR U25902 ( .A(n21291), .B(n21292), .Z(n21287) );
  NAND U25903 ( .A(n21293), .B(n21294), .Z(n21280) );
  OR U25904 ( .A(n21295), .B(n21296), .Z(n21294) );
  OR U25905 ( .A(n21297), .B(n21298), .Z(n21293) );
  NOR U25906 ( .A(n21299), .B(n21300), .Z(n21281) );
  ANDN U25907 ( .B(n21301), .A(n21302), .Z(n21275) );
  XNOR U25908 ( .A(n21268), .B(n21303), .Z(n21274) );
  XNOR U25909 ( .A(n21267), .B(n21269), .Z(n21303) );
  NAND U25910 ( .A(n21304), .B(n21305), .Z(n21269) );
  OR U25911 ( .A(n21306), .B(n21307), .Z(n21305) );
  OR U25912 ( .A(n21308), .B(n21309), .Z(n21304) );
  NAND U25913 ( .A(n21310), .B(n21311), .Z(n21267) );
  OR U25914 ( .A(n21312), .B(n21313), .Z(n21311) );
  OR U25915 ( .A(n21314), .B(n21315), .Z(n21310) );
  ANDN U25916 ( .B(n21316), .A(n21317), .Z(n21268) );
  IV U25917 ( .A(n21318), .Z(n21316) );
  ANDN U25918 ( .B(n21319), .A(n21320), .Z(n21260) );
  XOR U25919 ( .A(n21246), .B(n21321), .Z(n21258) );
  XOR U25920 ( .A(n21247), .B(n21248), .Z(n21321) );
  XOR U25921 ( .A(n21253), .B(n21322), .Z(n21248) );
  XOR U25922 ( .A(n21252), .B(n21255), .Z(n21322) );
  IV U25923 ( .A(n21254), .Z(n21255) );
  NAND U25924 ( .A(n21323), .B(n21324), .Z(n21254) );
  OR U25925 ( .A(n21325), .B(n21326), .Z(n21324) );
  OR U25926 ( .A(n21327), .B(n21328), .Z(n21323) );
  NAND U25927 ( .A(n21329), .B(n21330), .Z(n21252) );
  OR U25928 ( .A(n21331), .B(n21332), .Z(n21330) );
  OR U25929 ( .A(n21333), .B(n21334), .Z(n21329) );
  NOR U25930 ( .A(n21335), .B(n21336), .Z(n21253) );
  ANDN U25931 ( .B(n21337), .A(n21338), .Z(n21247) );
  IV U25932 ( .A(n21339), .Z(n21337) );
  XNOR U25933 ( .A(n21240), .B(n21340), .Z(n21246) );
  XNOR U25934 ( .A(n21239), .B(n21241), .Z(n21340) );
  NAND U25935 ( .A(n21341), .B(n21342), .Z(n21241) );
  OR U25936 ( .A(n21343), .B(n21344), .Z(n21342) );
  OR U25937 ( .A(n21345), .B(n21346), .Z(n21341) );
  NAND U25938 ( .A(n21347), .B(n21348), .Z(n21239) );
  OR U25939 ( .A(n21349), .B(n21350), .Z(n21348) );
  OR U25940 ( .A(n21351), .B(n21352), .Z(n21347) );
  ANDN U25941 ( .B(n21353), .A(n21354), .Z(n21240) );
  IV U25942 ( .A(n21355), .Z(n21353) );
  XNOR U25943 ( .A(n21320), .B(n21319), .Z(N28409) );
  XOR U25944 ( .A(n21339), .B(n21338), .Z(n21319) );
  XNOR U25945 ( .A(n21354), .B(n21355), .Z(n21338) );
  XNOR U25946 ( .A(n21349), .B(n21350), .Z(n21355) );
  XNOR U25947 ( .A(n21351), .B(n21352), .Z(n21350) );
  XNOR U25948 ( .A(y[964]), .B(x[964]), .Z(n21352) );
  XNOR U25949 ( .A(y[965]), .B(x[965]), .Z(n21351) );
  XNOR U25950 ( .A(y[963]), .B(x[963]), .Z(n21349) );
  XNOR U25951 ( .A(n21343), .B(n21344), .Z(n21354) );
  XNOR U25952 ( .A(y[960]), .B(x[960]), .Z(n21344) );
  XNOR U25953 ( .A(n21345), .B(n21346), .Z(n21343) );
  XNOR U25954 ( .A(y[961]), .B(x[961]), .Z(n21346) );
  XNOR U25955 ( .A(y[962]), .B(x[962]), .Z(n21345) );
  XNOR U25956 ( .A(n21336), .B(n21335), .Z(n21339) );
  XNOR U25957 ( .A(n21331), .B(n21332), .Z(n21335) );
  XNOR U25958 ( .A(y[957]), .B(x[957]), .Z(n21332) );
  XNOR U25959 ( .A(n21333), .B(n21334), .Z(n21331) );
  XNOR U25960 ( .A(y[958]), .B(x[958]), .Z(n21334) );
  XNOR U25961 ( .A(y[959]), .B(x[959]), .Z(n21333) );
  XNOR U25962 ( .A(n21325), .B(n21326), .Z(n21336) );
  XNOR U25963 ( .A(y[954]), .B(x[954]), .Z(n21326) );
  XNOR U25964 ( .A(n21327), .B(n21328), .Z(n21325) );
  XNOR U25965 ( .A(y[955]), .B(x[955]), .Z(n21328) );
  XNOR U25966 ( .A(y[956]), .B(x[956]), .Z(n21327) );
  XOR U25967 ( .A(n21301), .B(n21302), .Z(n21320) );
  XNOR U25968 ( .A(n21317), .B(n21318), .Z(n21302) );
  XNOR U25969 ( .A(n21312), .B(n21313), .Z(n21318) );
  XNOR U25970 ( .A(n21314), .B(n21315), .Z(n21313) );
  XNOR U25971 ( .A(y[952]), .B(x[952]), .Z(n21315) );
  XNOR U25972 ( .A(y[953]), .B(x[953]), .Z(n21314) );
  XNOR U25973 ( .A(y[951]), .B(x[951]), .Z(n21312) );
  XNOR U25974 ( .A(n21306), .B(n21307), .Z(n21317) );
  XNOR U25975 ( .A(y[948]), .B(x[948]), .Z(n21307) );
  XNOR U25976 ( .A(n21308), .B(n21309), .Z(n21306) );
  XNOR U25977 ( .A(y[949]), .B(x[949]), .Z(n21309) );
  XNOR U25978 ( .A(y[950]), .B(x[950]), .Z(n21308) );
  XOR U25979 ( .A(n21300), .B(n21299), .Z(n21301) );
  XNOR U25980 ( .A(n21295), .B(n21296), .Z(n21299) );
  XNOR U25981 ( .A(y[945]), .B(x[945]), .Z(n21296) );
  XNOR U25982 ( .A(n21297), .B(n21298), .Z(n21295) );
  XNOR U25983 ( .A(y[946]), .B(x[946]), .Z(n21298) );
  XNOR U25984 ( .A(y[947]), .B(x[947]), .Z(n21297) );
  XNOR U25985 ( .A(n21289), .B(n21290), .Z(n21300) );
  XNOR U25986 ( .A(y[942]), .B(x[942]), .Z(n21290) );
  XNOR U25987 ( .A(n21291), .B(n21292), .Z(n21289) );
  XNOR U25988 ( .A(y[943]), .B(x[943]), .Z(n21292) );
  XNOR U25989 ( .A(y[944]), .B(x[944]), .Z(n21291) );
  NAND U25990 ( .A(n21356), .B(n21357), .Z(N28401) );
  NANDN U25991 ( .A(n21358), .B(n21359), .Z(n21357) );
  OR U25992 ( .A(n21360), .B(n21361), .Z(n21359) );
  NAND U25993 ( .A(n21360), .B(n21361), .Z(n21356) );
  XOR U25994 ( .A(n21360), .B(n21362), .Z(N28400) );
  XNOR U25995 ( .A(n21358), .B(n21361), .Z(n21362) );
  AND U25996 ( .A(n21363), .B(n21364), .Z(n21361) );
  NANDN U25997 ( .A(n21365), .B(n21366), .Z(n21364) );
  NANDN U25998 ( .A(n21367), .B(n21368), .Z(n21366) );
  NANDN U25999 ( .A(n21368), .B(n21367), .Z(n21363) );
  NAND U26000 ( .A(n21369), .B(n21370), .Z(n21358) );
  NANDN U26001 ( .A(n21371), .B(n21372), .Z(n21370) );
  OR U26002 ( .A(n21373), .B(n21374), .Z(n21372) );
  NAND U26003 ( .A(n21374), .B(n21373), .Z(n21369) );
  AND U26004 ( .A(n21375), .B(n21376), .Z(n21360) );
  NANDN U26005 ( .A(n21377), .B(n21378), .Z(n21376) );
  NANDN U26006 ( .A(n21379), .B(n21380), .Z(n21378) );
  NANDN U26007 ( .A(n21380), .B(n21379), .Z(n21375) );
  XOR U26008 ( .A(n21374), .B(n21381), .Z(N28399) );
  XOR U26009 ( .A(n21371), .B(n21373), .Z(n21381) );
  XNOR U26010 ( .A(n21367), .B(n21382), .Z(n21373) );
  XNOR U26011 ( .A(n21365), .B(n21368), .Z(n21382) );
  NAND U26012 ( .A(n21383), .B(n21384), .Z(n21368) );
  NAND U26013 ( .A(n21385), .B(n21386), .Z(n21384) );
  OR U26014 ( .A(n21387), .B(n21388), .Z(n21385) );
  NANDN U26015 ( .A(n21389), .B(n21387), .Z(n21383) );
  IV U26016 ( .A(n21388), .Z(n21389) );
  NAND U26017 ( .A(n21390), .B(n21391), .Z(n21365) );
  NAND U26018 ( .A(n21392), .B(n21393), .Z(n21391) );
  NANDN U26019 ( .A(n21394), .B(n21395), .Z(n21392) );
  NANDN U26020 ( .A(n21395), .B(n21394), .Z(n21390) );
  AND U26021 ( .A(n21396), .B(n21397), .Z(n21367) );
  NAND U26022 ( .A(n21398), .B(n21399), .Z(n21397) );
  OR U26023 ( .A(n21400), .B(n21401), .Z(n21398) );
  NANDN U26024 ( .A(n21402), .B(n21400), .Z(n21396) );
  NAND U26025 ( .A(n21403), .B(n21404), .Z(n21371) );
  NANDN U26026 ( .A(n21405), .B(n21406), .Z(n21404) );
  OR U26027 ( .A(n21407), .B(n21408), .Z(n21406) );
  NANDN U26028 ( .A(n21409), .B(n21407), .Z(n21403) );
  IV U26029 ( .A(n21408), .Z(n21409) );
  XNOR U26030 ( .A(n21379), .B(n21410), .Z(n21374) );
  XNOR U26031 ( .A(n21377), .B(n21380), .Z(n21410) );
  NAND U26032 ( .A(n21411), .B(n21412), .Z(n21380) );
  NAND U26033 ( .A(n21413), .B(n21414), .Z(n21412) );
  OR U26034 ( .A(n21415), .B(n21416), .Z(n21413) );
  NANDN U26035 ( .A(n21417), .B(n21415), .Z(n21411) );
  IV U26036 ( .A(n21416), .Z(n21417) );
  NAND U26037 ( .A(n21418), .B(n21419), .Z(n21377) );
  NAND U26038 ( .A(n21420), .B(n21421), .Z(n21419) );
  NANDN U26039 ( .A(n21422), .B(n21423), .Z(n21420) );
  NANDN U26040 ( .A(n21423), .B(n21422), .Z(n21418) );
  AND U26041 ( .A(n21424), .B(n21425), .Z(n21379) );
  NAND U26042 ( .A(n21426), .B(n21427), .Z(n21425) );
  OR U26043 ( .A(n21428), .B(n21429), .Z(n21426) );
  NANDN U26044 ( .A(n21430), .B(n21428), .Z(n21424) );
  XNOR U26045 ( .A(n21405), .B(n21431), .Z(N28398) );
  XOR U26046 ( .A(n21407), .B(n21408), .Z(n21431) );
  XNOR U26047 ( .A(n21421), .B(n21432), .Z(n21408) );
  XOR U26048 ( .A(n21422), .B(n21423), .Z(n21432) );
  XOR U26049 ( .A(n21428), .B(n21433), .Z(n21423) );
  XOR U26050 ( .A(n21427), .B(n21430), .Z(n21433) );
  IV U26051 ( .A(n21429), .Z(n21430) );
  NAND U26052 ( .A(n21434), .B(n21435), .Z(n21429) );
  OR U26053 ( .A(n21436), .B(n21437), .Z(n21435) );
  OR U26054 ( .A(n21438), .B(n21439), .Z(n21434) );
  NAND U26055 ( .A(n21440), .B(n21441), .Z(n21427) );
  OR U26056 ( .A(n21442), .B(n21443), .Z(n21441) );
  OR U26057 ( .A(n21444), .B(n21445), .Z(n21440) );
  NOR U26058 ( .A(n21446), .B(n21447), .Z(n21428) );
  ANDN U26059 ( .B(n21448), .A(n21449), .Z(n21422) );
  XNOR U26060 ( .A(n21415), .B(n21450), .Z(n21421) );
  XNOR U26061 ( .A(n21414), .B(n21416), .Z(n21450) );
  NAND U26062 ( .A(n21451), .B(n21452), .Z(n21416) );
  OR U26063 ( .A(n21453), .B(n21454), .Z(n21452) );
  OR U26064 ( .A(n21455), .B(n21456), .Z(n21451) );
  NAND U26065 ( .A(n21457), .B(n21458), .Z(n21414) );
  OR U26066 ( .A(n21459), .B(n21460), .Z(n21458) );
  OR U26067 ( .A(n21461), .B(n21462), .Z(n21457) );
  ANDN U26068 ( .B(n21463), .A(n21464), .Z(n21415) );
  IV U26069 ( .A(n21465), .Z(n21463) );
  ANDN U26070 ( .B(n21466), .A(n21467), .Z(n21407) );
  XOR U26071 ( .A(n21393), .B(n21468), .Z(n21405) );
  XOR U26072 ( .A(n21394), .B(n21395), .Z(n21468) );
  XOR U26073 ( .A(n21400), .B(n21469), .Z(n21395) );
  XOR U26074 ( .A(n21399), .B(n21402), .Z(n21469) );
  IV U26075 ( .A(n21401), .Z(n21402) );
  NAND U26076 ( .A(n21470), .B(n21471), .Z(n21401) );
  OR U26077 ( .A(n21472), .B(n21473), .Z(n21471) );
  OR U26078 ( .A(n21474), .B(n21475), .Z(n21470) );
  NAND U26079 ( .A(n21476), .B(n21477), .Z(n21399) );
  OR U26080 ( .A(n21478), .B(n21479), .Z(n21477) );
  OR U26081 ( .A(n21480), .B(n21481), .Z(n21476) );
  NOR U26082 ( .A(n21482), .B(n21483), .Z(n21400) );
  ANDN U26083 ( .B(n21484), .A(n21485), .Z(n21394) );
  IV U26084 ( .A(n21486), .Z(n21484) );
  XNOR U26085 ( .A(n21387), .B(n21487), .Z(n21393) );
  XNOR U26086 ( .A(n21386), .B(n21388), .Z(n21487) );
  NAND U26087 ( .A(n21488), .B(n21489), .Z(n21388) );
  OR U26088 ( .A(n21490), .B(n21491), .Z(n21489) );
  OR U26089 ( .A(n21492), .B(n21493), .Z(n21488) );
  NAND U26090 ( .A(n21494), .B(n21495), .Z(n21386) );
  OR U26091 ( .A(n21496), .B(n21497), .Z(n21495) );
  OR U26092 ( .A(n21498), .B(n21499), .Z(n21494) );
  ANDN U26093 ( .B(n21500), .A(n21501), .Z(n21387) );
  IV U26094 ( .A(n21502), .Z(n21500) );
  XNOR U26095 ( .A(n21467), .B(n21466), .Z(N28397) );
  XOR U26096 ( .A(n21486), .B(n21485), .Z(n21466) );
  XNOR U26097 ( .A(n21501), .B(n21502), .Z(n21485) );
  XNOR U26098 ( .A(n21496), .B(n21497), .Z(n21502) );
  XNOR U26099 ( .A(n21498), .B(n21499), .Z(n21497) );
  XNOR U26100 ( .A(y[940]), .B(x[940]), .Z(n21499) );
  XNOR U26101 ( .A(y[941]), .B(x[941]), .Z(n21498) );
  XNOR U26102 ( .A(y[939]), .B(x[939]), .Z(n21496) );
  XNOR U26103 ( .A(n21490), .B(n21491), .Z(n21501) );
  XNOR U26104 ( .A(y[936]), .B(x[936]), .Z(n21491) );
  XNOR U26105 ( .A(n21492), .B(n21493), .Z(n21490) );
  XNOR U26106 ( .A(y[937]), .B(x[937]), .Z(n21493) );
  XNOR U26107 ( .A(y[938]), .B(x[938]), .Z(n21492) );
  XNOR U26108 ( .A(n21483), .B(n21482), .Z(n21486) );
  XNOR U26109 ( .A(n21478), .B(n21479), .Z(n21482) );
  XNOR U26110 ( .A(y[933]), .B(x[933]), .Z(n21479) );
  XNOR U26111 ( .A(n21480), .B(n21481), .Z(n21478) );
  XNOR U26112 ( .A(y[934]), .B(x[934]), .Z(n21481) );
  XNOR U26113 ( .A(y[935]), .B(x[935]), .Z(n21480) );
  XNOR U26114 ( .A(n21472), .B(n21473), .Z(n21483) );
  XNOR U26115 ( .A(y[930]), .B(x[930]), .Z(n21473) );
  XNOR U26116 ( .A(n21474), .B(n21475), .Z(n21472) );
  XNOR U26117 ( .A(y[931]), .B(x[931]), .Z(n21475) );
  XNOR U26118 ( .A(y[932]), .B(x[932]), .Z(n21474) );
  XOR U26119 ( .A(n21448), .B(n21449), .Z(n21467) );
  XNOR U26120 ( .A(n21464), .B(n21465), .Z(n21449) );
  XNOR U26121 ( .A(n21459), .B(n21460), .Z(n21465) );
  XNOR U26122 ( .A(n21461), .B(n21462), .Z(n21460) );
  XNOR U26123 ( .A(y[928]), .B(x[928]), .Z(n21462) );
  XNOR U26124 ( .A(y[929]), .B(x[929]), .Z(n21461) );
  XNOR U26125 ( .A(y[927]), .B(x[927]), .Z(n21459) );
  XNOR U26126 ( .A(n21453), .B(n21454), .Z(n21464) );
  XNOR U26127 ( .A(y[924]), .B(x[924]), .Z(n21454) );
  XNOR U26128 ( .A(n21455), .B(n21456), .Z(n21453) );
  XNOR U26129 ( .A(y[925]), .B(x[925]), .Z(n21456) );
  XNOR U26130 ( .A(y[926]), .B(x[926]), .Z(n21455) );
  XOR U26131 ( .A(n21447), .B(n21446), .Z(n21448) );
  XNOR U26132 ( .A(n21442), .B(n21443), .Z(n21446) );
  XNOR U26133 ( .A(y[921]), .B(x[921]), .Z(n21443) );
  XNOR U26134 ( .A(n21444), .B(n21445), .Z(n21442) );
  XNOR U26135 ( .A(y[922]), .B(x[922]), .Z(n21445) );
  XNOR U26136 ( .A(y[923]), .B(x[923]), .Z(n21444) );
  XNOR U26137 ( .A(n21436), .B(n21437), .Z(n21447) );
  XNOR U26138 ( .A(y[918]), .B(x[918]), .Z(n21437) );
  XNOR U26139 ( .A(n21438), .B(n21439), .Z(n21436) );
  XNOR U26140 ( .A(y[919]), .B(x[919]), .Z(n21439) );
  XNOR U26141 ( .A(y[920]), .B(x[920]), .Z(n21438) );
  NAND U26142 ( .A(n21503), .B(n21504), .Z(N28389) );
  NANDN U26143 ( .A(n21505), .B(n21506), .Z(n21504) );
  OR U26144 ( .A(n21507), .B(n21508), .Z(n21506) );
  NAND U26145 ( .A(n21507), .B(n21508), .Z(n21503) );
  XOR U26146 ( .A(n21507), .B(n21509), .Z(N28388) );
  XNOR U26147 ( .A(n21505), .B(n21508), .Z(n21509) );
  AND U26148 ( .A(n21510), .B(n21511), .Z(n21508) );
  NANDN U26149 ( .A(n21512), .B(n21513), .Z(n21511) );
  NANDN U26150 ( .A(n21514), .B(n21515), .Z(n21513) );
  NANDN U26151 ( .A(n21515), .B(n21514), .Z(n21510) );
  NAND U26152 ( .A(n21516), .B(n21517), .Z(n21505) );
  NANDN U26153 ( .A(n21518), .B(n21519), .Z(n21517) );
  OR U26154 ( .A(n21520), .B(n21521), .Z(n21519) );
  NAND U26155 ( .A(n21521), .B(n21520), .Z(n21516) );
  AND U26156 ( .A(n21522), .B(n21523), .Z(n21507) );
  NANDN U26157 ( .A(n21524), .B(n21525), .Z(n21523) );
  NANDN U26158 ( .A(n21526), .B(n21527), .Z(n21525) );
  NANDN U26159 ( .A(n21527), .B(n21526), .Z(n21522) );
  XOR U26160 ( .A(n21521), .B(n21528), .Z(N28387) );
  XOR U26161 ( .A(n21518), .B(n21520), .Z(n21528) );
  XNOR U26162 ( .A(n21514), .B(n21529), .Z(n21520) );
  XNOR U26163 ( .A(n21512), .B(n21515), .Z(n21529) );
  NAND U26164 ( .A(n21530), .B(n21531), .Z(n21515) );
  NAND U26165 ( .A(n21532), .B(n21533), .Z(n21531) );
  OR U26166 ( .A(n21534), .B(n21535), .Z(n21532) );
  NANDN U26167 ( .A(n21536), .B(n21534), .Z(n21530) );
  IV U26168 ( .A(n21535), .Z(n21536) );
  NAND U26169 ( .A(n21537), .B(n21538), .Z(n21512) );
  NAND U26170 ( .A(n21539), .B(n21540), .Z(n21538) );
  NANDN U26171 ( .A(n21541), .B(n21542), .Z(n21539) );
  NANDN U26172 ( .A(n21542), .B(n21541), .Z(n21537) );
  AND U26173 ( .A(n21543), .B(n21544), .Z(n21514) );
  NAND U26174 ( .A(n21545), .B(n21546), .Z(n21544) );
  OR U26175 ( .A(n21547), .B(n21548), .Z(n21545) );
  NANDN U26176 ( .A(n21549), .B(n21547), .Z(n21543) );
  NAND U26177 ( .A(n21550), .B(n21551), .Z(n21518) );
  NANDN U26178 ( .A(n21552), .B(n21553), .Z(n21551) );
  OR U26179 ( .A(n21554), .B(n21555), .Z(n21553) );
  NANDN U26180 ( .A(n21556), .B(n21554), .Z(n21550) );
  IV U26181 ( .A(n21555), .Z(n21556) );
  XNOR U26182 ( .A(n21526), .B(n21557), .Z(n21521) );
  XNOR U26183 ( .A(n21524), .B(n21527), .Z(n21557) );
  NAND U26184 ( .A(n21558), .B(n21559), .Z(n21527) );
  NAND U26185 ( .A(n21560), .B(n21561), .Z(n21559) );
  OR U26186 ( .A(n21562), .B(n21563), .Z(n21560) );
  NANDN U26187 ( .A(n21564), .B(n21562), .Z(n21558) );
  IV U26188 ( .A(n21563), .Z(n21564) );
  NAND U26189 ( .A(n21565), .B(n21566), .Z(n21524) );
  NAND U26190 ( .A(n21567), .B(n21568), .Z(n21566) );
  NANDN U26191 ( .A(n21569), .B(n21570), .Z(n21567) );
  NANDN U26192 ( .A(n21570), .B(n21569), .Z(n21565) );
  AND U26193 ( .A(n21571), .B(n21572), .Z(n21526) );
  NAND U26194 ( .A(n21573), .B(n21574), .Z(n21572) );
  OR U26195 ( .A(n21575), .B(n21576), .Z(n21573) );
  NANDN U26196 ( .A(n21577), .B(n21575), .Z(n21571) );
  XNOR U26197 ( .A(n21552), .B(n21578), .Z(N28386) );
  XOR U26198 ( .A(n21554), .B(n21555), .Z(n21578) );
  XNOR U26199 ( .A(n21568), .B(n21579), .Z(n21555) );
  XOR U26200 ( .A(n21569), .B(n21570), .Z(n21579) );
  XOR U26201 ( .A(n21575), .B(n21580), .Z(n21570) );
  XOR U26202 ( .A(n21574), .B(n21577), .Z(n21580) );
  IV U26203 ( .A(n21576), .Z(n21577) );
  NAND U26204 ( .A(n21581), .B(n21582), .Z(n21576) );
  OR U26205 ( .A(n21583), .B(n21584), .Z(n21582) );
  OR U26206 ( .A(n21585), .B(n21586), .Z(n21581) );
  NAND U26207 ( .A(n21587), .B(n21588), .Z(n21574) );
  OR U26208 ( .A(n21589), .B(n21590), .Z(n21588) );
  OR U26209 ( .A(n21591), .B(n21592), .Z(n21587) );
  NOR U26210 ( .A(n21593), .B(n21594), .Z(n21575) );
  ANDN U26211 ( .B(n21595), .A(n21596), .Z(n21569) );
  XNOR U26212 ( .A(n21562), .B(n21597), .Z(n21568) );
  XNOR U26213 ( .A(n21561), .B(n21563), .Z(n21597) );
  NAND U26214 ( .A(n21598), .B(n21599), .Z(n21563) );
  OR U26215 ( .A(n21600), .B(n21601), .Z(n21599) );
  OR U26216 ( .A(n21602), .B(n21603), .Z(n21598) );
  NAND U26217 ( .A(n21604), .B(n21605), .Z(n21561) );
  OR U26218 ( .A(n21606), .B(n21607), .Z(n21605) );
  OR U26219 ( .A(n21608), .B(n21609), .Z(n21604) );
  ANDN U26220 ( .B(n21610), .A(n21611), .Z(n21562) );
  IV U26221 ( .A(n21612), .Z(n21610) );
  ANDN U26222 ( .B(n21613), .A(n21614), .Z(n21554) );
  XOR U26223 ( .A(n21540), .B(n21615), .Z(n21552) );
  XOR U26224 ( .A(n21541), .B(n21542), .Z(n21615) );
  XOR U26225 ( .A(n21547), .B(n21616), .Z(n21542) );
  XOR U26226 ( .A(n21546), .B(n21549), .Z(n21616) );
  IV U26227 ( .A(n21548), .Z(n21549) );
  NAND U26228 ( .A(n21617), .B(n21618), .Z(n21548) );
  OR U26229 ( .A(n21619), .B(n21620), .Z(n21618) );
  OR U26230 ( .A(n21621), .B(n21622), .Z(n21617) );
  NAND U26231 ( .A(n21623), .B(n21624), .Z(n21546) );
  OR U26232 ( .A(n21625), .B(n21626), .Z(n21624) );
  OR U26233 ( .A(n21627), .B(n21628), .Z(n21623) );
  NOR U26234 ( .A(n21629), .B(n21630), .Z(n21547) );
  ANDN U26235 ( .B(n21631), .A(n21632), .Z(n21541) );
  IV U26236 ( .A(n21633), .Z(n21631) );
  XNOR U26237 ( .A(n21534), .B(n21634), .Z(n21540) );
  XNOR U26238 ( .A(n21533), .B(n21535), .Z(n21634) );
  NAND U26239 ( .A(n21635), .B(n21636), .Z(n21535) );
  OR U26240 ( .A(n21637), .B(n21638), .Z(n21636) );
  OR U26241 ( .A(n21639), .B(n21640), .Z(n21635) );
  NAND U26242 ( .A(n21641), .B(n21642), .Z(n21533) );
  OR U26243 ( .A(n21643), .B(n21644), .Z(n21642) );
  OR U26244 ( .A(n21645), .B(n21646), .Z(n21641) );
  ANDN U26245 ( .B(n21647), .A(n21648), .Z(n21534) );
  IV U26246 ( .A(n21649), .Z(n21647) );
  XNOR U26247 ( .A(n21614), .B(n21613), .Z(N28385) );
  XOR U26248 ( .A(n21633), .B(n21632), .Z(n21613) );
  XNOR U26249 ( .A(n21648), .B(n21649), .Z(n21632) );
  XNOR U26250 ( .A(n21643), .B(n21644), .Z(n21649) );
  XNOR U26251 ( .A(n21645), .B(n21646), .Z(n21644) );
  XNOR U26252 ( .A(y[916]), .B(x[916]), .Z(n21646) );
  XNOR U26253 ( .A(y[917]), .B(x[917]), .Z(n21645) );
  XNOR U26254 ( .A(y[915]), .B(x[915]), .Z(n21643) );
  XNOR U26255 ( .A(n21637), .B(n21638), .Z(n21648) );
  XNOR U26256 ( .A(y[912]), .B(x[912]), .Z(n21638) );
  XNOR U26257 ( .A(n21639), .B(n21640), .Z(n21637) );
  XNOR U26258 ( .A(y[913]), .B(x[913]), .Z(n21640) );
  XNOR U26259 ( .A(y[914]), .B(x[914]), .Z(n21639) );
  XNOR U26260 ( .A(n21630), .B(n21629), .Z(n21633) );
  XNOR U26261 ( .A(n21625), .B(n21626), .Z(n21629) );
  XNOR U26262 ( .A(y[909]), .B(x[909]), .Z(n21626) );
  XNOR U26263 ( .A(n21627), .B(n21628), .Z(n21625) );
  XNOR U26264 ( .A(y[910]), .B(x[910]), .Z(n21628) );
  XNOR U26265 ( .A(y[911]), .B(x[911]), .Z(n21627) );
  XNOR U26266 ( .A(n21619), .B(n21620), .Z(n21630) );
  XNOR U26267 ( .A(y[906]), .B(x[906]), .Z(n21620) );
  XNOR U26268 ( .A(n21621), .B(n21622), .Z(n21619) );
  XNOR U26269 ( .A(y[907]), .B(x[907]), .Z(n21622) );
  XNOR U26270 ( .A(y[908]), .B(x[908]), .Z(n21621) );
  XOR U26271 ( .A(n21595), .B(n21596), .Z(n21614) );
  XNOR U26272 ( .A(n21611), .B(n21612), .Z(n21596) );
  XNOR U26273 ( .A(n21606), .B(n21607), .Z(n21612) );
  XNOR U26274 ( .A(n21608), .B(n21609), .Z(n21607) );
  XNOR U26275 ( .A(y[904]), .B(x[904]), .Z(n21609) );
  XNOR U26276 ( .A(y[905]), .B(x[905]), .Z(n21608) );
  XNOR U26277 ( .A(y[903]), .B(x[903]), .Z(n21606) );
  XNOR U26278 ( .A(n21600), .B(n21601), .Z(n21611) );
  XNOR U26279 ( .A(y[900]), .B(x[900]), .Z(n21601) );
  XNOR U26280 ( .A(n21602), .B(n21603), .Z(n21600) );
  XNOR U26281 ( .A(y[901]), .B(x[901]), .Z(n21603) );
  XNOR U26282 ( .A(y[902]), .B(x[902]), .Z(n21602) );
  XOR U26283 ( .A(n21594), .B(n21593), .Z(n21595) );
  XNOR U26284 ( .A(n21589), .B(n21590), .Z(n21593) );
  XNOR U26285 ( .A(y[897]), .B(x[897]), .Z(n21590) );
  XNOR U26286 ( .A(n21591), .B(n21592), .Z(n21589) );
  XNOR U26287 ( .A(y[898]), .B(x[898]), .Z(n21592) );
  XNOR U26288 ( .A(y[899]), .B(x[899]), .Z(n21591) );
  XNOR U26289 ( .A(n21583), .B(n21584), .Z(n21594) );
  XNOR U26290 ( .A(y[894]), .B(x[894]), .Z(n21584) );
  XNOR U26291 ( .A(n21585), .B(n21586), .Z(n21583) );
  XNOR U26292 ( .A(y[895]), .B(x[895]), .Z(n21586) );
  XNOR U26293 ( .A(y[896]), .B(x[896]), .Z(n21585) );
  NAND U26294 ( .A(n21650), .B(n21651), .Z(N28377) );
  NANDN U26295 ( .A(n21652), .B(n21653), .Z(n21651) );
  OR U26296 ( .A(n21654), .B(n21655), .Z(n21653) );
  NAND U26297 ( .A(n21654), .B(n21655), .Z(n21650) );
  XOR U26298 ( .A(n21654), .B(n21656), .Z(N28376) );
  XNOR U26299 ( .A(n21652), .B(n21655), .Z(n21656) );
  AND U26300 ( .A(n21657), .B(n21658), .Z(n21655) );
  NANDN U26301 ( .A(n21659), .B(n21660), .Z(n21658) );
  NANDN U26302 ( .A(n21661), .B(n21662), .Z(n21660) );
  NANDN U26303 ( .A(n21662), .B(n21661), .Z(n21657) );
  NAND U26304 ( .A(n21663), .B(n21664), .Z(n21652) );
  NANDN U26305 ( .A(n21665), .B(n21666), .Z(n21664) );
  OR U26306 ( .A(n21667), .B(n21668), .Z(n21666) );
  NAND U26307 ( .A(n21668), .B(n21667), .Z(n21663) );
  AND U26308 ( .A(n21669), .B(n21670), .Z(n21654) );
  NANDN U26309 ( .A(n21671), .B(n21672), .Z(n21670) );
  NANDN U26310 ( .A(n21673), .B(n21674), .Z(n21672) );
  NANDN U26311 ( .A(n21674), .B(n21673), .Z(n21669) );
  XOR U26312 ( .A(n21668), .B(n21675), .Z(N28375) );
  XOR U26313 ( .A(n21665), .B(n21667), .Z(n21675) );
  XNOR U26314 ( .A(n21661), .B(n21676), .Z(n21667) );
  XNOR U26315 ( .A(n21659), .B(n21662), .Z(n21676) );
  NAND U26316 ( .A(n21677), .B(n21678), .Z(n21662) );
  NAND U26317 ( .A(n21679), .B(n21680), .Z(n21678) );
  OR U26318 ( .A(n21681), .B(n21682), .Z(n21679) );
  NANDN U26319 ( .A(n21683), .B(n21681), .Z(n21677) );
  IV U26320 ( .A(n21682), .Z(n21683) );
  NAND U26321 ( .A(n21684), .B(n21685), .Z(n21659) );
  NAND U26322 ( .A(n21686), .B(n21687), .Z(n21685) );
  NANDN U26323 ( .A(n21688), .B(n21689), .Z(n21686) );
  NANDN U26324 ( .A(n21689), .B(n21688), .Z(n21684) );
  AND U26325 ( .A(n21690), .B(n21691), .Z(n21661) );
  NAND U26326 ( .A(n21692), .B(n21693), .Z(n21691) );
  OR U26327 ( .A(n21694), .B(n21695), .Z(n21692) );
  NANDN U26328 ( .A(n21696), .B(n21694), .Z(n21690) );
  NAND U26329 ( .A(n21697), .B(n21698), .Z(n21665) );
  NANDN U26330 ( .A(n21699), .B(n21700), .Z(n21698) );
  OR U26331 ( .A(n21701), .B(n21702), .Z(n21700) );
  NANDN U26332 ( .A(n21703), .B(n21701), .Z(n21697) );
  IV U26333 ( .A(n21702), .Z(n21703) );
  XNOR U26334 ( .A(n21673), .B(n21704), .Z(n21668) );
  XNOR U26335 ( .A(n21671), .B(n21674), .Z(n21704) );
  NAND U26336 ( .A(n21705), .B(n21706), .Z(n21674) );
  NAND U26337 ( .A(n21707), .B(n21708), .Z(n21706) );
  OR U26338 ( .A(n21709), .B(n21710), .Z(n21707) );
  NANDN U26339 ( .A(n21711), .B(n21709), .Z(n21705) );
  IV U26340 ( .A(n21710), .Z(n21711) );
  NAND U26341 ( .A(n21712), .B(n21713), .Z(n21671) );
  NAND U26342 ( .A(n21714), .B(n21715), .Z(n21713) );
  NANDN U26343 ( .A(n21716), .B(n21717), .Z(n21714) );
  NANDN U26344 ( .A(n21717), .B(n21716), .Z(n21712) );
  AND U26345 ( .A(n21718), .B(n21719), .Z(n21673) );
  NAND U26346 ( .A(n21720), .B(n21721), .Z(n21719) );
  OR U26347 ( .A(n21722), .B(n21723), .Z(n21720) );
  NANDN U26348 ( .A(n21724), .B(n21722), .Z(n21718) );
  XNOR U26349 ( .A(n21699), .B(n21725), .Z(N28374) );
  XOR U26350 ( .A(n21701), .B(n21702), .Z(n21725) );
  XNOR U26351 ( .A(n21715), .B(n21726), .Z(n21702) );
  XOR U26352 ( .A(n21716), .B(n21717), .Z(n21726) );
  XOR U26353 ( .A(n21722), .B(n21727), .Z(n21717) );
  XOR U26354 ( .A(n21721), .B(n21724), .Z(n21727) );
  IV U26355 ( .A(n21723), .Z(n21724) );
  NAND U26356 ( .A(n21728), .B(n21729), .Z(n21723) );
  OR U26357 ( .A(n21730), .B(n21731), .Z(n21729) );
  OR U26358 ( .A(n21732), .B(n21733), .Z(n21728) );
  NAND U26359 ( .A(n21734), .B(n21735), .Z(n21721) );
  OR U26360 ( .A(n21736), .B(n21737), .Z(n21735) );
  OR U26361 ( .A(n21738), .B(n21739), .Z(n21734) );
  NOR U26362 ( .A(n21740), .B(n21741), .Z(n21722) );
  ANDN U26363 ( .B(n21742), .A(n21743), .Z(n21716) );
  XNOR U26364 ( .A(n21709), .B(n21744), .Z(n21715) );
  XNOR U26365 ( .A(n21708), .B(n21710), .Z(n21744) );
  NAND U26366 ( .A(n21745), .B(n21746), .Z(n21710) );
  OR U26367 ( .A(n21747), .B(n21748), .Z(n21746) );
  OR U26368 ( .A(n21749), .B(n21750), .Z(n21745) );
  NAND U26369 ( .A(n21751), .B(n21752), .Z(n21708) );
  OR U26370 ( .A(n21753), .B(n21754), .Z(n21752) );
  OR U26371 ( .A(n21755), .B(n21756), .Z(n21751) );
  ANDN U26372 ( .B(n21757), .A(n21758), .Z(n21709) );
  IV U26373 ( .A(n21759), .Z(n21757) );
  ANDN U26374 ( .B(n21760), .A(n21761), .Z(n21701) );
  XOR U26375 ( .A(n21687), .B(n21762), .Z(n21699) );
  XOR U26376 ( .A(n21688), .B(n21689), .Z(n21762) );
  XOR U26377 ( .A(n21694), .B(n21763), .Z(n21689) );
  XOR U26378 ( .A(n21693), .B(n21696), .Z(n21763) );
  IV U26379 ( .A(n21695), .Z(n21696) );
  NAND U26380 ( .A(n21764), .B(n21765), .Z(n21695) );
  OR U26381 ( .A(n21766), .B(n21767), .Z(n21765) );
  OR U26382 ( .A(n21768), .B(n21769), .Z(n21764) );
  NAND U26383 ( .A(n21770), .B(n21771), .Z(n21693) );
  OR U26384 ( .A(n21772), .B(n21773), .Z(n21771) );
  OR U26385 ( .A(n21774), .B(n21775), .Z(n21770) );
  NOR U26386 ( .A(n21776), .B(n21777), .Z(n21694) );
  ANDN U26387 ( .B(n21778), .A(n21779), .Z(n21688) );
  IV U26388 ( .A(n21780), .Z(n21778) );
  XNOR U26389 ( .A(n21681), .B(n21781), .Z(n21687) );
  XNOR U26390 ( .A(n21680), .B(n21682), .Z(n21781) );
  NAND U26391 ( .A(n21782), .B(n21783), .Z(n21682) );
  OR U26392 ( .A(n21784), .B(n21785), .Z(n21783) );
  OR U26393 ( .A(n21786), .B(n21787), .Z(n21782) );
  NAND U26394 ( .A(n21788), .B(n21789), .Z(n21680) );
  OR U26395 ( .A(n21790), .B(n21791), .Z(n21789) );
  OR U26396 ( .A(n21792), .B(n21793), .Z(n21788) );
  ANDN U26397 ( .B(n21794), .A(n21795), .Z(n21681) );
  IV U26398 ( .A(n21796), .Z(n21794) );
  XNOR U26399 ( .A(n21761), .B(n21760), .Z(N28373) );
  XOR U26400 ( .A(n21780), .B(n21779), .Z(n21760) );
  XNOR U26401 ( .A(n21795), .B(n21796), .Z(n21779) );
  XNOR U26402 ( .A(n21790), .B(n21791), .Z(n21796) );
  XNOR U26403 ( .A(n21792), .B(n21793), .Z(n21791) );
  XNOR U26404 ( .A(y[892]), .B(x[892]), .Z(n21793) );
  XNOR U26405 ( .A(y[893]), .B(x[893]), .Z(n21792) );
  XNOR U26406 ( .A(y[891]), .B(x[891]), .Z(n21790) );
  XNOR U26407 ( .A(n21784), .B(n21785), .Z(n21795) );
  XNOR U26408 ( .A(y[888]), .B(x[888]), .Z(n21785) );
  XNOR U26409 ( .A(n21786), .B(n21787), .Z(n21784) );
  XNOR U26410 ( .A(y[889]), .B(x[889]), .Z(n21787) );
  XNOR U26411 ( .A(y[890]), .B(x[890]), .Z(n21786) );
  XNOR U26412 ( .A(n21777), .B(n21776), .Z(n21780) );
  XNOR U26413 ( .A(n21772), .B(n21773), .Z(n21776) );
  XNOR U26414 ( .A(y[885]), .B(x[885]), .Z(n21773) );
  XNOR U26415 ( .A(n21774), .B(n21775), .Z(n21772) );
  XNOR U26416 ( .A(y[886]), .B(x[886]), .Z(n21775) );
  XNOR U26417 ( .A(y[887]), .B(x[887]), .Z(n21774) );
  XNOR U26418 ( .A(n21766), .B(n21767), .Z(n21777) );
  XNOR U26419 ( .A(y[882]), .B(x[882]), .Z(n21767) );
  XNOR U26420 ( .A(n21768), .B(n21769), .Z(n21766) );
  XNOR U26421 ( .A(y[883]), .B(x[883]), .Z(n21769) );
  XNOR U26422 ( .A(y[884]), .B(x[884]), .Z(n21768) );
  XOR U26423 ( .A(n21742), .B(n21743), .Z(n21761) );
  XNOR U26424 ( .A(n21758), .B(n21759), .Z(n21743) );
  XNOR U26425 ( .A(n21753), .B(n21754), .Z(n21759) );
  XNOR U26426 ( .A(n21755), .B(n21756), .Z(n21754) );
  XNOR U26427 ( .A(y[880]), .B(x[880]), .Z(n21756) );
  XNOR U26428 ( .A(y[881]), .B(x[881]), .Z(n21755) );
  XNOR U26429 ( .A(y[879]), .B(x[879]), .Z(n21753) );
  XNOR U26430 ( .A(n21747), .B(n21748), .Z(n21758) );
  XNOR U26431 ( .A(y[876]), .B(x[876]), .Z(n21748) );
  XNOR U26432 ( .A(n21749), .B(n21750), .Z(n21747) );
  XNOR U26433 ( .A(y[877]), .B(x[877]), .Z(n21750) );
  XNOR U26434 ( .A(y[878]), .B(x[878]), .Z(n21749) );
  XOR U26435 ( .A(n21741), .B(n21740), .Z(n21742) );
  XNOR U26436 ( .A(n21736), .B(n21737), .Z(n21740) );
  XNOR U26437 ( .A(y[873]), .B(x[873]), .Z(n21737) );
  XNOR U26438 ( .A(n21738), .B(n21739), .Z(n21736) );
  XNOR U26439 ( .A(y[874]), .B(x[874]), .Z(n21739) );
  XNOR U26440 ( .A(y[875]), .B(x[875]), .Z(n21738) );
  XNOR U26441 ( .A(n21730), .B(n21731), .Z(n21741) );
  XNOR U26442 ( .A(y[870]), .B(x[870]), .Z(n21731) );
  XNOR U26443 ( .A(n21732), .B(n21733), .Z(n21730) );
  XNOR U26444 ( .A(y[871]), .B(x[871]), .Z(n21733) );
  XNOR U26445 ( .A(y[872]), .B(x[872]), .Z(n21732) );
  NAND U26446 ( .A(n21797), .B(n21798), .Z(N28365) );
  NANDN U26447 ( .A(n21799), .B(n21800), .Z(n21798) );
  OR U26448 ( .A(n21801), .B(n21802), .Z(n21800) );
  NAND U26449 ( .A(n21801), .B(n21802), .Z(n21797) );
  XOR U26450 ( .A(n21801), .B(n21803), .Z(N28364) );
  XNOR U26451 ( .A(n21799), .B(n21802), .Z(n21803) );
  AND U26452 ( .A(n21804), .B(n21805), .Z(n21802) );
  NANDN U26453 ( .A(n21806), .B(n21807), .Z(n21805) );
  NANDN U26454 ( .A(n21808), .B(n21809), .Z(n21807) );
  NANDN U26455 ( .A(n21809), .B(n21808), .Z(n21804) );
  NAND U26456 ( .A(n21810), .B(n21811), .Z(n21799) );
  NANDN U26457 ( .A(n21812), .B(n21813), .Z(n21811) );
  OR U26458 ( .A(n21814), .B(n21815), .Z(n21813) );
  NAND U26459 ( .A(n21815), .B(n21814), .Z(n21810) );
  AND U26460 ( .A(n21816), .B(n21817), .Z(n21801) );
  NANDN U26461 ( .A(n21818), .B(n21819), .Z(n21817) );
  NANDN U26462 ( .A(n21820), .B(n21821), .Z(n21819) );
  NANDN U26463 ( .A(n21821), .B(n21820), .Z(n21816) );
  XOR U26464 ( .A(n21815), .B(n21822), .Z(N28363) );
  XOR U26465 ( .A(n21812), .B(n21814), .Z(n21822) );
  XNOR U26466 ( .A(n21808), .B(n21823), .Z(n21814) );
  XNOR U26467 ( .A(n21806), .B(n21809), .Z(n21823) );
  NAND U26468 ( .A(n21824), .B(n21825), .Z(n21809) );
  NAND U26469 ( .A(n21826), .B(n21827), .Z(n21825) );
  OR U26470 ( .A(n21828), .B(n21829), .Z(n21826) );
  NANDN U26471 ( .A(n21830), .B(n21828), .Z(n21824) );
  IV U26472 ( .A(n21829), .Z(n21830) );
  NAND U26473 ( .A(n21831), .B(n21832), .Z(n21806) );
  NAND U26474 ( .A(n21833), .B(n21834), .Z(n21832) );
  NANDN U26475 ( .A(n21835), .B(n21836), .Z(n21833) );
  NANDN U26476 ( .A(n21836), .B(n21835), .Z(n21831) );
  AND U26477 ( .A(n21837), .B(n21838), .Z(n21808) );
  NAND U26478 ( .A(n21839), .B(n21840), .Z(n21838) );
  OR U26479 ( .A(n21841), .B(n21842), .Z(n21839) );
  NANDN U26480 ( .A(n21843), .B(n21841), .Z(n21837) );
  NAND U26481 ( .A(n21844), .B(n21845), .Z(n21812) );
  NANDN U26482 ( .A(n21846), .B(n21847), .Z(n21845) );
  OR U26483 ( .A(n21848), .B(n21849), .Z(n21847) );
  NANDN U26484 ( .A(n21850), .B(n21848), .Z(n21844) );
  IV U26485 ( .A(n21849), .Z(n21850) );
  XNOR U26486 ( .A(n21820), .B(n21851), .Z(n21815) );
  XNOR U26487 ( .A(n21818), .B(n21821), .Z(n21851) );
  NAND U26488 ( .A(n21852), .B(n21853), .Z(n21821) );
  NAND U26489 ( .A(n21854), .B(n21855), .Z(n21853) );
  OR U26490 ( .A(n21856), .B(n21857), .Z(n21854) );
  NANDN U26491 ( .A(n21858), .B(n21856), .Z(n21852) );
  IV U26492 ( .A(n21857), .Z(n21858) );
  NAND U26493 ( .A(n21859), .B(n21860), .Z(n21818) );
  NAND U26494 ( .A(n21861), .B(n21862), .Z(n21860) );
  NANDN U26495 ( .A(n21863), .B(n21864), .Z(n21861) );
  NANDN U26496 ( .A(n21864), .B(n21863), .Z(n21859) );
  AND U26497 ( .A(n21865), .B(n21866), .Z(n21820) );
  NAND U26498 ( .A(n21867), .B(n21868), .Z(n21866) );
  OR U26499 ( .A(n21869), .B(n21870), .Z(n21867) );
  NANDN U26500 ( .A(n21871), .B(n21869), .Z(n21865) );
  XNOR U26501 ( .A(n21846), .B(n21872), .Z(N28362) );
  XOR U26502 ( .A(n21848), .B(n21849), .Z(n21872) );
  XNOR U26503 ( .A(n21862), .B(n21873), .Z(n21849) );
  XOR U26504 ( .A(n21863), .B(n21864), .Z(n21873) );
  XOR U26505 ( .A(n21869), .B(n21874), .Z(n21864) );
  XOR U26506 ( .A(n21868), .B(n21871), .Z(n21874) );
  IV U26507 ( .A(n21870), .Z(n21871) );
  NAND U26508 ( .A(n21875), .B(n21876), .Z(n21870) );
  OR U26509 ( .A(n21877), .B(n21878), .Z(n21876) );
  OR U26510 ( .A(n21879), .B(n21880), .Z(n21875) );
  NAND U26511 ( .A(n21881), .B(n21882), .Z(n21868) );
  OR U26512 ( .A(n21883), .B(n21884), .Z(n21882) );
  OR U26513 ( .A(n21885), .B(n21886), .Z(n21881) );
  NOR U26514 ( .A(n21887), .B(n21888), .Z(n21869) );
  ANDN U26515 ( .B(n21889), .A(n21890), .Z(n21863) );
  XNOR U26516 ( .A(n21856), .B(n21891), .Z(n21862) );
  XNOR U26517 ( .A(n21855), .B(n21857), .Z(n21891) );
  NAND U26518 ( .A(n21892), .B(n21893), .Z(n21857) );
  OR U26519 ( .A(n21894), .B(n21895), .Z(n21893) );
  OR U26520 ( .A(n21896), .B(n21897), .Z(n21892) );
  NAND U26521 ( .A(n21898), .B(n21899), .Z(n21855) );
  OR U26522 ( .A(n21900), .B(n21901), .Z(n21899) );
  OR U26523 ( .A(n21902), .B(n21903), .Z(n21898) );
  ANDN U26524 ( .B(n21904), .A(n21905), .Z(n21856) );
  IV U26525 ( .A(n21906), .Z(n21904) );
  ANDN U26526 ( .B(n21907), .A(n21908), .Z(n21848) );
  XOR U26527 ( .A(n21834), .B(n21909), .Z(n21846) );
  XOR U26528 ( .A(n21835), .B(n21836), .Z(n21909) );
  XOR U26529 ( .A(n21841), .B(n21910), .Z(n21836) );
  XOR U26530 ( .A(n21840), .B(n21843), .Z(n21910) );
  IV U26531 ( .A(n21842), .Z(n21843) );
  NAND U26532 ( .A(n21911), .B(n21912), .Z(n21842) );
  OR U26533 ( .A(n21913), .B(n21914), .Z(n21912) );
  OR U26534 ( .A(n21915), .B(n21916), .Z(n21911) );
  NAND U26535 ( .A(n21917), .B(n21918), .Z(n21840) );
  OR U26536 ( .A(n21919), .B(n21920), .Z(n21918) );
  OR U26537 ( .A(n21921), .B(n21922), .Z(n21917) );
  NOR U26538 ( .A(n21923), .B(n21924), .Z(n21841) );
  ANDN U26539 ( .B(n21925), .A(n21926), .Z(n21835) );
  IV U26540 ( .A(n21927), .Z(n21925) );
  XNOR U26541 ( .A(n21828), .B(n21928), .Z(n21834) );
  XNOR U26542 ( .A(n21827), .B(n21829), .Z(n21928) );
  NAND U26543 ( .A(n21929), .B(n21930), .Z(n21829) );
  OR U26544 ( .A(n21931), .B(n21932), .Z(n21930) );
  OR U26545 ( .A(n21933), .B(n21934), .Z(n21929) );
  NAND U26546 ( .A(n21935), .B(n21936), .Z(n21827) );
  OR U26547 ( .A(n21937), .B(n21938), .Z(n21936) );
  OR U26548 ( .A(n21939), .B(n21940), .Z(n21935) );
  ANDN U26549 ( .B(n21941), .A(n21942), .Z(n21828) );
  IV U26550 ( .A(n21943), .Z(n21941) );
  XNOR U26551 ( .A(n21908), .B(n21907), .Z(N28361) );
  XOR U26552 ( .A(n21927), .B(n21926), .Z(n21907) );
  XNOR U26553 ( .A(n21942), .B(n21943), .Z(n21926) );
  XNOR U26554 ( .A(n21937), .B(n21938), .Z(n21943) );
  XNOR U26555 ( .A(n21939), .B(n21940), .Z(n21938) );
  XNOR U26556 ( .A(y[868]), .B(x[868]), .Z(n21940) );
  XNOR U26557 ( .A(y[869]), .B(x[869]), .Z(n21939) );
  XNOR U26558 ( .A(y[867]), .B(x[867]), .Z(n21937) );
  XNOR U26559 ( .A(n21931), .B(n21932), .Z(n21942) );
  XNOR U26560 ( .A(y[864]), .B(x[864]), .Z(n21932) );
  XNOR U26561 ( .A(n21933), .B(n21934), .Z(n21931) );
  XNOR U26562 ( .A(y[865]), .B(x[865]), .Z(n21934) );
  XNOR U26563 ( .A(y[866]), .B(x[866]), .Z(n21933) );
  XNOR U26564 ( .A(n21924), .B(n21923), .Z(n21927) );
  XNOR U26565 ( .A(n21919), .B(n21920), .Z(n21923) );
  XNOR U26566 ( .A(y[861]), .B(x[861]), .Z(n21920) );
  XNOR U26567 ( .A(n21921), .B(n21922), .Z(n21919) );
  XNOR U26568 ( .A(y[862]), .B(x[862]), .Z(n21922) );
  XNOR U26569 ( .A(y[863]), .B(x[863]), .Z(n21921) );
  XNOR U26570 ( .A(n21913), .B(n21914), .Z(n21924) );
  XNOR U26571 ( .A(y[858]), .B(x[858]), .Z(n21914) );
  XNOR U26572 ( .A(n21915), .B(n21916), .Z(n21913) );
  XNOR U26573 ( .A(y[859]), .B(x[859]), .Z(n21916) );
  XNOR U26574 ( .A(y[860]), .B(x[860]), .Z(n21915) );
  XOR U26575 ( .A(n21889), .B(n21890), .Z(n21908) );
  XNOR U26576 ( .A(n21905), .B(n21906), .Z(n21890) );
  XNOR U26577 ( .A(n21900), .B(n21901), .Z(n21906) );
  XNOR U26578 ( .A(n21902), .B(n21903), .Z(n21901) );
  XNOR U26579 ( .A(y[856]), .B(x[856]), .Z(n21903) );
  XNOR U26580 ( .A(y[857]), .B(x[857]), .Z(n21902) );
  XNOR U26581 ( .A(y[855]), .B(x[855]), .Z(n21900) );
  XNOR U26582 ( .A(n21894), .B(n21895), .Z(n21905) );
  XNOR U26583 ( .A(y[852]), .B(x[852]), .Z(n21895) );
  XNOR U26584 ( .A(n21896), .B(n21897), .Z(n21894) );
  XNOR U26585 ( .A(y[853]), .B(x[853]), .Z(n21897) );
  XNOR U26586 ( .A(y[854]), .B(x[854]), .Z(n21896) );
  XOR U26587 ( .A(n21888), .B(n21887), .Z(n21889) );
  XNOR U26588 ( .A(n21883), .B(n21884), .Z(n21887) );
  XNOR U26589 ( .A(y[849]), .B(x[849]), .Z(n21884) );
  XNOR U26590 ( .A(n21885), .B(n21886), .Z(n21883) );
  XNOR U26591 ( .A(y[850]), .B(x[850]), .Z(n21886) );
  XNOR U26592 ( .A(y[851]), .B(x[851]), .Z(n21885) );
  XNOR U26593 ( .A(n21877), .B(n21878), .Z(n21888) );
  XNOR U26594 ( .A(y[846]), .B(x[846]), .Z(n21878) );
  XNOR U26595 ( .A(n21879), .B(n21880), .Z(n21877) );
  XNOR U26596 ( .A(y[847]), .B(x[847]), .Z(n21880) );
  XNOR U26597 ( .A(y[848]), .B(x[848]), .Z(n21879) );
  NAND U26598 ( .A(n21944), .B(n21945), .Z(N28353) );
  NANDN U26599 ( .A(n21946), .B(n21947), .Z(n21945) );
  OR U26600 ( .A(n21948), .B(n21949), .Z(n21947) );
  NAND U26601 ( .A(n21948), .B(n21949), .Z(n21944) );
  XOR U26602 ( .A(n21948), .B(n21950), .Z(N28352) );
  XNOR U26603 ( .A(n21946), .B(n21949), .Z(n21950) );
  AND U26604 ( .A(n21951), .B(n21952), .Z(n21949) );
  NANDN U26605 ( .A(n21953), .B(n21954), .Z(n21952) );
  NANDN U26606 ( .A(n21955), .B(n21956), .Z(n21954) );
  NANDN U26607 ( .A(n21956), .B(n21955), .Z(n21951) );
  NAND U26608 ( .A(n21957), .B(n21958), .Z(n21946) );
  NANDN U26609 ( .A(n21959), .B(n21960), .Z(n21958) );
  OR U26610 ( .A(n21961), .B(n21962), .Z(n21960) );
  NAND U26611 ( .A(n21962), .B(n21961), .Z(n21957) );
  AND U26612 ( .A(n21963), .B(n21964), .Z(n21948) );
  NANDN U26613 ( .A(n21965), .B(n21966), .Z(n21964) );
  NANDN U26614 ( .A(n21967), .B(n21968), .Z(n21966) );
  NANDN U26615 ( .A(n21968), .B(n21967), .Z(n21963) );
  XOR U26616 ( .A(n21962), .B(n21969), .Z(N28351) );
  XOR U26617 ( .A(n21959), .B(n21961), .Z(n21969) );
  XNOR U26618 ( .A(n21955), .B(n21970), .Z(n21961) );
  XNOR U26619 ( .A(n21953), .B(n21956), .Z(n21970) );
  NAND U26620 ( .A(n21971), .B(n21972), .Z(n21956) );
  NAND U26621 ( .A(n21973), .B(n21974), .Z(n21972) );
  OR U26622 ( .A(n21975), .B(n21976), .Z(n21973) );
  NANDN U26623 ( .A(n21977), .B(n21975), .Z(n21971) );
  IV U26624 ( .A(n21976), .Z(n21977) );
  NAND U26625 ( .A(n21978), .B(n21979), .Z(n21953) );
  NAND U26626 ( .A(n21980), .B(n21981), .Z(n21979) );
  NANDN U26627 ( .A(n21982), .B(n21983), .Z(n21980) );
  NANDN U26628 ( .A(n21983), .B(n21982), .Z(n21978) );
  AND U26629 ( .A(n21984), .B(n21985), .Z(n21955) );
  NAND U26630 ( .A(n21986), .B(n21987), .Z(n21985) );
  OR U26631 ( .A(n21988), .B(n21989), .Z(n21986) );
  NANDN U26632 ( .A(n21990), .B(n21988), .Z(n21984) );
  NAND U26633 ( .A(n21991), .B(n21992), .Z(n21959) );
  NANDN U26634 ( .A(n21993), .B(n21994), .Z(n21992) );
  OR U26635 ( .A(n21995), .B(n21996), .Z(n21994) );
  NANDN U26636 ( .A(n21997), .B(n21995), .Z(n21991) );
  IV U26637 ( .A(n21996), .Z(n21997) );
  XNOR U26638 ( .A(n21967), .B(n21998), .Z(n21962) );
  XNOR U26639 ( .A(n21965), .B(n21968), .Z(n21998) );
  NAND U26640 ( .A(n21999), .B(n22000), .Z(n21968) );
  NAND U26641 ( .A(n22001), .B(n22002), .Z(n22000) );
  OR U26642 ( .A(n22003), .B(n22004), .Z(n22001) );
  NANDN U26643 ( .A(n22005), .B(n22003), .Z(n21999) );
  IV U26644 ( .A(n22004), .Z(n22005) );
  NAND U26645 ( .A(n22006), .B(n22007), .Z(n21965) );
  NAND U26646 ( .A(n22008), .B(n22009), .Z(n22007) );
  NANDN U26647 ( .A(n22010), .B(n22011), .Z(n22008) );
  NANDN U26648 ( .A(n22011), .B(n22010), .Z(n22006) );
  AND U26649 ( .A(n22012), .B(n22013), .Z(n21967) );
  NAND U26650 ( .A(n22014), .B(n22015), .Z(n22013) );
  OR U26651 ( .A(n22016), .B(n22017), .Z(n22014) );
  NANDN U26652 ( .A(n22018), .B(n22016), .Z(n22012) );
  XNOR U26653 ( .A(n21993), .B(n22019), .Z(N28350) );
  XOR U26654 ( .A(n21995), .B(n21996), .Z(n22019) );
  XNOR U26655 ( .A(n22009), .B(n22020), .Z(n21996) );
  XOR U26656 ( .A(n22010), .B(n22011), .Z(n22020) );
  XOR U26657 ( .A(n22016), .B(n22021), .Z(n22011) );
  XOR U26658 ( .A(n22015), .B(n22018), .Z(n22021) );
  IV U26659 ( .A(n22017), .Z(n22018) );
  NAND U26660 ( .A(n22022), .B(n22023), .Z(n22017) );
  OR U26661 ( .A(n22024), .B(n22025), .Z(n22023) );
  OR U26662 ( .A(n22026), .B(n22027), .Z(n22022) );
  NAND U26663 ( .A(n22028), .B(n22029), .Z(n22015) );
  OR U26664 ( .A(n22030), .B(n22031), .Z(n22029) );
  OR U26665 ( .A(n22032), .B(n22033), .Z(n22028) );
  NOR U26666 ( .A(n22034), .B(n22035), .Z(n22016) );
  ANDN U26667 ( .B(n22036), .A(n22037), .Z(n22010) );
  XNOR U26668 ( .A(n22003), .B(n22038), .Z(n22009) );
  XNOR U26669 ( .A(n22002), .B(n22004), .Z(n22038) );
  NAND U26670 ( .A(n22039), .B(n22040), .Z(n22004) );
  OR U26671 ( .A(n22041), .B(n22042), .Z(n22040) );
  OR U26672 ( .A(n22043), .B(n22044), .Z(n22039) );
  NAND U26673 ( .A(n22045), .B(n22046), .Z(n22002) );
  OR U26674 ( .A(n22047), .B(n22048), .Z(n22046) );
  OR U26675 ( .A(n22049), .B(n22050), .Z(n22045) );
  ANDN U26676 ( .B(n22051), .A(n22052), .Z(n22003) );
  IV U26677 ( .A(n22053), .Z(n22051) );
  ANDN U26678 ( .B(n22054), .A(n22055), .Z(n21995) );
  XOR U26679 ( .A(n21981), .B(n22056), .Z(n21993) );
  XOR U26680 ( .A(n21982), .B(n21983), .Z(n22056) );
  XOR U26681 ( .A(n21988), .B(n22057), .Z(n21983) );
  XOR U26682 ( .A(n21987), .B(n21990), .Z(n22057) );
  IV U26683 ( .A(n21989), .Z(n21990) );
  NAND U26684 ( .A(n22058), .B(n22059), .Z(n21989) );
  OR U26685 ( .A(n22060), .B(n22061), .Z(n22059) );
  OR U26686 ( .A(n22062), .B(n22063), .Z(n22058) );
  NAND U26687 ( .A(n22064), .B(n22065), .Z(n21987) );
  OR U26688 ( .A(n22066), .B(n22067), .Z(n22065) );
  OR U26689 ( .A(n22068), .B(n22069), .Z(n22064) );
  NOR U26690 ( .A(n22070), .B(n22071), .Z(n21988) );
  ANDN U26691 ( .B(n22072), .A(n22073), .Z(n21982) );
  IV U26692 ( .A(n22074), .Z(n22072) );
  XNOR U26693 ( .A(n21975), .B(n22075), .Z(n21981) );
  XNOR U26694 ( .A(n21974), .B(n21976), .Z(n22075) );
  NAND U26695 ( .A(n22076), .B(n22077), .Z(n21976) );
  OR U26696 ( .A(n22078), .B(n22079), .Z(n22077) );
  OR U26697 ( .A(n22080), .B(n22081), .Z(n22076) );
  NAND U26698 ( .A(n22082), .B(n22083), .Z(n21974) );
  OR U26699 ( .A(n22084), .B(n22085), .Z(n22083) );
  OR U26700 ( .A(n22086), .B(n22087), .Z(n22082) );
  ANDN U26701 ( .B(n22088), .A(n22089), .Z(n21975) );
  IV U26702 ( .A(n22090), .Z(n22088) );
  XNOR U26703 ( .A(n22055), .B(n22054), .Z(N28349) );
  XOR U26704 ( .A(n22074), .B(n22073), .Z(n22054) );
  XNOR U26705 ( .A(n22089), .B(n22090), .Z(n22073) );
  XNOR U26706 ( .A(n22084), .B(n22085), .Z(n22090) );
  XNOR U26707 ( .A(n22086), .B(n22087), .Z(n22085) );
  XNOR U26708 ( .A(y[844]), .B(x[844]), .Z(n22087) );
  XNOR U26709 ( .A(y[845]), .B(x[845]), .Z(n22086) );
  XNOR U26710 ( .A(y[843]), .B(x[843]), .Z(n22084) );
  XNOR U26711 ( .A(n22078), .B(n22079), .Z(n22089) );
  XNOR U26712 ( .A(y[840]), .B(x[840]), .Z(n22079) );
  XNOR U26713 ( .A(n22080), .B(n22081), .Z(n22078) );
  XNOR U26714 ( .A(y[841]), .B(x[841]), .Z(n22081) );
  XNOR U26715 ( .A(y[842]), .B(x[842]), .Z(n22080) );
  XNOR U26716 ( .A(n22071), .B(n22070), .Z(n22074) );
  XNOR U26717 ( .A(n22066), .B(n22067), .Z(n22070) );
  XNOR U26718 ( .A(y[837]), .B(x[837]), .Z(n22067) );
  XNOR U26719 ( .A(n22068), .B(n22069), .Z(n22066) );
  XNOR U26720 ( .A(y[838]), .B(x[838]), .Z(n22069) );
  XNOR U26721 ( .A(y[839]), .B(x[839]), .Z(n22068) );
  XNOR U26722 ( .A(n22060), .B(n22061), .Z(n22071) );
  XNOR U26723 ( .A(y[834]), .B(x[834]), .Z(n22061) );
  XNOR U26724 ( .A(n22062), .B(n22063), .Z(n22060) );
  XNOR U26725 ( .A(y[835]), .B(x[835]), .Z(n22063) );
  XNOR U26726 ( .A(y[836]), .B(x[836]), .Z(n22062) );
  XOR U26727 ( .A(n22036), .B(n22037), .Z(n22055) );
  XNOR U26728 ( .A(n22052), .B(n22053), .Z(n22037) );
  XNOR U26729 ( .A(n22047), .B(n22048), .Z(n22053) );
  XNOR U26730 ( .A(n22049), .B(n22050), .Z(n22048) );
  XNOR U26731 ( .A(y[832]), .B(x[832]), .Z(n22050) );
  XNOR U26732 ( .A(y[833]), .B(x[833]), .Z(n22049) );
  XNOR U26733 ( .A(y[831]), .B(x[831]), .Z(n22047) );
  XNOR U26734 ( .A(n22041), .B(n22042), .Z(n22052) );
  XNOR U26735 ( .A(y[828]), .B(x[828]), .Z(n22042) );
  XNOR U26736 ( .A(n22043), .B(n22044), .Z(n22041) );
  XNOR U26737 ( .A(y[829]), .B(x[829]), .Z(n22044) );
  XNOR U26738 ( .A(y[830]), .B(x[830]), .Z(n22043) );
  XOR U26739 ( .A(n22035), .B(n22034), .Z(n22036) );
  XNOR U26740 ( .A(n22030), .B(n22031), .Z(n22034) );
  XNOR U26741 ( .A(y[825]), .B(x[825]), .Z(n22031) );
  XNOR U26742 ( .A(n22032), .B(n22033), .Z(n22030) );
  XNOR U26743 ( .A(y[826]), .B(x[826]), .Z(n22033) );
  XNOR U26744 ( .A(y[827]), .B(x[827]), .Z(n22032) );
  XNOR U26745 ( .A(n22024), .B(n22025), .Z(n22035) );
  XNOR U26746 ( .A(y[822]), .B(x[822]), .Z(n22025) );
  XNOR U26747 ( .A(n22026), .B(n22027), .Z(n22024) );
  XNOR U26748 ( .A(y[823]), .B(x[823]), .Z(n22027) );
  XNOR U26749 ( .A(y[824]), .B(x[824]), .Z(n22026) );
  NAND U26750 ( .A(n22091), .B(n22092), .Z(N28341) );
  NANDN U26751 ( .A(n22093), .B(n22094), .Z(n22092) );
  OR U26752 ( .A(n22095), .B(n22096), .Z(n22094) );
  NAND U26753 ( .A(n22095), .B(n22096), .Z(n22091) );
  XOR U26754 ( .A(n22095), .B(n22097), .Z(N28340) );
  XNOR U26755 ( .A(n22093), .B(n22096), .Z(n22097) );
  AND U26756 ( .A(n22098), .B(n22099), .Z(n22096) );
  NANDN U26757 ( .A(n22100), .B(n22101), .Z(n22099) );
  NANDN U26758 ( .A(n22102), .B(n22103), .Z(n22101) );
  NANDN U26759 ( .A(n22103), .B(n22102), .Z(n22098) );
  NAND U26760 ( .A(n22104), .B(n22105), .Z(n22093) );
  NANDN U26761 ( .A(n22106), .B(n22107), .Z(n22105) );
  OR U26762 ( .A(n22108), .B(n22109), .Z(n22107) );
  NAND U26763 ( .A(n22109), .B(n22108), .Z(n22104) );
  AND U26764 ( .A(n22110), .B(n22111), .Z(n22095) );
  NANDN U26765 ( .A(n22112), .B(n22113), .Z(n22111) );
  NANDN U26766 ( .A(n22114), .B(n22115), .Z(n22113) );
  NANDN U26767 ( .A(n22115), .B(n22114), .Z(n22110) );
  XOR U26768 ( .A(n22109), .B(n22116), .Z(N28339) );
  XOR U26769 ( .A(n22106), .B(n22108), .Z(n22116) );
  XNOR U26770 ( .A(n22102), .B(n22117), .Z(n22108) );
  XNOR U26771 ( .A(n22100), .B(n22103), .Z(n22117) );
  NAND U26772 ( .A(n22118), .B(n22119), .Z(n22103) );
  NAND U26773 ( .A(n22120), .B(n22121), .Z(n22119) );
  OR U26774 ( .A(n22122), .B(n22123), .Z(n22120) );
  NANDN U26775 ( .A(n22124), .B(n22122), .Z(n22118) );
  IV U26776 ( .A(n22123), .Z(n22124) );
  NAND U26777 ( .A(n22125), .B(n22126), .Z(n22100) );
  NAND U26778 ( .A(n22127), .B(n22128), .Z(n22126) );
  NANDN U26779 ( .A(n22129), .B(n22130), .Z(n22127) );
  NANDN U26780 ( .A(n22130), .B(n22129), .Z(n22125) );
  AND U26781 ( .A(n22131), .B(n22132), .Z(n22102) );
  NAND U26782 ( .A(n22133), .B(n22134), .Z(n22132) );
  OR U26783 ( .A(n22135), .B(n22136), .Z(n22133) );
  NANDN U26784 ( .A(n22137), .B(n22135), .Z(n22131) );
  NAND U26785 ( .A(n22138), .B(n22139), .Z(n22106) );
  NANDN U26786 ( .A(n22140), .B(n22141), .Z(n22139) );
  OR U26787 ( .A(n22142), .B(n22143), .Z(n22141) );
  NANDN U26788 ( .A(n22144), .B(n22142), .Z(n22138) );
  IV U26789 ( .A(n22143), .Z(n22144) );
  XNOR U26790 ( .A(n22114), .B(n22145), .Z(n22109) );
  XNOR U26791 ( .A(n22112), .B(n22115), .Z(n22145) );
  NAND U26792 ( .A(n22146), .B(n22147), .Z(n22115) );
  NAND U26793 ( .A(n22148), .B(n22149), .Z(n22147) );
  OR U26794 ( .A(n22150), .B(n22151), .Z(n22148) );
  NANDN U26795 ( .A(n22152), .B(n22150), .Z(n22146) );
  IV U26796 ( .A(n22151), .Z(n22152) );
  NAND U26797 ( .A(n22153), .B(n22154), .Z(n22112) );
  NAND U26798 ( .A(n22155), .B(n22156), .Z(n22154) );
  NANDN U26799 ( .A(n22157), .B(n22158), .Z(n22155) );
  NANDN U26800 ( .A(n22158), .B(n22157), .Z(n22153) );
  AND U26801 ( .A(n22159), .B(n22160), .Z(n22114) );
  NAND U26802 ( .A(n22161), .B(n22162), .Z(n22160) );
  OR U26803 ( .A(n22163), .B(n22164), .Z(n22161) );
  NANDN U26804 ( .A(n22165), .B(n22163), .Z(n22159) );
  XNOR U26805 ( .A(n22140), .B(n22166), .Z(N28338) );
  XOR U26806 ( .A(n22142), .B(n22143), .Z(n22166) );
  XNOR U26807 ( .A(n22156), .B(n22167), .Z(n22143) );
  XOR U26808 ( .A(n22157), .B(n22158), .Z(n22167) );
  XOR U26809 ( .A(n22163), .B(n22168), .Z(n22158) );
  XOR U26810 ( .A(n22162), .B(n22165), .Z(n22168) );
  IV U26811 ( .A(n22164), .Z(n22165) );
  NAND U26812 ( .A(n22169), .B(n22170), .Z(n22164) );
  OR U26813 ( .A(n22171), .B(n22172), .Z(n22170) );
  OR U26814 ( .A(n22173), .B(n22174), .Z(n22169) );
  NAND U26815 ( .A(n22175), .B(n22176), .Z(n22162) );
  OR U26816 ( .A(n22177), .B(n22178), .Z(n22176) );
  OR U26817 ( .A(n22179), .B(n22180), .Z(n22175) );
  NOR U26818 ( .A(n22181), .B(n22182), .Z(n22163) );
  ANDN U26819 ( .B(n22183), .A(n22184), .Z(n22157) );
  XNOR U26820 ( .A(n22150), .B(n22185), .Z(n22156) );
  XNOR U26821 ( .A(n22149), .B(n22151), .Z(n22185) );
  NAND U26822 ( .A(n22186), .B(n22187), .Z(n22151) );
  OR U26823 ( .A(n22188), .B(n22189), .Z(n22187) );
  OR U26824 ( .A(n22190), .B(n22191), .Z(n22186) );
  NAND U26825 ( .A(n22192), .B(n22193), .Z(n22149) );
  OR U26826 ( .A(n22194), .B(n22195), .Z(n22193) );
  OR U26827 ( .A(n22196), .B(n22197), .Z(n22192) );
  ANDN U26828 ( .B(n22198), .A(n22199), .Z(n22150) );
  IV U26829 ( .A(n22200), .Z(n22198) );
  ANDN U26830 ( .B(n22201), .A(n22202), .Z(n22142) );
  XOR U26831 ( .A(n22128), .B(n22203), .Z(n22140) );
  XOR U26832 ( .A(n22129), .B(n22130), .Z(n22203) );
  XOR U26833 ( .A(n22135), .B(n22204), .Z(n22130) );
  XOR U26834 ( .A(n22134), .B(n22137), .Z(n22204) );
  IV U26835 ( .A(n22136), .Z(n22137) );
  NAND U26836 ( .A(n22205), .B(n22206), .Z(n22136) );
  OR U26837 ( .A(n22207), .B(n22208), .Z(n22206) );
  OR U26838 ( .A(n22209), .B(n22210), .Z(n22205) );
  NAND U26839 ( .A(n22211), .B(n22212), .Z(n22134) );
  OR U26840 ( .A(n22213), .B(n22214), .Z(n22212) );
  OR U26841 ( .A(n22215), .B(n22216), .Z(n22211) );
  NOR U26842 ( .A(n22217), .B(n22218), .Z(n22135) );
  ANDN U26843 ( .B(n22219), .A(n22220), .Z(n22129) );
  IV U26844 ( .A(n22221), .Z(n22219) );
  XNOR U26845 ( .A(n22122), .B(n22222), .Z(n22128) );
  XNOR U26846 ( .A(n22121), .B(n22123), .Z(n22222) );
  NAND U26847 ( .A(n22223), .B(n22224), .Z(n22123) );
  OR U26848 ( .A(n22225), .B(n22226), .Z(n22224) );
  OR U26849 ( .A(n22227), .B(n22228), .Z(n22223) );
  NAND U26850 ( .A(n22229), .B(n22230), .Z(n22121) );
  OR U26851 ( .A(n22231), .B(n22232), .Z(n22230) );
  OR U26852 ( .A(n22233), .B(n22234), .Z(n22229) );
  ANDN U26853 ( .B(n22235), .A(n22236), .Z(n22122) );
  IV U26854 ( .A(n22237), .Z(n22235) );
  XNOR U26855 ( .A(n22202), .B(n22201), .Z(N28337) );
  XOR U26856 ( .A(n22221), .B(n22220), .Z(n22201) );
  XNOR U26857 ( .A(n22236), .B(n22237), .Z(n22220) );
  XNOR U26858 ( .A(n22231), .B(n22232), .Z(n22237) );
  XNOR U26859 ( .A(n22233), .B(n22234), .Z(n22232) );
  XNOR U26860 ( .A(y[820]), .B(x[820]), .Z(n22234) );
  XNOR U26861 ( .A(y[821]), .B(x[821]), .Z(n22233) );
  XNOR U26862 ( .A(y[819]), .B(x[819]), .Z(n22231) );
  XNOR U26863 ( .A(n22225), .B(n22226), .Z(n22236) );
  XNOR U26864 ( .A(y[816]), .B(x[816]), .Z(n22226) );
  XNOR U26865 ( .A(n22227), .B(n22228), .Z(n22225) );
  XNOR U26866 ( .A(y[817]), .B(x[817]), .Z(n22228) );
  XNOR U26867 ( .A(y[818]), .B(x[818]), .Z(n22227) );
  XNOR U26868 ( .A(n22218), .B(n22217), .Z(n22221) );
  XNOR U26869 ( .A(n22213), .B(n22214), .Z(n22217) );
  XNOR U26870 ( .A(y[813]), .B(x[813]), .Z(n22214) );
  XNOR U26871 ( .A(n22215), .B(n22216), .Z(n22213) );
  XNOR U26872 ( .A(y[814]), .B(x[814]), .Z(n22216) );
  XNOR U26873 ( .A(y[815]), .B(x[815]), .Z(n22215) );
  XNOR U26874 ( .A(n22207), .B(n22208), .Z(n22218) );
  XNOR U26875 ( .A(y[810]), .B(x[810]), .Z(n22208) );
  XNOR U26876 ( .A(n22209), .B(n22210), .Z(n22207) );
  XNOR U26877 ( .A(y[811]), .B(x[811]), .Z(n22210) );
  XNOR U26878 ( .A(y[812]), .B(x[812]), .Z(n22209) );
  XOR U26879 ( .A(n22183), .B(n22184), .Z(n22202) );
  XNOR U26880 ( .A(n22199), .B(n22200), .Z(n22184) );
  XNOR U26881 ( .A(n22194), .B(n22195), .Z(n22200) );
  XNOR U26882 ( .A(n22196), .B(n22197), .Z(n22195) );
  XNOR U26883 ( .A(y[808]), .B(x[808]), .Z(n22197) );
  XNOR U26884 ( .A(y[809]), .B(x[809]), .Z(n22196) );
  XNOR U26885 ( .A(y[807]), .B(x[807]), .Z(n22194) );
  XNOR U26886 ( .A(n22188), .B(n22189), .Z(n22199) );
  XNOR U26887 ( .A(y[804]), .B(x[804]), .Z(n22189) );
  XNOR U26888 ( .A(n22190), .B(n22191), .Z(n22188) );
  XNOR U26889 ( .A(y[805]), .B(x[805]), .Z(n22191) );
  XNOR U26890 ( .A(y[806]), .B(x[806]), .Z(n22190) );
  XOR U26891 ( .A(n22182), .B(n22181), .Z(n22183) );
  XNOR U26892 ( .A(n22177), .B(n22178), .Z(n22181) );
  XNOR U26893 ( .A(y[801]), .B(x[801]), .Z(n22178) );
  XNOR U26894 ( .A(n22179), .B(n22180), .Z(n22177) );
  XNOR U26895 ( .A(y[802]), .B(x[802]), .Z(n22180) );
  XNOR U26896 ( .A(y[803]), .B(x[803]), .Z(n22179) );
  XNOR U26897 ( .A(n22171), .B(n22172), .Z(n22182) );
  XNOR U26898 ( .A(y[798]), .B(x[798]), .Z(n22172) );
  XNOR U26899 ( .A(n22173), .B(n22174), .Z(n22171) );
  XNOR U26900 ( .A(y[799]), .B(x[799]), .Z(n22174) );
  XNOR U26901 ( .A(y[800]), .B(x[800]), .Z(n22173) );
  NAND U26902 ( .A(n22238), .B(n22239), .Z(N28329) );
  NANDN U26903 ( .A(n22240), .B(n22241), .Z(n22239) );
  OR U26904 ( .A(n22242), .B(n22243), .Z(n22241) );
  NAND U26905 ( .A(n22242), .B(n22243), .Z(n22238) );
  XOR U26906 ( .A(n22242), .B(n22244), .Z(N28328) );
  XNOR U26907 ( .A(n22240), .B(n22243), .Z(n22244) );
  AND U26908 ( .A(n22245), .B(n22246), .Z(n22243) );
  NANDN U26909 ( .A(n22247), .B(n22248), .Z(n22246) );
  NANDN U26910 ( .A(n22249), .B(n22250), .Z(n22248) );
  NANDN U26911 ( .A(n22250), .B(n22249), .Z(n22245) );
  NAND U26912 ( .A(n22251), .B(n22252), .Z(n22240) );
  NANDN U26913 ( .A(n22253), .B(n22254), .Z(n22252) );
  OR U26914 ( .A(n22255), .B(n22256), .Z(n22254) );
  NAND U26915 ( .A(n22256), .B(n22255), .Z(n22251) );
  AND U26916 ( .A(n22257), .B(n22258), .Z(n22242) );
  NANDN U26917 ( .A(n22259), .B(n22260), .Z(n22258) );
  NANDN U26918 ( .A(n22261), .B(n22262), .Z(n22260) );
  NANDN U26919 ( .A(n22262), .B(n22261), .Z(n22257) );
  XOR U26920 ( .A(n22256), .B(n22263), .Z(N28327) );
  XOR U26921 ( .A(n22253), .B(n22255), .Z(n22263) );
  XNOR U26922 ( .A(n22249), .B(n22264), .Z(n22255) );
  XNOR U26923 ( .A(n22247), .B(n22250), .Z(n22264) );
  NAND U26924 ( .A(n22265), .B(n22266), .Z(n22250) );
  NAND U26925 ( .A(n22267), .B(n22268), .Z(n22266) );
  OR U26926 ( .A(n22269), .B(n22270), .Z(n22267) );
  NANDN U26927 ( .A(n22271), .B(n22269), .Z(n22265) );
  IV U26928 ( .A(n22270), .Z(n22271) );
  NAND U26929 ( .A(n22272), .B(n22273), .Z(n22247) );
  NAND U26930 ( .A(n22274), .B(n22275), .Z(n22273) );
  NANDN U26931 ( .A(n22276), .B(n22277), .Z(n22274) );
  NANDN U26932 ( .A(n22277), .B(n22276), .Z(n22272) );
  AND U26933 ( .A(n22278), .B(n22279), .Z(n22249) );
  NAND U26934 ( .A(n22280), .B(n22281), .Z(n22279) );
  OR U26935 ( .A(n22282), .B(n22283), .Z(n22280) );
  NANDN U26936 ( .A(n22284), .B(n22282), .Z(n22278) );
  NAND U26937 ( .A(n22285), .B(n22286), .Z(n22253) );
  NANDN U26938 ( .A(n22287), .B(n22288), .Z(n22286) );
  OR U26939 ( .A(n22289), .B(n22290), .Z(n22288) );
  NANDN U26940 ( .A(n22291), .B(n22289), .Z(n22285) );
  IV U26941 ( .A(n22290), .Z(n22291) );
  XNOR U26942 ( .A(n22261), .B(n22292), .Z(n22256) );
  XNOR U26943 ( .A(n22259), .B(n22262), .Z(n22292) );
  NAND U26944 ( .A(n22293), .B(n22294), .Z(n22262) );
  NAND U26945 ( .A(n22295), .B(n22296), .Z(n22294) );
  OR U26946 ( .A(n22297), .B(n22298), .Z(n22295) );
  NANDN U26947 ( .A(n22299), .B(n22297), .Z(n22293) );
  IV U26948 ( .A(n22298), .Z(n22299) );
  NAND U26949 ( .A(n22300), .B(n22301), .Z(n22259) );
  NAND U26950 ( .A(n22302), .B(n22303), .Z(n22301) );
  NANDN U26951 ( .A(n22304), .B(n22305), .Z(n22302) );
  NANDN U26952 ( .A(n22305), .B(n22304), .Z(n22300) );
  AND U26953 ( .A(n22306), .B(n22307), .Z(n22261) );
  NAND U26954 ( .A(n22308), .B(n22309), .Z(n22307) );
  OR U26955 ( .A(n22310), .B(n22311), .Z(n22308) );
  NANDN U26956 ( .A(n22312), .B(n22310), .Z(n22306) );
  XNOR U26957 ( .A(n22287), .B(n22313), .Z(N28326) );
  XOR U26958 ( .A(n22289), .B(n22290), .Z(n22313) );
  XNOR U26959 ( .A(n22303), .B(n22314), .Z(n22290) );
  XOR U26960 ( .A(n22304), .B(n22305), .Z(n22314) );
  XOR U26961 ( .A(n22310), .B(n22315), .Z(n22305) );
  XOR U26962 ( .A(n22309), .B(n22312), .Z(n22315) );
  IV U26963 ( .A(n22311), .Z(n22312) );
  NAND U26964 ( .A(n22316), .B(n22317), .Z(n22311) );
  OR U26965 ( .A(n22318), .B(n22319), .Z(n22317) );
  OR U26966 ( .A(n22320), .B(n22321), .Z(n22316) );
  NAND U26967 ( .A(n22322), .B(n22323), .Z(n22309) );
  OR U26968 ( .A(n22324), .B(n22325), .Z(n22323) );
  OR U26969 ( .A(n22326), .B(n22327), .Z(n22322) );
  NOR U26970 ( .A(n22328), .B(n22329), .Z(n22310) );
  ANDN U26971 ( .B(n22330), .A(n22331), .Z(n22304) );
  XNOR U26972 ( .A(n22297), .B(n22332), .Z(n22303) );
  XNOR U26973 ( .A(n22296), .B(n22298), .Z(n22332) );
  NAND U26974 ( .A(n22333), .B(n22334), .Z(n22298) );
  OR U26975 ( .A(n22335), .B(n22336), .Z(n22334) );
  OR U26976 ( .A(n22337), .B(n22338), .Z(n22333) );
  NAND U26977 ( .A(n22339), .B(n22340), .Z(n22296) );
  OR U26978 ( .A(n22341), .B(n22342), .Z(n22340) );
  OR U26979 ( .A(n22343), .B(n22344), .Z(n22339) );
  ANDN U26980 ( .B(n22345), .A(n22346), .Z(n22297) );
  IV U26981 ( .A(n22347), .Z(n22345) );
  ANDN U26982 ( .B(n22348), .A(n22349), .Z(n22289) );
  XOR U26983 ( .A(n22275), .B(n22350), .Z(n22287) );
  XOR U26984 ( .A(n22276), .B(n22277), .Z(n22350) );
  XOR U26985 ( .A(n22282), .B(n22351), .Z(n22277) );
  XOR U26986 ( .A(n22281), .B(n22284), .Z(n22351) );
  IV U26987 ( .A(n22283), .Z(n22284) );
  NAND U26988 ( .A(n22352), .B(n22353), .Z(n22283) );
  OR U26989 ( .A(n22354), .B(n22355), .Z(n22353) );
  OR U26990 ( .A(n22356), .B(n22357), .Z(n22352) );
  NAND U26991 ( .A(n22358), .B(n22359), .Z(n22281) );
  OR U26992 ( .A(n22360), .B(n22361), .Z(n22359) );
  OR U26993 ( .A(n22362), .B(n22363), .Z(n22358) );
  NOR U26994 ( .A(n22364), .B(n22365), .Z(n22282) );
  ANDN U26995 ( .B(n22366), .A(n22367), .Z(n22276) );
  IV U26996 ( .A(n22368), .Z(n22366) );
  XNOR U26997 ( .A(n22269), .B(n22369), .Z(n22275) );
  XNOR U26998 ( .A(n22268), .B(n22270), .Z(n22369) );
  NAND U26999 ( .A(n22370), .B(n22371), .Z(n22270) );
  OR U27000 ( .A(n22372), .B(n22373), .Z(n22371) );
  OR U27001 ( .A(n22374), .B(n22375), .Z(n22370) );
  NAND U27002 ( .A(n22376), .B(n22377), .Z(n22268) );
  OR U27003 ( .A(n22378), .B(n22379), .Z(n22377) );
  OR U27004 ( .A(n22380), .B(n22381), .Z(n22376) );
  ANDN U27005 ( .B(n22382), .A(n22383), .Z(n22269) );
  IV U27006 ( .A(n22384), .Z(n22382) );
  XNOR U27007 ( .A(n22349), .B(n22348), .Z(N28325) );
  XOR U27008 ( .A(n22368), .B(n22367), .Z(n22348) );
  XNOR U27009 ( .A(n22383), .B(n22384), .Z(n22367) );
  XNOR U27010 ( .A(n22378), .B(n22379), .Z(n22384) );
  XNOR U27011 ( .A(n22380), .B(n22381), .Z(n22379) );
  XNOR U27012 ( .A(y[796]), .B(x[796]), .Z(n22381) );
  XNOR U27013 ( .A(y[797]), .B(x[797]), .Z(n22380) );
  XNOR U27014 ( .A(y[795]), .B(x[795]), .Z(n22378) );
  XNOR U27015 ( .A(n22372), .B(n22373), .Z(n22383) );
  XNOR U27016 ( .A(y[792]), .B(x[792]), .Z(n22373) );
  XNOR U27017 ( .A(n22374), .B(n22375), .Z(n22372) );
  XNOR U27018 ( .A(y[793]), .B(x[793]), .Z(n22375) );
  XNOR U27019 ( .A(y[794]), .B(x[794]), .Z(n22374) );
  XNOR U27020 ( .A(n22365), .B(n22364), .Z(n22368) );
  XNOR U27021 ( .A(n22360), .B(n22361), .Z(n22364) );
  XNOR U27022 ( .A(y[789]), .B(x[789]), .Z(n22361) );
  XNOR U27023 ( .A(n22362), .B(n22363), .Z(n22360) );
  XNOR U27024 ( .A(y[790]), .B(x[790]), .Z(n22363) );
  XNOR U27025 ( .A(y[791]), .B(x[791]), .Z(n22362) );
  XNOR U27026 ( .A(n22354), .B(n22355), .Z(n22365) );
  XNOR U27027 ( .A(y[786]), .B(x[786]), .Z(n22355) );
  XNOR U27028 ( .A(n22356), .B(n22357), .Z(n22354) );
  XNOR U27029 ( .A(y[787]), .B(x[787]), .Z(n22357) );
  XNOR U27030 ( .A(y[788]), .B(x[788]), .Z(n22356) );
  XOR U27031 ( .A(n22330), .B(n22331), .Z(n22349) );
  XNOR U27032 ( .A(n22346), .B(n22347), .Z(n22331) );
  XNOR U27033 ( .A(n22341), .B(n22342), .Z(n22347) );
  XNOR U27034 ( .A(n22343), .B(n22344), .Z(n22342) );
  XNOR U27035 ( .A(y[784]), .B(x[784]), .Z(n22344) );
  XNOR U27036 ( .A(y[785]), .B(x[785]), .Z(n22343) );
  XNOR U27037 ( .A(y[783]), .B(x[783]), .Z(n22341) );
  XNOR U27038 ( .A(n22335), .B(n22336), .Z(n22346) );
  XNOR U27039 ( .A(y[780]), .B(x[780]), .Z(n22336) );
  XNOR U27040 ( .A(n22337), .B(n22338), .Z(n22335) );
  XNOR U27041 ( .A(y[781]), .B(x[781]), .Z(n22338) );
  XNOR U27042 ( .A(y[782]), .B(x[782]), .Z(n22337) );
  XOR U27043 ( .A(n22329), .B(n22328), .Z(n22330) );
  XNOR U27044 ( .A(n22324), .B(n22325), .Z(n22328) );
  XNOR U27045 ( .A(y[777]), .B(x[777]), .Z(n22325) );
  XNOR U27046 ( .A(n22326), .B(n22327), .Z(n22324) );
  XNOR U27047 ( .A(y[778]), .B(x[778]), .Z(n22327) );
  XNOR U27048 ( .A(y[779]), .B(x[779]), .Z(n22326) );
  XNOR U27049 ( .A(n22318), .B(n22319), .Z(n22329) );
  XNOR U27050 ( .A(y[774]), .B(x[774]), .Z(n22319) );
  XNOR U27051 ( .A(n22320), .B(n22321), .Z(n22318) );
  XNOR U27052 ( .A(y[775]), .B(x[775]), .Z(n22321) );
  XNOR U27053 ( .A(y[776]), .B(x[776]), .Z(n22320) );
  NAND U27054 ( .A(n22385), .B(n22386), .Z(N28317) );
  NANDN U27055 ( .A(n22387), .B(n22388), .Z(n22386) );
  OR U27056 ( .A(n22389), .B(n22390), .Z(n22388) );
  NAND U27057 ( .A(n22389), .B(n22390), .Z(n22385) );
  XOR U27058 ( .A(n22389), .B(n22391), .Z(N28316) );
  XNOR U27059 ( .A(n22387), .B(n22390), .Z(n22391) );
  AND U27060 ( .A(n22392), .B(n22393), .Z(n22390) );
  NANDN U27061 ( .A(n22394), .B(n22395), .Z(n22393) );
  NANDN U27062 ( .A(n22396), .B(n22397), .Z(n22395) );
  NANDN U27063 ( .A(n22397), .B(n22396), .Z(n22392) );
  NAND U27064 ( .A(n22398), .B(n22399), .Z(n22387) );
  NANDN U27065 ( .A(n22400), .B(n22401), .Z(n22399) );
  OR U27066 ( .A(n22402), .B(n22403), .Z(n22401) );
  NAND U27067 ( .A(n22403), .B(n22402), .Z(n22398) );
  AND U27068 ( .A(n22404), .B(n22405), .Z(n22389) );
  NANDN U27069 ( .A(n22406), .B(n22407), .Z(n22405) );
  NANDN U27070 ( .A(n22408), .B(n22409), .Z(n22407) );
  NANDN U27071 ( .A(n22409), .B(n22408), .Z(n22404) );
  XOR U27072 ( .A(n22403), .B(n22410), .Z(N28315) );
  XOR U27073 ( .A(n22400), .B(n22402), .Z(n22410) );
  XNOR U27074 ( .A(n22396), .B(n22411), .Z(n22402) );
  XNOR U27075 ( .A(n22394), .B(n22397), .Z(n22411) );
  NAND U27076 ( .A(n22412), .B(n22413), .Z(n22397) );
  NAND U27077 ( .A(n22414), .B(n22415), .Z(n22413) );
  OR U27078 ( .A(n22416), .B(n22417), .Z(n22414) );
  NANDN U27079 ( .A(n22418), .B(n22416), .Z(n22412) );
  IV U27080 ( .A(n22417), .Z(n22418) );
  NAND U27081 ( .A(n22419), .B(n22420), .Z(n22394) );
  NAND U27082 ( .A(n22421), .B(n22422), .Z(n22420) );
  NANDN U27083 ( .A(n22423), .B(n22424), .Z(n22421) );
  NANDN U27084 ( .A(n22424), .B(n22423), .Z(n22419) );
  AND U27085 ( .A(n22425), .B(n22426), .Z(n22396) );
  NAND U27086 ( .A(n22427), .B(n22428), .Z(n22426) );
  OR U27087 ( .A(n22429), .B(n22430), .Z(n22427) );
  NANDN U27088 ( .A(n22431), .B(n22429), .Z(n22425) );
  NAND U27089 ( .A(n22432), .B(n22433), .Z(n22400) );
  NANDN U27090 ( .A(n22434), .B(n22435), .Z(n22433) );
  OR U27091 ( .A(n22436), .B(n22437), .Z(n22435) );
  NANDN U27092 ( .A(n22438), .B(n22436), .Z(n22432) );
  IV U27093 ( .A(n22437), .Z(n22438) );
  XNOR U27094 ( .A(n22408), .B(n22439), .Z(n22403) );
  XNOR U27095 ( .A(n22406), .B(n22409), .Z(n22439) );
  NAND U27096 ( .A(n22440), .B(n22441), .Z(n22409) );
  NAND U27097 ( .A(n22442), .B(n22443), .Z(n22441) );
  OR U27098 ( .A(n22444), .B(n22445), .Z(n22442) );
  NANDN U27099 ( .A(n22446), .B(n22444), .Z(n22440) );
  IV U27100 ( .A(n22445), .Z(n22446) );
  NAND U27101 ( .A(n22447), .B(n22448), .Z(n22406) );
  NAND U27102 ( .A(n22449), .B(n22450), .Z(n22448) );
  NANDN U27103 ( .A(n22451), .B(n22452), .Z(n22449) );
  NANDN U27104 ( .A(n22452), .B(n22451), .Z(n22447) );
  AND U27105 ( .A(n22453), .B(n22454), .Z(n22408) );
  NAND U27106 ( .A(n22455), .B(n22456), .Z(n22454) );
  OR U27107 ( .A(n22457), .B(n22458), .Z(n22455) );
  NANDN U27108 ( .A(n22459), .B(n22457), .Z(n22453) );
  XNOR U27109 ( .A(n22434), .B(n22460), .Z(N28314) );
  XOR U27110 ( .A(n22436), .B(n22437), .Z(n22460) );
  XNOR U27111 ( .A(n22450), .B(n22461), .Z(n22437) );
  XOR U27112 ( .A(n22451), .B(n22452), .Z(n22461) );
  XOR U27113 ( .A(n22457), .B(n22462), .Z(n22452) );
  XOR U27114 ( .A(n22456), .B(n22459), .Z(n22462) );
  IV U27115 ( .A(n22458), .Z(n22459) );
  NAND U27116 ( .A(n22463), .B(n22464), .Z(n22458) );
  OR U27117 ( .A(n22465), .B(n22466), .Z(n22464) );
  OR U27118 ( .A(n22467), .B(n22468), .Z(n22463) );
  NAND U27119 ( .A(n22469), .B(n22470), .Z(n22456) );
  OR U27120 ( .A(n22471), .B(n22472), .Z(n22470) );
  OR U27121 ( .A(n22473), .B(n22474), .Z(n22469) );
  NOR U27122 ( .A(n22475), .B(n22476), .Z(n22457) );
  ANDN U27123 ( .B(n22477), .A(n22478), .Z(n22451) );
  XNOR U27124 ( .A(n22444), .B(n22479), .Z(n22450) );
  XNOR U27125 ( .A(n22443), .B(n22445), .Z(n22479) );
  NAND U27126 ( .A(n22480), .B(n22481), .Z(n22445) );
  OR U27127 ( .A(n22482), .B(n22483), .Z(n22481) );
  OR U27128 ( .A(n22484), .B(n22485), .Z(n22480) );
  NAND U27129 ( .A(n22486), .B(n22487), .Z(n22443) );
  OR U27130 ( .A(n22488), .B(n22489), .Z(n22487) );
  OR U27131 ( .A(n22490), .B(n22491), .Z(n22486) );
  ANDN U27132 ( .B(n22492), .A(n22493), .Z(n22444) );
  IV U27133 ( .A(n22494), .Z(n22492) );
  ANDN U27134 ( .B(n22495), .A(n22496), .Z(n22436) );
  XOR U27135 ( .A(n22422), .B(n22497), .Z(n22434) );
  XOR U27136 ( .A(n22423), .B(n22424), .Z(n22497) );
  XOR U27137 ( .A(n22429), .B(n22498), .Z(n22424) );
  XOR U27138 ( .A(n22428), .B(n22431), .Z(n22498) );
  IV U27139 ( .A(n22430), .Z(n22431) );
  NAND U27140 ( .A(n22499), .B(n22500), .Z(n22430) );
  OR U27141 ( .A(n22501), .B(n22502), .Z(n22500) );
  OR U27142 ( .A(n22503), .B(n22504), .Z(n22499) );
  NAND U27143 ( .A(n22505), .B(n22506), .Z(n22428) );
  OR U27144 ( .A(n22507), .B(n22508), .Z(n22506) );
  OR U27145 ( .A(n22509), .B(n22510), .Z(n22505) );
  NOR U27146 ( .A(n22511), .B(n22512), .Z(n22429) );
  ANDN U27147 ( .B(n22513), .A(n22514), .Z(n22423) );
  IV U27148 ( .A(n22515), .Z(n22513) );
  XNOR U27149 ( .A(n22416), .B(n22516), .Z(n22422) );
  XNOR U27150 ( .A(n22415), .B(n22417), .Z(n22516) );
  NAND U27151 ( .A(n22517), .B(n22518), .Z(n22417) );
  OR U27152 ( .A(n22519), .B(n22520), .Z(n22518) );
  OR U27153 ( .A(n22521), .B(n22522), .Z(n22517) );
  NAND U27154 ( .A(n22523), .B(n22524), .Z(n22415) );
  OR U27155 ( .A(n22525), .B(n22526), .Z(n22524) );
  OR U27156 ( .A(n22527), .B(n22528), .Z(n22523) );
  ANDN U27157 ( .B(n22529), .A(n22530), .Z(n22416) );
  IV U27158 ( .A(n22531), .Z(n22529) );
  XNOR U27159 ( .A(n22496), .B(n22495), .Z(N28313) );
  XOR U27160 ( .A(n22515), .B(n22514), .Z(n22495) );
  XNOR U27161 ( .A(n22530), .B(n22531), .Z(n22514) );
  XNOR U27162 ( .A(n22525), .B(n22526), .Z(n22531) );
  XNOR U27163 ( .A(n22527), .B(n22528), .Z(n22526) );
  XNOR U27164 ( .A(y[772]), .B(x[772]), .Z(n22528) );
  XNOR U27165 ( .A(y[773]), .B(x[773]), .Z(n22527) );
  XNOR U27166 ( .A(y[771]), .B(x[771]), .Z(n22525) );
  XNOR U27167 ( .A(n22519), .B(n22520), .Z(n22530) );
  XNOR U27168 ( .A(y[768]), .B(x[768]), .Z(n22520) );
  XNOR U27169 ( .A(n22521), .B(n22522), .Z(n22519) );
  XNOR U27170 ( .A(y[769]), .B(x[769]), .Z(n22522) );
  XNOR U27171 ( .A(y[770]), .B(x[770]), .Z(n22521) );
  XNOR U27172 ( .A(n22512), .B(n22511), .Z(n22515) );
  XNOR U27173 ( .A(n22507), .B(n22508), .Z(n22511) );
  XNOR U27174 ( .A(y[765]), .B(x[765]), .Z(n22508) );
  XNOR U27175 ( .A(n22509), .B(n22510), .Z(n22507) );
  XNOR U27176 ( .A(y[766]), .B(x[766]), .Z(n22510) );
  XNOR U27177 ( .A(y[767]), .B(x[767]), .Z(n22509) );
  XNOR U27178 ( .A(n22501), .B(n22502), .Z(n22512) );
  XNOR U27179 ( .A(y[762]), .B(x[762]), .Z(n22502) );
  XNOR U27180 ( .A(n22503), .B(n22504), .Z(n22501) );
  XNOR U27181 ( .A(y[763]), .B(x[763]), .Z(n22504) );
  XNOR U27182 ( .A(y[764]), .B(x[764]), .Z(n22503) );
  XOR U27183 ( .A(n22477), .B(n22478), .Z(n22496) );
  XNOR U27184 ( .A(n22493), .B(n22494), .Z(n22478) );
  XNOR U27185 ( .A(n22488), .B(n22489), .Z(n22494) );
  XNOR U27186 ( .A(n22490), .B(n22491), .Z(n22489) );
  XNOR U27187 ( .A(y[760]), .B(x[760]), .Z(n22491) );
  XNOR U27188 ( .A(y[761]), .B(x[761]), .Z(n22490) );
  XNOR U27189 ( .A(y[759]), .B(x[759]), .Z(n22488) );
  XNOR U27190 ( .A(n22482), .B(n22483), .Z(n22493) );
  XNOR U27191 ( .A(y[756]), .B(x[756]), .Z(n22483) );
  XNOR U27192 ( .A(n22484), .B(n22485), .Z(n22482) );
  XNOR U27193 ( .A(y[757]), .B(x[757]), .Z(n22485) );
  XNOR U27194 ( .A(y[758]), .B(x[758]), .Z(n22484) );
  XOR U27195 ( .A(n22476), .B(n22475), .Z(n22477) );
  XNOR U27196 ( .A(n22471), .B(n22472), .Z(n22475) );
  XNOR U27197 ( .A(y[753]), .B(x[753]), .Z(n22472) );
  XNOR U27198 ( .A(n22473), .B(n22474), .Z(n22471) );
  XNOR U27199 ( .A(y[754]), .B(x[754]), .Z(n22474) );
  XNOR U27200 ( .A(y[755]), .B(x[755]), .Z(n22473) );
  XNOR U27201 ( .A(n22465), .B(n22466), .Z(n22476) );
  XNOR U27202 ( .A(y[750]), .B(x[750]), .Z(n22466) );
  XNOR U27203 ( .A(n22467), .B(n22468), .Z(n22465) );
  XNOR U27204 ( .A(y[751]), .B(x[751]), .Z(n22468) );
  XNOR U27205 ( .A(y[752]), .B(x[752]), .Z(n22467) );
  NAND U27206 ( .A(n22532), .B(n22533), .Z(N28305) );
  NANDN U27207 ( .A(n22534), .B(n22535), .Z(n22533) );
  OR U27208 ( .A(n22536), .B(n22537), .Z(n22535) );
  NAND U27209 ( .A(n22536), .B(n22537), .Z(n22532) );
  XOR U27210 ( .A(n22536), .B(n22538), .Z(N28304) );
  XNOR U27211 ( .A(n22534), .B(n22537), .Z(n22538) );
  AND U27212 ( .A(n22539), .B(n22540), .Z(n22537) );
  NANDN U27213 ( .A(n22541), .B(n22542), .Z(n22540) );
  NANDN U27214 ( .A(n22543), .B(n22544), .Z(n22542) );
  NANDN U27215 ( .A(n22544), .B(n22543), .Z(n22539) );
  NAND U27216 ( .A(n22545), .B(n22546), .Z(n22534) );
  NANDN U27217 ( .A(n22547), .B(n22548), .Z(n22546) );
  OR U27218 ( .A(n22549), .B(n22550), .Z(n22548) );
  NAND U27219 ( .A(n22550), .B(n22549), .Z(n22545) );
  AND U27220 ( .A(n22551), .B(n22552), .Z(n22536) );
  NANDN U27221 ( .A(n22553), .B(n22554), .Z(n22552) );
  NANDN U27222 ( .A(n22555), .B(n22556), .Z(n22554) );
  NANDN U27223 ( .A(n22556), .B(n22555), .Z(n22551) );
  XOR U27224 ( .A(n22550), .B(n22557), .Z(N28303) );
  XOR U27225 ( .A(n22547), .B(n22549), .Z(n22557) );
  XNOR U27226 ( .A(n22543), .B(n22558), .Z(n22549) );
  XNOR U27227 ( .A(n22541), .B(n22544), .Z(n22558) );
  NAND U27228 ( .A(n22559), .B(n22560), .Z(n22544) );
  NAND U27229 ( .A(n22561), .B(n22562), .Z(n22560) );
  OR U27230 ( .A(n22563), .B(n22564), .Z(n22561) );
  NANDN U27231 ( .A(n22565), .B(n22563), .Z(n22559) );
  IV U27232 ( .A(n22564), .Z(n22565) );
  NAND U27233 ( .A(n22566), .B(n22567), .Z(n22541) );
  NAND U27234 ( .A(n22568), .B(n22569), .Z(n22567) );
  NANDN U27235 ( .A(n22570), .B(n22571), .Z(n22568) );
  NANDN U27236 ( .A(n22571), .B(n22570), .Z(n22566) );
  AND U27237 ( .A(n22572), .B(n22573), .Z(n22543) );
  NAND U27238 ( .A(n22574), .B(n22575), .Z(n22573) );
  OR U27239 ( .A(n22576), .B(n22577), .Z(n22574) );
  NANDN U27240 ( .A(n22578), .B(n22576), .Z(n22572) );
  NAND U27241 ( .A(n22579), .B(n22580), .Z(n22547) );
  NANDN U27242 ( .A(n22581), .B(n22582), .Z(n22580) );
  OR U27243 ( .A(n22583), .B(n22584), .Z(n22582) );
  NANDN U27244 ( .A(n22585), .B(n22583), .Z(n22579) );
  IV U27245 ( .A(n22584), .Z(n22585) );
  XNOR U27246 ( .A(n22555), .B(n22586), .Z(n22550) );
  XNOR U27247 ( .A(n22553), .B(n22556), .Z(n22586) );
  NAND U27248 ( .A(n22587), .B(n22588), .Z(n22556) );
  NAND U27249 ( .A(n22589), .B(n22590), .Z(n22588) );
  OR U27250 ( .A(n22591), .B(n22592), .Z(n22589) );
  NANDN U27251 ( .A(n22593), .B(n22591), .Z(n22587) );
  IV U27252 ( .A(n22592), .Z(n22593) );
  NAND U27253 ( .A(n22594), .B(n22595), .Z(n22553) );
  NAND U27254 ( .A(n22596), .B(n22597), .Z(n22595) );
  NANDN U27255 ( .A(n22598), .B(n22599), .Z(n22596) );
  NANDN U27256 ( .A(n22599), .B(n22598), .Z(n22594) );
  AND U27257 ( .A(n22600), .B(n22601), .Z(n22555) );
  NAND U27258 ( .A(n22602), .B(n22603), .Z(n22601) );
  OR U27259 ( .A(n22604), .B(n22605), .Z(n22602) );
  NANDN U27260 ( .A(n22606), .B(n22604), .Z(n22600) );
  XNOR U27261 ( .A(n22581), .B(n22607), .Z(N28302) );
  XOR U27262 ( .A(n22583), .B(n22584), .Z(n22607) );
  XNOR U27263 ( .A(n22597), .B(n22608), .Z(n22584) );
  XOR U27264 ( .A(n22598), .B(n22599), .Z(n22608) );
  XOR U27265 ( .A(n22604), .B(n22609), .Z(n22599) );
  XOR U27266 ( .A(n22603), .B(n22606), .Z(n22609) );
  IV U27267 ( .A(n22605), .Z(n22606) );
  NAND U27268 ( .A(n22610), .B(n22611), .Z(n22605) );
  OR U27269 ( .A(n22612), .B(n22613), .Z(n22611) );
  OR U27270 ( .A(n22614), .B(n22615), .Z(n22610) );
  NAND U27271 ( .A(n22616), .B(n22617), .Z(n22603) );
  OR U27272 ( .A(n22618), .B(n22619), .Z(n22617) );
  OR U27273 ( .A(n22620), .B(n22621), .Z(n22616) );
  NOR U27274 ( .A(n22622), .B(n22623), .Z(n22604) );
  ANDN U27275 ( .B(n22624), .A(n22625), .Z(n22598) );
  XNOR U27276 ( .A(n22591), .B(n22626), .Z(n22597) );
  XNOR U27277 ( .A(n22590), .B(n22592), .Z(n22626) );
  NAND U27278 ( .A(n22627), .B(n22628), .Z(n22592) );
  OR U27279 ( .A(n22629), .B(n22630), .Z(n22628) );
  OR U27280 ( .A(n22631), .B(n22632), .Z(n22627) );
  NAND U27281 ( .A(n22633), .B(n22634), .Z(n22590) );
  OR U27282 ( .A(n22635), .B(n22636), .Z(n22634) );
  OR U27283 ( .A(n22637), .B(n22638), .Z(n22633) );
  ANDN U27284 ( .B(n22639), .A(n22640), .Z(n22591) );
  IV U27285 ( .A(n22641), .Z(n22639) );
  ANDN U27286 ( .B(n22642), .A(n22643), .Z(n22583) );
  XOR U27287 ( .A(n22569), .B(n22644), .Z(n22581) );
  XOR U27288 ( .A(n22570), .B(n22571), .Z(n22644) );
  XOR U27289 ( .A(n22576), .B(n22645), .Z(n22571) );
  XOR U27290 ( .A(n22575), .B(n22578), .Z(n22645) );
  IV U27291 ( .A(n22577), .Z(n22578) );
  NAND U27292 ( .A(n22646), .B(n22647), .Z(n22577) );
  OR U27293 ( .A(n22648), .B(n22649), .Z(n22647) );
  OR U27294 ( .A(n22650), .B(n22651), .Z(n22646) );
  NAND U27295 ( .A(n22652), .B(n22653), .Z(n22575) );
  OR U27296 ( .A(n22654), .B(n22655), .Z(n22653) );
  OR U27297 ( .A(n22656), .B(n22657), .Z(n22652) );
  NOR U27298 ( .A(n22658), .B(n22659), .Z(n22576) );
  ANDN U27299 ( .B(n22660), .A(n22661), .Z(n22570) );
  IV U27300 ( .A(n22662), .Z(n22660) );
  XNOR U27301 ( .A(n22563), .B(n22663), .Z(n22569) );
  XNOR U27302 ( .A(n22562), .B(n22564), .Z(n22663) );
  NAND U27303 ( .A(n22664), .B(n22665), .Z(n22564) );
  OR U27304 ( .A(n22666), .B(n22667), .Z(n22665) );
  OR U27305 ( .A(n22668), .B(n22669), .Z(n22664) );
  NAND U27306 ( .A(n22670), .B(n22671), .Z(n22562) );
  OR U27307 ( .A(n22672), .B(n22673), .Z(n22671) );
  OR U27308 ( .A(n22674), .B(n22675), .Z(n22670) );
  ANDN U27309 ( .B(n22676), .A(n22677), .Z(n22563) );
  IV U27310 ( .A(n22678), .Z(n22676) );
  XNOR U27311 ( .A(n22643), .B(n22642), .Z(N28301) );
  XOR U27312 ( .A(n22662), .B(n22661), .Z(n22642) );
  XNOR U27313 ( .A(n22677), .B(n22678), .Z(n22661) );
  XNOR U27314 ( .A(n22672), .B(n22673), .Z(n22678) );
  XNOR U27315 ( .A(n22674), .B(n22675), .Z(n22673) );
  XNOR U27316 ( .A(y[748]), .B(x[748]), .Z(n22675) );
  XNOR U27317 ( .A(y[749]), .B(x[749]), .Z(n22674) );
  XNOR U27318 ( .A(y[747]), .B(x[747]), .Z(n22672) );
  XNOR U27319 ( .A(n22666), .B(n22667), .Z(n22677) );
  XNOR U27320 ( .A(y[744]), .B(x[744]), .Z(n22667) );
  XNOR U27321 ( .A(n22668), .B(n22669), .Z(n22666) );
  XNOR U27322 ( .A(y[745]), .B(x[745]), .Z(n22669) );
  XNOR U27323 ( .A(y[746]), .B(x[746]), .Z(n22668) );
  XNOR U27324 ( .A(n22659), .B(n22658), .Z(n22662) );
  XNOR U27325 ( .A(n22654), .B(n22655), .Z(n22658) );
  XNOR U27326 ( .A(y[741]), .B(x[741]), .Z(n22655) );
  XNOR U27327 ( .A(n22656), .B(n22657), .Z(n22654) );
  XNOR U27328 ( .A(y[742]), .B(x[742]), .Z(n22657) );
  XNOR U27329 ( .A(y[743]), .B(x[743]), .Z(n22656) );
  XNOR U27330 ( .A(n22648), .B(n22649), .Z(n22659) );
  XNOR U27331 ( .A(y[738]), .B(x[738]), .Z(n22649) );
  XNOR U27332 ( .A(n22650), .B(n22651), .Z(n22648) );
  XNOR U27333 ( .A(y[739]), .B(x[739]), .Z(n22651) );
  XNOR U27334 ( .A(y[740]), .B(x[740]), .Z(n22650) );
  XOR U27335 ( .A(n22624), .B(n22625), .Z(n22643) );
  XNOR U27336 ( .A(n22640), .B(n22641), .Z(n22625) );
  XNOR U27337 ( .A(n22635), .B(n22636), .Z(n22641) );
  XNOR U27338 ( .A(n22637), .B(n22638), .Z(n22636) );
  XNOR U27339 ( .A(y[736]), .B(x[736]), .Z(n22638) );
  XNOR U27340 ( .A(y[737]), .B(x[737]), .Z(n22637) );
  XNOR U27341 ( .A(y[735]), .B(x[735]), .Z(n22635) );
  XNOR U27342 ( .A(n22629), .B(n22630), .Z(n22640) );
  XNOR U27343 ( .A(y[732]), .B(x[732]), .Z(n22630) );
  XNOR U27344 ( .A(n22631), .B(n22632), .Z(n22629) );
  XNOR U27345 ( .A(y[733]), .B(x[733]), .Z(n22632) );
  XNOR U27346 ( .A(y[734]), .B(x[734]), .Z(n22631) );
  XOR U27347 ( .A(n22623), .B(n22622), .Z(n22624) );
  XNOR U27348 ( .A(n22618), .B(n22619), .Z(n22622) );
  XNOR U27349 ( .A(y[729]), .B(x[729]), .Z(n22619) );
  XNOR U27350 ( .A(n22620), .B(n22621), .Z(n22618) );
  XNOR U27351 ( .A(y[730]), .B(x[730]), .Z(n22621) );
  XNOR U27352 ( .A(y[731]), .B(x[731]), .Z(n22620) );
  XNOR U27353 ( .A(n22612), .B(n22613), .Z(n22623) );
  XNOR U27354 ( .A(y[726]), .B(x[726]), .Z(n22613) );
  XNOR U27355 ( .A(n22614), .B(n22615), .Z(n22612) );
  XNOR U27356 ( .A(y[727]), .B(x[727]), .Z(n22615) );
  XNOR U27357 ( .A(y[728]), .B(x[728]), .Z(n22614) );
  NAND U27358 ( .A(n22679), .B(n22680), .Z(N28293) );
  NANDN U27359 ( .A(n22681), .B(n22682), .Z(n22680) );
  OR U27360 ( .A(n22683), .B(n22684), .Z(n22682) );
  NAND U27361 ( .A(n22683), .B(n22684), .Z(n22679) );
  XOR U27362 ( .A(n22683), .B(n22685), .Z(N28292) );
  XNOR U27363 ( .A(n22681), .B(n22684), .Z(n22685) );
  AND U27364 ( .A(n22686), .B(n22687), .Z(n22684) );
  NANDN U27365 ( .A(n22688), .B(n22689), .Z(n22687) );
  NANDN U27366 ( .A(n22690), .B(n22691), .Z(n22689) );
  NANDN U27367 ( .A(n22691), .B(n22690), .Z(n22686) );
  NAND U27368 ( .A(n22692), .B(n22693), .Z(n22681) );
  NANDN U27369 ( .A(n22694), .B(n22695), .Z(n22693) );
  OR U27370 ( .A(n22696), .B(n22697), .Z(n22695) );
  NAND U27371 ( .A(n22697), .B(n22696), .Z(n22692) );
  AND U27372 ( .A(n22698), .B(n22699), .Z(n22683) );
  NANDN U27373 ( .A(n22700), .B(n22701), .Z(n22699) );
  NANDN U27374 ( .A(n22702), .B(n22703), .Z(n22701) );
  NANDN U27375 ( .A(n22703), .B(n22702), .Z(n22698) );
  XOR U27376 ( .A(n22697), .B(n22704), .Z(N28291) );
  XOR U27377 ( .A(n22694), .B(n22696), .Z(n22704) );
  XNOR U27378 ( .A(n22690), .B(n22705), .Z(n22696) );
  XNOR U27379 ( .A(n22688), .B(n22691), .Z(n22705) );
  NAND U27380 ( .A(n22706), .B(n22707), .Z(n22691) );
  NAND U27381 ( .A(n22708), .B(n22709), .Z(n22707) );
  OR U27382 ( .A(n22710), .B(n22711), .Z(n22708) );
  NANDN U27383 ( .A(n22712), .B(n22710), .Z(n22706) );
  IV U27384 ( .A(n22711), .Z(n22712) );
  NAND U27385 ( .A(n22713), .B(n22714), .Z(n22688) );
  NAND U27386 ( .A(n22715), .B(n22716), .Z(n22714) );
  NANDN U27387 ( .A(n22717), .B(n22718), .Z(n22715) );
  NANDN U27388 ( .A(n22718), .B(n22717), .Z(n22713) );
  AND U27389 ( .A(n22719), .B(n22720), .Z(n22690) );
  NAND U27390 ( .A(n22721), .B(n22722), .Z(n22720) );
  OR U27391 ( .A(n22723), .B(n22724), .Z(n22721) );
  NANDN U27392 ( .A(n22725), .B(n22723), .Z(n22719) );
  NAND U27393 ( .A(n22726), .B(n22727), .Z(n22694) );
  NANDN U27394 ( .A(n22728), .B(n22729), .Z(n22727) );
  OR U27395 ( .A(n22730), .B(n22731), .Z(n22729) );
  NANDN U27396 ( .A(n22732), .B(n22730), .Z(n22726) );
  IV U27397 ( .A(n22731), .Z(n22732) );
  XNOR U27398 ( .A(n22702), .B(n22733), .Z(n22697) );
  XNOR U27399 ( .A(n22700), .B(n22703), .Z(n22733) );
  NAND U27400 ( .A(n22734), .B(n22735), .Z(n22703) );
  NAND U27401 ( .A(n22736), .B(n22737), .Z(n22735) );
  OR U27402 ( .A(n22738), .B(n22739), .Z(n22736) );
  NANDN U27403 ( .A(n22740), .B(n22738), .Z(n22734) );
  IV U27404 ( .A(n22739), .Z(n22740) );
  NAND U27405 ( .A(n22741), .B(n22742), .Z(n22700) );
  NAND U27406 ( .A(n22743), .B(n22744), .Z(n22742) );
  NANDN U27407 ( .A(n22745), .B(n22746), .Z(n22743) );
  NANDN U27408 ( .A(n22746), .B(n22745), .Z(n22741) );
  AND U27409 ( .A(n22747), .B(n22748), .Z(n22702) );
  NAND U27410 ( .A(n22749), .B(n22750), .Z(n22748) );
  OR U27411 ( .A(n22751), .B(n22752), .Z(n22749) );
  NANDN U27412 ( .A(n22753), .B(n22751), .Z(n22747) );
  XNOR U27413 ( .A(n22728), .B(n22754), .Z(N28290) );
  XOR U27414 ( .A(n22730), .B(n22731), .Z(n22754) );
  XNOR U27415 ( .A(n22744), .B(n22755), .Z(n22731) );
  XOR U27416 ( .A(n22745), .B(n22746), .Z(n22755) );
  XOR U27417 ( .A(n22751), .B(n22756), .Z(n22746) );
  XOR U27418 ( .A(n22750), .B(n22753), .Z(n22756) );
  IV U27419 ( .A(n22752), .Z(n22753) );
  NAND U27420 ( .A(n22757), .B(n22758), .Z(n22752) );
  OR U27421 ( .A(n22759), .B(n22760), .Z(n22758) );
  OR U27422 ( .A(n22761), .B(n22762), .Z(n22757) );
  NAND U27423 ( .A(n22763), .B(n22764), .Z(n22750) );
  OR U27424 ( .A(n22765), .B(n22766), .Z(n22764) );
  OR U27425 ( .A(n22767), .B(n22768), .Z(n22763) );
  NOR U27426 ( .A(n22769), .B(n22770), .Z(n22751) );
  ANDN U27427 ( .B(n22771), .A(n22772), .Z(n22745) );
  XNOR U27428 ( .A(n22738), .B(n22773), .Z(n22744) );
  XNOR U27429 ( .A(n22737), .B(n22739), .Z(n22773) );
  NAND U27430 ( .A(n22774), .B(n22775), .Z(n22739) );
  OR U27431 ( .A(n22776), .B(n22777), .Z(n22775) );
  OR U27432 ( .A(n22778), .B(n22779), .Z(n22774) );
  NAND U27433 ( .A(n22780), .B(n22781), .Z(n22737) );
  OR U27434 ( .A(n22782), .B(n22783), .Z(n22781) );
  OR U27435 ( .A(n22784), .B(n22785), .Z(n22780) );
  ANDN U27436 ( .B(n22786), .A(n22787), .Z(n22738) );
  IV U27437 ( .A(n22788), .Z(n22786) );
  ANDN U27438 ( .B(n22789), .A(n22790), .Z(n22730) );
  XOR U27439 ( .A(n22716), .B(n22791), .Z(n22728) );
  XOR U27440 ( .A(n22717), .B(n22718), .Z(n22791) );
  XOR U27441 ( .A(n22723), .B(n22792), .Z(n22718) );
  XOR U27442 ( .A(n22722), .B(n22725), .Z(n22792) );
  IV U27443 ( .A(n22724), .Z(n22725) );
  NAND U27444 ( .A(n22793), .B(n22794), .Z(n22724) );
  OR U27445 ( .A(n22795), .B(n22796), .Z(n22794) );
  OR U27446 ( .A(n22797), .B(n22798), .Z(n22793) );
  NAND U27447 ( .A(n22799), .B(n22800), .Z(n22722) );
  OR U27448 ( .A(n22801), .B(n22802), .Z(n22800) );
  OR U27449 ( .A(n22803), .B(n22804), .Z(n22799) );
  NOR U27450 ( .A(n22805), .B(n22806), .Z(n22723) );
  ANDN U27451 ( .B(n22807), .A(n22808), .Z(n22717) );
  IV U27452 ( .A(n22809), .Z(n22807) );
  XNOR U27453 ( .A(n22710), .B(n22810), .Z(n22716) );
  XNOR U27454 ( .A(n22709), .B(n22711), .Z(n22810) );
  NAND U27455 ( .A(n22811), .B(n22812), .Z(n22711) );
  OR U27456 ( .A(n22813), .B(n22814), .Z(n22812) );
  OR U27457 ( .A(n22815), .B(n22816), .Z(n22811) );
  NAND U27458 ( .A(n22817), .B(n22818), .Z(n22709) );
  OR U27459 ( .A(n22819), .B(n22820), .Z(n22818) );
  OR U27460 ( .A(n22821), .B(n22822), .Z(n22817) );
  ANDN U27461 ( .B(n22823), .A(n22824), .Z(n22710) );
  IV U27462 ( .A(n22825), .Z(n22823) );
  XNOR U27463 ( .A(n22790), .B(n22789), .Z(N28289) );
  XOR U27464 ( .A(n22809), .B(n22808), .Z(n22789) );
  XNOR U27465 ( .A(n22824), .B(n22825), .Z(n22808) );
  XNOR U27466 ( .A(n22819), .B(n22820), .Z(n22825) );
  XNOR U27467 ( .A(n22821), .B(n22822), .Z(n22820) );
  XNOR U27468 ( .A(y[724]), .B(x[724]), .Z(n22822) );
  XNOR U27469 ( .A(y[725]), .B(x[725]), .Z(n22821) );
  XNOR U27470 ( .A(y[723]), .B(x[723]), .Z(n22819) );
  XNOR U27471 ( .A(n22813), .B(n22814), .Z(n22824) );
  XNOR U27472 ( .A(y[720]), .B(x[720]), .Z(n22814) );
  XNOR U27473 ( .A(n22815), .B(n22816), .Z(n22813) );
  XNOR U27474 ( .A(y[721]), .B(x[721]), .Z(n22816) );
  XNOR U27475 ( .A(y[722]), .B(x[722]), .Z(n22815) );
  XNOR U27476 ( .A(n22806), .B(n22805), .Z(n22809) );
  XNOR U27477 ( .A(n22801), .B(n22802), .Z(n22805) );
  XNOR U27478 ( .A(y[717]), .B(x[717]), .Z(n22802) );
  XNOR U27479 ( .A(n22803), .B(n22804), .Z(n22801) );
  XNOR U27480 ( .A(y[718]), .B(x[718]), .Z(n22804) );
  XNOR U27481 ( .A(y[719]), .B(x[719]), .Z(n22803) );
  XNOR U27482 ( .A(n22795), .B(n22796), .Z(n22806) );
  XNOR U27483 ( .A(y[714]), .B(x[714]), .Z(n22796) );
  XNOR U27484 ( .A(n22797), .B(n22798), .Z(n22795) );
  XNOR U27485 ( .A(y[715]), .B(x[715]), .Z(n22798) );
  XNOR U27486 ( .A(y[716]), .B(x[716]), .Z(n22797) );
  XOR U27487 ( .A(n22771), .B(n22772), .Z(n22790) );
  XNOR U27488 ( .A(n22787), .B(n22788), .Z(n22772) );
  XNOR U27489 ( .A(n22782), .B(n22783), .Z(n22788) );
  XNOR U27490 ( .A(n22784), .B(n22785), .Z(n22783) );
  XNOR U27491 ( .A(y[712]), .B(x[712]), .Z(n22785) );
  XNOR U27492 ( .A(y[713]), .B(x[713]), .Z(n22784) );
  XNOR U27493 ( .A(y[711]), .B(x[711]), .Z(n22782) );
  XNOR U27494 ( .A(n22776), .B(n22777), .Z(n22787) );
  XNOR U27495 ( .A(y[708]), .B(x[708]), .Z(n22777) );
  XNOR U27496 ( .A(n22778), .B(n22779), .Z(n22776) );
  XNOR U27497 ( .A(y[709]), .B(x[709]), .Z(n22779) );
  XNOR U27498 ( .A(y[710]), .B(x[710]), .Z(n22778) );
  XOR U27499 ( .A(n22770), .B(n22769), .Z(n22771) );
  XNOR U27500 ( .A(n22765), .B(n22766), .Z(n22769) );
  XNOR U27501 ( .A(y[705]), .B(x[705]), .Z(n22766) );
  XNOR U27502 ( .A(n22767), .B(n22768), .Z(n22765) );
  XNOR U27503 ( .A(y[706]), .B(x[706]), .Z(n22768) );
  XNOR U27504 ( .A(y[707]), .B(x[707]), .Z(n22767) );
  XNOR U27505 ( .A(n22759), .B(n22760), .Z(n22770) );
  XNOR U27506 ( .A(y[702]), .B(x[702]), .Z(n22760) );
  XNOR U27507 ( .A(n22761), .B(n22762), .Z(n22759) );
  XNOR U27508 ( .A(y[703]), .B(x[703]), .Z(n22762) );
  XNOR U27509 ( .A(y[704]), .B(x[704]), .Z(n22761) );
  NAND U27510 ( .A(n22826), .B(n22827), .Z(N28281) );
  NANDN U27511 ( .A(n22828), .B(n22829), .Z(n22827) );
  OR U27512 ( .A(n22830), .B(n22831), .Z(n22829) );
  NAND U27513 ( .A(n22830), .B(n22831), .Z(n22826) );
  XOR U27514 ( .A(n22830), .B(n22832), .Z(N28280) );
  XNOR U27515 ( .A(n22828), .B(n22831), .Z(n22832) );
  AND U27516 ( .A(n22833), .B(n22834), .Z(n22831) );
  NANDN U27517 ( .A(n22835), .B(n22836), .Z(n22834) );
  NANDN U27518 ( .A(n22837), .B(n22838), .Z(n22836) );
  NANDN U27519 ( .A(n22838), .B(n22837), .Z(n22833) );
  NAND U27520 ( .A(n22839), .B(n22840), .Z(n22828) );
  NANDN U27521 ( .A(n22841), .B(n22842), .Z(n22840) );
  OR U27522 ( .A(n22843), .B(n22844), .Z(n22842) );
  NAND U27523 ( .A(n22844), .B(n22843), .Z(n22839) );
  AND U27524 ( .A(n22845), .B(n22846), .Z(n22830) );
  NANDN U27525 ( .A(n22847), .B(n22848), .Z(n22846) );
  NANDN U27526 ( .A(n22849), .B(n22850), .Z(n22848) );
  NANDN U27527 ( .A(n22850), .B(n22849), .Z(n22845) );
  XOR U27528 ( .A(n22844), .B(n22851), .Z(N28279) );
  XOR U27529 ( .A(n22841), .B(n22843), .Z(n22851) );
  XNOR U27530 ( .A(n22837), .B(n22852), .Z(n22843) );
  XNOR U27531 ( .A(n22835), .B(n22838), .Z(n22852) );
  NAND U27532 ( .A(n22853), .B(n22854), .Z(n22838) );
  NAND U27533 ( .A(n22855), .B(n22856), .Z(n22854) );
  OR U27534 ( .A(n22857), .B(n22858), .Z(n22855) );
  NANDN U27535 ( .A(n22859), .B(n22857), .Z(n22853) );
  IV U27536 ( .A(n22858), .Z(n22859) );
  NAND U27537 ( .A(n22860), .B(n22861), .Z(n22835) );
  NAND U27538 ( .A(n22862), .B(n22863), .Z(n22861) );
  NANDN U27539 ( .A(n22864), .B(n22865), .Z(n22862) );
  NANDN U27540 ( .A(n22865), .B(n22864), .Z(n22860) );
  AND U27541 ( .A(n22866), .B(n22867), .Z(n22837) );
  NAND U27542 ( .A(n22868), .B(n22869), .Z(n22867) );
  OR U27543 ( .A(n22870), .B(n22871), .Z(n22868) );
  NANDN U27544 ( .A(n22872), .B(n22870), .Z(n22866) );
  NAND U27545 ( .A(n22873), .B(n22874), .Z(n22841) );
  NANDN U27546 ( .A(n22875), .B(n22876), .Z(n22874) );
  OR U27547 ( .A(n22877), .B(n22878), .Z(n22876) );
  NANDN U27548 ( .A(n22879), .B(n22877), .Z(n22873) );
  IV U27549 ( .A(n22878), .Z(n22879) );
  XNOR U27550 ( .A(n22849), .B(n22880), .Z(n22844) );
  XNOR U27551 ( .A(n22847), .B(n22850), .Z(n22880) );
  NAND U27552 ( .A(n22881), .B(n22882), .Z(n22850) );
  NAND U27553 ( .A(n22883), .B(n22884), .Z(n22882) );
  OR U27554 ( .A(n22885), .B(n22886), .Z(n22883) );
  NANDN U27555 ( .A(n22887), .B(n22885), .Z(n22881) );
  IV U27556 ( .A(n22886), .Z(n22887) );
  NAND U27557 ( .A(n22888), .B(n22889), .Z(n22847) );
  NAND U27558 ( .A(n22890), .B(n22891), .Z(n22889) );
  NANDN U27559 ( .A(n22892), .B(n22893), .Z(n22890) );
  NANDN U27560 ( .A(n22893), .B(n22892), .Z(n22888) );
  AND U27561 ( .A(n22894), .B(n22895), .Z(n22849) );
  NAND U27562 ( .A(n22896), .B(n22897), .Z(n22895) );
  OR U27563 ( .A(n22898), .B(n22899), .Z(n22896) );
  NANDN U27564 ( .A(n22900), .B(n22898), .Z(n22894) );
  XNOR U27565 ( .A(n22875), .B(n22901), .Z(N28278) );
  XOR U27566 ( .A(n22877), .B(n22878), .Z(n22901) );
  XNOR U27567 ( .A(n22891), .B(n22902), .Z(n22878) );
  XOR U27568 ( .A(n22892), .B(n22893), .Z(n22902) );
  XOR U27569 ( .A(n22898), .B(n22903), .Z(n22893) );
  XOR U27570 ( .A(n22897), .B(n22900), .Z(n22903) );
  IV U27571 ( .A(n22899), .Z(n22900) );
  NAND U27572 ( .A(n22904), .B(n22905), .Z(n22899) );
  OR U27573 ( .A(n22906), .B(n22907), .Z(n22905) );
  OR U27574 ( .A(n22908), .B(n22909), .Z(n22904) );
  NAND U27575 ( .A(n22910), .B(n22911), .Z(n22897) );
  OR U27576 ( .A(n22912), .B(n22913), .Z(n22911) );
  OR U27577 ( .A(n22914), .B(n22915), .Z(n22910) );
  NOR U27578 ( .A(n22916), .B(n22917), .Z(n22898) );
  ANDN U27579 ( .B(n22918), .A(n22919), .Z(n22892) );
  XNOR U27580 ( .A(n22885), .B(n22920), .Z(n22891) );
  XNOR U27581 ( .A(n22884), .B(n22886), .Z(n22920) );
  NAND U27582 ( .A(n22921), .B(n22922), .Z(n22886) );
  OR U27583 ( .A(n22923), .B(n22924), .Z(n22922) );
  OR U27584 ( .A(n22925), .B(n22926), .Z(n22921) );
  NAND U27585 ( .A(n22927), .B(n22928), .Z(n22884) );
  OR U27586 ( .A(n22929), .B(n22930), .Z(n22928) );
  OR U27587 ( .A(n22931), .B(n22932), .Z(n22927) );
  ANDN U27588 ( .B(n22933), .A(n22934), .Z(n22885) );
  IV U27589 ( .A(n22935), .Z(n22933) );
  ANDN U27590 ( .B(n22936), .A(n22937), .Z(n22877) );
  XOR U27591 ( .A(n22863), .B(n22938), .Z(n22875) );
  XOR U27592 ( .A(n22864), .B(n22865), .Z(n22938) );
  XOR U27593 ( .A(n22870), .B(n22939), .Z(n22865) );
  XOR U27594 ( .A(n22869), .B(n22872), .Z(n22939) );
  IV U27595 ( .A(n22871), .Z(n22872) );
  NAND U27596 ( .A(n22940), .B(n22941), .Z(n22871) );
  OR U27597 ( .A(n22942), .B(n22943), .Z(n22941) );
  OR U27598 ( .A(n22944), .B(n22945), .Z(n22940) );
  NAND U27599 ( .A(n22946), .B(n22947), .Z(n22869) );
  OR U27600 ( .A(n22948), .B(n22949), .Z(n22947) );
  OR U27601 ( .A(n22950), .B(n22951), .Z(n22946) );
  NOR U27602 ( .A(n22952), .B(n22953), .Z(n22870) );
  ANDN U27603 ( .B(n22954), .A(n22955), .Z(n22864) );
  IV U27604 ( .A(n22956), .Z(n22954) );
  XNOR U27605 ( .A(n22857), .B(n22957), .Z(n22863) );
  XNOR U27606 ( .A(n22856), .B(n22858), .Z(n22957) );
  NAND U27607 ( .A(n22958), .B(n22959), .Z(n22858) );
  OR U27608 ( .A(n22960), .B(n22961), .Z(n22959) );
  OR U27609 ( .A(n22962), .B(n22963), .Z(n22958) );
  NAND U27610 ( .A(n22964), .B(n22965), .Z(n22856) );
  OR U27611 ( .A(n22966), .B(n22967), .Z(n22965) );
  OR U27612 ( .A(n22968), .B(n22969), .Z(n22964) );
  ANDN U27613 ( .B(n22970), .A(n22971), .Z(n22857) );
  IV U27614 ( .A(n22972), .Z(n22970) );
  XNOR U27615 ( .A(n22937), .B(n22936), .Z(N28277) );
  XOR U27616 ( .A(n22956), .B(n22955), .Z(n22936) );
  XNOR U27617 ( .A(n22971), .B(n22972), .Z(n22955) );
  XNOR U27618 ( .A(n22966), .B(n22967), .Z(n22972) );
  XNOR U27619 ( .A(n22968), .B(n22969), .Z(n22967) );
  XNOR U27620 ( .A(y[700]), .B(x[700]), .Z(n22969) );
  XNOR U27621 ( .A(y[701]), .B(x[701]), .Z(n22968) );
  XNOR U27622 ( .A(y[699]), .B(x[699]), .Z(n22966) );
  XNOR U27623 ( .A(n22960), .B(n22961), .Z(n22971) );
  XNOR U27624 ( .A(y[696]), .B(x[696]), .Z(n22961) );
  XNOR U27625 ( .A(n22962), .B(n22963), .Z(n22960) );
  XNOR U27626 ( .A(y[697]), .B(x[697]), .Z(n22963) );
  XNOR U27627 ( .A(y[698]), .B(x[698]), .Z(n22962) );
  XNOR U27628 ( .A(n22953), .B(n22952), .Z(n22956) );
  XNOR U27629 ( .A(n22948), .B(n22949), .Z(n22952) );
  XNOR U27630 ( .A(y[693]), .B(x[693]), .Z(n22949) );
  XNOR U27631 ( .A(n22950), .B(n22951), .Z(n22948) );
  XNOR U27632 ( .A(y[694]), .B(x[694]), .Z(n22951) );
  XNOR U27633 ( .A(y[695]), .B(x[695]), .Z(n22950) );
  XNOR U27634 ( .A(n22942), .B(n22943), .Z(n22953) );
  XNOR U27635 ( .A(y[690]), .B(x[690]), .Z(n22943) );
  XNOR U27636 ( .A(n22944), .B(n22945), .Z(n22942) );
  XNOR U27637 ( .A(y[691]), .B(x[691]), .Z(n22945) );
  XNOR U27638 ( .A(y[692]), .B(x[692]), .Z(n22944) );
  XOR U27639 ( .A(n22918), .B(n22919), .Z(n22937) );
  XNOR U27640 ( .A(n22934), .B(n22935), .Z(n22919) );
  XNOR U27641 ( .A(n22929), .B(n22930), .Z(n22935) );
  XNOR U27642 ( .A(n22931), .B(n22932), .Z(n22930) );
  XNOR U27643 ( .A(y[688]), .B(x[688]), .Z(n22932) );
  XNOR U27644 ( .A(y[689]), .B(x[689]), .Z(n22931) );
  XNOR U27645 ( .A(y[687]), .B(x[687]), .Z(n22929) );
  XNOR U27646 ( .A(n22923), .B(n22924), .Z(n22934) );
  XNOR U27647 ( .A(y[684]), .B(x[684]), .Z(n22924) );
  XNOR U27648 ( .A(n22925), .B(n22926), .Z(n22923) );
  XNOR U27649 ( .A(y[685]), .B(x[685]), .Z(n22926) );
  XNOR U27650 ( .A(y[686]), .B(x[686]), .Z(n22925) );
  XOR U27651 ( .A(n22917), .B(n22916), .Z(n22918) );
  XNOR U27652 ( .A(n22912), .B(n22913), .Z(n22916) );
  XNOR U27653 ( .A(y[681]), .B(x[681]), .Z(n22913) );
  XNOR U27654 ( .A(n22914), .B(n22915), .Z(n22912) );
  XNOR U27655 ( .A(y[682]), .B(x[682]), .Z(n22915) );
  XNOR U27656 ( .A(y[683]), .B(x[683]), .Z(n22914) );
  XNOR U27657 ( .A(n22906), .B(n22907), .Z(n22917) );
  XNOR U27658 ( .A(y[678]), .B(x[678]), .Z(n22907) );
  XNOR U27659 ( .A(n22908), .B(n22909), .Z(n22906) );
  XNOR U27660 ( .A(y[679]), .B(x[679]), .Z(n22909) );
  XNOR U27661 ( .A(y[680]), .B(x[680]), .Z(n22908) );
  NAND U27662 ( .A(n22973), .B(n22974), .Z(N28269) );
  NANDN U27663 ( .A(n22975), .B(n22976), .Z(n22974) );
  OR U27664 ( .A(n22977), .B(n22978), .Z(n22976) );
  NAND U27665 ( .A(n22977), .B(n22978), .Z(n22973) );
  XOR U27666 ( .A(n22977), .B(n22979), .Z(N28268) );
  XNOR U27667 ( .A(n22975), .B(n22978), .Z(n22979) );
  AND U27668 ( .A(n22980), .B(n22981), .Z(n22978) );
  NANDN U27669 ( .A(n22982), .B(n22983), .Z(n22981) );
  NANDN U27670 ( .A(n22984), .B(n22985), .Z(n22983) );
  NANDN U27671 ( .A(n22985), .B(n22984), .Z(n22980) );
  NAND U27672 ( .A(n22986), .B(n22987), .Z(n22975) );
  NANDN U27673 ( .A(n22988), .B(n22989), .Z(n22987) );
  OR U27674 ( .A(n22990), .B(n22991), .Z(n22989) );
  NAND U27675 ( .A(n22991), .B(n22990), .Z(n22986) );
  AND U27676 ( .A(n22992), .B(n22993), .Z(n22977) );
  NANDN U27677 ( .A(n22994), .B(n22995), .Z(n22993) );
  NANDN U27678 ( .A(n22996), .B(n22997), .Z(n22995) );
  NANDN U27679 ( .A(n22997), .B(n22996), .Z(n22992) );
  XOR U27680 ( .A(n22991), .B(n22998), .Z(N28267) );
  XOR U27681 ( .A(n22988), .B(n22990), .Z(n22998) );
  XNOR U27682 ( .A(n22984), .B(n22999), .Z(n22990) );
  XNOR U27683 ( .A(n22982), .B(n22985), .Z(n22999) );
  NAND U27684 ( .A(n23000), .B(n23001), .Z(n22985) );
  NAND U27685 ( .A(n23002), .B(n23003), .Z(n23001) );
  OR U27686 ( .A(n23004), .B(n23005), .Z(n23002) );
  NANDN U27687 ( .A(n23006), .B(n23004), .Z(n23000) );
  IV U27688 ( .A(n23005), .Z(n23006) );
  NAND U27689 ( .A(n23007), .B(n23008), .Z(n22982) );
  NAND U27690 ( .A(n23009), .B(n23010), .Z(n23008) );
  NANDN U27691 ( .A(n23011), .B(n23012), .Z(n23009) );
  NANDN U27692 ( .A(n23012), .B(n23011), .Z(n23007) );
  AND U27693 ( .A(n23013), .B(n23014), .Z(n22984) );
  NAND U27694 ( .A(n23015), .B(n23016), .Z(n23014) );
  OR U27695 ( .A(n23017), .B(n23018), .Z(n23015) );
  NANDN U27696 ( .A(n23019), .B(n23017), .Z(n23013) );
  NAND U27697 ( .A(n23020), .B(n23021), .Z(n22988) );
  NANDN U27698 ( .A(n23022), .B(n23023), .Z(n23021) );
  OR U27699 ( .A(n23024), .B(n23025), .Z(n23023) );
  NANDN U27700 ( .A(n23026), .B(n23024), .Z(n23020) );
  IV U27701 ( .A(n23025), .Z(n23026) );
  XNOR U27702 ( .A(n22996), .B(n23027), .Z(n22991) );
  XNOR U27703 ( .A(n22994), .B(n22997), .Z(n23027) );
  NAND U27704 ( .A(n23028), .B(n23029), .Z(n22997) );
  NAND U27705 ( .A(n23030), .B(n23031), .Z(n23029) );
  OR U27706 ( .A(n23032), .B(n23033), .Z(n23030) );
  NANDN U27707 ( .A(n23034), .B(n23032), .Z(n23028) );
  IV U27708 ( .A(n23033), .Z(n23034) );
  NAND U27709 ( .A(n23035), .B(n23036), .Z(n22994) );
  NAND U27710 ( .A(n23037), .B(n23038), .Z(n23036) );
  NANDN U27711 ( .A(n23039), .B(n23040), .Z(n23037) );
  NANDN U27712 ( .A(n23040), .B(n23039), .Z(n23035) );
  AND U27713 ( .A(n23041), .B(n23042), .Z(n22996) );
  NAND U27714 ( .A(n23043), .B(n23044), .Z(n23042) );
  OR U27715 ( .A(n23045), .B(n23046), .Z(n23043) );
  NANDN U27716 ( .A(n23047), .B(n23045), .Z(n23041) );
  XNOR U27717 ( .A(n23022), .B(n23048), .Z(N28266) );
  XOR U27718 ( .A(n23024), .B(n23025), .Z(n23048) );
  XNOR U27719 ( .A(n23038), .B(n23049), .Z(n23025) );
  XOR U27720 ( .A(n23039), .B(n23040), .Z(n23049) );
  XOR U27721 ( .A(n23045), .B(n23050), .Z(n23040) );
  XOR U27722 ( .A(n23044), .B(n23047), .Z(n23050) );
  IV U27723 ( .A(n23046), .Z(n23047) );
  NAND U27724 ( .A(n23051), .B(n23052), .Z(n23046) );
  OR U27725 ( .A(n23053), .B(n23054), .Z(n23052) );
  OR U27726 ( .A(n23055), .B(n23056), .Z(n23051) );
  NAND U27727 ( .A(n23057), .B(n23058), .Z(n23044) );
  OR U27728 ( .A(n23059), .B(n23060), .Z(n23058) );
  OR U27729 ( .A(n23061), .B(n23062), .Z(n23057) );
  NOR U27730 ( .A(n23063), .B(n23064), .Z(n23045) );
  ANDN U27731 ( .B(n23065), .A(n23066), .Z(n23039) );
  XNOR U27732 ( .A(n23032), .B(n23067), .Z(n23038) );
  XNOR U27733 ( .A(n23031), .B(n23033), .Z(n23067) );
  NAND U27734 ( .A(n23068), .B(n23069), .Z(n23033) );
  OR U27735 ( .A(n23070), .B(n23071), .Z(n23069) );
  OR U27736 ( .A(n23072), .B(n23073), .Z(n23068) );
  NAND U27737 ( .A(n23074), .B(n23075), .Z(n23031) );
  OR U27738 ( .A(n23076), .B(n23077), .Z(n23075) );
  OR U27739 ( .A(n23078), .B(n23079), .Z(n23074) );
  ANDN U27740 ( .B(n23080), .A(n23081), .Z(n23032) );
  IV U27741 ( .A(n23082), .Z(n23080) );
  ANDN U27742 ( .B(n23083), .A(n23084), .Z(n23024) );
  XOR U27743 ( .A(n23010), .B(n23085), .Z(n23022) );
  XOR U27744 ( .A(n23011), .B(n23012), .Z(n23085) );
  XOR U27745 ( .A(n23017), .B(n23086), .Z(n23012) );
  XOR U27746 ( .A(n23016), .B(n23019), .Z(n23086) );
  IV U27747 ( .A(n23018), .Z(n23019) );
  NAND U27748 ( .A(n23087), .B(n23088), .Z(n23018) );
  OR U27749 ( .A(n23089), .B(n23090), .Z(n23088) );
  OR U27750 ( .A(n23091), .B(n23092), .Z(n23087) );
  NAND U27751 ( .A(n23093), .B(n23094), .Z(n23016) );
  OR U27752 ( .A(n23095), .B(n23096), .Z(n23094) );
  OR U27753 ( .A(n23097), .B(n23098), .Z(n23093) );
  NOR U27754 ( .A(n23099), .B(n23100), .Z(n23017) );
  ANDN U27755 ( .B(n23101), .A(n23102), .Z(n23011) );
  IV U27756 ( .A(n23103), .Z(n23101) );
  XNOR U27757 ( .A(n23004), .B(n23104), .Z(n23010) );
  XNOR U27758 ( .A(n23003), .B(n23005), .Z(n23104) );
  NAND U27759 ( .A(n23105), .B(n23106), .Z(n23005) );
  OR U27760 ( .A(n23107), .B(n23108), .Z(n23106) );
  OR U27761 ( .A(n23109), .B(n23110), .Z(n23105) );
  NAND U27762 ( .A(n23111), .B(n23112), .Z(n23003) );
  OR U27763 ( .A(n23113), .B(n23114), .Z(n23112) );
  OR U27764 ( .A(n23115), .B(n23116), .Z(n23111) );
  ANDN U27765 ( .B(n23117), .A(n23118), .Z(n23004) );
  IV U27766 ( .A(n23119), .Z(n23117) );
  XNOR U27767 ( .A(n23084), .B(n23083), .Z(N28265) );
  XOR U27768 ( .A(n23103), .B(n23102), .Z(n23083) );
  XNOR U27769 ( .A(n23118), .B(n23119), .Z(n23102) );
  XNOR U27770 ( .A(n23113), .B(n23114), .Z(n23119) );
  XNOR U27771 ( .A(n23115), .B(n23116), .Z(n23114) );
  XNOR U27772 ( .A(y[676]), .B(x[676]), .Z(n23116) );
  XNOR U27773 ( .A(y[677]), .B(x[677]), .Z(n23115) );
  XNOR U27774 ( .A(y[675]), .B(x[675]), .Z(n23113) );
  XNOR U27775 ( .A(n23107), .B(n23108), .Z(n23118) );
  XNOR U27776 ( .A(y[672]), .B(x[672]), .Z(n23108) );
  XNOR U27777 ( .A(n23109), .B(n23110), .Z(n23107) );
  XNOR U27778 ( .A(y[673]), .B(x[673]), .Z(n23110) );
  XNOR U27779 ( .A(y[674]), .B(x[674]), .Z(n23109) );
  XNOR U27780 ( .A(n23100), .B(n23099), .Z(n23103) );
  XNOR U27781 ( .A(n23095), .B(n23096), .Z(n23099) );
  XNOR U27782 ( .A(y[669]), .B(x[669]), .Z(n23096) );
  XNOR U27783 ( .A(n23097), .B(n23098), .Z(n23095) );
  XNOR U27784 ( .A(y[670]), .B(x[670]), .Z(n23098) );
  XNOR U27785 ( .A(y[671]), .B(x[671]), .Z(n23097) );
  XNOR U27786 ( .A(n23089), .B(n23090), .Z(n23100) );
  XNOR U27787 ( .A(y[666]), .B(x[666]), .Z(n23090) );
  XNOR U27788 ( .A(n23091), .B(n23092), .Z(n23089) );
  XNOR U27789 ( .A(y[667]), .B(x[667]), .Z(n23092) );
  XNOR U27790 ( .A(y[668]), .B(x[668]), .Z(n23091) );
  XOR U27791 ( .A(n23065), .B(n23066), .Z(n23084) );
  XNOR U27792 ( .A(n23081), .B(n23082), .Z(n23066) );
  XNOR U27793 ( .A(n23076), .B(n23077), .Z(n23082) );
  XNOR U27794 ( .A(n23078), .B(n23079), .Z(n23077) );
  XNOR U27795 ( .A(y[664]), .B(x[664]), .Z(n23079) );
  XNOR U27796 ( .A(y[665]), .B(x[665]), .Z(n23078) );
  XNOR U27797 ( .A(y[663]), .B(x[663]), .Z(n23076) );
  XNOR U27798 ( .A(n23070), .B(n23071), .Z(n23081) );
  XNOR U27799 ( .A(y[660]), .B(x[660]), .Z(n23071) );
  XNOR U27800 ( .A(n23072), .B(n23073), .Z(n23070) );
  XNOR U27801 ( .A(y[661]), .B(x[661]), .Z(n23073) );
  XNOR U27802 ( .A(y[662]), .B(x[662]), .Z(n23072) );
  XOR U27803 ( .A(n23064), .B(n23063), .Z(n23065) );
  XNOR U27804 ( .A(n23059), .B(n23060), .Z(n23063) );
  XNOR U27805 ( .A(y[657]), .B(x[657]), .Z(n23060) );
  XNOR U27806 ( .A(n23061), .B(n23062), .Z(n23059) );
  XNOR U27807 ( .A(y[658]), .B(x[658]), .Z(n23062) );
  XNOR U27808 ( .A(y[659]), .B(x[659]), .Z(n23061) );
  XNOR U27809 ( .A(n23053), .B(n23054), .Z(n23064) );
  XNOR U27810 ( .A(y[654]), .B(x[654]), .Z(n23054) );
  XNOR U27811 ( .A(n23055), .B(n23056), .Z(n23053) );
  XNOR U27812 ( .A(y[655]), .B(x[655]), .Z(n23056) );
  XNOR U27813 ( .A(y[656]), .B(x[656]), .Z(n23055) );
  NAND U27814 ( .A(n23120), .B(n23121), .Z(N28257) );
  NANDN U27815 ( .A(n23122), .B(n23123), .Z(n23121) );
  OR U27816 ( .A(n23124), .B(n23125), .Z(n23123) );
  NAND U27817 ( .A(n23124), .B(n23125), .Z(n23120) );
  XOR U27818 ( .A(n23124), .B(n23126), .Z(N28256) );
  XNOR U27819 ( .A(n23122), .B(n23125), .Z(n23126) );
  AND U27820 ( .A(n23127), .B(n23128), .Z(n23125) );
  NANDN U27821 ( .A(n23129), .B(n23130), .Z(n23128) );
  NANDN U27822 ( .A(n23131), .B(n23132), .Z(n23130) );
  NANDN U27823 ( .A(n23132), .B(n23131), .Z(n23127) );
  NAND U27824 ( .A(n23133), .B(n23134), .Z(n23122) );
  NANDN U27825 ( .A(n23135), .B(n23136), .Z(n23134) );
  OR U27826 ( .A(n23137), .B(n23138), .Z(n23136) );
  NAND U27827 ( .A(n23138), .B(n23137), .Z(n23133) );
  AND U27828 ( .A(n23139), .B(n23140), .Z(n23124) );
  NANDN U27829 ( .A(n23141), .B(n23142), .Z(n23140) );
  NANDN U27830 ( .A(n23143), .B(n23144), .Z(n23142) );
  NANDN U27831 ( .A(n23144), .B(n23143), .Z(n23139) );
  XOR U27832 ( .A(n23138), .B(n23145), .Z(N28255) );
  XOR U27833 ( .A(n23135), .B(n23137), .Z(n23145) );
  XNOR U27834 ( .A(n23131), .B(n23146), .Z(n23137) );
  XNOR U27835 ( .A(n23129), .B(n23132), .Z(n23146) );
  NAND U27836 ( .A(n23147), .B(n23148), .Z(n23132) );
  NAND U27837 ( .A(n23149), .B(n23150), .Z(n23148) );
  OR U27838 ( .A(n23151), .B(n23152), .Z(n23149) );
  NANDN U27839 ( .A(n23153), .B(n23151), .Z(n23147) );
  IV U27840 ( .A(n23152), .Z(n23153) );
  NAND U27841 ( .A(n23154), .B(n23155), .Z(n23129) );
  NAND U27842 ( .A(n23156), .B(n23157), .Z(n23155) );
  NANDN U27843 ( .A(n23158), .B(n23159), .Z(n23156) );
  NANDN U27844 ( .A(n23159), .B(n23158), .Z(n23154) );
  AND U27845 ( .A(n23160), .B(n23161), .Z(n23131) );
  NAND U27846 ( .A(n23162), .B(n23163), .Z(n23161) );
  OR U27847 ( .A(n23164), .B(n23165), .Z(n23162) );
  NANDN U27848 ( .A(n23166), .B(n23164), .Z(n23160) );
  NAND U27849 ( .A(n23167), .B(n23168), .Z(n23135) );
  NANDN U27850 ( .A(n23169), .B(n23170), .Z(n23168) );
  OR U27851 ( .A(n23171), .B(n23172), .Z(n23170) );
  NANDN U27852 ( .A(n23173), .B(n23171), .Z(n23167) );
  IV U27853 ( .A(n23172), .Z(n23173) );
  XNOR U27854 ( .A(n23143), .B(n23174), .Z(n23138) );
  XNOR U27855 ( .A(n23141), .B(n23144), .Z(n23174) );
  NAND U27856 ( .A(n23175), .B(n23176), .Z(n23144) );
  NAND U27857 ( .A(n23177), .B(n23178), .Z(n23176) );
  OR U27858 ( .A(n23179), .B(n23180), .Z(n23177) );
  NANDN U27859 ( .A(n23181), .B(n23179), .Z(n23175) );
  IV U27860 ( .A(n23180), .Z(n23181) );
  NAND U27861 ( .A(n23182), .B(n23183), .Z(n23141) );
  NAND U27862 ( .A(n23184), .B(n23185), .Z(n23183) );
  NANDN U27863 ( .A(n23186), .B(n23187), .Z(n23184) );
  NANDN U27864 ( .A(n23187), .B(n23186), .Z(n23182) );
  AND U27865 ( .A(n23188), .B(n23189), .Z(n23143) );
  NAND U27866 ( .A(n23190), .B(n23191), .Z(n23189) );
  OR U27867 ( .A(n23192), .B(n23193), .Z(n23190) );
  NANDN U27868 ( .A(n23194), .B(n23192), .Z(n23188) );
  XNOR U27869 ( .A(n23169), .B(n23195), .Z(N28254) );
  XOR U27870 ( .A(n23171), .B(n23172), .Z(n23195) );
  XNOR U27871 ( .A(n23185), .B(n23196), .Z(n23172) );
  XOR U27872 ( .A(n23186), .B(n23187), .Z(n23196) );
  XOR U27873 ( .A(n23192), .B(n23197), .Z(n23187) );
  XOR U27874 ( .A(n23191), .B(n23194), .Z(n23197) );
  IV U27875 ( .A(n23193), .Z(n23194) );
  NAND U27876 ( .A(n23198), .B(n23199), .Z(n23193) );
  OR U27877 ( .A(n23200), .B(n23201), .Z(n23199) );
  OR U27878 ( .A(n23202), .B(n23203), .Z(n23198) );
  NAND U27879 ( .A(n23204), .B(n23205), .Z(n23191) );
  OR U27880 ( .A(n23206), .B(n23207), .Z(n23205) );
  OR U27881 ( .A(n23208), .B(n23209), .Z(n23204) );
  NOR U27882 ( .A(n23210), .B(n23211), .Z(n23192) );
  ANDN U27883 ( .B(n23212), .A(n23213), .Z(n23186) );
  XNOR U27884 ( .A(n23179), .B(n23214), .Z(n23185) );
  XNOR U27885 ( .A(n23178), .B(n23180), .Z(n23214) );
  NAND U27886 ( .A(n23215), .B(n23216), .Z(n23180) );
  OR U27887 ( .A(n23217), .B(n23218), .Z(n23216) );
  OR U27888 ( .A(n23219), .B(n23220), .Z(n23215) );
  NAND U27889 ( .A(n23221), .B(n23222), .Z(n23178) );
  OR U27890 ( .A(n23223), .B(n23224), .Z(n23222) );
  OR U27891 ( .A(n23225), .B(n23226), .Z(n23221) );
  ANDN U27892 ( .B(n23227), .A(n23228), .Z(n23179) );
  IV U27893 ( .A(n23229), .Z(n23227) );
  ANDN U27894 ( .B(n23230), .A(n23231), .Z(n23171) );
  XOR U27895 ( .A(n23157), .B(n23232), .Z(n23169) );
  XOR U27896 ( .A(n23158), .B(n23159), .Z(n23232) );
  XOR U27897 ( .A(n23164), .B(n23233), .Z(n23159) );
  XOR U27898 ( .A(n23163), .B(n23166), .Z(n23233) );
  IV U27899 ( .A(n23165), .Z(n23166) );
  NAND U27900 ( .A(n23234), .B(n23235), .Z(n23165) );
  OR U27901 ( .A(n23236), .B(n23237), .Z(n23235) );
  OR U27902 ( .A(n23238), .B(n23239), .Z(n23234) );
  NAND U27903 ( .A(n23240), .B(n23241), .Z(n23163) );
  OR U27904 ( .A(n23242), .B(n23243), .Z(n23241) );
  OR U27905 ( .A(n23244), .B(n23245), .Z(n23240) );
  NOR U27906 ( .A(n23246), .B(n23247), .Z(n23164) );
  ANDN U27907 ( .B(n23248), .A(n23249), .Z(n23158) );
  IV U27908 ( .A(n23250), .Z(n23248) );
  XNOR U27909 ( .A(n23151), .B(n23251), .Z(n23157) );
  XNOR U27910 ( .A(n23150), .B(n23152), .Z(n23251) );
  NAND U27911 ( .A(n23252), .B(n23253), .Z(n23152) );
  OR U27912 ( .A(n23254), .B(n23255), .Z(n23253) );
  OR U27913 ( .A(n23256), .B(n23257), .Z(n23252) );
  NAND U27914 ( .A(n23258), .B(n23259), .Z(n23150) );
  OR U27915 ( .A(n23260), .B(n23261), .Z(n23259) );
  OR U27916 ( .A(n23262), .B(n23263), .Z(n23258) );
  ANDN U27917 ( .B(n23264), .A(n23265), .Z(n23151) );
  IV U27918 ( .A(n23266), .Z(n23264) );
  XNOR U27919 ( .A(n23231), .B(n23230), .Z(N28253) );
  XOR U27920 ( .A(n23250), .B(n23249), .Z(n23230) );
  XNOR U27921 ( .A(n23265), .B(n23266), .Z(n23249) );
  XNOR U27922 ( .A(n23260), .B(n23261), .Z(n23266) );
  XNOR U27923 ( .A(n23262), .B(n23263), .Z(n23261) );
  XNOR U27924 ( .A(y[652]), .B(x[652]), .Z(n23263) );
  XNOR U27925 ( .A(y[653]), .B(x[653]), .Z(n23262) );
  XNOR U27926 ( .A(y[651]), .B(x[651]), .Z(n23260) );
  XNOR U27927 ( .A(n23254), .B(n23255), .Z(n23265) );
  XNOR U27928 ( .A(y[648]), .B(x[648]), .Z(n23255) );
  XNOR U27929 ( .A(n23256), .B(n23257), .Z(n23254) );
  XNOR U27930 ( .A(y[649]), .B(x[649]), .Z(n23257) );
  XNOR U27931 ( .A(y[650]), .B(x[650]), .Z(n23256) );
  XNOR U27932 ( .A(n23247), .B(n23246), .Z(n23250) );
  XNOR U27933 ( .A(n23242), .B(n23243), .Z(n23246) );
  XNOR U27934 ( .A(y[645]), .B(x[645]), .Z(n23243) );
  XNOR U27935 ( .A(n23244), .B(n23245), .Z(n23242) );
  XNOR U27936 ( .A(y[646]), .B(x[646]), .Z(n23245) );
  XNOR U27937 ( .A(y[647]), .B(x[647]), .Z(n23244) );
  XNOR U27938 ( .A(n23236), .B(n23237), .Z(n23247) );
  XNOR U27939 ( .A(y[642]), .B(x[642]), .Z(n23237) );
  XNOR U27940 ( .A(n23238), .B(n23239), .Z(n23236) );
  XNOR U27941 ( .A(y[643]), .B(x[643]), .Z(n23239) );
  XNOR U27942 ( .A(y[644]), .B(x[644]), .Z(n23238) );
  XOR U27943 ( .A(n23212), .B(n23213), .Z(n23231) );
  XNOR U27944 ( .A(n23228), .B(n23229), .Z(n23213) );
  XNOR U27945 ( .A(n23223), .B(n23224), .Z(n23229) );
  XNOR U27946 ( .A(n23225), .B(n23226), .Z(n23224) );
  XNOR U27947 ( .A(y[640]), .B(x[640]), .Z(n23226) );
  XNOR U27948 ( .A(y[641]), .B(x[641]), .Z(n23225) );
  XNOR U27949 ( .A(y[639]), .B(x[639]), .Z(n23223) );
  XNOR U27950 ( .A(n23217), .B(n23218), .Z(n23228) );
  XNOR U27951 ( .A(y[636]), .B(x[636]), .Z(n23218) );
  XNOR U27952 ( .A(n23219), .B(n23220), .Z(n23217) );
  XNOR U27953 ( .A(y[637]), .B(x[637]), .Z(n23220) );
  XNOR U27954 ( .A(y[638]), .B(x[638]), .Z(n23219) );
  XOR U27955 ( .A(n23211), .B(n23210), .Z(n23212) );
  XNOR U27956 ( .A(n23206), .B(n23207), .Z(n23210) );
  XNOR U27957 ( .A(y[633]), .B(x[633]), .Z(n23207) );
  XNOR U27958 ( .A(n23208), .B(n23209), .Z(n23206) );
  XNOR U27959 ( .A(y[634]), .B(x[634]), .Z(n23209) );
  XNOR U27960 ( .A(y[635]), .B(x[635]), .Z(n23208) );
  XNOR U27961 ( .A(n23200), .B(n23201), .Z(n23211) );
  XNOR U27962 ( .A(y[630]), .B(x[630]), .Z(n23201) );
  XNOR U27963 ( .A(n23202), .B(n23203), .Z(n23200) );
  XNOR U27964 ( .A(y[631]), .B(x[631]), .Z(n23203) );
  XNOR U27965 ( .A(y[632]), .B(x[632]), .Z(n23202) );
  NAND U27966 ( .A(n23267), .B(n23268), .Z(N28245) );
  NANDN U27967 ( .A(n23269), .B(n23270), .Z(n23268) );
  OR U27968 ( .A(n23271), .B(n23272), .Z(n23270) );
  NAND U27969 ( .A(n23271), .B(n23272), .Z(n23267) );
  XOR U27970 ( .A(n23271), .B(n23273), .Z(N28244) );
  XNOR U27971 ( .A(n23269), .B(n23272), .Z(n23273) );
  AND U27972 ( .A(n23274), .B(n23275), .Z(n23272) );
  NANDN U27973 ( .A(n23276), .B(n23277), .Z(n23275) );
  NANDN U27974 ( .A(n23278), .B(n23279), .Z(n23277) );
  NANDN U27975 ( .A(n23279), .B(n23278), .Z(n23274) );
  NAND U27976 ( .A(n23280), .B(n23281), .Z(n23269) );
  NANDN U27977 ( .A(n23282), .B(n23283), .Z(n23281) );
  OR U27978 ( .A(n23284), .B(n23285), .Z(n23283) );
  NAND U27979 ( .A(n23285), .B(n23284), .Z(n23280) );
  AND U27980 ( .A(n23286), .B(n23287), .Z(n23271) );
  NANDN U27981 ( .A(n23288), .B(n23289), .Z(n23287) );
  NANDN U27982 ( .A(n23290), .B(n23291), .Z(n23289) );
  NANDN U27983 ( .A(n23291), .B(n23290), .Z(n23286) );
  XOR U27984 ( .A(n23285), .B(n23292), .Z(N28243) );
  XOR U27985 ( .A(n23282), .B(n23284), .Z(n23292) );
  XNOR U27986 ( .A(n23278), .B(n23293), .Z(n23284) );
  XNOR U27987 ( .A(n23276), .B(n23279), .Z(n23293) );
  NAND U27988 ( .A(n23294), .B(n23295), .Z(n23279) );
  NAND U27989 ( .A(n23296), .B(n23297), .Z(n23295) );
  OR U27990 ( .A(n23298), .B(n23299), .Z(n23296) );
  NANDN U27991 ( .A(n23300), .B(n23298), .Z(n23294) );
  IV U27992 ( .A(n23299), .Z(n23300) );
  NAND U27993 ( .A(n23301), .B(n23302), .Z(n23276) );
  NAND U27994 ( .A(n23303), .B(n23304), .Z(n23302) );
  NANDN U27995 ( .A(n23305), .B(n23306), .Z(n23303) );
  NANDN U27996 ( .A(n23306), .B(n23305), .Z(n23301) );
  AND U27997 ( .A(n23307), .B(n23308), .Z(n23278) );
  NAND U27998 ( .A(n23309), .B(n23310), .Z(n23308) );
  OR U27999 ( .A(n23311), .B(n23312), .Z(n23309) );
  NANDN U28000 ( .A(n23313), .B(n23311), .Z(n23307) );
  NAND U28001 ( .A(n23314), .B(n23315), .Z(n23282) );
  NANDN U28002 ( .A(n23316), .B(n23317), .Z(n23315) );
  OR U28003 ( .A(n23318), .B(n23319), .Z(n23317) );
  NANDN U28004 ( .A(n23320), .B(n23318), .Z(n23314) );
  IV U28005 ( .A(n23319), .Z(n23320) );
  XNOR U28006 ( .A(n23290), .B(n23321), .Z(n23285) );
  XNOR U28007 ( .A(n23288), .B(n23291), .Z(n23321) );
  NAND U28008 ( .A(n23322), .B(n23323), .Z(n23291) );
  NAND U28009 ( .A(n23324), .B(n23325), .Z(n23323) );
  OR U28010 ( .A(n23326), .B(n23327), .Z(n23324) );
  NANDN U28011 ( .A(n23328), .B(n23326), .Z(n23322) );
  IV U28012 ( .A(n23327), .Z(n23328) );
  NAND U28013 ( .A(n23329), .B(n23330), .Z(n23288) );
  NAND U28014 ( .A(n23331), .B(n23332), .Z(n23330) );
  NANDN U28015 ( .A(n23333), .B(n23334), .Z(n23331) );
  NANDN U28016 ( .A(n23334), .B(n23333), .Z(n23329) );
  AND U28017 ( .A(n23335), .B(n23336), .Z(n23290) );
  NAND U28018 ( .A(n23337), .B(n23338), .Z(n23336) );
  OR U28019 ( .A(n23339), .B(n23340), .Z(n23337) );
  NANDN U28020 ( .A(n23341), .B(n23339), .Z(n23335) );
  XNOR U28021 ( .A(n23316), .B(n23342), .Z(N28242) );
  XOR U28022 ( .A(n23318), .B(n23319), .Z(n23342) );
  XNOR U28023 ( .A(n23332), .B(n23343), .Z(n23319) );
  XOR U28024 ( .A(n23333), .B(n23334), .Z(n23343) );
  XOR U28025 ( .A(n23339), .B(n23344), .Z(n23334) );
  XOR U28026 ( .A(n23338), .B(n23341), .Z(n23344) );
  IV U28027 ( .A(n23340), .Z(n23341) );
  NAND U28028 ( .A(n23345), .B(n23346), .Z(n23340) );
  OR U28029 ( .A(n23347), .B(n23348), .Z(n23346) );
  OR U28030 ( .A(n23349), .B(n23350), .Z(n23345) );
  NAND U28031 ( .A(n23351), .B(n23352), .Z(n23338) );
  OR U28032 ( .A(n23353), .B(n23354), .Z(n23352) );
  OR U28033 ( .A(n23355), .B(n23356), .Z(n23351) );
  NOR U28034 ( .A(n23357), .B(n23358), .Z(n23339) );
  ANDN U28035 ( .B(n23359), .A(n23360), .Z(n23333) );
  XNOR U28036 ( .A(n23326), .B(n23361), .Z(n23332) );
  XNOR U28037 ( .A(n23325), .B(n23327), .Z(n23361) );
  NAND U28038 ( .A(n23362), .B(n23363), .Z(n23327) );
  OR U28039 ( .A(n23364), .B(n23365), .Z(n23363) );
  OR U28040 ( .A(n23366), .B(n23367), .Z(n23362) );
  NAND U28041 ( .A(n23368), .B(n23369), .Z(n23325) );
  OR U28042 ( .A(n23370), .B(n23371), .Z(n23369) );
  OR U28043 ( .A(n23372), .B(n23373), .Z(n23368) );
  ANDN U28044 ( .B(n23374), .A(n23375), .Z(n23326) );
  IV U28045 ( .A(n23376), .Z(n23374) );
  ANDN U28046 ( .B(n23377), .A(n23378), .Z(n23318) );
  XOR U28047 ( .A(n23304), .B(n23379), .Z(n23316) );
  XOR U28048 ( .A(n23305), .B(n23306), .Z(n23379) );
  XOR U28049 ( .A(n23311), .B(n23380), .Z(n23306) );
  XOR U28050 ( .A(n23310), .B(n23313), .Z(n23380) );
  IV U28051 ( .A(n23312), .Z(n23313) );
  NAND U28052 ( .A(n23381), .B(n23382), .Z(n23312) );
  OR U28053 ( .A(n23383), .B(n23384), .Z(n23382) );
  OR U28054 ( .A(n23385), .B(n23386), .Z(n23381) );
  NAND U28055 ( .A(n23387), .B(n23388), .Z(n23310) );
  OR U28056 ( .A(n23389), .B(n23390), .Z(n23388) );
  OR U28057 ( .A(n23391), .B(n23392), .Z(n23387) );
  NOR U28058 ( .A(n23393), .B(n23394), .Z(n23311) );
  ANDN U28059 ( .B(n23395), .A(n23396), .Z(n23305) );
  IV U28060 ( .A(n23397), .Z(n23395) );
  XNOR U28061 ( .A(n23298), .B(n23398), .Z(n23304) );
  XNOR U28062 ( .A(n23297), .B(n23299), .Z(n23398) );
  NAND U28063 ( .A(n23399), .B(n23400), .Z(n23299) );
  OR U28064 ( .A(n23401), .B(n23402), .Z(n23400) );
  OR U28065 ( .A(n23403), .B(n23404), .Z(n23399) );
  NAND U28066 ( .A(n23405), .B(n23406), .Z(n23297) );
  OR U28067 ( .A(n23407), .B(n23408), .Z(n23406) );
  OR U28068 ( .A(n23409), .B(n23410), .Z(n23405) );
  ANDN U28069 ( .B(n23411), .A(n23412), .Z(n23298) );
  IV U28070 ( .A(n23413), .Z(n23411) );
  XNOR U28071 ( .A(n23378), .B(n23377), .Z(N28241) );
  XOR U28072 ( .A(n23397), .B(n23396), .Z(n23377) );
  XNOR U28073 ( .A(n23412), .B(n23413), .Z(n23396) );
  XNOR U28074 ( .A(n23407), .B(n23408), .Z(n23413) );
  XNOR U28075 ( .A(n23409), .B(n23410), .Z(n23408) );
  XNOR U28076 ( .A(y[628]), .B(x[628]), .Z(n23410) );
  XNOR U28077 ( .A(y[629]), .B(x[629]), .Z(n23409) );
  XNOR U28078 ( .A(y[627]), .B(x[627]), .Z(n23407) );
  XNOR U28079 ( .A(n23401), .B(n23402), .Z(n23412) );
  XNOR U28080 ( .A(y[624]), .B(x[624]), .Z(n23402) );
  XNOR U28081 ( .A(n23403), .B(n23404), .Z(n23401) );
  XNOR U28082 ( .A(y[625]), .B(x[625]), .Z(n23404) );
  XNOR U28083 ( .A(y[626]), .B(x[626]), .Z(n23403) );
  XNOR U28084 ( .A(n23394), .B(n23393), .Z(n23397) );
  XNOR U28085 ( .A(n23389), .B(n23390), .Z(n23393) );
  XNOR U28086 ( .A(y[621]), .B(x[621]), .Z(n23390) );
  XNOR U28087 ( .A(n23391), .B(n23392), .Z(n23389) );
  XNOR U28088 ( .A(y[622]), .B(x[622]), .Z(n23392) );
  XNOR U28089 ( .A(y[623]), .B(x[623]), .Z(n23391) );
  XNOR U28090 ( .A(n23383), .B(n23384), .Z(n23394) );
  XNOR U28091 ( .A(y[618]), .B(x[618]), .Z(n23384) );
  XNOR U28092 ( .A(n23385), .B(n23386), .Z(n23383) );
  XNOR U28093 ( .A(y[619]), .B(x[619]), .Z(n23386) );
  XNOR U28094 ( .A(y[620]), .B(x[620]), .Z(n23385) );
  XOR U28095 ( .A(n23359), .B(n23360), .Z(n23378) );
  XNOR U28096 ( .A(n23375), .B(n23376), .Z(n23360) );
  XNOR U28097 ( .A(n23370), .B(n23371), .Z(n23376) );
  XNOR U28098 ( .A(n23372), .B(n23373), .Z(n23371) );
  XNOR U28099 ( .A(y[616]), .B(x[616]), .Z(n23373) );
  XNOR U28100 ( .A(y[617]), .B(x[617]), .Z(n23372) );
  XNOR U28101 ( .A(y[615]), .B(x[615]), .Z(n23370) );
  XNOR U28102 ( .A(n23364), .B(n23365), .Z(n23375) );
  XNOR U28103 ( .A(y[612]), .B(x[612]), .Z(n23365) );
  XNOR U28104 ( .A(n23366), .B(n23367), .Z(n23364) );
  XNOR U28105 ( .A(y[613]), .B(x[613]), .Z(n23367) );
  XNOR U28106 ( .A(y[614]), .B(x[614]), .Z(n23366) );
  XOR U28107 ( .A(n23358), .B(n23357), .Z(n23359) );
  XNOR U28108 ( .A(n23353), .B(n23354), .Z(n23357) );
  XNOR U28109 ( .A(y[609]), .B(x[609]), .Z(n23354) );
  XNOR U28110 ( .A(n23355), .B(n23356), .Z(n23353) );
  XNOR U28111 ( .A(y[610]), .B(x[610]), .Z(n23356) );
  XNOR U28112 ( .A(y[611]), .B(x[611]), .Z(n23355) );
  XNOR U28113 ( .A(n23347), .B(n23348), .Z(n23358) );
  XNOR U28114 ( .A(y[606]), .B(x[606]), .Z(n23348) );
  XNOR U28115 ( .A(n23349), .B(n23350), .Z(n23347) );
  XNOR U28116 ( .A(y[607]), .B(x[607]), .Z(n23350) );
  XNOR U28117 ( .A(y[608]), .B(x[608]), .Z(n23349) );
  NAND U28118 ( .A(n23414), .B(n23415), .Z(N28233) );
  NANDN U28119 ( .A(n23416), .B(n23417), .Z(n23415) );
  OR U28120 ( .A(n23418), .B(n23419), .Z(n23417) );
  NAND U28121 ( .A(n23418), .B(n23419), .Z(n23414) );
  XOR U28122 ( .A(n23418), .B(n23420), .Z(N28232) );
  XNOR U28123 ( .A(n23416), .B(n23419), .Z(n23420) );
  AND U28124 ( .A(n23421), .B(n23422), .Z(n23419) );
  NANDN U28125 ( .A(n23423), .B(n23424), .Z(n23422) );
  NANDN U28126 ( .A(n23425), .B(n23426), .Z(n23424) );
  NANDN U28127 ( .A(n23426), .B(n23425), .Z(n23421) );
  NAND U28128 ( .A(n23427), .B(n23428), .Z(n23416) );
  NANDN U28129 ( .A(n23429), .B(n23430), .Z(n23428) );
  OR U28130 ( .A(n23431), .B(n23432), .Z(n23430) );
  NAND U28131 ( .A(n23432), .B(n23431), .Z(n23427) );
  AND U28132 ( .A(n23433), .B(n23434), .Z(n23418) );
  NANDN U28133 ( .A(n23435), .B(n23436), .Z(n23434) );
  NANDN U28134 ( .A(n23437), .B(n23438), .Z(n23436) );
  NANDN U28135 ( .A(n23438), .B(n23437), .Z(n23433) );
  XOR U28136 ( .A(n23432), .B(n23439), .Z(N28231) );
  XOR U28137 ( .A(n23429), .B(n23431), .Z(n23439) );
  XNOR U28138 ( .A(n23425), .B(n23440), .Z(n23431) );
  XNOR U28139 ( .A(n23423), .B(n23426), .Z(n23440) );
  NAND U28140 ( .A(n23441), .B(n23442), .Z(n23426) );
  NAND U28141 ( .A(n23443), .B(n23444), .Z(n23442) );
  OR U28142 ( .A(n23445), .B(n23446), .Z(n23443) );
  NANDN U28143 ( .A(n23447), .B(n23445), .Z(n23441) );
  IV U28144 ( .A(n23446), .Z(n23447) );
  NAND U28145 ( .A(n23448), .B(n23449), .Z(n23423) );
  NAND U28146 ( .A(n23450), .B(n23451), .Z(n23449) );
  NANDN U28147 ( .A(n23452), .B(n23453), .Z(n23450) );
  NANDN U28148 ( .A(n23453), .B(n23452), .Z(n23448) );
  AND U28149 ( .A(n23454), .B(n23455), .Z(n23425) );
  NAND U28150 ( .A(n23456), .B(n23457), .Z(n23455) );
  OR U28151 ( .A(n23458), .B(n23459), .Z(n23456) );
  NANDN U28152 ( .A(n23460), .B(n23458), .Z(n23454) );
  NAND U28153 ( .A(n23461), .B(n23462), .Z(n23429) );
  NANDN U28154 ( .A(n23463), .B(n23464), .Z(n23462) );
  OR U28155 ( .A(n23465), .B(n23466), .Z(n23464) );
  NANDN U28156 ( .A(n23467), .B(n23465), .Z(n23461) );
  IV U28157 ( .A(n23466), .Z(n23467) );
  XNOR U28158 ( .A(n23437), .B(n23468), .Z(n23432) );
  XNOR U28159 ( .A(n23435), .B(n23438), .Z(n23468) );
  NAND U28160 ( .A(n23469), .B(n23470), .Z(n23438) );
  NAND U28161 ( .A(n23471), .B(n23472), .Z(n23470) );
  OR U28162 ( .A(n23473), .B(n23474), .Z(n23471) );
  NANDN U28163 ( .A(n23475), .B(n23473), .Z(n23469) );
  IV U28164 ( .A(n23474), .Z(n23475) );
  NAND U28165 ( .A(n23476), .B(n23477), .Z(n23435) );
  NAND U28166 ( .A(n23478), .B(n23479), .Z(n23477) );
  NANDN U28167 ( .A(n23480), .B(n23481), .Z(n23478) );
  NANDN U28168 ( .A(n23481), .B(n23480), .Z(n23476) );
  AND U28169 ( .A(n23482), .B(n23483), .Z(n23437) );
  NAND U28170 ( .A(n23484), .B(n23485), .Z(n23483) );
  OR U28171 ( .A(n23486), .B(n23487), .Z(n23484) );
  NANDN U28172 ( .A(n23488), .B(n23486), .Z(n23482) );
  XNOR U28173 ( .A(n23463), .B(n23489), .Z(N28230) );
  XOR U28174 ( .A(n23465), .B(n23466), .Z(n23489) );
  XNOR U28175 ( .A(n23479), .B(n23490), .Z(n23466) );
  XOR U28176 ( .A(n23480), .B(n23481), .Z(n23490) );
  XOR U28177 ( .A(n23486), .B(n23491), .Z(n23481) );
  XOR U28178 ( .A(n23485), .B(n23488), .Z(n23491) );
  IV U28179 ( .A(n23487), .Z(n23488) );
  NAND U28180 ( .A(n23492), .B(n23493), .Z(n23487) );
  OR U28181 ( .A(n23494), .B(n23495), .Z(n23493) );
  OR U28182 ( .A(n23496), .B(n23497), .Z(n23492) );
  NAND U28183 ( .A(n23498), .B(n23499), .Z(n23485) );
  OR U28184 ( .A(n23500), .B(n23501), .Z(n23499) );
  OR U28185 ( .A(n23502), .B(n23503), .Z(n23498) );
  NOR U28186 ( .A(n23504), .B(n23505), .Z(n23486) );
  ANDN U28187 ( .B(n23506), .A(n23507), .Z(n23480) );
  XNOR U28188 ( .A(n23473), .B(n23508), .Z(n23479) );
  XNOR U28189 ( .A(n23472), .B(n23474), .Z(n23508) );
  NAND U28190 ( .A(n23509), .B(n23510), .Z(n23474) );
  OR U28191 ( .A(n23511), .B(n23512), .Z(n23510) );
  OR U28192 ( .A(n23513), .B(n23514), .Z(n23509) );
  NAND U28193 ( .A(n23515), .B(n23516), .Z(n23472) );
  OR U28194 ( .A(n23517), .B(n23518), .Z(n23516) );
  OR U28195 ( .A(n23519), .B(n23520), .Z(n23515) );
  ANDN U28196 ( .B(n23521), .A(n23522), .Z(n23473) );
  IV U28197 ( .A(n23523), .Z(n23521) );
  ANDN U28198 ( .B(n23524), .A(n23525), .Z(n23465) );
  XOR U28199 ( .A(n23451), .B(n23526), .Z(n23463) );
  XOR U28200 ( .A(n23452), .B(n23453), .Z(n23526) );
  XOR U28201 ( .A(n23458), .B(n23527), .Z(n23453) );
  XOR U28202 ( .A(n23457), .B(n23460), .Z(n23527) );
  IV U28203 ( .A(n23459), .Z(n23460) );
  NAND U28204 ( .A(n23528), .B(n23529), .Z(n23459) );
  OR U28205 ( .A(n23530), .B(n23531), .Z(n23529) );
  OR U28206 ( .A(n23532), .B(n23533), .Z(n23528) );
  NAND U28207 ( .A(n23534), .B(n23535), .Z(n23457) );
  OR U28208 ( .A(n23536), .B(n23537), .Z(n23535) );
  OR U28209 ( .A(n23538), .B(n23539), .Z(n23534) );
  NOR U28210 ( .A(n23540), .B(n23541), .Z(n23458) );
  ANDN U28211 ( .B(n23542), .A(n23543), .Z(n23452) );
  IV U28212 ( .A(n23544), .Z(n23542) );
  XNOR U28213 ( .A(n23445), .B(n23545), .Z(n23451) );
  XNOR U28214 ( .A(n23444), .B(n23446), .Z(n23545) );
  NAND U28215 ( .A(n23546), .B(n23547), .Z(n23446) );
  OR U28216 ( .A(n23548), .B(n23549), .Z(n23547) );
  OR U28217 ( .A(n23550), .B(n23551), .Z(n23546) );
  NAND U28218 ( .A(n23552), .B(n23553), .Z(n23444) );
  OR U28219 ( .A(n23554), .B(n23555), .Z(n23553) );
  OR U28220 ( .A(n23556), .B(n23557), .Z(n23552) );
  ANDN U28221 ( .B(n23558), .A(n23559), .Z(n23445) );
  IV U28222 ( .A(n23560), .Z(n23558) );
  XNOR U28223 ( .A(n23525), .B(n23524), .Z(N28229) );
  XOR U28224 ( .A(n23544), .B(n23543), .Z(n23524) );
  XNOR U28225 ( .A(n23559), .B(n23560), .Z(n23543) );
  XNOR U28226 ( .A(n23554), .B(n23555), .Z(n23560) );
  XNOR U28227 ( .A(n23556), .B(n23557), .Z(n23555) );
  XNOR U28228 ( .A(y[604]), .B(x[604]), .Z(n23557) );
  XNOR U28229 ( .A(y[605]), .B(x[605]), .Z(n23556) );
  XNOR U28230 ( .A(y[603]), .B(x[603]), .Z(n23554) );
  XNOR U28231 ( .A(n23548), .B(n23549), .Z(n23559) );
  XNOR U28232 ( .A(y[600]), .B(x[600]), .Z(n23549) );
  XNOR U28233 ( .A(n23550), .B(n23551), .Z(n23548) );
  XNOR U28234 ( .A(y[601]), .B(x[601]), .Z(n23551) );
  XNOR U28235 ( .A(y[602]), .B(x[602]), .Z(n23550) );
  XNOR U28236 ( .A(n23541), .B(n23540), .Z(n23544) );
  XNOR U28237 ( .A(n23536), .B(n23537), .Z(n23540) );
  XNOR U28238 ( .A(y[597]), .B(x[597]), .Z(n23537) );
  XNOR U28239 ( .A(n23538), .B(n23539), .Z(n23536) );
  XNOR U28240 ( .A(y[598]), .B(x[598]), .Z(n23539) );
  XNOR U28241 ( .A(y[599]), .B(x[599]), .Z(n23538) );
  XNOR U28242 ( .A(n23530), .B(n23531), .Z(n23541) );
  XNOR U28243 ( .A(y[594]), .B(x[594]), .Z(n23531) );
  XNOR U28244 ( .A(n23532), .B(n23533), .Z(n23530) );
  XNOR U28245 ( .A(y[595]), .B(x[595]), .Z(n23533) );
  XNOR U28246 ( .A(y[596]), .B(x[596]), .Z(n23532) );
  XOR U28247 ( .A(n23506), .B(n23507), .Z(n23525) );
  XNOR U28248 ( .A(n23522), .B(n23523), .Z(n23507) );
  XNOR U28249 ( .A(n23517), .B(n23518), .Z(n23523) );
  XNOR U28250 ( .A(n23519), .B(n23520), .Z(n23518) );
  XNOR U28251 ( .A(y[592]), .B(x[592]), .Z(n23520) );
  XNOR U28252 ( .A(y[593]), .B(x[593]), .Z(n23519) );
  XNOR U28253 ( .A(y[591]), .B(x[591]), .Z(n23517) );
  XNOR U28254 ( .A(n23511), .B(n23512), .Z(n23522) );
  XNOR U28255 ( .A(y[588]), .B(x[588]), .Z(n23512) );
  XNOR U28256 ( .A(n23513), .B(n23514), .Z(n23511) );
  XNOR U28257 ( .A(y[589]), .B(x[589]), .Z(n23514) );
  XNOR U28258 ( .A(y[590]), .B(x[590]), .Z(n23513) );
  XOR U28259 ( .A(n23505), .B(n23504), .Z(n23506) );
  XNOR U28260 ( .A(n23500), .B(n23501), .Z(n23504) );
  XNOR U28261 ( .A(y[585]), .B(x[585]), .Z(n23501) );
  XNOR U28262 ( .A(n23502), .B(n23503), .Z(n23500) );
  XNOR U28263 ( .A(y[586]), .B(x[586]), .Z(n23503) );
  XNOR U28264 ( .A(y[587]), .B(x[587]), .Z(n23502) );
  XNOR U28265 ( .A(n23494), .B(n23495), .Z(n23505) );
  XNOR U28266 ( .A(y[582]), .B(x[582]), .Z(n23495) );
  XNOR U28267 ( .A(n23496), .B(n23497), .Z(n23494) );
  XNOR U28268 ( .A(y[583]), .B(x[583]), .Z(n23497) );
  XNOR U28269 ( .A(y[584]), .B(x[584]), .Z(n23496) );
  NAND U28270 ( .A(n23561), .B(n23562), .Z(N28221) );
  NANDN U28271 ( .A(n23563), .B(n23564), .Z(n23562) );
  OR U28272 ( .A(n23565), .B(n23566), .Z(n23564) );
  NAND U28273 ( .A(n23565), .B(n23566), .Z(n23561) );
  XOR U28274 ( .A(n23565), .B(n23567), .Z(N28220) );
  XNOR U28275 ( .A(n23563), .B(n23566), .Z(n23567) );
  AND U28276 ( .A(n23568), .B(n23569), .Z(n23566) );
  NANDN U28277 ( .A(n23570), .B(n23571), .Z(n23569) );
  NANDN U28278 ( .A(n23572), .B(n23573), .Z(n23571) );
  NANDN U28279 ( .A(n23573), .B(n23572), .Z(n23568) );
  NAND U28280 ( .A(n23574), .B(n23575), .Z(n23563) );
  NANDN U28281 ( .A(n23576), .B(n23577), .Z(n23575) );
  OR U28282 ( .A(n23578), .B(n23579), .Z(n23577) );
  NAND U28283 ( .A(n23579), .B(n23578), .Z(n23574) );
  AND U28284 ( .A(n23580), .B(n23581), .Z(n23565) );
  NANDN U28285 ( .A(n23582), .B(n23583), .Z(n23581) );
  NANDN U28286 ( .A(n23584), .B(n23585), .Z(n23583) );
  NANDN U28287 ( .A(n23585), .B(n23584), .Z(n23580) );
  XOR U28288 ( .A(n23579), .B(n23586), .Z(N28219) );
  XOR U28289 ( .A(n23576), .B(n23578), .Z(n23586) );
  XNOR U28290 ( .A(n23572), .B(n23587), .Z(n23578) );
  XNOR U28291 ( .A(n23570), .B(n23573), .Z(n23587) );
  NAND U28292 ( .A(n23588), .B(n23589), .Z(n23573) );
  NAND U28293 ( .A(n23590), .B(n23591), .Z(n23589) );
  OR U28294 ( .A(n23592), .B(n23593), .Z(n23590) );
  NANDN U28295 ( .A(n23594), .B(n23592), .Z(n23588) );
  IV U28296 ( .A(n23593), .Z(n23594) );
  NAND U28297 ( .A(n23595), .B(n23596), .Z(n23570) );
  NAND U28298 ( .A(n23597), .B(n23598), .Z(n23596) );
  NANDN U28299 ( .A(n23599), .B(n23600), .Z(n23597) );
  NANDN U28300 ( .A(n23600), .B(n23599), .Z(n23595) );
  AND U28301 ( .A(n23601), .B(n23602), .Z(n23572) );
  NAND U28302 ( .A(n23603), .B(n23604), .Z(n23602) );
  OR U28303 ( .A(n23605), .B(n23606), .Z(n23603) );
  NANDN U28304 ( .A(n23607), .B(n23605), .Z(n23601) );
  NAND U28305 ( .A(n23608), .B(n23609), .Z(n23576) );
  NANDN U28306 ( .A(n23610), .B(n23611), .Z(n23609) );
  OR U28307 ( .A(n23612), .B(n23613), .Z(n23611) );
  NANDN U28308 ( .A(n23614), .B(n23612), .Z(n23608) );
  IV U28309 ( .A(n23613), .Z(n23614) );
  XNOR U28310 ( .A(n23584), .B(n23615), .Z(n23579) );
  XNOR U28311 ( .A(n23582), .B(n23585), .Z(n23615) );
  NAND U28312 ( .A(n23616), .B(n23617), .Z(n23585) );
  NAND U28313 ( .A(n23618), .B(n23619), .Z(n23617) );
  OR U28314 ( .A(n23620), .B(n23621), .Z(n23618) );
  NANDN U28315 ( .A(n23622), .B(n23620), .Z(n23616) );
  IV U28316 ( .A(n23621), .Z(n23622) );
  NAND U28317 ( .A(n23623), .B(n23624), .Z(n23582) );
  NAND U28318 ( .A(n23625), .B(n23626), .Z(n23624) );
  NANDN U28319 ( .A(n23627), .B(n23628), .Z(n23625) );
  NANDN U28320 ( .A(n23628), .B(n23627), .Z(n23623) );
  AND U28321 ( .A(n23629), .B(n23630), .Z(n23584) );
  NAND U28322 ( .A(n23631), .B(n23632), .Z(n23630) );
  OR U28323 ( .A(n23633), .B(n23634), .Z(n23631) );
  NANDN U28324 ( .A(n23635), .B(n23633), .Z(n23629) );
  XNOR U28325 ( .A(n23610), .B(n23636), .Z(N28218) );
  XOR U28326 ( .A(n23612), .B(n23613), .Z(n23636) );
  XNOR U28327 ( .A(n23626), .B(n23637), .Z(n23613) );
  XOR U28328 ( .A(n23627), .B(n23628), .Z(n23637) );
  XOR U28329 ( .A(n23633), .B(n23638), .Z(n23628) );
  XOR U28330 ( .A(n23632), .B(n23635), .Z(n23638) );
  IV U28331 ( .A(n23634), .Z(n23635) );
  NAND U28332 ( .A(n23639), .B(n23640), .Z(n23634) );
  OR U28333 ( .A(n23641), .B(n23642), .Z(n23640) );
  OR U28334 ( .A(n23643), .B(n23644), .Z(n23639) );
  NAND U28335 ( .A(n23645), .B(n23646), .Z(n23632) );
  OR U28336 ( .A(n23647), .B(n23648), .Z(n23646) );
  OR U28337 ( .A(n23649), .B(n23650), .Z(n23645) );
  NOR U28338 ( .A(n23651), .B(n23652), .Z(n23633) );
  ANDN U28339 ( .B(n23653), .A(n23654), .Z(n23627) );
  XNOR U28340 ( .A(n23620), .B(n23655), .Z(n23626) );
  XNOR U28341 ( .A(n23619), .B(n23621), .Z(n23655) );
  NAND U28342 ( .A(n23656), .B(n23657), .Z(n23621) );
  OR U28343 ( .A(n23658), .B(n23659), .Z(n23657) );
  OR U28344 ( .A(n23660), .B(n23661), .Z(n23656) );
  NAND U28345 ( .A(n23662), .B(n23663), .Z(n23619) );
  OR U28346 ( .A(n23664), .B(n23665), .Z(n23663) );
  OR U28347 ( .A(n23666), .B(n23667), .Z(n23662) );
  ANDN U28348 ( .B(n23668), .A(n23669), .Z(n23620) );
  IV U28349 ( .A(n23670), .Z(n23668) );
  ANDN U28350 ( .B(n23671), .A(n23672), .Z(n23612) );
  XOR U28351 ( .A(n23598), .B(n23673), .Z(n23610) );
  XOR U28352 ( .A(n23599), .B(n23600), .Z(n23673) );
  XOR U28353 ( .A(n23605), .B(n23674), .Z(n23600) );
  XOR U28354 ( .A(n23604), .B(n23607), .Z(n23674) );
  IV U28355 ( .A(n23606), .Z(n23607) );
  NAND U28356 ( .A(n23675), .B(n23676), .Z(n23606) );
  OR U28357 ( .A(n23677), .B(n23678), .Z(n23676) );
  OR U28358 ( .A(n23679), .B(n23680), .Z(n23675) );
  NAND U28359 ( .A(n23681), .B(n23682), .Z(n23604) );
  OR U28360 ( .A(n23683), .B(n23684), .Z(n23682) );
  OR U28361 ( .A(n23685), .B(n23686), .Z(n23681) );
  NOR U28362 ( .A(n23687), .B(n23688), .Z(n23605) );
  ANDN U28363 ( .B(n23689), .A(n23690), .Z(n23599) );
  IV U28364 ( .A(n23691), .Z(n23689) );
  XNOR U28365 ( .A(n23592), .B(n23692), .Z(n23598) );
  XNOR U28366 ( .A(n23591), .B(n23593), .Z(n23692) );
  NAND U28367 ( .A(n23693), .B(n23694), .Z(n23593) );
  OR U28368 ( .A(n23695), .B(n23696), .Z(n23694) );
  OR U28369 ( .A(n23697), .B(n23698), .Z(n23693) );
  NAND U28370 ( .A(n23699), .B(n23700), .Z(n23591) );
  OR U28371 ( .A(n23701), .B(n23702), .Z(n23700) );
  OR U28372 ( .A(n23703), .B(n23704), .Z(n23699) );
  ANDN U28373 ( .B(n23705), .A(n23706), .Z(n23592) );
  IV U28374 ( .A(n23707), .Z(n23705) );
  XNOR U28375 ( .A(n23672), .B(n23671), .Z(N28217) );
  XOR U28376 ( .A(n23691), .B(n23690), .Z(n23671) );
  XNOR U28377 ( .A(n23706), .B(n23707), .Z(n23690) );
  XNOR U28378 ( .A(n23701), .B(n23702), .Z(n23707) );
  XNOR U28379 ( .A(n23703), .B(n23704), .Z(n23702) );
  XNOR U28380 ( .A(y[580]), .B(x[580]), .Z(n23704) );
  XNOR U28381 ( .A(y[581]), .B(x[581]), .Z(n23703) );
  XNOR U28382 ( .A(y[579]), .B(x[579]), .Z(n23701) );
  XNOR U28383 ( .A(n23695), .B(n23696), .Z(n23706) );
  XNOR U28384 ( .A(y[576]), .B(x[576]), .Z(n23696) );
  XNOR U28385 ( .A(n23697), .B(n23698), .Z(n23695) );
  XNOR U28386 ( .A(y[577]), .B(x[577]), .Z(n23698) );
  XNOR U28387 ( .A(y[578]), .B(x[578]), .Z(n23697) );
  XNOR U28388 ( .A(n23688), .B(n23687), .Z(n23691) );
  XNOR U28389 ( .A(n23683), .B(n23684), .Z(n23687) );
  XNOR U28390 ( .A(y[573]), .B(x[573]), .Z(n23684) );
  XNOR U28391 ( .A(n23685), .B(n23686), .Z(n23683) );
  XNOR U28392 ( .A(y[574]), .B(x[574]), .Z(n23686) );
  XNOR U28393 ( .A(y[575]), .B(x[575]), .Z(n23685) );
  XNOR U28394 ( .A(n23677), .B(n23678), .Z(n23688) );
  XNOR U28395 ( .A(y[570]), .B(x[570]), .Z(n23678) );
  XNOR U28396 ( .A(n23679), .B(n23680), .Z(n23677) );
  XNOR U28397 ( .A(y[571]), .B(x[571]), .Z(n23680) );
  XNOR U28398 ( .A(y[572]), .B(x[572]), .Z(n23679) );
  XOR U28399 ( .A(n23653), .B(n23654), .Z(n23672) );
  XNOR U28400 ( .A(n23669), .B(n23670), .Z(n23654) );
  XNOR U28401 ( .A(n23664), .B(n23665), .Z(n23670) );
  XNOR U28402 ( .A(n23666), .B(n23667), .Z(n23665) );
  XNOR U28403 ( .A(y[568]), .B(x[568]), .Z(n23667) );
  XNOR U28404 ( .A(y[569]), .B(x[569]), .Z(n23666) );
  XNOR U28405 ( .A(y[567]), .B(x[567]), .Z(n23664) );
  XNOR U28406 ( .A(n23658), .B(n23659), .Z(n23669) );
  XNOR U28407 ( .A(y[564]), .B(x[564]), .Z(n23659) );
  XNOR U28408 ( .A(n23660), .B(n23661), .Z(n23658) );
  XNOR U28409 ( .A(y[565]), .B(x[565]), .Z(n23661) );
  XNOR U28410 ( .A(y[566]), .B(x[566]), .Z(n23660) );
  XOR U28411 ( .A(n23652), .B(n23651), .Z(n23653) );
  XNOR U28412 ( .A(n23647), .B(n23648), .Z(n23651) );
  XNOR U28413 ( .A(y[561]), .B(x[561]), .Z(n23648) );
  XNOR U28414 ( .A(n23649), .B(n23650), .Z(n23647) );
  XNOR U28415 ( .A(y[562]), .B(x[562]), .Z(n23650) );
  XNOR U28416 ( .A(y[563]), .B(x[563]), .Z(n23649) );
  XNOR U28417 ( .A(n23641), .B(n23642), .Z(n23652) );
  XNOR U28418 ( .A(y[558]), .B(x[558]), .Z(n23642) );
  XNOR U28419 ( .A(n23643), .B(n23644), .Z(n23641) );
  XNOR U28420 ( .A(y[559]), .B(x[559]), .Z(n23644) );
  XNOR U28421 ( .A(y[560]), .B(x[560]), .Z(n23643) );
  NAND U28422 ( .A(n23708), .B(n23709), .Z(N28209) );
  NANDN U28423 ( .A(n23710), .B(n23711), .Z(n23709) );
  OR U28424 ( .A(n23712), .B(n23713), .Z(n23711) );
  NAND U28425 ( .A(n23712), .B(n23713), .Z(n23708) );
  XOR U28426 ( .A(n23712), .B(n23714), .Z(N28208) );
  XNOR U28427 ( .A(n23710), .B(n23713), .Z(n23714) );
  AND U28428 ( .A(n23715), .B(n23716), .Z(n23713) );
  NANDN U28429 ( .A(n23717), .B(n23718), .Z(n23716) );
  NANDN U28430 ( .A(n23719), .B(n23720), .Z(n23718) );
  NANDN U28431 ( .A(n23720), .B(n23719), .Z(n23715) );
  NAND U28432 ( .A(n23721), .B(n23722), .Z(n23710) );
  NANDN U28433 ( .A(n23723), .B(n23724), .Z(n23722) );
  OR U28434 ( .A(n23725), .B(n23726), .Z(n23724) );
  NAND U28435 ( .A(n23726), .B(n23725), .Z(n23721) );
  AND U28436 ( .A(n23727), .B(n23728), .Z(n23712) );
  NANDN U28437 ( .A(n23729), .B(n23730), .Z(n23728) );
  NANDN U28438 ( .A(n23731), .B(n23732), .Z(n23730) );
  NANDN U28439 ( .A(n23732), .B(n23731), .Z(n23727) );
  XOR U28440 ( .A(n23726), .B(n23733), .Z(N28207) );
  XOR U28441 ( .A(n23723), .B(n23725), .Z(n23733) );
  XNOR U28442 ( .A(n23719), .B(n23734), .Z(n23725) );
  XNOR U28443 ( .A(n23717), .B(n23720), .Z(n23734) );
  NAND U28444 ( .A(n23735), .B(n23736), .Z(n23720) );
  NAND U28445 ( .A(n23737), .B(n23738), .Z(n23736) );
  OR U28446 ( .A(n23739), .B(n23740), .Z(n23737) );
  NANDN U28447 ( .A(n23741), .B(n23739), .Z(n23735) );
  IV U28448 ( .A(n23740), .Z(n23741) );
  NAND U28449 ( .A(n23742), .B(n23743), .Z(n23717) );
  NAND U28450 ( .A(n23744), .B(n23745), .Z(n23743) );
  NANDN U28451 ( .A(n23746), .B(n23747), .Z(n23744) );
  NANDN U28452 ( .A(n23747), .B(n23746), .Z(n23742) );
  AND U28453 ( .A(n23748), .B(n23749), .Z(n23719) );
  NAND U28454 ( .A(n23750), .B(n23751), .Z(n23749) );
  OR U28455 ( .A(n23752), .B(n23753), .Z(n23750) );
  NANDN U28456 ( .A(n23754), .B(n23752), .Z(n23748) );
  NAND U28457 ( .A(n23755), .B(n23756), .Z(n23723) );
  NANDN U28458 ( .A(n23757), .B(n23758), .Z(n23756) );
  OR U28459 ( .A(n23759), .B(n23760), .Z(n23758) );
  NANDN U28460 ( .A(n23761), .B(n23759), .Z(n23755) );
  IV U28461 ( .A(n23760), .Z(n23761) );
  XNOR U28462 ( .A(n23731), .B(n23762), .Z(n23726) );
  XNOR U28463 ( .A(n23729), .B(n23732), .Z(n23762) );
  NAND U28464 ( .A(n23763), .B(n23764), .Z(n23732) );
  NAND U28465 ( .A(n23765), .B(n23766), .Z(n23764) );
  OR U28466 ( .A(n23767), .B(n23768), .Z(n23765) );
  NANDN U28467 ( .A(n23769), .B(n23767), .Z(n23763) );
  IV U28468 ( .A(n23768), .Z(n23769) );
  NAND U28469 ( .A(n23770), .B(n23771), .Z(n23729) );
  NAND U28470 ( .A(n23772), .B(n23773), .Z(n23771) );
  NANDN U28471 ( .A(n23774), .B(n23775), .Z(n23772) );
  NANDN U28472 ( .A(n23775), .B(n23774), .Z(n23770) );
  AND U28473 ( .A(n23776), .B(n23777), .Z(n23731) );
  NAND U28474 ( .A(n23778), .B(n23779), .Z(n23777) );
  OR U28475 ( .A(n23780), .B(n23781), .Z(n23778) );
  NANDN U28476 ( .A(n23782), .B(n23780), .Z(n23776) );
  XNOR U28477 ( .A(n23757), .B(n23783), .Z(N28206) );
  XOR U28478 ( .A(n23759), .B(n23760), .Z(n23783) );
  XNOR U28479 ( .A(n23773), .B(n23784), .Z(n23760) );
  XOR U28480 ( .A(n23774), .B(n23775), .Z(n23784) );
  XOR U28481 ( .A(n23780), .B(n23785), .Z(n23775) );
  XOR U28482 ( .A(n23779), .B(n23782), .Z(n23785) );
  IV U28483 ( .A(n23781), .Z(n23782) );
  NAND U28484 ( .A(n23786), .B(n23787), .Z(n23781) );
  OR U28485 ( .A(n23788), .B(n23789), .Z(n23787) );
  OR U28486 ( .A(n23790), .B(n23791), .Z(n23786) );
  NAND U28487 ( .A(n23792), .B(n23793), .Z(n23779) );
  OR U28488 ( .A(n23794), .B(n23795), .Z(n23793) );
  OR U28489 ( .A(n23796), .B(n23797), .Z(n23792) );
  NOR U28490 ( .A(n23798), .B(n23799), .Z(n23780) );
  ANDN U28491 ( .B(n23800), .A(n23801), .Z(n23774) );
  XNOR U28492 ( .A(n23767), .B(n23802), .Z(n23773) );
  XNOR U28493 ( .A(n23766), .B(n23768), .Z(n23802) );
  NAND U28494 ( .A(n23803), .B(n23804), .Z(n23768) );
  OR U28495 ( .A(n23805), .B(n23806), .Z(n23804) );
  OR U28496 ( .A(n23807), .B(n23808), .Z(n23803) );
  NAND U28497 ( .A(n23809), .B(n23810), .Z(n23766) );
  OR U28498 ( .A(n23811), .B(n23812), .Z(n23810) );
  OR U28499 ( .A(n23813), .B(n23814), .Z(n23809) );
  ANDN U28500 ( .B(n23815), .A(n23816), .Z(n23767) );
  IV U28501 ( .A(n23817), .Z(n23815) );
  ANDN U28502 ( .B(n23818), .A(n23819), .Z(n23759) );
  XOR U28503 ( .A(n23745), .B(n23820), .Z(n23757) );
  XOR U28504 ( .A(n23746), .B(n23747), .Z(n23820) );
  XOR U28505 ( .A(n23752), .B(n23821), .Z(n23747) );
  XOR U28506 ( .A(n23751), .B(n23754), .Z(n23821) );
  IV U28507 ( .A(n23753), .Z(n23754) );
  NAND U28508 ( .A(n23822), .B(n23823), .Z(n23753) );
  OR U28509 ( .A(n23824), .B(n23825), .Z(n23823) );
  OR U28510 ( .A(n23826), .B(n23827), .Z(n23822) );
  NAND U28511 ( .A(n23828), .B(n23829), .Z(n23751) );
  OR U28512 ( .A(n23830), .B(n23831), .Z(n23829) );
  OR U28513 ( .A(n23832), .B(n23833), .Z(n23828) );
  NOR U28514 ( .A(n23834), .B(n23835), .Z(n23752) );
  ANDN U28515 ( .B(n23836), .A(n23837), .Z(n23746) );
  IV U28516 ( .A(n23838), .Z(n23836) );
  XNOR U28517 ( .A(n23739), .B(n23839), .Z(n23745) );
  XNOR U28518 ( .A(n23738), .B(n23740), .Z(n23839) );
  NAND U28519 ( .A(n23840), .B(n23841), .Z(n23740) );
  OR U28520 ( .A(n23842), .B(n23843), .Z(n23841) );
  OR U28521 ( .A(n23844), .B(n23845), .Z(n23840) );
  NAND U28522 ( .A(n23846), .B(n23847), .Z(n23738) );
  OR U28523 ( .A(n23848), .B(n23849), .Z(n23847) );
  OR U28524 ( .A(n23850), .B(n23851), .Z(n23846) );
  ANDN U28525 ( .B(n23852), .A(n23853), .Z(n23739) );
  IV U28526 ( .A(n23854), .Z(n23852) );
  XNOR U28527 ( .A(n23819), .B(n23818), .Z(N28205) );
  XOR U28528 ( .A(n23838), .B(n23837), .Z(n23818) );
  XNOR U28529 ( .A(n23853), .B(n23854), .Z(n23837) );
  XNOR U28530 ( .A(n23848), .B(n23849), .Z(n23854) );
  XNOR U28531 ( .A(n23850), .B(n23851), .Z(n23849) );
  XNOR U28532 ( .A(y[556]), .B(x[556]), .Z(n23851) );
  XNOR U28533 ( .A(y[557]), .B(x[557]), .Z(n23850) );
  XNOR U28534 ( .A(y[555]), .B(x[555]), .Z(n23848) );
  XNOR U28535 ( .A(n23842), .B(n23843), .Z(n23853) );
  XNOR U28536 ( .A(y[552]), .B(x[552]), .Z(n23843) );
  XNOR U28537 ( .A(n23844), .B(n23845), .Z(n23842) );
  XNOR U28538 ( .A(y[553]), .B(x[553]), .Z(n23845) );
  XNOR U28539 ( .A(y[554]), .B(x[554]), .Z(n23844) );
  XNOR U28540 ( .A(n23835), .B(n23834), .Z(n23838) );
  XNOR U28541 ( .A(n23830), .B(n23831), .Z(n23834) );
  XNOR U28542 ( .A(y[549]), .B(x[549]), .Z(n23831) );
  XNOR U28543 ( .A(n23832), .B(n23833), .Z(n23830) );
  XNOR U28544 ( .A(y[550]), .B(x[550]), .Z(n23833) );
  XNOR U28545 ( .A(y[551]), .B(x[551]), .Z(n23832) );
  XNOR U28546 ( .A(n23824), .B(n23825), .Z(n23835) );
  XNOR U28547 ( .A(y[546]), .B(x[546]), .Z(n23825) );
  XNOR U28548 ( .A(n23826), .B(n23827), .Z(n23824) );
  XNOR U28549 ( .A(y[547]), .B(x[547]), .Z(n23827) );
  XNOR U28550 ( .A(y[548]), .B(x[548]), .Z(n23826) );
  XOR U28551 ( .A(n23800), .B(n23801), .Z(n23819) );
  XNOR U28552 ( .A(n23816), .B(n23817), .Z(n23801) );
  XNOR U28553 ( .A(n23811), .B(n23812), .Z(n23817) );
  XNOR U28554 ( .A(n23813), .B(n23814), .Z(n23812) );
  XNOR U28555 ( .A(y[544]), .B(x[544]), .Z(n23814) );
  XNOR U28556 ( .A(y[545]), .B(x[545]), .Z(n23813) );
  XNOR U28557 ( .A(y[543]), .B(x[543]), .Z(n23811) );
  XNOR U28558 ( .A(n23805), .B(n23806), .Z(n23816) );
  XNOR U28559 ( .A(y[540]), .B(x[540]), .Z(n23806) );
  XNOR U28560 ( .A(n23807), .B(n23808), .Z(n23805) );
  XNOR U28561 ( .A(y[541]), .B(x[541]), .Z(n23808) );
  XNOR U28562 ( .A(y[542]), .B(x[542]), .Z(n23807) );
  XOR U28563 ( .A(n23799), .B(n23798), .Z(n23800) );
  XNOR U28564 ( .A(n23794), .B(n23795), .Z(n23798) );
  XNOR U28565 ( .A(y[537]), .B(x[537]), .Z(n23795) );
  XNOR U28566 ( .A(n23796), .B(n23797), .Z(n23794) );
  XNOR U28567 ( .A(y[538]), .B(x[538]), .Z(n23797) );
  XNOR U28568 ( .A(y[539]), .B(x[539]), .Z(n23796) );
  XNOR U28569 ( .A(n23788), .B(n23789), .Z(n23799) );
  XNOR U28570 ( .A(y[534]), .B(x[534]), .Z(n23789) );
  XNOR U28571 ( .A(n23790), .B(n23791), .Z(n23788) );
  XNOR U28572 ( .A(y[535]), .B(x[535]), .Z(n23791) );
  XNOR U28573 ( .A(y[536]), .B(x[536]), .Z(n23790) );
  NAND U28574 ( .A(n23855), .B(n23856), .Z(N28197) );
  NANDN U28575 ( .A(n23857), .B(n23858), .Z(n23856) );
  OR U28576 ( .A(n23859), .B(n23860), .Z(n23858) );
  NAND U28577 ( .A(n23859), .B(n23860), .Z(n23855) );
  XOR U28578 ( .A(n23859), .B(n23861), .Z(N28196) );
  XNOR U28579 ( .A(n23857), .B(n23860), .Z(n23861) );
  AND U28580 ( .A(n23862), .B(n23863), .Z(n23860) );
  NANDN U28581 ( .A(n23864), .B(n23865), .Z(n23863) );
  NANDN U28582 ( .A(n23866), .B(n23867), .Z(n23865) );
  NANDN U28583 ( .A(n23867), .B(n23866), .Z(n23862) );
  NAND U28584 ( .A(n23868), .B(n23869), .Z(n23857) );
  NANDN U28585 ( .A(n23870), .B(n23871), .Z(n23869) );
  OR U28586 ( .A(n23872), .B(n23873), .Z(n23871) );
  NAND U28587 ( .A(n23873), .B(n23872), .Z(n23868) );
  AND U28588 ( .A(n23874), .B(n23875), .Z(n23859) );
  NANDN U28589 ( .A(n23876), .B(n23877), .Z(n23875) );
  NANDN U28590 ( .A(n23878), .B(n23879), .Z(n23877) );
  NANDN U28591 ( .A(n23879), .B(n23878), .Z(n23874) );
  XOR U28592 ( .A(n23873), .B(n23880), .Z(N28195) );
  XOR U28593 ( .A(n23870), .B(n23872), .Z(n23880) );
  XNOR U28594 ( .A(n23866), .B(n23881), .Z(n23872) );
  XNOR U28595 ( .A(n23864), .B(n23867), .Z(n23881) );
  NAND U28596 ( .A(n23882), .B(n23883), .Z(n23867) );
  NAND U28597 ( .A(n23884), .B(n23885), .Z(n23883) );
  OR U28598 ( .A(n23886), .B(n23887), .Z(n23884) );
  NANDN U28599 ( .A(n23888), .B(n23886), .Z(n23882) );
  IV U28600 ( .A(n23887), .Z(n23888) );
  NAND U28601 ( .A(n23889), .B(n23890), .Z(n23864) );
  NAND U28602 ( .A(n23891), .B(n23892), .Z(n23890) );
  NANDN U28603 ( .A(n23893), .B(n23894), .Z(n23891) );
  NANDN U28604 ( .A(n23894), .B(n23893), .Z(n23889) );
  AND U28605 ( .A(n23895), .B(n23896), .Z(n23866) );
  NAND U28606 ( .A(n23897), .B(n23898), .Z(n23896) );
  OR U28607 ( .A(n23899), .B(n23900), .Z(n23897) );
  NANDN U28608 ( .A(n23901), .B(n23899), .Z(n23895) );
  NAND U28609 ( .A(n23902), .B(n23903), .Z(n23870) );
  NANDN U28610 ( .A(n23904), .B(n23905), .Z(n23903) );
  OR U28611 ( .A(n23906), .B(n23907), .Z(n23905) );
  NANDN U28612 ( .A(n23908), .B(n23906), .Z(n23902) );
  IV U28613 ( .A(n23907), .Z(n23908) );
  XNOR U28614 ( .A(n23878), .B(n23909), .Z(n23873) );
  XNOR U28615 ( .A(n23876), .B(n23879), .Z(n23909) );
  NAND U28616 ( .A(n23910), .B(n23911), .Z(n23879) );
  NAND U28617 ( .A(n23912), .B(n23913), .Z(n23911) );
  OR U28618 ( .A(n23914), .B(n23915), .Z(n23912) );
  NANDN U28619 ( .A(n23916), .B(n23914), .Z(n23910) );
  IV U28620 ( .A(n23915), .Z(n23916) );
  NAND U28621 ( .A(n23917), .B(n23918), .Z(n23876) );
  NAND U28622 ( .A(n23919), .B(n23920), .Z(n23918) );
  NANDN U28623 ( .A(n23921), .B(n23922), .Z(n23919) );
  NANDN U28624 ( .A(n23922), .B(n23921), .Z(n23917) );
  AND U28625 ( .A(n23923), .B(n23924), .Z(n23878) );
  NAND U28626 ( .A(n23925), .B(n23926), .Z(n23924) );
  OR U28627 ( .A(n23927), .B(n23928), .Z(n23925) );
  NANDN U28628 ( .A(n23929), .B(n23927), .Z(n23923) );
  XNOR U28629 ( .A(n23904), .B(n23930), .Z(N28194) );
  XOR U28630 ( .A(n23906), .B(n23907), .Z(n23930) );
  XNOR U28631 ( .A(n23920), .B(n23931), .Z(n23907) );
  XOR U28632 ( .A(n23921), .B(n23922), .Z(n23931) );
  XOR U28633 ( .A(n23927), .B(n23932), .Z(n23922) );
  XOR U28634 ( .A(n23926), .B(n23929), .Z(n23932) );
  IV U28635 ( .A(n23928), .Z(n23929) );
  NAND U28636 ( .A(n23933), .B(n23934), .Z(n23928) );
  OR U28637 ( .A(n23935), .B(n23936), .Z(n23934) );
  OR U28638 ( .A(n23937), .B(n23938), .Z(n23933) );
  NAND U28639 ( .A(n23939), .B(n23940), .Z(n23926) );
  OR U28640 ( .A(n23941), .B(n23942), .Z(n23940) );
  OR U28641 ( .A(n23943), .B(n23944), .Z(n23939) );
  NOR U28642 ( .A(n23945), .B(n23946), .Z(n23927) );
  ANDN U28643 ( .B(n23947), .A(n23948), .Z(n23921) );
  XNOR U28644 ( .A(n23914), .B(n23949), .Z(n23920) );
  XNOR U28645 ( .A(n23913), .B(n23915), .Z(n23949) );
  NAND U28646 ( .A(n23950), .B(n23951), .Z(n23915) );
  OR U28647 ( .A(n23952), .B(n23953), .Z(n23951) );
  OR U28648 ( .A(n23954), .B(n23955), .Z(n23950) );
  NAND U28649 ( .A(n23956), .B(n23957), .Z(n23913) );
  OR U28650 ( .A(n23958), .B(n23959), .Z(n23957) );
  OR U28651 ( .A(n23960), .B(n23961), .Z(n23956) );
  ANDN U28652 ( .B(n23962), .A(n23963), .Z(n23914) );
  IV U28653 ( .A(n23964), .Z(n23962) );
  ANDN U28654 ( .B(n23965), .A(n23966), .Z(n23906) );
  XOR U28655 ( .A(n23892), .B(n23967), .Z(n23904) );
  XOR U28656 ( .A(n23893), .B(n23894), .Z(n23967) );
  XOR U28657 ( .A(n23899), .B(n23968), .Z(n23894) );
  XOR U28658 ( .A(n23898), .B(n23901), .Z(n23968) );
  IV U28659 ( .A(n23900), .Z(n23901) );
  NAND U28660 ( .A(n23969), .B(n23970), .Z(n23900) );
  OR U28661 ( .A(n23971), .B(n23972), .Z(n23970) );
  OR U28662 ( .A(n23973), .B(n23974), .Z(n23969) );
  NAND U28663 ( .A(n23975), .B(n23976), .Z(n23898) );
  OR U28664 ( .A(n23977), .B(n23978), .Z(n23976) );
  OR U28665 ( .A(n23979), .B(n23980), .Z(n23975) );
  NOR U28666 ( .A(n23981), .B(n23982), .Z(n23899) );
  ANDN U28667 ( .B(n23983), .A(n23984), .Z(n23893) );
  IV U28668 ( .A(n23985), .Z(n23983) );
  XNOR U28669 ( .A(n23886), .B(n23986), .Z(n23892) );
  XNOR U28670 ( .A(n23885), .B(n23887), .Z(n23986) );
  NAND U28671 ( .A(n23987), .B(n23988), .Z(n23887) );
  OR U28672 ( .A(n23989), .B(n23990), .Z(n23988) );
  OR U28673 ( .A(n23991), .B(n23992), .Z(n23987) );
  NAND U28674 ( .A(n23993), .B(n23994), .Z(n23885) );
  OR U28675 ( .A(n23995), .B(n23996), .Z(n23994) );
  OR U28676 ( .A(n23997), .B(n23998), .Z(n23993) );
  ANDN U28677 ( .B(n23999), .A(n24000), .Z(n23886) );
  IV U28678 ( .A(n24001), .Z(n23999) );
  XNOR U28679 ( .A(n23966), .B(n23965), .Z(N28193) );
  XOR U28680 ( .A(n23985), .B(n23984), .Z(n23965) );
  XNOR U28681 ( .A(n24000), .B(n24001), .Z(n23984) );
  XNOR U28682 ( .A(n23995), .B(n23996), .Z(n24001) );
  XNOR U28683 ( .A(n23997), .B(n23998), .Z(n23996) );
  XNOR U28684 ( .A(y[532]), .B(x[532]), .Z(n23998) );
  XNOR U28685 ( .A(y[533]), .B(x[533]), .Z(n23997) );
  XNOR U28686 ( .A(y[531]), .B(x[531]), .Z(n23995) );
  XNOR U28687 ( .A(n23989), .B(n23990), .Z(n24000) );
  XNOR U28688 ( .A(y[528]), .B(x[528]), .Z(n23990) );
  XNOR U28689 ( .A(n23991), .B(n23992), .Z(n23989) );
  XNOR U28690 ( .A(y[529]), .B(x[529]), .Z(n23992) );
  XNOR U28691 ( .A(y[530]), .B(x[530]), .Z(n23991) );
  XNOR U28692 ( .A(n23982), .B(n23981), .Z(n23985) );
  XNOR U28693 ( .A(n23977), .B(n23978), .Z(n23981) );
  XNOR U28694 ( .A(y[525]), .B(x[525]), .Z(n23978) );
  XNOR U28695 ( .A(n23979), .B(n23980), .Z(n23977) );
  XNOR U28696 ( .A(y[526]), .B(x[526]), .Z(n23980) );
  XNOR U28697 ( .A(y[527]), .B(x[527]), .Z(n23979) );
  XNOR U28698 ( .A(n23971), .B(n23972), .Z(n23982) );
  XNOR U28699 ( .A(y[522]), .B(x[522]), .Z(n23972) );
  XNOR U28700 ( .A(n23973), .B(n23974), .Z(n23971) );
  XNOR U28701 ( .A(y[523]), .B(x[523]), .Z(n23974) );
  XNOR U28702 ( .A(y[524]), .B(x[524]), .Z(n23973) );
  XOR U28703 ( .A(n23947), .B(n23948), .Z(n23966) );
  XNOR U28704 ( .A(n23963), .B(n23964), .Z(n23948) );
  XNOR U28705 ( .A(n23958), .B(n23959), .Z(n23964) );
  XNOR U28706 ( .A(n23960), .B(n23961), .Z(n23959) );
  XNOR U28707 ( .A(y[520]), .B(x[520]), .Z(n23961) );
  XNOR U28708 ( .A(y[521]), .B(x[521]), .Z(n23960) );
  XNOR U28709 ( .A(y[519]), .B(x[519]), .Z(n23958) );
  XNOR U28710 ( .A(n23952), .B(n23953), .Z(n23963) );
  XNOR U28711 ( .A(y[516]), .B(x[516]), .Z(n23953) );
  XNOR U28712 ( .A(n23954), .B(n23955), .Z(n23952) );
  XNOR U28713 ( .A(y[517]), .B(x[517]), .Z(n23955) );
  XNOR U28714 ( .A(y[518]), .B(x[518]), .Z(n23954) );
  XOR U28715 ( .A(n23946), .B(n23945), .Z(n23947) );
  XNOR U28716 ( .A(n23941), .B(n23942), .Z(n23945) );
  XNOR U28717 ( .A(y[513]), .B(x[513]), .Z(n23942) );
  XNOR U28718 ( .A(n23943), .B(n23944), .Z(n23941) );
  XNOR U28719 ( .A(y[514]), .B(x[514]), .Z(n23944) );
  XNOR U28720 ( .A(y[515]), .B(x[515]), .Z(n23943) );
  XNOR U28721 ( .A(n23935), .B(n23936), .Z(n23946) );
  XNOR U28722 ( .A(y[510]), .B(x[510]), .Z(n23936) );
  XNOR U28723 ( .A(n23937), .B(n23938), .Z(n23935) );
  XNOR U28724 ( .A(y[511]), .B(x[511]), .Z(n23938) );
  XNOR U28725 ( .A(y[512]), .B(x[512]), .Z(n23937) );
  NAND U28726 ( .A(n24002), .B(n24003), .Z(N28185) );
  NANDN U28727 ( .A(n24004), .B(n24005), .Z(n24003) );
  OR U28728 ( .A(n24006), .B(n24007), .Z(n24005) );
  NAND U28729 ( .A(n24006), .B(n24007), .Z(n24002) );
  XOR U28730 ( .A(n24006), .B(n24008), .Z(N28184) );
  XNOR U28731 ( .A(n24004), .B(n24007), .Z(n24008) );
  AND U28732 ( .A(n24009), .B(n24010), .Z(n24007) );
  NANDN U28733 ( .A(n24011), .B(n24012), .Z(n24010) );
  NANDN U28734 ( .A(n24013), .B(n24014), .Z(n24012) );
  NANDN U28735 ( .A(n24014), .B(n24013), .Z(n24009) );
  NAND U28736 ( .A(n24015), .B(n24016), .Z(n24004) );
  NANDN U28737 ( .A(n24017), .B(n24018), .Z(n24016) );
  OR U28738 ( .A(n24019), .B(n24020), .Z(n24018) );
  NAND U28739 ( .A(n24020), .B(n24019), .Z(n24015) );
  AND U28740 ( .A(n24021), .B(n24022), .Z(n24006) );
  NANDN U28741 ( .A(n24023), .B(n24024), .Z(n24022) );
  NANDN U28742 ( .A(n24025), .B(n24026), .Z(n24024) );
  NANDN U28743 ( .A(n24026), .B(n24025), .Z(n24021) );
  XOR U28744 ( .A(n24020), .B(n24027), .Z(N28183) );
  XOR U28745 ( .A(n24017), .B(n24019), .Z(n24027) );
  XNOR U28746 ( .A(n24013), .B(n24028), .Z(n24019) );
  XNOR U28747 ( .A(n24011), .B(n24014), .Z(n24028) );
  NAND U28748 ( .A(n24029), .B(n24030), .Z(n24014) );
  NAND U28749 ( .A(n24031), .B(n24032), .Z(n24030) );
  OR U28750 ( .A(n24033), .B(n24034), .Z(n24031) );
  NANDN U28751 ( .A(n24035), .B(n24033), .Z(n24029) );
  IV U28752 ( .A(n24034), .Z(n24035) );
  NAND U28753 ( .A(n24036), .B(n24037), .Z(n24011) );
  NAND U28754 ( .A(n24038), .B(n24039), .Z(n24037) );
  NANDN U28755 ( .A(n24040), .B(n24041), .Z(n24038) );
  NANDN U28756 ( .A(n24041), .B(n24040), .Z(n24036) );
  AND U28757 ( .A(n24042), .B(n24043), .Z(n24013) );
  NAND U28758 ( .A(n24044), .B(n24045), .Z(n24043) );
  OR U28759 ( .A(n24046), .B(n24047), .Z(n24044) );
  NANDN U28760 ( .A(n24048), .B(n24046), .Z(n24042) );
  NAND U28761 ( .A(n24049), .B(n24050), .Z(n24017) );
  NANDN U28762 ( .A(n24051), .B(n24052), .Z(n24050) );
  OR U28763 ( .A(n24053), .B(n24054), .Z(n24052) );
  NANDN U28764 ( .A(n24055), .B(n24053), .Z(n24049) );
  IV U28765 ( .A(n24054), .Z(n24055) );
  XNOR U28766 ( .A(n24025), .B(n24056), .Z(n24020) );
  XNOR U28767 ( .A(n24023), .B(n24026), .Z(n24056) );
  NAND U28768 ( .A(n24057), .B(n24058), .Z(n24026) );
  NAND U28769 ( .A(n24059), .B(n24060), .Z(n24058) );
  OR U28770 ( .A(n24061), .B(n24062), .Z(n24059) );
  NANDN U28771 ( .A(n24063), .B(n24061), .Z(n24057) );
  IV U28772 ( .A(n24062), .Z(n24063) );
  NAND U28773 ( .A(n24064), .B(n24065), .Z(n24023) );
  NAND U28774 ( .A(n24066), .B(n24067), .Z(n24065) );
  NANDN U28775 ( .A(n24068), .B(n24069), .Z(n24066) );
  NANDN U28776 ( .A(n24069), .B(n24068), .Z(n24064) );
  AND U28777 ( .A(n24070), .B(n24071), .Z(n24025) );
  NAND U28778 ( .A(n24072), .B(n24073), .Z(n24071) );
  OR U28779 ( .A(n24074), .B(n24075), .Z(n24072) );
  NANDN U28780 ( .A(n24076), .B(n24074), .Z(n24070) );
  XNOR U28781 ( .A(n24051), .B(n24077), .Z(N28182) );
  XOR U28782 ( .A(n24053), .B(n24054), .Z(n24077) );
  XNOR U28783 ( .A(n24067), .B(n24078), .Z(n24054) );
  XOR U28784 ( .A(n24068), .B(n24069), .Z(n24078) );
  XOR U28785 ( .A(n24074), .B(n24079), .Z(n24069) );
  XOR U28786 ( .A(n24073), .B(n24076), .Z(n24079) );
  IV U28787 ( .A(n24075), .Z(n24076) );
  NAND U28788 ( .A(n24080), .B(n24081), .Z(n24075) );
  OR U28789 ( .A(n24082), .B(n24083), .Z(n24081) );
  OR U28790 ( .A(n24084), .B(n24085), .Z(n24080) );
  NAND U28791 ( .A(n24086), .B(n24087), .Z(n24073) );
  OR U28792 ( .A(n24088), .B(n24089), .Z(n24087) );
  OR U28793 ( .A(n24090), .B(n24091), .Z(n24086) );
  NOR U28794 ( .A(n24092), .B(n24093), .Z(n24074) );
  ANDN U28795 ( .B(n24094), .A(n24095), .Z(n24068) );
  XNOR U28796 ( .A(n24061), .B(n24096), .Z(n24067) );
  XNOR U28797 ( .A(n24060), .B(n24062), .Z(n24096) );
  NAND U28798 ( .A(n24097), .B(n24098), .Z(n24062) );
  OR U28799 ( .A(n24099), .B(n24100), .Z(n24098) );
  OR U28800 ( .A(n24101), .B(n24102), .Z(n24097) );
  NAND U28801 ( .A(n24103), .B(n24104), .Z(n24060) );
  OR U28802 ( .A(n24105), .B(n24106), .Z(n24104) );
  OR U28803 ( .A(n24107), .B(n24108), .Z(n24103) );
  ANDN U28804 ( .B(n24109), .A(n24110), .Z(n24061) );
  IV U28805 ( .A(n24111), .Z(n24109) );
  ANDN U28806 ( .B(n24112), .A(n24113), .Z(n24053) );
  XOR U28807 ( .A(n24039), .B(n24114), .Z(n24051) );
  XOR U28808 ( .A(n24040), .B(n24041), .Z(n24114) );
  XOR U28809 ( .A(n24046), .B(n24115), .Z(n24041) );
  XOR U28810 ( .A(n24045), .B(n24048), .Z(n24115) );
  IV U28811 ( .A(n24047), .Z(n24048) );
  NAND U28812 ( .A(n24116), .B(n24117), .Z(n24047) );
  OR U28813 ( .A(n24118), .B(n24119), .Z(n24117) );
  OR U28814 ( .A(n24120), .B(n24121), .Z(n24116) );
  NAND U28815 ( .A(n24122), .B(n24123), .Z(n24045) );
  OR U28816 ( .A(n24124), .B(n24125), .Z(n24123) );
  OR U28817 ( .A(n24126), .B(n24127), .Z(n24122) );
  NOR U28818 ( .A(n24128), .B(n24129), .Z(n24046) );
  ANDN U28819 ( .B(n24130), .A(n24131), .Z(n24040) );
  IV U28820 ( .A(n24132), .Z(n24130) );
  XNOR U28821 ( .A(n24033), .B(n24133), .Z(n24039) );
  XNOR U28822 ( .A(n24032), .B(n24034), .Z(n24133) );
  NAND U28823 ( .A(n24134), .B(n24135), .Z(n24034) );
  OR U28824 ( .A(n24136), .B(n24137), .Z(n24135) );
  OR U28825 ( .A(n24138), .B(n24139), .Z(n24134) );
  NAND U28826 ( .A(n24140), .B(n24141), .Z(n24032) );
  OR U28827 ( .A(n24142), .B(n24143), .Z(n24141) );
  OR U28828 ( .A(n24144), .B(n24145), .Z(n24140) );
  ANDN U28829 ( .B(n24146), .A(n24147), .Z(n24033) );
  IV U28830 ( .A(n24148), .Z(n24146) );
  XNOR U28831 ( .A(n24113), .B(n24112), .Z(N28181) );
  XOR U28832 ( .A(n24132), .B(n24131), .Z(n24112) );
  XNOR U28833 ( .A(n24147), .B(n24148), .Z(n24131) );
  XNOR U28834 ( .A(n24142), .B(n24143), .Z(n24148) );
  XNOR U28835 ( .A(n24144), .B(n24145), .Z(n24143) );
  XNOR U28836 ( .A(y[508]), .B(x[508]), .Z(n24145) );
  XNOR U28837 ( .A(y[509]), .B(x[509]), .Z(n24144) );
  XNOR U28838 ( .A(y[507]), .B(x[507]), .Z(n24142) );
  XNOR U28839 ( .A(n24136), .B(n24137), .Z(n24147) );
  XNOR U28840 ( .A(y[504]), .B(x[504]), .Z(n24137) );
  XNOR U28841 ( .A(n24138), .B(n24139), .Z(n24136) );
  XNOR U28842 ( .A(y[505]), .B(x[505]), .Z(n24139) );
  XNOR U28843 ( .A(y[506]), .B(x[506]), .Z(n24138) );
  XNOR U28844 ( .A(n24129), .B(n24128), .Z(n24132) );
  XNOR U28845 ( .A(n24124), .B(n24125), .Z(n24128) );
  XNOR U28846 ( .A(y[501]), .B(x[501]), .Z(n24125) );
  XNOR U28847 ( .A(n24126), .B(n24127), .Z(n24124) );
  XNOR U28848 ( .A(y[502]), .B(x[502]), .Z(n24127) );
  XNOR U28849 ( .A(y[503]), .B(x[503]), .Z(n24126) );
  XNOR U28850 ( .A(n24118), .B(n24119), .Z(n24129) );
  XNOR U28851 ( .A(y[498]), .B(x[498]), .Z(n24119) );
  XNOR U28852 ( .A(n24120), .B(n24121), .Z(n24118) );
  XNOR U28853 ( .A(y[499]), .B(x[499]), .Z(n24121) );
  XNOR U28854 ( .A(y[500]), .B(x[500]), .Z(n24120) );
  XOR U28855 ( .A(n24094), .B(n24095), .Z(n24113) );
  XNOR U28856 ( .A(n24110), .B(n24111), .Z(n24095) );
  XNOR U28857 ( .A(n24105), .B(n24106), .Z(n24111) );
  XNOR U28858 ( .A(n24107), .B(n24108), .Z(n24106) );
  XNOR U28859 ( .A(y[496]), .B(x[496]), .Z(n24108) );
  XNOR U28860 ( .A(y[497]), .B(x[497]), .Z(n24107) );
  XNOR U28861 ( .A(y[495]), .B(x[495]), .Z(n24105) );
  XNOR U28862 ( .A(n24099), .B(n24100), .Z(n24110) );
  XNOR U28863 ( .A(y[492]), .B(x[492]), .Z(n24100) );
  XNOR U28864 ( .A(n24101), .B(n24102), .Z(n24099) );
  XNOR U28865 ( .A(y[493]), .B(x[493]), .Z(n24102) );
  XNOR U28866 ( .A(y[494]), .B(x[494]), .Z(n24101) );
  XOR U28867 ( .A(n24093), .B(n24092), .Z(n24094) );
  XNOR U28868 ( .A(n24088), .B(n24089), .Z(n24092) );
  XNOR U28869 ( .A(y[489]), .B(x[489]), .Z(n24089) );
  XNOR U28870 ( .A(n24090), .B(n24091), .Z(n24088) );
  XNOR U28871 ( .A(y[490]), .B(x[490]), .Z(n24091) );
  XNOR U28872 ( .A(y[491]), .B(x[491]), .Z(n24090) );
  XNOR U28873 ( .A(n24082), .B(n24083), .Z(n24093) );
  XNOR U28874 ( .A(y[486]), .B(x[486]), .Z(n24083) );
  XNOR U28875 ( .A(n24084), .B(n24085), .Z(n24082) );
  XNOR U28876 ( .A(y[487]), .B(x[487]), .Z(n24085) );
  XNOR U28877 ( .A(y[488]), .B(x[488]), .Z(n24084) );
  NAND U28878 ( .A(n24149), .B(n24150), .Z(N28173) );
  NANDN U28879 ( .A(n24151), .B(n24152), .Z(n24150) );
  OR U28880 ( .A(n24153), .B(n24154), .Z(n24152) );
  NAND U28881 ( .A(n24153), .B(n24154), .Z(n24149) );
  XOR U28882 ( .A(n24153), .B(n24155), .Z(N28172) );
  XNOR U28883 ( .A(n24151), .B(n24154), .Z(n24155) );
  AND U28884 ( .A(n24156), .B(n24157), .Z(n24154) );
  NANDN U28885 ( .A(n24158), .B(n24159), .Z(n24157) );
  NANDN U28886 ( .A(n24160), .B(n24161), .Z(n24159) );
  NANDN U28887 ( .A(n24161), .B(n24160), .Z(n24156) );
  NAND U28888 ( .A(n24162), .B(n24163), .Z(n24151) );
  NANDN U28889 ( .A(n24164), .B(n24165), .Z(n24163) );
  OR U28890 ( .A(n24166), .B(n24167), .Z(n24165) );
  NAND U28891 ( .A(n24167), .B(n24166), .Z(n24162) );
  AND U28892 ( .A(n24168), .B(n24169), .Z(n24153) );
  NANDN U28893 ( .A(n24170), .B(n24171), .Z(n24169) );
  NANDN U28894 ( .A(n24172), .B(n24173), .Z(n24171) );
  NANDN U28895 ( .A(n24173), .B(n24172), .Z(n24168) );
  XOR U28896 ( .A(n24167), .B(n24174), .Z(N28171) );
  XOR U28897 ( .A(n24164), .B(n24166), .Z(n24174) );
  XNOR U28898 ( .A(n24160), .B(n24175), .Z(n24166) );
  XNOR U28899 ( .A(n24158), .B(n24161), .Z(n24175) );
  NAND U28900 ( .A(n24176), .B(n24177), .Z(n24161) );
  NAND U28901 ( .A(n24178), .B(n24179), .Z(n24177) );
  OR U28902 ( .A(n24180), .B(n24181), .Z(n24178) );
  NANDN U28903 ( .A(n24182), .B(n24180), .Z(n24176) );
  IV U28904 ( .A(n24181), .Z(n24182) );
  NAND U28905 ( .A(n24183), .B(n24184), .Z(n24158) );
  NAND U28906 ( .A(n24185), .B(n24186), .Z(n24184) );
  NANDN U28907 ( .A(n24187), .B(n24188), .Z(n24185) );
  NANDN U28908 ( .A(n24188), .B(n24187), .Z(n24183) );
  AND U28909 ( .A(n24189), .B(n24190), .Z(n24160) );
  NAND U28910 ( .A(n24191), .B(n24192), .Z(n24190) );
  OR U28911 ( .A(n24193), .B(n24194), .Z(n24191) );
  NANDN U28912 ( .A(n24195), .B(n24193), .Z(n24189) );
  NAND U28913 ( .A(n24196), .B(n24197), .Z(n24164) );
  NANDN U28914 ( .A(n24198), .B(n24199), .Z(n24197) );
  OR U28915 ( .A(n24200), .B(n24201), .Z(n24199) );
  NANDN U28916 ( .A(n24202), .B(n24200), .Z(n24196) );
  IV U28917 ( .A(n24201), .Z(n24202) );
  XNOR U28918 ( .A(n24172), .B(n24203), .Z(n24167) );
  XNOR U28919 ( .A(n24170), .B(n24173), .Z(n24203) );
  NAND U28920 ( .A(n24204), .B(n24205), .Z(n24173) );
  NAND U28921 ( .A(n24206), .B(n24207), .Z(n24205) );
  OR U28922 ( .A(n24208), .B(n24209), .Z(n24206) );
  NANDN U28923 ( .A(n24210), .B(n24208), .Z(n24204) );
  IV U28924 ( .A(n24209), .Z(n24210) );
  NAND U28925 ( .A(n24211), .B(n24212), .Z(n24170) );
  NAND U28926 ( .A(n24213), .B(n24214), .Z(n24212) );
  NANDN U28927 ( .A(n24215), .B(n24216), .Z(n24213) );
  NANDN U28928 ( .A(n24216), .B(n24215), .Z(n24211) );
  AND U28929 ( .A(n24217), .B(n24218), .Z(n24172) );
  NAND U28930 ( .A(n24219), .B(n24220), .Z(n24218) );
  OR U28931 ( .A(n24221), .B(n24222), .Z(n24219) );
  NANDN U28932 ( .A(n24223), .B(n24221), .Z(n24217) );
  XNOR U28933 ( .A(n24198), .B(n24224), .Z(N28170) );
  XOR U28934 ( .A(n24200), .B(n24201), .Z(n24224) );
  XNOR U28935 ( .A(n24214), .B(n24225), .Z(n24201) );
  XOR U28936 ( .A(n24215), .B(n24216), .Z(n24225) );
  XOR U28937 ( .A(n24221), .B(n24226), .Z(n24216) );
  XOR U28938 ( .A(n24220), .B(n24223), .Z(n24226) );
  IV U28939 ( .A(n24222), .Z(n24223) );
  NAND U28940 ( .A(n24227), .B(n24228), .Z(n24222) );
  OR U28941 ( .A(n24229), .B(n24230), .Z(n24228) );
  OR U28942 ( .A(n24231), .B(n24232), .Z(n24227) );
  NAND U28943 ( .A(n24233), .B(n24234), .Z(n24220) );
  OR U28944 ( .A(n24235), .B(n24236), .Z(n24234) );
  OR U28945 ( .A(n24237), .B(n24238), .Z(n24233) );
  NOR U28946 ( .A(n24239), .B(n24240), .Z(n24221) );
  ANDN U28947 ( .B(n24241), .A(n24242), .Z(n24215) );
  XNOR U28948 ( .A(n24208), .B(n24243), .Z(n24214) );
  XNOR U28949 ( .A(n24207), .B(n24209), .Z(n24243) );
  NAND U28950 ( .A(n24244), .B(n24245), .Z(n24209) );
  OR U28951 ( .A(n24246), .B(n24247), .Z(n24245) );
  OR U28952 ( .A(n24248), .B(n24249), .Z(n24244) );
  NAND U28953 ( .A(n24250), .B(n24251), .Z(n24207) );
  OR U28954 ( .A(n24252), .B(n24253), .Z(n24251) );
  OR U28955 ( .A(n24254), .B(n24255), .Z(n24250) );
  ANDN U28956 ( .B(n24256), .A(n24257), .Z(n24208) );
  IV U28957 ( .A(n24258), .Z(n24256) );
  ANDN U28958 ( .B(n24259), .A(n24260), .Z(n24200) );
  XOR U28959 ( .A(n24186), .B(n24261), .Z(n24198) );
  XOR U28960 ( .A(n24187), .B(n24188), .Z(n24261) );
  XOR U28961 ( .A(n24193), .B(n24262), .Z(n24188) );
  XOR U28962 ( .A(n24192), .B(n24195), .Z(n24262) );
  IV U28963 ( .A(n24194), .Z(n24195) );
  NAND U28964 ( .A(n24263), .B(n24264), .Z(n24194) );
  OR U28965 ( .A(n24265), .B(n24266), .Z(n24264) );
  OR U28966 ( .A(n24267), .B(n24268), .Z(n24263) );
  NAND U28967 ( .A(n24269), .B(n24270), .Z(n24192) );
  OR U28968 ( .A(n24271), .B(n24272), .Z(n24270) );
  OR U28969 ( .A(n24273), .B(n24274), .Z(n24269) );
  NOR U28970 ( .A(n24275), .B(n24276), .Z(n24193) );
  ANDN U28971 ( .B(n24277), .A(n24278), .Z(n24187) );
  IV U28972 ( .A(n24279), .Z(n24277) );
  XNOR U28973 ( .A(n24180), .B(n24280), .Z(n24186) );
  XNOR U28974 ( .A(n24179), .B(n24181), .Z(n24280) );
  NAND U28975 ( .A(n24281), .B(n24282), .Z(n24181) );
  OR U28976 ( .A(n24283), .B(n24284), .Z(n24282) );
  OR U28977 ( .A(n24285), .B(n24286), .Z(n24281) );
  NAND U28978 ( .A(n24287), .B(n24288), .Z(n24179) );
  OR U28979 ( .A(n24289), .B(n24290), .Z(n24288) );
  OR U28980 ( .A(n24291), .B(n24292), .Z(n24287) );
  ANDN U28981 ( .B(n24293), .A(n24294), .Z(n24180) );
  IV U28982 ( .A(n24295), .Z(n24293) );
  XNOR U28983 ( .A(n24260), .B(n24259), .Z(N28169) );
  XOR U28984 ( .A(n24279), .B(n24278), .Z(n24259) );
  XNOR U28985 ( .A(n24294), .B(n24295), .Z(n24278) );
  XNOR U28986 ( .A(n24289), .B(n24290), .Z(n24295) );
  XNOR U28987 ( .A(n24291), .B(n24292), .Z(n24290) );
  XNOR U28988 ( .A(y[484]), .B(x[484]), .Z(n24292) );
  XNOR U28989 ( .A(y[485]), .B(x[485]), .Z(n24291) );
  XNOR U28990 ( .A(y[483]), .B(x[483]), .Z(n24289) );
  XNOR U28991 ( .A(n24283), .B(n24284), .Z(n24294) );
  XNOR U28992 ( .A(y[480]), .B(x[480]), .Z(n24284) );
  XNOR U28993 ( .A(n24285), .B(n24286), .Z(n24283) );
  XNOR U28994 ( .A(y[481]), .B(x[481]), .Z(n24286) );
  XNOR U28995 ( .A(y[482]), .B(x[482]), .Z(n24285) );
  XNOR U28996 ( .A(n24276), .B(n24275), .Z(n24279) );
  XNOR U28997 ( .A(n24271), .B(n24272), .Z(n24275) );
  XNOR U28998 ( .A(y[477]), .B(x[477]), .Z(n24272) );
  XNOR U28999 ( .A(n24273), .B(n24274), .Z(n24271) );
  XNOR U29000 ( .A(y[478]), .B(x[478]), .Z(n24274) );
  XNOR U29001 ( .A(y[479]), .B(x[479]), .Z(n24273) );
  XNOR U29002 ( .A(n24265), .B(n24266), .Z(n24276) );
  XNOR U29003 ( .A(y[474]), .B(x[474]), .Z(n24266) );
  XNOR U29004 ( .A(n24267), .B(n24268), .Z(n24265) );
  XNOR U29005 ( .A(y[475]), .B(x[475]), .Z(n24268) );
  XNOR U29006 ( .A(y[476]), .B(x[476]), .Z(n24267) );
  XOR U29007 ( .A(n24241), .B(n24242), .Z(n24260) );
  XNOR U29008 ( .A(n24257), .B(n24258), .Z(n24242) );
  XNOR U29009 ( .A(n24252), .B(n24253), .Z(n24258) );
  XNOR U29010 ( .A(n24254), .B(n24255), .Z(n24253) );
  XNOR U29011 ( .A(y[472]), .B(x[472]), .Z(n24255) );
  XNOR U29012 ( .A(y[473]), .B(x[473]), .Z(n24254) );
  XNOR U29013 ( .A(y[471]), .B(x[471]), .Z(n24252) );
  XNOR U29014 ( .A(n24246), .B(n24247), .Z(n24257) );
  XNOR U29015 ( .A(y[468]), .B(x[468]), .Z(n24247) );
  XNOR U29016 ( .A(n24248), .B(n24249), .Z(n24246) );
  XNOR U29017 ( .A(y[469]), .B(x[469]), .Z(n24249) );
  XNOR U29018 ( .A(y[470]), .B(x[470]), .Z(n24248) );
  XOR U29019 ( .A(n24240), .B(n24239), .Z(n24241) );
  XNOR U29020 ( .A(n24235), .B(n24236), .Z(n24239) );
  XNOR U29021 ( .A(y[465]), .B(x[465]), .Z(n24236) );
  XNOR U29022 ( .A(n24237), .B(n24238), .Z(n24235) );
  XNOR U29023 ( .A(y[466]), .B(x[466]), .Z(n24238) );
  XNOR U29024 ( .A(y[467]), .B(x[467]), .Z(n24237) );
  XNOR U29025 ( .A(n24229), .B(n24230), .Z(n24240) );
  XNOR U29026 ( .A(y[462]), .B(x[462]), .Z(n24230) );
  XNOR U29027 ( .A(n24231), .B(n24232), .Z(n24229) );
  XNOR U29028 ( .A(y[463]), .B(x[463]), .Z(n24232) );
  XNOR U29029 ( .A(y[464]), .B(x[464]), .Z(n24231) );
  NAND U29030 ( .A(n24296), .B(n24297), .Z(N28161) );
  NANDN U29031 ( .A(n24298), .B(n24299), .Z(n24297) );
  OR U29032 ( .A(n24300), .B(n24301), .Z(n24299) );
  NAND U29033 ( .A(n24300), .B(n24301), .Z(n24296) );
  XOR U29034 ( .A(n24300), .B(n24302), .Z(N28160) );
  XNOR U29035 ( .A(n24298), .B(n24301), .Z(n24302) );
  AND U29036 ( .A(n24303), .B(n24304), .Z(n24301) );
  NANDN U29037 ( .A(n24305), .B(n24306), .Z(n24304) );
  NANDN U29038 ( .A(n24307), .B(n24308), .Z(n24306) );
  NANDN U29039 ( .A(n24308), .B(n24307), .Z(n24303) );
  NAND U29040 ( .A(n24309), .B(n24310), .Z(n24298) );
  NANDN U29041 ( .A(n24311), .B(n24312), .Z(n24310) );
  OR U29042 ( .A(n24313), .B(n24314), .Z(n24312) );
  NAND U29043 ( .A(n24314), .B(n24313), .Z(n24309) );
  AND U29044 ( .A(n24315), .B(n24316), .Z(n24300) );
  NANDN U29045 ( .A(n24317), .B(n24318), .Z(n24316) );
  NANDN U29046 ( .A(n24319), .B(n24320), .Z(n24318) );
  NANDN U29047 ( .A(n24320), .B(n24319), .Z(n24315) );
  XOR U29048 ( .A(n24314), .B(n24321), .Z(N28159) );
  XOR U29049 ( .A(n24311), .B(n24313), .Z(n24321) );
  XNOR U29050 ( .A(n24307), .B(n24322), .Z(n24313) );
  XNOR U29051 ( .A(n24305), .B(n24308), .Z(n24322) );
  NAND U29052 ( .A(n24323), .B(n24324), .Z(n24308) );
  NAND U29053 ( .A(n24325), .B(n24326), .Z(n24324) );
  OR U29054 ( .A(n24327), .B(n24328), .Z(n24325) );
  NANDN U29055 ( .A(n24329), .B(n24327), .Z(n24323) );
  IV U29056 ( .A(n24328), .Z(n24329) );
  NAND U29057 ( .A(n24330), .B(n24331), .Z(n24305) );
  NAND U29058 ( .A(n24332), .B(n24333), .Z(n24331) );
  NANDN U29059 ( .A(n24334), .B(n24335), .Z(n24332) );
  NANDN U29060 ( .A(n24335), .B(n24334), .Z(n24330) );
  AND U29061 ( .A(n24336), .B(n24337), .Z(n24307) );
  NAND U29062 ( .A(n24338), .B(n24339), .Z(n24337) );
  OR U29063 ( .A(n24340), .B(n24341), .Z(n24338) );
  NANDN U29064 ( .A(n24342), .B(n24340), .Z(n24336) );
  NAND U29065 ( .A(n24343), .B(n24344), .Z(n24311) );
  NANDN U29066 ( .A(n24345), .B(n24346), .Z(n24344) );
  OR U29067 ( .A(n24347), .B(n24348), .Z(n24346) );
  NANDN U29068 ( .A(n24349), .B(n24347), .Z(n24343) );
  IV U29069 ( .A(n24348), .Z(n24349) );
  XNOR U29070 ( .A(n24319), .B(n24350), .Z(n24314) );
  XNOR U29071 ( .A(n24317), .B(n24320), .Z(n24350) );
  NAND U29072 ( .A(n24351), .B(n24352), .Z(n24320) );
  NAND U29073 ( .A(n24353), .B(n24354), .Z(n24352) );
  OR U29074 ( .A(n24355), .B(n24356), .Z(n24353) );
  NANDN U29075 ( .A(n24357), .B(n24355), .Z(n24351) );
  IV U29076 ( .A(n24356), .Z(n24357) );
  NAND U29077 ( .A(n24358), .B(n24359), .Z(n24317) );
  NAND U29078 ( .A(n24360), .B(n24361), .Z(n24359) );
  NANDN U29079 ( .A(n24362), .B(n24363), .Z(n24360) );
  NANDN U29080 ( .A(n24363), .B(n24362), .Z(n24358) );
  AND U29081 ( .A(n24364), .B(n24365), .Z(n24319) );
  NAND U29082 ( .A(n24366), .B(n24367), .Z(n24365) );
  OR U29083 ( .A(n24368), .B(n24369), .Z(n24366) );
  NANDN U29084 ( .A(n24370), .B(n24368), .Z(n24364) );
  XNOR U29085 ( .A(n24345), .B(n24371), .Z(N28158) );
  XOR U29086 ( .A(n24347), .B(n24348), .Z(n24371) );
  XNOR U29087 ( .A(n24361), .B(n24372), .Z(n24348) );
  XOR U29088 ( .A(n24362), .B(n24363), .Z(n24372) );
  XOR U29089 ( .A(n24368), .B(n24373), .Z(n24363) );
  XOR U29090 ( .A(n24367), .B(n24370), .Z(n24373) );
  IV U29091 ( .A(n24369), .Z(n24370) );
  NAND U29092 ( .A(n24374), .B(n24375), .Z(n24369) );
  OR U29093 ( .A(n24376), .B(n24377), .Z(n24375) );
  OR U29094 ( .A(n24378), .B(n24379), .Z(n24374) );
  NAND U29095 ( .A(n24380), .B(n24381), .Z(n24367) );
  OR U29096 ( .A(n24382), .B(n24383), .Z(n24381) );
  OR U29097 ( .A(n24384), .B(n24385), .Z(n24380) );
  NOR U29098 ( .A(n24386), .B(n24387), .Z(n24368) );
  ANDN U29099 ( .B(n24388), .A(n24389), .Z(n24362) );
  XNOR U29100 ( .A(n24355), .B(n24390), .Z(n24361) );
  XNOR U29101 ( .A(n24354), .B(n24356), .Z(n24390) );
  NAND U29102 ( .A(n24391), .B(n24392), .Z(n24356) );
  OR U29103 ( .A(n24393), .B(n24394), .Z(n24392) );
  OR U29104 ( .A(n24395), .B(n24396), .Z(n24391) );
  NAND U29105 ( .A(n24397), .B(n24398), .Z(n24354) );
  OR U29106 ( .A(n24399), .B(n24400), .Z(n24398) );
  OR U29107 ( .A(n24401), .B(n24402), .Z(n24397) );
  ANDN U29108 ( .B(n24403), .A(n24404), .Z(n24355) );
  IV U29109 ( .A(n24405), .Z(n24403) );
  ANDN U29110 ( .B(n24406), .A(n24407), .Z(n24347) );
  XOR U29111 ( .A(n24333), .B(n24408), .Z(n24345) );
  XOR U29112 ( .A(n24334), .B(n24335), .Z(n24408) );
  XOR U29113 ( .A(n24340), .B(n24409), .Z(n24335) );
  XOR U29114 ( .A(n24339), .B(n24342), .Z(n24409) );
  IV U29115 ( .A(n24341), .Z(n24342) );
  NAND U29116 ( .A(n24410), .B(n24411), .Z(n24341) );
  OR U29117 ( .A(n24412), .B(n24413), .Z(n24411) );
  OR U29118 ( .A(n24414), .B(n24415), .Z(n24410) );
  NAND U29119 ( .A(n24416), .B(n24417), .Z(n24339) );
  OR U29120 ( .A(n24418), .B(n24419), .Z(n24417) );
  OR U29121 ( .A(n24420), .B(n24421), .Z(n24416) );
  NOR U29122 ( .A(n24422), .B(n24423), .Z(n24340) );
  ANDN U29123 ( .B(n24424), .A(n24425), .Z(n24334) );
  IV U29124 ( .A(n24426), .Z(n24424) );
  XNOR U29125 ( .A(n24327), .B(n24427), .Z(n24333) );
  XNOR U29126 ( .A(n24326), .B(n24328), .Z(n24427) );
  NAND U29127 ( .A(n24428), .B(n24429), .Z(n24328) );
  OR U29128 ( .A(n24430), .B(n24431), .Z(n24429) );
  OR U29129 ( .A(n24432), .B(n24433), .Z(n24428) );
  NAND U29130 ( .A(n24434), .B(n24435), .Z(n24326) );
  OR U29131 ( .A(n24436), .B(n24437), .Z(n24435) );
  OR U29132 ( .A(n24438), .B(n24439), .Z(n24434) );
  ANDN U29133 ( .B(n24440), .A(n24441), .Z(n24327) );
  IV U29134 ( .A(n24442), .Z(n24440) );
  XNOR U29135 ( .A(n24407), .B(n24406), .Z(N28157) );
  XOR U29136 ( .A(n24426), .B(n24425), .Z(n24406) );
  XNOR U29137 ( .A(n24441), .B(n24442), .Z(n24425) );
  XNOR U29138 ( .A(n24436), .B(n24437), .Z(n24442) );
  XNOR U29139 ( .A(n24438), .B(n24439), .Z(n24437) );
  XNOR U29140 ( .A(y[460]), .B(x[460]), .Z(n24439) );
  XNOR U29141 ( .A(y[461]), .B(x[461]), .Z(n24438) );
  XNOR U29142 ( .A(y[459]), .B(x[459]), .Z(n24436) );
  XNOR U29143 ( .A(n24430), .B(n24431), .Z(n24441) );
  XNOR U29144 ( .A(y[456]), .B(x[456]), .Z(n24431) );
  XNOR U29145 ( .A(n24432), .B(n24433), .Z(n24430) );
  XNOR U29146 ( .A(y[457]), .B(x[457]), .Z(n24433) );
  XNOR U29147 ( .A(y[458]), .B(x[458]), .Z(n24432) );
  XNOR U29148 ( .A(n24423), .B(n24422), .Z(n24426) );
  XNOR U29149 ( .A(n24418), .B(n24419), .Z(n24422) );
  XNOR U29150 ( .A(y[453]), .B(x[453]), .Z(n24419) );
  XNOR U29151 ( .A(n24420), .B(n24421), .Z(n24418) );
  XNOR U29152 ( .A(y[454]), .B(x[454]), .Z(n24421) );
  XNOR U29153 ( .A(y[455]), .B(x[455]), .Z(n24420) );
  XNOR U29154 ( .A(n24412), .B(n24413), .Z(n24423) );
  XNOR U29155 ( .A(y[450]), .B(x[450]), .Z(n24413) );
  XNOR U29156 ( .A(n24414), .B(n24415), .Z(n24412) );
  XNOR U29157 ( .A(y[451]), .B(x[451]), .Z(n24415) );
  XNOR U29158 ( .A(y[452]), .B(x[452]), .Z(n24414) );
  XOR U29159 ( .A(n24388), .B(n24389), .Z(n24407) );
  XNOR U29160 ( .A(n24404), .B(n24405), .Z(n24389) );
  XNOR U29161 ( .A(n24399), .B(n24400), .Z(n24405) );
  XNOR U29162 ( .A(n24401), .B(n24402), .Z(n24400) );
  XNOR U29163 ( .A(y[448]), .B(x[448]), .Z(n24402) );
  XNOR U29164 ( .A(y[449]), .B(x[449]), .Z(n24401) );
  XNOR U29165 ( .A(y[447]), .B(x[447]), .Z(n24399) );
  XNOR U29166 ( .A(n24393), .B(n24394), .Z(n24404) );
  XNOR U29167 ( .A(y[444]), .B(x[444]), .Z(n24394) );
  XNOR U29168 ( .A(n24395), .B(n24396), .Z(n24393) );
  XNOR U29169 ( .A(y[445]), .B(x[445]), .Z(n24396) );
  XNOR U29170 ( .A(y[446]), .B(x[446]), .Z(n24395) );
  XOR U29171 ( .A(n24387), .B(n24386), .Z(n24388) );
  XNOR U29172 ( .A(n24382), .B(n24383), .Z(n24386) );
  XNOR U29173 ( .A(y[441]), .B(x[441]), .Z(n24383) );
  XNOR U29174 ( .A(n24384), .B(n24385), .Z(n24382) );
  XNOR U29175 ( .A(y[442]), .B(x[442]), .Z(n24385) );
  XNOR U29176 ( .A(y[443]), .B(x[443]), .Z(n24384) );
  XNOR U29177 ( .A(n24376), .B(n24377), .Z(n24387) );
  XNOR U29178 ( .A(y[438]), .B(x[438]), .Z(n24377) );
  XNOR U29179 ( .A(n24378), .B(n24379), .Z(n24376) );
  XNOR U29180 ( .A(y[439]), .B(x[439]), .Z(n24379) );
  XNOR U29181 ( .A(y[440]), .B(x[440]), .Z(n24378) );
  NAND U29182 ( .A(n24443), .B(n24444), .Z(N28149) );
  NANDN U29183 ( .A(n24445), .B(n24446), .Z(n24444) );
  OR U29184 ( .A(n24447), .B(n24448), .Z(n24446) );
  NAND U29185 ( .A(n24447), .B(n24448), .Z(n24443) );
  XOR U29186 ( .A(n24447), .B(n24449), .Z(N28148) );
  XNOR U29187 ( .A(n24445), .B(n24448), .Z(n24449) );
  AND U29188 ( .A(n24450), .B(n24451), .Z(n24448) );
  NANDN U29189 ( .A(n24452), .B(n24453), .Z(n24451) );
  NANDN U29190 ( .A(n24454), .B(n24455), .Z(n24453) );
  NANDN U29191 ( .A(n24455), .B(n24454), .Z(n24450) );
  NAND U29192 ( .A(n24456), .B(n24457), .Z(n24445) );
  NANDN U29193 ( .A(n24458), .B(n24459), .Z(n24457) );
  OR U29194 ( .A(n24460), .B(n24461), .Z(n24459) );
  NAND U29195 ( .A(n24461), .B(n24460), .Z(n24456) );
  AND U29196 ( .A(n24462), .B(n24463), .Z(n24447) );
  NANDN U29197 ( .A(n24464), .B(n24465), .Z(n24463) );
  NANDN U29198 ( .A(n24466), .B(n24467), .Z(n24465) );
  NANDN U29199 ( .A(n24467), .B(n24466), .Z(n24462) );
  XOR U29200 ( .A(n24461), .B(n24468), .Z(N28147) );
  XOR U29201 ( .A(n24458), .B(n24460), .Z(n24468) );
  XNOR U29202 ( .A(n24454), .B(n24469), .Z(n24460) );
  XNOR U29203 ( .A(n24452), .B(n24455), .Z(n24469) );
  NAND U29204 ( .A(n24470), .B(n24471), .Z(n24455) );
  NAND U29205 ( .A(n24472), .B(n24473), .Z(n24471) );
  OR U29206 ( .A(n24474), .B(n24475), .Z(n24472) );
  NANDN U29207 ( .A(n24476), .B(n24474), .Z(n24470) );
  IV U29208 ( .A(n24475), .Z(n24476) );
  NAND U29209 ( .A(n24477), .B(n24478), .Z(n24452) );
  NAND U29210 ( .A(n24479), .B(n24480), .Z(n24478) );
  NANDN U29211 ( .A(n24481), .B(n24482), .Z(n24479) );
  NANDN U29212 ( .A(n24482), .B(n24481), .Z(n24477) );
  AND U29213 ( .A(n24483), .B(n24484), .Z(n24454) );
  NAND U29214 ( .A(n24485), .B(n24486), .Z(n24484) );
  OR U29215 ( .A(n24487), .B(n24488), .Z(n24485) );
  NANDN U29216 ( .A(n24489), .B(n24487), .Z(n24483) );
  NAND U29217 ( .A(n24490), .B(n24491), .Z(n24458) );
  NANDN U29218 ( .A(n24492), .B(n24493), .Z(n24491) );
  OR U29219 ( .A(n24494), .B(n24495), .Z(n24493) );
  NANDN U29220 ( .A(n24496), .B(n24494), .Z(n24490) );
  IV U29221 ( .A(n24495), .Z(n24496) );
  XNOR U29222 ( .A(n24466), .B(n24497), .Z(n24461) );
  XNOR U29223 ( .A(n24464), .B(n24467), .Z(n24497) );
  NAND U29224 ( .A(n24498), .B(n24499), .Z(n24467) );
  NAND U29225 ( .A(n24500), .B(n24501), .Z(n24499) );
  OR U29226 ( .A(n24502), .B(n24503), .Z(n24500) );
  NANDN U29227 ( .A(n24504), .B(n24502), .Z(n24498) );
  IV U29228 ( .A(n24503), .Z(n24504) );
  NAND U29229 ( .A(n24505), .B(n24506), .Z(n24464) );
  NAND U29230 ( .A(n24507), .B(n24508), .Z(n24506) );
  NANDN U29231 ( .A(n24509), .B(n24510), .Z(n24507) );
  NANDN U29232 ( .A(n24510), .B(n24509), .Z(n24505) );
  AND U29233 ( .A(n24511), .B(n24512), .Z(n24466) );
  NAND U29234 ( .A(n24513), .B(n24514), .Z(n24512) );
  OR U29235 ( .A(n24515), .B(n24516), .Z(n24513) );
  NANDN U29236 ( .A(n24517), .B(n24515), .Z(n24511) );
  XNOR U29237 ( .A(n24492), .B(n24518), .Z(N28146) );
  XOR U29238 ( .A(n24494), .B(n24495), .Z(n24518) );
  XNOR U29239 ( .A(n24508), .B(n24519), .Z(n24495) );
  XOR U29240 ( .A(n24509), .B(n24510), .Z(n24519) );
  XOR U29241 ( .A(n24515), .B(n24520), .Z(n24510) );
  XOR U29242 ( .A(n24514), .B(n24517), .Z(n24520) );
  IV U29243 ( .A(n24516), .Z(n24517) );
  NAND U29244 ( .A(n24521), .B(n24522), .Z(n24516) );
  OR U29245 ( .A(n24523), .B(n24524), .Z(n24522) );
  OR U29246 ( .A(n24525), .B(n24526), .Z(n24521) );
  NAND U29247 ( .A(n24527), .B(n24528), .Z(n24514) );
  OR U29248 ( .A(n24529), .B(n24530), .Z(n24528) );
  OR U29249 ( .A(n24531), .B(n24532), .Z(n24527) );
  NOR U29250 ( .A(n24533), .B(n24534), .Z(n24515) );
  ANDN U29251 ( .B(n24535), .A(n24536), .Z(n24509) );
  XNOR U29252 ( .A(n24502), .B(n24537), .Z(n24508) );
  XNOR U29253 ( .A(n24501), .B(n24503), .Z(n24537) );
  NAND U29254 ( .A(n24538), .B(n24539), .Z(n24503) );
  OR U29255 ( .A(n24540), .B(n24541), .Z(n24539) );
  OR U29256 ( .A(n24542), .B(n24543), .Z(n24538) );
  NAND U29257 ( .A(n24544), .B(n24545), .Z(n24501) );
  OR U29258 ( .A(n24546), .B(n24547), .Z(n24545) );
  OR U29259 ( .A(n24548), .B(n24549), .Z(n24544) );
  ANDN U29260 ( .B(n24550), .A(n24551), .Z(n24502) );
  IV U29261 ( .A(n24552), .Z(n24550) );
  ANDN U29262 ( .B(n24553), .A(n24554), .Z(n24494) );
  XOR U29263 ( .A(n24480), .B(n24555), .Z(n24492) );
  XOR U29264 ( .A(n24481), .B(n24482), .Z(n24555) );
  XOR U29265 ( .A(n24487), .B(n24556), .Z(n24482) );
  XOR U29266 ( .A(n24486), .B(n24489), .Z(n24556) );
  IV U29267 ( .A(n24488), .Z(n24489) );
  NAND U29268 ( .A(n24557), .B(n24558), .Z(n24488) );
  OR U29269 ( .A(n24559), .B(n24560), .Z(n24558) );
  OR U29270 ( .A(n24561), .B(n24562), .Z(n24557) );
  NAND U29271 ( .A(n24563), .B(n24564), .Z(n24486) );
  OR U29272 ( .A(n24565), .B(n24566), .Z(n24564) );
  OR U29273 ( .A(n24567), .B(n24568), .Z(n24563) );
  NOR U29274 ( .A(n24569), .B(n24570), .Z(n24487) );
  ANDN U29275 ( .B(n24571), .A(n24572), .Z(n24481) );
  IV U29276 ( .A(n24573), .Z(n24571) );
  XNOR U29277 ( .A(n24474), .B(n24574), .Z(n24480) );
  XNOR U29278 ( .A(n24473), .B(n24475), .Z(n24574) );
  NAND U29279 ( .A(n24575), .B(n24576), .Z(n24475) );
  OR U29280 ( .A(n24577), .B(n24578), .Z(n24576) );
  OR U29281 ( .A(n24579), .B(n24580), .Z(n24575) );
  NAND U29282 ( .A(n24581), .B(n24582), .Z(n24473) );
  OR U29283 ( .A(n24583), .B(n24584), .Z(n24582) );
  OR U29284 ( .A(n24585), .B(n24586), .Z(n24581) );
  ANDN U29285 ( .B(n24587), .A(n24588), .Z(n24474) );
  IV U29286 ( .A(n24589), .Z(n24587) );
  XNOR U29287 ( .A(n24554), .B(n24553), .Z(N28145) );
  XOR U29288 ( .A(n24573), .B(n24572), .Z(n24553) );
  XNOR U29289 ( .A(n24588), .B(n24589), .Z(n24572) );
  XNOR U29290 ( .A(n24583), .B(n24584), .Z(n24589) );
  XNOR U29291 ( .A(n24585), .B(n24586), .Z(n24584) );
  XNOR U29292 ( .A(y[436]), .B(x[436]), .Z(n24586) );
  XNOR U29293 ( .A(y[437]), .B(x[437]), .Z(n24585) );
  XNOR U29294 ( .A(y[435]), .B(x[435]), .Z(n24583) );
  XNOR U29295 ( .A(n24577), .B(n24578), .Z(n24588) );
  XNOR U29296 ( .A(y[432]), .B(x[432]), .Z(n24578) );
  XNOR U29297 ( .A(n24579), .B(n24580), .Z(n24577) );
  XNOR U29298 ( .A(y[433]), .B(x[433]), .Z(n24580) );
  XNOR U29299 ( .A(y[434]), .B(x[434]), .Z(n24579) );
  XNOR U29300 ( .A(n24570), .B(n24569), .Z(n24573) );
  XNOR U29301 ( .A(n24565), .B(n24566), .Z(n24569) );
  XNOR U29302 ( .A(y[429]), .B(x[429]), .Z(n24566) );
  XNOR U29303 ( .A(n24567), .B(n24568), .Z(n24565) );
  XNOR U29304 ( .A(y[430]), .B(x[430]), .Z(n24568) );
  XNOR U29305 ( .A(y[431]), .B(x[431]), .Z(n24567) );
  XNOR U29306 ( .A(n24559), .B(n24560), .Z(n24570) );
  XNOR U29307 ( .A(y[426]), .B(x[426]), .Z(n24560) );
  XNOR U29308 ( .A(n24561), .B(n24562), .Z(n24559) );
  XNOR U29309 ( .A(y[427]), .B(x[427]), .Z(n24562) );
  XNOR U29310 ( .A(y[428]), .B(x[428]), .Z(n24561) );
  XOR U29311 ( .A(n24535), .B(n24536), .Z(n24554) );
  XNOR U29312 ( .A(n24551), .B(n24552), .Z(n24536) );
  XNOR U29313 ( .A(n24546), .B(n24547), .Z(n24552) );
  XNOR U29314 ( .A(n24548), .B(n24549), .Z(n24547) );
  XNOR U29315 ( .A(y[424]), .B(x[424]), .Z(n24549) );
  XNOR U29316 ( .A(y[425]), .B(x[425]), .Z(n24548) );
  XNOR U29317 ( .A(y[423]), .B(x[423]), .Z(n24546) );
  XNOR U29318 ( .A(n24540), .B(n24541), .Z(n24551) );
  XNOR U29319 ( .A(y[420]), .B(x[420]), .Z(n24541) );
  XNOR U29320 ( .A(n24542), .B(n24543), .Z(n24540) );
  XNOR U29321 ( .A(y[421]), .B(x[421]), .Z(n24543) );
  XNOR U29322 ( .A(y[422]), .B(x[422]), .Z(n24542) );
  XOR U29323 ( .A(n24534), .B(n24533), .Z(n24535) );
  XNOR U29324 ( .A(n24529), .B(n24530), .Z(n24533) );
  XNOR U29325 ( .A(y[417]), .B(x[417]), .Z(n24530) );
  XNOR U29326 ( .A(n24531), .B(n24532), .Z(n24529) );
  XNOR U29327 ( .A(y[418]), .B(x[418]), .Z(n24532) );
  XNOR U29328 ( .A(y[419]), .B(x[419]), .Z(n24531) );
  XNOR U29329 ( .A(n24523), .B(n24524), .Z(n24534) );
  XNOR U29330 ( .A(y[414]), .B(x[414]), .Z(n24524) );
  XNOR U29331 ( .A(n24525), .B(n24526), .Z(n24523) );
  XNOR U29332 ( .A(y[415]), .B(x[415]), .Z(n24526) );
  XNOR U29333 ( .A(y[416]), .B(x[416]), .Z(n24525) );
  NAND U29334 ( .A(n24590), .B(n24591), .Z(N28137) );
  NANDN U29335 ( .A(n24592), .B(n24593), .Z(n24591) );
  OR U29336 ( .A(n24594), .B(n24595), .Z(n24593) );
  NAND U29337 ( .A(n24594), .B(n24595), .Z(n24590) );
  XOR U29338 ( .A(n24594), .B(n24596), .Z(N28136) );
  XNOR U29339 ( .A(n24592), .B(n24595), .Z(n24596) );
  AND U29340 ( .A(n24597), .B(n24598), .Z(n24595) );
  NANDN U29341 ( .A(n24599), .B(n24600), .Z(n24598) );
  NANDN U29342 ( .A(n24601), .B(n24602), .Z(n24600) );
  NANDN U29343 ( .A(n24602), .B(n24601), .Z(n24597) );
  NAND U29344 ( .A(n24603), .B(n24604), .Z(n24592) );
  NANDN U29345 ( .A(n24605), .B(n24606), .Z(n24604) );
  OR U29346 ( .A(n24607), .B(n24608), .Z(n24606) );
  NAND U29347 ( .A(n24608), .B(n24607), .Z(n24603) );
  AND U29348 ( .A(n24609), .B(n24610), .Z(n24594) );
  NANDN U29349 ( .A(n24611), .B(n24612), .Z(n24610) );
  NANDN U29350 ( .A(n24613), .B(n24614), .Z(n24612) );
  NANDN U29351 ( .A(n24614), .B(n24613), .Z(n24609) );
  XOR U29352 ( .A(n24608), .B(n24615), .Z(N28135) );
  XOR U29353 ( .A(n24605), .B(n24607), .Z(n24615) );
  XNOR U29354 ( .A(n24601), .B(n24616), .Z(n24607) );
  XNOR U29355 ( .A(n24599), .B(n24602), .Z(n24616) );
  NAND U29356 ( .A(n24617), .B(n24618), .Z(n24602) );
  NAND U29357 ( .A(n24619), .B(n24620), .Z(n24618) );
  OR U29358 ( .A(n24621), .B(n24622), .Z(n24619) );
  NANDN U29359 ( .A(n24623), .B(n24621), .Z(n24617) );
  IV U29360 ( .A(n24622), .Z(n24623) );
  NAND U29361 ( .A(n24624), .B(n24625), .Z(n24599) );
  NAND U29362 ( .A(n24626), .B(n24627), .Z(n24625) );
  NANDN U29363 ( .A(n24628), .B(n24629), .Z(n24626) );
  NANDN U29364 ( .A(n24629), .B(n24628), .Z(n24624) );
  AND U29365 ( .A(n24630), .B(n24631), .Z(n24601) );
  NAND U29366 ( .A(n24632), .B(n24633), .Z(n24631) );
  OR U29367 ( .A(n24634), .B(n24635), .Z(n24632) );
  NANDN U29368 ( .A(n24636), .B(n24634), .Z(n24630) );
  NAND U29369 ( .A(n24637), .B(n24638), .Z(n24605) );
  NANDN U29370 ( .A(n24639), .B(n24640), .Z(n24638) );
  OR U29371 ( .A(n24641), .B(n24642), .Z(n24640) );
  NANDN U29372 ( .A(n24643), .B(n24641), .Z(n24637) );
  IV U29373 ( .A(n24642), .Z(n24643) );
  XNOR U29374 ( .A(n24613), .B(n24644), .Z(n24608) );
  XNOR U29375 ( .A(n24611), .B(n24614), .Z(n24644) );
  NAND U29376 ( .A(n24645), .B(n24646), .Z(n24614) );
  NAND U29377 ( .A(n24647), .B(n24648), .Z(n24646) );
  OR U29378 ( .A(n24649), .B(n24650), .Z(n24647) );
  NANDN U29379 ( .A(n24651), .B(n24649), .Z(n24645) );
  IV U29380 ( .A(n24650), .Z(n24651) );
  NAND U29381 ( .A(n24652), .B(n24653), .Z(n24611) );
  NAND U29382 ( .A(n24654), .B(n24655), .Z(n24653) );
  NANDN U29383 ( .A(n24656), .B(n24657), .Z(n24654) );
  NANDN U29384 ( .A(n24657), .B(n24656), .Z(n24652) );
  AND U29385 ( .A(n24658), .B(n24659), .Z(n24613) );
  NAND U29386 ( .A(n24660), .B(n24661), .Z(n24659) );
  OR U29387 ( .A(n24662), .B(n24663), .Z(n24660) );
  NANDN U29388 ( .A(n24664), .B(n24662), .Z(n24658) );
  XNOR U29389 ( .A(n24639), .B(n24665), .Z(N28134) );
  XOR U29390 ( .A(n24641), .B(n24642), .Z(n24665) );
  XNOR U29391 ( .A(n24655), .B(n24666), .Z(n24642) );
  XOR U29392 ( .A(n24656), .B(n24657), .Z(n24666) );
  XOR U29393 ( .A(n24662), .B(n24667), .Z(n24657) );
  XOR U29394 ( .A(n24661), .B(n24664), .Z(n24667) );
  IV U29395 ( .A(n24663), .Z(n24664) );
  NAND U29396 ( .A(n24668), .B(n24669), .Z(n24663) );
  OR U29397 ( .A(n24670), .B(n24671), .Z(n24669) );
  OR U29398 ( .A(n24672), .B(n24673), .Z(n24668) );
  NAND U29399 ( .A(n24674), .B(n24675), .Z(n24661) );
  OR U29400 ( .A(n24676), .B(n24677), .Z(n24675) );
  OR U29401 ( .A(n24678), .B(n24679), .Z(n24674) );
  NOR U29402 ( .A(n24680), .B(n24681), .Z(n24662) );
  ANDN U29403 ( .B(n24682), .A(n24683), .Z(n24656) );
  XNOR U29404 ( .A(n24649), .B(n24684), .Z(n24655) );
  XNOR U29405 ( .A(n24648), .B(n24650), .Z(n24684) );
  NAND U29406 ( .A(n24685), .B(n24686), .Z(n24650) );
  OR U29407 ( .A(n24687), .B(n24688), .Z(n24686) );
  OR U29408 ( .A(n24689), .B(n24690), .Z(n24685) );
  NAND U29409 ( .A(n24691), .B(n24692), .Z(n24648) );
  OR U29410 ( .A(n24693), .B(n24694), .Z(n24692) );
  OR U29411 ( .A(n24695), .B(n24696), .Z(n24691) );
  ANDN U29412 ( .B(n24697), .A(n24698), .Z(n24649) );
  IV U29413 ( .A(n24699), .Z(n24697) );
  ANDN U29414 ( .B(n24700), .A(n24701), .Z(n24641) );
  XOR U29415 ( .A(n24627), .B(n24702), .Z(n24639) );
  XOR U29416 ( .A(n24628), .B(n24629), .Z(n24702) );
  XOR U29417 ( .A(n24634), .B(n24703), .Z(n24629) );
  XOR U29418 ( .A(n24633), .B(n24636), .Z(n24703) );
  IV U29419 ( .A(n24635), .Z(n24636) );
  NAND U29420 ( .A(n24704), .B(n24705), .Z(n24635) );
  OR U29421 ( .A(n24706), .B(n24707), .Z(n24705) );
  OR U29422 ( .A(n24708), .B(n24709), .Z(n24704) );
  NAND U29423 ( .A(n24710), .B(n24711), .Z(n24633) );
  OR U29424 ( .A(n24712), .B(n24713), .Z(n24711) );
  OR U29425 ( .A(n24714), .B(n24715), .Z(n24710) );
  NOR U29426 ( .A(n24716), .B(n24717), .Z(n24634) );
  ANDN U29427 ( .B(n24718), .A(n24719), .Z(n24628) );
  IV U29428 ( .A(n24720), .Z(n24718) );
  XNOR U29429 ( .A(n24621), .B(n24721), .Z(n24627) );
  XNOR U29430 ( .A(n24620), .B(n24622), .Z(n24721) );
  NAND U29431 ( .A(n24722), .B(n24723), .Z(n24622) );
  OR U29432 ( .A(n24724), .B(n24725), .Z(n24723) );
  OR U29433 ( .A(n24726), .B(n24727), .Z(n24722) );
  NAND U29434 ( .A(n24728), .B(n24729), .Z(n24620) );
  OR U29435 ( .A(n24730), .B(n24731), .Z(n24729) );
  OR U29436 ( .A(n24732), .B(n24733), .Z(n24728) );
  ANDN U29437 ( .B(n24734), .A(n24735), .Z(n24621) );
  IV U29438 ( .A(n24736), .Z(n24734) );
  XNOR U29439 ( .A(n24701), .B(n24700), .Z(N28133) );
  XOR U29440 ( .A(n24720), .B(n24719), .Z(n24700) );
  XNOR U29441 ( .A(n24735), .B(n24736), .Z(n24719) );
  XNOR U29442 ( .A(n24730), .B(n24731), .Z(n24736) );
  XNOR U29443 ( .A(n24732), .B(n24733), .Z(n24731) );
  XNOR U29444 ( .A(y[412]), .B(x[412]), .Z(n24733) );
  XNOR U29445 ( .A(y[413]), .B(x[413]), .Z(n24732) );
  XNOR U29446 ( .A(y[411]), .B(x[411]), .Z(n24730) );
  XNOR U29447 ( .A(n24724), .B(n24725), .Z(n24735) );
  XNOR U29448 ( .A(y[408]), .B(x[408]), .Z(n24725) );
  XNOR U29449 ( .A(n24726), .B(n24727), .Z(n24724) );
  XNOR U29450 ( .A(y[409]), .B(x[409]), .Z(n24727) );
  XNOR U29451 ( .A(y[410]), .B(x[410]), .Z(n24726) );
  XNOR U29452 ( .A(n24717), .B(n24716), .Z(n24720) );
  XNOR U29453 ( .A(n24712), .B(n24713), .Z(n24716) );
  XNOR U29454 ( .A(y[405]), .B(x[405]), .Z(n24713) );
  XNOR U29455 ( .A(n24714), .B(n24715), .Z(n24712) );
  XNOR U29456 ( .A(y[406]), .B(x[406]), .Z(n24715) );
  XNOR U29457 ( .A(y[407]), .B(x[407]), .Z(n24714) );
  XNOR U29458 ( .A(n24706), .B(n24707), .Z(n24717) );
  XNOR U29459 ( .A(y[402]), .B(x[402]), .Z(n24707) );
  XNOR U29460 ( .A(n24708), .B(n24709), .Z(n24706) );
  XNOR U29461 ( .A(y[403]), .B(x[403]), .Z(n24709) );
  XNOR U29462 ( .A(y[404]), .B(x[404]), .Z(n24708) );
  XOR U29463 ( .A(n24682), .B(n24683), .Z(n24701) );
  XNOR U29464 ( .A(n24698), .B(n24699), .Z(n24683) );
  XNOR U29465 ( .A(n24693), .B(n24694), .Z(n24699) );
  XNOR U29466 ( .A(n24695), .B(n24696), .Z(n24694) );
  XNOR U29467 ( .A(y[400]), .B(x[400]), .Z(n24696) );
  XNOR U29468 ( .A(y[401]), .B(x[401]), .Z(n24695) );
  XNOR U29469 ( .A(y[399]), .B(x[399]), .Z(n24693) );
  XNOR U29470 ( .A(n24687), .B(n24688), .Z(n24698) );
  XNOR U29471 ( .A(y[396]), .B(x[396]), .Z(n24688) );
  XNOR U29472 ( .A(n24689), .B(n24690), .Z(n24687) );
  XNOR U29473 ( .A(y[397]), .B(x[397]), .Z(n24690) );
  XNOR U29474 ( .A(y[398]), .B(x[398]), .Z(n24689) );
  XOR U29475 ( .A(n24681), .B(n24680), .Z(n24682) );
  XNOR U29476 ( .A(n24676), .B(n24677), .Z(n24680) );
  XNOR U29477 ( .A(y[393]), .B(x[393]), .Z(n24677) );
  XNOR U29478 ( .A(n24678), .B(n24679), .Z(n24676) );
  XNOR U29479 ( .A(y[394]), .B(x[394]), .Z(n24679) );
  XNOR U29480 ( .A(y[395]), .B(x[395]), .Z(n24678) );
  XNOR U29481 ( .A(n24670), .B(n24671), .Z(n24681) );
  XNOR U29482 ( .A(y[390]), .B(x[390]), .Z(n24671) );
  XNOR U29483 ( .A(n24672), .B(n24673), .Z(n24670) );
  XNOR U29484 ( .A(y[391]), .B(x[391]), .Z(n24673) );
  XNOR U29485 ( .A(y[392]), .B(x[392]), .Z(n24672) );
  NAND U29486 ( .A(n24737), .B(n24738), .Z(N28125) );
  NANDN U29487 ( .A(n24739), .B(n24740), .Z(n24738) );
  OR U29488 ( .A(n24741), .B(n24742), .Z(n24740) );
  NAND U29489 ( .A(n24741), .B(n24742), .Z(n24737) );
  XOR U29490 ( .A(n24741), .B(n24743), .Z(N28124) );
  XNOR U29491 ( .A(n24739), .B(n24742), .Z(n24743) );
  AND U29492 ( .A(n24744), .B(n24745), .Z(n24742) );
  NANDN U29493 ( .A(n24746), .B(n24747), .Z(n24745) );
  NANDN U29494 ( .A(n24748), .B(n24749), .Z(n24747) );
  NANDN U29495 ( .A(n24749), .B(n24748), .Z(n24744) );
  NAND U29496 ( .A(n24750), .B(n24751), .Z(n24739) );
  NANDN U29497 ( .A(n24752), .B(n24753), .Z(n24751) );
  OR U29498 ( .A(n24754), .B(n24755), .Z(n24753) );
  NAND U29499 ( .A(n24755), .B(n24754), .Z(n24750) );
  AND U29500 ( .A(n24756), .B(n24757), .Z(n24741) );
  NANDN U29501 ( .A(n24758), .B(n24759), .Z(n24757) );
  NANDN U29502 ( .A(n24760), .B(n24761), .Z(n24759) );
  NANDN U29503 ( .A(n24761), .B(n24760), .Z(n24756) );
  XOR U29504 ( .A(n24755), .B(n24762), .Z(N28123) );
  XOR U29505 ( .A(n24752), .B(n24754), .Z(n24762) );
  XNOR U29506 ( .A(n24748), .B(n24763), .Z(n24754) );
  XNOR U29507 ( .A(n24746), .B(n24749), .Z(n24763) );
  NAND U29508 ( .A(n24764), .B(n24765), .Z(n24749) );
  NAND U29509 ( .A(n24766), .B(n24767), .Z(n24765) );
  OR U29510 ( .A(n24768), .B(n24769), .Z(n24766) );
  NANDN U29511 ( .A(n24770), .B(n24768), .Z(n24764) );
  IV U29512 ( .A(n24769), .Z(n24770) );
  NAND U29513 ( .A(n24771), .B(n24772), .Z(n24746) );
  NAND U29514 ( .A(n24773), .B(n24774), .Z(n24772) );
  NANDN U29515 ( .A(n24775), .B(n24776), .Z(n24773) );
  NANDN U29516 ( .A(n24776), .B(n24775), .Z(n24771) );
  AND U29517 ( .A(n24777), .B(n24778), .Z(n24748) );
  NAND U29518 ( .A(n24779), .B(n24780), .Z(n24778) );
  OR U29519 ( .A(n24781), .B(n24782), .Z(n24779) );
  NANDN U29520 ( .A(n24783), .B(n24781), .Z(n24777) );
  NAND U29521 ( .A(n24784), .B(n24785), .Z(n24752) );
  NANDN U29522 ( .A(n24786), .B(n24787), .Z(n24785) );
  OR U29523 ( .A(n24788), .B(n24789), .Z(n24787) );
  NANDN U29524 ( .A(n24790), .B(n24788), .Z(n24784) );
  IV U29525 ( .A(n24789), .Z(n24790) );
  XNOR U29526 ( .A(n24760), .B(n24791), .Z(n24755) );
  XNOR U29527 ( .A(n24758), .B(n24761), .Z(n24791) );
  NAND U29528 ( .A(n24792), .B(n24793), .Z(n24761) );
  NAND U29529 ( .A(n24794), .B(n24795), .Z(n24793) );
  OR U29530 ( .A(n24796), .B(n24797), .Z(n24794) );
  NANDN U29531 ( .A(n24798), .B(n24796), .Z(n24792) );
  IV U29532 ( .A(n24797), .Z(n24798) );
  NAND U29533 ( .A(n24799), .B(n24800), .Z(n24758) );
  NAND U29534 ( .A(n24801), .B(n24802), .Z(n24800) );
  NANDN U29535 ( .A(n24803), .B(n24804), .Z(n24801) );
  NANDN U29536 ( .A(n24804), .B(n24803), .Z(n24799) );
  AND U29537 ( .A(n24805), .B(n24806), .Z(n24760) );
  NAND U29538 ( .A(n24807), .B(n24808), .Z(n24806) );
  OR U29539 ( .A(n24809), .B(n24810), .Z(n24807) );
  NANDN U29540 ( .A(n24811), .B(n24809), .Z(n24805) );
  XNOR U29541 ( .A(n24786), .B(n24812), .Z(N28122) );
  XOR U29542 ( .A(n24788), .B(n24789), .Z(n24812) );
  XNOR U29543 ( .A(n24802), .B(n24813), .Z(n24789) );
  XOR U29544 ( .A(n24803), .B(n24804), .Z(n24813) );
  XOR U29545 ( .A(n24809), .B(n24814), .Z(n24804) );
  XOR U29546 ( .A(n24808), .B(n24811), .Z(n24814) );
  IV U29547 ( .A(n24810), .Z(n24811) );
  NAND U29548 ( .A(n24815), .B(n24816), .Z(n24810) );
  OR U29549 ( .A(n24817), .B(n24818), .Z(n24816) );
  OR U29550 ( .A(n24819), .B(n24820), .Z(n24815) );
  NAND U29551 ( .A(n24821), .B(n24822), .Z(n24808) );
  OR U29552 ( .A(n24823), .B(n24824), .Z(n24822) );
  OR U29553 ( .A(n24825), .B(n24826), .Z(n24821) );
  NOR U29554 ( .A(n24827), .B(n24828), .Z(n24809) );
  ANDN U29555 ( .B(n24829), .A(n24830), .Z(n24803) );
  XNOR U29556 ( .A(n24796), .B(n24831), .Z(n24802) );
  XNOR U29557 ( .A(n24795), .B(n24797), .Z(n24831) );
  NAND U29558 ( .A(n24832), .B(n24833), .Z(n24797) );
  OR U29559 ( .A(n24834), .B(n24835), .Z(n24833) );
  OR U29560 ( .A(n24836), .B(n24837), .Z(n24832) );
  NAND U29561 ( .A(n24838), .B(n24839), .Z(n24795) );
  OR U29562 ( .A(n24840), .B(n24841), .Z(n24839) );
  OR U29563 ( .A(n24842), .B(n24843), .Z(n24838) );
  ANDN U29564 ( .B(n24844), .A(n24845), .Z(n24796) );
  IV U29565 ( .A(n24846), .Z(n24844) );
  ANDN U29566 ( .B(n24847), .A(n24848), .Z(n24788) );
  XOR U29567 ( .A(n24774), .B(n24849), .Z(n24786) );
  XOR U29568 ( .A(n24775), .B(n24776), .Z(n24849) );
  XOR U29569 ( .A(n24781), .B(n24850), .Z(n24776) );
  XOR U29570 ( .A(n24780), .B(n24783), .Z(n24850) );
  IV U29571 ( .A(n24782), .Z(n24783) );
  NAND U29572 ( .A(n24851), .B(n24852), .Z(n24782) );
  OR U29573 ( .A(n24853), .B(n24854), .Z(n24852) );
  OR U29574 ( .A(n24855), .B(n24856), .Z(n24851) );
  NAND U29575 ( .A(n24857), .B(n24858), .Z(n24780) );
  OR U29576 ( .A(n24859), .B(n24860), .Z(n24858) );
  OR U29577 ( .A(n24861), .B(n24862), .Z(n24857) );
  NOR U29578 ( .A(n24863), .B(n24864), .Z(n24781) );
  ANDN U29579 ( .B(n24865), .A(n24866), .Z(n24775) );
  IV U29580 ( .A(n24867), .Z(n24865) );
  XNOR U29581 ( .A(n24768), .B(n24868), .Z(n24774) );
  XNOR U29582 ( .A(n24767), .B(n24769), .Z(n24868) );
  NAND U29583 ( .A(n24869), .B(n24870), .Z(n24769) );
  OR U29584 ( .A(n24871), .B(n24872), .Z(n24870) );
  OR U29585 ( .A(n24873), .B(n24874), .Z(n24869) );
  NAND U29586 ( .A(n24875), .B(n24876), .Z(n24767) );
  OR U29587 ( .A(n24877), .B(n24878), .Z(n24876) );
  OR U29588 ( .A(n24879), .B(n24880), .Z(n24875) );
  ANDN U29589 ( .B(n24881), .A(n24882), .Z(n24768) );
  IV U29590 ( .A(n24883), .Z(n24881) );
  XNOR U29591 ( .A(n24848), .B(n24847), .Z(N28121) );
  XOR U29592 ( .A(n24867), .B(n24866), .Z(n24847) );
  XNOR U29593 ( .A(n24882), .B(n24883), .Z(n24866) );
  XNOR U29594 ( .A(n24877), .B(n24878), .Z(n24883) );
  XNOR U29595 ( .A(n24879), .B(n24880), .Z(n24878) );
  XNOR U29596 ( .A(y[388]), .B(x[388]), .Z(n24880) );
  XNOR U29597 ( .A(y[389]), .B(x[389]), .Z(n24879) );
  XNOR U29598 ( .A(y[387]), .B(x[387]), .Z(n24877) );
  XNOR U29599 ( .A(n24871), .B(n24872), .Z(n24882) );
  XNOR U29600 ( .A(y[384]), .B(x[384]), .Z(n24872) );
  XNOR U29601 ( .A(n24873), .B(n24874), .Z(n24871) );
  XNOR U29602 ( .A(y[385]), .B(x[385]), .Z(n24874) );
  XNOR U29603 ( .A(y[386]), .B(x[386]), .Z(n24873) );
  XNOR U29604 ( .A(n24864), .B(n24863), .Z(n24867) );
  XNOR U29605 ( .A(n24859), .B(n24860), .Z(n24863) );
  XNOR U29606 ( .A(y[381]), .B(x[381]), .Z(n24860) );
  XNOR U29607 ( .A(n24861), .B(n24862), .Z(n24859) );
  XNOR U29608 ( .A(y[382]), .B(x[382]), .Z(n24862) );
  XNOR U29609 ( .A(y[383]), .B(x[383]), .Z(n24861) );
  XNOR U29610 ( .A(n24853), .B(n24854), .Z(n24864) );
  XNOR U29611 ( .A(y[378]), .B(x[378]), .Z(n24854) );
  XNOR U29612 ( .A(n24855), .B(n24856), .Z(n24853) );
  XNOR U29613 ( .A(y[379]), .B(x[379]), .Z(n24856) );
  XNOR U29614 ( .A(y[380]), .B(x[380]), .Z(n24855) );
  XOR U29615 ( .A(n24829), .B(n24830), .Z(n24848) );
  XNOR U29616 ( .A(n24845), .B(n24846), .Z(n24830) );
  XNOR U29617 ( .A(n24840), .B(n24841), .Z(n24846) );
  XNOR U29618 ( .A(n24842), .B(n24843), .Z(n24841) );
  XNOR U29619 ( .A(y[376]), .B(x[376]), .Z(n24843) );
  XNOR U29620 ( .A(y[377]), .B(x[377]), .Z(n24842) );
  XNOR U29621 ( .A(y[375]), .B(x[375]), .Z(n24840) );
  XNOR U29622 ( .A(n24834), .B(n24835), .Z(n24845) );
  XNOR U29623 ( .A(y[372]), .B(x[372]), .Z(n24835) );
  XNOR U29624 ( .A(n24836), .B(n24837), .Z(n24834) );
  XNOR U29625 ( .A(y[373]), .B(x[373]), .Z(n24837) );
  XNOR U29626 ( .A(y[374]), .B(x[374]), .Z(n24836) );
  XOR U29627 ( .A(n24828), .B(n24827), .Z(n24829) );
  XNOR U29628 ( .A(n24823), .B(n24824), .Z(n24827) );
  XNOR U29629 ( .A(y[369]), .B(x[369]), .Z(n24824) );
  XNOR U29630 ( .A(n24825), .B(n24826), .Z(n24823) );
  XNOR U29631 ( .A(y[370]), .B(x[370]), .Z(n24826) );
  XNOR U29632 ( .A(y[371]), .B(x[371]), .Z(n24825) );
  XNOR U29633 ( .A(n24817), .B(n24818), .Z(n24828) );
  XNOR U29634 ( .A(y[366]), .B(x[366]), .Z(n24818) );
  XNOR U29635 ( .A(n24819), .B(n24820), .Z(n24817) );
  XNOR U29636 ( .A(y[367]), .B(x[367]), .Z(n24820) );
  XNOR U29637 ( .A(y[368]), .B(x[368]), .Z(n24819) );
  NAND U29638 ( .A(n24884), .B(n24885), .Z(N28113) );
  NANDN U29639 ( .A(n24886), .B(n24887), .Z(n24885) );
  OR U29640 ( .A(n24888), .B(n24889), .Z(n24887) );
  NAND U29641 ( .A(n24888), .B(n24889), .Z(n24884) );
  XOR U29642 ( .A(n24888), .B(n24890), .Z(N28112) );
  XNOR U29643 ( .A(n24886), .B(n24889), .Z(n24890) );
  AND U29644 ( .A(n24891), .B(n24892), .Z(n24889) );
  NANDN U29645 ( .A(n24893), .B(n24894), .Z(n24892) );
  NANDN U29646 ( .A(n24895), .B(n24896), .Z(n24894) );
  NANDN U29647 ( .A(n24896), .B(n24895), .Z(n24891) );
  NAND U29648 ( .A(n24897), .B(n24898), .Z(n24886) );
  NANDN U29649 ( .A(n24899), .B(n24900), .Z(n24898) );
  OR U29650 ( .A(n24901), .B(n24902), .Z(n24900) );
  NAND U29651 ( .A(n24902), .B(n24901), .Z(n24897) );
  AND U29652 ( .A(n24903), .B(n24904), .Z(n24888) );
  NANDN U29653 ( .A(n24905), .B(n24906), .Z(n24904) );
  NANDN U29654 ( .A(n24907), .B(n24908), .Z(n24906) );
  NANDN U29655 ( .A(n24908), .B(n24907), .Z(n24903) );
  XOR U29656 ( .A(n24902), .B(n24909), .Z(N28111) );
  XOR U29657 ( .A(n24899), .B(n24901), .Z(n24909) );
  XNOR U29658 ( .A(n24895), .B(n24910), .Z(n24901) );
  XNOR U29659 ( .A(n24893), .B(n24896), .Z(n24910) );
  NAND U29660 ( .A(n24911), .B(n24912), .Z(n24896) );
  NAND U29661 ( .A(n24913), .B(n24914), .Z(n24912) );
  OR U29662 ( .A(n24915), .B(n24916), .Z(n24913) );
  NANDN U29663 ( .A(n24917), .B(n24915), .Z(n24911) );
  IV U29664 ( .A(n24916), .Z(n24917) );
  NAND U29665 ( .A(n24918), .B(n24919), .Z(n24893) );
  NAND U29666 ( .A(n24920), .B(n24921), .Z(n24919) );
  NANDN U29667 ( .A(n24922), .B(n24923), .Z(n24920) );
  NANDN U29668 ( .A(n24923), .B(n24922), .Z(n24918) );
  AND U29669 ( .A(n24924), .B(n24925), .Z(n24895) );
  NAND U29670 ( .A(n24926), .B(n24927), .Z(n24925) );
  OR U29671 ( .A(n24928), .B(n24929), .Z(n24926) );
  NANDN U29672 ( .A(n24930), .B(n24928), .Z(n24924) );
  NAND U29673 ( .A(n24931), .B(n24932), .Z(n24899) );
  NANDN U29674 ( .A(n24933), .B(n24934), .Z(n24932) );
  OR U29675 ( .A(n24935), .B(n24936), .Z(n24934) );
  NANDN U29676 ( .A(n24937), .B(n24935), .Z(n24931) );
  IV U29677 ( .A(n24936), .Z(n24937) );
  XNOR U29678 ( .A(n24907), .B(n24938), .Z(n24902) );
  XNOR U29679 ( .A(n24905), .B(n24908), .Z(n24938) );
  NAND U29680 ( .A(n24939), .B(n24940), .Z(n24908) );
  NAND U29681 ( .A(n24941), .B(n24942), .Z(n24940) );
  OR U29682 ( .A(n24943), .B(n24944), .Z(n24941) );
  NANDN U29683 ( .A(n24945), .B(n24943), .Z(n24939) );
  IV U29684 ( .A(n24944), .Z(n24945) );
  NAND U29685 ( .A(n24946), .B(n24947), .Z(n24905) );
  NAND U29686 ( .A(n24948), .B(n24949), .Z(n24947) );
  NANDN U29687 ( .A(n24950), .B(n24951), .Z(n24948) );
  NANDN U29688 ( .A(n24951), .B(n24950), .Z(n24946) );
  AND U29689 ( .A(n24952), .B(n24953), .Z(n24907) );
  NAND U29690 ( .A(n24954), .B(n24955), .Z(n24953) );
  OR U29691 ( .A(n24956), .B(n24957), .Z(n24954) );
  NANDN U29692 ( .A(n24958), .B(n24956), .Z(n24952) );
  XNOR U29693 ( .A(n24933), .B(n24959), .Z(N28110) );
  XOR U29694 ( .A(n24935), .B(n24936), .Z(n24959) );
  XNOR U29695 ( .A(n24949), .B(n24960), .Z(n24936) );
  XOR U29696 ( .A(n24950), .B(n24951), .Z(n24960) );
  XOR U29697 ( .A(n24956), .B(n24961), .Z(n24951) );
  XOR U29698 ( .A(n24955), .B(n24958), .Z(n24961) );
  IV U29699 ( .A(n24957), .Z(n24958) );
  NAND U29700 ( .A(n24962), .B(n24963), .Z(n24957) );
  OR U29701 ( .A(n24964), .B(n24965), .Z(n24963) );
  OR U29702 ( .A(n24966), .B(n24967), .Z(n24962) );
  NAND U29703 ( .A(n24968), .B(n24969), .Z(n24955) );
  OR U29704 ( .A(n24970), .B(n24971), .Z(n24969) );
  OR U29705 ( .A(n24972), .B(n24973), .Z(n24968) );
  NOR U29706 ( .A(n24974), .B(n24975), .Z(n24956) );
  ANDN U29707 ( .B(n24976), .A(n24977), .Z(n24950) );
  XNOR U29708 ( .A(n24943), .B(n24978), .Z(n24949) );
  XNOR U29709 ( .A(n24942), .B(n24944), .Z(n24978) );
  NAND U29710 ( .A(n24979), .B(n24980), .Z(n24944) );
  OR U29711 ( .A(n24981), .B(n24982), .Z(n24980) );
  OR U29712 ( .A(n24983), .B(n24984), .Z(n24979) );
  NAND U29713 ( .A(n24985), .B(n24986), .Z(n24942) );
  OR U29714 ( .A(n24987), .B(n24988), .Z(n24986) );
  OR U29715 ( .A(n24989), .B(n24990), .Z(n24985) );
  ANDN U29716 ( .B(n24991), .A(n24992), .Z(n24943) );
  IV U29717 ( .A(n24993), .Z(n24991) );
  ANDN U29718 ( .B(n24994), .A(n24995), .Z(n24935) );
  XOR U29719 ( .A(n24921), .B(n24996), .Z(n24933) );
  XOR U29720 ( .A(n24922), .B(n24923), .Z(n24996) );
  XOR U29721 ( .A(n24928), .B(n24997), .Z(n24923) );
  XOR U29722 ( .A(n24927), .B(n24930), .Z(n24997) );
  IV U29723 ( .A(n24929), .Z(n24930) );
  NAND U29724 ( .A(n24998), .B(n24999), .Z(n24929) );
  OR U29725 ( .A(n25000), .B(n25001), .Z(n24999) );
  OR U29726 ( .A(n25002), .B(n25003), .Z(n24998) );
  NAND U29727 ( .A(n25004), .B(n25005), .Z(n24927) );
  OR U29728 ( .A(n25006), .B(n25007), .Z(n25005) );
  OR U29729 ( .A(n25008), .B(n25009), .Z(n25004) );
  NOR U29730 ( .A(n25010), .B(n25011), .Z(n24928) );
  ANDN U29731 ( .B(n25012), .A(n25013), .Z(n24922) );
  IV U29732 ( .A(n25014), .Z(n25012) );
  XNOR U29733 ( .A(n24915), .B(n25015), .Z(n24921) );
  XNOR U29734 ( .A(n24914), .B(n24916), .Z(n25015) );
  NAND U29735 ( .A(n25016), .B(n25017), .Z(n24916) );
  OR U29736 ( .A(n25018), .B(n25019), .Z(n25017) );
  OR U29737 ( .A(n25020), .B(n25021), .Z(n25016) );
  NAND U29738 ( .A(n25022), .B(n25023), .Z(n24914) );
  OR U29739 ( .A(n25024), .B(n25025), .Z(n25023) );
  OR U29740 ( .A(n25026), .B(n25027), .Z(n25022) );
  ANDN U29741 ( .B(n25028), .A(n25029), .Z(n24915) );
  IV U29742 ( .A(n25030), .Z(n25028) );
  XNOR U29743 ( .A(n24995), .B(n24994), .Z(N28109) );
  XOR U29744 ( .A(n25014), .B(n25013), .Z(n24994) );
  XNOR U29745 ( .A(n25029), .B(n25030), .Z(n25013) );
  XNOR U29746 ( .A(n25024), .B(n25025), .Z(n25030) );
  XNOR U29747 ( .A(n25026), .B(n25027), .Z(n25025) );
  XNOR U29748 ( .A(y[364]), .B(x[364]), .Z(n25027) );
  XNOR U29749 ( .A(y[365]), .B(x[365]), .Z(n25026) );
  XNOR U29750 ( .A(y[363]), .B(x[363]), .Z(n25024) );
  XNOR U29751 ( .A(n25018), .B(n25019), .Z(n25029) );
  XNOR U29752 ( .A(y[360]), .B(x[360]), .Z(n25019) );
  XNOR U29753 ( .A(n25020), .B(n25021), .Z(n25018) );
  XNOR U29754 ( .A(y[361]), .B(x[361]), .Z(n25021) );
  XNOR U29755 ( .A(y[362]), .B(x[362]), .Z(n25020) );
  XNOR U29756 ( .A(n25011), .B(n25010), .Z(n25014) );
  XNOR U29757 ( .A(n25006), .B(n25007), .Z(n25010) );
  XNOR U29758 ( .A(y[357]), .B(x[357]), .Z(n25007) );
  XNOR U29759 ( .A(n25008), .B(n25009), .Z(n25006) );
  XNOR U29760 ( .A(y[358]), .B(x[358]), .Z(n25009) );
  XNOR U29761 ( .A(y[359]), .B(x[359]), .Z(n25008) );
  XNOR U29762 ( .A(n25000), .B(n25001), .Z(n25011) );
  XNOR U29763 ( .A(y[354]), .B(x[354]), .Z(n25001) );
  XNOR U29764 ( .A(n25002), .B(n25003), .Z(n25000) );
  XNOR U29765 ( .A(y[355]), .B(x[355]), .Z(n25003) );
  XNOR U29766 ( .A(y[356]), .B(x[356]), .Z(n25002) );
  XOR U29767 ( .A(n24976), .B(n24977), .Z(n24995) );
  XNOR U29768 ( .A(n24992), .B(n24993), .Z(n24977) );
  XNOR U29769 ( .A(n24987), .B(n24988), .Z(n24993) );
  XNOR U29770 ( .A(n24989), .B(n24990), .Z(n24988) );
  XNOR U29771 ( .A(y[352]), .B(x[352]), .Z(n24990) );
  XNOR U29772 ( .A(y[353]), .B(x[353]), .Z(n24989) );
  XNOR U29773 ( .A(y[351]), .B(x[351]), .Z(n24987) );
  XNOR U29774 ( .A(n24981), .B(n24982), .Z(n24992) );
  XNOR U29775 ( .A(y[348]), .B(x[348]), .Z(n24982) );
  XNOR U29776 ( .A(n24983), .B(n24984), .Z(n24981) );
  XNOR U29777 ( .A(y[349]), .B(x[349]), .Z(n24984) );
  XNOR U29778 ( .A(y[350]), .B(x[350]), .Z(n24983) );
  XOR U29779 ( .A(n24975), .B(n24974), .Z(n24976) );
  XNOR U29780 ( .A(n24970), .B(n24971), .Z(n24974) );
  XNOR U29781 ( .A(y[345]), .B(x[345]), .Z(n24971) );
  XNOR U29782 ( .A(n24972), .B(n24973), .Z(n24970) );
  XNOR U29783 ( .A(y[346]), .B(x[346]), .Z(n24973) );
  XNOR U29784 ( .A(y[347]), .B(x[347]), .Z(n24972) );
  XNOR U29785 ( .A(n24964), .B(n24965), .Z(n24975) );
  XNOR U29786 ( .A(y[342]), .B(x[342]), .Z(n24965) );
  XNOR U29787 ( .A(n24966), .B(n24967), .Z(n24964) );
  XNOR U29788 ( .A(y[343]), .B(x[343]), .Z(n24967) );
  XNOR U29789 ( .A(y[344]), .B(x[344]), .Z(n24966) );
  NAND U29790 ( .A(n25031), .B(n25032), .Z(N28101) );
  NANDN U29791 ( .A(n25033), .B(n25034), .Z(n25032) );
  OR U29792 ( .A(n25035), .B(n25036), .Z(n25034) );
  NAND U29793 ( .A(n25035), .B(n25036), .Z(n25031) );
  XOR U29794 ( .A(n25035), .B(n25037), .Z(N28100) );
  XNOR U29795 ( .A(n25033), .B(n25036), .Z(n25037) );
  AND U29796 ( .A(n25038), .B(n25039), .Z(n25036) );
  NANDN U29797 ( .A(n25040), .B(n25041), .Z(n25039) );
  NANDN U29798 ( .A(n25042), .B(n25043), .Z(n25041) );
  NANDN U29799 ( .A(n25043), .B(n25042), .Z(n25038) );
  NAND U29800 ( .A(n25044), .B(n25045), .Z(n25033) );
  NANDN U29801 ( .A(n25046), .B(n25047), .Z(n25045) );
  OR U29802 ( .A(n25048), .B(n25049), .Z(n25047) );
  NAND U29803 ( .A(n25049), .B(n25048), .Z(n25044) );
  AND U29804 ( .A(n25050), .B(n25051), .Z(n25035) );
  NANDN U29805 ( .A(n25052), .B(n25053), .Z(n25051) );
  NANDN U29806 ( .A(n25054), .B(n25055), .Z(n25053) );
  NANDN U29807 ( .A(n25055), .B(n25054), .Z(n25050) );
  XOR U29808 ( .A(n25049), .B(n25056), .Z(N28099) );
  XOR U29809 ( .A(n25046), .B(n25048), .Z(n25056) );
  XNOR U29810 ( .A(n25042), .B(n25057), .Z(n25048) );
  XNOR U29811 ( .A(n25040), .B(n25043), .Z(n25057) );
  NAND U29812 ( .A(n25058), .B(n25059), .Z(n25043) );
  NAND U29813 ( .A(n25060), .B(n25061), .Z(n25059) );
  OR U29814 ( .A(n25062), .B(n25063), .Z(n25060) );
  NANDN U29815 ( .A(n25064), .B(n25062), .Z(n25058) );
  IV U29816 ( .A(n25063), .Z(n25064) );
  NAND U29817 ( .A(n25065), .B(n25066), .Z(n25040) );
  NAND U29818 ( .A(n25067), .B(n25068), .Z(n25066) );
  NANDN U29819 ( .A(n25069), .B(n25070), .Z(n25067) );
  NANDN U29820 ( .A(n25070), .B(n25069), .Z(n25065) );
  AND U29821 ( .A(n25071), .B(n25072), .Z(n25042) );
  NAND U29822 ( .A(n25073), .B(n25074), .Z(n25072) );
  OR U29823 ( .A(n25075), .B(n25076), .Z(n25073) );
  NANDN U29824 ( .A(n25077), .B(n25075), .Z(n25071) );
  NAND U29825 ( .A(n25078), .B(n25079), .Z(n25046) );
  NANDN U29826 ( .A(n25080), .B(n25081), .Z(n25079) );
  OR U29827 ( .A(n25082), .B(n25083), .Z(n25081) );
  NANDN U29828 ( .A(n25084), .B(n25082), .Z(n25078) );
  IV U29829 ( .A(n25083), .Z(n25084) );
  XNOR U29830 ( .A(n25054), .B(n25085), .Z(n25049) );
  XNOR U29831 ( .A(n25052), .B(n25055), .Z(n25085) );
  NAND U29832 ( .A(n25086), .B(n25087), .Z(n25055) );
  NAND U29833 ( .A(n25088), .B(n25089), .Z(n25087) );
  OR U29834 ( .A(n25090), .B(n25091), .Z(n25088) );
  NANDN U29835 ( .A(n25092), .B(n25090), .Z(n25086) );
  IV U29836 ( .A(n25091), .Z(n25092) );
  NAND U29837 ( .A(n25093), .B(n25094), .Z(n25052) );
  NAND U29838 ( .A(n25095), .B(n25096), .Z(n25094) );
  NANDN U29839 ( .A(n25097), .B(n25098), .Z(n25095) );
  NANDN U29840 ( .A(n25098), .B(n25097), .Z(n25093) );
  AND U29841 ( .A(n25099), .B(n25100), .Z(n25054) );
  NAND U29842 ( .A(n25101), .B(n25102), .Z(n25100) );
  OR U29843 ( .A(n25103), .B(n25104), .Z(n25101) );
  NANDN U29844 ( .A(n25105), .B(n25103), .Z(n25099) );
  XNOR U29845 ( .A(n25080), .B(n25106), .Z(N28098) );
  XOR U29846 ( .A(n25082), .B(n25083), .Z(n25106) );
  XNOR U29847 ( .A(n25096), .B(n25107), .Z(n25083) );
  XOR U29848 ( .A(n25097), .B(n25098), .Z(n25107) );
  XOR U29849 ( .A(n25103), .B(n25108), .Z(n25098) );
  XOR U29850 ( .A(n25102), .B(n25105), .Z(n25108) );
  IV U29851 ( .A(n25104), .Z(n25105) );
  NAND U29852 ( .A(n25109), .B(n25110), .Z(n25104) );
  OR U29853 ( .A(n25111), .B(n25112), .Z(n25110) );
  OR U29854 ( .A(n25113), .B(n25114), .Z(n25109) );
  NAND U29855 ( .A(n25115), .B(n25116), .Z(n25102) );
  OR U29856 ( .A(n25117), .B(n25118), .Z(n25116) );
  OR U29857 ( .A(n25119), .B(n25120), .Z(n25115) );
  NOR U29858 ( .A(n25121), .B(n25122), .Z(n25103) );
  ANDN U29859 ( .B(n25123), .A(n25124), .Z(n25097) );
  XNOR U29860 ( .A(n25090), .B(n25125), .Z(n25096) );
  XNOR U29861 ( .A(n25089), .B(n25091), .Z(n25125) );
  NAND U29862 ( .A(n25126), .B(n25127), .Z(n25091) );
  OR U29863 ( .A(n25128), .B(n25129), .Z(n25127) );
  OR U29864 ( .A(n25130), .B(n25131), .Z(n25126) );
  NAND U29865 ( .A(n25132), .B(n25133), .Z(n25089) );
  OR U29866 ( .A(n25134), .B(n25135), .Z(n25133) );
  OR U29867 ( .A(n25136), .B(n25137), .Z(n25132) );
  ANDN U29868 ( .B(n25138), .A(n25139), .Z(n25090) );
  IV U29869 ( .A(n25140), .Z(n25138) );
  ANDN U29870 ( .B(n25141), .A(n25142), .Z(n25082) );
  XOR U29871 ( .A(n25068), .B(n25143), .Z(n25080) );
  XOR U29872 ( .A(n25069), .B(n25070), .Z(n25143) );
  XOR U29873 ( .A(n25075), .B(n25144), .Z(n25070) );
  XOR U29874 ( .A(n25074), .B(n25077), .Z(n25144) );
  IV U29875 ( .A(n25076), .Z(n25077) );
  NAND U29876 ( .A(n25145), .B(n25146), .Z(n25076) );
  OR U29877 ( .A(n25147), .B(n25148), .Z(n25146) );
  OR U29878 ( .A(n25149), .B(n25150), .Z(n25145) );
  NAND U29879 ( .A(n25151), .B(n25152), .Z(n25074) );
  OR U29880 ( .A(n25153), .B(n25154), .Z(n25152) );
  OR U29881 ( .A(n25155), .B(n25156), .Z(n25151) );
  NOR U29882 ( .A(n25157), .B(n25158), .Z(n25075) );
  ANDN U29883 ( .B(n25159), .A(n25160), .Z(n25069) );
  IV U29884 ( .A(n25161), .Z(n25159) );
  XNOR U29885 ( .A(n25062), .B(n25162), .Z(n25068) );
  XNOR U29886 ( .A(n25061), .B(n25063), .Z(n25162) );
  NAND U29887 ( .A(n25163), .B(n25164), .Z(n25063) );
  OR U29888 ( .A(n25165), .B(n25166), .Z(n25164) );
  OR U29889 ( .A(n25167), .B(n25168), .Z(n25163) );
  NAND U29890 ( .A(n25169), .B(n25170), .Z(n25061) );
  OR U29891 ( .A(n25171), .B(n25172), .Z(n25170) );
  OR U29892 ( .A(n25173), .B(n25174), .Z(n25169) );
  ANDN U29893 ( .B(n25175), .A(n25176), .Z(n25062) );
  IV U29894 ( .A(n25177), .Z(n25175) );
  XNOR U29895 ( .A(n25142), .B(n25141), .Z(N28097) );
  XOR U29896 ( .A(n25161), .B(n25160), .Z(n25141) );
  XNOR U29897 ( .A(n25176), .B(n25177), .Z(n25160) );
  XNOR U29898 ( .A(n25171), .B(n25172), .Z(n25177) );
  XNOR U29899 ( .A(n25173), .B(n25174), .Z(n25172) );
  XNOR U29900 ( .A(y[340]), .B(x[340]), .Z(n25174) );
  XNOR U29901 ( .A(y[341]), .B(x[341]), .Z(n25173) );
  XNOR U29902 ( .A(y[339]), .B(x[339]), .Z(n25171) );
  XNOR U29903 ( .A(n25165), .B(n25166), .Z(n25176) );
  XNOR U29904 ( .A(y[336]), .B(x[336]), .Z(n25166) );
  XNOR U29905 ( .A(n25167), .B(n25168), .Z(n25165) );
  XNOR U29906 ( .A(y[337]), .B(x[337]), .Z(n25168) );
  XNOR U29907 ( .A(y[338]), .B(x[338]), .Z(n25167) );
  XNOR U29908 ( .A(n25158), .B(n25157), .Z(n25161) );
  XNOR U29909 ( .A(n25153), .B(n25154), .Z(n25157) );
  XNOR U29910 ( .A(y[333]), .B(x[333]), .Z(n25154) );
  XNOR U29911 ( .A(n25155), .B(n25156), .Z(n25153) );
  XNOR U29912 ( .A(y[334]), .B(x[334]), .Z(n25156) );
  XNOR U29913 ( .A(y[335]), .B(x[335]), .Z(n25155) );
  XNOR U29914 ( .A(n25147), .B(n25148), .Z(n25158) );
  XNOR U29915 ( .A(y[330]), .B(x[330]), .Z(n25148) );
  XNOR U29916 ( .A(n25149), .B(n25150), .Z(n25147) );
  XNOR U29917 ( .A(y[331]), .B(x[331]), .Z(n25150) );
  XNOR U29918 ( .A(y[332]), .B(x[332]), .Z(n25149) );
  XOR U29919 ( .A(n25123), .B(n25124), .Z(n25142) );
  XNOR U29920 ( .A(n25139), .B(n25140), .Z(n25124) );
  XNOR U29921 ( .A(n25134), .B(n25135), .Z(n25140) );
  XNOR U29922 ( .A(n25136), .B(n25137), .Z(n25135) );
  XNOR U29923 ( .A(y[328]), .B(x[328]), .Z(n25137) );
  XNOR U29924 ( .A(y[329]), .B(x[329]), .Z(n25136) );
  XNOR U29925 ( .A(y[327]), .B(x[327]), .Z(n25134) );
  XNOR U29926 ( .A(n25128), .B(n25129), .Z(n25139) );
  XNOR U29927 ( .A(y[324]), .B(x[324]), .Z(n25129) );
  XNOR U29928 ( .A(n25130), .B(n25131), .Z(n25128) );
  XNOR U29929 ( .A(y[325]), .B(x[325]), .Z(n25131) );
  XNOR U29930 ( .A(y[326]), .B(x[326]), .Z(n25130) );
  XOR U29931 ( .A(n25122), .B(n25121), .Z(n25123) );
  XNOR U29932 ( .A(n25117), .B(n25118), .Z(n25121) );
  XNOR U29933 ( .A(y[321]), .B(x[321]), .Z(n25118) );
  XNOR U29934 ( .A(n25119), .B(n25120), .Z(n25117) );
  XNOR U29935 ( .A(y[322]), .B(x[322]), .Z(n25120) );
  XNOR U29936 ( .A(y[323]), .B(x[323]), .Z(n25119) );
  XNOR U29937 ( .A(n25111), .B(n25112), .Z(n25122) );
  XNOR U29938 ( .A(y[318]), .B(x[318]), .Z(n25112) );
  XNOR U29939 ( .A(n25113), .B(n25114), .Z(n25111) );
  XNOR U29940 ( .A(y[319]), .B(x[319]), .Z(n25114) );
  XNOR U29941 ( .A(y[320]), .B(x[320]), .Z(n25113) );
  NAND U29942 ( .A(n25178), .B(n25179), .Z(N28089) );
  NANDN U29943 ( .A(n25180), .B(n25181), .Z(n25179) );
  OR U29944 ( .A(n25182), .B(n25183), .Z(n25181) );
  NAND U29945 ( .A(n25182), .B(n25183), .Z(n25178) );
  XOR U29946 ( .A(n25182), .B(n25184), .Z(N28088) );
  XNOR U29947 ( .A(n25180), .B(n25183), .Z(n25184) );
  AND U29948 ( .A(n25185), .B(n25186), .Z(n25183) );
  NANDN U29949 ( .A(n25187), .B(n25188), .Z(n25186) );
  NANDN U29950 ( .A(n25189), .B(n25190), .Z(n25188) );
  NANDN U29951 ( .A(n25190), .B(n25189), .Z(n25185) );
  NAND U29952 ( .A(n25191), .B(n25192), .Z(n25180) );
  NANDN U29953 ( .A(n25193), .B(n25194), .Z(n25192) );
  OR U29954 ( .A(n25195), .B(n25196), .Z(n25194) );
  NAND U29955 ( .A(n25196), .B(n25195), .Z(n25191) );
  AND U29956 ( .A(n25197), .B(n25198), .Z(n25182) );
  NANDN U29957 ( .A(n25199), .B(n25200), .Z(n25198) );
  NANDN U29958 ( .A(n25201), .B(n25202), .Z(n25200) );
  NANDN U29959 ( .A(n25202), .B(n25201), .Z(n25197) );
  XOR U29960 ( .A(n25196), .B(n25203), .Z(N28087) );
  XOR U29961 ( .A(n25193), .B(n25195), .Z(n25203) );
  XNOR U29962 ( .A(n25189), .B(n25204), .Z(n25195) );
  XNOR U29963 ( .A(n25187), .B(n25190), .Z(n25204) );
  NAND U29964 ( .A(n25205), .B(n25206), .Z(n25190) );
  NAND U29965 ( .A(n25207), .B(n25208), .Z(n25206) );
  OR U29966 ( .A(n25209), .B(n25210), .Z(n25207) );
  NANDN U29967 ( .A(n25211), .B(n25209), .Z(n25205) );
  IV U29968 ( .A(n25210), .Z(n25211) );
  NAND U29969 ( .A(n25212), .B(n25213), .Z(n25187) );
  NAND U29970 ( .A(n25214), .B(n25215), .Z(n25213) );
  NANDN U29971 ( .A(n25216), .B(n25217), .Z(n25214) );
  NANDN U29972 ( .A(n25217), .B(n25216), .Z(n25212) );
  AND U29973 ( .A(n25218), .B(n25219), .Z(n25189) );
  NAND U29974 ( .A(n25220), .B(n25221), .Z(n25219) );
  OR U29975 ( .A(n25222), .B(n25223), .Z(n25220) );
  NANDN U29976 ( .A(n25224), .B(n25222), .Z(n25218) );
  NAND U29977 ( .A(n25225), .B(n25226), .Z(n25193) );
  NANDN U29978 ( .A(n25227), .B(n25228), .Z(n25226) );
  OR U29979 ( .A(n25229), .B(n25230), .Z(n25228) );
  NANDN U29980 ( .A(n25231), .B(n25229), .Z(n25225) );
  IV U29981 ( .A(n25230), .Z(n25231) );
  XNOR U29982 ( .A(n25201), .B(n25232), .Z(n25196) );
  XNOR U29983 ( .A(n25199), .B(n25202), .Z(n25232) );
  NAND U29984 ( .A(n25233), .B(n25234), .Z(n25202) );
  NAND U29985 ( .A(n25235), .B(n25236), .Z(n25234) );
  OR U29986 ( .A(n25237), .B(n25238), .Z(n25235) );
  NANDN U29987 ( .A(n25239), .B(n25237), .Z(n25233) );
  IV U29988 ( .A(n25238), .Z(n25239) );
  NAND U29989 ( .A(n25240), .B(n25241), .Z(n25199) );
  NAND U29990 ( .A(n25242), .B(n25243), .Z(n25241) );
  NANDN U29991 ( .A(n25244), .B(n25245), .Z(n25242) );
  NANDN U29992 ( .A(n25245), .B(n25244), .Z(n25240) );
  AND U29993 ( .A(n25246), .B(n25247), .Z(n25201) );
  NAND U29994 ( .A(n25248), .B(n25249), .Z(n25247) );
  OR U29995 ( .A(n25250), .B(n25251), .Z(n25248) );
  NANDN U29996 ( .A(n25252), .B(n25250), .Z(n25246) );
  XNOR U29997 ( .A(n25227), .B(n25253), .Z(N28086) );
  XOR U29998 ( .A(n25229), .B(n25230), .Z(n25253) );
  XNOR U29999 ( .A(n25243), .B(n25254), .Z(n25230) );
  XOR U30000 ( .A(n25244), .B(n25245), .Z(n25254) );
  XOR U30001 ( .A(n25250), .B(n25255), .Z(n25245) );
  XOR U30002 ( .A(n25249), .B(n25252), .Z(n25255) );
  IV U30003 ( .A(n25251), .Z(n25252) );
  NAND U30004 ( .A(n25256), .B(n25257), .Z(n25251) );
  OR U30005 ( .A(n25258), .B(n25259), .Z(n25257) );
  OR U30006 ( .A(n25260), .B(n25261), .Z(n25256) );
  NAND U30007 ( .A(n25262), .B(n25263), .Z(n25249) );
  OR U30008 ( .A(n25264), .B(n25265), .Z(n25263) );
  OR U30009 ( .A(n25266), .B(n25267), .Z(n25262) );
  NOR U30010 ( .A(n25268), .B(n25269), .Z(n25250) );
  ANDN U30011 ( .B(n25270), .A(n25271), .Z(n25244) );
  XNOR U30012 ( .A(n25237), .B(n25272), .Z(n25243) );
  XNOR U30013 ( .A(n25236), .B(n25238), .Z(n25272) );
  NAND U30014 ( .A(n25273), .B(n25274), .Z(n25238) );
  OR U30015 ( .A(n25275), .B(n25276), .Z(n25274) );
  OR U30016 ( .A(n25277), .B(n25278), .Z(n25273) );
  NAND U30017 ( .A(n25279), .B(n25280), .Z(n25236) );
  OR U30018 ( .A(n25281), .B(n25282), .Z(n25280) );
  OR U30019 ( .A(n25283), .B(n25284), .Z(n25279) );
  ANDN U30020 ( .B(n25285), .A(n25286), .Z(n25237) );
  IV U30021 ( .A(n25287), .Z(n25285) );
  ANDN U30022 ( .B(n25288), .A(n25289), .Z(n25229) );
  XOR U30023 ( .A(n25215), .B(n25290), .Z(n25227) );
  XOR U30024 ( .A(n25216), .B(n25217), .Z(n25290) );
  XOR U30025 ( .A(n25222), .B(n25291), .Z(n25217) );
  XOR U30026 ( .A(n25221), .B(n25224), .Z(n25291) );
  IV U30027 ( .A(n25223), .Z(n25224) );
  NAND U30028 ( .A(n25292), .B(n25293), .Z(n25223) );
  OR U30029 ( .A(n25294), .B(n25295), .Z(n25293) );
  OR U30030 ( .A(n25296), .B(n25297), .Z(n25292) );
  NAND U30031 ( .A(n25298), .B(n25299), .Z(n25221) );
  OR U30032 ( .A(n25300), .B(n25301), .Z(n25299) );
  OR U30033 ( .A(n25302), .B(n25303), .Z(n25298) );
  NOR U30034 ( .A(n25304), .B(n25305), .Z(n25222) );
  ANDN U30035 ( .B(n25306), .A(n25307), .Z(n25216) );
  IV U30036 ( .A(n25308), .Z(n25306) );
  XNOR U30037 ( .A(n25209), .B(n25309), .Z(n25215) );
  XNOR U30038 ( .A(n25208), .B(n25210), .Z(n25309) );
  NAND U30039 ( .A(n25310), .B(n25311), .Z(n25210) );
  OR U30040 ( .A(n25312), .B(n25313), .Z(n25311) );
  OR U30041 ( .A(n25314), .B(n25315), .Z(n25310) );
  NAND U30042 ( .A(n25316), .B(n25317), .Z(n25208) );
  OR U30043 ( .A(n25318), .B(n25319), .Z(n25317) );
  OR U30044 ( .A(n25320), .B(n25321), .Z(n25316) );
  ANDN U30045 ( .B(n25322), .A(n25323), .Z(n25209) );
  IV U30046 ( .A(n25324), .Z(n25322) );
  XNOR U30047 ( .A(n25289), .B(n25288), .Z(N28085) );
  XOR U30048 ( .A(n25308), .B(n25307), .Z(n25288) );
  XNOR U30049 ( .A(n25323), .B(n25324), .Z(n25307) );
  XNOR U30050 ( .A(n25318), .B(n25319), .Z(n25324) );
  XNOR U30051 ( .A(n25320), .B(n25321), .Z(n25319) );
  XNOR U30052 ( .A(y[316]), .B(x[316]), .Z(n25321) );
  XNOR U30053 ( .A(y[317]), .B(x[317]), .Z(n25320) );
  XNOR U30054 ( .A(y[315]), .B(x[315]), .Z(n25318) );
  XNOR U30055 ( .A(n25312), .B(n25313), .Z(n25323) );
  XNOR U30056 ( .A(y[312]), .B(x[312]), .Z(n25313) );
  XNOR U30057 ( .A(n25314), .B(n25315), .Z(n25312) );
  XNOR U30058 ( .A(y[313]), .B(x[313]), .Z(n25315) );
  XNOR U30059 ( .A(y[314]), .B(x[314]), .Z(n25314) );
  XNOR U30060 ( .A(n25305), .B(n25304), .Z(n25308) );
  XNOR U30061 ( .A(n25300), .B(n25301), .Z(n25304) );
  XNOR U30062 ( .A(y[309]), .B(x[309]), .Z(n25301) );
  XNOR U30063 ( .A(n25302), .B(n25303), .Z(n25300) );
  XNOR U30064 ( .A(y[310]), .B(x[310]), .Z(n25303) );
  XNOR U30065 ( .A(y[311]), .B(x[311]), .Z(n25302) );
  XNOR U30066 ( .A(n25294), .B(n25295), .Z(n25305) );
  XNOR U30067 ( .A(y[306]), .B(x[306]), .Z(n25295) );
  XNOR U30068 ( .A(n25296), .B(n25297), .Z(n25294) );
  XNOR U30069 ( .A(y[307]), .B(x[307]), .Z(n25297) );
  XNOR U30070 ( .A(y[308]), .B(x[308]), .Z(n25296) );
  XOR U30071 ( .A(n25270), .B(n25271), .Z(n25289) );
  XNOR U30072 ( .A(n25286), .B(n25287), .Z(n25271) );
  XNOR U30073 ( .A(n25281), .B(n25282), .Z(n25287) );
  XNOR U30074 ( .A(n25283), .B(n25284), .Z(n25282) );
  XNOR U30075 ( .A(y[304]), .B(x[304]), .Z(n25284) );
  XNOR U30076 ( .A(y[305]), .B(x[305]), .Z(n25283) );
  XNOR U30077 ( .A(y[303]), .B(x[303]), .Z(n25281) );
  XNOR U30078 ( .A(n25275), .B(n25276), .Z(n25286) );
  XNOR U30079 ( .A(y[300]), .B(x[300]), .Z(n25276) );
  XNOR U30080 ( .A(n25277), .B(n25278), .Z(n25275) );
  XNOR U30081 ( .A(y[301]), .B(x[301]), .Z(n25278) );
  XNOR U30082 ( .A(y[302]), .B(x[302]), .Z(n25277) );
  XOR U30083 ( .A(n25269), .B(n25268), .Z(n25270) );
  XNOR U30084 ( .A(n25264), .B(n25265), .Z(n25268) );
  XNOR U30085 ( .A(y[297]), .B(x[297]), .Z(n25265) );
  XNOR U30086 ( .A(n25266), .B(n25267), .Z(n25264) );
  XNOR U30087 ( .A(y[298]), .B(x[298]), .Z(n25267) );
  XNOR U30088 ( .A(y[299]), .B(x[299]), .Z(n25266) );
  XNOR U30089 ( .A(n25258), .B(n25259), .Z(n25269) );
  XNOR U30090 ( .A(y[294]), .B(x[294]), .Z(n25259) );
  XNOR U30091 ( .A(n25260), .B(n25261), .Z(n25258) );
  XNOR U30092 ( .A(y[295]), .B(x[295]), .Z(n25261) );
  XNOR U30093 ( .A(y[296]), .B(x[296]), .Z(n25260) );
  NAND U30094 ( .A(n25325), .B(n25326), .Z(N28077) );
  NANDN U30095 ( .A(n25327), .B(n25328), .Z(n25326) );
  OR U30096 ( .A(n25329), .B(n25330), .Z(n25328) );
  NAND U30097 ( .A(n25329), .B(n25330), .Z(n25325) );
  XOR U30098 ( .A(n25329), .B(n25331), .Z(N28076) );
  XNOR U30099 ( .A(n25327), .B(n25330), .Z(n25331) );
  AND U30100 ( .A(n25332), .B(n25333), .Z(n25330) );
  NANDN U30101 ( .A(n25334), .B(n25335), .Z(n25333) );
  NANDN U30102 ( .A(n25336), .B(n25337), .Z(n25335) );
  NANDN U30103 ( .A(n25337), .B(n25336), .Z(n25332) );
  NAND U30104 ( .A(n25338), .B(n25339), .Z(n25327) );
  NANDN U30105 ( .A(n25340), .B(n25341), .Z(n25339) );
  OR U30106 ( .A(n25342), .B(n25343), .Z(n25341) );
  NAND U30107 ( .A(n25343), .B(n25342), .Z(n25338) );
  AND U30108 ( .A(n25344), .B(n25345), .Z(n25329) );
  NANDN U30109 ( .A(n25346), .B(n25347), .Z(n25345) );
  NANDN U30110 ( .A(n25348), .B(n25349), .Z(n25347) );
  NANDN U30111 ( .A(n25349), .B(n25348), .Z(n25344) );
  XOR U30112 ( .A(n25343), .B(n25350), .Z(N28075) );
  XOR U30113 ( .A(n25340), .B(n25342), .Z(n25350) );
  XNOR U30114 ( .A(n25336), .B(n25351), .Z(n25342) );
  XNOR U30115 ( .A(n25334), .B(n25337), .Z(n25351) );
  NAND U30116 ( .A(n25352), .B(n25353), .Z(n25337) );
  NAND U30117 ( .A(n25354), .B(n25355), .Z(n25353) );
  OR U30118 ( .A(n25356), .B(n25357), .Z(n25354) );
  NANDN U30119 ( .A(n25358), .B(n25356), .Z(n25352) );
  IV U30120 ( .A(n25357), .Z(n25358) );
  NAND U30121 ( .A(n25359), .B(n25360), .Z(n25334) );
  NAND U30122 ( .A(n25361), .B(n25362), .Z(n25360) );
  NANDN U30123 ( .A(n25363), .B(n25364), .Z(n25361) );
  NANDN U30124 ( .A(n25364), .B(n25363), .Z(n25359) );
  AND U30125 ( .A(n25365), .B(n25366), .Z(n25336) );
  NAND U30126 ( .A(n25367), .B(n25368), .Z(n25366) );
  OR U30127 ( .A(n25369), .B(n25370), .Z(n25367) );
  NANDN U30128 ( .A(n25371), .B(n25369), .Z(n25365) );
  NAND U30129 ( .A(n25372), .B(n25373), .Z(n25340) );
  NANDN U30130 ( .A(n25374), .B(n25375), .Z(n25373) );
  OR U30131 ( .A(n25376), .B(n25377), .Z(n25375) );
  NANDN U30132 ( .A(n25378), .B(n25376), .Z(n25372) );
  IV U30133 ( .A(n25377), .Z(n25378) );
  XNOR U30134 ( .A(n25348), .B(n25379), .Z(n25343) );
  XNOR U30135 ( .A(n25346), .B(n25349), .Z(n25379) );
  NAND U30136 ( .A(n25380), .B(n25381), .Z(n25349) );
  NAND U30137 ( .A(n25382), .B(n25383), .Z(n25381) );
  OR U30138 ( .A(n25384), .B(n25385), .Z(n25382) );
  NANDN U30139 ( .A(n25386), .B(n25384), .Z(n25380) );
  IV U30140 ( .A(n25385), .Z(n25386) );
  NAND U30141 ( .A(n25387), .B(n25388), .Z(n25346) );
  NAND U30142 ( .A(n25389), .B(n25390), .Z(n25388) );
  NANDN U30143 ( .A(n25391), .B(n25392), .Z(n25389) );
  NANDN U30144 ( .A(n25392), .B(n25391), .Z(n25387) );
  AND U30145 ( .A(n25393), .B(n25394), .Z(n25348) );
  NAND U30146 ( .A(n25395), .B(n25396), .Z(n25394) );
  OR U30147 ( .A(n25397), .B(n25398), .Z(n25395) );
  NANDN U30148 ( .A(n25399), .B(n25397), .Z(n25393) );
  XNOR U30149 ( .A(n25374), .B(n25400), .Z(N28074) );
  XOR U30150 ( .A(n25376), .B(n25377), .Z(n25400) );
  XNOR U30151 ( .A(n25390), .B(n25401), .Z(n25377) );
  XOR U30152 ( .A(n25391), .B(n25392), .Z(n25401) );
  XOR U30153 ( .A(n25397), .B(n25402), .Z(n25392) );
  XOR U30154 ( .A(n25396), .B(n25399), .Z(n25402) );
  IV U30155 ( .A(n25398), .Z(n25399) );
  NAND U30156 ( .A(n25403), .B(n25404), .Z(n25398) );
  OR U30157 ( .A(n25405), .B(n25406), .Z(n25404) );
  OR U30158 ( .A(n25407), .B(n25408), .Z(n25403) );
  NAND U30159 ( .A(n25409), .B(n25410), .Z(n25396) );
  OR U30160 ( .A(n25411), .B(n25412), .Z(n25410) );
  OR U30161 ( .A(n25413), .B(n25414), .Z(n25409) );
  NOR U30162 ( .A(n25415), .B(n25416), .Z(n25397) );
  ANDN U30163 ( .B(n25417), .A(n25418), .Z(n25391) );
  XNOR U30164 ( .A(n25384), .B(n25419), .Z(n25390) );
  XNOR U30165 ( .A(n25383), .B(n25385), .Z(n25419) );
  NAND U30166 ( .A(n25420), .B(n25421), .Z(n25385) );
  OR U30167 ( .A(n25422), .B(n25423), .Z(n25421) );
  OR U30168 ( .A(n25424), .B(n25425), .Z(n25420) );
  NAND U30169 ( .A(n25426), .B(n25427), .Z(n25383) );
  OR U30170 ( .A(n25428), .B(n25429), .Z(n25427) );
  OR U30171 ( .A(n25430), .B(n25431), .Z(n25426) );
  ANDN U30172 ( .B(n25432), .A(n25433), .Z(n25384) );
  IV U30173 ( .A(n25434), .Z(n25432) );
  ANDN U30174 ( .B(n25435), .A(n25436), .Z(n25376) );
  XOR U30175 ( .A(n25362), .B(n25437), .Z(n25374) );
  XOR U30176 ( .A(n25363), .B(n25364), .Z(n25437) );
  XOR U30177 ( .A(n25369), .B(n25438), .Z(n25364) );
  XOR U30178 ( .A(n25368), .B(n25371), .Z(n25438) );
  IV U30179 ( .A(n25370), .Z(n25371) );
  NAND U30180 ( .A(n25439), .B(n25440), .Z(n25370) );
  OR U30181 ( .A(n25441), .B(n25442), .Z(n25440) );
  OR U30182 ( .A(n25443), .B(n25444), .Z(n25439) );
  NAND U30183 ( .A(n25445), .B(n25446), .Z(n25368) );
  OR U30184 ( .A(n25447), .B(n25448), .Z(n25446) );
  OR U30185 ( .A(n25449), .B(n25450), .Z(n25445) );
  NOR U30186 ( .A(n25451), .B(n25452), .Z(n25369) );
  ANDN U30187 ( .B(n25453), .A(n25454), .Z(n25363) );
  IV U30188 ( .A(n25455), .Z(n25453) );
  XNOR U30189 ( .A(n25356), .B(n25456), .Z(n25362) );
  XNOR U30190 ( .A(n25355), .B(n25357), .Z(n25456) );
  NAND U30191 ( .A(n25457), .B(n25458), .Z(n25357) );
  OR U30192 ( .A(n25459), .B(n25460), .Z(n25458) );
  OR U30193 ( .A(n25461), .B(n25462), .Z(n25457) );
  NAND U30194 ( .A(n25463), .B(n25464), .Z(n25355) );
  OR U30195 ( .A(n25465), .B(n25466), .Z(n25464) );
  OR U30196 ( .A(n25467), .B(n25468), .Z(n25463) );
  ANDN U30197 ( .B(n25469), .A(n25470), .Z(n25356) );
  IV U30198 ( .A(n25471), .Z(n25469) );
  XNOR U30199 ( .A(n25436), .B(n25435), .Z(N28073) );
  XOR U30200 ( .A(n25455), .B(n25454), .Z(n25435) );
  XNOR U30201 ( .A(n25470), .B(n25471), .Z(n25454) );
  XNOR U30202 ( .A(n25465), .B(n25466), .Z(n25471) );
  XNOR U30203 ( .A(n25467), .B(n25468), .Z(n25466) );
  XNOR U30204 ( .A(y[292]), .B(x[292]), .Z(n25468) );
  XNOR U30205 ( .A(y[293]), .B(x[293]), .Z(n25467) );
  XNOR U30206 ( .A(y[291]), .B(x[291]), .Z(n25465) );
  XNOR U30207 ( .A(n25459), .B(n25460), .Z(n25470) );
  XNOR U30208 ( .A(y[288]), .B(x[288]), .Z(n25460) );
  XNOR U30209 ( .A(n25461), .B(n25462), .Z(n25459) );
  XNOR U30210 ( .A(y[289]), .B(x[289]), .Z(n25462) );
  XNOR U30211 ( .A(y[290]), .B(x[290]), .Z(n25461) );
  XNOR U30212 ( .A(n25452), .B(n25451), .Z(n25455) );
  XNOR U30213 ( .A(n25447), .B(n25448), .Z(n25451) );
  XNOR U30214 ( .A(y[285]), .B(x[285]), .Z(n25448) );
  XNOR U30215 ( .A(n25449), .B(n25450), .Z(n25447) );
  XNOR U30216 ( .A(y[286]), .B(x[286]), .Z(n25450) );
  XNOR U30217 ( .A(y[287]), .B(x[287]), .Z(n25449) );
  XNOR U30218 ( .A(n25441), .B(n25442), .Z(n25452) );
  XNOR U30219 ( .A(y[282]), .B(x[282]), .Z(n25442) );
  XNOR U30220 ( .A(n25443), .B(n25444), .Z(n25441) );
  XNOR U30221 ( .A(y[283]), .B(x[283]), .Z(n25444) );
  XNOR U30222 ( .A(y[284]), .B(x[284]), .Z(n25443) );
  XOR U30223 ( .A(n25417), .B(n25418), .Z(n25436) );
  XNOR U30224 ( .A(n25433), .B(n25434), .Z(n25418) );
  XNOR U30225 ( .A(n25428), .B(n25429), .Z(n25434) );
  XNOR U30226 ( .A(n25430), .B(n25431), .Z(n25429) );
  XNOR U30227 ( .A(y[280]), .B(x[280]), .Z(n25431) );
  XNOR U30228 ( .A(y[281]), .B(x[281]), .Z(n25430) );
  XNOR U30229 ( .A(y[279]), .B(x[279]), .Z(n25428) );
  XNOR U30230 ( .A(n25422), .B(n25423), .Z(n25433) );
  XNOR U30231 ( .A(y[276]), .B(x[276]), .Z(n25423) );
  XNOR U30232 ( .A(n25424), .B(n25425), .Z(n25422) );
  XNOR U30233 ( .A(y[277]), .B(x[277]), .Z(n25425) );
  XNOR U30234 ( .A(y[278]), .B(x[278]), .Z(n25424) );
  XOR U30235 ( .A(n25416), .B(n25415), .Z(n25417) );
  XNOR U30236 ( .A(n25411), .B(n25412), .Z(n25415) );
  XNOR U30237 ( .A(y[273]), .B(x[273]), .Z(n25412) );
  XNOR U30238 ( .A(n25413), .B(n25414), .Z(n25411) );
  XNOR U30239 ( .A(y[274]), .B(x[274]), .Z(n25414) );
  XNOR U30240 ( .A(y[275]), .B(x[275]), .Z(n25413) );
  XNOR U30241 ( .A(n25405), .B(n25406), .Z(n25416) );
  XNOR U30242 ( .A(y[270]), .B(x[270]), .Z(n25406) );
  XNOR U30243 ( .A(n25407), .B(n25408), .Z(n25405) );
  XNOR U30244 ( .A(y[271]), .B(x[271]), .Z(n25408) );
  XNOR U30245 ( .A(y[272]), .B(x[272]), .Z(n25407) );
  NAND U30246 ( .A(n25472), .B(n25473), .Z(N28065) );
  NANDN U30247 ( .A(n25474), .B(n25475), .Z(n25473) );
  OR U30248 ( .A(n25476), .B(n25477), .Z(n25475) );
  NAND U30249 ( .A(n25476), .B(n25477), .Z(n25472) );
  XOR U30250 ( .A(n25476), .B(n25478), .Z(N28064) );
  XNOR U30251 ( .A(n25474), .B(n25477), .Z(n25478) );
  AND U30252 ( .A(n25479), .B(n25480), .Z(n25477) );
  NANDN U30253 ( .A(n25481), .B(n25482), .Z(n25480) );
  NANDN U30254 ( .A(n25483), .B(n25484), .Z(n25482) );
  NANDN U30255 ( .A(n25484), .B(n25483), .Z(n25479) );
  NAND U30256 ( .A(n25485), .B(n25486), .Z(n25474) );
  NANDN U30257 ( .A(n25487), .B(n25488), .Z(n25486) );
  OR U30258 ( .A(n25489), .B(n25490), .Z(n25488) );
  NAND U30259 ( .A(n25490), .B(n25489), .Z(n25485) );
  AND U30260 ( .A(n25491), .B(n25492), .Z(n25476) );
  NANDN U30261 ( .A(n25493), .B(n25494), .Z(n25492) );
  NANDN U30262 ( .A(n25495), .B(n25496), .Z(n25494) );
  NANDN U30263 ( .A(n25496), .B(n25495), .Z(n25491) );
  XOR U30264 ( .A(n25490), .B(n25497), .Z(N28063) );
  XOR U30265 ( .A(n25487), .B(n25489), .Z(n25497) );
  XNOR U30266 ( .A(n25483), .B(n25498), .Z(n25489) );
  XNOR U30267 ( .A(n25481), .B(n25484), .Z(n25498) );
  NAND U30268 ( .A(n25499), .B(n25500), .Z(n25484) );
  NAND U30269 ( .A(n25501), .B(n25502), .Z(n25500) );
  OR U30270 ( .A(n25503), .B(n25504), .Z(n25501) );
  NANDN U30271 ( .A(n25505), .B(n25503), .Z(n25499) );
  IV U30272 ( .A(n25504), .Z(n25505) );
  NAND U30273 ( .A(n25506), .B(n25507), .Z(n25481) );
  NAND U30274 ( .A(n25508), .B(n25509), .Z(n25507) );
  NANDN U30275 ( .A(n25510), .B(n25511), .Z(n25508) );
  NANDN U30276 ( .A(n25511), .B(n25510), .Z(n25506) );
  AND U30277 ( .A(n25512), .B(n25513), .Z(n25483) );
  NAND U30278 ( .A(n25514), .B(n25515), .Z(n25513) );
  OR U30279 ( .A(n25516), .B(n25517), .Z(n25514) );
  NANDN U30280 ( .A(n25518), .B(n25516), .Z(n25512) );
  NAND U30281 ( .A(n25519), .B(n25520), .Z(n25487) );
  NANDN U30282 ( .A(n25521), .B(n25522), .Z(n25520) );
  OR U30283 ( .A(n25523), .B(n25524), .Z(n25522) );
  NANDN U30284 ( .A(n25525), .B(n25523), .Z(n25519) );
  IV U30285 ( .A(n25524), .Z(n25525) );
  XNOR U30286 ( .A(n25495), .B(n25526), .Z(n25490) );
  XNOR U30287 ( .A(n25493), .B(n25496), .Z(n25526) );
  NAND U30288 ( .A(n25527), .B(n25528), .Z(n25496) );
  NAND U30289 ( .A(n25529), .B(n25530), .Z(n25528) );
  OR U30290 ( .A(n25531), .B(n25532), .Z(n25529) );
  NANDN U30291 ( .A(n25533), .B(n25531), .Z(n25527) );
  IV U30292 ( .A(n25532), .Z(n25533) );
  NAND U30293 ( .A(n25534), .B(n25535), .Z(n25493) );
  NAND U30294 ( .A(n25536), .B(n25537), .Z(n25535) );
  NANDN U30295 ( .A(n25538), .B(n25539), .Z(n25536) );
  NANDN U30296 ( .A(n25539), .B(n25538), .Z(n25534) );
  AND U30297 ( .A(n25540), .B(n25541), .Z(n25495) );
  NAND U30298 ( .A(n25542), .B(n25543), .Z(n25541) );
  OR U30299 ( .A(n25544), .B(n25545), .Z(n25542) );
  NANDN U30300 ( .A(n25546), .B(n25544), .Z(n25540) );
  XNOR U30301 ( .A(n25521), .B(n25547), .Z(N28062) );
  XOR U30302 ( .A(n25523), .B(n25524), .Z(n25547) );
  XNOR U30303 ( .A(n25537), .B(n25548), .Z(n25524) );
  XOR U30304 ( .A(n25538), .B(n25539), .Z(n25548) );
  XOR U30305 ( .A(n25544), .B(n25549), .Z(n25539) );
  XOR U30306 ( .A(n25543), .B(n25546), .Z(n25549) );
  IV U30307 ( .A(n25545), .Z(n25546) );
  NAND U30308 ( .A(n25550), .B(n25551), .Z(n25545) );
  OR U30309 ( .A(n25552), .B(n25553), .Z(n25551) );
  OR U30310 ( .A(n25554), .B(n25555), .Z(n25550) );
  NAND U30311 ( .A(n25556), .B(n25557), .Z(n25543) );
  OR U30312 ( .A(n25558), .B(n25559), .Z(n25557) );
  OR U30313 ( .A(n25560), .B(n25561), .Z(n25556) );
  NOR U30314 ( .A(n25562), .B(n25563), .Z(n25544) );
  ANDN U30315 ( .B(n25564), .A(n25565), .Z(n25538) );
  XNOR U30316 ( .A(n25531), .B(n25566), .Z(n25537) );
  XNOR U30317 ( .A(n25530), .B(n25532), .Z(n25566) );
  NAND U30318 ( .A(n25567), .B(n25568), .Z(n25532) );
  OR U30319 ( .A(n25569), .B(n25570), .Z(n25568) );
  OR U30320 ( .A(n25571), .B(n25572), .Z(n25567) );
  NAND U30321 ( .A(n25573), .B(n25574), .Z(n25530) );
  OR U30322 ( .A(n25575), .B(n25576), .Z(n25574) );
  OR U30323 ( .A(n25577), .B(n25578), .Z(n25573) );
  ANDN U30324 ( .B(n25579), .A(n25580), .Z(n25531) );
  IV U30325 ( .A(n25581), .Z(n25579) );
  ANDN U30326 ( .B(n25582), .A(n25583), .Z(n25523) );
  XOR U30327 ( .A(n25509), .B(n25584), .Z(n25521) );
  XOR U30328 ( .A(n25510), .B(n25511), .Z(n25584) );
  XOR U30329 ( .A(n25516), .B(n25585), .Z(n25511) );
  XOR U30330 ( .A(n25515), .B(n25518), .Z(n25585) );
  IV U30331 ( .A(n25517), .Z(n25518) );
  NAND U30332 ( .A(n25586), .B(n25587), .Z(n25517) );
  OR U30333 ( .A(n25588), .B(n25589), .Z(n25587) );
  OR U30334 ( .A(n25590), .B(n25591), .Z(n25586) );
  NAND U30335 ( .A(n25592), .B(n25593), .Z(n25515) );
  OR U30336 ( .A(n25594), .B(n25595), .Z(n25593) );
  OR U30337 ( .A(n25596), .B(n25597), .Z(n25592) );
  NOR U30338 ( .A(n25598), .B(n25599), .Z(n25516) );
  ANDN U30339 ( .B(n25600), .A(n25601), .Z(n25510) );
  IV U30340 ( .A(n25602), .Z(n25600) );
  XNOR U30341 ( .A(n25503), .B(n25603), .Z(n25509) );
  XNOR U30342 ( .A(n25502), .B(n25504), .Z(n25603) );
  NAND U30343 ( .A(n25604), .B(n25605), .Z(n25504) );
  OR U30344 ( .A(n25606), .B(n25607), .Z(n25605) );
  OR U30345 ( .A(n25608), .B(n25609), .Z(n25604) );
  NAND U30346 ( .A(n25610), .B(n25611), .Z(n25502) );
  OR U30347 ( .A(n25612), .B(n25613), .Z(n25611) );
  OR U30348 ( .A(n25614), .B(n25615), .Z(n25610) );
  ANDN U30349 ( .B(n25616), .A(n25617), .Z(n25503) );
  IV U30350 ( .A(n25618), .Z(n25616) );
  XNOR U30351 ( .A(n25583), .B(n25582), .Z(N28061) );
  XOR U30352 ( .A(n25602), .B(n25601), .Z(n25582) );
  XNOR U30353 ( .A(n25617), .B(n25618), .Z(n25601) );
  XNOR U30354 ( .A(n25612), .B(n25613), .Z(n25618) );
  XNOR U30355 ( .A(n25614), .B(n25615), .Z(n25613) );
  XNOR U30356 ( .A(y[268]), .B(x[268]), .Z(n25615) );
  XNOR U30357 ( .A(y[269]), .B(x[269]), .Z(n25614) );
  XNOR U30358 ( .A(y[267]), .B(x[267]), .Z(n25612) );
  XNOR U30359 ( .A(n25606), .B(n25607), .Z(n25617) );
  XNOR U30360 ( .A(y[264]), .B(x[264]), .Z(n25607) );
  XNOR U30361 ( .A(n25608), .B(n25609), .Z(n25606) );
  XNOR U30362 ( .A(y[265]), .B(x[265]), .Z(n25609) );
  XNOR U30363 ( .A(y[266]), .B(x[266]), .Z(n25608) );
  XNOR U30364 ( .A(n25599), .B(n25598), .Z(n25602) );
  XNOR U30365 ( .A(n25594), .B(n25595), .Z(n25598) );
  XNOR U30366 ( .A(y[261]), .B(x[261]), .Z(n25595) );
  XNOR U30367 ( .A(n25596), .B(n25597), .Z(n25594) );
  XNOR U30368 ( .A(y[262]), .B(x[262]), .Z(n25597) );
  XNOR U30369 ( .A(y[263]), .B(x[263]), .Z(n25596) );
  XNOR U30370 ( .A(n25588), .B(n25589), .Z(n25599) );
  XNOR U30371 ( .A(y[258]), .B(x[258]), .Z(n25589) );
  XNOR U30372 ( .A(n25590), .B(n25591), .Z(n25588) );
  XNOR U30373 ( .A(y[259]), .B(x[259]), .Z(n25591) );
  XNOR U30374 ( .A(y[260]), .B(x[260]), .Z(n25590) );
  XOR U30375 ( .A(n25564), .B(n25565), .Z(n25583) );
  XNOR U30376 ( .A(n25580), .B(n25581), .Z(n25565) );
  XNOR U30377 ( .A(n25575), .B(n25576), .Z(n25581) );
  XNOR U30378 ( .A(n25577), .B(n25578), .Z(n25576) );
  XNOR U30379 ( .A(y[256]), .B(x[256]), .Z(n25578) );
  XNOR U30380 ( .A(y[257]), .B(x[257]), .Z(n25577) );
  XNOR U30381 ( .A(y[255]), .B(x[255]), .Z(n25575) );
  XNOR U30382 ( .A(n25569), .B(n25570), .Z(n25580) );
  XNOR U30383 ( .A(y[252]), .B(x[252]), .Z(n25570) );
  XNOR U30384 ( .A(n25571), .B(n25572), .Z(n25569) );
  XNOR U30385 ( .A(y[253]), .B(x[253]), .Z(n25572) );
  XNOR U30386 ( .A(y[254]), .B(x[254]), .Z(n25571) );
  XOR U30387 ( .A(n25563), .B(n25562), .Z(n25564) );
  XNOR U30388 ( .A(n25558), .B(n25559), .Z(n25562) );
  XNOR U30389 ( .A(y[249]), .B(x[249]), .Z(n25559) );
  XNOR U30390 ( .A(n25560), .B(n25561), .Z(n25558) );
  XNOR U30391 ( .A(y[250]), .B(x[250]), .Z(n25561) );
  XNOR U30392 ( .A(y[251]), .B(x[251]), .Z(n25560) );
  XNOR U30393 ( .A(n25552), .B(n25553), .Z(n25563) );
  XNOR U30394 ( .A(y[246]), .B(x[246]), .Z(n25553) );
  XNOR U30395 ( .A(n25554), .B(n25555), .Z(n25552) );
  XNOR U30396 ( .A(y[247]), .B(x[247]), .Z(n25555) );
  XNOR U30397 ( .A(y[248]), .B(x[248]), .Z(n25554) );
  NAND U30398 ( .A(n25619), .B(n25620), .Z(N28053) );
  NANDN U30399 ( .A(n25621), .B(n25622), .Z(n25620) );
  OR U30400 ( .A(n25623), .B(n25624), .Z(n25622) );
  NAND U30401 ( .A(n25623), .B(n25624), .Z(n25619) );
  XOR U30402 ( .A(n25623), .B(n25625), .Z(N28052) );
  XNOR U30403 ( .A(n25621), .B(n25624), .Z(n25625) );
  AND U30404 ( .A(n25626), .B(n25627), .Z(n25624) );
  NANDN U30405 ( .A(n25628), .B(n25629), .Z(n25627) );
  NANDN U30406 ( .A(n25630), .B(n25631), .Z(n25629) );
  NANDN U30407 ( .A(n25631), .B(n25630), .Z(n25626) );
  NAND U30408 ( .A(n25632), .B(n25633), .Z(n25621) );
  NANDN U30409 ( .A(n25634), .B(n25635), .Z(n25633) );
  OR U30410 ( .A(n25636), .B(n25637), .Z(n25635) );
  NAND U30411 ( .A(n25637), .B(n25636), .Z(n25632) );
  AND U30412 ( .A(n25638), .B(n25639), .Z(n25623) );
  NANDN U30413 ( .A(n25640), .B(n25641), .Z(n25639) );
  NANDN U30414 ( .A(n25642), .B(n25643), .Z(n25641) );
  NANDN U30415 ( .A(n25643), .B(n25642), .Z(n25638) );
  XOR U30416 ( .A(n25637), .B(n25644), .Z(N28051) );
  XOR U30417 ( .A(n25634), .B(n25636), .Z(n25644) );
  XNOR U30418 ( .A(n25630), .B(n25645), .Z(n25636) );
  XNOR U30419 ( .A(n25628), .B(n25631), .Z(n25645) );
  NAND U30420 ( .A(n25646), .B(n25647), .Z(n25631) );
  NAND U30421 ( .A(n25648), .B(n25649), .Z(n25647) );
  OR U30422 ( .A(n25650), .B(n25651), .Z(n25648) );
  NANDN U30423 ( .A(n25652), .B(n25650), .Z(n25646) );
  IV U30424 ( .A(n25651), .Z(n25652) );
  NAND U30425 ( .A(n25653), .B(n25654), .Z(n25628) );
  NAND U30426 ( .A(n25655), .B(n25656), .Z(n25654) );
  NANDN U30427 ( .A(n25657), .B(n25658), .Z(n25655) );
  NANDN U30428 ( .A(n25658), .B(n25657), .Z(n25653) );
  AND U30429 ( .A(n25659), .B(n25660), .Z(n25630) );
  NAND U30430 ( .A(n25661), .B(n25662), .Z(n25660) );
  OR U30431 ( .A(n25663), .B(n25664), .Z(n25661) );
  NANDN U30432 ( .A(n25665), .B(n25663), .Z(n25659) );
  NAND U30433 ( .A(n25666), .B(n25667), .Z(n25634) );
  NANDN U30434 ( .A(n25668), .B(n25669), .Z(n25667) );
  OR U30435 ( .A(n25670), .B(n25671), .Z(n25669) );
  NANDN U30436 ( .A(n25672), .B(n25670), .Z(n25666) );
  IV U30437 ( .A(n25671), .Z(n25672) );
  XNOR U30438 ( .A(n25642), .B(n25673), .Z(n25637) );
  XNOR U30439 ( .A(n25640), .B(n25643), .Z(n25673) );
  NAND U30440 ( .A(n25674), .B(n25675), .Z(n25643) );
  NAND U30441 ( .A(n25676), .B(n25677), .Z(n25675) );
  OR U30442 ( .A(n25678), .B(n25679), .Z(n25676) );
  NANDN U30443 ( .A(n25680), .B(n25678), .Z(n25674) );
  IV U30444 ( .A(n25679), .Z(n25680) );
  NAND U30445 ( .A(n25681), .B(n25682), .Z(n25640) );
  NAND U30446 ( .A(n25683), .B(n25684), .Z(n25682) );
  NANDN U30447 ( .A(n25685), .B(n25686), .Z(n25683) );
  NANDN U30448 ( .A(n25686), .B(n25685), .Z(n25681) );
  AND U30449 ( .A(n25687), .B(n25688), .Z(n25642) );
  NAND U30450 ( .A(n25689), .B(n25690), .Z(n25688) );
  OR U30451 ( .A(n25691), .B(n25692), .Z(n25689) );
  NANDN U30452 ( .A(n25693), .B(n25691), .Z(n25687) );
  XNOR U30453 ( .A(n25668), .B(n25694), .Z(N28050) );
  XOR U30454 ( .A(n25670), .B(n25671), .Z(n25694) );
  XNOR U30455 ( .A(n25684), .B(n25695), .Z(n25671) );
  XOR U30456 ( .A(n25685), .B(n25686), .Z(n25695) );
  XOR U30457 ( .A(n25691), .B(n25696), .Z(n25686) );
  XOR U30458 ( .A(n25690), .B(n25693), .Z(n25696) );
  IV U30459 ( .A(n25692), .Z(n25693) );
  NAND U30460 ( .A(n25697), .B(n25698), .Z(n25692) );
  OR U30461 ( .A(n25699), .B(n25700), .Z(n25698) );
  OR U30462 ( .A(n25701), .B(n25702), .Z(n25697) );
  NAND U30463 ( .A(n25703), .B(n25704), .Z(n25690) );
  OR U30464 ( .A(n25705), .B(n25706), .Z(n25704) );
  OR U30465 ( .A(n25707), .B(n25708), .Z(n25703) );
  NOR U30466 ( .A(n25709), .B(n25710), .Z(n25691) );
  ANDN U30467 ( .B(n25711), .A(n25712), .Z(n25685) );
  XNOR U30468 ( .A(n25678), .B(n25713), .Z(n25684) );
  XNOR U30469 ( .A(n25677), .B(n25679), .Z(n25713) );
  NAND U30470 ( .A(n25714), .B(n25715), .Z(n25679) );
  OR U30471 ( .A(n25716), .B(n25717), .Z(n25715) );
  OR U30472 ( .A(n25718), .B(n25719), .Z(n25714) );
  NAND U30473 ( .A(n25720), .B(n25721), .Z(n25677) );
  OR U30474 ( .A(n25722), .B(n25723), .Z(n25721) );
  OR U30475 ( .A(n25724), .B(n25725), .Z(n25720) );
  ANDN U30476 ( .B(n25726), .A(n25727), .Z(n25678) );
  IV U30477 ( .A(n25728), .Z(n25726) );
  ANDN U30478 ( .B(n25729), .A(n25730), .Z(n25670) );
  XOR U30479 ( .A(n25656), .B(n25731), .Z(n25668) );
  XOR U30480 ( .A(n25657), .B(n25658), .Z(n25731) );
  XOR U30481 ( .A(n25663), .B(n25732), .Z(n25658) );
  XOR U30482 ( .A(n25662), .B(n25665), .Z(n25732) );
  IV U30483 ( .A(n25664), .Z(n25665) );
  NAND U30484 ( .A(n25733), .B(n25734), .Z(n25664) );
  OR U30485 ( .A(n25735), .B(n25736), .Z(n25734) );
  OR U30486 ( .A(n25737), .B(n25738), .Z(n25733) );
  NAND U30487 ( .A(n25739), .B(n25740), .Z(n25662) );
  OR U30488 ( .A(n25741), .B(n25742), .Z(n25740) );
  OR U30489 ( .A(n25743), .B(n25744), .Z(n25739) );
  NOR U30490 ( .A(n25745), .B(n25746), .Z(n25663) );
  ANDN U30491 ( .B(n25747), .A(n25748), .Z(n25657) );
  IV U30492 ( .A(n25749), .Z(n25747) );
  XNOR U30493 ( .A(n25650), .B(n25750), .Z(n25656) );
  XNOR U30494 ( .A(n25649), .B(n25651), .Z(n25750) );
  NAND U30495 ( .A(n25751), .B(n25752), .Z(n25651) );
  OR U30496 ( .A(n25753), .B(n25754), .Z(n25752) );
  OR U30497 ( .A(n25755), .B(n25756), .Z(n25751) );
  NAND U30498 ( .A(n25757), .B(n25758), .Z(n25649) );
  OR U30499 ( .A(n25759), .B(n25760), .Z(n25758) );
  OR U30500 ( .A(n25761), .B(n25762), .Z(n25757) );
  ANDN U30501 ( .B(n25763), .A(n25764), .Z(n25650) );
  IV U30502 ( .A(n25765), .Z(n25763) );
  XNOR U30503 ( .A(n25730), .B(n25729), .Z(N28049) );
  XOR U30504 ( .A(n25749), .B(n25748), .Z(n25729) );
  XNOR U30505 ( .A(n25764), .B(n25765), .Z(n25748) );
  XNOR U30506 ( .A(n25759), .B(n25760), .Z(n25765) );
  XNOR U30507 ( .A(n25761), .B(n25762), .Z(n25760) );
  XNOR U30508 ( .A(y[244]), .B(x[244]), .Z(n25762) );
  XNOR U30509 ( .A(y[245]), .B(x[245]), .Z(n25761) );
  XNOR U30510 ( .A(y[243]), .B(x[243]), .Z(n25759) );
  XNOR U30511 ( .A(n25753), .B(n25754), .Z(n25764) );
  XNOR U30512 ( .A(y[240]), .B(x[240]), .Z(n25754) );
  XNOR U30513 ( .A(n25755), .B(n25756), .Z(n25753) );
  XNOR U30514 ( .A(y[241]), .B(x[241]), .Z(n25756) );
  XNOR U30515 ( .A(y[242]), .B(x[242]), .Z(n25755) );
  XNOR U30516 ( .A(n25746), .B(n25745), .Z(n25749) );
  XNOR U30517 ( .A(n25741), .B(n25742), .Z(n25745) );
  XNOR U30518 ( .A(y[237]), .B(x[237]), .Z(n25742) );
  XNOR U30519 ( .A(n25743), .B(n25744), .Z(n25741) );
  XNOR U30520 ( .A(y[238]), .B(x[238]), .Z(n25744) );
  XNOR U30521 ( .A(y[239]), .B(x[239]), .Z(n25743) );
  XNOR U30522 ( .A(n25735), .B(n25736), .Z(n25746) );
  XNOR U30523 ( .A(y[234]), .B(x[234]), .Z(n25736) );
  XNOR U30524 ( .A(n25737), .B(n25738), .Z(n25735) );
  XNOR U30525 ( .A(y[235]), .B(x[235]), .Z(n25738) );
  XNOR U30526 ( .A(y[236]), .B(x[236]), .Z(n25737) );
  XOR U30527 ( .A(n25711), .B(n25712), .Z(n25730) );
  XNOR U30528 ( .A(n25727), .B(n25728), .Z(n25712) );
  XNOR U30529 ( .A(n25722), .B(n25723), .Z(n25728) );
  XNOR U30530 ( .A(n25724), .B(n25725), .Z(n25723) );
  XNOR U30531 ( .A(y[232]), .B(x[232]), .Z(n25725) );
  XNOR U30532 ( .A(y[233]), .B(x[233]), .Z(n25724) );
  XNOR U30533 ( .A(y[231]), .B(x[231]), .Z(n25722) );
  XNOR U30534 ( .A(n25716), .B(n25717), .Z(n25727) );
  XNOR U30535 ( .A(y[228]), .B(x[228]), .Z(n25717) );
  XNOR U30536 ( .A(n25718), .B(n25719), .Z(n25716) );
  XNOR U30537 ( .A(y[229]), .B(x[229]), .Z(n25719) );
  XNOR U30538 ( .A(y[230]), .B(x[230]), .Z(n25718) );
  XOR U30539 ( .A(n25710), .B(n25709), .Z(n25711) );
  XNOR U30540 ( .A(n25705), .B(n25706), .Z(n25709) );
  XNOR U30541 ( .A(y[225]), .B(x[225]), .Z(n25706) );
  XNOR U30542 ( .A(n25707), .B(n25708), .Z(n25705) );
  XNOR U30543 ( .A(y[226]), .B(x[226]), .Z(n25708) );
  XNOR U30544 ( .A(y[227]), .B(x[227]), .Z(n25707) );
  XNOR U30545 ( .A(n25699), .B(n25700), .Z(n25710) );
  XNOR U30546 ( .A(y[222]), .B(x[222]), .Z(n25700) );
  XNOR U30547 ( .A(n25701), .B(n25702), .Z(n25699) );
  XNOR U30548 ( .A(y[223]), .B(x[223]), .Z(n25702) );
  XNOR U30549 ( .A(y[224]), .B(x[224]), .Z(n25701) );
  NAND U30550 ( .A(n25766), .B(n25767), .Z(N28041) );
  NANDN U30551 ( .A(n25768), .B(n25769), .Z(n25767) );
  OR U30552 ( .A(n25770), .B(n25771), .Z(n25769) );
  NAND U30553 ( .A(n25770), .B(n25771), .Z(n25766) );
  XOR U30554 ( .A(n25770), .B(n25772), .Z(N28040) );
  XNOR U30555 ( .A(n25768), .B(n25771), .Z(n25772) );
  AND U30556 ( .A(n25773), .B(n25774), .Z(n25771) );
  NANDN U30557 ( .A(n25775), .B(n25776), .Z(n25774) );
  NANDN U30558 ( .A(n25777), .B(n25778), .Z(n25776) );
  NANDN U30559 ( .A(n25778), .B(n25777), .Z(n25773) );
  NAND U30560 ( .A(n25779), .B(n25780), .Z(n25768) );
  NANDN U30561 ( .A(n25781), .B(n25782), .Z(n25780) );
  OR U30562 ( .A(n25783), .B(n25784), .Z(n25782) );
  NAND U30563 ( .A(n25784), .B(n25783), .Z(n25779) );
  AND U30564 ( .A(n25785), .B(n25786), .Z(n25770) );
  NANDN U30565 ( .A(n25787), .B(n25788), .Z(n25786) );
  NANDN U30566 ( .A(n25789), .B(n25790), .Z(n25788) );
  NANDN U30567 ( .A(n25790), .B(n25789), .Z(n25785) );
  XOR U30568 ( .A(n25784), .B(n25791), .Z(N28039) );
  XOR U30569 ( .A(n25781), .B(n25783), .Z(n25791) );
  XNOR U30570 ( .A(n25777), .B(n25792), .Z(n25783) );
  XNOR U30571 ( .A(n25775), .B(n25778), .Z(n25792) );
  NAND U30572 ( .A(n25793), .B(n25794), .Z(n25778) );
  NAND U30573 ( .A(n25795), .B(n25796), .Z(n25794) );
  OR U30574 ( .A(n25797), .B(n25798), .Z(n25795) );
  NANDN U30575 ( .A(n25799), .B(n25797), .Z(n25793) );
  IV U30576 ( .A(n25798), .Z(n25799) );
  NAND U30577 ( .A(n25800), .B(n25801), .Z(n25775) );
  NAND U30578 ( .A(n25802), .B(n25803), .Z(n25801) );
  NANDN U30579 ( .A(n25804), .B(n25805), .Z(n25802) );
  NANDN U30580 ( .A(n25805), .B(n25804), .Z(n25800) );
  AND U30581 ( .A(n25806), .B(n25807), .Z(n25777) );
  NAND U30582 ( .A(n25808), .B(n25809), .Z(n25807) );
  OR U30583 ( .A(n25810), .B(n25811), .Z(n25808) );
  NANDN U30584 ( .A(n25812), .B(n25810), .Z(n25806) );
  NAND U30585 ( .A(n25813), .B(n25814), .Z(n25781) );
  NANDN U30586 ( .A(n25815), .B(n25816), .Z(n25814) );
  OR U30587 ( .A(n25817), .B(n25818), .Z(n25816) );
  NANDN U30588 ( .A(n25819), .B(n25817), .Z(n25813) );
  IV U30589 ( .A(n25818), .Z(n25819) );
  XNOR U30590 ( .A(n25789), .B(n25820), .Z(n25784) );
  XNOR U30591 ( .A(n25787), .B(n25790), .Z(n25820) );
  NAND U30592 ( .A(n25821), .B(n25822), .Z(n25790) );
  NAND U30593 ( .A(n25823), .B(n25824), .Z(n25822) );
  OR U30594 ( .A(n25825), .B(n25826), .Z(n25823) );
  NANDN U30595 ( .A(n25827), .B(n25825), .Z(n25821) );
  IV U30596 ( .A(n25826), .Z(n25827) );
  NAND U30597 ( .A(n25828), .B(n25829), .Z(n25787) );
  NAND U30598 ( .A(n25830), .B(n25831), .Z(n25829) );
  NANDN U30599 ( .A(n25832), .B(n25833), .Z(n25830) );
  NANDN U30600 ( .A(n25833), .B(n25832), .Z(n25828) );
  AND U30601 ( .A(n25834), .B(n25835), .Z(n25789) );
  NAND U30602 ( .A(n25836), .B(n25837), .Z(n25835) );
  OR U30603 ( .A(n25838), .B(n25839), .Z(n25836) );
  NANDN U30604 ( .A(n25840), .B(n25838), .Z(n25834) );
  XNOR U30605 ( .A(n25815), .B(n25841), .Z(N28038) );
  XOR U30606 ( .A(n25817), .B(n25818), .Z(n25841) );
  XNOR U30607 ( .A(n25831), .B(n25842), .Z(n25818) );
  XOR U30608 ( .A(n25832), .B(n25833), .Z(n25842) );
  XOR U30609 ( .A(n25838), .B(n25843), .Z(n25833) );
  XOR U30610 ( .A(n25837), .B(n25840), .Z(n25843) );
  IV U30611 ( .A(n25839), .Z(n25840) );
  NAND U30612 ( .A(n25844), .B(n25845), .Z(n25839) );
  OR U30613 ( .A(n25846), .B(n25847), .Z(n25845) );
  OR U30614 ( .A(n25848), .B(n25849), .Z(n25844) );
  NAND U30615 ( .A(n25850), .B(n25851), .Z(n25837) );
  OR U30616 ( .A(n25852), .B(n25853), .Z(n25851) );
  OR U30617 ( .A(n25854), .B(n25855), .Z(n25850) );
  NOR U30618 ( .A(n25856), .B(n25857), .Z(n25838) );
  ANDN U30619 ( .B(n25858), .A(n25859), .Z(n25832) );
  XNOR U30620 ( .A(n25825), .B(n25860), .Z(n25831) );
  XNOR U30621 ( .A(n25824), .B(n25826), .Z(n25860) );
  NAND U30622 ( .A(n25861), .B(n25862), .Z(n25826) );
  OR U30623 ( .A(n25863), .B(n25864), .Z(n25862) );
  OR U30624 ( .A(n25865), .B(n25866), .Z(n25861) );
  NAND U30625 ( .A(n25867), .B(n25868), .Z(n25824) );
  OR U30626 ( .A(n25869), .B(n25870), .Z(n25868) );
  OR U30627 ( .A(n25871), .B(n25872), .Z(n25867) );
  ANDN U30628 ( .B(n25873), .A(n25874), .Z(n25825) );
  IV U30629 ( .A(n25875), .Z(n25873) );
  ANDN U30630 ( .B(n25876), .A(n25877), .Z(n25817) );
  XOR U30631 ( .A(n25803), .B(n25878), .Z(n25815) );
  XOR U30632 ( .A(n25804), .B(n25805), .Z(n25878) );
  XOR U30633 ( .A(n25810), .B(n25879), .Z(n25805) );
  XOR U30634 ( .A(n25809), .B(n25812), .Z(n25879) );
  IV U30635 ( .A(n25811), .Z(n25812) );
  NAND U30636 ( .A(n25880), .B(n25881), .Z(n25811) );
  OR U30637 ( .A(n25882), .B(n25883), .Z(n25881) );
  OR U30638 ( .A(n25884), .B(n25885), .Z(n25880) );
  NAND U30639 ( .A(n25886), .B(n25887), .Z(n25809) );
  OR U30640 ( .A(n25888), .B(n25889), .Z(n25887) );
  OR U30641 ( .A(n25890), .B(n25891), .Z(n25886) );
  NOR U30642 ( .A(n25892), .B(n25893), .Z(n25810) );
  ANDN U30643 ( .B(n25894), .A(n25895), .Z(n25804) );
  IV U30644 ( .A(n25896), .Z(n25894) );
  XNOR U30645 ( .A(n25797), .B(n25897), .Z(n25803) );
  XNOR U30646 ( .A(n25796), .B(n25798), .Z(n25897) );
  NAND U30647 ( .A(n25898), .B(n25899), .Z(n25798) );
  OR U30648 ( .A(n25900), .B(n25901), .Z(n25899) );
  OR U30649 ( .A(n25902), .B(n25903), .Z(n25898) );
  NAND U30650 ( .A(n25904), .B(n25905), .Z(n25796) );
  OR U30651 ( .A(n25906), .B(n25907), .Z(n25905) );
  OR U30652 ( .A(n25908), .B(n25909), .Z(n25904) );
  ANDN U30653 ( .B(n25910), .A(n25911), .Z(n25797) );
  IV U30654 ( .A(n25912), .Z(n25910) );
  XNOR U30655 ( .A(n25877), .B(n25876), .Z(N28037) );
  XOR U30656 ( .A(n25896), .B(n25895), .Z(n25876) );
  XNOR U30657 ( .A(n25911), .B(n25912), .Z(n25895) );
  XNOR U30658 ( .A(n25906), .B(n25907), .Z(n25912) );
  XNOR U30659 ( .A(n25908), .B(n25909), .Z(n25907) );
  XNOR U30660 ( .A(y[220]), .B(x[220]), .Z(n25909) );
  XNOR U30661 ( .A(y[221]), .B(x[221]), .Z(n25908) );
  XNOR U30662 ( .A(y[219]), .B(x[219]), .Z(n25906) );
  XNOR U30663 ( .A(n25900), .B(n25901), .Z(n25911) );
  XNOR U30664 ( .A(y[216]), .B(x[216]), .Z(n25901) );
  XNOR U30665 ( .A(n25902), .B(n25903), .Z(n25900) );
  XNOR U30666 ( .A(y[217]), .B(x[217]), .Z(n25903) );
  XNOR U30667 ( .A(y[218]), .B(x[218]), .Z(n25902) );
  XNOR U30668 ( .A(n25893), .B(n25892), .Z(n25896) );
  XNOR U30669 ( .A(n25888), .B(n25889), .Z(n25892) );
  XNOR U30670 ( .A(y[213]), .B(x[213]), .Z(n25889) );
  XNOR U30671 ( .A(n25890), .B(n25891), .Z(n25888) );
  XNOR U30672 ( .A(y[214]), .B(x[214]), .Z(n25891) );
  XNOR U30673 ( .A(y[215]), .B(x[215]), .Z(n25890) );
  XNOR U30674 ( .A(n25882), .B(n25883), .Z(n25893) );
  XNOR U30675 ( .A(y[210]), .B(x[210]), .Z(n25883) );
  XNOR U30676 ( .A(n25884), .B(n25885), .Z(n25882) );
  XNOR U30677 ( .A(y[211]), .B(x[211]), .Z(n25885) );
  XNOR U30678 ( .A(y[212]), .B(x[212]), .Z(n25884) );
  XOR U30679 ( .A(n25858), .B(n25859), .Z(n25877) );
  XNOR U30680 ( .A(n25874), .B(n25875), .Z(n25859) );
  XNOR U30681 ( .A(n25869), .B(n25870), .Z(n25875) );
  XNOR U30682 ( .A(n25871), .B(n25872), .Z(n25870) );
  XNOR U30683 ( .A(y[208]), .B(x[208]), .Z(n25872) );
  XNOR U30684 ( .A(y[209]), .B(x[209]), .Z(n25871) );
  XNOR U30685 ( .A(y[207]), .B(x[207]), .Z(n25869) );
  XNOR U30686 ( .A(n25863), .B(n25864), .Z(n25874) );
  XNOR U30687 ( .A(y[204]), .B(x[204]), .Z(n25864) );
  XNOR U30688 ( .A(n25865), .B(n25866), .Z(n25863) );
  XNOR U30689 ( .A(y[205]), .B(x[205]), .Z(n25866) );
  XNOR U30690 ( .A(y[206]), .B(x[206]), .Z(n25865) );
  XOR U30691 ( .A(n25857), .B(n25856), .Z(n25858) );
  XNOR U30692 ( .A(n25852), .B(n25853), .Z(n25856) );
  XNOR U30693 ( .A(y[201]), .B(x[201]), .Z(n25853) );
  XNOR U30694 ( .A(n25854), .B(n25855), .Z(n25852) );
  XNOR U30695 ( .A(y[202]), .B(x[202]), .Z(n25855) );
  XNOR U30696 ( .A(y[203]), .B(x[203]), .Z(n25854) );
  XNOR U30697 ( .A(n25846), .B(n25847), .Z(n25857) );
  XNOR U30698 ( .A(y[198]), .B(x[198]), .Z(n25847) );
  XNOR U30699 ( .A(n25848), .B(n25849), .Z(n25846) );
  XNOR U30700 ( .A(y[199]), .B(x[199]), .Z(n25849) );
  XNOR U30701 ( .A(y[200]), .B(x[200]), .Z(n25848) );
  NAND U30702 ( .A(n25913), .B(n25914), .Z(N28029) );
  NANDN U30703 ( .A(n25915), .B(n25916), .Z(n25914) );
  OR U30704 ( .A(n25917), .B(n25918), .Z(n25916) );
  NAND U30705 ( .A(n25917), .B(n25918), .Z(n25913) );
  XOR U30706 ( .A(n25917), .B(n25919), .Z(N28028) );
  XNOR U30707 ( .A(n25915), .B(n25918), .Z(n25919) );
  AND U30708 ( .A(n25920), .B(n25921), .Z(n25918) );
  NANDN U30709 ( .A(n25922), .B(n25923), .Z(n25921) );
  NANDN U30710 ( .A(n25924), .B(n25925), .Z(n25923) );
  NANDN U30711 ( .A(n25925), .B(n25924), .Z(n25920) );
  NAND U30712 ( .A(n25926), .B(n25927), .Z(n25915) );
  NANDN U30713 ( .A(n25928), .B(n25929), .Z(n25927) );
  OR U30714 ( .A(n25930), .B(n25931), .Z(n25929) );
  NAND U30715 ( .A(n25931), .B(n25930), .Z(n25926) );
  AND U30716 ( .A(n25932), .B(n25933), .Z(n25917) );
  NANDN U30717 ( .A(n25934), .B(n25935), .Z(n25933) );
  NANDN U30718 ( .A(n25936), .B(n25937), .Z(n25935) );
  NANDN U30719 ( .A(n25937), .B(n25936), .Z(n25932) );
  XOR U30720 ( .A(n25931), .B(n25938), .Z(N28027) );
  XOR U30721 ( .A(n25928), .B(n25930), .Z(n25938) );
  XNOR U30722 ( .A(n25924), .B(n25939), .Z(n25930) );
  XNOR U30723 ( .A(n25922), .B(n25925), .Z(n25939) );
  NAND U30724 ( .A(n25940), .B(n25941), .Z(n25925) );
  NAND U30725 ( .A(n25942), .B(n25943), .Z(n25941) );
  OR U30726 ( .A(n25944), .B(n25945), .Z(n25942) );
  NANDN U30727 ( .A(n25946), .B(n25944), .Z(n25940) );
  IV U30728 ( .A(n25945), .Z(n25946) );
  NAND U30729 ( .A(n25947), .B(n25948), .Z(n25922) );
  NAND U30730 ( .A(n25949), .B(n25950), .Z(n25948) );
  NANDN U30731 ( .A(n25951), .B(n25952), .Z(n25949) );
  NANDN U30732 ( .A(n25952), .B(n25951), .Z(n25947) );
  AND U30733 ( .A(n25953), .B(n25954), .Z(n25924) );
  NAND U30734 ( .A(n25955), .B(n25956), .Z(n25954) );
  OR U30735 ( .A(n25957), .B(n25958), .Z(n25955) );
  NANDN U30736 ( .A(n25959), .B(n25957), .Z(n25953) );
  NAND U30737 ( .A(n25960), .B(n25961), .Z(n25928) );
  NANDN U30738 ( .A(n25962), .B(n25963), .Z(n25961) );
  OR U30739 ( .A(n25964), .B(n25965), .Z(n25963) );
  NANDN U30740 ( .A(n25966), .B(n25964), .Z(n25960) );
  IV U30741 ( .A(n25965), .Z(n25966) );
  XNOR U30742 ( .A(n25936), .B(n25967), .Z(n25931) );
  XNOR U30743 ( .A(n25934), .B(n25937), .Z(n25967) );
  NAND U30744 ( .A(n25968), .B(n25969), .Z(n25937) );
  NAND U30745 ( .A(n25970), .B(n25971), .Z(n25969) );
  OR U30746 ( .A(n25972), .B(n25973), .Z(n25970) );
  NANDN U30747 ( .A(n25974), .B(n25972), .Z(n25968) );
  IV U30748 ( .A(n25973), .Z(n25974) );
  NAND U30749 ( .A(n25975), .B(n25976), .Z(n25934) );
  NAND U30750 ( .A(n25977), .B(n25978), .Z(n25976) );
  NANDN U30751 ( .A(n25979), .B(n25980), .Z(n25977) );
  NANDN U30752 ( .A(n25980), .B(n25979), .Z(n25975) );
  AND U30753 ( .A(n25981), .B(n25982), .Z(n25936) );
  NAND U30754 ( .A(n25983), .B(n25984), .Z(n25982) );
  OR U30755 ( .A(n25985), .B(n25986), .Z(n25983) );
  NANDN U30756 ( .A(n25987), .B(n25985), .Z(n25981) );
  XNOR U30757 ( .A(n25962), .B(n25988), .Z(N28026) );
  XOR U30758 ( .A(n25964), .B(n25965), .Z(n25988) );
  XNOR U30759 ( .A(n25978), .B(n25989), .Z(n25965) );
  XOR U30760 ( .A(n25979), .B(n25980), .Z(n25989) );
  XOR U30761 ( .A(n25985), .B(n25990), .Z(n25980) );
  XOR U30762 ( .A(n25984), .B(n25987), .Z(n25990) );
  IV U30763 ( .A(n25986), .Z(n25987) );
  NAND U30764 ( .A(n25991), .B(n25992), .Z(n25986) );
  OR U30765 ( .A(n25993), .B(n25994), .Z(n25992) );
  OR U30766 ( .A(n25995), .B(n25996), .Z(n25991) );
  NAND U30767 ( .A(n25997), .B(n25998), .Z(n25984) );
  OR U30768 ( .A(n25999), .B(n26000), .Z(n25998) );
  OR U30769 ( .A(n26001), .B(n26002), .Z(n25997) );
  NOR U30770 ( .A(n26003), .B(n26004), .Z(n25985) );
  ANDN U30771 ( .B(n26005), .A(n26006), .Z(n25979) );
  XNOR U30772 ( .A(n25972), .B(n26007), .Z(n25978) );
  XNOR U30773 ( .A(n25971), .B(n25973), .Z(n26007) );
  NAND U30774 ( .A(n26008), .B(n26009), .Z(n25973) );
  OR U30775 ( .A(n26010), .B(n26011), .Z(n26009) );
  OR U30776 ( .A(n26012), .B(n26013), .Z(n26008) );
  NAND U30777 ( .A(n26014), .B(n26015), .Z(n25971) );
  OR U30778 ( .A(n26016), .B(n26017), .Z(n26015) );
  OR U30779 ( .A(n26018), .B(n26019), .Z(n26014) );
  ANDN U30780 ( .B(n26020), .A(n26021), .Z(n25972) );
  IV U30781 ( .A(n26022), .Z(n26020) );
  ANDN U30782 ( .B(n26023), .A(n26024), .Z(n25964) );
  XOR U30783 ( .A(n25950), .B(n26025), .Z(n25962) );
  XOR U30784 ( .A(n25951), .B(n25952), .Z(n26025) );
  XOR U30785 ( .A(n25957), .B(n26026), .Z(n25952) );
  XOR U30786 ( .A(n25956), .B(n25959), .Z(n26026) );
  IV U30787 ( .A(n25958), .Z(n25959) );
  NAND U30788 ( .A(n26027), .B(n26028), .Z(n25958) );
  OR U30789 ( .A(n26029), .B(n26030), .Z(n26028) );
  OR U30790 ( .A(n26031), .B(n26032), .Z(n26027) );
  NAND U30791 ( .A(n26033), .B(n26034), .Z(n25956) );
  OR U30792 ( .A(n26035), .B(n26036), .Z(n26034) );
  OR U30793 ( .A(n26037), .B(n26038), .Z(n26033) );
  NOR U30794 ( .A(n26039), .B(n26040), .Z(n25957) );
  ANDN U30795 ( .B(n26041), .A(n26042), .Z(n25951) );
  IV U30796 ( .A(n26043), .Z(n26041) );
  XNOR U30797 ( .A(n25944), .B(n26044), .Z(n25950) );
  XNOR U30798 ( .A(n25943), .B(n25945), .Z(n26044) );
  NAND U30799 ( .A(n26045), .B(n26046), .Z(n25945) );
  OR U30800 ( .A(n26047), .B(n26048), .Z(n26046) );
  OR U30801 ( .A(n26049), .B(n26050), .Z(n26045) );
  NAND U30802 ( .A(n26051), .B(n26052), .Z(n25943) );
  OR U30803 ( .A(n26053), .B(n26054), .Z(n26052) );
  OR U30804 ( .A(n26055), .B(n26056), .Z(n26051) );
  ANDN U30805 ( .B(n26057), .A(n26058), .Z(n25944) );
  IV U30806 ( .A(n26059), .Z(n26057) );
  XNOR U30807 ( .A(n26024), .B(n26023), .Z(N28025) );
  XOR U30808 ( .A(n26043), .B(n26042), .Z(n26023) );
  XNOR U30809 ( .A(n26058), .B(n26059), .Z(n26042) );
  XNOR U30810 ( .A(n26053), .B(n26054), .Z(n26059) );
  XNOR U30811 ( .A(n26055), .B(n26056), .Z(n26054) );
  XNOR U30812 ( .A(y[196]), .B(x[196]), .Z(n26056) );
  XNOR U30813 ( .A(y[197]), .B(x[197]), .Z(n26055) );
  XNOR U30814 ( .A(y[195]), .B(x[195]), .Z(n26053) );
  XNOR U30815 ( .A(n26047), .B(n26048), .Z(n26058) );
  XNOR U30816 ( .A(y[192]), .B(x[192]), .Z(n26048) );
  XNOR U30817 ( .A(n26049), .B(n26050), .Z(n26047) );
  XNOR U30818 ( .A(y[193]), .B(x[193]), .Z(n26050) );
  XNOR U30819 ( .A(y[194]), .B(x[194]), .Z(n26049) );
  XNOR U30820 ( .A(n26040), .B(n26039), .Z(n26043) );
  XNOR U30821 ( .A(n26035), .B(n26036), .Z(n26039) );
  XNOR U30822 ( .A(y[189]), .B(x[189]), .Z(n26036) );
  XNOR U30823 ( .A(n26037), .B(n26038), .Z(n26035) );
  XNOR U30824 ( .A(y[190]), .B(x[190]), .Z(n26038) );
  XNOR U30825 ( .A(y[191]), .B(x[191]), .Z(n26037) );
  XNOR U30826 ( .A(n26029), .B(n26030), .Z(n26040) );
  XNOR U30827 ( .A(y[186]), .B(x[186]), .Z(n26030) );
  XNOR U30828 ( .A(n26031), .B(n26032), .Z(n26029) );
  XNOR U30829 ( .A(y[187]), .B(x[187]), .Z(n26032) );
  XNOR U30830 ( .A(y[188]), .B(x[188]), .Z(n26031) );
  XOR U30831 ( .A(n26005), .B(n26006), .Z(n26024) );
  XNOR U30832 ( .A(n26021), .B(n26022), .Z(n26006) );
  XNOR U30833 ( .A(n26016), .B(n26017), .Z(n26022) );
  XNOR U30834 ( .A(n26018), .B(n26019), .Z(n26017) );
  XNOR U30835 ( .A(y[184]), .B(x[184]), .Z(n26019) );
  XNOR U30836 ( .A(y[185]), .B(x[185]), .Z(n26018) );
  XNOR U30837 ( .A(y[183]), .B(x[183]), .Z(n26016) );
  XNOR U30838 ( .A(n26010), .B(n26011), .Z(n26021) );
  XNOR U30839 ( .A(y[180]), .B(x[180]), .Z(n26011) );
  XNOR U30840 ( .A(n26012), .B(n26013), .Z(n26010) );
  XNOR U30841 ( .A(y[181]), .B(x[181]), .Z(n26013) );
  XNOR U30842 ( .A(y[182]), .B(x[182]), .Z(n26012) );
  XOR U30843 ( .A(n26004), .B(n26003), .Z(n26005) );
  XNOR U30844 ( .A(n25999), .B(n26000), .Z(n26003) );
  XNOR U30845 ( .A(y[177]), .B(x[177]), .Z(n26000) );
  XNOR U30846 ( .A(n26001), .B(n26002), .Z(n25999) );
  XNOR U30847 ( .A(y[178]), .B(x[178]), .Z(n26002) );
  XNOR U30848 ( .A(y[179]), .B(x[179]), .Z(n26001) );
  XNOR U30849 ( .A(n25993), .B(n25994), .Z(n26004) );
  XNOR U30850 ( .A(y[174]), .B(x[174]), .Z(n25994) );
  XNOR U30851 ( .A(n25995), .B(n25996), .Z(n25993) );
  XNOR U30852 ( .A(y[175]), .B(x[175]), .Z(n25996) );
  XNOR U30853 ( .A(y[176]), .B(x[176]), .Z(n25995) );
  NAND U30854 ( .A(n26060), .B(n26061), .Z(N28017) );
  NANDN U30855 ( .A(n26062), .B(n26063), .Z(n26061) );
  OR U30856 ( .A(n26064), .B(n26065), .Z(n26063) );
  NAND U30857 ( .A(n26064), .B(n26065), .Z(n26060) );
  XOR U30858 ( .A(n26064), .B(n26066), .Z(N28016) );
  XNOR U30859 ( .A(n26062), .B(n26065), .Z(n26066) );
  AND U30860 ( .A(n26067), .B(n26068), .Z(n26065) );
  NANDN U30861 ( .A(n26069), .B(n26070), .Z(n26068) );
  NANDN U30862 ( .A(n26071), .B(n26072), .Z(n26070) );
  NANDN U30863 ( .A(n26072), .B(n26071), .Z(n26067) );
  NAND U30864 ( .A(n26073), .B(n26074), .Z(n26062) );
  NANDN U30865 ( .A(n26075), .B(n26076), .Z(n26074) );
  OR U30866 ( .A(n26077), .B(n26078), .Z(n26076) );
  NAND U30867 ( .A(n26078), .B(n26077), .Z(n26073) );
  AND U30868 ( .A(n26079), .B(n26080), .Z(n26064) );
  NANDN U30869 ( .A(n26081), .B(n26082), .Z(n26080) );
  NANDN U30870 ( .A(n26083), .B(n26084), .Z(n26082) );
  NANDN U30871 ( .A(n26084), .B(n26083), .Z(n26079) );
  XOR U30872 ( .A(n26078), .B(n26085), .Z(N28015) );
  XOR U30873 ( .A(n26075), .B(n26077), .Z(n26085) );
  XNOR U30874 ( .A(n26071), .B(n26086), .Z(n26077) );
  XNOR U30875 ( .A(n26069), .B(n26072), .Z(n26086) );
  NAND U30876 ( .A(n26087), .B(n26088), .Z(n26072) );
  NAND U30877 ( .A(n26089), .B(n26090), .Z(n26088) );
  OR U30878 ( .A(n26091), .B(n26092), .Z(n26089) );
  NANDN U30879 ( .A(n26093), .B(n26091), .Z(n26087) );
  IV U30880 ( .A(n26092), .Z(n26093) );
  NAND U30881 ( .A(n26094), .B(n26095), .Z(n26069) );
  NAND U30882 ( .A(n26096), .B(n26097), .Z(n26095) );
  NANDN U30883 ( .A(n26098), .B(n26099), .Z(n26096) );
  NANDN U30884 ( .A(n26099), .B(n26098), .Z(n26094) );
  AND U30885 ( .A(n26100), .B(n26101), .Z(n26071) );
  NAND U30886 ( .A(n26102), .B(n26103), .Z(n26101) );
  OR U30887 ( .A(n26104), .B(n26105), .Z(n26102) );
  NANDN U30888 ( .A(n26106), .B(n26104), .Z(n26100) );
  NAND U30889 ( .A(n26107), .B(n26108), .Z(n26075) );
  NANDN U30890 ( .A(n26109), .B(n26110), .Z(n26108) );
  OR U30891 ( .A(n26111), .B(n26112), .Z(n26110) );
  NANDN U30892 ( .A(n26113), .B(n26111), .Z(n26107) );
  IV U30893 ( .A(n26112), .Z(n26113) );
  XNOR U30894 ( .A(n26083), .B(n26114), .Z(n26078) );
  XNOR U30895 ( .A(n26081), .B(n26084), .Z(n26114) );
  NAND U30896 ( .A(n26115), .B(n26116), .Z(n26084) );
  NAND U30897 ( .A(n26117), .B(n26118), .Z(n26116) );
  OR U30898 ( .A(n26119), .B(n26120), .Z(n26117) );
  NANDN U30899 ( .A(n26121), .B(n26119), .Z(n26115) );
  IV U30900 ( .A(n26120), .Z(n26121) );
  NAND U30901 ( .A(n26122), .B(n26123), .Z(n26081) );
  NAND U30902 ( .A(n26124), .B(n26125), .Z(n26123) );
  NANDN U30903 ( .A(n26126), .B(n26127), .Z(n26124) );
  NANDN U30904 ( .A(n26127), .B(n26126), .Z(n26122) );
  AND U30905 ( .A(n26128), .B(n26129), .Z(n26083) );
  NAND U30906 ( .A(n26130), .B(n26131), .Z(n26129) );
  OR U30907 ( .A(n26132), .B(n26133), .Z(n26130) );
  NANDN U30908 ( .A(n26134), .B(n26132), .Z(n26128) );
  XNOR U30909 ( .A(n26109), .B(n26135), .Z(N28014) );
  XOR U30910 ( .A(n26111), .B(n26112), .Z(n26135) );
  XNOR U30911 ( .A(n26125), .B(n26136), .Z(n26112) );
  XOR U30912 ( .A(n26126), .B(n26127), .Z(n26136) );
  XOR U30913 ( .A(n26132), .B(n26137), .Z(n26127) );
  XOR U30914 ( .A(n26131), .B(n26134), .Z(n26137) );
  IV U30915 ( .A(n26133), .Z(n26134) );
  NAND U30916 ( .A(n26138), .B(n26139), .Z(n26133) );
  OR U30917 ( .A(n26140), .B(n26141), .Z(n26139) );
  OR U30918 ( .A(n26142), .B(n26143), .Z(n26138) );
  NAND U30919 ( .A(n26144), .B(n26145), .Z(n26131) );
  OR U30920 ( .A(n26146), .B(n26147), .Z(n26145) );
  OR U30921 ( .A(n26148), .B(n26149), .Z(n26144) );
  NOR U30922 ( .A(n26150), .B(n26151), .Z(n26132) );
  ANDN U30923 ( .B(n26152), .A(n26153), .Z(n26126) );
  XNOR U30924 ( .A(n26119), .B(n26154), .Z(n26125) );
  XNOR U30925 ( .A(n26118), .B(n26120), .Z(n26154) );
  NAND U30926 ( .A(n26155), .B(n26156), .Z(n26120) );
  OR U30927 ( .A(n26157), .B(n26158), .Z(n26156) );
  OR U30928 ( .A(n26159), .B(n26160), .Z(n26155) );
  NAND U30929 ( .A(n26161), .B(n26162), .Z(n26118) );
  OR U30930 ( .A(n26163), .B(n26164), .Z(n26162) );
  OR U30931 ( .A(n26165), .B(n26166), .Z(n26161) );
  ANDN U30932 ( .B(n26167), .A(n26168), .Z(n26119) );
  IV U30933 ( .A(n26169), .Z(n26167) );
  ANDN U30934 ( .B(n26170), .A(n26171), .Z(n26111) );
  XOR U30935 ( .A(n26097), .B(n26172), .Z(n26109) );
  XOR U30936 ( .A(n26098), .B(n26099), .Z(n26172) );
  XOR U30937 ( .A(n26104), .B(n26173), .Z(n26099) );
  XOR U30938 ( .A(n26103), .B(n26106), .Z(n26173) );
  IV U30939 ( .A(n26105), .Z(n26106) );
  NAND U30940 ( .A(n26174), .B(n26175), .Z(n26105) );
  OR U30941 ( .A(n26176), .B(n26177), .Z(n26175) );
  OR U30942 ( .A(n26178), .B(n26179), .Z(n26174) );
  NAND U30943 ( .A(n26180), .B(n26181), .Z(n26103) );
  OR U30944 ( .A(n26182), .B(n26183), .Z(n26181) );
  OR U30945 ( .A(n26184), .B(n26185), .Z(n26180) );
  NOR U30946 ( .A(n26186), .B(n26187), .Z(n26104) );
  ANDN U30947 ( .B(n26188), .A(n26189), .Z(n26098) );
  IV U30948 ( .A(n26190), .Z(n26188) );
  XNOR U30949 ( .A(n26091), .B(n26191), .Z(n26097) );
  XNOR U30950 ( .A(n26090), .B(n26092), .Z(n26191) );
  NAND U30951 ( .A(n26192), .B(n26193), .Z(n26092) );
  OR U30952 ( .A(n26194), .B(n26195), .Z(n26193) );
  OR U30953 ( .A(n26196), .B(n26197), .Z(n26192) );
  NAND U30954 ( .A(n26198), .B(n26199), .Z(n26090) );
  OR U30955 ( .A(n26200), .B(n26201), .Z(n26199) );
  OR U30956 ( .A(n26202), .B(n26203), .Z(n26198) );
  ANDN U30957 ( .B(n26204), .A(n26205), .Z(n26091) );
  IV U30958 ( .A(n26206), .Z(n26204) );
  XNOR U30959 ( .A(n26171), .B(n26170), .Z(N28013) );
  XOR U30960 ( .A(n26190), .B(n26189), .Z(n26170) );
  XNOR U30961 ( .A(n26205), .B(n26206), .Z(n26189) );
  XNOR U30962 ( .A(n26200), .B(n26201), .Z(n26206) );
  XNOR U30963 ( .A(n26202), .B(n26203), .Z(n26201) );
  XNOR U30964 ( .A(y[172]), .B(x[172]), .Z(n26203) );
  XNOR U30965 ( .A(y[173]), .B(x[173]), .Z(n26202) );
  XNOR U30966 ( .A(y[171]), .B(x[171]), .Z(n26200) );
  XNOR U30967 ( .A(n26194), .B(n26195), .Z(n26205) );
  XNOR U30968 ( .A(y[168]), .B(x[168]), .Z(n26195) );
  XNOR U30969 ( .A(n26196), .B(n26197), .Z(n26194) );
  XNOR U30970 ( .A(y[169]), .B(x[169]), .Z(n26197) );
  XNOR U30971 ( .A(y[170]), .B(x[170]), .Z(n26196) );
  XNOR U30972 ( .A(n26187), .B(n26186), .Z(n26190) );
  XNOR U30973 ( .A(n26182), .B(n26183), .Z(n26186) );
  XNOR U30974 ( .A(y[165]), .B(x[165]), .Z(n26183) );
  XNOR U30975 ( .A(n26184), .B(n26185), .Z(n26182) );
  XNOR U30976 ( .A(y[166]), .B(x[166]), .Z(n26185) );
  XNOR U30977 ( .A(y[167]), .B(x[167]), .Z(n26184) );
  XNOR U30978 ( .A(n26176), .B(n26177), .Z(n26187) );
  XNOR U30979 ( .A(y[162]), .B(x[162]), .Z(n26177) );
  XNOR U30980 ( .A(n26178), .B(n26179), .Z(n26176) );
  XNOR U30981 ( .A(y[163]), .B(x[163]), .Z(n26179) );
  XNOR U30982 ( .A(y[164]), .B(x[164]), .Z(n26178) );
  XOR U30983 ( .A(n26152), .B(n26153), .Z(n26171) );
  XNOR U30984 ( .A(n26168), .B(n26169), .Z(n26153) );
  XNOR U30985 ( .A(n26163), .B(n26164), .Z(n26169) );
  XNOR U30986 ( .A(n26165), .B(n26166), .Z(n26164) );
  XNOR U30987 ( .A(y[160]), .B(x[160]), .Z(n26166) );
  XNOR U30988 ( .A(y[161]), .B(x[161]), .Z(n26165) );
  XNOR U30989 ( .A(y[159]), .B(x[159]), .Z(n26163) );
  XNOR U30990 ( .A(n26157), .B(n26158), .Z(n26168) );
  XNOR U30991 ( .A(y[156]), .B(x[156]), .Z(n26158) );
  XNOR U30992 ( .A(n26159), .B(n26160), .Z(n26157) );
  XNOR U30993 ( .A(y[157]), .B(x[157]), .Z(n26160) );
  XNOR U30994 ( .A(y[158]), .B(x[158]), .Z(n26159) );
  XOR U30995 ( .A(n26151), .B(n26150), .Z(n26152) );
  XNOR U30996 ( .A(n26146), .B(n26147), .Z(n26150) );
  XNOR U30997 ( .A(y[153]), .B(x[153]), .Z(n26147) );
  XNOR U30998 ( .A(n26148), .B(n26149), .Z(n26146) );
  XNOR U30999 ( .A(y[154]), .B(x[154]), .Z(n26149) );
  XNOR U31000 ( .A(y[155]), .B(x[155]), .Z(n26148) );
  XNOR U31001 ( .A(n26140), .B(n26141), .Z(n26151) );
  XNOR U31002 ( .A(y[150]), .B(x[150]), .Z(n26141) );
  XNOR U31003 ( .A(n26142), .B(n26143), .Z(n26140) );
  XNOR U31004 ( .A(y[151]), .B(x[151]), .Z(n26143) );
  XNOR U31005 ( .A(y[152]), .B(x[152]), .Z(n26142) );
  NAND U31006 ( .A(n26207), .B(n26208), .Z(N28005) );
  NANDN U31007 ( .A(n26209), .B(n26210), .Z(n26208) );
  OR U31008 ( .A(n26211), .B(n26212), .Z(n26210) );
  NAND U31009 ( .A(n26211), .B(n26212), .Z(n26207) );
  XOR U31010 ( .A(n26211), .B(n26213), .Z(N28004) );
  XNOR U31011 ( .A(n26209), .B(n26212), .Z(n26213) );
  AND U31012 ( .A(n26214), .B(n26215), .Z(n26212) );
  NANDN U31013 ( .A(n26216), .B(n26217), .Z(n26215) );
  NANDN U31014 ( .A(n26218), .B(n26219), .Z(n26217) );
  NANDN U31015 ( .A(n26219), .B(n26218), .Z(n26214) );
  NAND U31016 ( .A(n26220), .B(n26221), .Z(n26209) );
  NANDN U31017 ( .A(n26222), .B(n26223), .Z(n26221) );
  OR U31018 ( .A(n26224), .B(n26225), .Z(n26223) );
  NAND U31019 ( .A(n26225), .B(n26224), .Z(n26220) );
  AND U31020 ( .A(n26226), .B(n26227), .Z(n26211) );
  NANDN U31021 ( .A(n26228), .B(n26229), .Z(n26227) );
  NANDN U31022 ( .A(n26230), .B(n26231), .Z(n26229) );
  NANDN U31023 ( .A(n26231), .B(n26230), .Z(n26226) );
  XOR U31024 ( .A(n26225), .B(n26232), .Z(N28003) );
  XOR U31025 ( .A(n26222), .B(n26224), .Z(n26232) );
  XNOR U31026 ( .A(n26218), .B(n26233), .Z(n26224) );
  XNOR U31027 ( .A(n26216), .B(n26219), .Z(n26233) );
  NAND U31028 ( .A(n26234), .B(n26235), .Z(n26219) );
  NAND U31029 ( .A(n26236), .B(n26237), .Z(n26235) );
  OR U31030 ( .A(n26238), .B(n26239), .Z(n26236) );
  NANDN U31031 ( .A(n26240), .B(n26238), .Z(n26234) );
  IV U31032 ( .A(n26239), .Z(n26240) );
  NAND U31033 ( .A(n26241), .B(n26242), .Z(n26216) );
  NAND U31034 ( .A(n26243), .B(n26244), .Z(n26242) );
  NANDN U31035 ( .A(n26245), .B(n26246), .Z(n26243) );
  NANDN U31036 ( .A(n26246), .B(n26245), .Z(n26241) );
  AND U31037 ( .A(n26247), .B(n26248), .Z(n26218) );
  NAND U31038 ( .A(n26249), .B(n26250), .Z(n26248) );
  OR U31039 ( .A(n26251), .B(n26252), .Z(n26249) );
  NANDN U31040 ( .A(n26253), .B(n26251), .Z(n26247) );
  NAND U31041 ( .A(n26254), .B(n26255), .Z(n26222) );
  NANDN U31042 ( .A(n26256), .B(n26257), .Z(n26255) );
  OR U31043 ( .A(n26258), .B(n26259), .Z(n26257) );
  NANDN U31044 ( .A(n26260), .B(n26258), .Z(n26254) );
  IV U31045 ( .A(n26259), .Z(n26260) );
  XNOR U31046 ( .A(n26230), .B(n26261), .Z(n26225) );
  XNOR U31047 ( .A(n26228), .B(n26231), .Z(n26261) );
  NAND U31048 ( .A(n26262), .B(n26263), .Z(n26231) );
  NAND U31049 ( .A(n26264), .B(n26265), .Z(n26263) );
  OR U31050 ( .A(n26266), .B(n26267), .Z(n26264) );
  NANDN U31051 ( .A(n26268), .B(n26266), .Z(n26262) );
  IV U31052 ( .A(n26267), .Z(n26268) );
  NAND U31053 ( .A(n26269), .B(n26270), .Z(n26228) );
  NAND U31054 ( .A(n26271), .B(n26272), .Z(n26270) );
  NANDN U31055 ( .A(n26273), .B(n26274), .Z(n26271) );
  NANDN U31056 ( .A(n26274), .B(n26273), .Z(n26269) );
  AND U31057 ( .A(n26275), .B(n26276), .Z(n26230) );
  NAND U31058 ( .A(n26277), .B(n26278), .Z(n26276) );
  OR U31059 ( .A(n26279), .B(n26280), .Z(n26277) );
  NANDN U31060 ( .A(n26281), .B(n26279), .Z(n26275) );
  XNOR U31061 ( .A(n26256), .B(n26282), .Z(N28002) );
  XOR U31062 ( .A(n26258), .B(n26259), .Z(n26282) );
  XNOR U31063 ( .A(n26272), .B(n26283), .Z(n26259) );
  XOR U31064 ( .A(n26273), .B(n26274), .Z(n26283) );
  XOR U31065 ( .A(n26279), .B(n26284), .Z(n26274) );
  XOR U31066 ( .A(n26278), .B(n26281), .Z(n26284) );
  IV U31067 ( .A(n26280), .Z(n26281) );
  NAND U31068 ( .A(n26285), .B(n26286), .Z(n26280) );
  OR U31069 ( .A(n26287), .B(n26288), .Z(n26286) );
  OR U31070 ( .A(n26289), .B(n26290), .Z(n26285) );
  NAND U31071 ( .A(n26291), .B(n26292), .Z(n26278) );
  OR U31072 ( .A(n26293), .B(n26294), .Z(n26292) );
  OR U31073 ( .A(n26295), .B(n26296), .Z(n26291) );
  NOR U31074 ( .A(n26297), .B(n26298), .Z(n26279) );
  ANDN U31075 ( .B(n26299), .A(n26300), .Z(n26273) );
  XNOR U31076 ( .A(n26266), .B(n26301), .Z(n26272) );
  XNOR U31077 ( .A(n26265), .B(n26267), .Z(n26301) );
  NAND U31078 ( .A(n26302), .B(n26303), .Z(n26267) );
  OR U31079 ( .A(n26304), .B(n26305), .Z(n26303) );
  OR U31080 ( .A(n26306), .B(n26307), .Z(n26302) );
  NAND U31081 ( .A(n26308), .B(n26309), .Z(n26265) );
  OR U31082 ( .A(n26310), .B(n26311), .Z(n26309) );
  OR U31083 ( .A(n26312), .B(n26313), .Z(n26308) );
  ANDN U31084 ( .B(n26314), .A(n26315), .Z(n26266) );
  IV U31085 ( .A(n26316), .Z(n26314) );
  ANDN U31086 ( .B(n26317), .A(n26318), .Z(n26258) );
  XOR U31087 ( .A(n26244), .B(n26319), .Z(n26256) );
  XOR U31088 ( .A(n26245), .B(n26246), .Z(n26319) );
  XOR U31089 ( .A(n26251), .B(n26320), .Z(n26246) );
  XOR U31090 ( .A(n26250), .B(n26253), .Z(n26320) );
  IV U31091 ( .A(n26252), .Z(n26253) );
  NAND U31092 ( .A(n26321), .B(n26322), .Z(n26252) );
  OR U31093 ( .A(n26323), .B(n26324), .Z(n26322) );
  OR U31094 ( .A(n26325), .B(n26326), .Z(n26321) );
  NAND U31095 ( .A(n26327), .B(n26328), .Z(n26250) );
  OR U31096 ( .A(n26329), .B(n26330), .Z(n26328) );
  OR U31097 ( .A(n26331), .B(n26332), .Z(n26327) );
  NOR U31098 ( .A(n26333), .B(n26334), .Z(n26251) );
  ANDN U31099 ( .B(n26335), .A(n26336), .Z(n26245) );
  IV U31100 ( .A(n26337), .Z(n26335) );
  XNOR U31101 ( .A(n26238), .B(n26338), .Z(n26244) );
  XNOR U31102 ( .A(n26237), .B(n26239), .Z(n26338) );
  NAND U31103 ( .A(n26339), .B(n26340), .Z(n26239) );
  OR U31104 ( .A(n26341), .B(n26342), .Z(n26340) );
  OR U31105 ( .A(n26343), .B(n26344), .Z(n26339) );
  NAND U31106 ( .A(n26345), .B(n26346), .Z(n26237) );
  OR U31107 ( .A(n26347), .B(n26348), .Z(n26346) );
  OR U31108 ( .A(n26349), .B(n26350), .Z(n26345) );
  ANDN U31109 ( .B(n26351), .A(n26352), .Z(n26238) );
  IV U31110 ( .A(n26353), .Z(n26351) );
  XNOR U31111 ( .A(n26318), .B(n26317), .Z(N28001) );
  XOR U31112 ( .A(n26337), .B(n26336), .Z(n26317) );
  XNOR U31113 ( .A(n26352), .B(n26353), .Z(n26336) );
  XNOR U31114 ( .A(n26347), .B(n26348), .Z(n26353) );
  XNOR U31115 ( .A(n26349), .B(n26350), .Z(n26348) );
  XNOR U31116 ( .A(y[148]), .B(x[148]), .Z(n26350) );
  XNOR U31117 ( .A(y[149]), .B(x[149]), .Z(n26349) );
  XNOR U31118 ( .A(y[147]), .B(x[147]), .Z(n26347) );
  XNOR U31119 ( .A(n26341), .B(n26342), .Z(n26352) );
  XNOR U31120 ( .A(y[144]), .B(x[144]), .Z(n26342) );
  XNOR U31121 ( .A(n26343), .B(n26344), .Z(n26341) );
  XNOR U31122 ( .A(y[145]), .B(x[145]), .Z(n26344) );
  XNOR U31123 ( .A(y[146]), .B(x[146]), .Z(n26343) );
  XNOR U31124 ( .A(n26334), .B(n26333), .Z(n26337) );
  XNOR U31125 ( .A(n26329), .B(n26330), .Z(n26333) );
  XNOR U31126 ( .A(y[141]), .B(x[141]), .Z(n26330) );
  XNOR U31127 ( .A(n26331), .B(n26332), .Z(n26329) );
  XNOR U31128 ( .A(y[142]), .B(x[142]), .Z(n26332) );
  XNOR U31129 ( .A(y[143]), .B(x[143]), .Z(n26331) );
  XNOR U31130 ( .A(n26323), .B(n26324), .Z(n26334) );
  XNOR U31131 ( .A(y[138]), .B(x[138]), .Z(n26324) );
  XNOR U31132 ( .A(n26325), .B(n26326), .Z(n26323) );
  XNOR U31133 ( .A(y[139]), .B(x[139]), .Z(n26326) );
  XNOR U31134 ( .A(y[140]), .B(x[140]), .Z(n26325) );
  XOR U31135 ( .A(n26299), .B(n26300), .Z(n26318) );
  XNOR U31136 ( .A(n26315), .B(n26316), .Z(n26300) );
  XNOR U31137 ( .A(n26310), .B(n26311), .Z(n26316) );
  XNOR U31138 ( .A(n26312), .B(n26313), .Z(n26311) );
  XNOR U31139 ( .A(y[136]), .B(x[136]), .Z(n26313) );
  XNOR U31140 ( .A(y[137]), .B(x[137]), .Z(n26312) );
  XNOR U31141 ( .A(y[135]), .B(x[135]), .Z(n26310) );
  XNOR U31142 ( .A(n26304), .B(n26305), .Z(n26315) );
  XNOR U31143 ( .A(y[132]), .B(x[132]), .Z(n26305) );
  XNOR U31144 ( .A(n26306), .B(n26307), .Z(n26304) );
  XNOR U31145 ( .A(y[133]), .B(x[133]), .Z(n26307) );
  XNOR U31146 ( .A(y[134]), .B(x[134]), .Z(n26306) );
  XOR U31147 ( .A(n26298), .B(n26297), .Z(n26299) );
  XNOR U31148 ( .A(n26293), .B(n26294), .Z(n26297) );
  XNOR U31149 ( .A(y[129]), .B(x[129]), .Z(n26294) );
  XNOR U31150 ( .A(n26295), .B(n26296), .Z(n26293) );
  XNOR U31151 ( .A(y[130]), .B(x[130]), .Z(n26296) );
  XNOR U31152 ( .A(y[131]), .B(x[131]), .Z(n26295) );
  XNOR U31153 ( .A(n26287), .B(n26288), .Z(n26298) );
  XNOR U31154 ( .A(y[126]), .B(x[126]), .Z(n26288) );
  XNOR U31155 ( .A(n26289), .B(n26290), .Z(n26287) );
  XNOR U31156 ( .A(y[127]), .B(x[127]), .Z(n26290) );
  XNOR U31157 ( .A(y[128]), .B(x[128]), .Z(n26289) );
  NAND U31158 ( .A(n26354), .B(n26355), .Z(N27993) );
  NANDN U31159 ( .A(n26356), .B(n26357), .Z(n26355) );
  OR U31160 ( .A(n26358), .B(n26359), .Z(n26357) );
  NAND U31161 ( .A(n26358), .B(n26359), .Z(n26354) );
  XOR U31162 ( .A(n26358), .B(n26360), .Z(N27992) );
  XNOR U31163 ( .A(n26356), .B(n26359), .Z(n26360) );
  AND U31164 ( .A(n26361), .B(n26362), .Z(n26359) );
  NANDN U31165 ( .A(n26363), .B(n26364), .Z(n26362) );
  NANDN U31166 ( .A(n26365), .B(n26366), .Z(n26364) );
  NANDN U31167 ( .A(n26366), .B(n26365), .Z(n26361) );
  NAND U31168 ( .A(n26367), .B(n26368), .Z(n26356) );
  NANDN U31169 ( .A(n26369), .B(n26370), .Z(n26368) );
  OR U31170 ( .A(n26371), .B(n26372), .Z(n26370) );
  NAND U31171 ( .A(n26372), .B(n26371), .Z(n26367) );
  AND U31172 ( .A(n26373), .B(n26374), .Z(n26358) );
  NANDN U31173 ( .A(n26375), .B(n26376), .Z(n26374) );
  NANDN U31174 ( .A(n26377), .B(n26378), .Z(n26376) );
  NANDN U31175 ( .A(n26378), .B(n26377), .Z(n26373) );
  XOR U31176 ( .A(n26372), .B(n26379), .Z(N27991) );
  XOR U31177 ( .A(n26369), .B(n26371), .Z(n26379) );
  XNOR U31178 ( .A(n26365), .B(n26380), .Z(n26371) );
  XNOR U31179 ( .A(n26363), .B(n26366), .Z(n26380) );
  NAND U31180 ( .A(n26381), .B(n26382), .Z(n26366) );
  NAND U31181 ( .A(n26383), .B(n26384), .Z(n26382) );
  OR U31182 ( .A(n26385), .B(n26386), .Z(n26383) );
  NANDN U31183 ( .A(n26387), .B(n26385), .Z(n26381) );
  IV U31184 ( .A(n26386), .Z(n26387) );
  NAND U31185 ( .A(n26388), .B(n26389), .Z(n26363) );
  NAND U31186 ( .A(n26390), .B(n26391), .Z(n26389) );
  NANDN U31187 ( .A(n26392), .B(n26393), .Z(n26390) );
  NANDN U31188 ( .A(n26393), .B(n26392), .Z(n26388) );
  AND U31189 ( .A(n26394), .B(n26395), .Z(n26365) );
  NAND U31190 ( .A(n26396), .B(n26397), .Z(n26395) );
  OR U31191 ( .A(n26398), .B(n26399), .Z(n26396) );
  NANDN U31192 ( .A(n26400), .B(n26398), .Z(n26394) );
  NAND U31193 ( .A(n26401), .B(n26402), .Z(n26369) );
  NANDN U31194 ( .A(n26403), .B(n26404), .Z(n26402) );
  OR U31195 ( .A(n26405), .B(n26406), .Z(n26404) );
  NANDN U31196 ( .A(n26407), .B(n26405), .Z(n26401) );
  IV U31197 ( .A(n26406), .Z(n26407) );
  XNOR U31198 ( .A(n26377), .B(n26408), .Z(n26372) );
  XNOR U31199 ( .A(n26375), .B(n26378), .Z(n26408) );
  NAND U31200 ( .A(n26409), .B(n26410), .Z(n26378) );
  NAND U31201 ( .A(n26411), .B(n26412), .Z(n26410) );
  OR U31202 ( .A(n26413), .B(n26414), .Z(n26411) );
  NANDN U31203 ( .A(n26415), .B(n26413), .Z(n26409) );
  IV U31204 ( .A(n26414), .Z(n26415) );
  NAND U31205 ( .A(n26416), .B(n26417), .Z(n26375) );
  NAND U31206 ( .A(n26418), .B(n26419), .Z(n26417) );
  NANDN U31207 ( .A(n26420), .B(n26421), .Z(n26418) );
  NANDN U31208 ( .A(n26421), .B(n26420), .Z(n26416) );
  AND U31209 ( .A(n26422), .B(n26423), .Z(n26377) );
  NAND U31210 ( .A(n26424), .B(n26425), .Z(n26423) );
  OR U31211 ( .A(n26426), .B(n26427), .Z(n26424) );
  NANDN U31212 ( .A(n26428), .B(n26426), .Z(n26422) );
  XNOR U31213 ( .A(n26403), .B(n26429), .Z(N27990) );
  XOR U31214 ( .A(n26405), .B(n26406), .Z(n26429) );
  XNOR U31215 ( .A(n26419), .B(n26430), .Z(n26406) );
  XOR U31216 ( .A(n26420), .B(n26421), .Z(n26430) );
  XOR U31217 ( .A(n26426), .B(n26431), .Z(n26421) );
  XOR U31218 ( .A(n26425), .B(n26428), .Z(n26431) );
  IV U31219 ( .A(n26427), .Z(n26428) );
  NAND U31220 ( .A(n26432), .B(n26433), .Z(n26427) );
  OR U31221 ( .A(n26434), .B(n26435), .Z(n26433) );
  OR U31222 ( .A(n26436), .B(n26437), .Z(n26432) );
  NAND U31223 ( .A(n26438), .B(n26439), .Z(n26425) );
  OR U31224 ( .A(n26440), .B(n26441), .Z(n26439) );
  OR U31225 ( .A(n26442), .B(n26443), .Z(n26438) );
  NOR U31226 ( .A(n26444), .B(n26445), .Z(n26426) );
  ANDN U31227 ( .B(n26446), .A(n26447), .Z(n26420) );
  XNOR U31228 ( .A(n26413), .B(n26448), .Z(n26419) );
  XNOR U31229 ( .A(n26412), .B(n26414), .Z(n26448) );
  NAND U31230 ( .A(n26449), .B(n26450), .Z(n26414) );
  OR U31231 ( .A(n26451), .B(n26452), .Z(n26450) );
  OR U31232 ( .A(n26453), .B(n26454), .Z(n26449) );
  NAND U31233 ( .A(n26455), .B(n26456), .Z(n26412) );
  OR U31234 ( .A(n26457), .B(n26458), .Z(n26456) );
  OR U31235 ( .A(n26459), .B(n26460), .Z(n26455) );
  ANDN U31236 ( .B(n26461), .A(n26462), .Z(n26413) );
  IV U31237 ( .A(n26463), .Z(n26461) );
  ANDN U31238 ( .B(n26464), .A(n26465), .Z(n26405) );
  XOR U31239 ( .A(n26391), .B(n26466), .Z(n26403) );
  XOR U31240 ( .A(n26392), .B(n26393), .Z(n26466) );
  XOR U31241 ( .A(n26398), .B(n26467), .Z(n26393) );
  XOR U31242 ( .A(n26397), .B(n26400), .Z(n26467) );
  IV U31243 ( .A(n26399), .Z(n26400) );
  NAND U31244 ( .A(n26468), .B(n26469), .Z(n26399) );
  OR U31245 ( .A(n26470), .B(n26471), .Z(n26469) );
  OR U31246 ( .A(n26472), .B(n26473), .Z(n26468) );
  NAND U31247 ( .A(n26474), .B(n26475), .Z(n26397) );
  OR U31248 ( .A(n26476), .B(n26477), .Z(n26475) );
  OR U31249 ( .A(n26478), .B(n26479), .Z(n26474) );
  NOR U31250 ( .A(n26480), .B(n26481), .Z(n26398) );
  ANDN U31251 ( .B(n26482), .A(n26483), .Z(n26392) );
  IV U31252 ( .A(n26484), .Z(n26482) );
  XNOR U31253 ( .A(n26385), .B(n26485), .Z(n26391) );
  XNOR U31254 ( .A(n26384), .B(n26386), .Z(n26485) );
  NAND U31255 ( .A(n26486), .B(n26487), .Z(n26386) );
  OR U31256 ( .A(n26488), .B(n26489), .Z(n26487) );
  OR U31257 ( .A(n26490), .B(n26491), .Z(n26486) );
  NAND U31258 ( .A(n26492), .B(n26493), .Z(n26384) );
  OR U31259 ( .A(n26494), .B(n26495), .Z(n26493) );
  OR U31260 ( .A(n26496), .B(n26497), .Z(n26492) );
  ANDN U31261 ( .B(n26498), .A(n26499), .Z(n26385) );
  IV U31262 ( .A(n26500), .Z(n26498) );
  XNOR U31263 ( .A(n26465), .B(n26464), .Z(N27989) );
  XOR U31264 ( .A(n26484), .B(n26483), .Z(n26464) );
  XNOR U31265 ( .A(n26499), .B(n26500), .Z(n26483) );
  XNOR U31266 ( .A(n26494), .B(n26495), .Z(n26500) );
  XNOR U31267 ( .A(n26496), .B(n26497), .Z(n26495) );
  XNOR U31268 ( .A(y[124]), .B(x[124]), .Z(n26497) );
  XNOR U31269 ( .A(y[125]), .B(x[125]), .Z(n26496) );
  XNOR U31270 ( .A(y[123]), .B(x[123]), .Z(n26494) );
  XNOR U31271 ( .A(n26488), .B(n26489), .Z(n26499) );
  XNOR U31272 ( .A(y[120]), .B(x[120]), .Z(n26489) );
  XNOR U31273 ( .A(n26490), .B(n26491), .Z(n26488) );
  XNOR U31274 ( .A(y[121]), .B(x[121]), .Z(n26491) );
  XNOR U31275 ( .A(y[122]), .B(x[122]), .Z(n26490) );
  XNOR U31276 ( .A(n26481), .B(n26480), .Z(n26484) );
  XNOR U31277 ( .A(n26476), .B(n26477), .Z(n26480) );
  XNOR U31278 ( .A(y[117]), .B(x[117]), .Z(n26477) );
  XNOR U31279 ( .A(n26478), .B(n26479), .Z(n26476) );
  XNOR U31280 ( .A(y[118]), .B(x[118]), .Z(n26479) );
  XNOR U31281 ( .A(y[119]), .B(x[119]), .Z(n26478) );
  XNOR U31282 ( .A(n26470), .B(n26471), .Z(n26481) );
  XNOR U31283 ( .A(y[114]), .B(x[114]), .Z(n26471) );
  XNOR U31284 ( .A(n26472), .B(n26473), .Z(n26470) );
  XNOR U31285 ( .A(y[115]), .B(x[115]), .Z(n26473) );
  XNOR U31286 ( .A(y[116]), .B(x[116]), .Z(n26472) );
  XOR U31287 ( .A(n26446), .B(n26447), .Z(n26465) );
  XNOR U31288 ( .A(n26462), .B(n26463), .Z(n26447) );
  XNOR U31289 ( .A(n26457), .B(n26458), .Z(n26463) );
  XNOR U31290 ( .A(n26459), .B(n26460), .Z(n26458) );
  XNOR U31291 ( .A(y[112]), .B(x[112]), .Z(n26460) );
  XNOR U31292 ( .A(y[113]), .B(x[113]), .Z(n26459) );
  XNOR U31293 ( .A(y[111]), .B(x[111]), .Z(n26457) );
  XNOR U31294 ( .A(n26451), .B(n26452), .Z(n26462) );
  XNOR U31295 ( .A(y[108]), .B(x[108]), .Z(n26452) );
  XNOR U31296 ( .A(n26453), .B(n26454), .Z(n26451) );
  XNOR U31297 ( .A(y[109]), .B(x[109]), .Z(n26454) );
  XNOR U31298 ( .A(y[110]), .B(x[110]), .Z(n26453) );
  XOR U31299 ( .A(n26445), .B(n26444), .Z(n26446) );
  XNOR U31300 ( .A(n26440), .B(n26441), .Z(n26444) );
  XNOR U31301 ( .A(y[105]), .B(x[105]), .Z(n26441) );
  XNOR U31302 ( .A(n26442), .B(n26443), .Z(n26440) );
  XNOR U31303 ( .A(y[106]), .B(x[106]), .Z(n26443) );
  XNOR U31304 ( .A(y[107]), .B(x[107]), .Z(n26442) );
  XNOR U31305 ( .A(n26434), .B(n26435), .Z(n26445) );
  XNOR U31306 ( .A(y[102]), .B(x[102]), .Z(n26435) );
  XNOR U31307 ( .A(n26436), .B(n26437), .Z(n26434) );
  XNOR U31308 ( .A(y[103]), .B(x[103]), .Z(n26437) );
  XNOR U31309 ( .A(y[104]), .B(x[104]), .Z(n26436) );
  NAND U31310 ( .A(n26501), .B(n26502), .Z(N27981) );
  NANDN U31311 ( .A(n26503), .B(n26504), .Z(n26502) );
  OR U31312 ( .A(n26505), .B(n26506), .Z(n26504) );
  NAND U31313 ( .A(n26505), .B(n26506), .Z(n26501) );
  XOR U31314 ( .A(n26505), .B(n26507), .Z(N27980) );
  XNOR U31315 ( .A(n26503), .B(n26506), .Z(n26507) );
  AND U31316 ( .A(n26508), .B(n26509), .Z(n26506) );
  NANDN U31317 ( .A(n26510), .B(n26511), .Z(n26509) );
  NANDN U31318 ( .A(n26512), .B(n26513), .Z(n26511) );
  NANDN U31319 ( .A(n26513), .B(n26512), .Z(n26508) );
  NAND U31320 ( .A(n26514), .B(n26515), .Z(n26503) );
  NANDN U31321 ( .A(n26516), .B(n26517), .Z(n26515) );
  OR U31322 ( .A(n26518), .B(n26519), .Z(n26517) );
  NAND U31323 ( .A(n26519), .B(n26518), .Z(n26514) );
  AND U31324 ( .A(n26520), .B(n26521), .Z(n26505) );
  NANDN U31325 ( .A(n26522), .B(n26523), .Z(n26521) );
  NANDN U31326 ( .A(n26524), .B(n26525), .Z(n26523) );
  NANDN U31327 ( .A(n26525), .B(n26524), .Z(n26520) );
  XOR U31328 ( .A(n26519), .B(n26526), .Z(N27979) );
  XOR U31329 ( .A(n26516), .B(n26518), .Z(n26526) );
  XNOR U31330 ( .A(n26512), .B(n26527), .Z(n26518) );
  XNOR U31331 ( .A(n26510), .B(n26513), .Z(n26527) );
  NAND U31332 ( .A(n26528), .B(n26529), .Z(n26513) );
  NAND U31333 ( .A(n26530), .B(n26531), .Z(n26529) );
  OR U31334 ( .A(n26532), .B(n26533), .Z(n26530) );
  NANDN U31335 ( .A(n26534), .B(n26532), .Z(n26528) );
  IV U31336 ( .A(n26533), .Z(n26534) );
  NAND U31337 ( .A(n26535), .B(n26536), .Z(n26510) );
  NAND U31338 ( .A(n26537), .B(n26538), .Z(n26536) );
  NANDN U31339 ( .A(n26539), .B(n26540), .Z(n26537) );
  NANDN U31340 ( .A(n26540), .B(n26539), .Z(n26535) );
  AND U31341 ( .A(n26541), .B(n26542), .Z(n26512) );
  NAND U31342 ( .A(n26543), .B(n26544), .Z(n26542) );
  OR U31343 ( .A(n26545), .B(n26546), .Z(n26543) );
  NANDN U31344 ( .A(n26547), .B(n26545), .Z(n26541) );
  NAND U31345 ( .A(n26548), .B(n26549), .Z(n26516) );
  NANDN U31346 ( .A(n26550), .B(n26551), .Z(n26549) );
  OR U31347 ( .A(n26552), .B(n26553), .Z(n26551) );
  NANDN U31348 ( .A(n26554), .B(n26552), .Z(n26548) );
  IV U31349 ( .A(n26553), .Z(n26554) );
  XNOR U31350 ( .A(n26524), .B(n26555), .Z(n26519) );
  XNOR U31351 ( .A(n26522), .B(n26525), .Z(n26555) );
  NAND U31352 ( .A(n26556), .B(n26557), .Z(n26525) );
  NAND U31353 ( .A(n26558), .B(n26559), .Z(n26557) );
  OR U31354 ( .A(n26560), .B(n26561), .Z(n26558) );
  NANDN U31355 ( .A(n26562), .B(n26560), .Z(n26556) );
  IV U31356 ( .A(n26561), .Z(n26562) );
  NAND U31357 ( .A(n26563), .B(n26564), .Z(n26522) );
  NAND U31358 ( .A(n26565), .B(n26566), .Z(n26564) );
  NANDN U31359 ( .A(n26567), .B(n26568), .Z(n26565) );
  NANDN U31360 ( .A(n26568), .B(n26567), .Z(n26563) );
  AND U31361 ( .A(n26569), .B(n26570), .Z(n26524) );
  NAND U31362 ( .A(n26571), .B(n26572), .Z(n26570) );
  OR U31363 ( .A(n26573), .B(n26574), .Z(n26571) );
  NANDN U31364 ( .A(n26575), .B(n26573), .Z(n26569) );
  XNOR U31365 ( .A(n26550), .B(n26576), .Z(N27978) );
  XOR U31366 ( .A(n26552), .B(n26553), .Z(n26576) );
  XNOR U31367 ( .A(n26566), .B(n26577), .Z(n26553) );
  XOR U31368 ( .A(n26567), .B(n26568), .Z(n26577) );
  XOR U31369 ( .A(n26573), .B(n26578), .Z(n26568) );
  XOR U31370 ( .A(n26572), .B(n26575), .Z(n26578) );
  IV U31371 ( .A(n26574), .Z(n26575) );
  NAND U31372 ( .A(n26579), .B(n26580), .Z(n26574) );
  OR U31373 ( .A(n26581), .B(n26582), .Z(n26580) );
  OR U31374 ( .A(n26583), .B(n26584), .Z(n26579) );
  NAND U31375 ( .A(n26585), .B(n26586), .Z(n26572) );
  OR U31376 ( .A(n26587), .B(n26588), .Z(n26586) );
  OR U31377 ( .A(n26589), .B(n26590), .Z(n26585) );
  NOR U31378 ( .A(n26591), .B(n26592), .Z(n26573) );
  ANDN U31379 ( .B(n26593), .A(n26594), .Z(n26567) );
  XNOR U31380 ( .A(n26560), .B(n26595), .Z(n26566) );
  XNOR U31381 ( .A(n26559), .B(n26561), .Z(n26595) );
  NAND U31382 ( .A(n26596), .B(n26597), .Z(n26561) );
  OR U31383 ( .A(n26598), .B(n26599), .Z(n26597) );
  OR U31384 ( .A(n26600), .B(n26601), .Z(n26596) );
  NAND U31385 ( .A(n26602), .B(n26603), .Z(n26559) );
  OR U31386 ( .A(n26604), .B(n26605), .Z(n26603) );
  OR U31387 ( .A(n26606), .B(n26607), .Z(n26602) );
  ANDN U31388 ( .B(n26608), .A(n26609), .Z(n26560) );
  IV U31389 ( .A(n26610), .Z(n26608) );
  ANDN U31390 ( .B(n26611), .A(n26612), .Z(n26552) );
  XOR U31391 ( .A(n26538), .B(n26613), .Z(n26550) );
  XOR U31392 ( .A(n26539), .B(n26540), .Z(n26613) );
  XOR U31393 ( .A(n26545), .B(n26614), .Z(n26540) );
  XOR U31394 ( .A(n26544), .B(n26547), .Z(n26614) );
  IV U31395 ( .A(n26546), .Z(n26547) );
  NAND U31396 ( .A(n26615), .B(n26616), .Z(n26546) );
  OR U31397 ( .A(n26617), .B(n26618), .Z(n26616) );
  OR U31398 ( .A(n26619), .B(n26620), .Z(n26615) );
  NAND U31399 ( .A(n26621), .B(n26622), .Z(n26544) );
  OR U31400 ( .A(n26623), .B(n26624), .Z(n26622) );
  OR U31401 ( .A(n26625), .B(n26626), .Z(n26621) );
  NOR U31402 ( .A(n26627), .B(n26628), .Z(n26545) );
  ANDN U31403 ( .B(n26629), .A(n26630), .Z(n26539) );
  IV U31404 ( .A(n26631), .Z(n26629) );
  XNOR U31405 ( .A(n26532), .B(n26632), .Z(n26538) );
  XNOR U31406 ( .A(n26531), .B(n26533), .Z(n26632) );
  NAND U31407 ( .A(n26633), .B(n26634), .Z(n26533) );
  OR U31408 ( .A(n26635), .B(n26636), .Z(n26634) );
  OR U31409 ( .A(n26637), .B(n26638), .Z(n26633) );
  NAND U31410 ( .A(n26639), .B(n26640), .Z(n26531) );
  OR U31411 ( .A(n26641), .B(n26642), .Z(n26640) );
  OR U31412 ( .A(n26643), .B(n26644), .Z(n26639) );
  ANDN U31413 ( .B(n26645), .A(n26646), .Z(n26532) );
  IV U31414 ( .A(n26647), .Z(n26645) );
  XNOR U31415 ( .A(n26612), .B(n26611), .Z(N27977) );
  XOR U31416 ( .A(n26631), .B(n26630), .Z(n26611) );
  XNOR U31417 ( .A(n26646), .B(n26647), .Z(n26630) );
  XNOR U31418 ( .A(n26641), .B(n26642), .Z(n26647) );
  XNOR U31419 ( .A(n26643), .B(n26644), .Z(n26642) );
  XNOR U31420 ( .A(y[100]), .B(x[100]), .Z(n26644) );
  XNOR U31421 ( .A(y[101]), .B(x[101]), .Z(n26643) );
  XNOR U31422 ( .A(y[99]), .B(x[99]), .Z(n26641) );
  XNOR U31423 ( .A(n26635), .B(n26636), .Z(n26646) );
  XNOR U31424 ( .A(y[96]), .B(x[96]), .Z(n26636) );
  XNOR U31425 ( .A(n26637), .B(n26638), .Z(n26635) );
  XNOR U31426 ( .A(y[97]), .B(x[97]), .Z(n26638) );
  XNOR U31427 ( .A(y[98]), .B(x[98]), .Z(n26637) );
  XNOR U31428 ( .A(n26628), .B(n26627), .Z(n26631) );
  XNOR U31429 ( .A(n26623), .B(n26624), .Z(n26627) );
  XNOR U31430 ( .A(y[93]), .B(x[93]), .Z(n26624) );
  XNOR U31431 ( .A(n26625), .B(n26626), .Z(n26623) );
  XNOR U31432 ( .A(y[94]), .B(x[94]), .Z(n26626) );
  XNOR U31433 ( .A(y[95]), .B(x[95]), .Z(n26625) );
  XNOR U31434 ( .A(n26617), .B(n26618), .Z(n26628) );
  XNOR U31435 ( .A(y[90]), .B(x[90]), .Z(n26618) );
  XNOR U31436 ( .A(n26619), .B(n26620), .Z(n26617) );
  XNOR U31437 ( .A(y[91]), .B(x[91]), .Z(n26620) );
  XNOR U31438 ( .A(y[92]), .B(x[92]), .Z(n26619) );
  XOR U31439 ( .A(n26593), .B(n26594), .Z(n26612) );
  XNOR U31440 ( .A(n26609), .B(n26610), .Z(n26594) );
  XNOR U31441 ( .A(n26604), .B(n26605), .Z(n26610) );
  XNOR U31442 ( .A(n26606), .B(n26607), .Z(n26605) );
  XNOR U31443 ( .A(y[88]), .B(x[88]), .Z(n26607) );
  XNOR U31444 ( .A(y[89]), .B(x[89]), .Z(n26606) );
  XNOR U31445 ( .A(y[87]), .B(x[87]), .Z(n26604) );
  XNOR U31446 ( .A(n26598), .B(n26599), .Z(n26609) );
  XNOR U31447 ( .A(y[84]), .B(x[84]), .Z(n26599) );
  XNOR U31448 ( .A(n26600), .B(n26601), .Z(n26598) );
  XNOR U31449 ( .A(y[85]), .B(x[85]), .Z(n26601) );
  XNOR U31450 ( .A(y[86]), .B(x[86]), .Z(n26600) );
  XOR U31451 ( .A(n26592), .B(n26591), .Z(n26593) );
  XNOR U31452 ( .A(n26587), .B(n26588), .Z(n26591) );
  XNOR U31453 ( .A(y[81]), .B(x[81]), .Z(n26588) );
  XNOR U31454 ( .A(n26589), .B(n26590), .Z(n26587) );
  XNOR U31455 ( .A(y[82]), .B(x[82]), .Z(n26590) );
  XNOR U31456 ( .A(y[83]), .B(x[83]), .Z(n26589) );
  XNOR U31457 ( .A(n26581), .B(n26582), .Z(n26592) );
  XNOR U31458 ( .A(y[78]), .B(x[78]), .Z(n26582) );
  XNOR U31459 ( .A(n26583), .B(n26584), .Z(n26581) );
  XNOR U31460 ( .A(y[79]), .B(x[79]), .Z(n26584) );
  XNOR U31461 ( .A(y[80]), .B(x[80]), .Z(n26583) );
  NAND U31462 ( .A(n26648), .B(n26649), .Z(N27969) );
  NANDN U31463 ( .A(n26650), .B(n26651), .Z(n26649) );
  OR U31464 ( .A(n26652), .B(n26653), .Z(n26651) );
  NAND U31465 ( .A(n26652), .B(n26653), .Z(n26648) );
  XOR U31466 ( .A(n26652), .B(n26654), .Z(N27968) );
  XNOR U31467 ( .A(n26650), .B(n26653), .Z(n26654) );
  AND U31468 ( .A(n26655), .B(n26656), .Z(n26653) );
  NANDN U31469 ( .A(n26657), .B(n26658), .Z(n26656) );
  NANDN U31470 ( .A(n26659), .B(n26660), .Z(n26658) );
  NANDN U31471 ( .A(n26660), .B(n26659), .Z(n26655) );
  NAND U31472 ( .A(n26661), .B(n26662), .Z(n26650) );
  NANDN U31473 ( .A(n26663), .B(n26664), .Z(n26662) );
  OR U31474 ( .A(n26665), .B(n26666), .Z(n26664) );
  NAND U31475 ( .A(n26666), .B(n26665), .Z(n26661) );
  AND U31476 ( .A(n26667), .B(n26668), .Z(n26652) );
  NANDN U31477 ( .A(n26669), .B(n26670), .Z(n26668) );
  NANDN U31478 ( .A(n26671), .B(n26672), .Z(n26670) );
  NANDN U31479 ( .A(n26672), .B(n26671), .Z(n26667) );
  XOR U31480 ( .A(n26666), .B(n26673), .Z(N27967) );
  XOR U31481 ( .A(n26663), .B(n26665), .Z(n26673) );
  XNOR U31482 ( .A(n26659), .B(n26674), .Z(n26665) );
  XNOR U31483 ( .A(n26657), .B(n26660), .Z(n26674) );
  NAND U31484 ( .A(n26675), .B(n26676), .Z(n26660) );
  NAND U31485 ( .A(n26677), .B(n26678), .Z(n26676) );
  OR U31486 ( .A(n26679), .B(n26680), .Z(n26677) );
  NANDN U31487 ( .A(n26681), .B(n26679), .Z(n26675) );
  IV U31488 ( .A(n26680), .Z(n26681) );
  NAND U31489 ( .A(n26682), .B(n26683), .Z(n26657) );
  NAND U31490 ( .A(n26684), .B(n26685), .Z(n26683) );
  NANDN U31491 ( .A(n26686), .B(n26687), .Z(n26684) );
  NANDN U31492 ( .A(n26687), .B(n26686), .Z(n26682) );
  AND U31493 ( .A(n26688), .B(n26689), .Z(n26659) );
  NAND U31494 ( .A(n26690), .B(n26691), .Z(n26689) );
  OR U31495 ( .A(n26692), .B(n26693), .Z(n26690) );
  NANDN U31496 ( .A(n26694), .B(n26692), .Z(n26688) );
  NAND U31497 ( .A(n26695), .B(n26696), .Z(n26663) );
  NANDN U31498 ( .A(n26697), .B(n26698), .Z(n26696) );
  OR U31499 ( .A(n26699), .B(n26700), .Z(n26698) );
  NANDN U31500 ( .A(n26701), .B(n26699), .Z(n26695) );
  IV U31501 ( .A(n26700), .Z(n26701) );
  XNOR U31502 ( .A(n26671), .B(n26702), .Z(n26666) );
  XNOR U31503 ( .A(n26669), .B(n26672), .Z(n26702) );
  NAND U31504 ( .A(n26703), .B(n26704), .Z(n26672) );
  NAND U31505 ( .A(n26705), .B(n26706), .Z(n26704) );
  OR U31506 ( .A(n26707), .B(n26708), .Z(n26705) );
  NANDN U31507 ( .A(n26709), .B(n26707), .Z(n26703) );
  IV U31508 ( .A(n26708), .Z(n26709) );
  NAND U31509 ( .A(n26710), .B(n26711), .Z(n26669) );
  NAND U31510 ( .A(n26712), .B(n26713), .Z(n26711) );
  NANDN U31511 ( .A(n26714), .B(n26715), .Z(n26712) );
  NANDN U31512 ( .A(n26715), .B(n26714), .Z(n26710) );
  AND U31513 ( .A(n26716), .B(n26717), .Z(n26671) );
  NAND U31514 ( .A(n26718), .B(n26719), .Z(n26717) );
  OR U31515 ( .A(n26720), .B(n26721), .Z(n26718) );
  NANDN U31516 ( .A(n26722), .B(n26720), .Z(n26716) );
  XNOR U31517 ( .A(n26697), .B(n26723), .Z(N27966) );
  XOR U31518 ( .A(n26699), .B(n26700), .Z(n26723) );
  XNOR U31519 ( .A(n26713), .B(n26724), .Z(n26700) );
  XOR U31520 ( .A(n26714), .B(n26715), .Z(n26724) );
  XOR U31521 ( .A(n26720), .B(n26725), .Z(n26715) );
  XOR U31522 ( .A(n26719), .B(n26722), .Z(n26725) );
  IV U31523 ( .A(n26721), .Z(n26722) );
  NAND U31524 ( .A(n26726), .B(n26727), .Z(n26721) );
  OR U31525 ( .A(n26728), .B(n26729), .Z(n26727) );
  OR U31526 ( .A(n26730), .B(n26731), .Z(n26726) );
  NAND U31527 ( .A(n26732), .B(n26733), .Z(n26719) );
  OR U31528 ( .A(n26734), .B(n26735), .Z(n26733) );
  OR U31529 ( .A(n26736), .B(n26737), .Z(n26732) );
  NOR U31530 ( .A(n26738), .B(n26739), .Z(n26720) );
  ANDN U31531 ( .B(n26740), .A(n26741), .Z(n26714) );
  XNOR U31532 ( .A(n26707), .B(n26742), .Z(n26713) );
  XNOR U31533 ( .A(n26706), .B(n26708), .Z(n26742) );
  NAND U31534 ( .A(n26743), .B(n26744), .Z(n26708) );
  OR U31535 ( .A(n26745), .B(n26746), .Z(n26744) );
  OR U31536 ( .A(n26747), .B(n26748), .Z(n26743) );
  NAND U31537 ( .A(n26749), .B(n26750), .Z(n26706) );
  OR U31538 ( .A(n26751), .B(n26752), .Z(n26750) );
  OR U31539 ( .A(n26753), .B(n26754), .Z(n26749) );
  ANDN U31540 ( .B(n26755), .A(n26756), .Z(n26707) );
  IV U31541 ( .A(n26757), .Z(n26755) );
  ANDN U31542 ( .B(n26758), .A(n26759), .Z(n26699) );
  XOR U31543 ( .A(n26685), .B(n26760), .Z(n26697) );
  XOR U31544 ( .A(n26686), .B(n26687), .Z(n26760) );
  XOR U31545 ( .A(n26692), .B(n26761), .Z(n26687) );
  XOR U31546 ( .A(n26691), .B(n26694), .Z(n26761) );
  IV U31547 ( .A(n26693), .Z(n26694) );
  NAND U31548 ( .A(n26762), .B(n26763), .Z(n26693) );
  OR U31549 ( .A(n26764), .B(n26765), .Z(n26763) );
  OR U31550 ( .A(n26766), .B(n26767), .Z(n26762) );
  NAND U31551 ( .A(n26768), .B(n26769), .Z(n26691) );
  OR U31552 ( .A(n26770), .B(n26771), .Z(n26769) );
  OR U31553 ( .A(n26772), .B(n26773), .Z(n26768) );
  NOR U31554 ( .A(n26774), .B(n26775), .Z(n26692) );
  ANDN U31555 ( .B(n26776), .A(n26777), .Z(n26686) );
  IV U31556 ( .A(n26778), .Z(n26776) );
  XNOR U31557 ( .A(n26679), .B(n26779), .Z(n26685) );
  XNOR U31558 ( .A(n26678), .B(n26680), .Z(n26779) );
  NAND U31559 ( .A(n26780), .B(n26781), .Z(n26680) );
  OR U31560 ( .A(n26782), .B(n26783), .Z(n26781) );
  OR U31561 ( .A(n26784), .B(n26785), .Z(n26780) );
  NAND U31562 ( .A(n26786), .B(n26787), .Z(n26678) );
  OR U31563 ( .A(n26788), .B(n26789), .Z(n26787) );
  OR U31564 ( .A(n26790), .B(n26791), .Z(n26786) );
  ANDN U31565 ( .B(n26792), .A(n26793), .Z(n26679) );
  IV U31566 ( .A(n26794), .Z(n26792) );
  XNOR U31567 ( .A(n26759), .B(n26758), .Z(N27965) );
  XOR U31568 ( .A(n26778), .B(n26777), .Z(n26758) );
  XNOR U31569 ( .A(n26793), .B(n26794), .Z(n26777) );
  XNOR U31570 ( .A(n26788), .B(n26789), .Z(n26794) );
  XNOR U31571 ( .A(n26790), .B(n26791), .Z(n26789) );
  XNOR U31572 ( .A(y[76]), .B(x[76]), .Z(n26791) );
  XNOR U31573 ( .A(y[77]), .B(x[77]), .Z(n26790) );
  XNOR U31574 ( .A(y[75]), .B(x[75]), .Z(n26788) );
  XNOR U31575 ( .A(n26782), .B(n26783), .Z(n26793) );
  XNOR U31576 ( .A(y[72]), .B(x[72]), .Z(n26783) );
  XNOR U31577 ( .A(n26784), .B(n26785), .Z(n26782) );
  XNOR U31578 ( .A(y[73]), .B(x[73]), .Z(n26785) );
  XNOR U31579 ( .A(y[74]), .B(x[74]), .Z(n26784) );
  XNOR U31580 ( .A(n26775), .B(n26774), .Z(n26778) );
  XNOR U31581 ( .A(n26770), .B(n26771), .Z(n26774) );
  XNOR U31582 ( .A(y[69]), .B(x[69]), .Z(n26771) );
  XNOR U31583 ( .A(n26772), .B(n26773), .Z(n26770) );
  XNOR U31584 ( .A(y[70]), .B(x[70]), .Z(n26773) );
  XNOR U31585 ( .A(y[71]), .B(x[71]), .Z(n26772) );
  XNOR U31586 ( .A(n26764), .B(n26765), .Z(n26775) );
  XNOR U31587 ( .A(y[66]), .B(x[66]), .Z(n26765) );
  XNOR U31588 ( .A(n26766), .B(n26767), .Z(n26764) );
  XNOR U31589 ( .A(y[67]), .B(x[67]), .Z(n26767) );
  XNOR U31590 ( .A(y[68]), .B(x[68]), .Z(n26766) );
  XOR U31591 ( .A(n26740), .B(n26741), .Z(n26759) );
  XNOR U31592 ( .A(n26756), .B(n26757), .Z(n26741) );
  XNOR U31593 ( .A(n26751), .B(n26752), .Z(n26757) );
  XNOR U31594 ( .A(n26753), .B(n26754), .Z(n26752) );
  XNOR U31595 ( .A(y[64]), .B(x[64]), .Z(n26754) );
  XNOR U31596 ( .A(y[65]), .B(x[65]), .Z(n26753) );
  XNOR U31597 ( .A(y[63]), .B(x[63]), .Z(n26751) );
  XNOR U31598 ( .A(n26745), .B(n26746), .Z(n26756) );
  XNOR U31599 ( .A(y[60]), .B(x[60]), .Z(n26746) );
  XNOR U31600 ( .A(n26747), .B(n26748), .Z(n26745) );
  XNOR U31601 ( .A(y[61]), .B(x[61]), .Z(n26748) );
  XNOR U31602 ( .A(y[62]), .B(x[62]), .Z(n26747) );
  XOR U31603 ( .A(n26739), .B(n26738), .Z(n26740) );
  XNOR U31604 ( .A(n26734), .B(n26735), .Z(n26738) );
  XNOR U31605 ( .A(y[57]), .B(x[57]), .Z(n26735) );
  XNOR U31606 ( .A(n26736), .B(n26737), .Z(n26734) );
  XNOR U31607 ( .A(y[58]), .B(x[58]), .Z(n26737) );
  XNOR U31608 ( .A(y[59]), .B(x[59]), .Z(n26736) );
  XNOR U31609 ( .A(n26728), .B(n26729), .Z(n26739) );
  XNOR U31610 ( .A(y[54]), .B(x[54]), .Z(n26729) );
  XNOR U31611 ( .A(n26730), .B(n26731), .Z(n26728) );
  XNOR U31612 ( .A(y[55]), .B(x[55]), .Z(n26731) );
  XNOR U31613 ( .A(y[56]), .B(x[56]), .Z(n26730) );
  NAND U31614 ( .A(n26795), .B(n26796), .Z(N27957) );
  NANDN U31615 ( .A(n26797), .B(n26798), .Z(n26796) );
  OR U31616 ( .A(n26799), .B(n26800), .Z(n26798) );
  NAND U31617 ( .A(n26799), .B(n26800), .Z(n26795) );
  XOR U31618 ( .A(n26799), .B(n26801), .Z(N27956) );
  XNOR U31619 ( .A(n26797), .B(n26800), .Z(n26801) );
  AND U31620 ( .A(n26802), .B(n26803), .Z(n26800) );
  NANDN U31621 ( .A(n26804), .B(n26805), .Z(n26803) );
  NANDN U31622 ( .A(n26806), .B(n26807), .Z(n26805) );
  NANDN U31623 ( .A(n26807), .B(n26806), .Z(n26802) );
  NAND U31624 ( .A(n26808), .B(n26809), .Z(n26797) );
  NANDN U31625 ( .A(n26810), .B(n26811), .Z(n26809) );
  OR U31626 ( .A(n26812), .B(n26813), .Z(n26811) );
  NAND U31627 ( .A(n26813), .B(n26812), .Z(n26808) );
  AND U31628 ( .A(n26814), .B(n26815), .Z(n26799) );
  NANDN U31629 ( .A(n26816), .B(n26817), .Z(n26815) );
  NANDN U31630 ( .A(n26818), .B(n26819), .Z(n26817) );
  NANDN U31631 ( .A(n26819), .B(n26818), .Z(n26814) );
  XOR U31632 ( .A(n26813), .B(n26820), .Z(N27955) );
  XOR U31633 ( .A(n26810), .B(n26812), .Z(n26820) );
  XNOR U31634 ( .A(n26806), .B(n26821), .Z(n26812) );
  XNOR U31635 ( .A(n26804), .B(n26807), .Z(n26821) );
  NAND U31636 ( .A(n26822), .B(n26823), .Z(n26807) );
  NAND U31637 ( .A(n26824), .B(n26825), .Z(n26823) );
  OR U31638 ( .A(n26826), .B(n26827), .Z(n26824) );
  NANDN U31639 ( .A(n26828), .B(n26826), .Z(n26822) );
  IV U31640 ( .A(n26827), .Z(n26828) );
  NAND U31641 ( .A(n26829), .B(n26830), .Z(n26804) );
  NAND U31642 ( .A(n26831), .B(n26832), .Z(n26830) );
  NANDN U31643 ( .A(n26833), .B(n26834), .Z(n26831) );
  NANDN U31644 ( .A(n26834), .B(n26833), .Z(n26829) );
  AND U31645 ( .A(n26835), .B(n26836), .Z(n26806) );
  NAND U31646 ( .A(n26837), .B(n26838), .Z(n26836) );
  OR U31647 ( .A(n26839), .B(n26840), .Z(n26837) );
  NANDN U31648 ( .A(n26841), .B(n26839), .Z(n26835) );
  NAND U31649 ( .A(n26842), .B(n26843), .Z(n26810) );
  NANDN U31650 ( .A(n26844), .B(n26845), .Z(n26843) );
  OR U31651 ( .A(n26846), .B(n26847), .Z(n26845) );
  NANDN U31652 ( .A(n26848), .B(n26846), .Z(n26842) );
  IV U31653 ( .A(n26847), .Z(n26848) );
  XNOR U31654 ( .A(n26818), .B(n26849), .Z(n26813) );
  XNOR U31655 ( .A(n26816), .B(n26819), .Z(n26849) );
  NAND U31656 ( .A(n26850), .B(n26851), .Z(n26819) );
  NAND U31657 ( .A(n26852), .B(n26853), .Z(n26851) );
  OR U31658 ( .A(n26854), .B(n26855), .Z(n26852) );
  NANDN U31659 ( .A(n26856), .B(n26854), .Z(n26850) );
  IV U31660 ( .A(n26855), .Z(n26856) );
  NAND U31661 ( .A(n26857), .B(n26858), .Z(n26816) );
  NAND U31662 ( .A(n26859), .B(n26860), .Z(n26858) );
  NANDN U31663 ( .A(n26861), .B(n26862), .Z(n26859) );
  NANDN U31664 ( .A(n26862), .B(n26861), .Z(n26857) );
  AND U31665 ( .A(n26863), .B(n26864), .Z(n26818) );
  NAND U31666 ( .A(n26865), .B(n26866), .Z(n26864) );
  OR U31667 ( .A(n26867), .B(n26868), .Z(n26865) );
  NANDN U31668 ( .A(n26869), .B(n26867), .Z(n26863) );
  XNOR U31669 ( .A(n26844), .B(n26870), .Z(N27954) );
  XOR U31670 ( .A(n26846), .B(n26847), .Z(n26870) );
  XNOR U31671 ( .A(n26860), .B(n26871), .Z(n26847) );
  XOR U31672 ( .A(n26861), .B(n26862), .Z(n26871) );
  XOR U31673 ( .A(n26867), .B(n26872), .Z(n26862) );
  XOR U31674 ( .A(n26866), .B(n26869), .Z(n26872) );
  IV U31675 ( .A(n26868), .Z(n26869) );
  NAND U31676 ( .A(n26873), .B(n26874), .Z(n26868) );
  OR U31677 ( .A(n26875), .B(n26876), .Z(n26874) );
  OR U31678 ( .A(n26877), .B(n26878), .Z(n26873) );
  NAND U31679 ( .A(n26879), .B(n26880), .Z(n26866) );
  OR U31680 ( .A(n26881), .B(n26882), .Z(n26880) );
  OR U31681 ( .A(n26883), .B(n26884), .Z(n26879) );
  NOR U31682 ( .A(n26885), .B(n26886), .Z(n26867) );
  ANDN U31683 ( .B(n26887), .A(n26888), .Z(n26861) );
  XNOR U31684 ( .A(n26854), .B(n26889), .Z(n26860) );
  XNOR U31685 ( .A(n26853), .B(n26855), .Z(n26889) );
  NAND U31686 ( .A(n26890), .B(n26891), .Z(n26855) );
  OR U31687 ( .A(n26892), .B(n26893), .Z(n26891) );
  OR U31688 ( .A(n26894), .B(n26895), .Z(n26890) );
  NAND U31689 ( .A(n26896), .B(n26897), .Z(n26853) );
  OR U31690 ( .A(n26898), .B(n26899), .Z(n26897) );
  OR U31691 ( .A(n26900), .B(n26901), .Z(n26896) );
  ANDN U31692 ( .B(n26902), .A(n26903), .Z(n26854) );
  IV U31693 ( .A(n26904), .Z(n26902) );
  ANDN U31694 ( .B(n26905), .A(n26906), .Z(n26846) );
  XOR U31695 ( .A(n26832), .B(n26907), .Z(n26844) );
  XOR U31696 ( .A(n26833), .B(n26834), .Z(n26907) );
  XOR U31697 ( .A(n26839), .B(n26908), .Z(n26834) );
  XOR U31698 ( .A(n26838), .B(n26841), .Z(n26908) );
  IV U31699 ( .A(n26840), .Z(n26841) );
  NAND U31700 ( .A(n26909), .B(n26910), .Z(n26840) );
  OR U31701 ( .A(n26911), .B(n26912), .Z(n26910) );
  OR U31702 ( .A(n26913), .B(n26914), .Z(n26909) );
  NAND U31703 ( .A(n26915), .B(n26916), .Z(n26838) );
  OR U31704 ( .A(n26917), .B(n26918), .Z(n26916) );
  OR U31705 ( .A(n26919), .B(n26920), .Z(n26915) );
  NOR U31706 ( .A(n26921), .B(n26922), .Z(n26839) );
  ANDN U31707 ( .B(n26923), .A(n26924), .Z(n26833) );
  IV U31708 ( .A(n26925), .Z(n26923) );
  XNOR U31709 ( .A(n26826), .B(n26926), .Z(n26832) );
  XNOR U31710 ( .A(n26825), .B(n26827), .Z(n26926) );
  NAND U31711 ( .A(n26927), .B(n26928), .Z(n26827) );
  OR U31712 ( .A(n26929), .B(n26930), .Z(n26928) );
  OR U31713 ( .A(n26931), .B(n26932), .Z(n26927) );
  NAND U31714 ( .A(n26933), .B(n26934), .Z(n26825) );
  OR U31715 ( .A(n26935), .B(n26936), .Z(n26934) );
  OR U31716 ( .A(n26937), .B(n26938), .Z(n26933) );
  ANDN U31717 ( .B(n26939), .A(n26940), .Z(n26826) );
  IV U31718 ( .A(n26941), .Z(n26939) );
  XNOR U31719 ( .A(n26906), .B(n26905), .Z(N27953) );
  XOR U31720 ( .A(n26925), .B(n26924), .Z(n26905) );
  XNOR U31721 ( .A(n26940), .B(n26941), .Z(n26924) );
  XNOR U31722 ( .A(n26935), .B(n26936), .Z(n26941) );
  XNOR U31723 ( .A(n26937), .B(n26938), .Z(n26936) );
  XNOR U31724 ( .A(y[52]), .B(x[52]), .Z(n26938) );
  XNOR U31725 ( .A(y[53]), .B(x[53]), .Z(n26937) );
  XNOR U31726 ( .A(y[51]), .B(x[51]), .Z(n26935) );
  XNOR U31727 ( .A(n26929), .B(n26930), .Z(n26940) );
  XNOR U31728 ( .A(y[48]), .B(x[48]), .Z(n26930) );
  XNOR U31729 ( .A(n26931), .B(n26932), .Z(n26929) );
  XNOR U31730 ( .A(y[49]), .B(x[49]), .Z(n26932) );
  XNOR U31731 ( .A(y[50]), .B(x[50]), .Z(n26931) );
  XNOR U31732 ( .A(n26922), .B(n26921), .Z(n26925) );
  XNOR U31733 ( .A(n26917), .B(n26918), .Z(n26921) );
  XNOR U31734 ( .A(y[45]), .B(x[45]), .Z(n26918) );
  XNOR U31735 ( .A(n26919), .B(n26920), .Z(n26917) );
  XNOR U31736 ( .A(y[46]), .B(x[46]), .Z(n26920) );
  XNOR U31737 ( .A(y[47]), .B(x[47]), .Z(n26919) );
  XNOR U31738 ( .A(n26911), .B(n26912), .Z(n26922) );
  XNOR U31739 ( .A(y[42]), .B(x[42]), .Z(n26912) );
  XNOR U31740 ( .A(n26913), .B(n26914), .Z(n26911) );
  XNOR U31741 ( .A(y[43]), .B(x[43]), .Z(n26914) );
  XNOR U31742 ( .A(y[44]), .B(x[44]), .Z(n26913) );
  XOR U31743 ( .A(n26887), .B(n26888), .Z(n26906) );
  XNOR U31744 ( .A(n26903), .B(n26904), .Z(n26888) );
  XNOR U31745 ( .A(n26898), .B(n26899), .Z(n26904) );
  XNOR U31746 ( .A(n26900), .B(n26901), .Z(n26899) );
  XNOR U31747 ( .A(y[40]), .B(x[40]), .Z(n26901) );
  XNOR U31748 ( .A(y[41]), .B(x[41]), .Z(n26900) );
  XNOR U31749 ( .A(y[39]), .B(x[39]), .Z(n26898) );
  XNOR U31750 ( .A(n26892), .B(n26893), .Z(n26903) );
  XNOR U31751 ( .A(y[36]), .B(x[36]), .Z(n26893) );
  XNOR U31752 ( .A(n26894), .B(n26895), .Z(n26892) );
  XNOR U31753 ( .A(y[37]), .B(x[37]), .Z(n26895) );
  XNOR U31754 ( .A(y[38]), .B(x[38]), .Z(n26894) );
  XOR U31755 ( .A(n26886), .B(n26885), .Z(n26887) );
  XNOR U31756 ( .A(n26881), .B(n26882), .Z(n26885) );
  XNOR U31757 ( .A(y[33]), .B(x[33]), .Z(n26882) );
  XNOR U31758 ( .A(n26883), .B(n26884), .Z(n26881) );
  XNOR U31759 ( .A(y[34]), .B(x[34]), .Z(n26884) );
  XNOR U31760 ( .A(y[35]), .B(x[35]), .Z(n26883) );
  XNOR U31761 ( .A(n26875), .B(n26876), .Z(n26886) );
  XNOR U31762 ( .A(y[30]), .B(x[30]), .Z(n26876) );
  XNOR U31763 ( .A(n26877), .B(n26878), .Z(n26875) );
  XNOR U31764 ( .A(y[31]), .B(x[31]), .Z(n26878) );
  XNOR U31765 ( .A(y[32]), .B(x[32]), .Z(n26877) );
  NAND U31766 ( .A(n26942), .B(n26943), .Z(N27945) );
  NANDN U31767 ( .A(n26944), .B(n26945), .Z(n26943) );
  OR U31768 ( .A(n26946), .B(n26947), .Z(n26945) );
  NAND U31769 ( .A(n26946), .B(n26947), .Z(n26942) );
  XOR U31770 ( .A(n26946), .B(n26948), .Z(N27944) );
  XNOR U31771 ( .A(n26944), .B(n26947), .Z(n26948) );
  AND U31772 ( .A(n26949), .B(n26950), .Z(n26947) );
  NANDN U31773 ( .A(n26951), .B(n26952), .Z(n26950) );
  NANDN U31774 ( .A(n26953), .B(n26954), .Z(n26952) );
  NANDN U31775 ( .A(n26954), .B(n26953), .Z(n26949) );
  NAND U31776 ( .A(n26955), .B(n26956), .Z(n26944) );
  NANDN U31777 ( .A(n26957), .B(n26958), .Z(n26956) );
  OR U31778 ( .A(n26959), .B(n26960), .Z(n26958) );
  NAND U31779 ( .A(n26960), .B(n26959), .Z(n26955) );
  AND U31780 ( .A(n26961), .B(n26962), .Z(n26946) );
  NANDN U31781 ( .A(n26963), .B(n26964), .Z(n26962) );
  NANDN U31782 ( .A(n26965), .B(n26966), .Z(n26964) );
  NANDN U31783 ( .A(n26966), .B(n26965), .Z(n26961) );
  XOR U31784 ( .A(n26960), .B(n26967), .Z(N27943) );
  XOR U31785 ( .A(n26957), .B(n26959), .Z(n26967) );
  XNOR U31786 ( .A(n26953), .B(n26968), .Z(n26959) );
  XNOR U31787 ( .A(n26951), .B(n26954), .Z(n26968) );
  NAND U31788 ( .A(n26969), .B(n26970), .Z(n26954) );
  NAND U31789 ( .A(n26971), .B(n26972), .Z(n26970) );
  OR U31790 ( .A(n26973), .B(n26974), .Z(n26971) );
  NANDN U31791 ( .A(n26975), .B(n26973), .Z(n26969) );
  IV U31792 ( .A(n26974), .Z(n26975) );
  NAND U31793 ( .A(n26976), .B(n26977), .Z(n26951) );
  NAND U31794 ( .A(n26978), .B(n26979), .Z(n26977) );
  NANDN U31795 ( .A(n26980), .B(n26981), .Z(n26978) );
  NANDN U31796 ( .A(n26981), .B(n26980), .Z(n26976) );
  AND U31797 ( .A(n26982), .B(n26983), .Z(n26953) );
  NAND U31798 ( .A(n26984), .B(n26985), .Z(n26983) );
  OR U31799 ( .A(n26986), .B(n26987), .Z(n26984) );
  NANDN U31800 ( .A(n26988), .B(n26986), .Z(n26982) );
  NAND U31801 ( .A(n26989), .B(n26990), .Z(n26957) );
  NANDN U31802 ( .A(n26991), .B(n26992), .Z(n26990) );
  OR U31803 ( .A(n26993), .B(n26994), .Z(n26992) );
  NANDN U31804 ( .A(n26995), .B(n26993), .Z(n26989) );
  IV U31805 ( .A(n26994), .Z(n26995) );
  XNOR U31806 ( .A(n26965), .B(n26996), .Z(n26960) );
  XNOR U31807 ( .A(n26963), .B(n26966), .Z(n26996) );
  NAND U31808 ( .A(n26997), .B(n26998), .Z(n26966) );
  NAND U31809 ( .A(n26999), .B(n27000), .Z(n26998) );
  OR U31810 ( .A(n27001), .B(n27002), .Z(n26999) );
  NANDN U31811 ( .A(n27003), .B(n27001), .Z(n26997) );
  IV U31812 ( .A(n27002), .Z(n27003) );
  NAND U31813 ( .A(n27004), .B(n27005), .Z(n26963) );
  NAND U31814 ( .A(n27006), .B(n27007), .Z(n27005) );
  NANDN U31815 ( .A(n27008), .B(n27009), .Z(n27006) );
  NANDN U31816 ( .A(n27009), .B(n27008), .Z(n27004) );
  AND U31817 ( .A(n27010), .B(n27011), .Z(n26965) );
  NAND U31818 ( .A(n27012), .B(n27013), .Z(n27011) );
  OR U31819 ( .A(n27014), .B(n27015), .Z(n27012) );
  NANDN U31820 ( .A(n27016), .B(n27014), .Z(n27010) );
  IV U31821 ( .A(n27015), .Z(n27016) );
  XNOR U31822 ( .A(n26991), .B(n27017), .Z(N27942) );
  XOR U31823 ( .A(n26993), .B(n26994), .Z(n27017) );
  XNOR U31824 ( .A(n27007), .B(n27018), .Z(n26994) );
  XOR U31825 ( .A(n27008), .B(n27009), .Z(n27018) );
  XOR U31826 ( .A(n27014), .B(n27019), .Z(n27009) );
  XNOR U31827 ( .A(n27013), .B(n27015), .Z(n27019) );
  NAND U31828 ( .A(n27020), .B(n27021), .Z(n27015) );
  OR U31829 ( .A(n27022), .B(n27023), .Z(n27021) );
  IV U31830 ( .A(n27024), .Z(n27023) );
  OR U31831 ( .A(n27025), .B(n27026), .Z(n27020) );
  NAND U31832 ( .A(n27027), .B(n27028), .Z(n27013) );
  OR U31833 ( .A(n27029), .B(n27030), .Z(n27028) );
  OR U31834 ( .A(n27031), .B(n27032), .Z(n27027) );
  ANDN U31835 ( .B(n27033), .A(n27034), .Z(n27014) );
  IV U31836 ( .A(n27035), .Z(n27033) );
  NOR U31837 ( .A(n27036), .B(n27037), .Z(n27008) );
  XNOR U31838 ( .A(n27001), .B(n27038), .Z(n27007) );
  XNOR U31839 ( .A(n27000), .B(n27002), .Z(n27038) );
  NAND U31840 ( .A(n27039), .B(n27040), .Z(n27002) );
  OR U31841 ( .A(n27041), .B(n27042), .Z(n27040) );
  OR U31842 ( .A(n27043), .B(n27044), .Z(n27039) );
  NAND U31843 ( .A(n27045), .B(n27046), .Z(n27000) );
  OR U31844 ( .A(n27047), .B(n27048), .Z(n27046) );
  OR U31845 ( .A(n27049), .B(n27050), .Z(n27045) );
  ANDN U31846 ( .B(n27051), .A(n27052), .Z(n27001) );
  IV U31847 ( .A(n27053), .Z(n27051) );
  ANDN U31848 ( .B(n27054), .A(n27055), .Z(n26993) );
  XOR U31849 ( .A(n26979), .B(n27056), .Z(n26991) );
  XOR U31850 ( .A(n26980), .B(n26981), .Z(n27056) );
  XOR U31851 ( .A(n26986), .B(n27057), .Z(n26981) );
  XOR U31852 ( .A(n26985), .B(n26988), .Z(n27057) );
  IV U31853 ( .A(n26987), .Z(n26988) );
  NAND U31854 ( .A(n27058), .B(n27059), .Z(n26987) );
  OR U31855 ( .A(n27060), .B(n27061), .Z(n27059) );
  OR U31856 ( .A(n27062), .B(n27063), .Z(n27058) );
  NAND U31857 ( .A(n27064), .B(n27065), .Z(n26985) );
  OR U31858 ( .A(n27066), .B(n27067), .Z(n27065) );
  OR U31859 ( .A(n27068), .B(n27069), .Z(n27064) );
  NOR U31860 ( .A(n27070), .B(n27071), .Z(n26986) );
  ANDN U31861 ( .B(n27072), .A(n27073), .Z(n26980) );
  IV U31862 ( .A(n27074), .Z(n27072) );
  XNOR U31863 ( .A(n26973), .B(n27075), .Z(n26979) );
  XNOR U31864 ( .A(n26972), .B(n26974), .Z(n27075) );
  NAND U31865 ( .A(n27076), .B(n27077), .Z(n26974) );
  OR U31866 ( .A(n27078), .B(n27079), .Z(n27077) );
  OR U31867 ( .A(n27080), .B(n27081), .Z(n27076) );
  NAND U31868 ( .A(n27082), .B(n27083), .Z(n26972) );
  OR U31869 ( .A(n27084), .B(n27085), .Z(n27083) );
  OR U31870 ( .A(n27086), .B(n27087), .Z(n27082) );
  ANDN U31871 ( .B(n27088), .A(n27089), .Z(n26973) );
  IV U31872 ( .A(n27090), .Z(n27088) );
  XNOR U31873 ( .A(n27055), .B(n27054), .Z(N27941) );
  XOR U31874 ( .A(n27074), .B(n27073), .Z(n27054) );
  XNOR U31875 ( .A(n27089), .B(n27090), .Z(n27073) );
  XNOR U31876 ( .A(n27084), .B(n27085), .Z(n27090) );
  XNOR U31877 ( .A(n27086), .B(n27087), .Z(n27085) );
  XNOR U31878 ( .A(y[28]), .B(x[28]), .Z(n27087) );
  XNOR U31879 ( .A(y[29]), .B(x[29]), .Z(n27086) );
  XNOR U31880 ( .A(y[27]), .B(x[27]), .Z(n27084) );
  XNOR U31881 ( .A(n27078), .B(n27079), .Z(n27089) );
  XNOR U31882 ( .A(y[24]), .B(x[24]), .Z(n27079) );
  XNOR U31883 ( .A(n27080), .B(n27081), .Z(n27078) );
  XNOR U31884 ( .A(y[25]), .B(x[25]), .Z(n27081) );
  XNOR U31885 ( .A(y[26]), .B(x[26]), .Z(n27080) );
  XNOR U31886 ( .A(n27071), .B(n27070), .Z(n27074) );
  XNOR U31887 ( .A(n27066), .B(n27067), .Z(n27070) );
  XNOR U31888 ( .A(y[21]), .B(x[21]), .Z(n27067) );
  XNOR U31889 ( .A(n27068), .B(n27069), .Z(n27066) );
  XNOR U31890 ( .A(y[22]), .B(x[22]), .Z(n27069) );
  XNOR U31891 ( .A(y[23]), .B(x[23]), .Z(n27068) );
  XNOR U31892 ( .A(n27060), .B(n27061), .Z(n27071) );
  XNOR U31893 ( .A(y[18]), .B(x[18]), .Z(n27061) );
  XNOR U31894 ( .A(n27062), .B(n27063), .Z(n27060) );
  XNOR U31895 ( .A(y[19]), .B(x[19]), .Z(n27063) );
  XNOR U31896 ( .A(y[20]), .B(x[20]), .Z(n27062) );
  XNOR U31897 ( .A(n27036), .B(n27037), .Z(n27055) );
  XNOR U31898 ( .A(n27052), .B(n27053), .Z(n27037) );
  XNOR U31899 ( .A(n27047), .B(n27048), .Z(n27053) );
  XNOR U31900 ( .A(n27049), .B(n27050), .Z(n27048) );
  XNOR U31901 ( .A(y[16]), .B(x[16]), .Z(n27050) );
  XNOR U31902 ( .A(y[17]), .B(x[17]), .Z(n27049) );
  XNOR U31903 ( .A(y[15]), .B(x[15]), .Z(n27047) );
  XNOR U31904 ( .A(n27041), .B(n27042), .Z(n27052) );
  XNOR U31905 ( .A(y[12]), .B(x[12]), .Z(n27042) );
  XNOR U31906 ( .A(n27043), .B(n27044), .Z(n27041) );
  XNOR U31907 ( .A(y[13]), .B(x[13]), .Z(n27044) );
  XNOR U31908 ( .A(y[14]), .B(x[14]), .Z(n27043) );
  XNOR U31909 ( .A(n27035), .B(n27034), .Z(n27036) );
  XNOR U31910 ( .A(n27029), .B(n27030), .Z(n27034) );
  XNOR U31911 ( .A(y[9]), .B(x[9]), .Z(n27030) );
  XNOR U31912 ( .A(n27031), .B(n27032), .Z(n27029) );
  XNOR U31913 ( .A(y[10]), .B(x[10]), .Z(n27032) );
  XNOR U31914 ( .A(y[11]), .B(x[11]), .Z(n27031) );
  XOR U31915 ( .A(n27022), .B(n27024), .Z(n27035) );
  XOR U31916 ( .A(n27025), .B(n27026), .Z(n27024) );
  XNOR U31917 ( .A(y[7]), .B(x[7]), .Z(n27026) );
  XNOR U31918 ( .A(y[8]), .B(x[8]), .Z(n27025) );
  XNOR U31919 ( .A(y[6]), .B(x[6]), .Z(n27022) );
  ANDN U31920 ( .B(n27091), .A(n27092), .Z(N27933) );
  XNOR U31921 ( .A(n27092), .B(n27091), .Z(N27932) );
  ANDN U31922 ( .B(n27093), .A(n27094), .Z(n27091) );
  NAND U31923 ( .A(n27095), .B(n27096), .Z(n27092) );
  NANDN U31924 ( .A(n27097), .B(n27098), .Z(n27096) );
  OR U31925 ( .A(n27099), .B(n27100), .Z(n27098) );
  NAND U31926 ( .A(n27099), .B(n27100), .Z(n27095) );
  XNOR U31927 ( .A(n27099), .B(n27101), .Z(N27931) );
  XNOR U31928 ( .A(n27097), .B(n27100), .Z(n27101) );
  AND U31929 ( .A(n27102), .B(n27103), .Z(n27100) );
  NAND U31930 ( .A(n27104), .B(n27105), .Z(n27103) );
  OR U31931 ( .A(n27106), .B(n27107), .Z(n27104) );
  NANDN U31932 ( .A(n27108), .B(n27106), .Z(n27102) );
  IV U31933 ( .A(n27107), .Z(n27108) );
  NAND U31934 ( .A(n27109), .B(n27110), .Z(n27097) );
  NANDN U31935 ( .A(n27111), .B(n27112), .Z(n27110) );
  OR U31936 ( .A(n27113), .B(n27114), .Z(n27112) );
  NAND U31937 ( .A(n27114), .B(n27113), .Z(n27109) );
  XOR U31938 ( .A(n27094), .B(n27093), .Z(n27099) );
  NAND U31939 ( .A(n27115), .B(n27116), .Z(n27093) );
  OR U31940 ( .A(n27117), .B(n27118), .Z(n27116) );
  OR U31941 ( .A(n27119), .B(n27120), .Z(n27115) );
  AND U31942 ( .A(n27121), .B(n27122), .Z(n27094) );
  NAND U31943 ( .A(n27123), .B(n27124), .Z(n27122) );
  NAND U31944 ( .A(n27125), .B(n27126), .Z(n27123) );
  OR U31945 ( .A(n27125), .B(n27126), .Z(n27121) );
  XNOR U31946 ( .A(n27111), .B(n27127), .Z(N27930) );
  XOR U31947 ( .A(n27113), .B(n27114), .Z(n27127) );
  XNOR U31948 ( .A(n27106), .B(n27128), .Z(n27114) );
  XNOR U31949 ( .A(n27105), .B(n27107), .Z(n27128) );
  NAND U31950 ( .A(n27129), .B(n27130), .Z(n27107) );
  OR U31951 ( .A(n27131), .B(n27132), .Z(n27130) );
  OR U31952 ( .A(n27133), .B(n27134), .Z(n27129) );
  NAND U31953 ( .A(n27135), .B(n27136), .Z(n27105) );
  OR U31954 ( .A(n27137), .B(n27138), .Z(n27136) );
  OR U31955 ( .A(n27139), .B(n27140), .Z(n27135) );
  ANDN U31956 ( .B(n27141), .A(n27142), .Z(n27106) );
  IV U31957 ( .A(n27143), .Z(n27141) );
  ANDN U31958 ( .B(n27144), .A(n27145), .Z(n27113) );
  XNOR U31959 ( .A(n27124), .B(n27146), .Z(n27111) );
  XOR U31960 ( .A(n27126), .B(n27125), .Z(n27146) );
  OR U31961 ( .A(n27147), .B(n27148), .Z(n27125) );
  AND U31962 ( .A(n27149), .B(n27150), .Z(n27126) );
  OR U31963 ( .A(n27151), .B(n27152), .Z(n27150) );
  OR U31964 ( .A(n27153), .B(n27154), .Z(n27149) );
  XOR U31965 ( .A(n27117), .B(n27118), .Z(n27124) );
  XOR U31966 ( .A(n27155), .B(n27119), .Z(n27118) );
  AND U31967 ( .A(n27156), .B(n27157), .Z(n27119) );
  OR U31968 ( .A(n27158), .B(n27159), .Z(n27157) );
  OR U31969 ( .A(n27160), .B(n27161), .Z(n27156) );
  IV U31970 ( .A(n27120), .Z(n27155) );
  AND U31971 ( .A(n27162), .B(n27163), .Z(n27120) );
  NANDN U31972 ( .A(n27164), .B(n27165), .Z(n27163) );
  OR U31973 ( .A(n27166), .B(n27167), .Z(n27162) );
  AND U31974 ( .A(n27168), .B(n27169), .Z(n27117) );
  NANDN U31975 ( .A(n27170), .B(n27171), .Z(n27169) );
  NANDN U31976 ( .A(n27172), .B(n27173), .Z(n27168) );
  XNOR U31977 ( .A(n27145), .B(n27144), .Z(N27929) );
  XOR U31978 ( .A(n27148), .B(n27147), .Z(n27144) );
  XOR U31979 ( .A(n27170), .B(n27171), .Z(n27147) );
  XNOR U31980 ( .A(n27172), .B(n27173), .Z(n27171) );
  XOR U31981 ( .A(n27159), .B(n27158), .Z(n27173) );
  XNOR U31982 ( .A(y[0]), .B(x[0]), .Z(n27158) );
  XNOR U31983 ( .A(n27161), .B(n27160), .Z(n27159) );
  XNOR U31984 ( .A(y[1]), .B(x[1]), .Z(n27160) );
  XNOR U31985 ( .A(y[2]), .B(x[2]), .Z(n27161) );
  XOR U31986 ( .A(n27165), .B(n27164), .Z(n27172) );
  XNOR U31987 ( .A(y[3]), .B(x[3]), .Z(n27164) );
  XOR U31988 ( .A(n27167), .B(n27166), .Z(n27165) );
  XNOR U31989 ( .A(y[4]), .B(x[4]), .Z(n27166) );
  XNOR U31990 ( .A(y[5]), .B(x[5]), .Z(n27167) );
  XNOR U31991 ( .A(y[3999]), .B(x[3999]), .Z(n27170) );
  XNOR U31992 ( .A(n27151), .B(n27152), .Z(n27148) );
  XNOR U31993 ( .A(y[3996]), .B(x[3996]), .Z(n27152) );
  XNOR U31994 ( .A(n27153), .B(n27154), .Z(n27151) );
  XNOR U31995 ( .A(y[3997]), .B(x[3997]), .Z(n27154) );
  XNOR U31996 ( .A(y[3998]), .B(x[3998]), .Z(n27153) );
  XNOR U31997 ( .A(n27142), .B(n27143), .Z(n27145) );
  XNOR U31998 ( .A(n27137), .B(n27138), .Z(n27143) );
  XNOR U31999 ( .A(n27139), .B(n27140), .Z(n27138) );
  XNOR U32000 ( .A(y[3994]), .B(x[3994]), .Z(n27140) );
  XNOR U32001 ( .A(y[3995]), .B(x[3995]), .Z(n27139) );
  XNOR U32002 ( .A(y[3993]), .B(x[3993]), .Z(n27137) );
  XNOR U32003 ( .A(n27131), .B(n27132), .Z(n27142) );
  XNOR U32004 ( .A(y[3990]), .B(x[3990]), .Z(n27132) );
  XNOR U32005 ( .A(n27133), .B(n27134), .Z(n27131) );
  XNOR U32006 ( .A(y[3991]), .B(x[3991]), .Z(n27134) );
  XNOR U32007 ( .A(y[3992]), .B(x[3992]), .Z(n27133) );
endmodule

