
module sha3_seq_CC12 ( clk, rst, in, out );
  input [575:0] in;
  output [1599:0] out;
  input clk, rst;
  wire   init, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
         n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
         n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
         n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
         n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877,
         n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
         n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
         n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901,
         n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
         n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917,
         n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
         n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
         n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941,
         n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
         n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
         n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965,
         n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973,
         n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
         n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
         n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
         n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
         n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013,
         n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021,
         n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
         n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037,
         n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045,
         n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
         n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
         n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
         n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
         n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085,
         n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093,
         n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
         n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
         n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117,
         n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125,
         n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133,
         n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
         n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
         n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
         n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165,
         n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173,
         n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
         n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
         n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197,
         n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
         n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213,
         n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
         n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
         n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
         n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
         n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
         n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
         n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
         n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
         n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
         n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
         n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
         n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325,
         n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
         n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
         n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
         n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
         n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
         n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
         n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
         n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
         n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
         n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
         n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
         n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
         n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
         n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
         n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
         n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
         n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
         n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
         n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
         n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
         n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
         n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
         n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
         n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
         n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
         n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
         n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
         n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
         n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
         n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
         n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
         n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
         n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
         n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
         n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
         n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
         n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
         n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
         n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
         n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
         n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
         n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
         n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
         n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
         n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
         n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
         n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
         n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
         n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069,
         n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
         n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
         n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
         n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
         n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
         n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
         n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
         n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133,
         n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
         n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
         n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
         n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165,
         n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
         n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
         n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189,
         n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
         n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205,
         n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
         n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
         n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
         n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237,
         n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245,
         n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
         n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261,
         n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
         n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277,
         n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285,
         n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293,
         n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301,
         n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309,
         n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317,
         n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325,
         n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333,
         n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341,
         n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349,
         n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357,
         n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
         n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373,
         n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
         n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389,
         n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397,
         n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405,
         n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
         n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
         n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429,
         n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
         n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445,
         n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453,
         n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461,
         n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469,
         n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477,
         n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485,
         n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493,
         n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501,
         n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509,
         n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
         n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525,
         n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533,
         n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541,
         n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549,
         n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557,
         n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565,
         n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573,
         n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
         n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589,
         n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597,
         n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605,
         n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
         n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621,
         n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629,
         n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637,
         n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645,
         n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
         n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661,
         n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
         n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677,
         n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
         n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693,
         n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701,
         n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
         n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
         n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
         n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
         n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
         n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
         n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
         n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765,
         n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
         n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
         n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789,
         n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
         n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
         n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
         n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
         n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
         n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
         n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
         n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
         n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
         n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997;
  wire   [11:0] rc_i;
  wire   [1599:0] round_reg;

  DFF init_reg ( .D(1'b1), .CLK(clk), .RST(rst), .I(1'b0), .Q(init) );
  DFF \rc_i_reg[0]  ( .D(n1038), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[0])
         );
  DFF \rc_i_reg[1]  ( .D(rc_i[0]), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[1])
         );
  DFF \rc_i_reg[2]  ( .D(rc_i[1]), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[2])
         );
  DFF \rc_i_reg[3]  ( .D(rc_i[2]), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[3])
         );
  DFF \rc_i_reg[4]  ( .D(rc_i[3]), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[4])
         );
  DFF \rc_i_reg[5]  ( .D(rc_i[4]), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[5])
         );
  DFF \rc_i_reg[6]  ( .D(rc_i[5]), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[6])
         );
  DFF \rc_i_reg[7]  ( .D(rc_i[6]), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[7])
         );
  DFF \rc_i_reg[8]  ( .D(rc_i[7]), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[8])
         );
  DFF \rc_i_reg[9]  ( .D(rc_i[8]), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[9])
         );
  DFF \rc_i_reg[10]  ( .D(rc_i[9]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        rc_i[10]) );
  DFF \rc_i_reg[11]  ( .D(rc_i[10]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        rc_i[11]) );
  DFF \round_reg_reg[0]  ( .D(out[0]), .CLK(clk), .RST(rst), .I(in[0]), .Q(
        round_reg[0]) );
  DFF \round_reg_reg[1]  ( .D(out[1]), .CLK(clk), .RST(rst), .I(in[1]), .Q(
        round_reg[1]) );
  DFF \round_reg_reg[2]  ( .D(out[2]), .CLK(clk), .RST(rst), .I(in[2]), .Q(
        round_reg[2]) );
  DFF \round_reg_reg[3]  ( .D(out[3]), .CLK(clk), .RST(rst), .I(in[3]), .Q(
        round_reg[3]) );
  DFF \round_reg_reg[4]  ( .D(out[4]), .CLK(clk), .RST(rst), .I(in[4]), .Q(
        round_reg[4]) );
  DFF \round_reg_reg[5]  ( .D(out[5]), .CLK(clk), .RST(rst), .I(in[5]), .Q(
        round_reg[5]) );
  DFF \round_reg_reg[6]  ( .D(out[6]), .CLK(clk), .RST(rst), .I(in[6]), .Q(
        round_reg[6]) );
  DFF \round_reg_reg[7]  ( .D(out[7]), .CLK(clk), .RST(rst), .I(in[7]), .Q(
        round_reg[7]) );
  DFF \round_reg_reg[8]  ( .D(out[8]), .CLK(clk), .RST(rst), .I(in[8]), .Q(
        round_reg[8]) );
  DFF \round_reg_reg[9]  ( .D(out[9]), .CLK(clk), .RST(rst), .I(in[9]), .Q(
        round_reg[9]) );
  DFF \round_reg_reg[10]  ( .D(out[10]), .CLK(clk), .RST(rst), .I(in[10]), .Q(
        round_reg[10]) );
  DFF \round_reg_reg[11]  ( .D(out[11]), .CLK(clk), .RST(rst), .I(in[11]), .Q(
        round_reg[11]) );
  DFF \round_reg_reg[12]  ( .D(out[12]), .CLK(clk), .RST(rst), .I(in[12]), .Q(
        round_reg[12]) );
  DFF \round_reg_reg[13]  ( .D(out[13]), .CLK(clk), .RST(rst), .I(in[13]), .Q(
        round_reg[13]) );
  DFF \round_reg_reg[14]  ( .D(out[14]), .CLK(clk), .RST(rst), .I(in[14]), .Q(
        round_reg[14]) );
  DFF \round_reg_reg[15]  ( .D(out[15]), .CLK(clk), .RST(rst), .I(in[15]), .Q(
        round_reg[15]) );
  DFF \round_reg_reg[16]  ( .D(out[16]), .CLK(clk), .RST(rst), .I(in[16]), .Q(
        round_reg[16]) );
  DFF \round_reg_reg[17]  ( .D(out[17]), .CLK(clk), .RST(rst), .I(in[17]), .Q(
        round_reg[17]) );
  DFF \round_reg_reg[18]  ( .D(out[18]), .CLK(clk), .RST(rst), .I(in[18]), .Q(
        round_reg[18]) );
  DFF \round_reg_reg[19]  ( .D(out[19]), .CLK(clk), .RST(rst), .I(in[19]), .Q(
        round_reg[19]) );
  DFF \round_reg_reg[20]  ( .D(out[20]), .CLK(clk), .RST(rst), .I(in[20]), .Q(
        round_reg[20]) );
  DFF \round_reg_reg[21]  ( .D(out[21]), .CLK(clk), .RST(rst), .I(in[21]), .Q(
        round_reg[21]) );
  DFF \round_reg_reg[22]  ( .D(out[22]), .CLK(clk), .RST(rst), .I(in[22]), .Q(
        round_reg[22]) );
  DFF \round_reg_reg[23]  ( .D(out[23]), .CLK(clk), .RST(rst), .I(in[23]), .Q(
        round_reg[23]) );
  DFF \round_reg_reg[24]  ( .D(out[24]), .CLK(clk), .RST(rst), .I(in[24]), .Q(
        round_reg[24]) );
  DFF \round_reg_reg[25]  ( .D(out[25]), .CLK(clk), .RST(rst), .I(in[25]), .Q(
        round_reg[25]) );
  DFF \round_reg_reg[26]  ( .D(out[26]), .CLK(clk), .RST(rst), .I(in[26]), .Q(
        round_reg[26]) );
  DFF \round_reg_reg[27]  ( .D(out[27]), .CLK(clk), .RST(rst), .I(in[27]), .Q(
        round_reg[27]) );
  DFF \round_reg_reg[28]  ( .D(out[28]), .CLK(clk), .RST(rst), .I(in[28]), .Q(
        round_reg[28]) );
  DFF \round_reg_reg[29]  ( .D(out[29]), .CLK(clk), .RST(rst), .I(in[29]), .Q(
        round_reg[29]) );
  DFF \round_reg_reg[30]  ( .D(out[30]), .CLK(clk), .RST(rst), .I(in[30]), .Q(
        round_reg[30]) );
  DFF \round_reg_reg[31]  ( .D(out[31]), .CLK(clk), .RST(rst), .I(in[31]), .Q(
        round_reg[31]) );
  DFF \round_reg_reg[32]  ( .D(out[32]), .CLK(clk), .RST(rst), .I(in[32]), .Q(
        round_reg[32]) );
  DFF \round_reg_reg[33]  ( .D(out[33]), .CLK(clk), .RST(rst), .I(in[33]), .Q(
        round_reg[33]) );
  DFF \round_reg_reg[34]  ( .D(out[34]), .CLK(clk), .RST(rst), .I(in[34]), .Q(
        round_reg[34]) );
  DFF \round_reg_reg[35]  ( .D(out[35]), .CLK(clk), .RST(rst), .I(in[35]), .Q(
        round_reg[35]) );
  DFF \round_reg_reg[36]  ( .D(out[36]), .CLK(clk), .RST(rst), .I(in[36]), .Q(
        round_reg[36]) );
  DFF \round_reg_reg[37]  ( .D(out[37]), .CLK(clk), .RST(rst), .I(in[37]), .Q(
        round_reg[37]) );
  DFF \round_reg_reg[38]  ( .D(out[38]), .CLK(clk), .RST(rst), .I(in[38]), .Q(
        round_reg[38]) );
  DFF \round_reg_reg[39]  ( .D(out[39]), .CLK(clk), .RST(rst), .I(in[39]), .Q(
        round_reg[39]) );
  DFF \round_reg_reg[40]  ( .D(out[40]), .CLK(clk), .RST(rst), .I(in[40]), .Q(
        round_reg[40]) );
  DFF \round_reg_reg[41]  ( .D(out[41]), .CLK(clk), .RST(rst), .I(in[41]), .Q(
        round_reg[41]) );
  DFF \round_reg_reg[42]  ( .D(out[42]), .CLK(clk), .RST(rst), .I(in[42]), .Q(
        round_reg[42]) );
  DFF \round_reg_reg[43]  ( .D(out[43]), .CLK(clk), .RST(rst), .I(in[43]), .Q(
        round_reg[43]) );
  DFF \round_reg_reg[44]  ( .D(out[44]), .CLK(clk), .RST(rst), .I(in[44]), .Q(
        round_reg[44]) );
  DFF \round_reg_reg[45]  ( .D(out[45]), .CLK(clk), .RST(rst), .I(in[45]), .Q(
        round_reg[45]) );
  DFF \round_reg_reg[46]  ( .D(out[46]), .CLK(clk), .RST(rst), .I(in[46]), .Q(
        round_reg[46]) );
  DFF \round_reg_reg[47]  ( .D(out[47]), .CLK(clk), .RST(rst), .I(in[47]), .Q(
        round_reg[47]) );
  DFF \round_reg_reg[48]  ( .D(out[48]), .CLK(clk), .RST(rst), .I(in[48]), .Q(
        round_reg[48]) );
  DFF \round_reg_reg[49]  ( .D(out[49]), .CLK(clk), .RST(rst), .I(in[49]), .Q(
        round_reg[49]) );
  DFF \round_reg_reg[50]  ( .D(out[50]), .CLK(clk), .RST(rst), .I(in[50]), .Q(
        round_reg[50]) );
  DFF \round_reg_reg[51]  ( .D(out[51]), .CLK(clk), .RST(rst), .I(in[51]), .Q(
        round_reg[51]) );
  DFF \round_reg_reg[52]  ( .D(out[52]), .CLK(clk), .RST(rst), .I(in[52]), .Q(
        round_reg[52]) );
  DFF \round_reg_reg[53]  ( .D(out[53]), .CLK(clk), .RST(rst), .I(in[53]), .Q(
        round_reg[53]) );
  DFF \round_reg_reg[54]  ( .D(out[54]), .CLK(clk), .RST(rst), .I(in[54]), .Q(
        round_reg[54]) );
  DFF \round_reg_reg[55]  ( .D(out[55]), .CLK(clk), .RST(rst), .I(in[55]), .Q(
        round_reg[55]) );
  DFF \round_reg_reg[56]  ( .D(out[56]), .CLK(clk), .RST(rst), .I(in[56]), .Q(
        round_reg[56]) );
  DFF \round_reg_reg[57]  ( .D(out[57]), .CLK(clk), .RST(rst), .I(in[57]), .Q(
        round_reg[57]) );
  DFF \round_reg_reg[58]  ( .D(out[58]), .CLK(clk), .RST(rst), .I(in[58]), .Q(
        round_reg[58]) );
  DFF \round_reg_reg[59]  ( .D(out[59]), .CLK(clk), .RST(rst), .I(in[59]), .Q(
        round_reg[59]) );
  DFF \round_reg_reg[60]  ( .D(out[60]), .CLK(clk), .RST(rst), .I(in[60]), .Q(
        round_reg[60]) );
  DFF \round_reg_reg[61]  ( .D(out[61]), .CLK(clk), .RST(rst), .I(in[61]), .Q(
        round_reg[61]) );
  DFF \round_reg_reg[62]  ( .D(out[62]), .CLK(clk), .RST(rst), .I(in[62]), .Q(
        round_reg[62]) );
  DFF \round_reg_reg[63]  ( .D(out[63]), .CLK(clk), .RST(rst), .I(in[63]), .Q(
        round_reg[63]) );
  DFF \round_reg_reg[64]  ( .D(out[64]), .CLK(clk), .RST(rst), .I(in[64]), .Q(
        round_reg[64]) );
  DFF \round_reg_reg[65]  ( .D(out[65]), .CLK(clk), .RST(rst), .I(in[65]), .Q(
        round_reg[65]) );
  DFF \round_reg_reg[66]  ( .D(out[66]), .CLK(clk), .RST(rst), .I(in[66]), .Q(
        round_reg[66]) );
  DFF \round_reg_reg[67]  ( .D(out[67]), .CLK(clk), .RST(rst), .I(in[67]), .Q(
        round_reg[67]) );
  DFF \round_reg_reg[68]  ( .D(out[68]), .CLK(clk), .RST(rst), .I(in[68]), .Q(
        round_reg[68]) );
  DFF \round_reg_reg[69]  ( .D(out[69]), .CLK(clk), .RST(rst), .I(in[69]), .Q(
        round_reg[69]) );
  DFF \round_reg_reg[70]  ( .D(out[70]), .CLK(clk), .RST(rst), .I(in[70]), .Q(
        round_reg[70]) );
  DFF \round_reg_reg[71]  ( .D(out[71]), .CLK(clk), .RST(rst), .I(in[71]), .Q(
        round_reg[71]) );
  DFF \round_reg_reg[72]  ( .D(out[72]), .CLK(clk), .RST(rst), .I(in[72]), .Q(
        round_reg[72]) );
  DFF \round_reg_reg[73]  ( .D(out[73]), .CLK(clk), .RST(rst), .I(in[73]), .Q(
        round_reg[73]) );
  DFF \round_reg_reg[74]  ( .D(out[74]), .CLK(clk), .RST(rst), .I(in[74]), .Q(
        round_reg[74]) );
  DFF \round_reg_reg[75]  ( .D(out[75]), .CLK(clk), .RST(rst), .I(in[75]), .Q(
        round_reg[75]) );
  DFF \round_reg_reg[76]  ( .D(out[76]), .CLK(clk), .RST(rst), .I(in[76]), .Q(
        round_reg[76]) );
  DFF \round_reg_reg[77]  ( .D(out[77]), .CLK(clk), .RST(rst), .I(in[77]), .Q(
        round_reg[77]) );
  DFF \round_reg_reg[78]  ( .D(out[78]), .CLK(clk), .RST(rst), .I(in[78]), .Q(
        round_reg[78]) );
  DFF \round_reg_reg[79]  ( .D(out[79]), .CLK(clk), .RST(rst), .I(in[79]), .Q(
        round_reg[79]) );
  DFF \round_reg_reg[80]  ( .D(out[80]), .CLK(clk), .RST(rst), .I(in[80]), .Q(
        round_reg[80]) );
  DFF \round_reg_reg[81]  ( .D(out[81]), .CLK(clk), .RST(rst), .I(in[81]), .Q(
        round_reg[81]) );
  DFF \round_reg_reg[82]  ( .D(out[82]), .CLK(clk), .RST(rst), .I(in[82]), .Q(
        round_reg[82]) );
  DFF \round_reg_reg[83]  ( .D(out[83]), .CLK(clk), .RST(rst), .I(in[83]), .Q(
        round_reg[83]) );
  DFF \round_reg_reg[84]  ( .D(out[84]), .CLK(clk), .RST(rst), .I(in[84]), .Q(
        round_reg[84]) );
  DFF \round_reg_reg[85]  ( .D(out[85]), .CLK(clk), .RST(rst), .I(in[85]), .Q(
        round_reg[85]) );
  DFF \round_reg_reg[86]  ( .D(out[86]), .CLK(clk), .RST(rst), .I(in[86]), .Q(
        round_reg[86]) );
  DFF \round_reg_reg[87]  ( .D(out[87]), .CLK(clk), .RST(rst), .I(in[87]), .Q(
        round_reg[87]) );
  DFF \round_reg_reg[88]  ( .D(out[88]), .CLK(clk), .RST(rst), .I(in[88]), .Q(
        round_reg[88]) );
  DFF \round_reg_reg[89]  ( .D(out[89]), .CLK(clk), .RST(rst), .I(in[89]), .Q(
        round_reg[89]) );
  DFF \round_reg_reg[90]  ( .D(out[90]), .CLK(clk), .RST(rst), .I(in[90]), .Q(
        round_reg[90]) );
  DFF \round_reg_reg[91]  ( .D(out[91]), .CLK(clk), .RST(rst), .I(in[91]), .Q(
        round_reg[91]) );
  DFF \round_reg_reg[92]  ( .D(out[92]), .CLK(clk), .RST(rst), .I(in[92]), .Q(
        round_reg[92]) );
  DFF \round_reg_reg[93]  ( .D(out[93]), .CLK(clk), .RST(rst), .I(in[93]), .Q(
        round_reg[93]) );
  DFF \round_reg_reg[94]  ( .D(out[94]), .CLK(clk), .RST(rst), .I(in[94]), .Q(
        round_reg[94]) );
  DFF \round_reg_reg[95]  ( .D(out[95]), .CLK(clk), .RST(rst), .I(in[95]), .Q(
        round_reg[95]) );
  DFF \round_reg_reg[96]  ( .D(out[96]), .CLK(clk), .RST(rst), .I(in[96]), .Q(
        round_reg[96]) );
  DFF \round_reg_reg[97]  ( .D(out[97]), .CLK(clk), .RST(rst), .I(in[97]), .Q(
        round_reg[97]) );
  DFF \round_reg_reg[98]  ( .D(out[98]), .CLK(clk), .RST(rst), .I(in[98]), .Q(
        round_reg[98]) );
  DFF \round_reg_reg[99]  ( .D(out[99]), .CLK(clk), .RST(rst), .I(in[99]), .Q(
        round_reg[99]) );
  DFF \round_reg_reg[100]  ( .D(out[100]), .CLK(clk), .RST(rst), .I(in[100]), 
        .Q(round_reg[100]) );
  DFF \round_reg_reg[101]  ( .D(out[101]), .CLK(clk), .RST(rst), .I(in[101]), 
        .Q(round_reg[101]) );
  DFF \round_reg_reg[102]  ( .D(out[102]), .CLK(clk), .RST(rst), .I(in[102]), 
        .Q(round_reg[102]) );
  DFF \round_reg_reg[103]  ( .D(out[103]), .CLK(clk), .RST(rst), .I(in[103]), 
        .Q(round_reg[103]) );
  DFF \round_reg_reg[104]  ( .D(out[104]), .CLK(clk), .RST(rst), .I(in[104]), 
        .Q(round_reg[104]) );
  DFF \round_reg_reg[105]  ( .D(out[105]), .CLK(clk), .RST(rst), .I(in[105]), 
        .Q(round_reg[105]) );
  DFF \round_reg_reg[106]  ( .D(out[106]), .CLK(clk), .RST(rst), .I(in[106]), 
        .Q(round_reg[106]) );
  DFF \round_reg_reg[107]  ( .D(out[107]), .CLK(clk), .RST(rst), .I(in[107]), 
        .Q(round_reg[107]) );
  DFF \round_reg_reg[108]  ( .D(out[108]), .CLK(clk), .RST(rst), .I(in[108]), 
        .Q(round_reg[108]) );
  DFF \round_reg_reg[109]  ( .D(out[109]), .CLK(clk), .RST(rst), .I(in[109]), 
        .Q(round_reg[109]) );
  DFF \round_reg_reg[110]  ( .D(out[110]), .CLK(clk), .RST(rst), .I(in[110]), 
        .Q(round_reg[110]) );
  DFF \round_reg_reg[111]  ( .D(out[111]), .CLK(clk), .RST(rst), .I(in[111]), 
        .Q(round_reg[111]) );
  DFF \round_reg_reg[112]  ( .D(out[112]), .CLK(clk), .RST(rst), .I(in[112]), 
        .Q(round_reg[112]) );
  DFF \round_reg_reg[113]  ( .D(out[113]), .CLK(clk), .RST(rst), .I(in[113]), 
        .Q(round_reg[113]) );
  DFF \round_reg_reg[114]  ( .D(out[114]), .CLK(clk), .RST(rst), .I(in[114]), 
        .Q(round_reg[114]) );
  DFF \round_reg_reg[115]  ( .D(out[115]), .CLK(clk), .RST(rst), .I(in[115]), 
        .Q(round_reg[115]) );
  DFF \round_reg_reg[116]  ( .D(out[116]), .CLK(clk), .RST(rst), .I(in[116]), 
        .Q(round_reg[116]) );
  DFF \round_reg_reg[117]  ( .D(out[117]), .CLK(clk), .RST(rst), .I(in[117]), 
        .Q(round_reg[117]) );
  DFF \round_reg_reg[118]  ( .D(out[118]), .CLK(clk), .RST(rst), .I(in[118]), 
        .Q(round_reg[118]) );
  DFF \round_reg_reg[119]  ( .D(out[119]), .CLK(clk), .RST(rst), .I(in[119]), 
        .Q(round_reg[119]) );
  DFF \round_reg_reg[120]  ( .D(out[120]), .CLK(clk), .RST(rst), .I(in[120]), 
        .Q(round_reg[120]) );
  DFF \round_reg_reg[121]  ( .D(out[121]), .CLK(clk), .RST(rst), .I(in[121]), 
        .Q(round_reg[121]) );
  DFF \round_reg_reg[122]  ( .D(out[122]), .CLK(clk), .RST(rst), .I(in[122]), 
        .Q(round_reg[122]) );
  DFF \round_reg_reg[123]  ( .D(out[123]), .CLK(clk), .RST(rst), .I(in[123]), 
        .Q(round_reg[123]) );
  DFF \round_reg_reg[124]  ( .D(out[124]), .CLK(clk), .RST(rst), .I(in[124]), 
        .Q(round_reg[124]) );
  DFF \round_reg_reg[125]  ( .D(out[125]), .CLK(clk), .RST(rst), .I(in[125]), 
        .Q(round_reg[125]) );
  DFF \round_reg_reg[126]  ( .D(out[126]), .CLK(clk), .RST(rst), .I(in[126]), 
        .Q(round_reg[126]) );
  DFF \round_reg_reg[127]  ( .D(out[127]), .CLK(clk), .RST(rst), .I(in[127]), 
        .Q(round_reg[127]) );
  DFF \round_reg_reg[128]  ( .D(out[128]), .CLK(clk), .RST(rst), .I(in[128]), 
        .Q(round_reg[128]) );
  DFF \round_reg_reg[129]  ( .D(out[129]), .CLK(clk), .RST(rst), .I(in[129]), 
        .Q(round_reg[129]) );
  DFF \round_reg_reg[130]  ( .D(out[130]), .CLK(clk), .RST(rst), .I(in[130]), 
        .Q(round_reg[130]) );
  DFF \round_reg_reg[131]  ( .D(out[131]), .CLK(clk), .RST(rst), .I(in[131]), 
        .Q(round_reg[131]) );
  DFF \round_reg_reg[132]  ( .D(out[132]), .CLK(clk), .RST(rst), .I(in[132]), 
        .Q(round_reg[132]) );
  DFF \round_reg_reg[133]  ( .D(out[133]), .CLK(clk), .RST(rst), .I(in[133]), 
        .Q(round_reg[133]) );
  DFF \round_reg_reg[134]  ( .D(out[134]), .CLK(clk), .RST(rst), .I(in[134]), 
        .Q(round_reg[134]) );
  DFF \round_reg_reg[135]  ( .D(out[135]), .CLK(clk), .RST(rst), .I(in[135]), 
        .Q(round_reg[135]) );
  DFF \round_reg_reg[136]  ( .D(out[136]), .CLK(clk), .RST(rst), .I(in[136]), 
        .Q(round_reg[136]) );
  DFF \round_reg_reg[137]  ( .D(out[137]), .CLK(clk), .RST(rst), .I(in[137]), 
        .Q(round_reg[137]) );
  DFF \round_reg_reg[138]  ( .D(out[138]), .CLK(clk), .RST(rst), .I(in[138]), 
        .Q(round_reg[138]) );
  DFF \round_reg_reg[139]  ( .D(out[139]), .CLK(clk), .RST(rst), .I(in[139]), 
        .Q(round_reg[139]) );
  DFF \round_reg_reg[140]  ( .D(out[140]), .CLK(clk), .RST(rst), .I(in[140]), 
        .Q(round_reg[140]) );
  DFF \round_reg_reg[141]  ( .D(out[141]), .CLK(clk), .RST(rst), .I(in[141]), 
        .Q(round_reg[141]) );
  DFF \round_reg_reg[142]  ( .D(out[142]), .CLK(clk), .RST(rst), .I(in[142]), 
        .Q(round_reg[142]) );
  DFF \round_reg_reg[143]  ( .D(out[143]), .CLK(clk), .RST(rst), .I(in[143]), 
        .Q(round_reg[143]) );
  DFF \round_reg_reg[144]  ( .D(out[144]), .CLK(clk), .RST(rst), .I(in[144]), 
        .Q(round_reg[144]) );
  DFF \round_reg_reg[145]  ( .D(out[145]), .CLK(clk), .RST(rst), .I(in[145]), 
        .Q(round_reg[145]) );
  DFF \round_reg_reg[146]  ( .D(out[146]), .CLK(clk), .RST(rst), .I(in[146]), 
        .Q(round_reg[146]) );
  DFF \round_reg_reg[147]  ( .D(out[147]), .CLK(clk), .RST(rst), .I(in[147]), 
        .Q(round_reg[147]) );
  DFF \round_reg_reg[148]  ( .D(out[148]), .CLK(clk), .RST(rst), .I(in[148]), 
        .Q(round_reg[148]) );
  DFF \round_reg_reg[149]  ( .D(out[149]), .CLK(clk), .RST(rst), .I(in[149]), 
        .Q(round_reg[149]) );
  DFF \round_reg_reg[150]  ( .D(out[150]), .CLK(clk), .RST(rst), .I(in[150]), 
        .Q(round_reg[150]) );
  DFF \round_reg_reg[151]  ( .D(out[151]), .CLK(clk), .RST(rst), .I(in[151]), 
        .Q(round_reg[151]) );
  DFF \round_reg_reg[152]  ( .D(out[152]), .CLK(clk), .RST(rst), .I(in[152]), 
        .Q(round_reg[152]) );
  DFF \round_reg_reg[153]  ( .D(out[153]), .CLK(clk), .RST(rst), .I(in[153]), 
        .Q(round_reg[153]) );
  DFF \round_reg_reg[154]  ( .D(out[154]), .CLK(clk), .RST(rst), .I(in[154]), 
        .Q(round_reg[154]) );
  DFF \round_reg_reg[155]  ( .D(out[155]), .CLK(clk), .RST(rst), .I(in[155]), 
        .Q(round_reg[155]) );
  DFF \round_reg_reg[156]  ( .D(out[156]), .CLK(clk), .RST(rst), .I(in[156]), 
        .Q(round_reg[156]) );
  DFF \round_reg_reg[157]  ( .D(out[157]), .CLK(clk), .RST(rst), .I(in[157]), 
        .Q(round_reg[157]) );
  DFF \round_reg_reg[158]  ( .D(out[158]), .CLK(clk), .RST(rst), .I(in[158]), 
        .Q(round_reg[158]) );
  DFF \round_reg_reg[159]  ( .D(out[159]), .CLK(clk), .RST(rst), .I(in[159]), 
        .Q(round_reg[159]) );
  DFF \round_reg_reg[160]  ( .D(out[160]), .CLK(clk), .RST(rst), .I(in[160]), 
        .Q(round_reg[160]) );
  DFF \round_reg_reg[161]  ( .D(out[161]), .CLK(clk), .RST(rst), .I(in[161]), 
        .Q(round_reg[161]) );
  DFF \round_reg_reg[162]  ( .D(out[162]), .CLK(clk), .RST(rst), .I(in[162]), 
        .Q(round_reg[162]) );
  DFF \round_reg_reg[163]  ( .D(out[163]), .CLK(clk), .RST(rst), .I(in[163]), 
        .Q(round_reg[163]) );
  DFF \round_reg_reg[164]  ( .D(out[164]), .CLK(clk), .RST(rst), .I(in[164]), 
        .Q(round_reg[164]) );
  DFF \round_reg_reg[165]  ( .D(out[165]), .CLK(clk), .RST(rst), .I(in[165]), 
        .Q(round_reg[165]) );
  DFF \round_reg_reg[166]  ( .D(out[166]), .CLK(clk), .RST(rst), .I(in[166]), 
        .Q(round_reg[166]) );
  DFF \round_reg_reg[167]  ( .D(out[167]), .CLK(clk), .RST(rst), .I(in[167]), 
        .Q(round_reg[167]) );
  DFF \round_reg_reg[168]  ( .D(out[168]), .CLK(clk), .RST(rst), .I(in[168]), 
        .Q(round_reg[168]) );
  DFF \round_reg_reg[169]  ( .D(out[169]), .CLK(clk), .RST(rst), .I(in[169]), 
        .Q(round_reg[169]) );
  DFF \round_reg_reg[170]  ( .D(out[170]), .CLK(clk), .RST(rst), .I(in[170]), 
        .Q(round_reg[170]) );
  DFF \round_reg_reg[171]  ( .D(out[171]), .CLK(clk), .RST(rst), .I(in[171]), 
        .Q(round_reg[171]) );
  DFF \round_reg_reg[172]  ( .D(out[172]), .CLK(clk), .RST(rst), .I(in[172]), 
        .Q(round_reg[172]) );
  DFF \round_reg_reg[173]  ( .D(out[173]), .CLK(clk), .RST(rst), .I(in[173]), 
        .Q(round_reg[173]) );
  DFF \round_reg_reg[174]  ( .D(out[174]), .CLK(clk), .RST(rst), .I(in[174]), 
        .Q(round_reg[174]) );
  DFF \round_reg_reg[175]  ( .D(out[175]), .CLK(clk), .RST(rst), .I(in[175]), 
        .Q(round_reg[175]) );
  DFF \round_reg_reg[176]  ( .D(out[176]), .CLK(clk), .RST(rst), .I(in[176]), 
        .Q(round_reg[176]) );
  DFF \round_reg_reg[177]  ( .D(out[177]), .CLK(clk), .RST(rst), .I(in[177]), 
        .Q(round_reg[177]) );
  DFF \round_reg_reg[178]  ( .D(out[178]), .CLK(clk), .RST(rst), .I(in[178]), 
        .Q(round_reg[178]) );
  DFF \round_reg_reg[179]  ( .D(out[179]), .CLK(clk), .RST(rst), .I(in[179]), 
        .Q(round_reg[179]) );
  DFF \round_reg_reg[180]  ( .D(out[180]), .CLK(clk), .RST(rst), .I(in[180]), 
        .Q(round_reg[180]) );
  DFF \round_reg_reg[181]  ( .D(out[181]), .CLK(clk), .RST(rst), .I(in[181]), 
        .Q(round_reg[181]) );
  DFF \round_reg_reg[182]  ( .D(out[182]), .CLK(clk), .RST(rst), .I(in[182]), 
        .Q(round_reg[182]) );
  DFF \round_reg_reg[183]  ( .D(out[183]), .CLK(clk), .RST(rst), .I(in[183]), 
        .Q(round_reg[183]) );
  DFF \round_reg_reg[184]  ( .D(out[184]), .CLK(clk), .RST(rst), .I(in[184]), 
        .Q(round_reg[184]) );
  DFF \round_reg_reg[185]  ( .D(out[185]), .CLK(clk), .RST(rst), .I(in[185]), 
        .Q(round_reg[185]) );
  DFF \round_reg_reg[186]  ( .D(out[186]), .CLK(clk), .RST(rst), .I(in[186]), 
        .Q(round_reg[186]) );
  DFF \round_reg_reg[187]  ( .D(out[187]), .CLK(clk), .RST(rst), .I(in[187]), 
        .Q(round_reg[187]) );
  DFF \round_reg_reg[188]  ( .D(out[188]), .CLK(clk), .RST(rst), .I(in[188]), 
        .Q(round_reg[188]) );
  DFF \round_reg_reg[189]  ( .D(out[189]), .CLK(clk), .RST(rst), .I(in[189]), 
        .Q(round_reg[189]) );
  DFF \round_reg_reg[190]  ( .D(out[190]), .CLK(clk), .RST(rst), .I(in[190]), 
        .Q(round_reg[190]) );
  DFF \round_reg_reg[191]  ( .D(out[191]), .CLK(clk), .RST(rst), .I(in[191]), 
        .Q(round_reg[191]) );
  DFF \round_reg_reg[192]  ( .D(out[192]), .CLK(clk), .RST(rst), .I(in[192]), 
        .Q(round_reg[192]) );
  DFF \round_reg_reg[193]  ( .D(out[193]), .CLK(clk), .RST(rst), .I(in[193]), 
        .Q(round_reg[193]) );
  DFF \round_reg_reg[194]  ( .D(out[194]), .CLK(clk), .RST(rst), .I(in[194]), 
        .Q(round_reg[194]) );
  DFF \round_reg_reg[195]  ( .D(out[195]), .CLK(clk), .RST(rst), .I(in[195]), 
        .Q(round_reg[195]) );
  DFF \round_reg_reg[196]  ( .D(out[196]), .CLK(clk), .RST(rst), .I(in[196]), 
        .Q(round_reg[196]) );
  DFF \round_reg_reg[197]  ( .D(out[197]), .CLK(clk), .RST(rst), .I(in[197]), 
        .Q(round_reg[197]) );
  DFF \round_reg_reg[198]  ( .D(out[198]), .CLK(clk), .RST(rst), .I(in[198]), 
        .Q(round_reg[198]) );
  DFF \round_reg_reg[199]  ( .D(out[199]), .CLK(clk), .RST(rst), .I(in[199]), 
        .Q(round_reg[199]) );
  DFF \round_reg_reg[200]  ( .D(out[200]), .CLK(clk), .RST(rst), .I(in[200]), 
        .Q(round_reg[200]) );
  DFF \round_reg_reg[201]  ( .D(out[201]), .CLK(clk), .RST(rst), .I(in[201]), 
        .Q(round_reg[201]) );
  DFF \round_reg_reg[202]  ( .D(out[202]), .CLK(clk), .RST(rst), .I(in[202]), 
        .Q(round_reg[202]) );
  DFF \round_reg_reg[203]  ( .D(out[203]), .CLK(clk), .RST(rst), .I(in[203]), 
        .Q(round_reg[203]) );
  DFF \round_reg_reg[204]  ( .D(out[204]), .CLK(clk), .RST(rst), .I(in[204]), 
        .Q(round_reg[204]) );
  DFF \round_reg_reg[205]  ( .D(out[205]), .CLK(clk), .RST(rst), .I(in[205]), 
        .Q(round_reg[205]) );
  DFF \round_reg_reg[206]  ( .D(out[206]), .CLK(clk), .RST(rst), .I(in[206]), 
        .Q(round_reg[206]) );
  DFF \round_reg_reg[207]  ( .D(out[207]), .CLK(clk), .RST(rst), .I(in[207]), 
        .Q(round_reg[207]) );
  DFF \round_reg_reg[208]  ( .D(out[208]), .CLK(clk), .RST(rst), .I(in[208]), 
        .Q(round_reg[208]) );
  DFF \round_reg_reg[209]  ( .D(out[209]), .CLK(clk), .RST(rst), .I(in[209]), 
        .Q(round_reg[209]) );
  DFF \round_reg_reg[210]  ( .D(out[210]), .CLK(clk), .RST(rst), .I(in[210]), 
        .Q(round_reg[210]) );
  DFF \round_reg_reg[211]  ( .D(out[211]), .CLK(clk), .RST(rst), .I(in[211]), 
        .Q(round_reg[211]) );
  DFF \round_reg_reg[212]  ( .D(out[212]), .CLK(clk), .RST(rst), .I(in[212]), 
        .Q(round_reg[212]) );
  DFF \round_reg_reg[213]  ( .D(out[213]), .CLK(clk), .RST(rst), .I(in[213]), 
        .Q(round_reg[213]) );
  DFF \round_reg_reg[214]  ( .D(out[214]), .CLK(clk), .RST(rst), .I(in[214]), 
        .Q(round_reg[214]) );
  DFF \round_reg_reg[215]  ( .D(out[215]), .CLK(clk), .RST(rst), .I(in[215]), 
        .Q(round_reg[215]) );
  DFF \round_reg_reg[216]  ( .D(out[216]), .CLK(clk), .RST(rst), .I(in[216]), 
        .Q(round_reg[216]) );
  DFF \round_reg_reg[217]  ( .D(out[217]), .CLK(clk), .RST(rst), .I(in[217]), 
        .Q(round_reg[217]) );
  DFF \round_reg_reg[218]  ( .D(out[218]), .CLK(clk), .RST(rst), .I(in[218]), 
        .Q(round_reg[218]) );
  DFF \round_reg_reg[219]  ( .D(out[219]), .CLK(clk), .RST(rst), .I(in[219]), 
        .Q(round_reg[219]) );
  DFF \round_reg_reg[220]  ( .D(out[220]), .CLK(clk), .RST(rst), .I(in[220]), 
        .Q(round_reg[220]) );
  DFF \round_reg_reg[221]  ( .D(out[221]), .CLK(clk), .RST(rst), .I(in[221]), 
        .Q(round_reg[221]) );
  DFF \round_reg_reg[222]  ( .D(out[222]), .CLK(clk), .RST(rst), .I(in[222]), 
        .Q(round_reg[222]) );
  DFF \round_reg_reg[223]  ( .D(out[223]), .CLK(clk), .RST(rst), .I(in[223]), 
        .Q(round_reg[223]) );
  DFF \round_reg_reg[224]  ( .D(out[224]), .CLK(clk), .RST(rst), .I(in[224]), 
        .Q(round_reg[224]) );
  DFF \round_reg_reg[225]  ( .D(out[225]), .CLK(clk), .RST(rst), .I(in[225]), 
        .Q(round_reg[225]) );
  DFF \round_reg_reg[226]  ( .D(out[226]), .CLK(clk), .RST(rst), .I(in[226]), 
        .Q(round_reg[226]) );
  DFF \round_reg_reg[227]  ( .D(out[227]), .CLK(clk), .RST(rst), .I(in[227]), 
        .Q(round_reg[227]) );
  DFF \round_reg_reg[228]  ( .D(out[228]), .CLK(clk), .RST(rst), .I(in[228]), 
        .Q(round_reg[228]) );
  DFF \round_reg_reg[229]  ( .D(out[229]), .CLK(clk), .RST(rst), .I(in[229]), 
        .Q(round_reg[229]) );
  DFF \round_reg_reg[230]  ( .D(out[230]), .CLK(clk), .RST(rst), .I(in[230]), 
        .Q(round_reg[230]) );
  DFF \round_reg_reg[231]  ( .D(out[231]), .CLK(clk), .RST(rst), .I(in[231]), 
        .Q(round_reg[231]) );
  DFF \round_reg_reg[232]  ( .D(out[232]), .CLK(clk), .RST(rst), .I(in[232]), 
        .Q(round_reg[232]) );
  DFF \round_reg_reg[233]  ( .D(out[233]), .CLK(clk), .RST(rst), .I(in[233]), 
        .Q(round_reg[233]) );
  DFF \round_reg_reg[234]  ( .D(out[234]), .CLK(clk), .RST(rst), .I(in[234]), 
        .Q(round_reg[234]) );
  DFF \round_reg_reg[235]  ( .D(out[235]), .CLK(clk), .RST(rst), .I(in[235]), 
        .Q(round_reg[235]) );
  DFF \round_reg_reg[236]  ( .D(out[236]), .CLK(clk), .RST(rst), .I(in[236]), 
        .Q(round_reg[236]) );
  DFF \round_reg_reg[237]  ( .D(out[237]), .CLK(clk), .RST(rst), .I(in[237]), 
        .Q(round_reg[237]) );
  DFF \round_reg_reg[238]  ( .D(out[238]), .CLK(clk), .RST(rst), .I(in[238]), 
        .Q(round_reg[238]) );
  DFF \round_reg_reg[239]  ( .D(out[239]), .CLK(clk), .RST(rst), .I(in[239]), 
        .Q(round_reg[239]) );
  DFF \round_reg_reg[240]  ( .D(out[240]), .CLK(clk), .RST(rst), .I(in[240]), 
        .Q(round_reg[240]) );
  DFF \round_reg_reg[241]  ( .D(out[241]), .CLK(clk), .RST(rst), .I(in[241]), 
        .Q(round_reg[241]) );
  DFF \round_reg_reg[242]  ( .D(out[242]), .CLK(clk), .RST(rst), .I(in[242]), 
        .Q(round_reg[242]) );
  DFF \round_reg_reg[243]  ( .D(out[243]), .CLK(clk), .RST(rst), .I(in[243]), 
        .Q(round_reg[243]) );
  DFF \round_reg_reg[244]  ( .D(out[244]), .CLK(clk), .RST(rst), .I(in[244]), 
        .Q(round_reg[244]) );
  DFF \round_reg_reg[245]  ( .D(out[245]), .CLK(clk), .RST(rst), .I(in[245]), 
        .Q(round_reg[245]) );
  DFF \round_reg_reg[246]  ( .D(out[246]), .CLK(clk), .RST(rst), .I(in[246]), 
        .Q(round_reg[246]) );
  DFF \round_reg_reg[247]  ( .D(out[247]), .CLK(clk), .RST(rst), .I(in[247]), 
        .Q(round_reg[247]) );
  DFF \round_reg_reg[248]  ( .D(out[248]), .CLK(clk), .RST(rst), .I(in[248]), 
        .Q(round_reg[248]) );
  DFF \round_reg_reg[249]  ( .D(out[249]), .CLK(clk), .RST(rst), .I(in[249]), 
        .Q(round_reg[249]) );
  DFF \round_reg_reg[250]  ( .D(out[250]), .CLK(clk), .RST(rst), .I(in[250]), 
        .Q(round_reg[250]) );
  DFF \round_reg_reg[251]  ( .D(out[251]), .CLK(clk), .RST(rst), .I(in[251]), 
        .Q(round_reg[251]) );
  DFF \round_reg_reg[252]  ( .D(out[252]), .CLK(clk), .RST(rst), .I(in[252]), 
        .Q(round_reg[252]) );
  DFF \round_reg_reg[253]  ( .D(out[253]), .CLK(clk), .RST(rst), .I(in[253]), 
        .Q(round_reg[253]) );
  DFF \round_reg_reg[254]  ( .D(out[254]), .CLK(clk), .RST(rst), .I(in[254]), 
        .Q(round_reg[254]) );
  DFF \round_reg_reg[255]  ( .D(out[255]), .CLK(clk), .RST(rst), .I(in[255]), 
        .Q(round_reg[255]) );
  DFF \round_reg_reg[256]  ( .D(out[256]), .CLK(clk), .RST(rst), .I(in[256]), 
        .Q(round_reg[256]) );
  DFF \round_reg_reg[257]  ( .D(out[257]), .CLK(clk), .RST(rst), .I(in[257]), 
        .Q(round_reg[257]) );
  DFF \round_reg_reg[258]  ( .D(out[258]), .CLK(clk), .RST(rst), .I(in[258]), 
        .Q(round_reg[258]) );
  DFF \round_reg_reg[259]  ( .D(out[259]), .CLK(clk), .RST(rst), .I(in[259]), 
        .Q(round_reg[259]) );
  DFF \round_reg_reg[260]  ( .D(out[260]), .CLK(clk), .RST(rst), .I(in[260]), 
        .Q(round_reg[260]) );
  DFF \round_reg_reg[261]  ( .D(out[261]), .CLK(clk), .RST(rst), .I(in[261]), 
        .Q(round_reg[261]) );
  DFF \round_reg_reg[262]  ( .D(out[262]), .CLK(clk), .RST(rst), .I(in[262]), 
        .Q(round_reg[262]) );
  DFF \round_reg_reg[263]  ( .D(out[263]), .CLK(clk), .RST(rst), .I(in[263]), 
        .Q(round_reg[263]) );
  DFF \round_reg_reg[264]  ( .D(out[264]), .CLK(clk), .RST(rst), .I(in[264]), 
        .Q(round_reg[264]) );
  DFF \round_reg_reg[265]  ( .D(out[265]), .CLK(clk), .RST(rst), .I(in[265]), 
        .Q(round_reg[265]) );
  DFF \round_reg_reg[266]  ( .D(out[266]), .CLK(clk), .RST(rst), .I(in[266]), 
        .Q(round_reg[266]) );
  DFF \round_reg_reg[267]  ( .D(out[267]), .CLK(clk), .RST(rst), .I(in[267]), 
        .Q(round_reg[267]) );
  DFF \round_reg_reg[268]  ( .D(out[268]), .CLK(clk), .RST(rst), .I(in[268]), 
        .Q(round_reg[268]) );
  DFF \round_reg_reg[269]  ( .D(out[269]), .CLK(clk), .RST(rst), .I(in[269]), 
        .Q(round_reg[269]) );
  DFF \round_reg_reg[270]  ( .D(out[270]), .CLK(clk), .RST(rst), .I(in[270]), 
        .Q(round_reg[270]) );
  DFF \round_reg_reg[271]  ( .D(out[271]), .CLK(clk), .RST(rst), .I(in[271]), 
        .Q(round_reg[271]) );
  DFF \round_reg_reg[272]  ( .D(out[272]), .CLK(clk), .RST(rst), .I(in[272]), 
        .Q(round_reg[272]) );
  DFF \round_reg_reg[273]  ( .D(out[273]), .CLK(clk), .RST(rst), .I(in[273]), 
        .Q(round_reg[273]) );
  DFF \round_reg_reg[274]  ( .D(out[274]), .CLK(clk), .RST(rst), .I(in[274]), 
        .Q(round_reg[274]) );
  DFF \round_reg_reg[275]  ( .D(out[275]), .CLK(clk), .RST(rst), .I(in[275]), 
        .Q(round_reg[275]) );
  DFF \round_reg_reg[276]  ( .D(out[276]), .CLK(clk), .RST(rst), .I(in[276]), 
        .Q(round_reg[276]) );
  DFF \round_reg_reg[277]  ( .D(out[277]), .CLK(clk), .RST(rst), .I(in[277]), 
        .Q(round_reg[277]) );
  DFF \round_reg_reg[278]  ( .D(out[278]), .CLK(clk), .RST(rst), .I(in[278]), 
        .Q(round_reg[278]) );
  DFF \round_reg_reg[279]  ( .D(out[279]), .CLK(clk), .RST(rst), .I(in[279]), 
        .Q(round_reg[279]) );
  DFF \round_reg_reg[280]  ( .D(out[280]), .CLK(clk), .RST(rst), .I(in[280]), 
        .Q(round_reg[280]) );
  DFF \round_reg_reg[281]  ( .D(out[281]), .CLK(clk), .RST(rst), .I(in[281]), 
        .Q(round_reg[281]) );
  DFF \round_reg_reg[282]  ( .D(out[282]), .CLK(clk), .RST(rst), .I(in[282]), 
        .Q(round_reg[282]) );
  DFF \round_reg_reg[283]  ( .D(out[283]), .CLK(clk), .RST(rst), .I(in[283]), 
        .Q(round_reg[283]) );
  DFF \round_reg_reg[284]  ( .D(out[284]), .CLK(clk), .RST(rst), .I(in[284]), 
        .Q(round_reg[284]) );
  DFF \round_reg_reg[285]  ( .D(out[285]), .CLK(clk), .RST(rst), .I(in[285]), 
        .Q(round_reg[285]) );
  DFF \round_reg_reg[286]  ( .D(out[286]), .CLK(clk), .RST(rst), .I(in[286]), 
        .Q(round_reg[286]) );
  DFF \round_reg_reg[287]  ( .D(out[287]), .CLK(clk), .RST(rst), .I(in[287]), 
        .Q(round_reg[287]) );
  DFF \round_reg_reg[288]  ( .D(out[288]), .CLK(clk), .RST(rst), .I(in[288]), 
        .Q(round_reg[288]) );
  DFF \round_reg_reg[289]  ( .D(out[289]), .CLK(clk), .RST(rst), .I(in[289]), 
        .Q(round_reg[289]) );
  DFF \round_reg_reg[290]  ( .D(out[290]), .CLK(clk), .RST(rst), .I(in[290]), 
        .Q(round_reg[290]) );
  DFF \round_reg_reg[291]  ( .D(out[291]), .CLK(clk), .RST(rst), .I(in[291]), 
        .Q(round_reg[291]) );
  DFF \round_reg_reg[292]  ( .D(out[292]), .CLK(clk), .RST(rst), .I(in[292]), 
        .Q(round_reg[292]) );
  DFF \round_reg_reg[293]  ( .D(out[293]), .CLK(clk), .RST(rst), .I(in[293]), 
        .Q(round_reg[293]) );
  DFF \round_reg_reg[294]  ( .D(out[294]), .CLK(clk), .RST(rst), .I(in[294]), 
        .Q(round_reg[294]) );
  DFF \round_reg_reg[295]  ( .D(out[295]), .CLK(clk), .RST(rst), .I(in[295]), 
        .Q(round_reg[295]) );
  DFF \round_reg_reg[296]  ( .D(out[296]), .CLK(clk), .RST(rst), .I(in[296]), 
        .Q(round_reg[296]) );
  DFF \round_reg_reg[297]  ( .D(out[297]), .CLK(clk), .RST(rst), .I(in[297]), 
        .Q(round_reg[297]) );
  DFF \round_reg_reg[298]  ( .D(out[298]), .CLK(clk), .RST(rst), .I(in[298]), 
        .Q(round_reg[298]) );
  DFF \round_reg_reg[299]  ( .D(out[299]), .CLK(clk), .RST(rst), .I(in[299]), 
        .Q(round_reg[299]) );
  DFF \round_reg_reg[300]  ( .D(out[300]), .CLK(clk), .RST(rst), .I(in[300]), 
        .Q(round_reg[300]) );
  DFF \round_reg_reg[301]  ( .D(out[301]), .CLK(clk), .RST(rst), .I(in[301]), 
        .Q(round_reg[301]) );
  DFF \round_reg_reg[302]  ( .D(out[302]), .CLK(clk), .RST(rst), .I(in[302]), 
        .Q(round_reg[302]) );
  DFF \round_reg_reg[303]  ( .D(out[303]), .CLK(clk), .RST(rst), .I(in[303]), 
        .Q(round_reg[303]) );
  DFF \round_reg_reg[304]  ( .D(out[304]), .CLK(clk), .RST(rst), .I(in[304]), 
        .Q(round_reg[304]) );
  DFF \round_reg_reg[305]  ( .D(out[305]), .CLK(clk), .RST(rst), .I(in[305]), 
        .Q(round_reg[305]) );
  DFF \round_reg_reg[306]  ( .D(out[306]), .CLK(clk), .RST(rst), .I(in[306]), 
        .Q(round_reg[306]) );
  DFF \round_reg_reg[307]  ( .D(out[307]), .CLK(clk), .RST(rst), .I(in[307]), 
        .Q(round_reg[307]) );
  DFF \round_reg_reg[308]  ( .D(out[308]), .CLK(clk), .RST(rst), .I(in[308]), 
        .Q(round_reg[308]) );
  DFF \round_reg_reg[309]  ( .D(out[309]), .CLK(clk), .RST(rst), .I(in[309]), 
        .Q(round_reg[309]) );
  DFF \round_reg_reg[310]  ( .D(out[310]), .CLK(clk), .RST(rst), .I(in[310]), 
        .Q(round_reg[310]) );
  DFF \round_reg_reg[311]  ( .D(out[311]), .CLK(clk), .RST(rst), .I(in[311]), 
        .Q(round_reg[311]) );
  DFF \round_reg_reg[312]  ( .D(out[312]), .CLK(clk), .RST(rst), .I(in[312]), 
        .Q(round_reg[312]) );
  DFF \round_reg_reg[313]  ( .D(out[313]), .CLK(clk), .RST(rst), .I(in[313]), 
        .Q(round_reg[313]) );
  DFF \round_reg_reg[314]  ( .D(out[314]), .CLK(clk), .RST(rst), .I(in[314]), 
        .Q(round_reg[314]) );
  DFF \round_reg_reg[315]  ( .D(out[315]), .CLK(clk), .RST(rst), .I(in[315]), 
        .Q(round_reg[315]) );
  DFF \round_reg_reg[316]  ( .D(out[316]), .CLK(clk), .RST(rst), .I(in[316]), 
        .Q(round_reg[316]) );
  DFF \round_reg_reg[317]  ( .D(out[317]), .CLK(clk), .RST(rst), .I(in[317]), 
        .Q(round_reg[317]) );
  DFF \round_reg_reg[318]  ( .D(out[318]), .CLK(clk), .RST(rst), .I(in[318]), 
        .Q(round_reg[318]) );
  DFF \round_reg_reg[319]  ( .D(out[319]), .CLK(clk), .RST(rst), .I(in[319]), 
        .Q(round_reg[319]) );
  DFF \round_reg_reg[320]  ( .D(out[320]), .CLK(clk), .RST(rst), .I(in[320]), 
        .Q(round_reg[320]) );
  DFF \round_reg_reg[321]  ( .D(out[321]), .CLK(clk), .RST(rst), .I(in[321]), 
        .Q(round_reg[321]) );
  DFF \round_reg_reg[322]  ( .D(out[322]), .CLK(clk), .RST(rst), .I(in[322]), 
        .Q(round_reg[322]) );
  DFF \round_reg_reg[323]  ( .D(out[323]), .CLK(clk), .RST(rst), .I(in[323]), 
        .Q(round_reg[323]) );
  DFF \round_reg_reg[324]  ( .D(out[324]), .CLK(clk), .RST(rst), .I(in[324]), 
        .Q(round_reg[324]) );
  DFF \round_reg_reg[325]  ( .D(out[325]), .CLK(clk), .RST(rst), .I(in[325]), 
        .Q(round_reg[325]) );
  DFF \round_reg_reg[326]  ( .D(out[326]), .CLK(clk), .RST(rst), .I(in[326]), 
        .Q(round_reg[326]) );
  DFF \round_reg_reg[327]  ( .D(out[327]), .CLK(clk), .RST(rst), .I(in[327]), 
        .Q(round_reg[327]) );
  DFF \round_reg_reg[328]  ( .D(out[328]), .CLK(clk), .RST(rst), .I(in[328]), 
        .Q(round_reg[328]) );
  DFF \round_reg_reg[329]  ( .D(out[329]), .CLK(clk), .RST(rst), .I(in[329]), 
        .Q(round_reg[329]) );
  DFF \round_reg_reg[330]  ( .D(out[330]), .CLK(clk), .RST(rst), .I(in[330]), 
        .Q(round_reg[330]) );
  DFF \round_reg_reg[331]  ( .D(out[331]), .CLK(clk), .RST(rst), .I(in[331]), 
        .Q(round_reg[331]) );
  DFF \round_reg_reg[332]  ( .D(out[332]), .CLK(clk), .RST(rst), .I(in[332]), 
        .Q(round_reg[332]) );
  DFF \round_reg_reg[333]  ( .D(out[333]), .CLK(clk), .RST(rst), .I(in[333]), 
        .Q(round_reg[333]) );
  DFF \round_reg_reg[334]  ( .D(out[334]), .CLK(clk), .RST(rst), .I(in[334]), 
        .Q(round_reg[334]) );
  DFF \round_reg_reg[335]  ( .D(out[335]), .CLK(clk), .RST(rst), .I(in[335]), 
        .Q(round_reg[335]) );
  DFF \round_reg_reg[336]  ( .D(out[336]), .CLK(clk), .RST(rst), .I(in[336]), 
        .Q(round_reg[336]) );
  DFF \round_reg_reg[337]  ( .D(out[337]), .CLK(clk), .RST(rst), .I(in[337]), 
        .Q(round_reg[337]) );
  DFF \round_reg_reg[338]  ( .D(out[338]), .CLK(clk), .RST(rst), .I(in[338]), 
        .Q(round_reg[338]) );
  DFF \round_reg_reg[339]  ( .D(out[339]), .CLK(clk), .RST(rst), .I(in[339]), 
        .Q(round_reg[339]) );
  DFF \round_reg_reg[340]  ( .D(out[340]), .CLK(clk), .RST(rst), .I(in[340]), 
        .Q(round_reg[340]) );
  DFF \round_reg_reg[341]  ( .D(out[341]), .CLK(clk), .RST(rst), .I(in[341]), 
        .Q(round_reg[341]) );
  DFF \round_reg_reg[342]  ( .D(out[342]), .CLK(clk), .RST(rst), .I(in[342]), 
        .Q(round_reg[342]) );
  DFF \round_reg_reg[343]  ( .D(out[343]), .CLK(clk), .RST(rst), .I(in[343]), 
        .Q(round_reg[343]) );
  DFF \round_reg_reg[344]  ( .D(out[344]), .CLK(clk), .RST(rst), .I(in[344]), 
        .Q(round_reg[344]) );
  DFF \round_reg_reg[345]  ( .D(out[345]), .CLK(clk), .RST(rst), .I(in[345]), 
        .Q(round_reg[345]) );
  DFF \round_reg_reg[346]  ( .D(out[346]), .CLK(clk), .RST(rst), .I(in[346]), 
        .Q(round_reg[346]) );
  DFF \round_reg_reg[347]  ( .D(out[347]), .CLK(clk), .RST(rst), .I(in[347]), 
        .Q(round_reg[347]) );
  DFF \round_reg_reg[348]  ( .D(out[348]), .CLK(clk), .RST(rst), .I(in[348]), 
        .Q(round_reg[348]) );
  DFF \round_reg_reg[349]  ( .D(out[349]), .CLK(clk), .RST(rst), .I(in[349]), 
        .Q(round_reg[349]) );
  DFF \round_reg_reg[350]  ( .D(out[350]), .CLK(clk), .RST(rst), .I(in[350]), 
        .Q(round_reg[350]) );
  DFF \round_reg_reg[351]  ( .D(out[351]), .CLK(clk), .RST(rst), .I(in[351]), 
        .Q(round_reg[351]) );
  DFF \round_reg_reg[352]  ( .D(out[352]), .CLK(clk), .RST(rst), .I(in[352]), 
        .Q(round_reg[352]) );
  DFF \round_reg_reg[353]  ( .D(out[353]), .CLK(clk), .RST(rst), .I(in[353]), 
        .Q(round_reg[353]) );
  DFF \round_reg_reg[354]  ( .D(out[354]), .CLK(clk), .RST(rst), .I(in[354]), 
        .Q(round_reg[354]) );
  DFF \round_reg_reg[355]  ( .D(out[355]), .CLK(clk), .RST(rst), .I(in[355]), 
        .Q(round_reg[355]) );
  DFF \round_reg_reg[356]  ( .D(out[356]), .CLK(clk), .RST(rst), .I(in[356]), 
        .Q(round_reg[356]) );
  DFF \round_reg_reg[357]  ( .D(out[357]), .CLK(clk), .RST(rst), .I(in[357]), 
        .Q(round_reg[357]) );
  DFF \round_reg_reg[358]  ( .D(out[358]), .CLK(clk), .RST(rst), .I(in[358]), 
        .Q(round_reg[358]) );
  DFF \round_reg_reg[359]  ( .D(out[359]), .CLK(clk), .RST(rst), .I(in[359]), 
        .Q(round_reg[359]) );
  DFF \round_reg_reg[360]  ( .D(out[360]), .CLK(clk), .RST(rst), .I(in[360]), 
        .Q(round_reg[360]) );
  DFF \round_reg_reg[361]  ( .D(out[361]), .CLK(clk), .RST(rst), .I(in[361]), 
        .Q(round_reg[361]) );
  DFF \round_reg_reg[362]  ( .D(out[362]), .CLK(clk), .RST(rst), .I(in[362]), 
        .Q(round_reg[362]) );
  DFF \round_reg_reg[363]  ( .D(out[363]), .CLK(clk), .RST(rst), .I(in[363]), 
        .Q(round_reg[363]) );
  DFF \round_reg_reg[364]  ( .D(out[364]), .CLK(clk), .RST(rst), .I(in[364]), 
        .Q(round_reg[364]) );
  DFF \round_reg_reg[365]  ( .D(out[365]), .CLK(clk), .RST(rst), .I(in[365]), 
        .Q(round_reg[365]) );
  DFF \round_reg_reg[366]  ( .D(out[366]), .CLK(clk), .RST(rst), .I(in[366]), 
        .Q(round_reg[366]) );
  DFF \round_reg_reg[367]  ( .D(out[367]), .CLK(clk), .RST(rst), .I(in[367]), 
        .Q(round_reg[367]) );
  DFF \round_reg_reg[368]  ( .D(out[368]), .CLK(clk), .RST(rst), .I(in[368]), 
        .Q(round_reg[368]) );
  DFF \round_reg_reg[369]  ( .D(out[369]), .CLK(clk), .RST(rst), .I(in[369]), 
        .Q(round_reg[369]) );
  DFF \round_reg_reg[370]  ( .D(out[370]), .CLK(clk), .RST(rst), .I(in[370]), 
        .Q(round_reg[370]) );
  DFF \round_reg_reg[371]  ( .D(out[371]), .CLK(clk), .RST(rst), .I(in[371]), 
        .Q(round_reg[371]) );
  DFF \round_reg_reg[372]  ( .D(out[372]), .CLK(clk), .RST(rst), .I(in[372]), 
        .Q(round_reg[372]) );
  DFF \round_reg_reg[373]  ( .D(out[373]), .CLK(clk), .RST(rst), .I(in[373]), 
        .Q(round_reg[373]) );
  DFF \round_reg_reg[374]  ( .D(out[374]), .CLK(clk), .RST(rst), .I(in[374]), 
        .Q(round_reg[374]) );
  DFF \round_reg_reg[375]  ( .D(out[375]), .CLK(clk), .RST(rst), .I(in[375]), 
        .Q(round_reg[375]) );
  DFF \round_reg_reg[376]  ( .D(out[376]), .CLK(clk), .RST(rst), .I(in[376]), 
        .Q(round_reg[376]) );
  DFF \round_reg_reg[377]  ( .D(out[377]), .CLK(clk), .RST(rst), .I(in[377]), 
        .Q(round_reg[377]) );
  DFF \round_reg_reg[378]  ( .D(out[378]), .CLK(clk), .RST(rst), .I(in[378]), 
        .Q(round_reg[378]) );
  DFF \round_reg_reg[379]  ( .D(out[379]), .CLK(clk), .RST(rst), .I(in[379]), 
        .Q(round_reg[379]) );
  DFF \round_reg_reg[380]  ( .D(out[380]), .CLK(clk), .RST(rst), .I(in[380]), 
        .Q(round_reg[380]) );
  DFF \round_reg_reg[381]  ( .D(out[381]), .CLK(clk), .RST(rst), .I(in[381]), 
        .Q(round_reg[381]) );
  DFF \round_reg_reg[382]  ( .D(out[382]), .CLK(clk), .RST(rst), .I(in[382]), 
        .Q(round_reg[382]) );
  DFF \round_reg_reg[383]  ( .D(out[383]), .CLK(clk), .RST(rst), .I(in[383]), 
        .Q(round_reg[383]) );
  DFF \round_reg_reg[384]  ( .D(out[384]), .CLK(clk), .RST(rst), .I(in[384]), 
        .Q(round_reg[384]) );
  DFF \round_reg_reg[385]  ( .D(out[385]), .CLK(clk), .RST(rst), .I(in[385]), 
        .Q(round_reg[385]) );
  DFF \round_reg_reg[386]  ( .D(out[386]), .CLK(clk), .RST(rst), .I(in[386]), 
        .Q(round_reg[386]) );
  DFF \round_reg_reg[387]  ( .D(out[387]), .CLK(clk), .RST(rst), .I(in[387]), 
        .Q(round_reg[387]) );
  DFF \round_reg_reg[388]  ( .D(out[388]), .CLK(clk), .RST(rst), .I(in[388]), 
        .Q(round_reg[388]) );
  DFF \round_reg_reg[389]  ( .D(out[389]), .CLK(clk), .RST(rst), .I(in[389]), 
        .Q(round_reg[389]) );
  DFF \round_reg_reg[390]  ( .D(out[390]), .CLK(clk), .RST(rst), .I(in[390]), 
        .Q(round_reg[390]) );
  DFF \round_reg_reg[391]  ( .D(out[391]), .CLK(clk), .RST(rst), .I(in[391]), 
        .Q(round_reg[391]) );
  DFF \round_reg_reg[392]  ( .D(out[392]), .CLK(clk), .RST(rst), .I(in[392]), 
        .Q(round_reg[392]) );
  DFF \round_reg_reg[393]  ( .D(out[393]), .CLK(clk), .RST(rst), .I(in[393]), 
        .Q(round_reg[393]) );
  DFF \round_reg_reg[394]  ( .D(out[394]), .CLK(clk), .RST(rst), .I(in[394]), 
        .Q(round_reg[394]) );
  DFF \round_reg_reg[395]  ( .D(out[395]), .CLK(clk), .RST(rst), .I(in[395]), 
        .Q(round_reg[395]) );
  DFF \round_reg_reg[396]  ( .D(out[396]), .CLK(clk), .RST(rst), .I(in[396]), 
        .Q(round_reg[396]) );
  DFF \round_reg_reg[397]  ( .D(out[397]), .CLK(clk), .RST(rst), .I(in[397]), 
        .Q(round_reg[397]) );
  DFF \round_reg_reg[398]  ( .D(out[398]), .CLK(clk), .RST(rst), .I(in[398]), 
        .Q(round_reg[398]) );
  DFF \round_reg_reg[399]  ( .D(out[399]), .CLK(clk), .RST(rst), .I(in[399]), 
        .Q(round_reg[399]) );
  DFF \round_reg_reg[400]  ( .D(out[400]), .CLK(clk), .RST(rst), .I(in[400]), 
        .Q(round_reg[400]) );
  DFF \round_reg_reg[401]  ( .D(out[401]), .CLK(clk), .RST(rst), .I(in[401]), 
        .Q(round_reg[401]) );
  DFF \round_reg_reg[402]  ( .D(out[402]), .CLK(clk), .RST(rst), .I(in[402]), 
        .Q(round_reg[402]) );
  DFF \round_reg_reg[403]  ( .D(out[403]), .CLK(clk), .RST(rst), .I(in[403]), 
        .Q(round_reg[403]) );
  DFF \round_reg_reg[404]  ( .D(out[404]), .CLK(clk), .RST(rst), .I(in[404]), 
        .Q(round_reg[404]) );
  DFF \round_reg_reg[405]  ( .D(out[405]), .CLK(clk), .RST(rst), .I(in[405]), 
        .Q(round_reg[405]) );
  DFF \round_reg_reg[406]  ( .D(out[406]), .CLK(clk), .RST(rst), .I(in[406]), 
        .Q(round_reg[406]) );
  DFF \round_reg_reg[407]  ( .D(out[407]), .CLK(clk), .RST(rst), .I(in[407]), 
        .Q(round_reg[407]) );
  DFF \round_reg_reg[408]  ( .D(out[408]), .CLK(clk), .RST(rst), .I(in[408]), 
        .Q(round_reg[408]) );
  DFF \round_reg_reg[409]  ( .D(out[409]), .CLK(clk), .RST(rst), .I(in[409]), 
        .Q(round_reg[409]) );
  DFF \round_reg_reg[410]  ( .D(out[410]), .CLK(clk), .RST(rst), .I(in[410]), 
        .Q(round_reg[410]) );
  DFF \round_reg_reg[411]  ( .D(out[411]), .CLK(clk), .RST(rst), .I(in[411]), 
        .Q(round_reg[411]) );
  DFF \round_reg_reg[412]  ( .D(out[412]), .CLK(clk), .RST(rst), .I(in[412]), 
        .Q(round_reg[412]) );
  DFF \round_reg_reg[413]  ( .D(out[413]), .CLK(clk), .RST(rst), .I(in[413]), 
        .Q(round_reg[413]) );
  DFF \round_reg_reg[414]  ( .D(out[414]), .CLK(clk), .RST(rst), .I(in[414]), 
        .Q(round_reg[414]) );
  DFF \round_reg_reg[415]  ( .D(out[415]), .CLK(clk), .RST(rst), .I(in[415]), 
        .Q(round_reg[415]) );
  DFF \round_reg_reg[416]  ( .D(out[416]), .CLK(clk), .RST(rst), .I(in[416]), 
        .Q(round_reg[416]) );
  DFF \round_reg_reg[417]  ( .D(out[417]), .CLK(clk), .RST(rst), .I(in[417]), 
        .Q(round_reg[417]) );
  DFF \round_reg_reg[418]  ( .D(out[418]), .CLK(clk), .RST(rst), .I(in[418]), 
        .Q(round_reg[418]) );
  DFF \round_reg_reg[419]  ( .D(out[419]), .CLK(clk), .RST(rst), .I(in[419]), 
        .Q(round_reg[419]) );
  DFF \round_reg_reg[420]  ( .D(out[420]), .CLK(clk), .RST(rst), .I(in[420]), 
        .Q(round_reg[420]) );
  DFF \round_reg_reg[421]  ( .D(out[421]), .CLK(clk), .RST(rst), .I(in[421]), 
        .Q(round_reg[421]) );
  DFF \round_reg_reg[422]  ( .D(out[422]), .CLK(clk), .RST(rst), .I(in[422]), 
        .Q(round_reg[422]) );
  DFF \round_reg_reg[423]  ( .D(out[423]), .CLK(clk), .RST(rst), .I(in[423]), 
        .Q(round_reg[423]) );
  DFF \round_reg_reg[424]  ( .D(out[424]), .CLK(clk), .RST(rst), .I(in[424]), 
        .Q(round_reg[424]) );
  DFF \round_reg_reg[425]  ( .D(out[425]), .CLK(clk), .RST(rst), .I(in[425]), 
        .Q(round_reg[425]) );
  DFF \round_reg_reg[426]  ( .D(out[426]), .CLK(clk), .RST(rst), .I(in[426]), 
        .Q(round_reg[426]) );
  DFF \round_reg_reg[427]  ( .D(out[427]), .CLK(clk), .RST(rst), .I(in[427]), 
        .Q(round_reg[427]) );
  DFF \round_reg_reg[428]  ( .D(out[428]), .CLK(clk), .RST(rst), .I(in[428]), 
        .Q(round_reg[428]) );
  DFF \round_reg_reg[429]  ( .D(out[429]), .CLK(clk), .RST(rst), .I(in[429]), 
        .Q(round_reg[429]) );
  DFF \round_reg_reg[430]  ( .D(out[430]), .CLK(clk), .RST(rst), .I(in[430]), 
        .Q(round_reg[430]) );
  DFF \round_reg_reg[431]  ( .D(out[431]), .CLK(clk), .RST(rst), .I(in[431]), 
        .Q(round_reg[431]) );
  DFF \round_reg_reg[432]  ( .D(out[432]), .CLK(clk), .RST(rst), .I(in[432]), 
        .Q(round_reg[432]) );
  DFF \round_reg_reg[433]  ( .D(out[433]), .CLK(clk), .RST(rst), .I(in[433]), 
        .Q(round_reg[433]) );
  DFF \round_reg_reg[434]  ( .D(out[434]), .CLK(clk), .RST(rst), .I(in[434]), 
        .Q(round_reg[434]) );
  DFF \round_reg_reg[435]  ( .D(out[435]), .CLK(clk), .RST(rst), .I(in[435]), 
        .Q(round_reg[435]) );
  DFF \round_reg_reg[436]  ( .D(out[436]), .CLK(clk), .RST(rst), .I(in[436]), 
        .Q(round_reg[436]) );
  DFF \round_reg_reg[437]  ( .D(out[437]), .CLK(clk), .RST(rst), .I(in[437]), 
        .Q(round_reg[437]) );
  DFF \round_reg_reg[438]  ( .D(out[438]), .CLK(clk), .RST(rst), .I(in[438]), 
        .Q(round_reg[438]) );
  DFF \round_reg_reg[439]  ( .D(out[439]), .CLK(clk), .RST(rst), .I(in[439]), 
        .Q(round_reg[439]) );
  DFF \round_reg_reg[440]  ( .D(out[440]), .CLK(clk), .RST(rst), .I(in[440]), 
        .Q(round_reg[440]) );
  DFF \round_reg_reg[441]  ( .D(out[441]), .CLK(clk), .RST(rst), .I(in[441]), 
        .Q(round_reg[441]) );
  DFF \round_reg_reg[442]  ( .D(out[442]), .CLK(clk), .RST(rst), .I(in[442]), 
        .Q(round_reg[442]) );
  DFF \round_reg_reg[443]  ( .D(out[443]), .CLK(clk), .RST(rst), .I(in[443]), 
        .Q(round_reg[443]) );
  DFF \round_reg_reg[444]  ( .D(out[444]), .CLK(clk), .RST(rst), .I(in[444]), 
        .Q(round_reg[444]) );
  DFF \round_reg_reg[445]  ( .D(out[445]), .CLK(clk), .RST(rst), .I(in[445]), 
        .Q(round_reg[445]) );
  DFF \round_reg_reg[446]  ( .D(out[446]), .CLK(clk), .RST(rst), .I(in[446]), 
        .Q(round_reg[446]) );
  DFF \round_reg_reg[447]  ( .D(out[447]), .CLK(clk), .RST(rst), .I(in[447]), 
        .Q(round_reg[447]) );
  DFF \round_reg_reg[448]  ( .D(out[448]), .CLK(clk), .RST(rst), .I(in[448]), 
        .Q(round_reg[448]) );
  DFF \round_reg_reg[449]  ( .D(out[449]), .CLK(clk), .RST(rst), .I(in[449]), 
        .Q(round_reg[449]) );
  DFF \round_reg_reg[450]  ( .D(out[450]), .CLK(clk), .RST(rst), .I(in[450]), 
        .Q(round_reg[450]) );
  DFF \round_reg_reg[451]  ( .D(out[451]), .CLK(clk), .RST(rst), .I(in[451]), 
        .Q(round_reg[451]) );
  DFF \round_reg_reg[452]  ( .D(out[452]), .CLK(clk), .RST(rst), .I(in[452]), 
        .Q(round_reg[452]) );
  DFF \round_reg_reg[453]  ( .D(out[453]), .CLK(clk), .RST(rst), .I(in[453]), 
        .Q(round_reg[453]) );
  DFF \round_reg_reg[454]  ( .D(out[454]), .CLK(clk), .RST(rst), .I(in[454]), 
        .Q(round_reg[454]) );
  DFF \round_reg_reg[455]  ( .D(out[455]), .CLK(clk), .RST(rst), .I(in[455]), 
        .Q(round_reg[455]) );
  DFF \round_reg_reg[456]  ( .D(out[456]), .CLK(clk), .RST(rst), .I(in[456]), 
        .Q(round_reg[456]) );
  DFF \round_reg_reg[457]  ( .D(out[457]), .CLK(clk), .RST(rst), .I(in[457]), 
        .Q(round_reg[457]) );
  DFF \round_reg_reg[458]  ( .D(out[458]), .CLK(clk), .RST(rst), .I(in[458]), 
        .Q(round_reg[458]) );
  DFF \round_reg_reg[459]  ( .D(out[459]), .CLK(clk), .RST(rst), .I(in[459]), 
        .Q(round_reg[459]) );
  DFF \round_reg_reg[460]  ( .D(out[460]), .CLK(clk), .RST(rst), .I(in[460]), 
        .Q(round_reg[460]) );
  DFF \round_reg_reg[461]  ( .D(out[461]), .CLK(clk), .RST(rst), .I(in[461]), 
        .Q(round_reg[461]) );
  DFF \round_reg_reg[462]  ( .D(out[462]), .CLK(clk), .RST(rst), .I(in[462]), 
        .Q(round_reg[462]) );
  DFF \round_reg_reg[463]  ( .D(out[463]), .CLK(clk), .RST(rst), .I(in[463]), 
        .Q(round_reg[463]) );
  DFF \round_reg_reg[464]  ( .D(out[464]), .CLK(clk), .RST(rst), .I(in[464]), 
        .Q(round_reg[464]) );
  DFF \round_reg_reg[465]  ( .D(out[465]), .CLK(clk), .RST(rst), .I(in[465]), 
        .Q(round_reg[465]) );
  DFF \round_reg_reg[466]  ( .D(out[466]), .CLK(clk), .RST(rst), .I(in[466]), 
        .Q(round_reg[466]) );
  DFF \round_reg_reg[467]  ( .D(out[467]), .CLK(clk), .RST(rst), .I(in[467]), 
        .Q(round_reg[467]) );
  DFF \round_reg_reg[468]  ( .D(out[468]), .CLK(clk), .RST(rst), .I(in[468]), 
        .Q(round_reg[468]) );
  DFF \round_reg_reg[469]  ( .D(out[469]), .CLK(clk), .RST(rst), .I(in[469]), 
        .Q(round_reg[469]) );
  DFF \round_reg_reg[470]  ( .D(out[470]), .CLK(clk), .RST(rst), .I(in[470]), 
        .Q(round_reg[470]) );
  DFF \round_reg_reg[471]  ( .D(out[471]), .CLK(clk), .RST(rst), .I(in[471]), 
        .Q(round_reg[471]) );
  DFF \round_reg_reg[472]  ( .D(out[472]), .CLK(clk), .RST(rst), .I(in[472]), 
        .Q(round_reg[472]) );
  DFF \round_reg_reg[473]  ( .D(out[473]), .CLK(clk), .RST(rst), .I(in[473]), 
        .Q(round_reg[473]) );
  DFF \round_reg_reg[474]  ( .D(out[474]), .CLK(clk), .RST(rst), .I(in[474]), 
        .Q(round_reg[474]) );
  DFF \round_reg_reg[475]  ( .D(out[475]), .CLK(clk), .RST(rst), .I(in[475]), 
        .Q(round_reg[475]) );
  DFF \round_reg_reg[476]  ( .D(out[476]), .CLK(clk), .RST(rst), .I(in[476]), 
        .Q(round_reg[476]) );
  DFF \round_reg_reg[477]  ( .D(out[477]), .CLK(clk), .RST(rst), .I(in[477]), 
        .Q(round_reg[477]) );
  DFF \round_reg_reg[478]  ( .D(out[478]), .CLK(clk), .RST(rst), .I(in[478]), 
        .Q(round_reg[478]) );
  DFF \round_reg_reg[479]  ( .D(out[479]), .CLK(clk), .RST(rst), .I(in[479]), 
        .Q(round_reg[479]) );
  DFF \round_reg_reg[480]  ( .D(out[480]), .CLK(clk), .RST(rst), .I(in[480]), 
        .Q(round_reg[480]) );
  DFF \round_reg_reg[481]  ( .D(out[481]), .CLK(clk), .RST(rst), .I(in[481]), 
        .Q(round_reg[481]) );
  DFF \round_reg_reg[482]  ( .D(out[482]), .CLK(clk), .RST(rst), .I(in[482]), 
        .Q(round_reg[482]) );
  DFF \round_reg_reg[483]  ( .D(out[483]), .CLK(clk), .RST(rst), .I(in[483]), 
        .Q(round_reg[483]) );
  DFF \round_reg_reg[484]  ( .D(out[484]), .CLK(clk), .RST(rst), .I(in[484]), 
        .Q(round_reg[484]) );
  DFF \round_reg_reg[485]  ( .D(out[485]), .CLK(clk), .RST(rst), .I(in[485]), 
        .Q(round_reg[485]) );
  DFF \round_reg_reg[486]  ( .D(out[486]), .CLK(clk), .RST(rst), .I(in[486]), 
        .Q(round_reg[486]) );
  DFF \round_reg_reg[487]  ( .D(out[487]), .CLK(clk), .RST(rst), .I(in[487]), 
        .Q(round_reg[487]) );
  DFF \round_reg_reg[488]  ( .D(out[488]), .CLK(clk), .RST(rst), .I(in[488]), 
        .Q(round_reg[488]) );
  DFF \round_reg_reg[489]  ( .D(out[489]), .CLK(clk), .RST(rst), .I(in[489]), 
        .Q(round_reg[489]) );
  DFF \round_reg_reg[490]  ( .D(out[490]), .CLK(clk), .RST(rst), .I(in[490]), 
        .Q(round_reg[490]) );
  DFF \round_reg_reg[491]  ( .D(out[491]), .CLK(clk), .RST(rst), .I(in[491]), 
        .Q(round_reg[491]) );
  DFF \round_reg_reg[492]  ( .D(out[492]), .CLK(clk), .RST(rst), .I(in[492]), 
        .Q(round_reg[492]) );
  DFF \round_reg_reg[493]  ( .D(out[493]), .CLK(clk), .RST(rst), .I(in[493]), 
        .Q(round_reg[493]) );
  DFF \round_reg_reg[494]  ( .D(out[494]), .CLK(clk), .RST(rst), .I(in[494]), 
        .Q(round_reg[494]) );
  DFF \round_reg_reg[495]  ( .D(out[495]), .CLK(clk), .RST(rst), .I(in[495]), 
        .Q(round_reg[495]) );
  DFF \round_reg_reg[496]  ( .D(out[496]), .CLK(clk), .RST(rst), .I(in[496]), 
        .Q(round_reg[496]) );
  DFF \round_reg_reg[497]  ( .D(out[497]), .CLK(clk), .RST(rst), .I(in[497]), 
        .Q(round_reg[497]) );
  DFF \round_reg_reg[498]  ( .D(out[498]), .CLK(clk), .RST(rst), .I(in[498]), 
        .Q(round_reg[498]) );
  DFF \round_reg_reg[499]  ( .D(out[499]), .CLK(clk), .RST(rst), .I(in[499]), 
        .Q(round_reg[499]) );
  DFF \round_reg_reg[500]  ( .D(out[500]), .CLK(clk), .RST(rst), .I(in[500]), 
        .Q(round_reg[500]) );
  DFF \round_reg_reg[501]  ( .D(out[501]), .CLK(clk), .RST(rst), .I(in[501]), 
        .Q(round_reg[501]) );
  DFF \round_reg_reg[502]  ( .D(out[502]), .CLK(clk), .RST(rst), .I(in[502]), 
        .Q(round_reg[502]) );
  DFF \round_reg_reg[503]  ( .D(out[503]), .CLK(clk), .RST(rst), .I(in[503]), 
        .Q(round_reg[503]) );
  DFF \round_reg_reg[504]  ( .D(out[504]), .CLK(clk), .RST(rst), .I(in[504]), 
        .Q(round_reg[504]) );
  DFF \round_reg_reg[505]  ( .D(out[505]), .CLK(clk), .RST(rst), .I(in[505]), 
        .Q(round_reg[505]) );
  DFF \round_reg_reg[506]  ( .D(out[506]), .CLK(clk), .RST(rst), .I(in[506]), 
        .Q(round_reg[506]) );
  DFF \round_reg_reg[507]  ( .D(out[507]), .CLK(clk), .RST(rst), .I(in[507]), 
        .Q(round_reg[507]) );
  DFF \round_reg_reg[508]  ( .D(out[508]), .CLK(clk), .RST(rst), .I(in[508]), 
        .Q(round_reg[508]) );
  DFF \round_reg_reg[509]  ( .D(out[509]), .CLK(clk), .RST(rst), .I(in[509]), 
        .Q(round_reg[509]) );
  DFF \round_reg_reg[510]  ( .D(out[510]), .CLK(clk), .RST(rst), .I(in[510]), 
        .Q(round_reg[510]) );
  DFF \round_reg_reg[511]  ( .D(out[511]), .CLK(clk), .RST(rst), .I(in[511]), 
        .Q(round_reg[511]) );
  DFF \round_reg_reg[512]  ( .D(out[512]), .CLK(clk), .RST(rst), .I(in[512]), 
        .Q(round_reg[512]) );
  DFF \round_reg_reg[513]  ( .D(out[513]), .CLK(clk), .RST(rst), .I(in[513]), 
        .Q(round_reg[513]) );
  DFF \round_reg_reg[514]  ( .D(out[514]), .CLK(clk), .RST(rst), .I(in[514]), 
        .Q(round_reg[514]) );
  DFF \round_reg_reg[515]  ( .D(out[515]), .CLK(clk), .RST(rst), .I(in[515]), 
        .Q(round_reg[515]) );
  DFF \round_reg_reg[516]  ( .D(out[516]), .CLK(clk), .RST(rst), .I(in[516]), 
        .Q(round_reg[516]) );
  DFF \round_reg_reg[517]  ( .D(out[517]), .CLK(clk), .RST(rst), .I(in[517]), 
        .Q(round_reg[517]) );
  DFF \round_reg_reg[518]  ( .D(out[518]), .CLK(clk), .RST(rst), .I(in[518]), 
        .Q(round_reg[518]) );
  DFF \round_reg_reg[519]  ( .D(out[519]), .CLK(clk), .RST(rst), .I(in[519]), 
        .Q(round_reg[519]) );
  DFF \round_reg_reg[520]  ( .D(out[520]), .CLK(clk), .RST(rst), .I(in[520]), 
        .Q(round_reg[520]) );
  DFF \round_reg_reg[521]  ( .D(out[521]), .CLK(clk), .RST(rst), .I(in[521]), 
        .Q(round_reg[521]) );
  DFF \round_reg_reg[522]  ( .D(out[522]), .CLK(clk), .RST(rst), .I(in[522]), 
        .Q(round_reg[522]) );
  DFF \round_reg_reg[523]  ( .D(out[523]), .CLK(clk), .RST(rst), .I(in[523]), 
        .Q(round_reg[523]) );
  DFF \round_reg_reg[524]  ( .D(out[524]), .CLK(clk), .RST(rst), .I(in[524]), 
        .Q(round_reg[524]) );
  DFF \round_reg_reg[525]  ( .D(out[525]), .CLK(clk), .RST(rst), .I(in[525]), 
        .Q(round_reg[525]) );
  DFF \round_reg_reg[526]  ( .D(out[526]), .CLK(clk), .RST(rst), .I(in[526]), 
        .Q(round_reg[526]) );
  DFF \round_reg_reg[527]  ( .D(out[527]), .CLK(clk), .RST(rst), .I(in[527]), 
        .Q(round_reg[527]) );
  DFF \round_reg_reg[528]  ( .D(out[528]), .CLK(clk), .RST(rst), .I(in[528]), 
        .Q(round_reg[528]) );
  DFF \round_reg_reg[529]  ( .D(out[529]), .CLK(clk), .RST(rst), .I(in[529]), 
        .Q(round_reg[529]) );
  DFF \round_reg_reg[530]  ( .D(out[530]), .CLK(clk), .RST(rst), .I(in[530]), 
        .Q(round_reg[530]) );
  DFF \round_reg_reg[531]  ( .D(out[531]), .CLK(clk), .RST(rst), .I(in[531]), 
        .Q(round_reg[531]) );
  DFF \round_reg_reg[532]  ( .D(out[532]), .CLK(clk), .RST(rst), .I(in[532]), 
        .Q(round_reg[532]) );
  DFF \round_reg_reg[533]  ( .D(out[533]), .CLK(clk), .RST(rst), .I(in[533]), 
        .Q(round_reg[533]) );
  DFF \round_reg_reg[534]  ( .D(out[534]), .CLK(clk), .RST(rst), .I(in[534]), 
        .Q(round_reg[534]) );
  DFF \round_reg_reg[535]  ( .D(out[535]), .CLK(clk), .RST(rst), .I(in[535]), 
        .Q(round_reg[535]) );
  DFF \round_reg_reg[536]  ( .D(out[536]), .CLK(clk), .RST(rst), .I(in[536]), 
        .Q(round_reg[536]) );
  DFF \round_reg_reg[537]  ( .D(out[537]), .CLK(clk), .RST(rst), .I(in[537]), 
        .Q(round_reg[537]) );
  DFF \round_reg_reg[538]  ( .D(out[538]), .CLK(clk), .RST(rst), .I(in[538]), 
        .Q(round_reg[538]) );
  DFF \round_reg_reg[539]  ( .D(out[539]), .CLK(clk), .RST(rst), .I(in[539]), 
        .Q(round_reg[539]) );
  DFF \round_reg_reg[540]  ( .D(out[540]), .CLK(clk), .RST(rst), .I(in[540]), 
        .Q(round_reg[540]) );
  DFF \round_reg_reg[541]  ( .D(out[541]), .CLK(clk), .RST(rst), .I(in[541]), 
        .Q(round_reg[541]) );
  DFF \round_reg_reg[542]  ( .D(out[542]), .CLK(clk), .RST(rst), .I(in[542]), 
        .Q(round_reg[542]) );
  DFF \round_reg_reg[543]  ( .D(out[543]), .CLK(clk), .RST(rst), .I(in[543]), 
        .Q(round_reg[543]) );
  DFF \round_reg_reg[544]  ( .D(out[544]), .CLK(clk), .RST(rst), .I(in[544]), 
        .Q(round_reg[544]) );
  DFF \round_reg_reg[545]  ( .D(out[545]), .CLK(clk), .RST(rst), .I(in[545]), 
        .Q(round_reg[545]) );
  DFF \round_reg_reg[546]  ( .D(out[546]), .CLK(clk), .RST(rst), .I(in[546]), 
        .Q(round_reg[546]) );
  DFF \round_reg_reg[547]  ( .D(out[547]), .CLK(clk), .RST(rst), .I(in[547]), 
        .Q(round_reg[547]) );
  DFF \round_reg_reg[548]  ( .D(out[548]), .CLK(clk), .RST(rst), .I(in[548]), 
        .Q(round_reg[548]) );
  DFF \round_reg_reg[549]  ( .D(out[549]), .CLK(clk), .RST(rst), .I(in[549]), 
        .Q(round_reg[549]) );
  DFF \round_reg_reg[550]  ( .D(out[550]), .CLK(clk), .RST(rst), .I(in[550]), 
        .Q(round_reg[550]) );
  DFF \round_reg_reg[551]  ( .D(out[551]), .CLK(clk), .RST(rst), .I(in[551]), 
        .Q(round_reg[551]) );
  DFF \round_reg_reg[552]  ( .D(out[552]), .CLK(clk), .RST(rst), .I(in[552]), 
        .Q(round_reg[552]) );
  DFF \round_reg_reg[553]  ( .D(out[553]), .CLK(clk), .RST(rst), .I(in[553]), 
        .Q(round_reg[553]) );
  DFF \round_reg_reg[554]  ( .D(out[554]), .CLK(clk), .RST(rst), .I(in[554]), 
        .Q(round_reg[554]) );
  DFF \round_reg_reg[555]  ( .D(out[555]), .CLK(clk), .RST(rst), .I(in[555]), 
        .Q(round_reg[555]) );
  DFF \round_reg_reg[556]  ( .D(out[556]), .CLK(clk), .RST(rst), .I(in[556]), 
        .Q(round_reg[556]) );
  DFF \round_reg_reg[557]  ( .D(out[557]), .CLK(clk), .RST(rst), .I(in[557]), 
        .Q(round_reg[557]) );
  DFF \round_reg_reg[558]  ( .D(out[558]), .CLK(clk), .RST(rst), .I(in[558]), 
        .Q(round_reg[558]) );
  DFF \round_reg_reg[559]  ( .D(out[559]), .CLK(clk), .RST(rst), .I(in[559]), 
        .Q(round_reg[559]) );
  DFF \round_reg_reg[560]  ( .D(out[560]), .CLK(clk), .RST(rst), .I(in[560]), 
        .Q(round_reg[560]) );
  DFF \round_reg_reg[561]  ( .D(out[561]), .CLK(clk), .RST(rst), .I(in[561]), 
        .Q(round_reg[561]) );
  DFF \round_reg_reg[562]  ( .D(out[562]), .CLK(clk), .RST(rst), .I(in[562]), 
        .Q(round_reg[562]) );
  DFF \round_reg_reg[563]  ( .D(out[563]), .CLK(clk), .RST(rst), .I(in[563]), 
        .Q(round_reg[563]) );
  DFF \round_reg_reg[564]  ( .D(out[564]), .CLK(clk), .RST(rst), .I(in[564]), 
        .Q(round_reg[564]) );
  DFF \round_reg_reg[565]  ( .D(out[565]), .CLK(clk), .RST(rst), .I(in[565]), 
        .Q(round_reg[565]) );
  DFF \round_reg_reg[566]  ( .D(out[566]), .CLK(clk), .RST(rst), .I(in[566]), 
        .Q(round_reg[566]) );
  DFF \round_reg_reg[567]  ( .D(out[567]), .CLK(clk), .RST(rst), .I(in[567]), 
        .Q(round_reg[567]) );
  DFF \round_reg_reg[568]  ( .D(out[568]), .CLK(clk), .RST(rst), .I(in[568]), 
        .Q(round_reg[568]) );
  DFF \round_reg_reg[569]  ( .D(out[569]), .CLK(clk), .RST(rst), .I(in[569]), 
        .Q(round_reg[569]) );
  DFF \round_reg_reg[570]  ( .D(out[570]), .CLK(clk), .RST(rst), .I(in[570]), 
        .Q(round_reg[570]) );
  DFF \round_reg_reg[571]  ( .D(out[571]), .CLK(clk), .RST(rst), .I(in[571]), 
        .Q(round_reg[571]) );
  DFF \round_reg_reg[572]  ( .D(out[572]), .CLK(clk), .RST(rst), .I(in[572]), 
        .Q(round_reg[572]) );
  DFF \round_reg_reg[573]  ( .D(out[573]), .CLK(clk), .RST(rst), .I(in[573]), 
        .Q(round_reg[573]) );
  DFF \round_reg_reg[574]  ( .D(out[574]), .CLK(clk), .RST(rst), .I(in[574]), 
        .Q(round_reg[574]) );
  DFF \round_reg_reg[575]  ( .D(out[575]), .CLK(clk), .RST(rst), .I(in[575]), 
        .Q(round_reg[575]) );
  DFF \round_reg_reg[576]  ( .D(out[576]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[576]) );
  DFF \round_reg_reg[577]  ( .D(out[577]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[577]) );
  DFF \round_reg_reg[578]  ( .D(out[578]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[578]) );
  DFF \round_reg_reg[579]  ( .D(out[579]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[579]) );
  DFF \round_reg_reg[580]  ( .D(out[580]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[580]) );
  DFF \round_reg_reg[581]  ( .D(out[581]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[581]) );
  DFF \round_reg_reg[582]  ( .D(out[582]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[582]) );
  DFF \round_reg_reg[583]  ( .D(out[583]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[583]) );
  DFF \round_reg_reg[584]  ( .D(out[584]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[584]) );
  DFF \round_reg_reg[585]  ( .D(out[585]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[585]) );
  DFF \round_reg_reg[586]  ( .D(out[586]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[586]) );
  DFF \round_reg_reg[587]  ( .D(out[587]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[587]) );
  DFF \round_reg_reg[588]  ( .D(out[588]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[588]) );
  DFF \round_reg_reg[589]  ( .D(out[589]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[589]) );
  DFF \round_reg_reg[590]  ( .D(out[590]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[590]) );
  DFF \round_reg_reg[591]  ( .D(out[591]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[591]) );
  DFF \round_reg_reg[592]  ( .D(out[592]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[592]) );
  DFF \round_reg_reg[593]  ( .D(out[593]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[593]) );
  DFF \round_reg_reg[594]  ( .D(out[594]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[594]) );
  DFF \round_reg_reg[595]  ( .D(out[595]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[595]) );
  DFF \round_reg_reg[596]  ( .D(out[596]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[596]) );
  DFF \round_reg_reg[597]  ( .D(out[597]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[597]) );
  DFF \round_reg_reg[598]  ( .D(out[598]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[598]) );
  DFF \round_reg_reg[599]  ( .D(out[599]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[599]) );
  DFF \round_reg_reg[600]  ( .D(out[600]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[600]) );
  DFF \round_reg_reg[601]  ( .D(out[601]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[601]) );
  DFF \round_reg_reg[602]  ( .D(out[602]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[602]) );
  DFF \round_reg_reg[603]  ( .D(out[603]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[603]) );
  DFF \round_reg_reg[604]  ( .D(out[604]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[604]) );
  DFF \round_reg_reg[605]  ( .D(out[605]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[605]) );
  DFF \round_reg_reg[606]  ( .D(out[606]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[606]) );
  DFF \round_reg_reg[607]  ( .D(out[607]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[607]) );
  DFF \round_reg_reg[608]  ( .D(out[608]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[608]) );
  DFF \round_reg_reg[609]  ( .D(out[609]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[609]) );
  DFF \round_reg_reg[610]  ( .D(out[610]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[610]) );
  DFF \round_reg_reg[611]  ( .D(out[611]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[611]) );
  DFF \round_reg_reg[612]  ( .D(out[612]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[612]) );
  DFF \round_reg_reg[613]  ( .D(out[613]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[613]) );
  DFF \round_reg_reg[614]  ( .D(out[614]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[614]) );
  DFF \round_reg_reg[615]  ( .D(out[615]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[615]) );
  DFF \round_reg_reg[616]  ( .D(out[616]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[616]) );
  DFF \round_reg_reg[617]  ( .D(out[617]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[617]) );
  DFF \round_reg_reg[618]  ( .D(out[618]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[618]) );
  DFF \round_reg_reg[619]  ( .D(out[619]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[619]) );
  DFF \round_reg_reg[620]  ( .D(out[620]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[620]) );
  DFF \round_reg_reg[621]  ( .D(out[621]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[621]) );
  DFF \round_reg_reg[622]  ( .D(out[622]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[622]) );
  DFF \round_reg_reg[623]  ( .D(out[623]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[623]) );
  DFF \round_reg_reg[624]  ( .D(out[624]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[624]) );
  DFF \round_reg_reg[625]  ( .D(out[625]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[625]) );
  DFF \round_reg_reg[626]  ( .D(out[626]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[626]) );
  DFF \round_reg_reg[627]  ( .D(out[627]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[627]) );
  DFF \round_reg_reg[628]  ( .D(out[628]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[628]) );
  DFF \round_reg_reg[629]  ( .D(out[629]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[629]) );
  DFF \round_reg_reg[630]  ( .D(out[630]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[630]) );
  DFF \round_reg_reg[631]  ( .D(out[631]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[631]) );
  DFF \round_reg_reg[632]  ( .D(out[632]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[632]) );
  DFF \round_reg_reg[633]  ( .D(out[633]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[633]) );
  DFF \round_reg_reg[634]  ( .D(out[634]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[634]) );
  DFF \round_reg_reg[635]  ( .D(out[635]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[635]) );
  DFF \round_reg_reg[636]  ( .D(out[636]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[636]) );
  DFF \round_reg_reg[637]  ( .D(out[637]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[637]) );
  DFF \round_reg_reg[638]  ( .D(out[638]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[638]) );
  DFF \round_reg_reg[639]  ( .D(out[639]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[639]) );
  DFF \round_reg_reg[640]  ( .D(out[640]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[640]) );
  DFF \round_reg_reg[641]  ( .D(out[641]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[641]) );
  DFF \round_reg_reg[642]  ( .D(out[642]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[642]) );
  DFF \round_reg_reg[643]  ( .D(out[643]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[643]) );
  DFF \round_reg_reg[644]  ( .D(out[644]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[644]) );
  DFF \round_reg_reg[645]  ( .D(out[645]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[645]) );
  DFF \round_reg_reg[646]  ( .D(out[646]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[646]) );
  DFF \round_reg_reg[647]  ( .D(out[647]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[647]) );
  DFF \round_reg_reg[648]  ( .D(out[648]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[648]) );
  DFF \round_reg_reg[649]  ( .D(out[649]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[649]) );
  DFF \round_reg_reg[650]  ( .D(out[650]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[650]) );
  DFF \round_reg_reg[651]  ( .D(out[651]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[651]) );
  DFF \round_reg_reg[652]  ( .D(out[652]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[652]) );
  DFF \round_reg_reg[653]  ( .D(out[653]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[653]) );
  DFF \round_reg_reg[654]  ( .D(out[654]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[654]) );
  DFF \round_reg_reg[655]  ( .D(out[655]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[655]) );
  DFF \round_reg_reg[656]  ( .D(out[656]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[656]) );
  DFF \round_reg_reg[657]  ( .D(out[657]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[657]) );
  DFF \round_reg_reg[658]  ( .D(out[658]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[658]) );
  DFF \round_reg_reg[659]  ( .D(out[659]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[659]) );
  DFF \round_reg_reg[660]  ( .D(out[660]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[660]) );
  DFF \round_reg_reg[661]  ( .D(out[661]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[661]) );
  DFF \round_reg_reg[662]  ( .D(out[662]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[662]) );
  DFF \round_reg_reg[663]  ( .D(out[663]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[663]) );
  DFF \round_reg_reg[664]  ( .D(out[664]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[664]) );
  DFF \round_reg_reg[665]  ( .D(out[665]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[665]) );
  DFF \round_reg_reg[666]  ( .D(out[666]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[666]) );
  DFF \round_reg_reg[667]  ( .D(out[667]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[667]) );
  DFF \round_reg_reg[668]  ( .D(out[668]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[668]) );
  DFF \round_reg_reg[669]  ( .D(out[669]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[669]) );
  DFF \round_reg_reg[670]  ( .D(out[670]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[670]) );
  DFF \round_reg_reg[671]  ( .D(out[671]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[671]) );
  DFF \round_reg_reg[672]  ( .D(out[672]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[672]) );
  DFF \round_reg_reg[673]  ( .D(out[673]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[673]) );
  DFF \round_reg_reg[674]  ( .D(out[674]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[674]) );
  DFF \round_reg_reg[675]  ( .D(out[675]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[675]) );
  DFF \round_reg_reg[676]  ( .D(out[676]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[676]) );
  DFF \round_reg_reg[677]  ( .D(out[677]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[677]) );
  DFF \round_reg_reg[678]  ( .D(out[678]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[678]) );
  DFF \round_reg_reg[679]  ( .D(out[679]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[679]) );
  DFF \round_reg_reg[680]  ( .D(out[680]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[680]) );
  DFF \round_reg_reg[681]  ( .D(out[681]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[681]) );
  DFF \round_reg_reg[682]  ( .D(out[682]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[682]) );
  DFF \round_reg_reg[683]  ( .D(out[683]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[683]) );
  DFF \round_reg_reg[684]  ( .D(out[684]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[684]) );
  DFF \round_reg_reg[685]  ( .D(out[685]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[685]) );
  DFF \round_reg_reg[686]  ( .D(out[686]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[686]) );
  DFF \round_reg_reg[687]  ( .D(out[687]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[687]) );
  DFF \round_reg_reg[688]  ( .D(out[688]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[688]) );
  DFF \round_reg_reg[689]  ( .D(out[689]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[689]) );
  DFF \round_reg_reg[690]  ( .D(out[690]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[690]) );
  DFF \round_reg_reg[691]  ( .D(out[691]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[691]) );
  DFF \round_reg_reg[692]  ( .D(out[692]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[692]) );
  DFF \round_reg_reg[693]  ( .D(out[693]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[693]) );
  DFF \round_reg_reg[694]  ( .D(out[694]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[694]) );
  DFF \round_reg_reg[695]  ( .D(out[695]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[695]) );
  DFF \round_reg_reg[696]  ( .D(out[696]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[696]) );
  DFF \round_reg_reg[697]  ( .D(out[697]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[697]) );
  DFF \round_reg_reg[698]  ( .D(out[698]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[698]) );
  DFF \round_reg_reg[699]  ( .D(out[699]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[699]) );
  DFF \round_reg_reg[700]  ( .D(out[700]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[700]) );
  DFF \round_reg_reg[701]  ( .D(out[701]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[701]) );
  DFF \round_reg_reg[702]  ( .D(out[702]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[702]) );
  DFF \round_reg_reg[703]  ( .D(out[703]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[703]) );
  DFF \round_reg_reg[704]  ( .D(out[704]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[704]) );
  DFF \round_reg_reg[705]  ( .D(out[705]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[705]) );
  DFF \round_reg_reg[706]  ( .D(out[706]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[706]) );
  DFF \round_reg_reg[707]  ( .D(out[707]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[707]) );
  DFF \round_reg_reg[708]  ( .D(out[708]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[708]) );
  DFF \round_reg_reg[709]  ( .D(out[709]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[709]) );
  DFF \round_reg_reg[710]  ( .D(out[710]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[710]) );
  DFF \round_reg_reg[711]  ( .D(out[711]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[711]) );
  DFF \round_reg_reg[712]  ( .D(out[712]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[712]) );
  DFF \round_reg_reg[713]  ( .D(out[713]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[713]) );
  DFF \round_reg_reg[714]  ( .D(out[714]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[714]) );
  DFF \round_reg_reg[715]  ( .D(out[715]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[715]) );
  DFF \round_reg_reg[716]  ( .D(out[716]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[716]) );
  DFF \round_reg_reg[717]  ( .D(out[717]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[717]) );
  DFF \round_reg_reg[718]  ( .D(out[718]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[718]) );
  DFF \round_reg_reg[719]  ( .D(out[719]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[719]) );
  DFF \round_reg_reg[720]  ( .D(out[720]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[720]) );
  DFF \round_reg_reg[721]  ( .D(out[721]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[721]) );
  DFF \round_reg_reg[722]  ( .D(out[722]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[722]) );
  DFF \round_reg_reg[723]  ( .D(out[723]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[723]) );
  DFF \round_reg_reg[724]  ( .D(out[724]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[724]) );
  DFF \round_reg_reg[725]  ( .D(out[725]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[725]) );
  DFF \round_reg_reg[726]  ( .D(out[726]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[726]) );
  DFF \round_reg_reg[727]  ( .D(out[727]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[727]) );
  DFF \round_reg_reg[728]  ( .D(out[728]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[728]) );
  DFF \round_reg_reg[729]  ( .D(out[729]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[729]) );
  DFF \round_reg_reg[730]  ( .D(out[730]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[730]) );
  DFF \round_reg_reg[731]  ( .D(out[731]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[731]) );
  DFF \round_reg_reg[732]  ( .D(out[732]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[732]) );
  DFF \round_reg_reg[733]  ( .D(out[733]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[733]) );
  DFF \round_reg_reg[734]  ( .D(out[734]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[734]) );
  DFF \round_reg_reg[735]  ( .D(out[735]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[735]) );
  DFF \round_reg_reg[736]  ( .D(out[736]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[736]) );
  DFF \round_reg_reg[737]  ( .D(out[737]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[737]) );
  DFF \round_reg_reg[738]  ( .D(out[738]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[738]) );
  DFF \round_reg_reg[739]  ( .D(out[739]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[739]) );
  DFF \round_reg_reg[740]  ( .D(out[740]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[740]) );
  DFF \round_reg_reg[741]  ( .D(out[741]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[741]) );
  DFF \round_reg_reg[742]  ( .D(out[742]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[742]) );
  DFF \round_reg_reg[743]  ( .D(out[743]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[743]) );
  DFF \round_reg_reg[744]  ( .D(out[744]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[744]) );
  DFF \round_reg_reg[745]  ( .D(out[745]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[745]) );
  DFF \round_reg_reg[746]  ( .D(out[746]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[746]) );
  DFF \round_reg_reg[747]  ( .D(out[747]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[747]) );
  DFF \round_reg_reg[748]  ( .D(out[748]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[748]) );
  DFF \round_reg_reg[749]  ( .D(out[749]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[749]) );
  DFF \round_reg_reg[750]  ( .D(out[750]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[750]) );
  DFF \round_reg_reg[751]  ( .D(out[751]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[751]) );
  DFF \round_reg_reg[752]  ( .D(out[752]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[752]) );
  DFF \round_reg_reg[753]  ( .D(out[753]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[753]) );
  DFF \round_reg_reg[754]  ( .D(out[754]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[754]) );
  DFF \round_reg_reg[755]  ( .D(out[755]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[755]) );
  DFF \round_reg_reg[756]  ( .D(out[756]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[756]) );
  DFF \round_reg_reg[757]  ( .D(out[757]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[757]) );
  DFF \round_reg_reg[758]  ( .D(out[758]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[758]) );
  DFF \round_reg_reg[759]  ( .D(out[759]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[759]) );
  DFF \round_reg_reg[760]  ( .D(out[760]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[760]) );
  DFF \round_reg_reg[761]  ( .D(out[761]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[761]) );
  DFF \round_reg_reg[762]  ( .D(out[762]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[762]) );
  DFF \round_reg_reg[763]  ( .D(out[763]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[763]) );
  DFF \round_reg_reg[764]  ( .D(out[764]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[764]) );
  DFF \round_reg_reg[765]  ( .D(out[765]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[765]) );
  DFF \round_reg_reg[766]  ( .D(out[766]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[766]) );
  DFF \round_reg_reg[767]  ( .D(out[767]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[767]) );
  DFF \round_reg_reg[768]  ( .D(out[768]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[768]) );
  DFF \round_reg_reg[769]  ( .D(out[769]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[769]) );
  DFF \round_reg_reg[770]  ( .D(out[770]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[770]) );
  DFF \round_reg_reg[771]  ( .D(out[771]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[771]) );
  DFF \round_reg_reg[772]  ( .D(out[772]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[772]) );
  DFF \round_reg_reg[773]  ( .D(out[773]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[773]) );
  DFF \round_reg_reg[774]  ( .D(out[774]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[774]) );
  DFF \round_reg_reg[775]  ( .D(out[775]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[775]) );
  DFF \round_reg_reg[776]  ( .D(out[776]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[776]) );
  DFF \round_reg_reg[777]  ( .D(out[777]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[777]) );
  DFF \round_reg_reg[778]  ( .D(out[778]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[778]) );
  DFF \round_reg_reg[779]  ( .D(out[779]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[779]) );
  DFF \round_reg_reg[780]  ( .D(out[780]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[780]) );
  DFF \round_reg_reg[781]  ( .D(out[781]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[781]) );
  DFF \round_reg_reg[782]  ( .D(out[782]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[782]) );
  DFF \round_reg_reg[783]  ( .D(out[783]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[783]) );
  DFF \round_reg_reg[784]  ( .D(out[784]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[784]) );
  DFF \round_reg_reg[785]  ( .D(out[785]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[785]) );
  DFF \round_reg_reg[786]  ( .D(out[786]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[786]) );
  DFF \round_reg_reg[787]  ( .D(out[787]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[787]) );
  DFF \round_reg_reg[788]  ( .D(out[788]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[788]) );
  DFF \round_reg_reg[789]  ( .D(out[789]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[789]) );
  DFF \round_reg_reg[790]  ( .D(out[790]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[790]) );
  DFF \round_reg_reg[791]  ( .D(out[791]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[791]) );
  DFF \round_reg_reg[792]  ( .D(out[792]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[792]) );
  DFF \round_reg_reg[793]  ( .D(out[793]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[793]) );
  DFF \round_reg_reg[794]  ( .D(out[794]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[794]) );
  DFF \round_reg_reg[795]  ( .D(out[795]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[795]) );
  DFF \round_reg_reg[796]  ( .D(out[796]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[796]) );
  DFF \round_reg_reg[797]  ( .D(out[797]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[797]) );
  DFF \round_reg_reg[798]  ( .D(out[798]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[798]) );
  DFF \round_reg_reg[799]  ( .D(out[799]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[799]) );
  DFF \round_reg_reg[800]  ( .D(out[800]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[800]) );
  DFF \round_reg_reg[801]  ( .D(out[801]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[801]) );
  DFF \round_reg_reg[802]  ( .D(out[802]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[802]) );
  DFF \round_reg_reg[803]  ( .D(out[803]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[803]) );
  DFF \round_reg_reg[804]  ( .D(out[804]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[804]) );
  DFF \round_reg_reg[805]  ( .D(out[805]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[805]) );
  DFF \round_reg_reg[806]  ( .D(out[806]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[806]) );
  DFF \round_reg_reg[807]  ( .D(out[807]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[807]) );
  DFF \round_reg_reg[808]  ( .D(out[808]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[808]) );
  DFF \round_reg_reg[809]  ( .D(out[809]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[809]) );
  DFF \round_reg_reg[810]  ( .D(out[810]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[810]) );
  DFF \round_reg_reg[811]  ( .D(out[811]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[811]) );
  DFF \round_reg_reg[812]  ( .D(out[812]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[812]) );
  DFF \round_reg_reg[813]  ( .D(out[813]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[813]) );
  DFF \round_reg_reg[814]  ( .D(out[814]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[814]) );
  DFF \round_reg_reg[815]  ( .D(out[815]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[815]) );
  DFF \round_reg_reg[816]  ( .D(out[816]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[816]) );
  DFF \round_reg_reg[817]  ( .D(out[817]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[817]) );
  DFF \round_reg_reg[818]  ( .D(out[818]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[818]) );
  DFF \round_reg_reg[819]  ( .D(out[819]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[819]) );
  DFF \round_reg_reg[820]  ( .D(out[820]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[820]) );
  DFF \round_reg_reg[821]  ( .D(out[821]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[821]) );
  DFF \round_reg_reg[822]  ( .D(out[822]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[822]) );
  DFF \round_reg_reg[823]  ( .D(out[823]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[823]) );
  DFF \round_reg_reg[824]  ( .D(out[824]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[824]) );
  DFF \round_reg_reg[825]  ( .D(out[825]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[825]) );
  DFF \round_reg_reg[826]  ( .D(out[826]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[826]) );
  DFF \round_reg_reg[827]  ( .D(out[827]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[827]) );
  DFF \round_reg_reg[828]  ( .D(out[828]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[828]) );
  DFF \round_reg_reg[829]  ( .D(out[829]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[829]) );
  DFF \round_reg_reg[830]  ( .D(out[830]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[830]) );
  DFF \round_reg_reg[831]  ( .D(out[831]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[831]) );
  DFF \round_reg_reg[832]  ( .D(out[832]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[832]) );
  DFF \round_reg_reg[833]  ( .D(out[833]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[833]) );
  DFF \round_reg_reg[834]  ( .D(out[834]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[834]) );
  DFF \round_reg_reg[835]  ( .D(out[835]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[835]) );
  DFF \round_reg_reg[836]  ( .D(out[836]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[836]) );
  DFF \round_reg_reg[837]  ( .D(out[837]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[837]) );
  DFF \round_reg_reg[838]  ( .D(out[838]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[838]) );
  DFF \round_reg_reg[839]  ( .D(out[839]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[839]) );
  DFF \round_reg_reg[840]  ( .D(out[840]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[840]) );
  DFF \round_reg_reg[841]  ( .D(out[841]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[841]) );
  DFF \round_reg_reg[842]  ( .D(out[842]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[842]) );
  DFF \round_reg_reg[843]  ( .D(out[843]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[843]) );
  DFF \round_reg_reg[844]  ( .D(out[844]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[844]) );
  DFF \round_reg_reg[845]  ( .D(out[845]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[845]) );
  DFF \round_reg_reg[846]  ( .D(out[846]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[846]) );
  DFF \round_reg_reg[847]  ( .D(out[847]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[847]) );
  DFF \round_reg_reg[848]  ( .D(out[848]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[848]) );
  DFF \round_reg_reg[849]  ( .D(out[849]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[849]) );
  DFF \round_reg_reg[850]  ( .D(out[850]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[850]) );
  DFF \round_reg_reg[851]  ( .D(out[851]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[851]) );
  DFF \round_reg_reg[852]  ( .D(out[852]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[852]) );
  DFF \round_reg_reg[853]  ( .D(out[853]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[853]) );
  DFF \round_reg_reg[854]  ( .D(out[854]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[854]) );
  DFF \round_reg_reg[855]  ( .D(out[855]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[855]) );
  DFF \round_reg_reg[856]  ( .D(out[856]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[856]) );
  DFF \round_reg_reg[857]  ( .D(out[857]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[857]) );
  DFF \round_reg_reg[858]  ( .D(out[858]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[858]) );
  DFF \round_reg_reg[859]  ( .D(out[859]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[859]) );
  DFF \round_reg_reg[860]  ( .D(out[860]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[860]) );
  DFF \round_reg_reg[861]  ( .D(out[861]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[861]) );
  DFF \round_reg_reg[862]  ( .D(out[862]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[862]) );
  DFF \round_reg_reg[863]  ( .D(out[863]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[863]) );
  DFF \round_reg_reg[864]  ( .D(out[864]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[864]) );
  DFF \round_reg_reg[865]  ( .D(out[865]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[865]) );
  DFF \round_reg_reg[866]  ( .D(out[866]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[866]) );
  DFF \round_reg_reg[867]  ( .D(out[867]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[867]) );
  DFF \round_reg_reg[868]  ( .D(out[868]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[868]) );
  DFF \round_reg_reg[869]  ( .D(out[869]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[869]) );
  DFF \round_reg_reg[870]  ( .D(out[870]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[870]) );
  DFF \round_reg_reg[871]  ( .D(out[871]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[871]) );
  DFF \round_reg_reg[872]  ( .D(out[872]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[872]) );
  DFF \round_reg_reg[873]  ( .D(out[873]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[873]) );
  DFF \round_reg_reg[874]  ( .D(out[874]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[874]) );
  DFF \round_reg_reg[875]  ( .D(out[875]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[875]) );
  DFF \round_reg_reg[876]  ( .D(out[876]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[876]) );
  DFF \round_reg_reg[877]  ( .D(out[877]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[877]) );
  DFF \round_reg_reg[878]  ( .D(out[878]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[878]) );
  DFF \round_reg_reg[879]  ( .D(out[879]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[879]) );
  DFF \round_reg_reg[880]  ( .D(out[880]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[880]) );
  DFF \round_reg_reg[881]  ( .D(out[881]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[881]) );
  DFF \round_reg_reg[882]  ( .D(out[882]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[882]) );
  DFF \round_reg_reg[883]  ( .D(out[883]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[883]) );
  DFF \round_reg_reg[884]  ( .D(out[884]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[884]) );
  DFF \round_reg_reg[885]  ( .D(out[885]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[885]) );
  DFF \round_reg_reg[886]  ( .D(out[886]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[886]) );
  DFF \round_reg_reg[887]  ( .D(out[887]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[887]) );
  DFF \round_reg_reg[888]  ( .D(out[888]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[888]) );
  DFF \round_reg_reg[889]  ( .D(out[889]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[889]) );
  DFF \round_reg_reg[890]  ( .D(out[890]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[890]) );
  DFF \round_reg_reg[891]  ( .D(out[891]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[891]) );
  DFF \round_reg_reg[892]  ( .D(out[892]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[892]) );
  DFF \round_reg_reg[893]  ( .D(out[893]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[893]) );
  DFF \round_reg_reg[894]  ( .D(out[894]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[894]) );
  DFF \round_reg_reg[895]  ( .D(out[895]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[895]) );
  DFF \round_reg_reg[896]  ( .D(out[896]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[896]) );
  DFF \round_reg_reg[897]  ( .D(out[897]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[897]) );
  DFF \round_reg_reg[898]  ( .D(out[898]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[898]) );
  DFF \round_reg_reg[899]  ( .D(out[899]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[899]) );
  DFF \round_reg_reg[900]  ( .D(out[900]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[900]) );
  DFF \round_reg_reg[901]  ( .D(out[901]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[901]) );
  DFF \round_reg_reg[902]  ( .D(out[902]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[902]) );
  DFF \round_reg_reg[903]  ( .D(out[903]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[903]) );
  DFF \round_reg_reg[904]  ( .D(out[904]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[904]) );
  DFF \round_reg_reg[905]  ( .D(out[905]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[905]) );
  DFF \round_reg_reg[906]  ( .D(out[906]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[906]) );
  DFF \round_reg_reg[907]  ( .D(out[907]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[907]) );
  DFF \round_reg_reg[908]  ( .D(out[908]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[908]) );
  DFF \round_reg_reg[909]  ( .D(out[909]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[909]) );
  DFF \round_reg_reg[910]  ( .D(out[910]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[910]) );
  DFF \round_reg_reg[911]  ( .D(out[911]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[911]) );
  DFF \round_reg_reg[912]  ( .D(out[912]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[912]) );
  DFF \round_reg_reg[913]  ( .D(out[913]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[913]) );
  DFF \round_reg_reg[914]  ( .D(out[914]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[914]) );
  DFF \round_reg_reg[915]  ( .D(out[915]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[915]) );
  DFF \round_reg_reg[916]  ( .D(out[916]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[916]) );
  DFF \round_reg_reg[917]  ( .D(out[917]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[917]) );
  DFF \round_reg_reg[918]  ( .D(out[918]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[918]) );
  DFF \round_reg_reg[919]  ( .D(out[919]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[919]) );
  DFF \round_reg_reg[920]  ( .D(out[920]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[920]) );
  DFF \round_reg_reg[921]  ( .D(out[921]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[921]) );
  DFF \round_reg_reg[922]  ( .D(out[922]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[922]) );
  DFF \round_reg_reg[923]  ( .D(out[923]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[923]) );
  DFF \round_reg_reg[924]  ( .D(out[924]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[924]) );
  DFF \round_reg_reg[925]  ( .D(out[925]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[925]) );
  DFF \round_reg_reg[926]  ( .D(out[926]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[926]) );
  DFF \round_reg_reg[927]  ( .D(out[927]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[927]) );
  DFF \round_reg_reg[928]  ( .D(out[928]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[928]) );
  DFF \round_reg_reg[929]  ( .D(out[929]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[929]) );
  DFF \round_reg_reg[930]  ( .D(out[930]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[930]) );
  DFF \round_reg_reg[931]  ( .D(out[931]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[931]) );
  DFF \round_reg_reg[932]  ( .D(out[932]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[932]) );
  DFF \round_reg_reg[933]  ( .D(out[933]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[933]) );
  DFF \round_reg_reg[934]  ( .D(out[934]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[934]) );
  DFF \round_reg_reg[935]  ( .D(out[935]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[935]) );
  DFF \round_reg_reg[936]  ( .D(out[936]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[936]) );
  DFF \round_reg_reg[937]  ( .D(out[937]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[937]) );
  DFF \round_reg_reg[938]  ( .D(out[938]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[938]) );
  DFF \round_reg_reg[939]  ( .D(out[939]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[939]) );
  DFF \round_reg_reg[940]  ( .D(out[940]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[940]) );
  DFF \round_reg_reg[941]  ( .D(out[941]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[941]) );
  DFF \round_reg_reg[942]  ( .D(out[942]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[942]) );
  DFF \round_reg_reg[943]  ( .D(out[943]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[943]) );
  DFF \round_reg_reg[944]  ( .D(out[944]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[944]) );
  DFF \round_reg_reg[945]  ( .D(out[945]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[945]) );
  DFF \round_reg_reg[946]  ( .D(out[946]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[946]) );
  DFF \round_reg_reg[947]  ( .D(out[947]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[947]) );
  DFF \round_reg_reg[948]  ( .D(out[948]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[948]) );
  DFF \round_reg_reg[949]  ( .D(out[949]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[949]) );
  DFF \round_reg_reg[950]  ( .D(out[950]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[950]) );
  DFF \round_reg_reg[951]  ( .D(out[951]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[951]) );
  DFF \round_reg_reg[952]  ( .D(out[952]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[952]) );
  DFF \round_reg_reg[953]  ( .D(out[953]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[953]) );
  DFF \round_reg_reg[954]  ( .D(out[954]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[954]) );
  DFF \round_reg_reg[955]  ( .D(out[955]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[955]) );
  DFF \round_reg_reg[956]  ( .D(out[956]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[956]) );
  DFF \round_reg_reg[957]  ( .D(out[957]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[957]) );
  DFF \round_reg_reg[958]  ( .D(out[958]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[958]) );
  DFF \round_reg_reg[959]  ( .D(out[959]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[959]) );
  DFF \round_reg_reg[960]  ( .D(out[960]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[960]) );
  DFF \round_reg_reg[961]  ( .D(out[961]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[961]) );
  DFF \round_reg_reg[962]  ( .D(out[962]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[962]) );
  DFF \round_reg_reg[963]  ( .D(out[963]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[963]) );
  DFF \round_reg_reg[964]  ( .D(out[964]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[964]) );
  DFF \round_reg_reg[965]  ( .D(out[965]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[965]) );
  DFF \round_reg_reg[966]  ( .D(out[966]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[966]) );
  DFF \round_reg_reg[967]  ( .D(out[967]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[967]) );
  DFF \round_reg_reg[968]  ( .D(out[968]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[968]) );
  DFF \round_reg_reg[969]  ( .D(out[969]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[969]) );
  DFF \round_reg_reg[970]  ( .D(out[970]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[970]) );
  DFF \round_reg_reg[971]  ( .D(out[971]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[971]) );
  DFF \round_reg_reg[972]  ( .D(out[972]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[972]) );
  DFF \round_reg_reg[973]  ( .D(out[973]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[973]) );
  DFF \round_reg_reg[974]  ( .D(out[974]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[974]) );
  DFF \round_reg_reg[975]  ( .D(out[975]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[975]) );
  DFF \round_reg_reg[976]  ( .D(out[976]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[976]) );
  DFF \round_reg_reg[977]  ( .D(out[977]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[977]) );
  DFF \round_reg_reg[978]  ( .D(out[978]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[978]) );
  DFF \round_reg_reg[979]  ( .D(out[979]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[979]) );
  DFF \round_reg_reg[980]  ( .D(out[980]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[980]) );
  DFF \round_reg_reg[981]  ( .D(out[981]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[981]) );
  DFF \round_reg_reg[982]  ( .D(out[982]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[982]) );
  DFF \round_reg_reg[983]  ( .D(out[983]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[983]) );
  DFF \round_reg_reg[984]  ( .D(out[984]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[984]) );
  DFF \round_reg_reg[985]  ( .D(out[985]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[985]) );
  DFF \round_reg_reg[986]  ( .D(out[986]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[986]) );
  DFF \round_reg_reg[987]  ( .D(out[987]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[987]) );
  DFF \round_reg_reg[988]  ( .D(out[988]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[988]) );
  DFF \round_reg_reg[989]  ( .D(out[989]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[989]) );
  DFF \round_reg_reg[990]  ( .D(out[990]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[990]) );
  DFF \round_reg_reg[991]  ( .D(out[991]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[991]) );
  DFF \round_reg_reg[992]  ( .D(out[992]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[992]) );
  DFF \round_reg_reg[993]  ( .D(out[993]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[993]) );
  DFF \round_reg_reg[994]  ( .D(out[994]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[994]) );
  DFF \round_reg_reg[995]  ( .D(out[995]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[995]) );
  DFF \round_reg_reg[996]  ( .D(out[996]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[996]) );
  DFF \round_reg_reg[997]  ( .D(out[997]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[997]) );
  DFF \round_reg_reg[998]  ( .D(out[998]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[998]) );
  DFF \round_reg_reg[999]  ( .D(out[999]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[999]) );
  DFF \round_reg_reg[1000]  ( .D(out[1000]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1000]) );
  DFF \round_reg_reg[1001]  ( .D(out[1001]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1001]) );
  DFF \round_reg_reg[1002]  ( .D(out[1002]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1002]) );
  DFF \round_reg_reg[1003]  ( .D(out[1003]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1003]) );
  DFF \round_reg_reg[1004]  ( .D(out[1004]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1004]) );
  DFF \round_reg_reg[1005]  ( .D(out[1005]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1005]) );
  DFF \round_reg_reg[1006]  ( .D(out[1006]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1006]) );
  DFF \round_reg_reg[1007]  ( .D(out[1007]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1007]) );
  DFF \round_reg_reg[1008]  ( .D(out[1008]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1008]) );
  DFF \round_reg_reg[1009]  ( .D(out[1009]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1009]) );
  DFF \round_reg_reg[1010]  ( .D(out[1010]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1010]) );
  DFF \round_reg_reg[1011]  ( .D(out[1011]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1011]) );
  DFF \round_reg_reg[1012]  ( .D(out[1012]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1012]) );
  DFF \round_reg_reg[1013]  ( .D(out[1013]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1013]) );
  DFF \round_reg_reg[1014]  ( .D(out[1014]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1014]) );
  DFF \round_reg_reg[1015]  ( .D(out[1015]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1015]) );
  DFF \round_reg_reg[1016]  ( .D(out[1016]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1016]) );
  DFF \round_reg_reg[1017]  ( .D(out[1017]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1017]) );
  DFF \round_reg_reg[1018]  ( .D(out[1018]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1018]) );
  DFF \round_reg_reg[1019]  ( .D(out[1019]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1019]) );
  DFF \round_reg_reg[1020]  ( .D(out[1020]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1020]) );
  DFF \round_reg_reg[1021]  ( .D(out[1021]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1021]) );
  DFF \round_reg_reg[1022]  ( .D(out[1022]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1022]) );
  DFF \round_reg_reg[1023]  ( .D(out[1023]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1023]) );
  DFF \round_reg_reg[1024]  ( .D(out[1024]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1024]) );
  DFF \round_reg_reg[1025]  ( .D(out[1025]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1025]) );
  DFF \round_reg_reg[1026]  ( .D(out[1026]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1026]) );
  DFF \round_reg_reg[1027]  ( .D(out[1027]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1027]) );
  DFF \round_reg_reg[1028]  ( .D(out[1028]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1028]) );
  DFF \round_reg_reg[1029]  ( .D(out[1029]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1029]) );
  DFF \round_reg_reg[1030]  ( .D(out[1030]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1030]) );
  DFF \round_reg_reg[1031]  ( .D(out[1031]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1031]) );
  DFF \round_reg_reg[1032]  ( .D(out[1032]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1032]) );
  DFF \round_reg_reg[1033]  ( .D(out[1033]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1033]) );
  DFF \round_reg_reg[1034]  ( .D(out[1034]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1034]) );
  DFF \round_reg_reg[1035]  ( .D(out[1035]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1035]) );
  DFF \round_reg_reg[1036]  ( .D(out[1036]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1036]) );
  DFF \round_reg_reg[1037]  ( .D(out[1037]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1037]) );
  DFF \round_reg_reg[1038]  ( .D(out[1038]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1038]) );
  DFF \round_reg_reg[1039]  ( .D(out[1039]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1039]) );
  DFF \round_reg_reg[1040]  ( .D(out[1040]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1040]) );
  DFF \round_reg_reg[1041]  ( .D(out[1041]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1041]) );
  DFF \round_reg_reg[1042]  ( .D(out[1042]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1042]) );
  DFF \round_reg_reg[1043]  ( .D(out[1043]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1043]) );
  DFF \round_reg_reg[1044]  ( .D(out[1044]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1044]) );
  DFF \round_reg_reg[1045]  ( .D(out[1045]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1045]) );
  DFF \round_reg_reg[1046]  ( .D(out[1046]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1046]) );
  DFF \round_reg_reg[1047]  ( .D(out[1047]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1047]) );
  DFF \round_reg_reg[1048]  ( .D(out[1048]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1048]) );
  DFF \round_reg_reg[1049]  ( .D(out[1049]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1049]) );
  DFF \round_reg_reg[1050]  ( .D(out[1050]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1050]) );
  DFF \round_reg_reg[1051]  ( .D(out[1051]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1051]) );
  DFF \round_reg_reg[1052]  ( .D(out[1052]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1052]) );
  DFF \round_reg_reg[1053]  ( .D(out[1053]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1053]) );
  DFF \round_reg_reg[1054]  ( .D(out[1054]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1054]) );
  DFF \round_reg_reg[1055]  ( .D(out[1055]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1055]) );
  DFF \round_reg_reg[1056]  ( .D(out[1056]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1056]) );
  DFF \round_reg_reg[1057]  ( .D(out[1057]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1057]) );
  DFF \round_reg_reg[1058]  ( .D(out[1058]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1058]) );
  DFF \round_reg_reg[1059]  ( .D(out[1059]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1059]) );
  DFF \round_reg_reg[1060]  ( .D(out[1060]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1060]) );
  DFF \round_reg_reg[1061]  ( .D(out[1061]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1061]) );
  DFF \round_reg_reg[1062]  ( .D(out[1062]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1062]) );
  DFF \round_reg_reg[1063]  ( .D(out[1063]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1063]) );
  DFF \round_reg_reg[1064]  ( .D(out[1064]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1064]) );
  DFF \round_reg_reg[1065]  ( .D(out[1065]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1065]) );
  DFF \round_reg_reg[1066]  ( .D(out[1066]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1066]) );
  DFF \round_reg_reg[1067]  ( .D(out[1067]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1067]) );
  DFF \round_reg_reg[1068]  ( .D(out[1068]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1068]) );
  DFF \round_reg_reg[1069]  ( .D(out[1069]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1069]) );
  DFF \round_reg_reg[1070]  ( .D(out[1070]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1070]) );
  DFF \round_reg_reg[1071]  ( .D(out[1071]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1071]) );
  DFF \round_reg_reg[1072]  ( .D(out[1072]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1072]) );
  DFF \round_reg_reg[1073]  ( .D(out[1073]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1073]) );
  DFF \round_reg_reg[1074]  ( .D(out[1074]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1074]) );
  DFF \round_reg_reg[1075]  ( .D(out[1075]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1075]) );
  DFF \round_reg_reg[1076]  ( .D(out[1076]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1076]) );
  DFF \round_reg_reg[1077]  ( .D(out[1077]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1077]) );
  DFF \round_reg_reg[1078]  ( .D(out[1078]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1078]) );
  DFF \round_reg_reg[1079]  ( .D(out[1079]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1079]) );
  DFF \round_reg_reg[1080]  ( .D(out[1080]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1080]) );
  DFF \round_reg_reg[1081]  ( .D(out[1081]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1081]) );
  DFF \round_reg_reg[1082]  ( .D(out[1082]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1082]) );
  DFF \round_reg_reg[1083]  ( .D(out[1083]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1083]) );
  DFF \round_reg_reg[1084]  ( .D(out[1084]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1084]) );
  DFF \round_reg_reg[1085]  ( .D(out[1085]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1085]) );
  DFF \round_reg_reg[1086]  ( .D(out[1086]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1086]) );
  DFF \round_reg_reg[1087]  ( .D(out[1087]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1087]) );
  DFF \round_reg_reg[1088]  ( .D(out[1088]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1088]) );
  DFF \round_reg_reg[1089]  ( .D(out[1089]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1089]) );
  DFF \round_reg_reg[1090]  ( .D(out[1090]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1090]) );
  DFF \round_reg_reg[1091]  ( .D(out[1091]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1091]) );
  DFF \round_reg_reg[1092]  ( .D(out[1092]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1092]) );
  DFF \round_reg_reg[1093]  ( .D(out[1093]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1093]) );
  DFF \round_reg_reg[1094]  ( .D(out[1094]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1094]) );
  DFF \round_reg_reg[1095]  ( .D(out[1095]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1095]) );
  DFF \round_reg_reg[1096]  ( .D(out[1096]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1096]) );
  DFF \round_reg_reg[1097]  ( .D(out[1097]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1097]) );
  DFF \round_reg_reg[1098]  ( .D(out[1098]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1098]) );
  DFF \round_reg_reg[1099]  ( .D(out[1099]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1099]) );
  DFF \round_reg_reg[1100]  ( .D(out[1100]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1100]) );
  DFF \round_reg_reg[1101]  ( .D(out[1101]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1101]) );
  DFF \round_reg_reg[1102]  ( .D(out[1102]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1102]) );
  DFF \round_reg_reg[1103]  ( .D(out[1103]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1103]) );
  DFF \round_reg_reg[1104]  ( .D(out[1104]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1104]) );
  DFF \round_reg_reg[1105]  ( .D(out[1105]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1105]) );
  DFF \round_reg_reg[1106]  ( .D(out[1106]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1106]) );
  DFF \round_reg_reg[1107]  ( .D(out[1107]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1107]) );
  DFF \round_reg_reg[1108]  ( .D(out[1108]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1108]) );
  DFF \round_reg_reg[1109]  ( .D(out[1109]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1109]) );
  DFF \round_reg_reg[1110]  ( .D(out[1110]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1110]) );
  DFF \round_reg_reg[1111]  ( .D(out[1111]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1111]) );
  DFF \round_reg_reg[1112]  ( .D(out[1112]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1112]) );
  DFF \round_reg_reg[1113]  ( .D(out[1113]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1113]) );
  DFF \round_reg_reg[1114]  ( .D(out[1114]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1114]) );
  DFF \round_reg_reg[1115]  ( .D(out[1115]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1115]) );
  DFF \round_reg_reg[1116]  ( .D(out[1116]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1116]) );
  DFF \round_reg_reg[1117]  ( .D(out[1117]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1117]) );
  DFF \round_reg_reg[1118]  ( .D(out[1118]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1118]) );
  DFF \round_reg_reg[1119]  ( .D(out[1119]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1119]) );
  DFF \round_reg_reg[1120]  ( .D(out[1120]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1120]) );
  DFF \round_reg_reg[1121]  ( .D(out[1121]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1121]) );
  DFF \round_reg_reg[1122]  ( .D(out[1122]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1122]) );
  DFF \round_reg_reg[1123]  ( .D(out[1123]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1123]) );
  DFF \round_reg_reg[1124]  ( .D(out[1124]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1124]) );
  DFF \round_reg_reg[1125]  ( .D(out[1125]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1125]) );
  DFF \round_reg_reg[1126]  ( .D(out[1126]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1126]) );
  DFF \round_reg_reg[1127]  ( .D(out[1127]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1127]) );
  DFF \round_reg_reg[1128]  ( .D(out[1128]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1128]) );
  DFF \round_reg_reg[1129]  ( .D(out[1129]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1129]) );
  DFF \round_reg_reg[1130]  ( .D(out[1130]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1130]) );
  DFF \round_reg_reg[1131]  ( .D(out[1131]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1131]) );
  DFF \round_reg_reg[1132]  ( .D(out[1132]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1132]) );
  DFF \round_reg_reg[1133]  ( .D(out[1133]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1133]) );
  DFF \round_reg_reg[1134]  ( .D(out[1134]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1134]) );
  DFF \round_reg_reg[1135]  ( .D(out[1135]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1135]) );
  DFF \round_reg_reg[1136]  ( .D(out[1136]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1136]) );
  DFF \round_reg_reg[1137]  ( .D(out[1137]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1137]) );
  DFF \round_reg_reg[1138]  ( .D(out[1138]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1138]) );
  DFF \round_reg_reg[1139]  ( .D(out[1139]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1139]) );
  DFF \round_reg_reg[1140]  ( .D(out[1140]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1140]) );
  DFF \round_reg_reg[1141]  ( .D(out[1141]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1141]) );
  DFF \round_reg_reg[1142]  ( .D(out[1142]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1142]) );
  DFF \round_reg_reg[1143]  ( .D(out[1143]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1143]) );
  DFF \round_reg_reg[1144]  ( .D(out[1144]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1144]) );
  DFF \round_reg_reg[1145]  ( .D(out[1145]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1145]) );
  DFF \round_reg_reg[1146]  ( .D(out[1146]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1146]) );
  DFF \round_reg_reg[1147]  ( .D(out[1147]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1147]) );
  DFF \round_reg_reg[1148]  ( .D(out[1148]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1148]) );
  DFF \round_reg_reg[1149]  ( .D(out[1149]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1149]) );
  DFF \round_reg_reg[1150]  ( .D(out[1150]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1150]) );
  DFF \round_reg_reg[1151]  ( .D(out[1151]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1151]) );
  DFF \round_reg_reg[1152]  ( .D(out[1152]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1152]) );
  DFF \round_reg_reg[1153]  ( .D(out[1153]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1153]) );
  DFF \round_reg_reg[1154]  ( .D(out[1154]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1154]) );
  DFF \round_reg_reg[1155]  ( .D(out[1155]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1155]) );
  DFF \round_reg_reg[1156]  ( .D(out[1156]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1156]) );
  DFF \round_reg_reg[1157]  ( .D(out[1157]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1157]) );
  DFF \round_reg_reg[1158]  ( .D(out[1158]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1158]) );
  DFF \round_reg_reg[1159]  ( .D(out[1159]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1159]) );
  DFF \round_reg_reg[1160]  ( .D(out[1160]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1160]) );
  DFF \round_reg_reg[1161]  ( .D(out[1161]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1161]) );
  DFF \round_reg_reg[1162]  ( .D(out[1162]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1162]) );
  DFF \round_reg_reg[1163]  ( .D(out[1163]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1163]) );
  DFF \round_reg_reg[1164]  ( .D(out[1164]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1164]) );
  DFF \round_reg_reg[1165]  ( .D(out[1165]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1165]) );
  DFF \round_reg_reg[1166]  ( .D(out[1166]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1166]) );
  DFF \round_reg_reg[1167]  ( .D(out[1167]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1167]) );
  DFF \round_reg_reg[1168]  ( .D(out[1168]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1168]) );
  DFF \round_reg_reg[1169]  ( .D(out[1169]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1169]) );
  DFF \round_reg_reg[1170]  ( .D(out[1170]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1170]) );
  DFF \round_reg_reg[1171]  ( .D(out[1171]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1171]) );
  DFF \round_reg_reg[1172]  ( .D(out[1172]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1172]) );
  DFF \round_reg_reg[1173]  ( .D(out[1173]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1173]) );
  DFF \round_reg_reg[1174]  ( .D(out[1174]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1174]) );
  DFF \round_reg_reg[1175]  ( .D(out[1175]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1175]) );
  DFF \round_reg_reg[1176]  ( .D(out[1176]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1176]) );
  DFF \round_reg_reg[1177]  ( .D(out[1177]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1177]) );
  DFF \round_reg_reg[1178]  ( .D(out[1178]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1178]) );
  DFF \round_reg_reg[1179]  ( .D(out[1179]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1179]) );
  DFF \round_reg_reg[1180]  ( .D(out[1180]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1180]) );
  DFF \round_reg_reg[1181]  ( .D(out[1181]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1181]) );
  DFF \round_reg_reg[1182]  ( .D(out[1182]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1182]) );
  DFF \round_reg_reg[1183]  ( .D(out[1183]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1183]) );
  DFF \round_reg_reg[1184]  ( .D(out[1184]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1184]) );
  DFF \round_reg_reg[1185]  ( .D(out[1185]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1185]) );
  DFF \round_reg_reg[1186]  ( .D(out[1186]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1186]) );
  DFF \round_reg_reg[1187]  ( .D(out[1187]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1187]) );
  DFF \round_reg_reg[1188]  ( .D(out[1188]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1188]) );
  DFF \round_reg_reg[1189]  ( .D(out[1189]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1189]) );
  DFF \round_reg_reg[1190]  ( .D(out[1190]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1190]) );
  DFF \round_reg_reg[1191]  ( .D(out[1191]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1191]) );
  DFF \round_reg_reg[1192]  ( .D(out[1192]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1192]) );
  DFF \round_reg_reg[1193]  ( .D(out[1193]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1193]) );
  DFF \round_reg_reg[1194]  ( .D(out[1194]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1194]) );
  DFF \round_reg_reg[1195]  ( .D(out[1195]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1195]) );
  DFF \round_reg_reg[1196]  ( .D(out[1196]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1196]) );
  DFF \round_reg_reg[1197]  ( .D(out[1197]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1197]) );
  DFF \round_reg_reg[1198]  ( .D(out[1198]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1198]) );
  DFF \round_reg_reg[1199]  ( .D(out[1199]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1199]) );
  DFF \round_reg_reg[1200]  ( .D(out[1200]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1200]) );
  DFF \round_reg_reg[1201]  ( .D(out[1201]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1201]) );
  DFF \round_reg_reg[1202]  ( .D(out[1202]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1202]) );
  DFF \round_reg_reg[1203]  ( .D(out[1203]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1203]) );
  DFF \round_reg_reg[1204]  ( .D(out[1204]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1204]) );
  DFF \round_reg_reg[1205]  ( .D(out[1205]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1205]) );
  DFF \round_reg_reg[1206]  ( .D(out[1206]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1206]) );
  DFF \round_reg_reg[1207]  ( .D(out[1207]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1207]) );
  DFF \round_reg_reg[1208]  ( .D(out[1208]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1208]) );
  DFF \round_reg_reg[1209]  ( .D(out[1209]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1209]) );
  DFF \round_reg_reg[1210]  ( .D(out[1210]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1210]) );
  DFF \round_reg_reg[1211]  ( .D(out[1211]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1211]) );
  DFF \round_reg_reg[1212]  ( .D(out[1212]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1212]) );
  DFF \round_reg_reg[1213]  ( .D(out[1213]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1213]) );
  DFF \round_reg_reg[1214]  ( .D(out[1214]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1214]) );
  DFF \round_reg_reg[1215]  ( .D(out[1215]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1215]) );
  DFF \round_reg_reg[1216]  ( .D(out[1216]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1216]) );
  DFF \round_reg_reg[1217]  ( .D(out[1217]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1217]) );
  DFF \round_reg_reg[1218]  ( .D(out[1218]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1218]) );
  DFF \round_reg_reg[1219]  ( .D(out[1219]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1219]) );
  DFF \round_reg_reg[1220]  ( .D(out[1220]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1220]) );
  DFF \round_reg_reg[1221]  ( .D(out[1221]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1221]) );
  DFF \round_reg_reg[1222]  ( .D(out[1222]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1222]) );
  DFF \round_reg_reg[1223]  ( .D(out[1223]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1223]) );
  DFF \round_reg_reg[1224]  ( .D(out[1224]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1224]) );
  DFF \round_reg_reg[1225]  ( .D(out[1225]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1225]) );
  DFF \round_reg_reg[1226]  ( .D(out[1226]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1226]) );
  DFF \round_reg_reg[1227]  ( .D(out[1227]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1227]) );
  DFF \round_reg_reg[1228]  ( .D(out[1228]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1228]) );
  DFF \round_reg_reg[1229]  ( .D(out[1229]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1229]) );
  DFF \round_reg_reg[1230]  ( .D(out[1230]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1230]) );
  DFF \round_reg_reg[1231]  ( .D(out[1231]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1231]) );
  DFF \round_reg_reg[1232]  ( .D(out[1232]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1232]) );
  DFF \round_reg_reg[1233]  ( .D(out[1233]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1233]) );
  DFF \round_reg_reg[1234]  ( .D(out[1234]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1234]) );
  DFF \round_reg_reg[1235]  ( .D(out[1235]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1235]) );
  DFF \round_reg_reg[1236]  ( .D(out[1236]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1236]) );
  DFF \round_reg_reg[1237]  ( .D(out[1237]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1237]) );
  DFF \round_reg_reg[1238]  ( .D(out[1238]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1238]) );
  DFF \round_reg_reg[1239]  ( .D(out[1239]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1239]) );
  DFF \round_reg_reg[1240]  ( .D(out[1240]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1240]) );
  DFF \round_reg_reg[1241]  ( .D(out[1241]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1241]) );
  DFF \round_reg_reg[1242]  ( .D(out[1242]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1242]) );
  DFF \round_reg_reg[1243]  ( .D(out[1243]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1243]) );
  DFF \round_reg_reg[1244]  ( .D(out[1244]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1244]) );
  DFF \round_reg_reg[1245]  ( .D(out[1245]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1245]) );
  DFF \round_reg_reg[1246]  ( .D(out[1246]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1246]) );
  DFF \round_reg_reg[1247]  ( .D(out[1247]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1247]) );
  DFF \round_reg_reg[1248]  ( .D(out[1248]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1248]) );
  DFF \round_reg_reg[1249]  ( .D(out[1249]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1249]) );
  DFF \round_reg_reg[1250]  ( .D(out[1250]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1250]) );
  DFF \round_reg_reg[1251]  ( .D(out[1251]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1251]) );
  DFF \round_reg_reg[1252]  ( .D(out[1252]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1252]) );
  DFF \round_reg_reg[1253]  ( .D(out[1253]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1253]) );
  DFF \round_reg_reg[1254]  ( .D(out[1254]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1254]) );
  DFF \round_reg_reg[1255]  ( .D(out[1255]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1255]) );
  DFF \round_reg_reg[1256]  ( .D(out[1256]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1256]) );
  DFF \round_reg_reg[1257]  ( .D(out[1257]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1257]) );
  DFF \round_reg_reg[1258]  ( .D(out[1258]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1258]) );
  DFF \round_reg_reg[1259]  ( .D(out[1259]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1259]) );
  DFF \round_reg_reg[1260]  ( .D(out[1260]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1260]) );
  DFF \round_reg_reg[1261]  ( .D(out[1261]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1261]) );
  DFF \round_reg_reg[1262]  ( .D(out[1262]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1262]) );
  DFF \round_reg_reg[1263]  ( .D(out[1263]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1263]) );
  DFF \round_reg_reg[1264]  ( .D(out[1264]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1264]) );
  DFF \round_reg_reg[1265]  ( .D(out[1265]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1265]) );
  DFF \round_reg_reg[1266]  ( .D(out[1266]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1266]) );
  DFF \round_reg_reg[1267]  ( .D(out[1267]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1267]) );
  DFF \round_reg_reg[1268]  ( .D(out[1268]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1268]) );
  DFF \round_reg_reg[1269]  ( .D(out[1269]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1269]) );
  DFF \round_reg_reg[1270]  ( .D(out[1270]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1270]) );
  DFF \round_reg_reg[1271]  ( .D(out[1271]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1271]) );
  DFF \round_reg_reg[1272]  ( .D(out[1272]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1272]) );
  DFF \round_reg_reg[1273]  ( .D(out[1273]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1273]) );
  DFF \round_reg_reg[1274]  ( .D(out[1274]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1274]) );
  DFF \round_reg_reg[1275]  ( .D(out[1275]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1275]) );
  DFF \round_reg_reg[1276]  ( .D(out[1276]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1276]) );
  DFF \round_reg_reg[1277]  ( .D(out[1277]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1277]) );
  DFF \round_reg_reg[1278]  ( .D(out[1278]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1278]) );
  DFF \round_reg_reg[1279]  ( .D(out[1279]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1279]) );
  DFF \round_reg_reg[1280]  ( .D(out[1280]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1280]) );
  DFF \round_reg_reg[1281]  ( .D(out[1281]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1281]) );
  DFF \round_reg_reg[1282]  ( .D(out[1282]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1282]) );
  DFF \round_reg_reg[1283]  ( .D(out[1283]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1283]) );
  DFF \round_reg_reg[1284]  ( .D(out[1284]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1284]) );
  DFF \round_reg_reg[1285]  ( .D(out[1285]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1285]) );
  DFF \round_reg_reg[1286]  ( .D(out[1286]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1286]) );
  DFF \round_reg_reg[1287]  ( .D(out[1287]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1287]) );
  DFF \round_reg_reg[1288]  ( .D(out[1288]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1288]) );
  DFF \round_reg_reg[1289]  ( .D(out[1289]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1289]) );
  DFF \round_reg_reg[1290]  ( .D(out[1290]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1290]) );
  DFF \round_reg_reg[1291]  ( .D(out[1291]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1291]) );
  DFF \round_reg_reg[1292]  ( .D(out[1292]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1292]) );
  DFF \round_reg_reg[1293]  ( .D(out[1293]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1293]) );
  DFF \round_reg_reg[1294]  ( .D(out[1294]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1294]) );
  DFF \round_reg_reg[1295]  ( .D(out[1295]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1295]) );
  DFF \round_reg_reg[1296]  ( .D(out[1296]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1296]) );
  DFF \round_reg_reg[1297]  ( .D(out[1297]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1297]) );
  DFF \round_reg_reg[1298]  ( .D(out[1298]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1298]) );
  DFF \round_reg_reg[1299]  ( .D(out[1299]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1299]) );
  DFF \round_reg_reg[1300]  ( .D(out[1300]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1300]) );
  DFF \round_reg_reg[1301]  ( .D(out[1301]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1301]) );
  DFF \round_reg_reg[1302]  ( .D(out[1302]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1302]) );
  DFF \round_reg_reg[1303]  ( .D(out[1303]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1303]) );
  DFF \round_reg_reg[1304]  ( .D(out[1304]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1304]) );
  DFF \round_reg_reg[1305]  ( .D(out[1305]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1305]) );
  DFF \round_reg_reg[1306]  ( .D(out[1306]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1306]) );
  DFF \round_reg_reg[1307]  ( .D(out[1307]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1307]) );
  DFF \round_reg_reg[1308]  ( .D(out[1308]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1308]) );
  DFF \round_reg_reg[1309]  ( .D(out[1309]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1309]) );
  DFF \round_reg_reg[1310]  ( .D(out[1310]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1310]) );
  DFF \round_reg_reg[1311]  ( .D(out[1311]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1311]) );
  DFF \round_reg_reg[1312]  ( .D(out[1312]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1312]) );
  DFF \round_reg_reg[1313]  ( .D(out[1313]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1313]) );
  DFF \round_reg_reg[1314]  ( .D(out[1314]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1314]) );
  DFF \round_reg_reg[1315]  ( .D(out[1315]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1315]) );
  DFF \round_reg_reg[1316]  ( .D(out[1316]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1316]) );
  DFF \round_reg_reg[1317]  ( .D(out[1317]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1317]) );
  DFF \round_reg_reg[1318]  ( .D(out[1318]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1318]) );
  DFF \round_reg_reg[1319]  ( .D(out[1319]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1319]) );
  DFF \round_reg_reg[1320]  ( .D(out[1320]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1320]) );
  DFF \round_reg_reg[1321]  ( .D(out[1321]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1321]) );
  DFF \round_reg_reg[1322]  ( .D(out[1322]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1322]) );
  DFF \round_reg_reg[1323]  ( .D(out[1323]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1323]) );
  DFF \round_reg_reg[1324]  ( .D(out[1324]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1324]) );
  DFF \round_reg_reg[1325]  ( .D(out[1325]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1325]) );
  DFF \round_reg_reg[1326]  ( .D(out[1326]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1326]) );
  DFF \round_reg_reg[1327]  ( .D(out[1327]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1327]) );
  DFF \round_reg_reg[1328]  ( .D(out[1328]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1328]) );
  DFF \round_reg_reg[1329]  ( .D(out[1329]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1329]) );
  DFF \round_reg_reg[1330]  ( .D(out[1330]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1330]) );
  DFF \round_reg_reg[1331]  ( .D(out[1331]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1331]) );
  DFF \round_reg_reg[1332]  ( .D(out[1332]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1332]) );
  DFF \round_reg_reg[1333]  ( .D(out[1333]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1333]) );
  DFF \round_reg_reg[1334]  ( .D(out[1334]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1334]) );
  DFF \round_reg_reg[1335]  ( .D(out[1335]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1335]) );
  DFF \round_reg_reg[1336]  ( .D(out[1336]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1336]) );
  DFF \round_reg_reg[1337]  ( .D(out[1337]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1337]) );
  DFF \round_reg_reg[1338]  ( .D(out[1338]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1338]) );
  DFF \round_reg_reg[1339]  ( .D(out[1339]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1339]) );
  DFF \round_reg_reg[1340]  ( .D(out[1340]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1340]) );
  DFF \round_reg_reg[1341]  ( .D(out[1341]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1341]) );
  DFF \round_reg_reg[1342]  ( .D(out[1342]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1342]) );
  DFF \round_reg_reg[1343]  ( .D(out[1343]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1343]) );
  DFF \round_reg_reg[1344]  ( .D(out[1344]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1344]) );
  DFF \round_reg_reg[1345]  ( .D(out[1345]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1345]) );
  DFF \round_reg_reg[1346]  ( .D(out[1346]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1346]) );
  DFF \round_reg_reg[1347]  ( .D(out[1347]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1347]) );
  DFF \round_reg_reg[1348]  ( .D(out[1348]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1348]) );
  DFF \round_reg_reg[1349]  ( .D(out[1349]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1349]) );
  DFF \round_reg_reg[1350]  ( .D(out[1350]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1350]) );
  DFF \round_reg_reg[1351]  ( .D(out[1351]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1351]) );
  DFF \round_reg_reg[1352]  ( .D(out[1352]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1352]) );
  DFF \round_reg_reg[1353]  ( .D(out[1353]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1353]) );
  DFF \round_reg_reg[1354]  ( .D(out[1354]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1354]) );
  DFF \round_reg_reg[1355]  ( .D(out[1355]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1355]) );
  DFF \round_reg_reg[1356]  ( .D(out[1356]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1356]) );
  DFF \round_reg_reg[1357]  ( .D(out[1357]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1357]) );
  DFF \round_reg_reg[1358]  ( .D(out[1358]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1358]) );
  DFF \round_reg_reg[1359]  ( .D(out[1359]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1359]) );
  DFF \round_reg_reg[1360]  ( .D(out[1360]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1360]) );
  DFF \round_reg_reg[1361]  ( .D(out[1361]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1361]) );
  DFF \round_reg_reg[1362]  ( .D(out[1362]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1362]) );
  DFF \round_reg_reg[1363]  ( .D(out[1363]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1363]) );
  DFF \round_reg_reg[1364]  ( .D(out[1364]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1364]) );
  DFF \round_reg_reg[1365]  ( .D(out[1365]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1365]) );
  DFF \round_reg_reg[1366]  ( .D(out[1366]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1366]) );
  DFF \round_reg_reg[1367]  ( .D(out[1367]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1367]) );
  DFF \round_reg_reg[1368]  ( .D(out[1368]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1368]) );
  DFF \round_reg_reg[1369]  ( .D(out[1369]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1369]) );
  DFF \round_reg_reg[1370]  ( .D(out[1370]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1370]) );
  DFF \round_reg_reg[1371]  ( .D(out[1371]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1371]) );
  DFF \round_reg_reg[1372]  ( .D(out[1372]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1372]) );
  DFF \round_reg_reg[1373]  ( .D(out[1373]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1373]) );
  DFF \round_reg_reg[1374]  ( .D(out[1374]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1374]) );
  DFF \round_reg_reg[1375]  ( .D(out[1375]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1375]) );
  DFF \round_reg_reg[1376]  ( .D(out[1376]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1376]) );
  DFF \round_reg_reg[1377]  ( .D(out[1377]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1377]) );
  DFF \round_reg_reg[1378]  ( .D(out[1378]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1378]) );
  DFF \round_reg_reg[1379]  ( .D(out[1379]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1379]) );
  DFF \round_reg_reg[1380]  ( .D(out[1380]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1380]) );
  DFF \round_reg_reg[1381]  ( .D(out[1381]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1381]) );
  DFF \round_reg_reg[1382]  ( .D(out[1382]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1382]) );
  DFF \round_reg_reg[1383]  ( .D(out[1383]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1383]) );
  DFF \round_reg_reg[1384]  ( .D(out[1384]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1384]) );
  DFF \round_reg_reg[1385]  ( .D(out[1385]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1385]) );
  DFF \round_reg_reg[1386]  ( .D(out[1386]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1386]) );
  DFF \round_reg_reg[1387]  ( .D(out[1387]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1387]) );
  DFF \round_reg_reg[1388]  ( .D(out[1388]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1388]) );
  DFF \round_reg_reg[1389]  ( .D(out[1389]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1389]) );
  DFF \round_reg_reg[1390]  ( .D(out[1390]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1390]) );
  DFF \round_reg_reg[1391]  ( .D(out[1391]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1391]) );
  DFF \round_reg_reg[1392]  ( .D(out[1392]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1392]) );
  DFF \round_reg_reg[1393]  ( .D(out[1393]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1393]) );
  DFF \round_reg_reg[1394]  ( .D(out[1394]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1394]) );
  DFF \round_reg_reg[1395]  ( .D(out[1395]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1395]) );
  DFF \round_reg_reg[1396]  ( .D(out[1396]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1396]) );
  DFF \round_reg_reg[1397]  ( .D(out[1397]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1397]) );
  DFF \round_reg_reg[1398]  ( .D(out[1398]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1398]) );
  DFF \round_reg_reg[1399]  ( .D(out[1399]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1399]) );
  DFF \round_reg_reg[1400]  ( .D(out[1400]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1400]) );
  DFF \round_reg_reg[1401]  ( .D(out[1401]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1401]) );
  DFF \round_reg_reg[1402]  ( .D(out[1402]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1402]) );
  DFF \round_reg_reg[1403]  ( .D(out[1403]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1403]) );
  DFF \round_reg_reg[1404]  ( .D(out[1404]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1404]) );
  DFF \round_reg_reg[1405]  ( .D(out[1405]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1405]) );
  DFF \round_reg_reg[1406]  ( .D(out[1406]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1406]) );
  DFF \round_reg_reg[1407]  ( .D(out[1407]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1407]) );
  DFF \round_reg_reg[1408]  ( .D(out[1408]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1408]) );
  DFF \round_reg_reg[1409]  ( .D(out[1409]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1409]) );
  DFF \round_reg_reg[1410]  ( .D(out[1410]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1410]) );
  DFF \round_reg_reg[1411]  ( .D(out[1411]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1411]) );
  DFF \round_reg_reg[1412]  ( .D(out[1412]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1412]) );
  DFF \round_reg_reg[1413]  ( .D(out[1413]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1413]) );
  DFF \round_reg_reg[1414]  ( .D(out[1414]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1414]) );
  DFF \round_reg_reg[1415]  ( .D(out[1415]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1415]) );
  DFF \round_reg_reg[1416]  ( .D(out[1416]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1416]) );
  DFF \round_reg_reg[1417]  ( .D(out[1417]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1417]) );
  DFF \round_reg_reg[1418]  ( .D(out[1418]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1418]) );
  DFF \round_reg_reg[1419]  ( .D(out[1419]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1419]) );
  DFF \round_reg_reg[1420]  ( .D(out[1420]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1420]) );
  DFF \round_reg_reg[1421]  ( .D(out[1421]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1421]) );
  DFF \round_reg_reg[1422]  ( .D(out[1422]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1422]) );
  DFF \round_reg_reg[1423]  ( .D(out[1423]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1423]) );
  DFF \round_reg_reg[1424]  ( .D(out[1424]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1424]) );
  DFF \round_reg_reg[1425]  ( .D(out[1425]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1425]) );
  DFF \round_reg_reg[1426]  ( .D(out[1426]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1426]) );
  DFF \round_reg_reg[1427]  ( .D(out[1427]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1427]) );
  DFF \round_reg_reg[1428]  ( .D(out[1428]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1428]) );
  DFF \round_reg_reg[1429]  ( .D(out[1429]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1429]) );
  DFF \round_reg_reg[1430]  ( .D(out[1430]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1430]) );
  DFF \round_reg_reg[1431]  ( .D(out[1431]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1431]) );
  DFF \round_reg_reg[1432]  ( .D(out[1432]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1432]) );
  DFF \round_reg_reg[1433]  ( .D(out[1433]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1433]) );
  DFF \round_reg_reg[1434]  ( .D(out[1434]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1434]) );
  DFF \round_reg_reg[1435]  ( .D(out[1435]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1435]) );
  DFF \round_reg_reg[1436]  ( .D(out[1436]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1436]) );
  DFF \round_reg_reg[1437]  ( .D(out[1437]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1437]) );
  DFF \round_reg_reg[1438]  ( .D(out[1438]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1438]) );
  DFF \round_reg_reg[1439]  ( .D(out[1439]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1439]) );
  DFF \round_reg_reg[1440]  ( .D(out[1440]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1440]) );
  DFF \round_reg_reg[1441]  ( .D(out[1441]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1441]) );
  DFF \round_reg_reg[1442]  ( .D(out[1442]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1442]) );
  DFF \round_reg_reg[1443]  ( .D(out[1443]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1443]) );
  DFF \round_reg_reg[1444]  ( .D(out[1444]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1444]) );
  DFF \round_reg_reg[1445]  ( .D(out[1445]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1445]) );
  DFF \round_reg_reg[1446]  ( .D(out[1446]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1446]) );
  DFF \round_reg_reg[1447]  ( .D(out[1447]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1447]) );
  DFF \round_reg_reg[1448]  ( .D(out[1448]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1448]) );
  DFF \round_reg_reg[1449]  ( .D(out[1449]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1449]) );
  DFF \round_reg_reg[1450]  ( .D(out[1450]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1450]) );
  DFF \round_reg_reg[1451]  ( .D(out[1451]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1451]) );
  DFF \round_reg_reg[1452]  ( .D(out[1452]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1452]) );
  DFF \round_reg_reg[1453]  ( .D(out[1453]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1453]) );
  DFF \round_reg_reg[1454]  ( .D(out[1454]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1454]) );
  DFF \round_reg_reg[1455]  ( .D(out[1455]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1455]) );
  DFF \round_reg_reg[1456]  ( .D(out[1456]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1456]) );
  DFF \round_reg_reg[1457]  ( .D(out[1457]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1457]) );
  DFF \round_reg_reg[1458]  ( .D(out[1458]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1458]) );
  DFF \round_reg_reg[1459]  ( .D(out[1459]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1459]) );
  DFF \round_reg_reg[1460]  ( .D(out[1460]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1460]) );
  DFF \round_reg_reg[1461]  ( .D(out[1461]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1461]) );
  DFF \round_reg_reg[1462]  ( .D(out[1462]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1462]) );
  DFF \round_reg_reg[1463]  ( .D(out[1463]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1463]) );
  DFF \round_reg_reg[1464]  ( .D(out[1464]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1464]) );
  DFF \round_reg_reg[1465]  ( .D(out[1465]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1465]) );
  DFF \round_reg_reg[1466]  ( .D(out[1466]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1466]) );
  DFF \round_reg_reg[1467]  ( .D(out[1467]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1467]) );
  DFF \round_reg_reg[1468]  ( .D(out[1468]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1468]) );
  DFF \round_reg_reg[1469]  ( .D(out[1469]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1469]) );
  DFF \round_reg_reg[1470]  ( .D(out[1470]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1470]) );
  DFF \round_reg_reg[1471]  ( .D(out[1471]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1471]) );
  DFF \round_reg_reg[1472]  ( .D(out[1472]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1472]) );
  DFF \round_reg_reg[1473]  ( .D(out[1473]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1473]) );
  DFF \round_reg_reg[1474]  ( .D(out[1474]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1474]) );
  DFF \round_reg_reg[1475]  ( .D(out[1475]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1475]) );
  DFF \round_reg_reg[1476]  ( .D(out[1476]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1476]) );
  DFF \round_reg_reg[1477]  ( .D(out[1477]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1477]) );
  DFF \round_reg_reg[1478]  ( .D(out[1478]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1478]) );
  DFF \round_reg_reg[1479]  ( .D(out[1479]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1479]) );
  DFF \round_reg_reg[1480]  ( .D(out[1480]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1480]) );
  DFF \round_reg_reg[1481]  ( .D(out[1481]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1481]) );
  DFF \round_reg_reg[1482]  ( .D(out[1482]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1482]) );
  DFF \round_reg_reg[1483]  ( .D(out[1483]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1483]) );
  DFF \round_reg_reg[1484]  ( .D(out[1484]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1484]) );
  DFF \round_reg_reg[1485]  ( .D(out[1485]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1485]) );
  DFF \round_reg_reg[1486]  ( .D(out[1486]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1486]) );
  DFF \round_reg_reg[1487]  ( .D(out[1487]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1487]) );
  DFF \round_reg_reg[1488]  ( .D(out[1488]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1488]) );
  DFF \round_reg_reg[1489]  ( .D(out[1489]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1489]) );
  DFF \round_reg_reg[1490]  ( .D(out[1490]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1490]) );
  DFF \round_reg_reg[1491]  ( .D(out[1491]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1491]) );
  DFF \round_reg_reg[1492]  ( .D(out[1492]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1492]) );
  DFF \round_reg_reg[1493]  ( .D(out[1493]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1493]) );
  DFF \round_reg_reg[1494]  ( .D(out[1494]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1494]) );
  DFF \round_reg_reg[1495]  ( .D(out[1495]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1495]) );
  DFF \round_reg_reg[1496]  ( .D(out[1496]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1496]) );
  DFF \round_reg_reg[1497]  ( .D(out[1497]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1497]) );
  DFF \round_reg_reg[1498]  ( .D(out[1498]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1498]) );
  DFF \round_reg_reg[1499]  ( .D(out[1499]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1499]) );
  DFF \round_reg_reg[1500]  ( .D(out[1500]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1500]) );
  DFF \round_reg_reg[1501]  ( .D(out[1501]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1501]) );
  DFF \round_reg_reg[1502]  ( .D(out[1502]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1502]) );
  DFF \round_reg_reg[1503]  ( .D(out[1503]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1503]) );
  DFF \round_reg_reg[1504]  ( .D(out[1504]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1504]) );
  DFF \round_reg_reg[1505]  ( .D(out[1505]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1505]) );
  DFF \round_reg_reg[1506]  ( .D(out[1506]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1506]) );
  DFF \round_reg_reg[1507]  ( .D(out[1507]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1507]) );
  DFF \round_reg_reg[1508]  ( .D(out[1508]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1508]) );
  DFF \round_reg_reg[1509]  ( .D(out[1509]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1509]) );
  DFF \round_reg_reg[1510]  ( .D(out[1510]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1510]) );
  DFF \round_reg_reg[1511]  ( .D(out[1511]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1511]) );
  DFF \round_reg_reg[1512]  ( .D(out[1512]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1512]) );
  DFF \round_reg_reg[1513]  ( .D(out[1513]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1513]) );
  DFF \round_reg_reg[1514]  ( .D(out[1514]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1514]) );
  DFF \round_reg_reg[1515]  ( .D(out[1515]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1515]) );
  DFF \round_reg_reg[1516]  ( .D(out[1516]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1516]) );
  DFF \round_reg_reg[1517]  ( .D(out[1517]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1517]) );
  DFF \round_reg_reg[1518]  ( .D(out[1518]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1518]) );
  DFF \round_reg_reg[1519]  ( .D(out[1519]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1519]) );
  DFF \round_reg_reg[1520]  ( .D(out[1520]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1520]) );
  DFF \round_reg_reg[1521]  ( .D(out[1521]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1521]) );
  DFF \round_reg_reg[1522]  ( .D(out[1522]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1522]) );
  DFF \round_reg_reg[1523]  ( .D(out[1523]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1523]) );
  DFF \round_reg_reg[1524]  ( .D(out[1524]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1524]) );
  DFF \round_reg_reg[1525]  ( .D(out[1525]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1525]) );
  DFF \round_reg_reg[1526]  ( .D(out[1526]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1526]) );
  DFF \round_reg_reg[1527]  ( .D(out[1527]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1527]) );
  DFF \round_reg_reg[1528]  ( .D(out[1528]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1528]) );
  DFF \round_reg_reg[1529]  ( .D(out[1529]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1529]) );
  DFF \round_reg_reg[1530]  ( .D(out[1530]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1530]) );
  DFF \round_reg_reg[1531]  ( .D(out[1531]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1531]) );
  DFF \round_reg_reg[1532]  ( .D(out[1532]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1532]) );
  DFF \round_reg_reg[1533]  ( .D(out[1533]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1533]) );
  DFF \round_reg_reg[1534]  ( .D(out[1534]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1534]) );
  DFF \round_reg_reg[1535]  ( .D(out[1535]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1535]) );
  DFF \round_reg_reg[1536]  ( .D(out[1536]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1536]) );
  DFF \round_reg_reg[1537]  ( .D(out[1537]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1537]) );
  DFF \round_reg_reg[1538]  ( .D(out[1538]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1538]) );
  DFF \round_reg_reg[1539]  ( .D(out[1539]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1539]) );
  DFF \round_reg_reg[1540]  ( .D(out[1540]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1540]) );
  DFF \round_reg_reg[1541]  ( .D(out[1541]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1541]) );
  DFF \round_reg_reg[1542]  ( .D(out[1542]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1542]) );
  DFF \round_reg_reg[1543]  ( .D(out[1543]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1543]) );
  DFF \round_reg_reg[1544]  ( .D(out[1544]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1544]) );
  DFF \round_reg_reg[1545]  ( .D(out[1545]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1545]) );
  DFF \round_reg_reg[1546]  ( .D(out[1546]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1546]) );
  DFF \round_reg_reg[1547]  ( .D(out[1547]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1547]) );
  DFF \round_reg_reg[1548]  ( .D(out[1548]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1548]) );
  DFF \round_reg_reg[1549]  ( .D(out[1549]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1549]) );
  DFF \round_reg_reg[1550]  ( .D(out[1550]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1550]) );
  DFF \round_reg_reg[1551]  ( .D(out[1551]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1551]) );
  DFF \round_reg_reg[1552]  ( .D(out[1552]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1552]) );
  DFF \round_reg_reg[1553]  ( .D(out[1553]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1553]) );
  DFF \round_reg_reg[1554]  ( .D(out[1554]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1554]) );
  DFF \round_reg_reg[1555]  ( .D(out[1555]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1555]) );
  DFF \round_reg_reg[1556]  ( .D(out[1556]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1556]) );
  DFF \round_reg_reg[1557]  ( .D(out[1557]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1557]) );
  DFF \round_reg_reg[1558]  ( .D(out[1558]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1558]) );
  DFF \round_reg_reg[1559]  ( .D(out[1559]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1559]) );
  DFF \round_reg_reg[1560]  ( .D(out[1560]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1560]) );
  DFF \round_reg_reg[1561]  ( .D(out[1561]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1561]) );
  DFF \round_reg_reg[1562]  ( .D(out[1562]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1562]) );
  DFF \round_reg_reg[1563]  ( .D(out[1563]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1563]) );
  DFF \round_reg_reg[1564]  ( .D(out[1564]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1564]) );
  DFF \round_reg_reg[1565]  ( .D(out[1565]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1565]) );
  DFF \round_reg_reg[1566]  ( .D(out[1566]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1566]) );
  DFF \round_reg_reg[1567]  ( .D(out[1567]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1567]) );
  DFF \round_reg_reg[1568]  ( .D(out[1568]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1568]) );
  DFF \round_reg_reg[1569]  ( .D(out[1569]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1569]) );
  DFF \round_reg_reg[1570]  ( .D(out[1570]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1570]) );
  DFF \round_reg_reg[1571]  ( .D(out[1571]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1571]) );
  DFF \round_reg_reg[1572]  ( .D(out[1572]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1572]) );
  DFF \round_reg_reg[1573]  ( .D(out[1573]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1573]) );
  DFF \round_reg_reg[1574]  ( .D(out[1574]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1574]) );
  DFF \round_reg_reg[1575]  ( .D(out[1575]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1575]) );
  DFF \round_reg_reg[1576]  ( .D(out[1576]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1576]) );
  DFF \round_reg_reg[1577]  ( .D(out[1577]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1577]) );
  DFF \round_reg_reg[1578]  ( .D(out[1578]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1578]) );
  DFF \round_reg_reg[1579]  ( .D(out[1579]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1579]) );
  DFF \round_reg_reg[1580]  ( .D(out[1580]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1580]) );
  DFF \round_reg_reg[1581]  ( .D(out[1581]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1581]) );
  DFF \round_reg_reg[1582]  ( .D(out[1582]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1582]) );
  DFF \round_reg_reg[1583]  ( .D(out[1583]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1583]) );
  DFF \round_reg_reg[1584]  ( .D(out[1584]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1584]) );
  DFF \round_reg_reg[1585]  ( .D(out[1585]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1585]) );
  DFF \round_reg_reg[1586]  ( .D(out[1586]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1586]) );
  DFF \round_reg_reg[1587]  ( .D(out[1587]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1587]) );
  DFF \round_reg_reg[1588]  ( .D(out[1588]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1588]) );
  DFF \round_reg_reg[1589]  ( .D(out[1589]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1589]) );
  DFF \round_reg_reg[1590]  ( .D(out[1590]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1590]) );
  DFF \round_reg_reg[1591]  ( .D(out[1591]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1591]) );
  DFF \round_reg_reg[1592]  ( .D(out[1592]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1592]) );
  DFF \round_reg_reg[1593]  ( .D(out[1593]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1593]) );
  DFF \round_reg_reg[1594]  ( .D(out[1594]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1594]) );
  DFF \round_reg_reg[1595]  ( .D(out[1595]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1595]) );
  DFF \round_reg_reg[1596]  ( .D(out[1596]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1596]) );
  DFF \round_reg_reg[1597]  ( .D(out[1597]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1597]) );
  DFF \round_reg_reg[1598]  ( .D(out[1598]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1598]) );
  DFF \round_reg_reg[1599]  ( .D(out[1599]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1599]) );
  NOR U1041 ( .A(n7973), .B(n7975), .Z(n10919) );
  XNOR U1042 ( .A(n6386), .B(n6511), .Z(n5165) );
  XNOR U1043 ( .A(n6390), .B(n6537), .Z(n5173) );
  XOR U1044 ( .A(n7534), .B(n6289), .Z(n2387) );
  XOR U1045 ( .A(n8896), .B(n8895), .Z(n2462) );
  XOR U1046 ( .A(n9015), .B(n9014), .Z(n2480) );
  XOR U1047 ( .A(n6350), .B(n9328), .Z(n1737) );
  XOR U1048 ( .A(n6358), .B(n9475), .Z(n1747) );
  ANDN U1049 ( .B(n4595), .A(n4596), .Z(n4593) );
  ANDN U1050 ( .B(n4368), .A(n4850), .Z(n5103) );
  ANDN U1051 ( .B(n4372), .A(n4853), .Z(n5105) );
  ANDN U1052 ( .B(n5679), .A(n5680), .Z(n5677) );
  XNOR U1053 ( .A(n1227), .B(n1228), .Z(out[958]) );
  XNOR U1054 ( .A(n1328), .B(n1329), .Z(out[934]) );
  XNOR U1055 ( .A(n1332), .B(n2077), .Z(out[933]) );
  XNOR U1056 ( .A(n11752), .B(n11751), .Z(n9779) );
  XOR U1057 ( .A(round_reg[709]), .B(n10293), .Z(n7898) );
  NOR U1058 ( .A(n7903), .B(n7905), .Z(n10833) );
  ANDN U1059 ( .B(n7013), .A(n7011), .Z(n7991) );
  XNOR U1060 ( .A(n6378), .B(n6459), .Z(n5159) );
  XNOR U1061 ( .A(n6382), .B(n6485), .Z(n5162) );
  XNOR U1062 ( .A(n9922), .B(n7875), .Z(n1853) );
  NOR U1063 ( .A(n10309), .B(n10374), .Z(n10964) );
  ANDN U1064 ( .B(n7788), .A(n7789), .Z(n7786) );
  XOR U1065 ( .A(n8779), .B(n8778), .Z(n2445) );
  XOR U1066 ( .A(n6338), .B(n9068), .Z(n1724) );
  XOR U1067 ( .A(n6370), .B(n9639), .Z(n1757) );
  ANDN U1068 ( .B(n4532), .A(n4533), .Z(n4530) );
  ANDN U1069 ( .B(n4571), .A(n4572), .Z(n4569) );
  ANDN U1070 ( .B(n4579), .A(n4580), .Z(n4577) );
  ANDN U1071 ( .B(n4591), .A(n4592), .Z(n4589) );
  ANDN U1072 ( .B(n4599), .A(n4600), .Z(n4597) );
  ANDN U1073 ( .B(n4682), .A(n4374), .Z(n4681) );
  ANDN U1074 ( .B(n4684), .A(n4378), .Z(n4683) );
  ANDN U1075 ( .B(n4738), .A(n4482), .Z(n4737) );
  ANDN U1076 ( .B(n4914), .A(n4720), .Z(n4912) );
  ANDN U1077 ( .B(n5683), .A(n5684), .Z(n5681) );
  ANDN U1078 ( .B(n1185), .A(n1186), .Z(n1183) );
  XNOR U1079 ( .A(n1282), .B(n2033), .Z(out[944]) );
  XNOR U1080 ( .A(n1286), .B(n2037), .Z(out[943]) );
  XNOR U1081 ( .A(n1294), .B(n2049), .Z(out[941]) );
  ANDN U1082 ( .B(n1322), .A(n1323), .Z(n1320) );
  ANDN U1083 ( .B(n1365), .A(n1366), .Z(n1363) );
  ANDN U1084 ( .B(n1664), .A(n1506), .Z(n1661) );
  ANDN U1085 ( .B(n1672), .A(n1508), .Z(n1669) );
  ANDN U1086 ( .B(n1729), .A(n1534), .Z(n1726) );
  ANDN U1087 ( .B(n1785), .A(n1560), .Z(n1782) );
  ANDN U1088 ( .B(n1789), .A(n1563), .Z(n1786) );
  ANDN U1089 ( .B(n1793), .A(n1569), .Z(n1790) );
  XNOR U1090 ( .A(n11150), .B(n11149), .Z(n9684) );
  XNOR U1091 ( .A(n10690), .B(n12080), .Z(n10384) );
  XNOR U1092 ( .A(n12528), .B(n11506), .Z(n11107) );
  XNOR U1093 ( .A(n11446), .B(n11445), .Z(n10291) );
  XNOR U1094 ( .A(n11013), .B(n11108), .Z(n9092) );
  XOR U1095 ( .A(n12578), .B(n12577), .Z(n9901) );
  XOR U1096 ( .A(round_reg[1379]), .B(n9928), .Z(n6996) );
  NOR U1097 ( .A(n9506), .B(n9507), .Z(n10276) );
  ANDN U1098 ( .B(n6764), .A(n6763), .Z(n7265) );
  ANDN U1099 ( .B(n7038), .A(n7036), .Z(n9290) );
  NOR U1100 ( .A(n7059), .B(n7061), .Z(n10088) );
  NOR U1101 ( .A(n8353), .B(n8352), .Z(n8350) );
  ANDN U1102 ( .B(n7831), .A(n7830), .Z(n10757) );
  NOR U1103 ( .A(n7897), .B(n7898), .Z(n10839) );
  NOR U1104 ( .A(n7967), .B(n7968), .Z(n10925) );
  ANDN U1105 ( .B(n6498), .A(n11370), .Z(n11447) );
  XNOR U1106 ( .A(n6398), .B(n6597), .Z(n5179) );
  XNOR U1107 ( .A(n12777), .B(n7750), .Z(n7732) );
  ANDN U1108 ( .B(n8478), .A(n8564), .Z(n8563) );
  ANDN U1109 ( .B(n6667), .A(n6668), .Z(n6665) );
  NOR U1110 ( .A(n8213), .B(n8173), .Z(n8212) );
  ANDN U1111 ( .B(n8541), .A(n8683), .Z(n8682) );
  NOR U1112 ( .A(n10731), .B(n8347), .Z(n10729) );
  ANDN U1113 ( .B(n7922), .A(n7920), .Z(n8969) );
  XOR U1114 ( .A(n6035), .B(n6034), .Z(n2191) );
  XOR U1115 ( .A(n6253), .B(n8020), .Z(n1946) );
  XOR U1116 ( .A(n6280), .B(n8252), .Z(n1971) );
  XOR U1117 ( .A(n2127), .B(n5942), .Z(n1061) );
  ANDN U1118 ( .B(n4548), .A(n4549), .Z(n4546) );
  ANDN U1119 ( .B(n4567), .A(n4568), .Z(n4560) );
  ANDN U1120 ( .B(n4583), .A(n4584), .Z(n4581) );
  ANDN U1121 ( .B(n4622), .A(n4623), .Z(n4620) );
  ANDN U1122 ( .B(n5657), .A(n5658), .Z(n5655) );
  ANDN U1123 ( .B(n5730), .A(n1054), .Z(n5729) );
  ANDN U1124 ( .B(n5737), .A(n1066), .Z(n5736) );
  ANDN U1125 ( .B(n5818), .A(n1174), .Z(n5817) );
  ANDN U1126 ( .B(n6259), .A(n5911), .Z(n6255) );
  XNOR U1127 ( .A(n1239), .B(n1989), .Z(out[955]) );
  XNOR U1128 ( .A(n1268), .B(n2018), .Z(out[948]) );
  XNOR U1129 ( .A(n1290), .B(n2041), .Z(out[942]) );
  XNOR U1130 ( .A(n1298), .B(n2053), .Z(out[940]) );
  ANDN U1131 ( .B(n1308), .A(n1309), .Z(n1306) );
  XNOR U1132 ( .A(n1310), .B(n1311), .Z(out[938]) );
  XNOR U1133 ( .A(n1315), .B(n1316), .Z(out[937]) );
  ANDN U1134 ( .B(n1345), .A(n1346), .Z(n1343) );
  ANDN U1135 ( .B(n1361), .A(n1362), .Z(n1359) );
  ANDN U1136 ( .B(n1369), .A(n1370), .Z(n1367) );
  ANDN U1137 ( .B(n1421), .A(n1422), .Z(n1419) );
  NOR U1138 ( .A(n1283), .B(n1739), .Z(n1537) );
  NOR U1139 ( .A(n1287), .B(n1744), .Z(n1543) );
  NOR U1140 ( .A(n1295), .B(n1754), .Z(n1547) );
  ANDN U1141 ( .B(n1631), .A(n1454), .Z(n1630) );
  ANDN U1142 ( .B(n1633), .A(n1458), .Z(n1632) );
  ANDN U1143 ( .B(n1635), .A(n1462), .Z(n1634) );
  NOR U1144 ( .A(n1793), .B(n2077), .Z(n2074) );
  NOR U1145 ( .A(n1829), .B(n1364), .Z(n2103) );
  ANDN U1146 ( .B(n3281), .A(n3075), .Z(n3279) );
  ANDN U1147 ( .B(n3285), .A(n3077), .Z(n3282) );
  ANDN U1148 ( .B(n3288), .A(n3083), .Z(n3286) );
  NOR U1149 ( .A(n3371), .B(n2939), .Z(n3553) );
  NOR U1150 ( .A(n3374), .B(n2943), .Z(n3556) );
  NOR U1151 ( .A(n3377), .B(n2947), .Z(n3563) );
  XNOR U1152 ( .A(n11717), .B(n12652), .Z(n11240) );
  XNOR U1153 ( .A(n11709), .B(n11416), .Z(n9824) );
  XNOR U1154 ( .A(n11585), .B(n11584), .Z(n9677) );
  XNOR U1155 ( .A(n12116), .B(n11854), .Z(n10042) );
  XOR U1156 ( .A(n11380), .B(n11379), .Z(n9749) );
  XNOR U1157 ( .A(n12633), .B(n12108), .Z(n9386) );
  XNOR U1158 ( .A(n12351), .B(n12350), .Z(n10923) );
  XNOR U1159 ( .A(n11004), .B(n11003), .Z(n9758) );
  XNOR U1160 ( .A(n11395), .B(n11394), .Z(n10601) );
  XNOR U1161 ( .A(n11496), .B(n11055), .Z(n9109) );
  XOR U1162 ( .A(n11456), .B(n11014), .Z(n9191) );
  XOR U1163 ( .A(n11032), .B(n11031), .Z(n9621) );
  XOR U1164 ( .A(round_reg[721]), .B(n9829), .Z(n8005) );
  XOR U1165 ( .A(round_reg[1410]), .B(n9859), .Z(n6983) );
  XOR U1166 ( .A(round_reg[234]), .B(n11048), .Z(n9032) );
  XOR U1167 ( .A(round_reg[15]), .B(n10504), .Z(n10234) );
  XOR U1168 ( .A(round_reg[8]), .B(n10492), .Z(n10816) );
  NOR U1169 ( .A(n7607), .B(n7546), .Z(n7606) );
  NOR U1170 ( .A(n6654), .B(n7140), .Z(n9114) );
  NOR U1171 ( .A(n7778), .B(n7779), .Z(n10661) );
  NOR U1172 ( .A(n8249), .B(n8248), .Z(n8246) );
  XNOR U1173 ( .A(n6094), .B(n6093), .Z(n5600) );
  NOR U1174 ( .A(n7243), .B(n8381), .Z(n10706) );
  ANDN U1175 ( .B(n9643), .A(n9644), .Z(n9641) );
  ANDN U1176 ( .B(n9291), .A(n10144), .Z(n12576) );
  ANDN U1177 ( .B(n10089), .A(n10229), .Z(n10316) );
  NOR U1178 ( .A(n9793), .B(n9743), .Z(n9791) );
  XNOR U1179 ( .A(n9629), .B(n7553), .Z(n7535) );
  XNOR U1180 ( .A(n9701), .B(n7605), .Z(n7588) );
  NOR U1181 ( .A(n6889), .B(n6891), .Z(n7543) );
  NOR U1182 ( .A(n7363), .B(n7364), .Z(n8414) );
  NOR U1183 ( .A(n7210), .B(n8327), .Z(n10620) );
  ANDN U1184 ( .B(n8914), .A(n8986), .Z(n8985) );
  ANDN U1185 ( .B(n7827), .A(n7826), .Z(n10756) );
  NOR U1186 ( .A(n7758), .B(n7665), .Z(n7757) );
  NOR U1187 ( .A(n9874), .B(n9875), .Z(n10675) );
  ANDN U1188 ( .B(n7078), .A(n7076), .Z(n10967) );
  ANDN U1189 ( .B(n8025), .A(n8026), .Z(n8023) );
  ANDN U1190 ( .B(n7793), .A(n7791), .Z(n8849) );
  ANDN U1191 ( .B(n6489), .A(n8703), .Z(n8701) );
  NOR U1192 ( .A(n7907), .B(n7908), .Z(n10831) );
  NOR U1193 ( .A(n7977), .B(n7978), .Z(n10917) );
  NOR U1194 ( .A(n7015), .B(n7016), .Z(n7987) );
  NOR U1195 ( .A(n7318), .B(n7319), .Z(n8363) );
  NOR U1196 ( .A(n7442), .B(n7444), .Z(n8470) );
  NOR U1197 ( .A(n9179), .B(n8004), .Z(n9177) );
  XOR U1198 ( .A(n6248), .B(n7912), .Z(n1941) );
  XOR U1199 ( .A(n6263), .B(n8137), .Z(n1957) );
  XOR U1200 ( .A(n6269), .B(n8198), .Z(n1966) );
  XOR U1201 ( .A(n6342), .B(n9144), .Z(n1728) );
  XOR U1202 ( .A(n6354), .B(n9398), .Z(n1742) );
  XOR U1203 ( .A(n6362), .B(n9558), .Z(n1752) );
  ANDN U1204 ( .B(n4345), .A(n4346), .Z(n4335) );
  ANDN U1205 ( .B(n4397), .A(n4398), .Z(n4395) );
  ANDN U1206 ( .B(n4516), .A(n4517), .Z(n4514) );
  ANDN U1207 ( .B(n4528), .A(n4529), .Z(n4526) );
  ANDN U1208 ( .B(n4544), .A(n4545), .Z(n4542) );
  ANDN U1209 ( .B(n4552), .A(n4553), .Z(n4550) );
  ANDN U1210 ( .B(n4556), .A(n4557), .Z(n4554) );
  ANDN U1211 ( .B(n4641), .A(n4642), .Z(n4639) );
  ANDN U1212 ( .B(n4650), .A(n4651), .Z(n4645) );
  ANDN U1213 ( .B(n4667), .A(n4358), .Z(n4666) );
  ANDN U1214 ( .B(n5021), .A(n4788), .Z(n5018) );
  ANDN U1215 ( .B(n5025), .A(n4790), .Z(n5022) );
  NOR U1216 ( .A(n4558), .B(n5013), .Z(n5245) );
  ANDN U1217 ( .B(n5675), .A(n5676), .Z(n5673) );
  ANDN U1218 ( .B(n5739), .A(n1070), .Z(n5738) );
  ANDN U1219 ( .B(n1189), .A(n1190), .Z(n1187) );
  XNOR U1220 ( .A(n1223), .B(n1224), .Z(out[959]) );
  XNOR U1221 ( .A(n1254), .B(n2006), .Z(out[951]) );
  XNOR U1222 ( .A(n1265), .B(n2014), .Z(out[949]) );
  XNOR U1223 ( .A(n1279), .B(n2029), .Z(out[945]) );
  XNOR U1224 ( .A(n1324), .B(n1325), .Z(out[935]) );
  ANDN U1225 ( .B(n1337), .A(n1338), .Z(n1335) );
  ANDN U1226 ( .B(n1341), .A(n1342), .Z(n1339) );
  ANDN U1227 ( .B(n1353), .A(n1354), .Z(n1351) );
  NOR U1228 ( .A(n1291), .B(n1749), .Z(n1545) );
  NOR U1229 ( .A(n1299), .B(n1759), .Z(n1549) );
  NOR U1230 ( .A(n1312), .B(n1768), .Z(n1553) );
  NOR U1231 ( .A(n1317), .B(n1777), .Z(n1555) );
  ANDN U1232 ( .B(n1599), .A(n1390), .Z(n1598) );
  ANDN U1233 ( .B(n1605), .A(n1406), .Z(n1604) );
  ANDN U1234 ( .B(n1607), .A(n1410), .Z(n1606) );
  ANDN U1235 ( .B(n1609), .A(n1414), .Z(n1608) );
  ANDN U1236 ( .B(n1725), .A(n1532), .Z(n1722) );
  ANDN U1237 ( .B(n1579), .A(n1813), .Z(n1810) );
  NOR U1238 ( .A(n1706), .B(n2010), .Z(n2007) );
  NOR U1239 ( .A(n1716), .B(n2018), .Z(n2015) );
  NOR U1240 ( .A(n1729), .B(n2025), .Z(n2022) );
  NOR U1241 ( .A(n1743), .B(n2037), .Z(n2034) );
  NOR U1242 ( .A(n1753), .B(n2049), .Z(n2046) );
  NOR U1243 ( .A(n1833), .B(n1368), .Z(n2106) );
  XNOR U1244 ( .A(n2908), .B(n3533), .Z(out[591]) );
  XNOR U1245 ( .A(n2911), .B(n3536), .Z(out[590]) );
  XNOR U1246 ( .A(n2918), .B(n3539), .Z(out[589]) );
  XNOR U1247 ( .A(n2921), .B(n3542), .Z(out[588]) );
  XNOR U1248 ( .A(n2924), .B(n3545), .Z(out[587]) );
  XNOR U1249 ( .A(n2931), .B(n3550), .Z(out[585]) );
  ANDN U1250 ( .B(n2991), .A(n2724), .Z(n2990) );
  ANDN U1251 ( .B(n2993), .A(n2728), .Z(n2992) );
  ANDN U1252 ( .B(n3035), .A(n2788), .Z(n3034) );
  ANDN U1253 ( .B(n3042), .A(n2800), .Z(n3041) );
  ANDN U1254 ( .B(n3044), .A(n2804), .Z(n3043) );
  ANDN U1255 ( .B(n3099), .A(n2887), .Z(n3098) );
  ANDN U1256 ( .B(n3103), .A(n2895), .Z(n3102) );
  ANDN U1257 ( .B(n3105), .A(n2899), .Z(n3104) );
  NOR U1258 ( .A(n3281), .B(n2846), .Z(n3484) );
  NOR U1259 ( .A(n3285), .B(n2850), .Z(n3487) );
  NOR U1260 ( .A(n3288), .B(n2854), .Z(n3490) );
  NOR U1261 ( .A(n3380), .B(n2951), .Z(n3565) );
  NOR U1262 ( .A(n1041), .B(n4197), .Z(n4008) );
  ANDN U1263 ( .B(n4021), .A(n2246), .Z(n4019) );
  ANDN U1264 ( .B(n4024), .A(n2870), .Z(n4022) );
  ANDN U1265 ( .B(n4027), .A(n3197), .Z(n4025) );
  ANDN U1266 ( .B(n4042), .A(n4043), .Z(n4040) );
  XNOR U1267 ( .A(n11714), .B(n11713), .Z(n11295) );
  XNOR U1268 ( .A(n11903), .B(n11285), .Z(n11133) );
  XNOR U1269 ( .A(n11492), .B(n11491), .Z(n10171) );
  XNOR U1270 ( .A(n12140), .B(n12370), .Z(n11341) );
  XOR U1271 ( .A(n11718), .B(n11717), .Z(n10522) );
  XNOR U1272 ( .A(n12054), .B(n11472), .Z(n10705) );
  XOR U1273 ( .A(n12598), .B(n11522), .Z(n9616) );
  XOR U1274 ( .A(n12753), .B(n12514), .Z(n9918) );
  XNOR U1275 ( .A(n11202), .B(n11485), .Z(n10688) );
  XOR U1276 ( .A(n11887), .B(n11662), .Z(n10674) );
  XNOR U1277 ( .A(n10847), .B(n11657), .Z(n9889) );
  XOR U1278 ( .A(n11399), .B(n11398), .Z(n10045) );
  XOR U1279 ( .A(n10540), .B(n11332), .Z(n9108) );
  XOR U1280 ( .A(n11070), .B(n11848), .Z(n9188) );
  XOR U1281 ( .A(round_reg[718]), .B(n9456), .Z(n9485) );
  XOR U1282 ( .A(round_reg[704]), .B(n10518), .Z(n8238) );
  XOR U1283 ( .A(round_reg[119]), .B(n11409), .Z(n8845) );
  XOR U1284 ( .A(round_reg[731]), .B(n10601), .Z(n7443) );
  XNOR U1285 ( .A(round_reg[744]), .B(n9632), .Z(n6952) );
  XOR U1286 ( .A(round_reg[1185]), .B(n10496), .Z(n6611) );
  XOR U1287 ( .A(round_reg[236]), .B(n10796), .Z(n8912) );
  XOR U1288 ( .A(round_reg[1311]), .B(n9554), .Z(n7108) );
  XOR U1289 ( .A(round_reg[782]), .B(n10529), .Z(n7158) );
  XNOR U1290 ( .A(round_reg[525]), .B(n10527), .Z(n8213) );
  NOR U1291 ( .A(n9001), .B(n6636), .Z(n8999) );
  NOR U1292 ( .A(n9173), .B(n8000), .Z(n9171) );
  XNOR U1293 ( .A(n6077), .B(n6076), .Z(n5585) );
  XNOR U1294 ( .A(n6083), .B(n6082), .Z(n5590) );
  XNOR U1295 ( .A(n6089), .B(n6088), .Z(n5595) );
  ANDN U1296 ( .B(n10053), .A(n10054), .Z(n10850) );
  ANDN U1297 ( .B(n10315), .A(n10314), .Z(n10387) );
  ANDN U1298 ( .B(n8317), .A(n10603), .Z(n10712) );
  NOR U1299 ( .A(n7124), .B(n6689), .Z(n9085) );
  ANDN U1300 ( .B(n10825), .A(n10824), .Z(n11909) );
  NOR U1301 ( .A(n7310), .B(n7311), .Z(n8361) );
  ANDN U1302 ( .B(n8794), .A(n8867), .Z(n8866) );
  ANDN U1303 ( .B(n7964), .A(n7963), .Z(n10924) );
  ANDN U1304 ( .B(n7121), .A(n7197), .Z(n7196) );
  NOR U1305 ( .A(n7561), .B(n7451), .Z(n7560) );
  NOR U1306 ( .A(n7613), .B(n7541), .Z(n7612) );
  NOR U1307 ( .A(n7683), .B(n7594), .Z(n7682) );
  NOR U1308 ( .A(n7820), .B(n7738), .Z(n7819) );
  NOR U1309 ( .A(n7887), .B(n7886), .Z(n7885) );
  ANDN U1310 ( .B(n7956), .A(n7957), .Z(n7954) );
  ANDN U1311 ( .B(n9293), .A(n10139), .Z(n12639) );
  ANDN U1312 ( .B(n8112), .A(n8113), .Z(n8111) );
  ANDN U1313 ( .B(n7801), .A(n7802), .Z(n7799) );
  ANDN U1314 ( .B(n6654), .A(n6655), .Z(n6652) );
  XNOR U1315 ( .A(n12029), .B(n12030), .Z(n3687) );
  ANDN U1316 ( .B(n7211), .A(n7209), .Z(n8262) );
  ANDN U1317 ( .B(n7239), .A(n7237), .Z(n8314) );
  ANDN U1318 ( .B(n7850), .A(n7851), .Z(n7848) );
  ANDN U1319 ( .B(n7917), .A(n7918), .Z(n7915) );
  ANDN U1320 ( .B(n8030), .A(n8028), .Z(n9029) );
  ANDN U1321 ( .B(n10200), .A(n7840), .Z(n10745) );
  ANDN U1322 ( .B(n6506), .A(n8711), .Z(n8709) );
  NOR U1323 ( .A(n6767), .B(n6768), .Z(n7256) );
  XNOR U1324 ( .A(n7669), .B(n7670), .Z(n4294) );
  NOR U1325 ( .A(n8611), .B(n8610), .Z(n8608) );
  NOR U1326 ( .A(n7040), .B(n7041), .Z(n9285) );
  NOR U1327 ( .A(n7063), .B(n7064), .Z(n10084) );
  NOR U1328 ( .A(n7086), .B(n7087), .Z(n10965) );
  ANDN U1329 ( .B(n7649), .A(n7650), .Z(n7647) );
  NOR U1330 ( .A(n8898), .B(n8899), .Z(n10836) );
  XOR U1331 ( .A(n6258), .B(n8071), .Z(n1951) );
  XOR U1332 ( .A(n6285), .B(n8304), .Z(n1658) );
  ANDN U1333 ( .B(n10594), .A(n10681), .Z(n10680) );
  XOR U1334 ( .A(n6346), .B(n9221), .Z(n1732) );
  ANDN U1335 ( .B(n4520), .A(n4521), .Z(n4518) );
  ANDN U1336 ( .B(n4536), .A(n4537), .Z(n4534) );
  ANDN U1337 ( .B(n4540), .A(n4541), .Z(n4538) );
  ANDN U1338 ( .B(n4610), .A(n4611), .Z(n4603) );
  ANDN U1339 ( .B(n4614), .A(n4615), .Z(n4612) );
  ANDN U1340 ( .B(n4618), .A(n4619), .Z(n4616) );
  ANDN U1341 ( .B(n4637), .A(n4638), .Z(n4630) );
  ANDN U1342 ( .B(n4658), .A(n4659), .Z(n4654) );
  ANDN U1343 ( .B(n5017), .A(n4786), .Z(n5015) );
  ANDN U1344 ( .B(n5667), .A(n5668), .Z(n5665) );
  ANDN U1345 ( .B(n5728), .A(n1050), .Z(n5727) );
  ANDN U1346 ( .B(n5789), .A(n1138), .Z(n5788) );
  ANDN U1347 ( .B(n6239), .A(n5890), .Z(n6235) );
  ANDN U1348 ( .B(n6249), .A(n5907), .Z(n6245) );
  ANDN U1349 ( .B(n6254), .A(n5909), .Z(n6250) );
  ANDN U1350 ( .B(n6281), .A(n5917), .Z(n6277) );
  ANDN U1351 ( .B(n6286), .A(n5919), .Z(n6282) );
  ANDN U1352 ( .B(n1357), .A(n1358), .Z(n1355) );
  ANDN U1353 ( .B(n1373), .A(n1374), .Z(n1371) );
  ANDN U1354 ( .B(n1377), .A(n1378), .Z(n1375) );
  ANDN U1355 ( .B(n1381), .A(n1382), .Z(n1379) );
  ANDN U1356 ( .B(n1385), .A(n1386), .Z(n1383) );
  XNOR U1357 ( .A(n1439), .B(n1440), .Z(out[909]) );
  ANDN U1358 ( .B(n1601), .A(n1398), .Z(n1600) );
  ANDN U1359 ( .B(n1603), .A(n1402), .Z(n1602) );
  NOR U1360 ( .A(n1681), .B(n1989), .Z(n1986) );
  NOR U1361 ( .A(n1701), .B(n2006), .Z(n2003) );
  NOR U1362 ( .A(n1711), .B(n2014), .Z(n2011) );
  NOR U1363 ( .A(n1733), .B(n2029), .Z(n2026) );
  NOR U1364 ( .A(n1738), .B(n2033), .Z(n2030) );
  NOR U1365 ( .A(n1748), .B(n2041), .Z(n2038) );
  NOR U1366 ( .A(n1758), .B(n2053), .Z(n2050) );
  XNOR U1367 ( .A(n2861), .B(n2862), .Z(out[601]) );
  ANDN U1368 ( .B(n3046), .A(n2808), .Z(n3045) );
  ANDN U1369 ( .B(n3101), .A(n2891), .Z(n3100) );
  NOR U1370 ( .A(n3274), .B(n2838), .Z(n3479) );
  NOR U1371 ( .A(n3331), .B(n3533), .Z(n3531) );
  NOR U1372 ( .A(n3335), .B(n3536), .Z(n3534) );
  NOR U1373 ( .A(n3340), .B(n3539), .Z(n3537) );
  NOR U1374 ( .A(n3345), .B(n3542), .Z(n3540) );
  NOR U1375 ( .A(n3354), .B(n3545), .Z(n3543) );
  NOR U1376 ( .A(n3364), .B(n3550), .Z(n3548) );
  NOR U1377 ( .A(n3368), .B(n2935), .Z(n3551) );
  ANDN U1378 ( .B(n3898), .A(n3350), .Z(n3897) );
  ANDN U1379 ( .B(n3900), .A(n3392), .Z(n3899) );
  ANDN U1380 ( .B(n3950), .A(n3951), .Z(n3949) );
  ANDN U1381 ( .B(n3953), .A(n3954), .Z(n3952) );
  NOR U1382 ( .A(n3525), .B(n4217), .Z(n4030) );
  ANDN U1383 ( .B(n4038), .A(n4039), .Z(n4036) );
  NOR U1384 ( .A(n3948), .B(n1348), .Z(n4155) );
  ANDN U1385 ( .B(n1719), .A(n3983), .Z(n4187) );
  NOR U1386 ( .A(n4021), .B(n2196), .Z(n4208) );
  ANDN U1387 ( .B(n2249), .A(n4024), .Z(n4210) );
  NOR U1388 ( .A(n4027), .B(n2323), .Z(n4213) );
  ANDN U1389 ( .B(n2826), .A(n4055), .Z(n4237) );
  NOR U1390 ( .A(n4058), .B(n2873), .Z(n4239) );
  NOR U1391 ( .A(n4066), .B(n2955), .Z(n4244) );
  NOR U1392 ( .A(n4069), .B(n2987), .Z(n4246) );
  NOR U1393 ( .A(n4072), .B(n3019), .Z(n4248) );
  ANDN U1394 ( .B(n1911), .A(n1912), .Z(n1909) );
  ANDN U1395 ( .B(n2001), .A(n2002), .Z(n1999) );
  ANDN U1396 ( .B(n2044), .A(n2045), .Z(n2042) );
  XNOR U1397 ( .A(n2618), .B(n2619), .Z(out[64]) );
  XNOR U1398 ( .A(n3130), .B(n3131), .Z(out[51]) );
  XNOR U1399 ( .A(n3158), .B(n3159), .Z(out[50]) );
  ANDN U1400 ( .B(n3497), .A(n3498), .Z(n3495) );
  ANDN U1401 ( .B(n3529), .A(n3530), .Z(n3527) );
  ANDN U1402 ( .B(n3561), .A(n3562), .Z(n3559) );
  ANDN U1403 ( .B(n3595), .A(n3596), .Z(n3593) );
  ANDN U1404 ( .B(n3639), .A(n3640), .Z(n3637) );
  ANDN U1405 ( .B(n3683), .A(n1046), .Z(n3682) );
  ANDN U1406 ( .B(n3726), .A(n1090), .Z(n3725) );
  ANDN U1407 ( .B(n3813), .A(n1178), .Z(n3812) );
  ANDN U1408 ( .B(n3855), .A(n1222), .Z(n3854) );
  ANDN U1409 ( .B(n1041), .A(n1042), .Z(n1039) );
  XOR U1410 ( .A(n1039), .B(n1040), .Z(out[9]) );
  XNOR U1411 ( .A(n1043), .B(n1044), .Z(out[99]) );
  AND U1412 ( .A(n1045), .B(n1046), .Z(n1043) );
  XNOR U1413 ( .A(n1047), .B(n1048), .Z(out[999]) );
  AND U1414 ( .A(n1049), .B(n1050), .Z(n1047) );
  XNOR U1415 ( .A(n1051), .B(n1052), .Z(out[998]) );
  AND U1416 ( .A(n1053), .B(n1054), .Z(n1051) );
  XNOR U1417 ( .A(n1055), .B(n1056), .Z(out[997]) );
  AND U1418 ( .A(n1057), .B(n1058), .Z(n1055) );
  XNOR U1419 ( .A(n1059), .B(n1060), .Z(out[996]) );
  AND U1420 ( .A(n1061), .B(n1062), .Z(n1059) );
  XNOR U1421 ( .A(n1063), .B(n1064), .Z(out[995]) );
  AND U1422 ( .A(n1065), .B(n1066), .Z(n1063) );
  XNOR U1423 ( .A(n1067), .B(n1068), .Z(out[994]) );
  AND U1424 ( .A(n1069), .B(n1070), .Z(n1067) );
  XNOR U1425 ( .A(n1071), .B(n1072), .Z(out[993]) );
  AND U1426 ( .A(n1073), .B(n1074), .Z(n1071) );
  XOR U1427 ( .A(n1075), .B(n1076), .Z(out[992]) );
  AND U1428 ( .A(n1077), .B(n1078), .Z(n1075) );
  XNOR U1429 ( .A(n1079), .B(n1080), .Z(out[991]) );
  AND U1430 ( .A(n1081), .B(n1082), .Z(n1079) );
  XNOR U1431 ( .A(n1083), .B(n1084), .Z(out[990]) );
  AND U1432 ( .A(n1085), .B(n1086), .Z(n1083) );
  XNOR U1433 ( .A(n1087), .B(n1088), .Z(out[98]) );
  AND U1434 ( .A(n1089), .B(n1090), .Z(n1087) );
  XNOR U1435 ( .A(n1091), .B(n1092), .Z(out[989]) );
  AND U1436 ( .A(n1093), .B(n1094), .Z(n1091) );
  XNOR U1437 ( .A(n1095), .B(n1096), .Z(out[988]) );
  AND U1438 ( .A(n1097), .B(n1098), .Z(n1095) );
  XNOR U1439 ( .A(n1099), .B(n1100), .Z(out[987]) );
  AND U1440 ( .A(n1101), .B(n1102), .Z(n1099) );
  XNOR U1441 ( .A(n1103), .B(n1104), .Z(out[986]) );
  AND U1442 ( .A(n1105), .B(n1106), .Z(n1103) );
  XNOR U1443 ( .A(n1107), .B(n1108), .Z(out[985]) );
  AND U1444 ( .A(n1109), .B(n1110), .Z(n1107) );
  XNOR U1445 ( .A(n1111), .B(n1112), .Z(out[984]) );
  AND U1446 ( .A(n1113), .B(n1114), .Z(n1111) );
  XNOR U1447 ( .A(n1115), .B(n1116), .Z(out[983]) );
  AND U1448 ( .A(n1117), .B(n1118), .Z(n1115) );
  XNOR U1449 ( .A(n1119), .B(n1120), .Z(out[982]) );
  AND U1450 ( .A(n1121), .B(n1122), .Z(n1119) );
  XNOR U1451 ( .A(n1123), .B(n1124), .Z(out[981]) );
  AND U1452 ( .A(n1125), .B(n1126), .Z(n1123) );
  XNOR U1453 ( .A(n1127), .B(n1128), .Z(out[980]) );
  AND U1454 ( .A(n1129), .B(n1130), .Z(n1127) );
  XOR U1455 ( .A(n1131), .B(n1132), .Z(out[97]) );
  ANDN U1456 ( .B(n1133), .A(n1134), .Z(n1131) );
  XNOR U1457 ( .A(n1135), .B(n1136), .Z(out[979]) );
  AND U1458 ( .A(n1137), .B(n1138), .Z(n1135) );
  XNOR U1459 ( .A(n1139), .B(n1140), .Z(out[978]) );
  AND U1460 ( .A(n1141), .B(n1142), .Z(n1139) );
  XNOR U1461 ( .A(n1143), .B(n1144), .Z(out[977]) );
  AND U1462 ( .A(n1145), .B(n1146), .Z(n1143) );
  XNOR U1463 ( .A(n1147), .B(n1148), .Z(out[976]) );
  AND U1464 ( .A(n1149), .B(n1150), .Z(n1147) );
  XNOR U1465 ( .A(n1151), .B(n1152), .Z(out[975]) );
  AND U1466 ( .A(n1153), .B(n1154), .Z(n1151) );
  XNOR U1467 ( .A(n1155), .B(n1156), .Z(out[974]) );
  AND U1468 ( .A(n1157), .B(n1158), .Z(n1155) );
  XOR U1469 ( .A(n1159), .B(n1160), .Z(out[973]) );
  AND U1470 ( .A(n1161), .B(n1162), .Z(n1159) );
  XNOR U1471 ( .A(n1163), .B(n1164), .Z(out[972]) );
  ANDN U1472 ( .B(n1165), .A(n1166), .Z(n1163) );
  XNOR U1473 ( .A(n1167), .B(n1168), .Z(out[971]) );
  ANDN U1474 ( .B(n1169), .A(n1170), .Z(n1167) );
  XNOR U1475 ( .A(n1171), .B(n1172), .Z(out[970]) );
  AND U1476 ( .A(n1173), .B(n1174), .Z(n1171) );
  XOR U1477 ( .A(n1175), .B(n1176), .Z(out[96]) );
  AND U1478 ( .A(n1177), .B(n1178), .Z(n1175) );
  XNOR U1479 ( .A(n1179), .B(n1180), .Z(out[969]) );
  ANDN U1480 ( .B(n1181), .A(n1182), .Z(n1179) );
  XOR U1481 ( .A(n1183), .B(n1184), .Z(out[968]) );
  XNOR U1482 ( .A(n1187), .B(n1188), .Z(out[967]) );
  XNOR U1483 ( .A(n1191), .B(n1192), .Z(out[966]) );
  ANDN U1484 ( .B(n1193), .A(n1194), .Z(n1191) );
  XNOR U1485 ( .A(n1195), .B(n1196), .Z(out[965]) );
  ANDN U1486 ( .B(n1197), .A(n1198), .Z(n1195) );
  XNOR U1487 ( .A(n1199), .B(n1200), .Z(out[964]) );
  ANDN U1488 ( .B(n1201), .A(n1202), .Z(n1199) );
  XNOR U1489 ( .A(n1203), .B(n1204), .Z(out[963]) );
  ANDN U1490 ( .B(n1205), .A(n1206), .Z(n1203) );
  XNOR U1491 ( .A(n1207), .B(n1208), .Z(out[962]) );
  ANDN U1492 ( .B(n1209), .A(n1210), .Z(n1207) );
  XNOR U1493 ( .A(n1211), .B(n1212), .Z(out[961]) );
  AND U1494 ( .A(n1213), .B(n1214), .Z(n1211) );
  XNOR U1495 ( .A(n1215), .B(n1216), .Z(out[960]) );
  ANDN U1496 ( .B(n1217), .A(n1218), .Z(n1215) );
  XOR U1497 ( .A(n1219), .B(n1220), .Z(out[95]) );
  AND U1498 ( .A(n1221), .B(n1222), .Z(n1219) );
  ANDN U1499 ( .B(n1225), .A(n1226), .Z(n1223) );
  ANDN U1500 ( .B(n1229), .A(n1230), .Z(n1227) );
  XNOR U1501 ( .A(n1231), .B(n1232), .Z(out[957]) );
  ANDN U1502 ( .B(n1233), .A(n1234), .Z(n1231) );
  XNOR U1503 ( .A(n1235), .B(n1236), .Z(out[956]) );
  ANDN U1504 ( .B(n1237), .A(n1238), .Z(n1235) );
  ANDN U1505 ( .B(n1240), .A(n1241), .Z(n1239) );
  XNOR U1506 ( .A(n1242), .B(n1243), .Z(out[954]) );
  ANDN U1507 ( .B(n1244), .A(n1245), .Z(n1242) );
  XNOR U1508 ( .A(n1246), .B(n1247), .Z(out[953]) );
  ANDN U1509 ( .B(n1248), .A(n1249), .Z(n1246) );
  XNOR U1510 ( .A(n1250), .B(n1251), .Z(out[952]) );
  ANDN U1511 ( .B(n1252), .A(n1253), .Z(n1250) );
  ANDN U1512 ( .B(n1255), .A(n1256), .Z(n1254) );
  XOR U1513 ( .A(n1257), .B(n1258), .Z(out[950]) );
  ANDN U1514 ( .B(n1259), .A(n1260), .Z(n1257) );
  XOR U1515 ( .A(n1261), .B(n1262), .Z(out[94]) );
  AND U1516 ( .A(n1263), .B(n1264), .Z(n1261) );
  ANDN U1517 ( .B(n1266), .A(n1267), .Z(n1265) );
  ANDN U1518 ( .B(n1269), .A(n1270), .Z(n1268) );
  XNOR U1519 ( .A(n1271), .B(n1272), .Z(out[947]) );
  ANDN U1520 ( .B(n1273), .A(n1274), .Z(n1271) );
  XOR U1521 ( .A(n1275), .B(n1276), .Z(out[946]) );
  ANDN U1522 ( .B(n1277), .A(n1278), .Z(n1275) );
  ANDN U1523 ( .B(n1280), .A(n1281), .Z(n1279) );
  AND U1524 ( .A(n1283), .B(n1284), .Z(n1282) );
  IV U1525 ( .A(n1285), .Z(n1284) );
  AND U1526 ( .A(n1287), .B(n1288), .Z(n1286) );
  IV U1527 ( .A(n1289), .Z(n1288) );
  AND U1528 ( .A(n1291), .B(n1292), .Z(n1290) );
  IV U1529 ( .A(n1293), .Z(n1292) );
  AND U1530 ( .A(n1295), .B(n1296), .Z(n1294) );
  IV U1531 ( .A(n1297), .Z(n1296) );
  AND U1532 ( .A(n1299), .B(n1300), .Z(n1298) );
  IV U1533 ( .A(n1301), .Z(n1300) );
  XOR U1534 ( .A(n1302), .B(n1303), .Z(out[93]) );
  AND U1535 ( .A(n1304), .B(n1305), .Z(n1302) );
  XNOR U1536 ( .A(n1306), .B(n1307), .Z(out[939]) );
  AND U1537 ( .A(n1312), .B(n1313), .Z(n1310) );
  IV U1538 ( .A(n1314), .Z(n1313) );
  AND U1539 ( .A(n1317), .B(n1318), .Z(n1315) );
  IV U1540 ( .A(n1319), .Z(n1318) );
  XNOR U1541 ( .A(n1320), .B(n1321), .Z(out[936]) );
  NOR U1542 ( .A(n1326), .B(n1327), .Z(n1324) );
  ANDN U1543 ( .B(n1330), .A(n1331), .Z(n1328) );
  ANDN U1544 ( .B(n1333), .A(n1334), .Z(n1332) );
  XNOR U1545 ( .A(n1335), .B(n1336), .Z(out[932]) );
  XNOR U1546 ( .A(n1339), .B(n1340), .Z(out[931]) );
  XOR U1547 ( .A(n1343), .B(n1344), .Z(out[930]) );
  XNOR U1548 ( .A(n1347), .B(n1348), .Z(out[92]) );
  AND U1549 ( .A(n1349), .B(n1350), .Z(n1347) );
  XOR U1550 ( .A(n1351), .B(n1352), .Z(out[929]) );
  XNOR U1551 ( .A(n1355), .B(n1356), .Z(out[928]) );
  XNOR U1552 ( .A(n1359), .B(n1360), .Z(out[927]) );
  XNOR U1553 ( .A(n1363), .B(n1364), .Z(out[926]) );
  XNOR U1554 ( .A(n1367), .B(n1368), .Z(out[925]) );
  XNOR U1555 ( .A(n1371), .B(n1372), .Z(out[924]) );
  XOR U1556 ( .A(n1375), .B(n1376), .Z(out[923]) );
  XOR U1557 ( .A(n1379), .B(n1380), .Z(out[922]) );
  XNOR U1558 ( .A(n1383), .B(n1384), .Z(out[921]) );
  XNOR U1559 ( .A(n1387), .B(n1388), .Z(out[920]) );
  AND U1560 ( .A(n1389), .B(n1390), .Z(n1387) );
  XOR U1561 ( .A(n1391), .B(n1392), .Z(out[91]) );
  AND U1562 ( .A(n1393), .B(n1394), .Z(n1391) );
  XOR U1563 ( .A(n1395), .B(n1396), .Z(out[919]) );
  AND U1564 ( .A(n1397), .B(n1398), .Z(n1395) );
  XOR U1565 ( .A(n1399), .B(n1400), .Z(out[918]) );
  AND U1566 ( .A(n1401), .B(n1402), .Z(n1399) );
  XOR U1567 ( .A(n1403), .B(n1404), .Z(out[917]) );
  AND U1568 ( .A(n1405), .B(n1406), .Z(n1403) );
  XOR U1569 ( .A(n1407), .B(n1408), .Z(out[916]) );
  AND U1570 ( .A(n1409), .B(n1410), .Z(n1407) );
  XOR U1571 ( .A(n1411), .B(n1412), .Z(out[915]) );
  AND U1572 ( .A(n1413), .B(n1414), .Z(n1411) );
  XNOR U1573 ( .A(n1415), .B(n1416), .Z(out[914]) );
  ANDN U1574 ( .B(n1417), .A(n1418), .Z(n1415) );
  XNOR U1575 ( .A(n1419), .B(n1420), .Z(out[913]) );
  XNOR U1576 ( .A(n1423), .B(n1424), .Z(out[912]) );
  AND U1577 ( .A(n1425), .B(n1426), .Z(n1423) );
  XNOR U1578 ( .A(n1427), .B(n1428), .Z(out[911]) );
  AND U1579 ( .A(n1429), .B(n1430), .Z(n1427) );
  XNOR U1580 ( .A(n1431), .B(n1432), .Z(out[910]) );
  AND U1581 ( .A(n1433), .B(n1434), .Z(n1431) );
  XOR U1582 ( .A(n1435), .B(n1436), .Z(out[90]) );
  AND U1583 ( .A(n1437), .B(n1438), .Z(n1435) );
  ANDN U1584 ( .B(n1441), .A(n1442), .Z(n1439) );
  XNOR U1585 ( .A(n1443), .B(n1444), .Z(out[908]) );
  ANDN U1586 ( .B(n1445), .A(n1446), .Z(n1443) );
  XNOR U1587 ( .A(n1447), .B(n1448), .Z(out[907]) );
  ANDN U1588 ( .B(n1449), .A(n1450), .Z(n1447) );
  XNOR U1589 ( .A(n1451), .B(n1452), .Z(out[906]) );
  AND U1590 ( .A(n1453), .B(n1454), .Z(n1451) );
  XNOR U1591 ( .A(n1455), .B(n1456), .Z(out[905]) );
  AND U1592 ( .A(n1457), .B(n1458), .Z(n1455) );
  XNOR U1593 ( .A(n1459), .B(n1460), .Z(out[904]) );
  AND U1594 ( .A(n1461), .B(n1462), .Z(n1459) );
  XNOR U1595 ( .A(n1463), .B(n1464), .Z(out[903]) );
  ANDN U1596 ( .B(n1465), .A(n1466), .Z(n1463) );
  XNOR U1597 ( .A(n1467), .B(n1468), .Z(out[902]) );
  ANDN U1598 ( .B(n1469), .A(n1470), .Z(n1467) );
  XNOR U1599 ( .A(n1471), .B(n1472), .Z(out[901]) );
  ANDN U1600 ( .B(n1473), .A(n1474), .Z(n1471) );
  XNOR U1601 ( .A(n1475), .B(n1476), .Z(out[900]) );
  ANDN U1602 ( .B(n1477), .A(n1478), .Z(n1475) );
  XNOR U1603 ( .A(n1479), .B(n1480), .Z(out[8]) );
  NOR U1604 ( .A(n1481), .B(n1482), .Z(n1479) );
  XOR U1605 ( .A(n1483), .B(n1484), .Z(out[89]) );
  AND U1606 ( .A(n1485), .B(n1486), .Z(n1483) );
  XNOR U1607 ( .A(n1487), .B(n1488), .Z(out[899]) );
  ANDN U1608 ( .B(n1489), .A(n1490), .Z(n1487) );
  XNOR U1609 ( .A(n1491), .B(n1492), .Z(out[898]) );
  ANDN U1610 ( .B(n1493), .A(n1494), .Z(n1491) );
  XNOR U1611 ( .A(n1495), .B(n1496), .Z(out[897]) );
  ANDN U1612 ( .B(n1497), .A(n1498), .Z(n1495) );
  XNOR U1613 ( .A(n1499), .B(n1500), .Z(out[896]) );
  ANDN U1614 ( .B(n1501), .A(n1502), .Z(n1499) );
  XNOR U1615 ( .A(n1503), .B(n1225), .Z(out[895]) );
  AND U1616 ( .A(n1226), .B(n1504), .Z(n1503) );
  XNOR U1617 ( .A(n1505), .B(n1229), .Z(out[894]) );
  AND U1618 ( .A(n1230), .B(n1506), .Z(n1505) );
  XNOR U1619 ( .A(n1507), .B(n1233), .Z(out[893]) );
  AND U1620 ( .A(n1234), .B(n1508), .Z(n1507) );
  XNOR U1621 ( .A(n1509), .B(n1237), .Z(out[892]) );
  AND U1622 ( .A(n1238), .B(n1510), .Z(n1509) );
  XNOR U1623 ( .A(n1511), .B(n1240), .Z(out[891]) );
  AND U1624 ( .A(n1241), .B(n1512), .Z(n1511) );
  XNOR U1625 ( .A(n1513), .B(n1244), .Z(out[890]) );
  AND U1626 ( .A(n1245), .B(n1514), .Z(n1513) );
  XOR U1627 ( .A(n1515), .B(n1516), .Z(out[88]) );
  AND U1628 ( .A(n1517), .B(n1518), .Z(n1515) );
  XNOR U1629 ( .A(n1519), .B(n1248), .Z(out[889]) );
  AND U1630 ( .A(n1249), .B(n1520), .Z(n1519) );
  XNOR U1631 ( .A(n1521), .B(n1252), .Z(out[888]) );
  AND U1632 ( .A(n1253), .B(n1522), .Z(n1521) );
  XNOR U1633 ( .A(n1523), .B(n1255), .Z(out[887]) );
  AND U1634 ( .A(n1256), .B(n1524), .Z(n1523) );
  XNOR U1635 ( .A(n1525), .B(n1259), .Z(out[886]) );
  AND U1636 ( .A(n1260), .B(n1526), .Z(n1525) );
  XNOR U1637 ( .A(n1527), .B(n1266), .Z(out[885]) );
  AND U1638 ( .A(n1267), .B(n1528), .Z(n1527) );
  XNOR U1639 ( .A(n1529), .B(n1269), .Z(out[884]) );
  AND U1640 ( .A(n1270), .B(n1530), .Z(n1529) );
  XNOR U1641 ( .A(n1531), .B(n1273), .Z(out[883]) );
  AND U1642 ( .A(n1274), .B(n1532), .Z(n1531) );
  XNOR U1643 ( .A(n1533), .B(n1277), .Z(out[882]) );
  AND U1644 ( .A(n1278), .B(n1534), .Z(n1533) );
  XNOR U1645 ( .A(n1535), .B(n1280), .Z(out[881]) );
  AND U1646 ( .A(n1281), .B(n1536), .Z(n1535) );
  XOR U1647 ( .A(n1537), .B(n1285), .Z(out[880]) );
  XOR U1648 ( .A(n1539), .B(n1540), .Z(out[87]) );
  AND U1649 ( .A(n1541), .B(n1542), .Z(n1539) );
  XOR U1650 ( .A(n1543), .B(n1289), .Z(out[879]) );
  XOR U1651 ( .A(n1545), .B(n1293), .Z(out[878]) );
  XOR U1652 ( .A(n1547), .B(n1297), .Z(out[877]) );
  XOR U1653 ( .A(n1549), .B(n1301), .Z(out[876]) );
  XOR U1654 ( .A(n1551), .B(n1309), .Z(out[875]) );
  NOR U1655 ( .A(n1552), .B(n1308), .Z(n1551) );
  XOR U1656 ( .A(n1553), .B(n1314), .Z(out[874]) );
  XOR U1657 ( .A(n1555), .B(n1319), .Z(out[873]) );
  XOR U1658 ( .A(n1557), .B(n1323), .Z(out[872]) );
  NOR U1659 ( .A(n1322), .B(n1558), .Z(n1557) );
  XOR U1660 ( .A(n1559), .B(n1327), .Z(out[871]) );
  AND U1661 ( .A(n1326), .B(n1560), .Z(n1559) );
  IV U1662 ( .A(n1561), .Z(n1326) );
  XNOR U1663 ( .A(n1562), .B(n1330), .Z(out[870]) );
  AND U1664 ( .A(n1331), .B(n1563), .Z(n1562) );
  XOR U1665 ( .A(n1564), .B(n1565), .Z(out[86]) );
  AND U1666 ( .A(n1566), .B(n1567), .Z(n1564) );
  XNOR U1667 ( .A(n1568), .B(n1333), .Z(out[869]) );
  AND U1668 ( .A(n1334), .B(n1569), .Z(n1568) );
  XOR U1669 ( .A(n1570), .B(n1338), .Z(out[868]) );
  NOR U1670 ( .A(n1571), .B(n1337), .Z(n1570) );
  XOR U1671 ( .A(n1572), .B(n1342), .Z(out[867]) );
  ANDN U1672 ( .B(n1573), .A(n1341), .Z(n1572) );
  XOR U1673 ( .A(n1574), .B(n1346), .Z(out[866]) );
  NOR U1674 ( .A(n1575), .B(n1345), .Z(n1574) );
  XOR U1675 ( .A(n1576), .B(n1354), .Z(out[865]) );
  NOR U1676 ( .A(n1577), .B(n1353), .Z(n1576) );
  XOR U1677 ( .A(n1578), .B(n1358), .Z(out[864]) );
  NOR U1678 ( .A(n1579), .B(n1357), .Z(n1578) );
  XOR U1679 ( .A(n1580), .B(n1362), .Z(out[863]) );
  NOR U1680 ( .A(n1581), .B(n1361), .Z(n1580) );
  XOR U1681 ( .A(n1582), .B(n1366), .Z(out[862]) );
  NOR U1682 ( .A(n1583), .B(n1365), .Z(n1582) );
  XOR U1683 ( .A(n1584), .B(n1370), .Z(out[861]) );
  NOR U1684 ( .A(n1585), .B(n1369), .Z(n1584) );
  XOR U1685 ( .A(n1586), .B(n1374), .Z(out[860]) );
  NOR U1686 ( .A(n1587), .B(n1373), .Z(n1586) );
  XOR U1687 ( .A(n1588), .B(n1589), .Z(out[85]) );
  AND U1688 ( .A(n1590), .B(n1591), .Z(n1588) );
  XOR U1689 ( .A(n1592), .B(n1378), .Z(out[859]) );
  ANDN U1690 ( .B(n1593), .A(n1377), .Z(n1592) );
  XOR U1691 ( .A(n1594), .B(n1382), .Z(out[858]) );
  ANDN U1692 ( .B(n1595), .A(n1381), .Z(n1594) );
  XOR U1693 ( .A(n1596), .B(n1386), .Z(out[857]) );
  ANDN U1694 ( .B(n1597), .A(n1385), .Z(n1596) );
  XNOR U1695 ( .A(n1598), .B(n1389), .Z(out[856]) );
  XNOR U1696 ( .A(n1600), .B(n1397), .Z(out[855]) );
  XNOR U1697 ( .A(n1602), .B(n1401), .Z(out[854]) );
  XNOR U1698 ( .A(n1604), .B(n1405), .Z(out[853]) );
  XNOR U1699 ( .A(n1606), .B(n1409), .Z(out[852]) );
  XNOR U1700 ( .A(n1608), .B(n1413), .Z(out[851]) );
  XNOR U1701 ( .A(n1610), .B(n1417), .Z(out[850]) );
  AND U1702 ( .A(n1418), .B(n1611), .Z(n1610) );
  XOR U1703 ( .A(n1612), .B(n1613), .Z(out[84]) );
  AND U1704 ( .A(n1614), .B(n1615), .Z(n1612) );
  XOR U1705 ( .A(n1616), .B(n1422), .Z(out[849]) );
  NOR U1706 ( .A(n1617), .B(n1421), .Z(n1616) );
  XNOR U1707 ( .A(n1618), .B(n1426), .Z(out[848]) );
  ANDN U1708 ( .B(n1619), .A(n1425), .Z(n1618) );
  XNOR U1709 ( .A(n1620), .B(n1430), .Z(out[847]) );
  NOR U1710 ( .A(n1621), .B(n1429), .Z(n1620) );
  XNOR U1711 ( .A(n1622), .B(n1434), .Z(out[846]) );
  NOR U1712 ( .A(n1623), .B(n1433), .Z(n1622) );
  XNOR U1713 ( .A(n1624), .B(n1441), .Z(out[845]) );
  AND U1714 ( .A(n1442), .B(n1625), .Z(n1624) );
  XNOR U1715 ( .A(n1626), .B(n1445), .Z(out[844]) );
  ANDN U1716 ( .B(n1446), .A(n1627), .Z(n1626) );
  XNOR U1717 ( .A(n1628), .B(n1449), .Z(out[843]) );
  AND U1718 ( .A(n1450), .B(n1629), .Z(n1628) );
  XNOR U1719 ( .A(n1630), .B(n1453), .Z(out[842]) );
  XNOR U1720 ( .A(n1632), .B(n1457), .Z(out[841]) );
  XNOR U1721 ( .A(n1634), .B(n1461), .Z(out[840]) );
  XNOR U1722 ( .A(n1636), .B(n1637), .Z(out[83]) );
  AND U1723 ( .A(n1638), .B(n1639), .Z(n1636) );
  XNOR U1724 ( .A(n1640), .B(n1465), .Z(out[839]) );
  AND U1725 ( .A(n1466), .B(n1641), .Z(n1640) );
  XNOR U1726 ( .A(n1642), .B(n1469), .Z(out[838]) );
  AND U1727 ( .A(n1470), .B(n1643), .Z(n1642) );
  XNOR U1728 ( .A(n1644), .B(n1473), .Z(out[837]) );
  AND U1729 ( .A(n1474), .B(n1645), .Z(n1644) );
  XNOR U1730 ( .A(n1646), .B(n1477), .Z(out[836]) );
  AND U1731 ( .A(n1478), .B(n1647), .Z(n1646) );
  XNOR U1732 ( .A(n1648), .B(n1489), .Z(out[835]) );
  AND U1733 ( .A(n1490), .B(n1649), .Z(n1648) );
  XNOR U1734 ( .A(n1650), .B(n1493), .Z(out[834]) );
  AND U1735 ( .A(n1494), .B(n1651), .Z(n1650) );
  XNOR U1736 ( .A(n1652), .B(n1497), .Z(out[833]) );
  AND U1737 ( .A(n1498), .B(n1653), .Z(n1652) );
  XNOR U1738 ( .A(n1654), .B(n1501), .Z(out[832]) );
  AND U1739 ( .A(n1502), .B(n1655), .Z(n1654) );
  XNOR U1740 ( .A(n1656), .B(n1226), .Z(out[831]) );
  XOR U1741 ( .A(n1657), .B(n1658), .Z(n1226) );
  AND U1742 ( .A(n1659), .B(n1660), .Z(n1656) );
  XNOR U1743 ( .A(n1661), .B(n1230), .Z(out[830]) );
  XOR U1744 ( .A(n1662), .B(n1663), .Z(n1230) );
  XNOR U1745 ( .A(n1665), .B(n1666), .Z(out[82]) );
  AND U1746 ( .A(n1667), .B(n1668), .Z(n1665) );
  XNOR U1747 ( .A(n1669), .B(n1234), .Z(out[829]) );
  XOR U1748 ( .A(n1670), .B(n1671), .Z(n1234) );
  XNOR U1749 ( .A(n1673), .B(n1238), .Z(out[828]) );
  XOR U1750 ( .A(n1674), .B(n1675), .Z(n1238) );
  AND U1751 ( .A(n1676), .B(n1677), .Z(n1673) );
  XNOR U1752 ( .A(n1678), .B(n1241), .Z(out[827]) );
  XNOR U1753 ( .A(n1679), .B(n1680), .Z(n1241) );
  AND U1754 ( .A(n1681), .B(n1682), .Z(n1678) );
  XNOR U1755 ( .A(n1683), .B(n1245), .Z(out[826]) );
  XNOR U1756 ( .A(n1684), .B(n1685), .Z(n1245) );
  AND U1757 ( .A(n1686), .B(n1687), .Z(n1683) );
  XNOR U1758 ( .A(n1688), .B(n1249), .Z(out[825]) );
  XOR U1759 ( .A(n1689), .B(n1690), .Z(n1249) );
  AND U1760 ( .A(n1691), .B(n1692), .Z(n1688) );
  XNOR U1761 ( .A(n1693), .B(n1253), .Z(out[824]) );
  XOR U1762 ( .A(n1694), .B(n1695), .Z(n1253) );
  AND U1763 ( .A(n1696), .B(n1697), .Z(n1693) );
  XNOR U1764 ( .A(n1698), .B(n1256), .Z(out[823]) );
  XNOR U1765 ( .A(n1699), .B(n1700), .Z(n1256) );
  AND U1766 ( .A(n1701), .B(n1702), .Z(n1698) );
  XNOR U1767 ( .A(n1703), .B(n1260), .Z(out[822]) );
  XNOR U1768 ( .A(n1704), .B(n1705), .Z(n1260) );
  AND U1769 ( .A(n1706), .B(n1707), .Z(n1703) );
  XNOR U1770 ( .A(n1708), .B(n1267), .Z(out[821]) );
  XNOR U1771 ( .A(n1709), .B(n1710), .Z(n1267) );
  AND U1772 ( .A(n1711), .B(n1712), .Z(n1708) );
  XNOR U1773 ( .A(n1713), .B(n1270), .Z(out[820]) );
  XNOR U1774 ( .A(n1714), .B(n1715), .Z(n1270) );
  AND U1775 ( .A(n1716), .B(n1717), .Z(n1713) );
  XOR U1776 ( .A(n1718), .B(n1719), .Z(out[81]) );
  NOR U1777 ( .A(n1720), .B(n1721), .Z(n1718) );
  XNOR U1778 ( .A(n1722), .B(n1274), .Z(out[819]) );
  XOR U1779 ( .A(n1723), .B(n1724), .Z(n1274) );
  XNOR U1780 ( .A(n1726), .B(n1278), .Z(out[818]) );
  XOR U1781 ( .A(n1727), .B(n1728), .Z(n1278) );
  XNOR U1782 ( .A(n1730), .B(n1281), .Z(out[817]) );
  XOR U1783 ( .A(n1731), .B(n1732), .Z(n1281) );
  AND U1784 ( .A(n1733), .B(n1734), .Z(n1730) );
  XOR U1785 ( .A(n1735), .B(n1283), .Z(out[816]) );
  XNOR U1786 ( .A(n1736), .B(n1737), .Z(n1283) );
  AND U1787 ( .A(n1738), .B(n1739), .Z(n1735) );
  XOR U1788 ( .A(n1740), .B(n1287), .Z(out[815]) );
  XNOR U1789 ( .A(n1741), .B(n1742), .Z(n1287) );
  AND U1790 ( .A(n1743), .B(n1744), .Z(n1740) );
  XOR U1791 ( .A(n1745), .B(n1291), .Z(out[814]) );
  XNOR U1792 ( .A(n1746), .B(n1747), .Z(n1291) );
  AND U1793 ( .A(n1748), .B(n1749), .Z(n1745) );
  XOR U1794 ( .A(n1750), .B(n1295), .Z(out[813]) );
  XNOR U1795 ( .A(n1751), .B(n1752), .Z(n1295) );
  AND U1796 ( .A(n1753), .B(n1754), .Z(n1750) );
  XOR U1797 ( .A(n1755), .B(n1299), .Z(out[812]) );
  XNOR U1798 ( .A(n1756), .B(n1757), .Z(n1299) );
  AND U1799 ( .A(n1758), .B(n1759), .Z(n1755) );
  XOR U1800 ( .A(n1760), .B(n1308), .Z(out[811]) );
  XOR U1801 ( .A(n1761), .B(n1762), .Z(n1308) );
  AND U1802 ( .A(n1552), .B(n1763), .Z(n1760) );
  XOR U1803 ( .A(n1764), .B(n1312), .Z(out[810]) );
  XOR U1804 ( .A(n1765), .B(n1766), .Z(n1312) );
  AND U1805 ( .A(n1767), .B(n1768), .Z(n1764) );
  XNOR U1806 ( .A(n1769), .B(n1770), .Z(out[80]) );
  AND U1807 ( .A(n1771), .B(n1772), .Z(n1769) );
  XOR U1808 ( .A(n1773), .B(n1317), .Z(out[809]) );
  XOR U1809 ( .A(n1774), .B(n1775), .Z(n1317) );
  AND U1810 ( .A(n1776), .B(n1777), .Z(n1773) );
  XOR U1811 ( .A(n1778), .B(n1322), .Z(out[808]) );
  XOR U1812 ( .A(n1779), .B(n1780), .Z(n1322) );
  AND U1813 ( .A(n1558), .B(n1781), .Z(n1778) );
  XOR U1814 ( .A(n1782), .B(n1561), .Z(out[807]) );
  XOR U1815 ( .A(n1783), .B(n1784), .Z(n1561) );
  XNOR U1816 ( .A(n1786), .B(n1331), .Z(out[806]) );
  XNOR U1817 ( .A(n1787), .B(n1788), .Z(n1331) );
  XNOR U1818 ( .A(n1790), .B(n1334), .Z(out[805]) );
  XNOR U1819 ( .A(n1791), .B(n1792), .Z(n1334) );
  XOR U1820 ( .A(n1794), .B(n1337), .Z(out[804]) );
  XNOR U1821 ( .A(n1795), .B(n1796), .Z(n1337) );
  AND U1822 ( .A(n1571), .B(n1797), .Z(n1794) );
  XOR U1823 ( .A(n1798), .B(n1341), .Z(out[803]) );
  XOR U1824 ( .A(n1799), .B(n1800), .Z(n1341) );
  ANDN U1825 ( .B(n1801), .A(n1573), .Z(n1798) );
  XOR U1826 ( .A(n1802), .B(n1345), .Z(out[802]) );
  XOR U1827 ( .A(n1803), .B(n1804), .Z(n1345) );
  AND U1828 ( .A(n1575), .B(n1805), .Z(n1802) );
  XOR U1829 ( .A(n1806), .B(n1353), .Z(out[801]) );
  XOR U1830 ( .A(n1807), .B(n1808), .Z(n1353) );
  AND U1831 ( .A(n1577), .B(n1809), .Z(n1806) );
  XOR U1832 ( .A(n1810), .B(n1357), .Z(out[800]) );
  XOR U1833 ( .A(n1811), .B(n1812), .Z(n1357) );
  XNOR U1834 ( .A(n1814), .B(n1815), .Z(out[7]) );
  NOR U1835 ( .A(n1816), .B(n1817), .Z(n1814) );
  XNOR U1836 ( .A(n1818), .B(n1819), .Z(out[79]) );
  AND U1837 ( .A(n1820), .B(n1821), .Z(n1818) );
  XOR U1838 ( .A(n1822), .B(n1361), .Z(out[799]) );
  XOR U1839 ( .A(n1823), .B(n1824), .Z(n1361) );
  AND U1840 ( .A(n1581), .B(n1825), .Z(n1822) );
  XOR U1841 ( .A(n1826), .B(n1365), .Z(out[798]) );
  XOR U1842 ( .A(n1827), .B(n1828), .Z(n1365) );
  AND U1843 ( .A(n1583), .B(n1829), .Z(n1826) );
  XOR U1844 ( .A(n1830), .B(n1369), .Z(out[797]) );
  XOR U1845 ( .A(n1831), .B(n1832), .Z(n1369) );
  AND U1846 ( .A(n1585), .B(n1833), .Z(n1830) );
  XOR U1847 ( .A(n1834), .B(n1373), .Z(out[796]) );
  XOR U1848 ( .A(n1835), .B(n1836), .Z(n1373) );
  AND U1849 ( .A(n1587), .B(n1837), .Z(n1834) );
  XOR U1850 ( .A(n1838), .B(n1377), .Z(out[795]) );
  XOR U1851 ( .A(n1839), .B(n1840), .Z(n1377) );
  NOR U1852 ( .A(n1841), .B(n1593), .Z(n1838) );
  XOR U1853 ( .A(n1842), .B(n1381), .Z(out[794]) );
  XOR U1854 ( .A(n1843), .B(n1844), .Z(n1381) );
  NOR U1855 ( .A(n1845), .B(n1595), .Z(n1842) );
  XOR U1856 ( .A(n1846), .B(n1385), .Z(out[793]) );
  XOR U1857 ( .A(n1847), .B(n1848), .Z(n1385) );
  AND U1858 ( .A(n1849), .B(n1850), .Z(n1846) );
  XOR U1859 ( .A(n1851), .B(n1390), .Z(out[792]) );
  XOR U1860 ( .A(n1852), .B(n1853), .Z(n1390) );
  ANDN U1861 ( .B(n1854), .A(n1599), .Z(n1851) );
  XOR U1862 ( .A(n1855), .B(n1398), .Z(out[791]) );
  XOR U1863 ( .A(n1856), .B(n1857), .Z(n1398) );
  NOR U1864 ( .A(n1858), .B(n1601), .Z(n1855) );
  XOR U1865 ( .A(n1859), .B(n1402), .Z(out[790]) );
  XOR U1866 ( .A(n1860), .B(n1861), .Z(n1402) );
  NOR U1867 ( .A(n1862), .B(n1603), .Z(n1859) );
  XNOR U1868 ( .A(n1863), .B(n1864), .Z(out[78]) );
  AND U1869 ( .A(n1865), .B(n1866), .Z(n1863) );
  XOR U1870 ( .A(n1867), .B(n1406), .Z(out[789]) );
  XOR U1871 ( .A(n1868), .B(n1869), .Z(n1406) );
  NOR U1872 ( .A(n1870), .B(n1605), .Z(n1867) );
  XOR U1873 ( .A(n1871), .B(n1410), .Z(out[788]) );
  XOR U1874 ( .A(n1872), .B(n1873), .Z(n1410) );
  NOR U1875 ( .A(n1874), .B(n1607), .Z(n1871) );
  XOR U1876 ( .A(n1875), .B(n1414), .Z(out[787]) );
  XOR U1877 ( .A(n1876), .B(n1877), .Z(n1414) );
  NOR U1878 ( .A(n1878), .B(n1609), .Z(n1875) );
  XNOR U1879 ( .A(n1879), .B(n1418), .Z(out[786]) );
  XNOR U1880 ( .A(n1880), .B(n1881), .Z(n1418) );
  AND U1881 ( .A(n1882), .B(n1883), .Z(n1879) );
  XOR U1882 ( .A(n1884), .B(n1421), .Z(out[785]) );
  XNOR U1883 ( .A(n1885), .B(n1886), .Z(n1421) );
  AND U1884 ( .A(n1617), .B(n1887), .Z(n1884) );
  XOR U1885 ( .A(n1888), .B(n1425), .Z(out[784]) );
  XNOR U1886 ( .A(n1889), .B(n1890), .Z(n1425) );
  ANDN U1887 ( .B(n1891), .A(n1619), .Z(n1888) );
  XOR U1888 ( .A(n1892), .B(n1429), .Z(out[783]) );
  XOR U1889 ( .A(n1893), .B(n1894), .Z(n1429) );
  AND U1890 ( .A(n1621), .B(n1895), .Z(n1892) );
  XOR U1891 ( .A(n1896), .B(n1433), .Z(out[782]) );
  XOR U1892 ( .A(n1897), .B(n1898), .Z(n1433) );
  AND U1893 ( .A(n1623), .B(n1899), .Z(n1896) );
  XNOR U1894 ( .A(n1900), .B(n1442), .Z(out[781]) );
  XNOR U1895 ( .A(n1901), .B(n1902), .Z(n1442) );
  AND U1896 ( .A(n1903), .B(n1904), .Z(n1900) );
  XNOR U1897 ( .A(n1905), .B(n1446), .Z(out[780]) );
  XNOR U1898 ( .A(n1906), .B(n1907), .Z(n1446) );
  AND U1899 ( .A(n1627), .B(n1908), .Z(n1905) );
  XNOR U1900 ( .A(n1909), .B(n1910), .Z(out[77]) );
  XNOR U1901 ( .A(n1913), .B(n1450), .Z(out[779]) );
  XNOR U1902 ( .A(n1914), .B(n1915), .Z(n1450) );
  AND U1903 ( .A(n1916), .B(n1917), .Z(n1913) );
  XOR U1904 ( .A(n1918), .B(n1454), .Z(out[778]) );
  XOR U1905 ( .A(n1919), .B(n1920), .Z(n1454) );
  ANDN U1906 ( .B(n1921), .A(n1631), .Z(n1918) );
  XOR U1907 ( .A(n1922), .B(n1458), .Z(out[777]) );
  XOR U1908 ( .A(n1923), .B(n1924), .Z(n1458) );
  ANDN U1909 ( .B(n1925), .A(n1633), .Z(n1922) );
  XOR U1910 ( .A(n1926), .B(n1462), .Z(out[776]) );
  XOR U1911 ( .A(n1927), .B(n1928), .Z(n1462) );
  ANDN U1912 ( .B(n1929), .A(n1635), .Z(n1926) );
  XNOR U1913 ( .A(n1930), .B(n1466), .Z(out[775]) );
  XNOR U1914 ( .A(n1931), .B(n1932), .Z(n1466) );
  AND U1915 ( .A(n1933), .B(n1934), .Z(n1930) );
  XNOR U1916 ( .A(n1935), .B(n1470), .Z(out[774]) );
  XNOR U1917 ( .A(n1936), .B(n1937), .Z(n1470) );
  AND U1918 ( .A(n1938), .B(n1939), .Z(n1935) );
  XNOR U1919 ( .A(n1940), .B(n1474), .Z(out[773]) );
  XNOR U1920 ( .A(n1941), .B(n1942), .Z(n1474) );
  AND U1921 ( .A(n1943), .B(n1944), .Z(n1940) );
  XNOR U1922 ( .A(n1945), .B(n1478), .Z(out[772]) );
  XNOR U1923 ( .A(n1946), .B(n1947), .Z(n1478) );
  AND U1924 ( .A(n1948), .B(n1949), .Z(n1945) );
  XNOR U1925 ( .A(n1950), .B(n1490), .Z(out[771]) );
  XOR U1926 ( .A(n1951), .B(n1952), .Z(n1490) );
  AND U1927 ( .A(n1953), .B(n1954), .Z(n1950) );
  XNOR U1928 ( .A(n1955), .B(n1494), .Z(out[770]) );
  XOR U1929 ( .A(n1956), .B(n1957), .Z(n1494) );
  AND U1930 ( .A(n1958), .B(n1959), .Z(n1955) );
  XNOR U1931 ( .A(n1960), .B(n1961), .Z(out[76]) );
  ANDN U1932 ( .B(n1962), .A(n1963), .Z(n1960) );
  XNOR U1933 ( .A(n1964), .B(n1498), .Z(out[769]) );
  XOR U1934 ( .A(n1965), .B(n1966), .Z(n1498) );
  AND U1935 ( .A(n1967), .B(n1968), .Z(n1964) );
  XNOR U1936 ( .A(n1969), .B(n1502), .Z(out[768]) );
  XOR U1937 ( .A(n1970), .B(n1971), .Z(n1502) );
  AND U1938 ( .A(n1972), .B(n1973), .Z(n1969) );
  XOR U1939 ( .A(n1974), .B(n1504), .Z(out[767]) );
  IV U1940 ( .A(n1660), .Z(n1504) );
  XOR U1941 ( .A(n1975), .B(n1976), .Z(n1660) );
  NOR U1942 ( .A(n1224), .B(n1659), .Z(n1974) );
  XOR U1943 ( .A(n1977), .B(n1506), .Z(out[766]) );
  XOR U1944 ( .A(n1978), .B(n1979), .Z(n1506) );
  NOR U1945 ( .A(n1228), .B(n1664), .Z(n1977) );
  XOR U1946 ( .A(n1980), .B(n1508), .Z(out[765]) );
  XOR U1947 ( .A(n1981), .B(n1982), .Z(n1508) );
  NOR U1948 ( .A(n1672), .B(n1232), .Z(n1980) );
  XOR U1949 ( .A(n1983), .B(n1510), .Z(out[764]) );
  IV U1950 ( .A(n1677), .Z(n1510) );
  XNOR U1951 ( .A(n1984), .B(n1985), .Z(n1677) );
  NOR U1952 ( .A(n1676), .B(n1236), .Z(n1983) );
  XOR U1953 ( .A(n1986), .B(n1512), .Z(out[763]) );
  IV U1954 ( .A(n1682), .Z(n1512) );
  XNOR U1955 ( .A(n1987), .B(n1988), .Z(n1682) );
  XOR U1956 ( .A(n1990), .B(n1514), .Z(out[762]) );
  IV U1957 ( .A(n1687), .Z(n1514) );
  XNOR U1958 ( .A(n1991), .B(n1992), .Z(n1687) );
  NOR U1959 ( .A(n1686), .B(n1243), .Z(n1990) );
  XOR U1960 ( .A(n1993), .B(n1520), .Z(out[761]) );
  IV U1961 ( .A(n1692), .Z(n1520) );
  XNOR U1962 ( .A(n1994), .B(n1995), .Z(n1692) );
  NOR U1963 ( .A(n1691), .B(n1247), .Z(n1993) );
  XOR U1964 ( .A(n1996), .B(n1522), .Z(out[760]) );
  IV U1965 ( .A(n1697), .Z(n1522) );
  XNOR U1966 ( .A(n1997), .B(n1998), .Z(n1697) );
  NOR U1967 ( .A(n1696), .B(n1251), .Z(n1996) );
  XNOR U1968 ( .A(n1999), .B(n2000), .Z(out[75]) );
  XOR U1969 ( .A(n2003), .B(n1524), .Z(out[759]) );
  IV U1970 ( .A(n1702), .Z(n1524) );
  XNOR U1971 ( .A(n2004), .B(n2005), .Z(n1702) );
  XOR U1972 ( .A(n2007), .B(n1526), .Z(out[758]) );
  IV U1973 ( .A(n1707), .Z(n1526) );
  XNOR U1974 ( .A(n2008), .B(n2009), .Z(n1707) );
  IV U1975 ( .A(n2010), .Z(n1258) );
  XOR U1976 ( .A(n2011), .B(n1528), .Z(out[757]) );
  IV U1977 ( .A(n1712), .Z(n1528) );
  XNOR U1978 ( .A(n2012), .B(n2013), .Z(n1712) );
  XOR U1979 ( .A(n2015), .B(n1530), .Z(out[756]) );
  IV U1980 ( .A(n1717), .Z(n1530) );
  XNOR U1981 ( .A(n2016), .B(n2017), .Z(n1717) );
  XOR U1982 ( .A(n2019), .B(n1532), .Z(out[755]) );
  XOR U1983 ( .A(n2020), .B(n2021), .Z(n1532) );
  NOR U1984 ( .A(n1725), .B(n1272), .Z(n2019) );
  XOR U1985 ( .A(n2022), .B(n1534), .Z(out[754]) );
  XOR U1986 ( .A(n2023), .B(n2024), .Z(n1534) );
  IV U1987 ( .A(n2025), .Z(n1276) );
  XOR U1988 ( .A(n2026), .B(n1536), .Z(out[753]) );
  IV U1989 ( .A(n1734), .Z(n1536) );
  XOR U1990 ( .A(n2027), .B(n2028), .Z(n1734) );
  XOR U1991 ( .A(n2030), .B(n1538), .Z(out[752]) );
  IV U1992 ( .A(n1739), .Z(n1538) );
  XOR U1993 ( .A(n2031), .B(n2032), .Z(n1739) );
  XOR U1994 ( .A(n2034), .B(n1544), .Z(out[751]) );
  IV U1995 ( .A(n1744), .Z(n1544) );
  XOR U1996 ( .A(n2035), .B(n2036), .Z(n1744) );
  XOR U1997 ( .A(n2038), .B(n1546), .Z(out[750]) );
  IV U1998 ( .A(n1749), .Z(n1546) );
  XOR U1999 ( .A(n2039), .B(n2040), .Z(n1749) );
  XNOR U2000 ( .A(n2042), .B(n2043), .Z(out[74]) );
  XOR U2001 ( .A(n2046), .B(n1548), .Z(out[749]) );
  IV U2002 ( .A(n1754), .Z(n1548) );
  XOR U2003 ( .A(n2047), .B(n2048), .Z(n1754) );
  XOR U2004 ( .A(n2050), .B(n1550), .Z(out[748]) );
  IV U2005 ( .A(n1759), .Z(n1550) );
  XOR U2006 ( .A(n2051), .B(n2052), .Z(n1759) );
  XNOR U2007 ( .A(n2054), .B(n1552), .Z(out[747]) );
  XOR U2008 ( .A(n2055), .B(n2056), .Z(n1552) );
  ANDN U2009 ( .B(n2057), .A(n1307), .Z(n2054) );
  XOR U2010 ( .A(n2058), .B(n1554), .Z(out[746]) );
  IV U2011 ( .A(n1768), .Z(n1554) );
  XOR U2012 ( .A(n2059), .B(n2060), .Z(n1768) );
  NOR U2013 ( .A(n1311), .B(n1767), .Z(n2058) );
  XOR U2014 ( .A(n2061), .B(n1556), .Z(out[745]) );
  IV U2015 ( .A(n1777), .Z(n1556) );
  XOR U2016 ( .A(n2062), .B(n2063), .Z(n1777) );
  NOR U2017 ( .A(n1316), .B(n1776), .Z(n2061) );
  XNOR U2018 ( .A(n2064), .B(n1558), .Z(out[744]) );
  XOR U2019 ( .A(n2065), .B(n2066), .Z(n1558) );
  ANDN U2020 ( .B(n2067), .A(n1321), .Z(n2064) );
  XOR U2021 ( .A(n2068), .B(n1560), .Z(out[743]) );
  XOR U2022 ( .A(n2069), .B(n2070), .Z(n1560) );
  NOR U2023 ( .A(n1325), .B(n1785), .Z(n2068) );
  XOR U2024 ( .A(n2071), .B(n1563), .Z(out[742]) );
  XOR U2025 ( .A(n2072), .B(n2073), .Z(n1563) );
  NOR U2026 ( .A(n1329), .B(n1789), .Z(n2071) );
  XOR U2027 ( .A(n2074), .B(n1569), .Z(out[741]) );
  XOR U2028 ( .A(n2075), .B(n2076), .Z(n1569) );
  XNOR U2029 ( .A(n2078), .B(n1571), .Z(out[740]) );
  XNOR U2030 ( .A(n2079), .B(n2080), .Z(n1571) );
  ANDN U2031 ( .B(n2081), .A(n1336), .Z(n2078) );
  XNOR U2032 ( .A(n2082), .B(n2083), .Z(out[73]) );
  AND U2033 ( .A(n1042), .B(n2084), .Z(n2082) );
  XOR U2034 ( .A(n2085), .B(n1573), .Z(out[739]) );
  XOR U2035 ( .A(n2086), .B(n2087), .Z(n1573) );
  NOR U2036 ( .A(n1801), .B(n1340), .Z(n2085) );
  XNOR U2037 ( .A(n2088), .B(n1575), .Z(out[738]) );
  XOR U2038 ( .A(n2089), .B(n2090), .Z(n1575) );
  AND U2039 ( .A(n1344), .B(n2091), .Z(n2088) );
  XNOR U2040 ( .A(n2092), .B(n1577), .Z(out[737]) );
  XOR U2041 ( .A(n2093), .B(n2094), .Z(n1577) );
  AND U2042 ( .A(n1352), .B(n2095), .Z(n2092) );
  XNOR U2043 ( .A(n2096), .B(n1579), .Z(out[736]) );
  XOR U2044 ( .A(n2097), .B(n2098), .Z(n1579) );
  ANDN U2045 ( .B(n1813), .A(n1356), .Z(n2096) );
  XNOR U2046 ( .A(n2099), .B(n1581), .Z(out[735]) );
  XOR U2047 ( .A(n2100), .B(n2101), .Z(n1581) );
  ANDN U2048 ( .B(n2102), .A(n1360), .Z(n2099) );
  XNOR U2049 ( .A(n2103), .B(n1583), .Z(out[734]) );
  XOR U2050 ( .A(n2104), .B(n2105), .Z(n1583) );
  XNOR U2051 ( .A(n2106), .B(n1585), .Z(out[733]) );
  XOR U2052 ( .A(n2107), .B(n2108), .Z(n1585) );
  XNOR U2053 ( .A(n2109), .B(n1587), .Z(out[732]) );
  XOR U2054 ( .A(n2110), .B(n2111), .Z(n1587) );
  ANDN U2055 ( .B(n2112), .A(n1372), .Z(n2109) );
  XOR U2056 ( .A(n2113), .B(n1593), .Z(out[731]) );
  XOR U2057 ( .A(n2114), .B(n2115), .Z(n1593) );
  AND U2058 ( .A(n1841), .B(n1376), .Z(n2113) );
  IV U2059 ( .A(n2116), .Z(n1376) );
  XOR U2060 ( .A(n2117), .B(n1595), .Z(out[730]) );
  XNOR U2061 ( .A(n2118), .B(n2119), .Z(n1595) );
  AND U2062 ( .A(n1845), .B(n1380), .Z(n2117) );
  IV U2063 ( .A(n2120), .Z(n1380) );
  XNOR U2064 ( .A(n2121), .B(n2122), .Z(out[72]) );
  AND U2065 ( .A(n1482), .B(n1480), .Z(n2121) );
  XOR U2066 ( .A(n2123), .B(n1597), .Z(out[729]) );
  IV U2067 ( .A(n1850), .Z(n1597) );
  XNOR U2068 ( .A(n2124), .B(n2125), .Z(n1850) );
  NOR U2069 ( .A(n1849), .B(n1384), .Z(n2123) );
  XOR U2070 ( .A(n2126), .B(n1599), .Z(out[728]) );
  XOR U2071 ( .A(n2127), .B(n2128), .Z(n1599) );
  ANDN U2072 ( .B(n2129), .A(n1388), .Z(n2126) );
  XOR U2073 ( .A(n2130), .B(n1601), .Z(out[727]) );
  XOR U2074 ( .A(n2131), .B(n2132), .Z(n1601) );
  AND U2075 ( .A(n1858), .B(n1396), .Z(n2130) );
  IV U2076 ( .A(n2133), .Z(n1396) );
  XOR U2077 ( .A(n2134), .B(n1603), .Z(out[726]) );
  XOR U2078 ( .A(n2135), .B(n2136), .Z(n1603) );
  AND U2079 ( .A(n1862), .B(n1400), .Z(n2134) );
  IV U2080 ( .A(n2137), .Z(n1400) );
  XOR U2081 ( .A(n2138), .B(n1605), .Z(out[725]) );
  XOR U2082 ( .A(n2139), .B(n2140), .Z(n1605) );
  AND U2083 ( .A(n1870), .B(n1404), .Z(n2138) );
  IV U2084 ( .A(n2141), .Z(n1404) );
  XOR U2085 ( .A(n2142), .B(n1607), .Z(out[724]) );
  XOR U2086 ( .A(n2143), .B(n2144), .Z(n1607) );
  AND U2087 ( .A(n1874), .B(n1408), .Z(n2142) );
  IV U2088 ( .A(n2145), .Z(n1408) );
  XOR U2089 ( .A(n2146), .B(n1609), .Z(out[723]) );
  XNOR U2090 ( .A(n2147), .B(n2148), .Z(n1609) );
  AND U2091 ( .A(n1878), .B(n1412), .Z(n2146) );
  IV U2092 ( .A(n2149), .Z(n1412) );
  XOR U2093 ( .A(n2150), .B(n1611), .Z(out[722]) );
  IV U2094 ( .A(n1883), .Z(n1611) );
  XOR U2095 ( .A(n2151), .B(n2152), .Z(n1883) );
  NOR U2096 ( .A(n1882), .B(n1416), .Z(n2150) );
  XNOR U2097 ( .A(n2153), .B(n1617), .Z(out[721]) );
  XNOR U2098 ( .A(n2154), .B(n2155), .Z(n1617) );
  ANDN U2099 ( .B(n2156), .A(n1420), .Z(n2153) );
  XOR U2100 ( .A(n2157), .B(n1619), .Z(out[720]) );
  XOR U2101 ( .A(n2158), .B(n2159), .Z(n1619) );
  NOR U2102 ( .A(n1891), .B(n1424), .Z(n2157) );
  XNOR U2103 ( .A(n2160), .B(n2161), .Z(out[71]) );
  AND U2104 ( .A(n1817), .B(n1815), .Z(n2160) );
  XNOR U2105 ( .A(n2162), .B(n1621), .Z(out[719]) );
  XNOR U2106 ( .A(n2163), .B(n2164), .Z(n1621) );
  ANDN U2107 ( .B(n2165), .A(n1428), .Z(n2162) );
  XNOR U2108 ( .A(n2166), .B(n1623), .Z(out[718]) );
  XNOR U2109 ( .A(n2167), .B(n2168), .Z(n1623) );
  ANDN U2110 ( .B(n2169), .A(n1432), .Z(n2166) );
  XOR U2111 ( .A(n2170), .B(n1625), .Z(out[717]) );
  IV U2112 ( .A(n1904), .Z(n1625) );
  XNOR U2113 ( .A(n2171), .B(n2172), .Z(n1904) );
  NOR U2114 ( .A(n1440), .B(n1903), .Z(n2170) );
  XNOR U2115 ( .A(n2173), .B(n1627), .Z(out[716]) );
  XOR U2116 ( .A(n2174), .B(n2175), .Z(n1627) );
  NOR U2117 ( .A(n1444), .B(n1908), .Z(n2173) );
  XOR U2118 ( .A(n2176), .B(n1629), .Z(out[715]) );
  IV U2119 ( .A(n1917), .Z(n1629) );
  XNOR U2120 ( .A(n2177), .B(n2178), .Z(n1917) );
  NOR U2121 ( .A(n1448), .B(n1916), .Z(n2176) );
  XOR U2122 ( .A(n2179), .B(n1631), .Z(out[714]) );
  XNOR U2123 ( .A(n2180), .B(n2181), .Z(n1631) );
  NOR U2124 ( .A(n1452), .B(n1921), .Z(n2179) );
  XOR U2125 ( .A(n2182), .B(n1633), .Z(out[713]) );
  XNOR U2126 ( .A(n2183), .B(n2184), .Z(n1633) );
  ANDN U2127 ( .B(n2185), .A(n1456), .Z(n2182) );
  XOR U2128 ( .A(n2186), .B(n1635), .Z(out[712]) );
  XNOR U2129 ( .A(n2187), .B(n2188), .Z(n1635) );
  NOR U2130 ( .A(n1929), .B(n1460), .Z(n2186) );
  XOR U2131 ( .A(n2189), .B(n1641), .Z(out[711]) );
  IV U2132 ( .A(n1934), .Z(n1641) );
  XNOR U2133 ( .A(n2190), .B(n2191), .Z(n1934) );
  NOR U2134 ( .A(n1933), .B(n1464), .Z(n2189) );
  XOR U2135 ( .A(n2192), .B(n1643), .Z(out[710]) );
  IV U2136 ( .A(n1939), .Z(n1643) );
  XOR U2137 ( .A(n2193), .B(n2194), .Z(n1939) );
  NOR U2138 ( .A(n1938), .B(n1468), .Z(n2192) );
  XNOR U2139 ( .A(n2195), .B(n2196), .Z(out[70]) );
  AND U2140 ( .A(n2197), .B(n2198), .Z(n2195) );
  XOR U2141 ( .A(n2199), .B(n1645), .Z(out[709]) );
  IV U2142 ( .A(n1944), .Z(n1645) );
  XOR U2143 ( .A(n2200), .B(n2201), .Z(n1944) );
  NOR U2144 ( .A(n1943), .B(n1472), .Z(n2199) );
  XOR U2145 ( .A(n2202), .B(n1647), .Z(out[708]) );
  IV U2146 ( .A(n1949), .Z(n1647) );
  XOR U2147 ( .A(n2203), .B(n2204), .Z(n1949) );
  NOR U2148 ( .A(n1948), .B(n1476), .Z(n2202) );
  XOR U2149 ( .A(n2205), .B(n1649), .Z(out[707]) );
  IV U2150 ( .A(n1954), .Z(n1649) );
  XNOR U2151 ( .A(n2206), .B(n2207), .Z(n1954) );
  NOR U2152 ( .A(n1953), .B(n1488), .Z(n2205) );
  XOR U2153 ( .A(n2208), .B(n1651), .Z(out[706]) );
  IV U2154 ( .A(n1959), .Z(n1651) );
  XOR U2155 ( .A(n2209), .B(n2210), .Z(n1959) );
  NOR U2156 ( .A(n1958), .B(n1492), .Z(n2208) );
  XOR U2157 ( .A(n2211), .B(n1653), .Z(out[705]) );
  IV U2158 ( .A(n1968), .Z(n1653) );
  XOR U2159 ( .A(n2212), .B(n2213), .Z(n1968) );
  NOR U2160 ( .A(n1967), .B(n1496), .Z(n2211) );
  XOR U2161 ( .A(n2214), .B(n1655), .Z(out[704]) );
  IV U2162 ( .A(n1973), .Z(n1655) );
  XOR U2163 ( .A(n2215), .B(n2216), .Z(n1973) );
  NOR U2164 ( .A(n1972), .B(n1500), .Z(n2214) );
  XOR U2165 ( .A(n2217), .B(n1659), .Z(out[703]) );
  XNOR U2166 ( .A(n2218), .B(n2219), .Z(n1659) );
  ANDN U2167 ( .B(n1224), .A(n1225), .Z(n2217) );
  XOR U2168 ( .A(n2220), .B(n2221), .Z(n1225) );
  XNOR U2169 ( .A(n2222), .B(n2223), .Z(n1224) );
  XOR U2170 ( .A(n2224), .B(n1664), .Z(out[702]) );
  XNOR U2171 ( .A(n2225), .B(n2226), .Z(n1664) );
  ANDN U2172 ( .B(n1228), .A(n1229), .Z(n2224) );
  XOR U2173 ( .A(n2227), .B(n2228), .Z(n1229) );
  XNOR U2174 ( .A(n2229), .B(n2230), .Z(n1228) );
  XOR U2175 ( .A(n2231), .B(n1672), .Z(out[701]) );
  XNOR U2176 ( .A(n2232), .B(n2233), .Z(n1672) );
  ANDN U2177 ( .B(n1232), .A(n1233), .Z(n2231) );
  XOR U2178 ( .A(n2234), .B(n2235), .Z(n1233) );
  XNOR U2179 ( .A(n2236), .B(n2237), .Z(n1232) );
  XOR U2180 ( .A(n2238), .B(n1676), .Z(out[700]) );
  XNOR U2181 ( .A(n2239), .B(n2240), .Z(n1676) );
  ANDN U2182 ( .B(n1236), .A(n1237), .Z(n2238) );
  XNOR U2183 ( .A(n2241), .B(n2242), .Z(n1237) );
  XNOR U2184 ( .A(n2243), .B(n2244), .Z(n1236) );
  XNOR U2185 ( .A(n2245), .B(n2197), .Z(out[6]) );
  AND U2186 ( .A(n2246), .B(n2247), .Z(n2245) );
  XOR U2187 ( .A(n2248), .B(n2249), .Z(out[69]) );
  ANDN U2188 ( .B(n2250), .A(n2251), .Z(n2248) );
  XOR U2189 ( .A(n2252), .B(n1681), .Z(out[699]) );
  XOR U2190 ( .A(n2253), .B(n2254), .Z(n1681) );
  ANDN U2191 ( .B(n1989), .A(n1240), .Z(n2252) );
  XNOR U2192 ( .A(n2255), .B(n2256), .Z(n1240) );
  XNOR U2193 ( .A(n2257), .B(n2258), .Z(n1989) );
  XOR U2194 ( .A(n2259), .B(n1686), .Z(out[698]) );
  XOR U2195 ( .A(n2260), .B(n2261), .Z(n1686) );
  ANDN U2196 ( .B(n1243), .A(n1244), .Z(n2259) );
  XNOR U2197 ( .A(n2262), .B(n2263), .Z(n1244) );
  XNOR U2198 ( .A(n2264), .B(n2265), .Z(n1243) );
  XOR U2199 ( .A(n2266), .B(n1691), .Z(out[697]) );
  XOR U2200 ( .A(n2267), .B(n2268), .Z(n1691) );
  ANDN U2201 ( .B(n1247), .A(n1248), .Z(n2266) );
  XNOR U2202 ( .A(n2269), .B(n2270), .Z(n1248) );
  XNOR U2203 ( .A(n2271), .B(n2272), .Z(n1247) );
  XOR U2204 ( .A(n2273), .B(n1696), .Z(out[696]) );
  XOR U2205 ( .A(n2274), .B(n2275), .Z(n1696) );
  ANDN U2206 ( .B(n1251), .A(n1252), .Z(n2273) );
  XNOR U2207 ( .A(n2276), .B(n2277), .Z(n1252) );
  XNOR U2208 ( .A(n2278), .B(n2279), .Z(n1251) );
  XOR U2209 ( .A(n2280), .B(n1701), .Z(out[695]) );
  XOR U2210 ( .A(n2281), .B(n2282), .Z(n1701) );
  ANDN U2211 ( .B(n2006), .A(n1255), .Z(n2280) );
  XNOR U2212 ( .A(n2283), .B(n2284), .Z(n1255) );
  XOR U2213 ( .A(n2285), .B(n2286), .Z(n2006) );
  XOR U2214 ( .A(n2287), .B(n1706), .Z(out[694]) );
  XOR U2215 ( .A(n2288), .B(n2289), .Z(n1706) );
  ANDN U2216 ( .B(n2010), .A(n1259), .Z(n2287) );
  XNOR U2217 ( .A(n2290), .B(n2291), .Z(n1259) );
  XOR U2218 ( .A(n2292), .B(n2293), .Z(n2010) );
  XOR U2219 ( .A(n2294), .B(n1711), .Z(out[693]) );
  XOR U2220 ( .A(n2295), .B(n2296), .Z(n1711) );
  ANDN U2221 ( .B(n2014), .A(n1266), .Z(n2294) );
  XNOR U2222 ( .A(n2297), .B(n2298), .Z(n1266) );
  XOR U2223 ( .A(n2299), .B(n2300), .Z(n2014) );
  XOR U2224 ( .A(n2301), .B(n1716), .Z(out[692]) );
  XOR U2225 ( .A(n2302), .B(n2303), .Z(n1716) );
  ANDN U2226 ( .B(n2018), .A(n1269), .Z(n2301) );
  XNOR U2227 ( .A(n2304), .B(n2305), .Z(n1269) );
  XOR U2228 ( .A(n2306), .B(n2307), .Z(n2018) );
  XOR U2229 ( .A(n2308), .B(n1725), .Z(out[691]) );
  XNOR U2230 ( .A(n2309), .B(n2310), .Z(n1725) );
  ANDN U2231 ( .B(n1272), .A(n1273), .Z(n2308) );
  XNOR U2232 ( .A(n2311), .B(n2312), .Z(n1273) );
  XOR U2233 ( .A(n2313), .B(n2314), .Z(n1272) );
  XOR U2234 ( .A(n2315), .B(n1729), .Z(out[690]) );
  XOR U2235 ( .A(n2316), .B(n2317), .Z(n1729) );
  ANDN U2236 ( .B(n2025), .A(n1277), .Z(n2315) );
  XNOR U2237 ( .A(n2318), .B(n2319), .Z(n1277) );
  XOR U2238 ( .A(n2320), .B(n2321), .Z(n2025) );
  XNOR U2239 ( .A(n2322), .B(n2323), .Z(out[68]) );
  AND U2240 ( .A(n2324), .B(n2325), .Z(n2322) );
  XOR U2241 ( .A(n2326), .B(n1733), .Z(out[689]) );
  XOR U2242 ( .A(n2327), .B(n2328), .Z(n1733) );
  ANDN U2243 ( .B(n2029), .A(n1280), .Z(n2326) );
  XNOR U2244 ( .A(n2329), .B(n2330), .Z(n1280) );
  XOR U2245 ( .A(n2331), .B(n2332), .Z(n2029) );
  XOR U2246 ( .A(n2333), .B(n1738), .Z(out[688]) );
  XOR U2247 ( .A(n2334), .B(n2335), .Z(n1738) );
  AND U2248 ( .A(n1285), .B(n2033), .Z(n2333) );
  XOR U2249 ( .A(n2336), .B(n2337), .Z(n2033) );
  XOR U2250 ( .A(n2338), .B(n2339), .Z(n1285) );
  XOR U2251 ( .A(n2340), .B(n1743), .Z(out[687]) );
  XOR U2252 ( .A(n2341), .B(n2342), .Z(n1743) );
  AND U2253 ( .A(n1289), .B(n2037), .Z(n2340) );
  XOR U2254 ( .A(n2343), .B(n2344), .Z(n2037) );
  XOR U2255 ( .A(n2345), .B(n2346), .Z(n1289) );
  XOR U2256 ( .A(n2347), .B(n1748), .Z(out[686]) );
  XOR U2257 ( .A(n2348), .B(n2349), .Z(n1748) );
  AND U2258 ( .A(n1293), .B(n2041), .Z(n2347) );
  XOR U2259 ( .A(n2350), .B(n2351), .Z(n2041) );
  XOR U2260 ( .A(n2352), .B(n2353), .Z(n1293) );
  XOR U2261 ( .A(n2354), .B(n1753), .Z(out[685]) );
  XOR U2262 ( .A(n2355), .B(n2356), .Z(n1753) );
  AND U2263 ( .A(n1297), .B(n2049), .Z(n2354) );
  XOR U2264 ( .A(n2357), .B(n2358), .Z(n2049) );
  XOR U2265 ( .A(n2359), .B(n2360), .Z(n1297) );
  XOR U2266 ( .A(n2361), .B(n1758), .Z(out[684]) );
  XOR U2267 ( .A(n2362), .B(n2363), .Z(n1758) );
  AND U2268 ( .A(n1301), .B(n2053), .Z(n2361) );
  XOR U2269 ( .A(n2364), .B(n2365), .Z(n2053) );
  XOR U2270 ( .A(n2366), .B(n2367), .Z(n1301) );
  XOR U2271 ( .A(n2368), .B(n1763), .Z(out[683]) );
  IV U2272 ( .A(n2057), .Z(n1763) );
  XOR U2273 ( .A(n2369), .B(n2370), .Z(n2057) );
  AND U2274 ( .A(n1307), .B(n1309), .Z(n2368) );
  XOR U2275 ( .A(n2371), .B(n2372), .Z(n1309) );
  XNOR U2276 ( .A(n2373), .B(n2374), .Z(n1307) );
  XOR U2277 ( .A(n2375), .B(n1767), .Z(out[682]) );
  XNOR U2278 ( .A(n2376), .B(n2377), .Z(n1767) );
  AND U2279 ( .A(n1314), .B(n1311), .Z(n2375) );
  XNOR U2280 ( .A(n2378), .B(n2379), .Z(n1311) );
  XOR U2281 ( .A(n2380), .B(n2381), .Z(n1314) );
  XOR U2282 ( .A(n2382), .B(n1776), .Z(out[681]) );
  XNOR U2283 ( .A(n2383), .B(n2384), .Z(n1776) );
  AND U2284 ( .A(n1319), .B(n1316), .Z(n2382) );
  XNOR U2285 ( .A(n2385), .B(n2386), .Z(n1316) );
  XOR U2286 ( .A(n2387), .B(n2388), .Z(n1319) );
  XOR U2287 ( .A(n2389), .B(n1781), .Z(out[680]) );
  IV U2288 ( .A(n2067), .Z(n1781) );
  XOR U2289 ( .A(n2390), .B(n2391), .Z(n2067) );
  AND U2290 ( .A(n1321), .B(n1323), .Z(n2389) );
  XOR U2291 ( .A(n2392), .B(n2393), .Z(n1323) );
  XNOR U2292 ( .A(n2394), .B(n2395), .Z(n1321) );
  XOR U2293 ( .A(n2396), .B(n2397), .Z(out[67]) );
  ANDN U2294 ( .B(n2398), .A(n2399), .Z(n2396) );
  XOR U2295 ( .A(n2400), .B(n1785), .Z(out[679]) );
  XNOR U2296 ( .A(n2401), .B(n2402), .Z(n1785) );
  AND U2297 ( .A(n1327), .B(n1325), .Z(n2400) );
  XNOR U2298 ( .A(n2403), .B(n2404), .Z(n1325) );
  XNOR U2299 ( .A(n2405), .B(n2406), .Z(n1327) );
  XOR U2300 ( .A(n2407), .B(n1789), .Z(out[678]) );
  XNOR U2301 ( .A(n2408), .B(n2409), .Z(n1789) );
  ANDN U2302 ( .B(n1329), .A(n1330), .Z(n2407) );
  XNOR U2303 ( .A(n2410), .B(n2411), .Z(n1330) );
  XNOR U2304 ( .A(n2412), .B(n2413), .Z(n1329) );
  XOR U2305 ( .A(n2414), .B(n1793), .Z(out[677]) );
  XOR U2306 ( .A(n2415), .B(n2416), .Z(n1793) );
  ANDN U2307 ( .B(n2077), .A(n1333), .Z(n2414) );
  XNOR U2308 ( .A(n2417), .B(n2418), .Z(n1333) );
  XNOR U2309 ( .A(n2419), .B(n2420), .Z(n2077) );
  XOR U2310 ( .A(n2421), .B(n1797), .Z(out[676]) );
  IV U2311 ( .A(n2081), .Z(n1797) );
  XOR U2312 ( .A(n2422), .B(n2423), .Z(n2081) );
  AND U2313 ( .A(n1336), .B(n1338), .Z(n2421) );
  XOR U2314 ( .A(n2424), .B(n2425), .Z(n1338) );
  XNOR U2315 ( .A(n2426), .B(n2427), .Z(n1336) );
  XOR U2316 ( .A(n2428), .B(n1801), .Z(out[675]) );
  XNOR U2317 ( .A(n2429), .B(n2430), .Z(n1801) );
  AND U2318 ( .A(n1340), .B(n1342), .Z(n2428) );
  XOR U2319 ( .A(n2431), .B(n2432), .Z(n1342) );
  XNOR U2320 ( .A(n2433), .B(n2434), .Z(n1340) );
  XOR U2321 ( .A(n2435), .B(n1805), .Z(out[674]) );
  IV U2322 ( .A(n2091), .Z(n1805) );
  XOR U2323 ( .A(n2436), .B(n2437), .Z(n2091) );
  ANDN U2324 ( .B(n1346), .A(n1344), .Z(n2435) );
  XOR U2325 ( .A(n2438), .B(n2439), .Z(n1344) );
  XOR U2326 ( .A(n2440), .B(n2441), .Z(n1346) );
  XOR U2327 ( .A(n2442), .B(n1809), .Z(out[673]) );
  IV U2328 ( .A(n2095), .Z(n1809) );
  XOR U2329 ( .A(n2443), .B(n2444), .Z(n2095) );
  ANDN U2330 ( .B(n1354), .A(n1352), .Z(n2442) );
  XOR U2331 ( .A(n2445), .B(n2446), .Z(n1352) );
  XOR U2332 ( .A(n2447), .B(n2448), .Z(n1354) );
  XNOR U2333 ( .A(n2449), .B(n1813), .Z(out[672]) );
  XOR U2334 ( .A(n2450), .B(n2451), .Z(n1813) );
  AND U2335 ( .A(n1356), .B(n1358), .Z(n2449) );
  XOR U2336 ( .A(n2452), .B(n2453), .Z(n1358) );
  XNOR U2337 ( .A(n2454), .B(n2455), .Z(n1356) );
  XOR U2338 ( .A(n2456), .B(n1825), .Z(out[671]) );
  IV U2339 ( .A(n2102), .Z(n1825) );
  XOR U2340 ( .A(n2457), .B(n2458), .Z(n2102) );
  AND U2341 ( .A(n1360), .B(n1362), .Z(n2456) );
  XOR U2342 ( .A(n2459), .B(n2460), .Z(n1362) );
  XOR U2343 ( .A(n2461), .B(n2462), .Z(n1360) );
  XOR U2344 ( .A(n2463), .B(n1829), .Z(out[670]) );
  XOR U2345 ( .A(n2464), .B(n2465), .Z(n1829) );
  AND U2346 ( .A(n1364), .B(n1366), .Z(n2463) );
  XOR U2347 ( .A(n2466), .B(n2467), .Z(n1366) );
  XOR U2348 ( .A(n2468), .B(n2469), .Z(n1364) );
  XOR U2349 ( .A(n2470), .B(n2471), .Z(out[66]) );
  ANDN U2350 ( .B(n2472), .A(n2473), .Z(n2470) );
  XOR U2351 ( .A(n2474), .B(n1833), .Z(out[669]) );
  XOR U2352 ( .A(n2475), .B(n2476), .Z(n1833) );
  AND U2353 ( .A(n1368), .B(n1370), .Z(n2474) );
  XOR U2354 ( .A(n2477), .B(n2478), .Z(n1370) );
  XOR U2355 ( .A(n2479), .B(n2480), .Z(n1368) );
  XOR U2356 ( .A(n2481), .B(n1837), .Z(out[668]) );
  IV U2357 ( .A(n2112), .Z(n1837) );
  XNOR U2358 ( .A(n2482), .B(n2483), .Z(n2112) );
  AND U2359 ( .A(n1372), .B(n1374), .Z(n2481) );
  XOR U2360 ( .A(n2484), .B(n2485), .Z(n1374) );
  XNOR U2361 ( .A(n2486), .B(n2487), .Z(n1372) );
  XNOR U2362 ( .A(n2488), .B(n1841), .Z(out[667]) );
  XOR U2363 ( .A(n2489), .B(n2490), .Z(n1841) );
  AND U2364 ( .A(n1378), .B(n2116), .Z(n2488) );
  XNOR U2365 ( .A(n2491), .B(n2492), .Z(n2116) );
  XOR U2366 ( .A(n2493), .B(n2494), .Z(n1378) );
  XNOR U2367 ( .A(n2495), .B(n1845), .Z(out[666]) );
  XOR U2368 ( .A(n2496), .B(n2497), .Z(n1845) );
  AND U2369 ( .A(n1382), .B(n2120), .Z(n2495) );
  XNOR U2370 ( .A(n2498), .B(n2499), .Z(n2120) );
  XOR U2371 ( .A(n2500), .B(n2501), .Z(n1382) );
  XOR U2372 ( .A(n2502), .B(n1849), .Z(out[665]) );
  XOR U2373 ( .A(n2503), .B(n2504), .Z(n1849) );
  AND U2374 ( .A(n1384), .B(n1386), .Z(n2502) );
  XOR U2375 ( .A(n2505), .B(n2506), .Z(n1386) );
  XNOR U2376 ( .A(n2507), .B(n2508), .Z(n1384) );
  XOR U2377 ( .A(n2509), .B(n1854), .Z(out[664]) );
  IV U2378 ( .A(n2129), .Z(n1854) );
  XOR U2379 ( .A(n2510), .B(n2511), .Z(n2129) );
  ANDN U2380 ( .B(n1388), .A(n1389), .Z(n2509) );
  XNOR U2381 ( .A(n2512), .B(n2513), .Z(n1389) );
  XNOR U2382 ( .A(n2514), .B(n2515), .Z(n1388) );
  XNOR U2383 ( .A(n2516), .B(n1858), .Z(out[663]) );
  XOR U2384 ( .A(n2517), .B(n2518), .Z(n1858) );
  ANDN U2385 ( .B(n2133), .A(n1397), .Z(n2516) );
  XOR U2386 ( .A(n2519), .B(n2520), .Z(n1397) );
  XNOR U2387 ( .A(n2521), .B(n2522), .Z(n2133) );
  XNOR U2388 ( .A(n2523), .B(n1862), .Z(out[662]) );
  XOR U2389 ( .A(n2524), .B(n2525), .Z(n1862) );
  ANDN U2390 ( .B(n2137), .A(n1401), .Z(n2523) );
  XOR U2391 ( .A(n2526), .B(n2527), .Z(n1401) );
  XNOR U2392 ( .A(n2528), .B(n2529), .Z(n2137) );
  XNOR U2393 ( .A(n2530), .B(n1870), .Z(out[661]) );
  XOR U2394 ( .A(n2531), .B(n2532), .Z(n1870) );
  ANDN U2395 ( .B(n2141), .A(n1405), .Z(n2530) );
  XOR U2396 ( .A(n2533), .B(n2534), .Z(n1405) );
  XNOR U2397 ( .A(n2535), .B(n2536), .Z(n2141) );
  XNOR U2398 ( .A(n2537), .B(n1874), .Z(out[660]) );
  XOR U2399 ( .A(n2538), .B(n2539), .Z(n1874) );
  ANDN U2400 ( .B(n2145), .A(n1409), .Z(n2537) );
  XOR U2401 ( .A(n2540), .B(n2541), .Z(n1409) );
  XNOR U2402 ( .A(n2542), .B(n2543), .Z(n2145) );
  XOR U2403 ( .A(n2544), .B(n2545), .Z(out[65]) );
  ANDN U2404 ( .B(n2546), .A(n2547), .Z(n2544) );
  XNOR U2405 ( .A(n2548), .B(n1878), .Z(out[659]) );
  XOR U2406 ( .A(n2549), .B(n2550), .Z(n1878) );
  ANDN U2407 ( .B(n2149), .A(n1413), .Z(n2548) );
  XOR U2408 ( .A(n2551), .B(n2552), .Z(n1413) );
  XOR U2409 ( .A(n2553), .B(n2554), .Z(n2149) );
  XOR U2410 ( .A(n2555), .B(n1882), .Z(out[658]) );
  XNOR U2411 ( .A(n2556), .B(n2557), .Z(n1882) );
  ANDN U2412 ( .B(n1416), .A(n1417), .Z(n2555) );
  XOR U2413 ( .A(n2558), .B(n2559), .Z(n1417) );
  XNOR U2414 ( .A(n2560), .B(n2561), .Z(n1416) );
  XOR U2415 ( .A(n2562), .B(n1887), .Z(out[657]) );
  IV U2416 ( .A(n2156), .Z(n1887) );
  XOR U2417 ( .A(n2563), .B(n2564), .Z(n2156) );
  AND U2418 ( .A(n1420), .B(n1422), .Z(n2562) );
  XOR U2419 ( .A(n2565), .B(n2566), .Z(n1422) );
  XOR U2420 ( .A(n2567), .B(n2568), .Z(n1420) );
  XOR U2421 ( .A(n2569), .B(n1891), .Z(out[656]) );
  XOR U2422 ( .A(n2570), .B(n2571), .Z(n1891) );
  ANDN U2423 ( .B(n1424), .A(n1426), .Z(n2569) );
  XNOR U2424 ( .A(n2572), .B(n2573), .Z(n1426) );
  XNOR U2425 ( .A(n2574), .B(n2575), .Z(n1424) );
  XOR U2426 ( .A(n2576), .B(n1895), .Z(out[655]) );
  IV U2427 ( .A(n2165), .Z(n1895) );
  XOR U2428 ( .A(n2577), .B(n2578), .Z(n2165) );
  ANDN U2429 ( .B(n1428), .A(n1430), .Z(n2576) );
  XNOR U2430 ( .A(n2579), .B(n2580), .Z(n1430) );
  XOR U2431 ( .A(n2581), .B(n2582), .Z(n1428) );
  XOR U2432 ( .A(n2583), .B(n1899), .Z(out[654]) );
  IV U2433 ( .A(n2169), .Z(n1899) );
  XOR U2434 ( .A(n2584), .B(n2585), .Z(n2169) );
  ANDN U2435 ( .B(n1432), .A(n1434), .Z(n2583) );
  XNOR U2436 ( .A(n2586), .B(n2587), .Z(n1434) );
  XOR U2437 ( .A(n2588), .B(n2589), .Z(n1432) );
  XOR U2438 ( .A(n2590), .B(n1903), .Z(out[653]) );
  XNOR U2439 ( .A(n2591), .B(n2592), .Z(n1903) );
  ANDN U2440 ( .B(n1440), .A(n1441), .Z(n2590) );
  XNOR U2441 ( .A(n2593), .B(n2594), .Z(n1441) );
  XOR U2442 ( .A(n2595), .B(n2596), .Z(n1440) );
  XOR U2443 ( .A(n2597), .B(n1908), .Z(out[652]) );
  XOR U2444 ( .A(n2598), .B(n2599), .Z(n1908) );
  ANDN U2445 ( .B(n1444), .A(n1445), .Z(n2597) );
  XNOR U2446 ( .A(n2600), .B(n2601), .Z(n1445) );
  XNOR U2447 ( .A(n2602), .B(n2603), .Z(n1444) );
  XOR U2448 ( .A(n2604), .B(n1916), .Z(out[651]) );
  XOR U2449 ( .A(n2605), .B(n2606), .Z(n1916) );
  ANDN U2450 ( .B(n1448), .A(n1449), .Z(n2604) );
  XNOR U2451 ( .A(n2607), .B(n2608), .Z(n1449) );
  XNOR U2452 ( .A(n2609), .B(n2610), .Z(n1448) );
  XOR U2453 ( .A(n2611), .B(n1921), .Z(out[650]) );
  XOR U2454 ( .A(n2612), .B(n2613), .Z(n1921) );
  ANDN U2455 ( .B(n1452), .A(n1453), .Z(n2611) );
  XNOR U2456 ( .A(n2614), .B(n2615), .Z(n1453) );
  XNOR U2457 ( .A(n2616), .B(n2617), .Z(n1452) );
  AND U2458 ( .A(n2620), .B(n2621), .Z(n2618) );
  IV U2459 ( .A(n2622), .Z(n2621) );
  XOR U2460 ( .A(n2623), .B(n1925), .Z(out[649]) );
  IV U2461 ( .A(n2185), .Z(n1925) );
  XOR U2462 ( .A(n2624), .B(n2625), .Z(n2185) );
  ANDN U2463 ( .B(n1456), .A(n1457), .Z(n2623) );
  XNOR U2464 ( .A(n2626), .B(n2627), .Z(n1457) );
  XNOR U2465 ( .A(n2628), .B(n2629), .Z(n1456) );
  XOR U2466 ( .A(n2630), .B(n1929), .Z(out[648]) );
  XOR U2467 ( .A(n2631), .B(n2632), .Z(n1929) );
  ANDN U2468 ( .B(n1460), .A(n1461), .Z(n2630) );
  XNOR U2469 ( .A(n2633), .B(n2634), .Z(n1461) );
  XNOR U2470 ( .A(n2635), .B(n2636), .Z(n1460) );
  XOR U2471 ( .A(n2637), .B(n1933), .Z(out[647]) );
  XNOR U2472 ( .A(n2638), .B(n2639), .Z(n1933) );
  ANDN U2473 ( .B(n1464), .A(n1465), .Z(n2637) );
  XNOR U2474 ( .A(n2640), .B(n2641), .Z(n1465) );
  XNOR U2475 ( .A(n2642), .B(n2643), .Z(n1464) );
  XOR U2476 ( .A(n2644), .B(n1938), .Z(out[646]) );
  XNOR U2477 ( .A(n2645), .B(n2646), .Z(n1938) );
  ANDN U2478 ( .B(n1468), .A(n1469), .Z(n2644) );
  XNOR U2479 ( .A(n2647), .B(n2648), .Z(n1469) );
  XNOR U2480 ( .A(n2649), .B(n2650), .Z(n1468) );
  XOR U2481 ( .A(n2651), .B(n1943), .Z(out[645]) );
  XNOR U2482 ( .A(n2652), .B(n2653), .Z(n1943) );
  ANDN U2483 ( .B(n1472), .A(n1473), .Z(n2651) );
  XNOR U2484 ( .A(n2654), .B(n2655), .Z(n1473) );
  XNOR U2485 ( .A(n2656), .B(n2657), .Z(n1472) );
  XOR U2486 ( .A(n2658), .B(n1948), .Z(out[644]) );
  XNOR U2487 ( .A(n2659), .B(n2660), .Z(n1948) );
  ANDN U2488 ( .B(n1476), .A(n1477), .Z(n2658) );
  XNOR U2489 ( .A(n2661), .B(n2662), .Z(n1477) );
  XNOR U2490 ( .A(n2663), .B(n2664), .Z(n1476) );
  XOR U2491 ( .A(n2665), .B(n1953), .Z(out[643]) );
  XNOR U2492 ( .A(n2666), .B(n2667), .Z(n1953) );
  ANDN U2493 ( .B(n1488), .A(n1489), .Z(n2665) );
  XNOR U2494 ( .A(n2668), .B(n2669), .Z(n1489) );
  XNOR U2495 ( .A(n2670), .B(n2671), .Z(n1488) );
  XOR U2496 ( .A(n2672), .B(n1958), .Z(out[642]) );
  XNOR U2497 ( .A(n2673), .B(n2674), .Z(n1958) );
  ANDN U2498 ( .B(n1492), .A(n1493), .Z(n2672) );
  XNOR U2499 ( .A(n2675), .B(n2676), .Z(n1493) );
  XNOR U2500 ( .A(n2677), .B(n2678), .Z(n1492) );
  XOR U2501 ( .A(n2679), .B(n1967), .Z(out[641]) );
  XNOR U2502 ( .A(n2680), .B(n2681), .Z(n1967) );
  ANDN U2503 ( .B(n1496), .A(n1497), .Z(n2679) );
  XNOR U2504 ( .A(n2682), .B(n2683), .Z(n1497) );
  XNOR U2505 ( .A(n2684), .B(n2685), .Z(n1496) );
  XOR U2506 ( .A(n2686), .B(n1972), .Z(out[640]) );
  XNOR U2507 ( .A(n2687), .B(n2688), .Z(n1972) );
  ANDN U2508 ( .B(n1500), .A(n1501), .Z(n2686) );
  XNOR U2509 ( .A(n2689), .B(n2690), .Z(n1501) );
  XNOR U2510 ( .A(n2691), .B(n2692), .Z(n1500) );
  XOR U2511 ( .A(n2693), .B(n2694), .Z(out[63]) );
  AND U2512 ( .A(n2695), .B(n2696), .Z(n2693) );
  XNOR U2513 ( .A(n2697), .B(n2698), .Z(out[639]) );
  ANDN U2514 ( .B(n2699), .A(n2700), .Z(n2697) );
  XNOR U2515 ( .A(n2701), .B(n2702), .Z(out[638]) );
  ANDN U2516 ( .B(n2703), .A(n2704), .Z(n2701) );
  XNOR U2517 ( .A(n2705), .B(n2706), .Z(out[637]) );
  ANDN U2518 ( .B(n2707), .A(n2708), .Z(n2705) );
  XNOR U2519 ( .A(n2709), .B(n2710), .Z(out[636]) );
  ANDN U2520 ( .B(n2711), .A(n2712), .Z(n2709) );
  XOR U2521 ( .A(n2713), .B(n2714), .Z(out[635]) );
  ANDN U2522 ( .B(n2715), .A(n2716), .Z(n2713) );
  XNOR U2523 ( .A(n2717), .B(n2718), .Z(out[634]) );
  ANDN U2524 ( .B(n2719), .A(n2720), .Z(n2717) );
  XNOR U2525 ( .A(n2721), .B(n2722), .Z(out[633]) );
  AND U2526 ( .A(n2723), .B(n2724), .Z(n2721) );
  XNOR U2527 ( .A(n2725), .B(n2726), .Z(out[632]) );
  AND U2528 ( .A(n2727), .B(n2728), .Z(n2725) );
  XNOR U2529 ( .A(n2729), .B(n2730), .Z(out[631]) );
  AND U2530 ( .A(n2731), .B(n2732), .Z(n2729) );
  XNOR U2531 ( .A(n2733), .B(n2734), .Z(out[630]) );
  AND U2532 ( .A(n2735), .B(n2736), .Z(n2733) );
  XOR U2533 ( .A(n2737), .B(n2738), .Z(out[62]) );
  AND U2534 ( .A(n2739), .B(n2740), .Z(n2737) );
  XNOR U2535 ( .A(n2741), .B(n2742), .Z(out[629]) );
  AND U2536 ( .A(n2743), .B(n2744), .Z(n2741) );
  XNOR U2537 ( .A(n2745), .B(n2746), .Z(out[628]) );
  AND U2538 ( .A(n2747), .B(n2748), .Z(n2745) );
  XNOR U2539 ( .A(n2749), .B(n2750), .Z(out[627]) );
  AND U2540 ( .A(n2751), .B(n2752), .Z(n2749) );
  XNOR U2541 ( .A(n2753), .B(n2754), .Z(out[626]) );
  AND U2542 ( .A(n2755), .B(n2756), .Z(n2753) );
  XNOR U2543 ( .A(n2757), .B(n2758), .Z(out[625]) );
  AND U2544 ( .A(n2759), .B(n2760), .Z(n2757) );
  XNOR U2545 ( .A(n2761), .B(n2762), .Z(out[624]) );
  AND U2546 ( .A(n2763), .B(n2764), .Z(n2761) );
  XNOR U2547 ( .A(n2765), .B(n2766), .Z(out[623]) );
  AND U2548 ( .A(n2767), .B(n2768), .Z(n2765) );
  XNOR U2549 ( .A(n2769), .B(n2770), .Z(out[622]) );
  AND U2550 ( .A(n2771), .B(n2772), .Z(n2769) );
  XNOR U2551 ( .A(n2773), .B(n2774), .Z(out[621]) );
  AND U2552 ( .A(n2775), .B(n2776), .Z(n2773) );
  XNOR U2553 ( .A(n2777), .B(n2778), .Z(out[620]) );
  AND U2554 ( .A(n2779), .B(n2780), .Z(n2777) );
  XOR U2555 ( .A(n2781), .B(n2782), .Z(out[61]) );
  AND U2556 ( .A(n2783), .B(n2784), .Z(n2781) );
  XNOR U2557 ( .A(n2785), .B(n2786), .Z(out[619]) );
  AND U2558 ( .A(n2787), .B(n2788), .Z(n2785) );
  XNOR U2559 ( .A(n2789), .B(n2790), .Z(out[618]) );
  AND U2560 ( .A(n2791), .B(n2792), .Z(n2789) );
  XNOR U2561 ( .A(n2793), .B(n2794), .Z(out[617]) );
  AND U2562 ( .A(n2795), .B(n2796), .Z(n2793) );
  XNOR U2563 ( .A(n2797), .B(n2798), .Z(out[616]) );
  AND U2564 ( .A(n2799), .B(n2800), .Z(n2797) );
  XNOR U2565 ( .A(n2801), .B(n2802), .Z(out[615]) );
  AND U2566 ( .A(n2803), .B(n2804), .Z(n2801) );
  XOR U2567 ( .A(n2805), .B(n2806), .Z(out[614]) );
  AND U2568 ( .A(n2807), .B(n2808), .Z(n2805) );
  XNOR U2569 ( .A(n2809), .B(n2810), .Z(out[613]) );
  AND U2570 ( .A(n2811), .B(n2812), .Z(n2809) );
  XNOR U2571 ( .A(n2813), .B(n2814), .Z(out[612]) );
  AND U2572 ( .A(n2815), .B(n2816), .Z(n2813) );
  XNOR U2573 ( .A(n2817), .B(n2818), .Z(out[611]) );
  AND U2574 ( .A(n2819), .B(n2820), .Z(n2817) );
  XNOR U2575 ( .A(n2821), .B(n2822), .Z(out[610]) );
  AND U2576 ( .A(n2823), .B(n2824), .Z(n2821) );
  XOR U2577 ( .A(n2825), .B(n2826), .Z(out[60]) );
  AND U2578 ( .A(n2827), .B(n2828), .Z(n2825) );
  XOR U2579 ( .A(n2829), .B(n2830), .Z(out[609]) );
  AND U2580 ( .A(n2831), .B(n2832), .Z(n2829) );
  XOR U2581 ( .A(n2833), .B(n2834), .Z(out[608]) );
  AND U2582 ( .A(n2835), .B(n2836), .Z(n2833) );
  XNOR U2583 ( .A(n2837), .B(n2838), .Z(out[607]) );
  ANDN U2584 ( .B(n2839), .A(n2840), .Z(n2837) );
  XOR U2585 ( .A(n2841), .B(n2842), .Z(out[606]) );
  AND U2586 ( .A(n2843), .B(n2844), .Z(n2841) );
  XNOR U2587 ( .A(n2845), .B(n2846), .Z(out[605]) );
  ANDN U2588 ( .B(n2847), .A(n2848), .Z(n2845) );
  XNOR U2589 ( .A(n2849), .B(n2850), .Z(out[604]) );
  ANDN U2590 ( .B(n2851), .A(n2852), .Z(n2849) );
  XNOR U2591 ( .A(n2853), .B(n2854), .Z(out[603]) );
  ANDN U2592 ( .B(n2855), .A(n2856), .Z(n2853) );
  XNOR U2593 ( .A(n2857), .B(n2858), .Z(out[602]) );
  AND U2594 ( .A(n2859), .B(n2860), .Z(n2857) );
  AND U2595 ( .A(n2863), .B(n2864), .Z(n2861) );
  XOR U2596 ( .A(n2865), .B(n2866), .Z(out[600]) );
  AND U2597 ( .A(n2867), .B(n2868), .Z(n2865) );
  XOR U2598 ( .A(n2869), .B(n2251), .Z(out[5]) );
  AND U2599 ( .A(n2870), .B(n2871), .Z(n2869) );
  XNOR U2600 ( .A(n2872), .B(n2873), .Z(out[59]) );
  AND U2601 ( .A(n2874), .B(n2875), .Z(n2872) );
  XOR U2602 ( .A(n2876), .B(n2877), .Z(out[599]) );
  AND U2603 ( .A(n2878), .B(n2879), .Z(n2876) );
  XOR U2604 ( .A(n2880), .B(n2881), .Z(out[598]) );
  AND U2605 ( .A(n2882), .B(n2883), .Z(n2880) );
  XOR U2606 ( .A(n2884), .B(n2885), .Z(out[597]) );
  AND U2607 ( .A(n2886), .B(n2887), .Z(n2884) );
  XOR U2608 ( .A(n2888), .B(n2889), .Z(out[596]) );
  AND U2609 ( .A(n2890), .B(n2891), .Z(n2888) );
  XNOR U2610 ( .A(n2892), .B(n2893), .Z(out[595]) );
  AND U2611 ( .A(n2894), .B(n2895), .Z(n2892) );
  XNOR U2612 ( .A(n2896), .B(n2897), .Z(out[594]) );
  AND U2613 ( .A(n2898), .B(n2899), .Z(n2896) );
  XNOR U2614 ( .A(n2900), .B(n2901), .Z(out[593]) );
  ANDN U2615 ( .B(n2902), .A(n2903), .Z(n2900) );
  XNOR U2616 ( .A(n2904), .B(n2905), .Z(out[592]) );
  ANDN U2617 ( .B(n2906), .A(n2907), .Z(n2904) );
  ANDN U2618 ( .B(n2909), .A(n2910), .Z(n2908) );
  ANDN U2619 ( .B(n2912), .A(n2913), .Z(n2911) );
  XNOR U2620 ( .A(n2914), .B(n2915), .Z(out[58]) );
  AND U2621 ( .A(n2916), .B(n2917), .Z(n2914) );
  AND U2622 ( .A(n2919), .B(n2920), .Z(n2918) );
  ANDN U2623 ( .B(n2922), .A(n2923), .Z(n2921) );
  AND U2624 ( .A(n2925), .B(n2926), .Z(n2924) );
  XNOR U2625 ( .A(n2927), .B(n2928), .Z(out[586]) );
  AND U2626 ( .A(n2929), .B(n2930), .Z(n2927) );
  AND U2627 ( .A(n2932), .B(n2933), .Z(n2931) );
  XNOR U2628 ( .A(n2934), .B(n2935), .Z(out[584]) );
  AND U2629 ( .A(n2936), .B(n2937), .Z(n2934) );
  XNOR U2630 ( .A(n2938), .B(n2939), .Z(out[583]) );
  AND U2631 ( .A(n2940), .B(n2941), .Z(n2938) );
  XNOR U2632 ( .A(n2942), .B(n2943), .Z(out[582]) );
  AND U2633 ( .A(n2944), .B(n2945), .Z(n2942) );
  XNOR U2634 ( .A(n2946), .B(n2947), .Z(out[581]) );
  AND U2635 ( .A(n2948), .B(n2949), .Z(n2946) );
  XNOR U2636 ( .A(n2950), .B(n2951), .Z(out[580]) );
  AND U2637 ( .A(n2952), .B(n2953), .Z(n2950) );
  XNOR U2638 ( .A(n2954), .B(n2955), .Z(out[57]) );
  AND U2639 ( .A(n2956), .B(n2957), .Z(n2954) );
  XNOR U2640 ( .A(n2958), .B(n2959), .Z(out[579]) );
  ANDN U2641 ( .B(n2960), .A(n2961), .Z(n2958) );
  XNOR U2642 ( .A(n2962), .B(n2963), .Z(out[578]) );
  ANDN U2643 ( .B(n2964), .A(n2965), .Z(n2962) );
  XNOR U2644 ( .A(n2966), .B(n2967), .Z(out[577]) );
  ANDN U2645 ( .B(n2968), .A(n2969), .Z(n2966) );
  XNOR U2646 ( .A(n2970), .B(n2971), .Z(out[576]) );
  ANDN U2647 ( .B(n2972), .A(n2973), .Z(n2970) );
  XNOR U2648 ( .A(n2974), .B(n2699), .Z(out[575]) );
  AND U2649 ( .A(n2700), .B(n2975), .Z(n2974) );
  XNOR U2650 ( .A(n2976), .B(n2703), .Z(out[574]) );
  AND U2651 ( .A(n2704), .B(n2977), .Z(n2976) );
  XNOR U2652 ( .A(n2978), .B(n2707), .Z(out[573]) );
  AND U2653 ( .A(n2708), .B(n2979), .Z(n2978) );
  XNOR U2654 ( .A(n2980), .B(n2711), .Z(out[572]) );
  AND U2655 ( .A(n2712), .B(n2981), .Z(n2980) );
  XNOR U2656 ( .A(n2982), .B(n2715), .Z(out[571]) );
  AND U2657 ( .A(n2716), .B(n2983), .Z(n2982) );
  XNOR U2658 ( .A(n2984), .B(n2719), .Z(out[570]) );
  AND U2659 ( .A(n2720), .B(n2985), .Z(n2984) );
  XNOR U2660 ( .A(n2986), .B(n2987), .Z(out[56]) );
  AND U2661 ( .A(n2988), .B(n2989), .Z(n2986) );
  XNOR U2662 ( .A(n2990), .B(n2723), .Z(out[569]) );
  XNOR U2663 ( .A(n2992), .B(n2727), .Z(out[568]) );
  XNOR U2664 ( .A(n2994), .B(n2731), .Z(out[567]) );
  AND U2665 ( .A(n2995), .B(n2996), .Z(n2994) );
  XNOR U2666 ( .A(n2997), .B(n2735), .Z(out[566]) );
  AND U2667 ( .A(n2998), .B(n2999), .Z(n2997) );
  XNOR U2668 ( .A(n3000), .B(n2743), .Z(out[565]) );
  AND U2669 ( .A(n3001), .B(n3002), .Z(n3000) );
  XNOR U2670 ( .A(n3003), .B(n2747), .Z(out[564]) );
  AND U2671 ( .A(n3004), .B(n3005), .Z(n3003) );
  XNOR U2672 ( .A(n3006), .B(n2751), .Z(out[563]) );
  AND U2673 ( .A(n3007), .B(n3008), .Z(n3006) );
  XNOR U2674 ( .A(n3009), .B(n2755), .Z(out[562]) );
  AND U2675 ( .A(n3010), .B(n3011), .Z(n3009) );
  XNOR U2676 ( .A(n3012), .B(n2759), .Z(out[561]) );
  AND U2677 ( .A(n3013), .B(n3014), .Z(n3012) );
  XNOR U2678 ( .A(n3015), .B(n2763), .Z(out[560]) );
  AND U2679 ( .A(n3016), .B(n3017), .Z(n3015) );
  XNOR U2680 ( .A(n3018), .B(n3019), .Z(out[55]) );
  AND U2681 ( .A(n3020), .B(n3021), .Z(n3018) );
  XNOR U2682 ( .A(n3022), .B(n2767), .Z(out[559]) );
  AND U2683 ( .A(n3023), .B(n3024), .Z(n3022) );
  XNOR U2684 ( .A(n3025), .B(n2771), .Z(out[558]) );
  AND U2685 ( .A(n3026), .B(n3027), .Z(n3025) );
  XNOR U2686 ( .A(n3028), .B(n2775), .Z(out[557]) );
  AND U2687 ( .A(n3029), .B(n3030), .Z(n3028) );
  XNOR U2688 ( .A(n3031), .B(n2779), .Z(out[556]) );
  AND U2689 ( .A(n3032), .B(n3033), .Z(n3031) );
  XNOR U2690 ( .A(n3034), .B(n2787), .Z(out[555]) );
  XNOR U2691 ( .A(n3036), .B(n2791), .Z(out[554]) );
  AND U2692 ( .A(n3037), .B(n3038), .Z(n3036) );
  XNOR U2693 ( .A(n3039), .B(n2796), .Z(out[553]) );
  ANDN U2694 ( .B(n3040), .A(n2795), .Z(n3039) );
  XNOR U2695 ( .A(n3041), .B(n2799), .Z(out[552]) );
  XNOR U2696 ( .A(n3043), .B(n2803), .Z(out[551]) );
  XNOR U2697 ( .A(n3045), .B(n2807), .Z(out[550]) );
  XNOR U2698 ( .A(n3047), .B(n3048), .Z(out[54]) );
  AND U2699 ( .A(n3049), .B(n3050), .Z(n3047) );
  XNOR U2700 ( .A(n3051), .B(n2811), .Z(out[549]) );
  AND U2701 ( .A(n3052), .B(n3053), .Z(n3051) );
  XNOR U2702 ( .A(n3054), .B(n2815), .Z(out[548]) );
  AND U2703 ( .A(n3055), .B(n3056), .Z(n3054) );
  XNOR U2704 ( .A(n3057), .B(n2819), .Z(out[547]) );
  AND U2705 ( .A(n3058), .B(n3059), .Z(n3057) );
  XNOR U2706 ( .A(n3060), .B(n2823), .Z(out[546]) );
  AND U2707 ( .A(n3061), .B(n3062), .Z(n3060) );
  XNOR U2708 ( .A(n3063), .B(n2831), .Z(out[545]) );
  AND U2709 ( .A(n3064), .B(n3065), .Z(n3063) );
  XNOR U2710 ( .A(n3066), .B(n2835), .Z(out[544]) );
  AND U2711 ( .A(n3067), .B(n3068), .Z(n3066) );
  XNOR U2712 ( .A(n3069), .B(n2839), .Z(out[543]) );
  AND U2713 ( .A(n2840), .B(n3070), .Z(n3069) );
  XNOR U2714 ( .A(n3071), .B(n2843), .Z(out[542]) );
  AND U2715 ( .A(n3072), .B(n3073), .Z(n3071) );
  XNOR U2716 ( .A(n3074), .B(n2847), .Z(out[541]) );
  AND U2717 ( .A(n2848), .B(n3075), .Z(n3074) );
  XNOR U2718 ( .A(n3076), .B(n2851), .Z(out[540]) );
  AND U2719 ( .A(n2852), .B(n3077), .Z(n3076) );
  XNOR U2720 ( .A(n3078), .B(n3079), .Z(out[53]) );
  AND U2721 ( .A(n3080), .B(n3081), .Z(n3078) );
  XNOR U2722 ( .A(n3082), .B(n2855), .Z(out[539]) );
  AND U2723 ( .A(n2856), .B(n3083), .Z(n3082) );
  XNOR U2724 ( .A(n3084), .B(n2859), .Z(out[538]) );
  AND U2725 ( .A(n3085), .B(n3086), .Z(n3084) );
  XNOR U2726 ( .A(n3087), .B(n2864), .Z(out[537]) );
  ANDN U2727 ( .B(n3088), .A(n2863), .Z(n3087) );
  XNOR U2728 ( .A(n3089), .B(n2867), .Z(out[536]) );
  AND U2729 ( .A(n3090), .B(n3091), .Z(n3089) );
  XNOR U2730 ( .A(n3092), .B(n2878), .Z(out[535]) );
  AND U2731 ( .A(n3093), .B(n3094), .Z(n3092) );
  XNOR U2732 ( .A(n3095), .B(n2882), .Z(out[534]) );
  AND U2733 ( .A(n3096), .B(n3097), .Z(n3095) );
  XNOR U2734 ( .A(n3098), .B(n2886), .Z(out[533]) );
  XNOR U2735 ( .A(n3100), .B(n2890), .Z(out[532]) );
  XNOR U2736 ( .A(n3102), .B(n2894), .Z(out[531]) );
  XNOR U2737 ( .A(n3104), .B(n2898), .Z(out[530]) );
  XNOR U2738 ( .A(n3106), .B(n3107), .Z(out[52]) );
  AND U2739 ( .A(n3108), .B(n3109), .Z(n3106) );
  XNOR U2740 ( .A(n3110), .B(n2902), .Z(out[529]) );
  AND U2741 ( .A(n2903), .B(n3111), .Z(n3110) );
  XNOR U2742 ( .A(n3112), .B(n2906), .Z(out[528]) );
  AND U2743 ( .A(n2907), .B(n3113), .Z(n3112) );
  XNOR U2744 ( .A(n3114), .B(n2909), .Z(out[527]) );
  AND U2745 ( .A(n2910), .B(n3115), .Z(n3114) );
  XNOR U2746 ( .A(n3116), .B(n2912), .Z(out[526]) );
  AND U2747 ( .A(n2913), .B(n3117), .Z(n3116) );
  XNOR U2748 ( .A(n3118), .B(n2920), .Z(out[525]) );
  ANDN U2749 ( .B(n3119), .A(n2919), .Z(n3118) );
  XNOR U2750 ( .A(n3120), .B(n2922), .Z(out[524]) );
  AND U2751 ( .A(n2923), .B(n3121), .Z(n3120) );
  XNOR U2752 ( .A(n3122), .B(n2926), .Z(out[523]) );
  ANDN U2753 ( .B(n3123), .A(n2925), .Z(n3122) );
  XNOR U2754 ( .A(n3124), .B(n2930), .Z(out[522]) );
  ANDN U2755 ( .B(n3125), .A(n2929), .Z(n3124) );
  XNOR U2756 ( .A(n3126), .B(n2933), .Z(out[521]) );
  ANDN U2757 ( .B(n3127), .A(n2932), .Z(n3126) );
  XNOR U2758 ( .A(n3128), .B(n2937), .Z(out[520]) );
  NOR U2759 ( .A(n3129), .B(n2936), .Z(n3128) );
  AND U2760 ( .A(n3132), .B(n3133), .Z(n3130) );
  XNOR U2761 ( .A(n3134), .B(n2941), .Z(out[519]) );
  NOR U2762 ( .A(n3135), .B(n2940), .Z(n3134) );
  XNOR U2763 ( .A(n3136), .B(n2945), .Z(out[518]) );
  NOR U2764 ( .A(n3137), .B(n2944), .Z(n3136) );
  XNOR U2765 ( .A(n3138), .B(n2949), .Z(out[517]) );
  NOR U2766 ( .A(n3139), .B(n2948), .Z(n3138) );
  XNOR U2767 ( .A(n3140), .B(n2953), .Z(out[516]) );
  NOR U2768 ( .A(n3141), .B(n2952), .Z(n3140) );
  XNOR U2769 ( .A(n3142), .B(n2960), .Z(out[515]) );
  AND U2770 ( .A(n2961), .B(n3143), .Z(n3142) );
  XNOR U2771 ( .A(n3144), .B(n2964), .Z(out[514]) );
  AND U2772 ( .A(n2965), .B(n3145), .Z(n3144) );
  XNOR U2773 ( .A(n3146), .B(n2968), .Z(out[513]) );
  AND U2774 ( .A(n2969), .B(n3147), .Z(n3146) );
  XNOR U2775 ( .A(n3148), .B(n2972), .Z(out[512]) );
  AND U2776 ( .A(n2973), .B(n3149), .Z(n3148) );
  XNOR U2777 ( .A(n3150), .B(n2700), .Z(out[511]) );
  XNOR U2778 ( .A(n3151), .B(n2293), .Z(n2700) );
  AND U2779 ( .A(n3152), .B(n3153), .Z(n3150) );
  XNOR U2780 ( .A(n3154), .B(n2704), .Z(out[510]) );
  XNOR U2781 ( .A(n3155), .B(n2300), .Z(n2704) );
  AND U2782 ( .A(n3156), .B(n3157), .Z(n3154) );
  AND U2783 ( .A(n3160), .B(n3161), .Z(n3158) );
  XNOR U2784 ( .A(n3162), .B(n2708), .Z(out[509]) );
  XNOR U2785 ( .A(n3163), .B(n2307), .Z(n2708) );
  AND U2786 ( .A(n3164), .B(n3165), .Z(n3162) );
  XNOR U2787 ( .A(n3166), .B(n2712), .Z(out[508]) );
  XNOR U2788 ( .A(n3167), .B(n2314), .Z(n2712) );
  AND U2789 ( .A(n3168), .B(n3169), .Z(n3166) );
  XNOR U2790 ( .A(n3170), .B(n2716), .Z(out[507]) );
  XNOR U2791 ( .A(n3171), .B(n2321), .Z(n2716) );
  AND U2792 ( .A(n3172), .B(n3173), .Z(n3170) );
  XNOR U2793 ( .A(n3174), .B(n2720), .Z(out[506]) );
  XNOR U2794 ( .A(n3175), .B(n2332), .Z(n2720) );
  AND U2795 ( .A(n3176), .B(n3177), .Z(n3174) );
  XOR U2796 ( .A(n3178), .B(n2724), .Z(out[505]) );
  XOR U2797 ( .A(n3179), .B(n2337), .Z(n2724) );
  ANDN U2798 ( .B(n3180), .A(n2991), .Z(n3178) );
  XOR U2799 ( .A(n3181), .B(n2728), .Z(out[504]) );
  XOR U2800 ( .A(n3182), .B(n2344), .Z(n2728) );
  ANDN U2801 ( .B(n3183), .A(n2993), .Z(n3181) );
  XOR U2802 ( .A(n3184), .B(n2732), .Z(out[503]) );
  IV U2803 ( .A(n2996), .Z(n2732) );
  XNOR U2804 ( .A(n3185), .B(n2351), .Z(n2996) );
  ANDN U2805 ( .B(n3186), .A(n2995), .Z(n3184) );
  XOR U2806 ( .A(n3187), .B(n2736), .Z(out[502]) );
  IV U2807 ( .A(n2999), .Z(n2736) );
  XNOR U2808 ( .A(n3188), .B(n2358), .Z(n2999) );
  ANDN U2809 ( .B(n3189), .A(n2998), .Z(n3187) );
  XOR U2810 ( .A(n3190), .B(n2744), .Z(out[501]) );
  IV U2811 ( .A(n3002), .Z(n2744) );
  XNOR U2812 ( .A(n3191), .B(n2365), .Z(n3002) );
  ANDN U2813 ( .B(n3192), .A(n3001), .Z(n3190) );
  XOR U2814 ( .A(n3193), .B(n2748), .Z(out[500]) );
  IV U2815 ( .A(n3005), .Z(n2748) );
  XNOR U2816 ( .A(n3194), .B(n2374), .Z(n3005) );
  ANDN U2817 ( .B(n3195), .A(n3004), .Z(n3193) );
  XNOR U2818 ( .A(n3196), .B(n2324), .Z(out[4]) );
  AND U2819 ( .A(n3197), .B(n3198), .Z(n3196) );
  XNOR U2820 ( .A(n3199), .B(n3200), .Z(out[49]) );
  AND U2821 ( .A(n3201), .B(n3202), .Z(n3199) );
  XOR U2822 ( .A(n3203), .B(n2752), .Z(out[499]) );
  IV U2823 ( .A(n3008), .Z(n2752) );
  XNOR U2824 ( .A(n3204), .B(n2379), .Z(n3008) );
  ANDN U2825 ( .B(n3205), .A(n3007), .Z(n3203) );
  XOR U2826 ( .A(n3206), .B(n2756), .Z(out[498]) );
  IV U2827 ( .A(n3011), .Z(n2756) );
  XNOR U2828 ( .A(n3207), .B(n2386), .Z(n3011) );
  ANDN U2829 ( .B(n3208), .A(n3010), .Z(n3206) );
  XOR U2830 ( .A(n3209), .B(n2760), .Z(out[497]) );
  IV U2831 ( .A(n3014), .Z(n2760) );
  XNOR U2832 ( .A(n3210), .B(n2395), .Z(n3014) );
  ANDN U2833 ( .B(n3211), .A(n3013), .Z(n3209) );
  XOR U2834 ( .A(n3212), .B(n2764), .Z(out[496]) );
  IV U2835 ( .A(n3017), .Z(n2764) );
  XNOR U2836 ( .A(n3213), .B(n2404), .Z(n3017) );
  ANDN U2837 ( .B(n3214), .A(n3016), .Z(n3212) );
  XOR U2838 ( .A(n3215), .B(n2768), .Z(out[495]) );
  IV U2839 ( .A(n3024), .Z(n2768) );
  XNOR U2840 ( .A(n3216), .B(n2413), .Z(n3024) );
  ANDN U2841 ( .B(n3217), .A(n3023), .Z(n3215) );
  XOR U2842 ( .A(n3218), .B(n2772), .Z(out[494]) );
  IV U2843 ( .A(n3027), .Z(n2772) );
  XNOR U2844 ( .A(n3219), .B(n2420), .Z(n3027) );
  ANDN U2845 ( .B(n3220), .A(n3026), .Z(n3218) );
  XOR U2846 ( .A(n3221), .B(n2776), .Z(out[493]) );
  IV U2847 ( .A(n3030), .Z(n2776) );
  XNOR U2848 ( .A(n3222), .B(n2427), .Z(n3030) );
  ANDN U2849 ( .B(n3223), .A(n3029), .Z(n3221) );
  XOR U2850 ( .A(n3224), .B(n2780), .Z(out[492]) );
  IV U2851 ( .A(n3033), .Z(n2780) );
  XNOR U2852 ( .A(n3225), .B(n2434), .Z(n3033) );
  ANDN U2853 ( .B(n3226), .A(n3032), .Z(n3224) );
  XOR U2854 ( .A(n3227), .B(n2788), .Z(out[491]) );
  XOR U2855 ( .A(n2438), .B(n3228), .Z(n2788) );
  ANDN U2856 ( .B(n3229), .A(n3035), .Z(n3227) );
  XOR U2857 ( .A(n3230), .B(n2792), .Z(out[490]) );
  IV U2858 ( .A(n3038), .Z(n2792) );
  XNOR U2859 ( .A(n2445), .B(n3231), .Z(n3038) );
  ANDN U2860 ( .B(n3232), .A(n3037), .Z(n3230) );
  XNOR U2861 ( .A(n3233), .B(n3234), .Z(out[48]) );
  AND U2862 ( .A(n3235), .B(n3236), .Z(n3233) );
  XOR U2863 ( .A(n3237), .B(n2795), .Z(out[489]) );
  XNOR U2864 ( .A(n3238), .B(n3239), .Z(n2795) );
  ANDN U2865 ( .B(n3240), .A(n3040), .Z(n3237) );
  XOR U2866 ( .A(n3241), .B(n2800), .Z(out[488]) );
  XNOR U2867 ( .A(n3242), .B(n2462), .Z(n2800) );
  ANDN U2868 ( .B(n3243), .A(n3042), .Z(n3241) );
  XOR U2869 ( .A(n3244), .B(n2804), .Z(out[487]) );
  XNOR U2870 ( .A(n3245), .B(n2469), .Z(n2804) );
  ANDN U2871 ( .B(n3246), .A(n3044), .Z(n3244) );
  XOR U2872 ( .A(n3247), .B(n2808), .Z(out[486]) );
  XNOR U2873 ( .A(n3248), .B(n2480), .Z(n2808) );
  ANDN U2874 ( .B(n3249), .A(n3046), .Z(n3247) );
  XOR U2875 ( .A(n3250), .B(n2812), .Z(out[485]) );
  IV U2876 ( .A(n3053), .Z(n2812) );
  XNOR U2877 ( .A(n3251), .B(n2487), .Z(n3053) );
  ANDN U2878 ( .B(n3252), .A(n3052), .Z(n3250) );
  XOR U2879 ( .A(n3253), .B(n2816), .Z(out[484]) );
  IV U2880 ( .A(n3056), .Z(n2816) );
  XNOR U2881 ( .A(n3254), .B(n2492), .Z(n3056) );
  ANDN U2882 ( .B(n3255), .A(n3055), .Z(n3253) );
  XOR U2883 ( .A(n3256), .B(n2820), .Z(out[483]) );
  IV U2884 ( .A(n3059), .Z(n2820) );
  XNOR U2885 ( .A(n3257), .B(n2499), .Z(n3059) );
  ANDN U2886 ( .B(n3258), .A(n3058), .Z(n3256) );
  XOR U2887 ( .A(n3259), .B(n2824), .Z(out[482]) );
  IV U2888 ( .A(n3062), .Z(n2824) );
  XNOR U2889 ( .A(n3260), .B(n2508), .Z(n3062) );
  ANDN U2890 ( .B(n3261), .A(n3061), .Z(n3259) );
  XOR U2891 ( .A(n3262), .B(n2832), .Z(out[481]) );
  IV U2892 ( .A(n3065), .Z(n2832) );
  XNOR U2893 ( .A(n3263), .B(n2515), .Z(n3065) );
  NOR U2894 ( .A(n3264), .B(n3064), .Z(n3262) );
  XOR U2895 ( .A(n3265), .B(n2836), .Z(out[480]) );
  IV U2896 ( .A(n3068), .Z(n2836) );
  XNOR U2897 ( .A(n3266), .B(n2522), .Z(n3068) );
  NOR U2898 ( .A(n3267), .B(n3067), .Z(n3265) );
  XNOR U2899 ( .A(n3268), .B(n3269), .Z(out[47]) );
  AND U2900 ( .A(n3270), .B(n3271), .Z(n3268) );
  XNOR U2901 ( .A(n3272), .B(n2840), .Z(out[479]) );
  XNOR U2902 ( .A(n3273), .B(n2529), .Z(n2840) );
  AND U2903 ( .A(n3274), .B(n3275), .Z(n3272) );
  XOR U2904 ( .A(n3276), .B(n2844), .Z(out[478]) );
  IV U2905 ( .A(n3073), .Z(n2844) );
  XNOR U2906 ( .A(n3277), .B(n2536), .Z(n3073) );
  NOR U2907 ( .A(n3278), .B(n3072), .Z(n3276) );
  XNOR U2908 ( .A(n3279), .B(n2848), .Z(out[477]) );
  XNOR U2909 ( .A(n3280), .B(n2543), .Z(n2848) );
  XNOR U2910 ( .A(n3282), .B(n2852), .Z(out[476]) );
  XNOR U2911 ( .A(n3283), .B(n3284), .Z(n2852) );
  XNOR U2912 ( .A(n3286), .B(n2856), .Z(out[475]) );
  XNOR U2913 ( .A(n3287), .B(n2561), .Z(n2856) );
  XOR U2914 ( .A(n3289), .B(n2860), .Z(out[474]) );
  IV U2915 ( .A(n3086), .Z(n2860) );
  XOR U2916 ( .A(n3290), .B(n2568), .Z(n3086) );
  NOR U2917 ( .A(n3291), .B(n3085), .Z(n3289) );
  XOR U2918 ( .A(n3292), .B(n2863), .Z(out[473]) );
  XOR U2919 ( .A(n3293), .B(n2575), .Z(n2863) );
  AND U2920 ( .A(n3294), .B(n3295), .Z(n3292) );
  XOR U2921 ( .A(n3296), .B(n2868), .Z(out[472]) );
  IV U2922 ( .A(n3091), .Z(n2868) );
  XOR U2923 ( .A(n3297), .B(n2582), .Z(n3091) );
  NOR U2924 ( .A(n3298), .B(n3090), .Z(n3296) );
  XOR U2925 ( .A(n3299), .B(n2879), .Z(out[471]) );
  IV U2926 ( .A(n3094), .Z(n2879) );
  XOR U2927 ( .A(n3300), .B(n2589), .Z(n3094) );
  NOR U2928 ( .A(n3301), .B(n3093), .Z(n3299) );
  XOR U2929 ( .A(n3302), .B(n2883), .Z(out[470]) );
  IV U2930 ( .A(n3097), .Z(n2883) );
  XOR U2931 ( .A(n3303), .B(n2596), .Z(n3097) );
  NOR U2932 ( .A(n3304), .B(n3096), .Z(n3302) );
  XOR U2933 ( .A(n3305), .B(n3306), .Z(out[46]) );
  AND U2934 ( .A(n3307), .B(n3308), .Z(n3305) );
  XOR U2935 ( .A(n3309), .B(n2887), .Z(out[469]) );
  XOR U2936 ( .A(n3310), .B(n2603), .Z(n2887) );
  NOR U2937 ( .A(n3311), .B(n3099), .Z(n3309) );
  XOR U2938 ( .A(n3312), .B(n2891), .Z(out[468]) );
  XOR U2939 ( .A(n3313), .B(n2610), .Z(n2891) );
  NOR U2940 ( .A(n3314), .B(n3101), .Z(n3312) );
  XOR U2941 ( .A(n3315), .B(n2895), .Z(out[467]) );
  XOR U2942 ( .A(n3316), .B(n2617), .Z(n2895) );
  NOR U2943 ( .A(n3317), .B(n3103), .Z(n3315) );
  XOR U2944 ( .A(n3318), .B(n2899), .Z(out[466]) );
  XOR U2945 ( .A(n3319), .B(n2629), .Z(n2899) );
  NOR U2946 ( .A(n3320), .B(n3105), .Z(n3318) );
  XNOR U2947 ( .A(n3321), .B(n2903), .Z(out[465]) );
  XNOR U2948 ( .A(n2635), .B(n3322), .Z(n2903) );
  AND U2949 ( .A(n3323), .B(n3324), .Z(n3321) );
  XNOR U2950 ( .A(n3325), .B(n2907), .Z(out[464]) );
  XNOR U2951 ( .A(n3326), .B(n2643), .Z(n2907) );
  AND U2952 ( .A(n3327), .B(n3328), .Z(n3325) );
  XNOR U2953 ( .A(n3329), .B(n2910), .Z(out[463]) );
  XNOR U2954 ( .A(n3330), .B(n2650), .Z(n2910) );
  AND U2955 ( .A(n3331), .B(n3332), .Z(n3329) );
  XNOR U2956 ( .A(n3333), .B(n2913), .Z(out[462]) );
  XNOR U2957 ( .A(n3334), .B(n2657), .Z(n2913) );
  AND U2958 ( .A(n3335), .B(n3336), .Z(n3333) );
  XOR U2959 ( .A(n3337), .B(n2919), .Z(out[461]) );
  XNOR U2960 ( .A(n3338), .B(n3339), .Z(n2919) );
  AND U2961 ( .A(n3340), .B(n3341), .Z(n3337) );
  XNOR U2962 ( .A(n3342), .B(n2923), .Z(out[460]) );
  XNOR U2963 ( .A(n3343), .B(n3344), .Z(n2923) );
  AND U2964 ( .A(n3345), .B(n3346), .Z(n3342) );
  XOR U2965 ( .A(n3347), .B(n3348), .Z(out[45]) );
  AND U2966 ( .A(n3349), .B(n3350), .Z(n3347) );
  XOR U2967 ( .A(n3351), .B(n2925), .Z(out[459]) );
  XNOR U2968 ( .A(n3352), .B(n3353), .Z(n2925) );
  AND U2969 ( .A(n3354), .B(n3355), .Z(n3351) );
  XOR U2970 ( .A(n3356), .B(n2929), .Z(out[458]) );
  XNOR U2971 ( .A(n3357), .B(n3358), .Z(n2929) );
  AND U2972 ( .A(n3359), .B(n3360), .Z(n3356) );
  XOR U2973 ( .A(n3361), .B(n2932), .Z(out[457]) );
  XNOR U2974 ( .A(n3362), .B(n3363), .Z(n2932) );
  AND U2975 ( .A(n3364), .B(n3365), .Z(n3361) );
  XOR U2976 ( .A(n3366), .B(n2936), .Z(out[456]) );
  XNOR U2977 ( .A(n2222), .B(n3367), .Z(n2936) );
  AND U2978 ( .A(n3129), .B(n3368), .Z(n3366) );
  XOR U2979 ( .A(n3369), .B(n2940), .Z(out[455]) );
  XNOR U2980 ( .A(n2229), .B(n3370), .Z(n2940) );
  AND U2981 ( .A(n3135), .B(n3371), .Z(n3369) );
  XOR U2982 ( .A(n3372), .B(n2944), .Z(out[454]) );
  XNOR U2983 ( .A(n2236), .B(n3373), .Z(n2944) );
  AND U2984 ( .A(n3137), .B(n3374), .Z(n3372) );
  XOR U2985 ( .A(n3375), .B(n2948), .Z(out[453]) );
  XNOR U2986 ( .A(n2243), .B(n3376), .Z(n2948) );
  AND U2987 ( .A(n3139), .B(n3377), .Z(n3375) );
  XOR U2988 ( .A(n3378), .B(n2952), .Z(out[452]) );
  XNOR U2989 ( .A(n2257), .B(n3379), .Z(n2952) );
  AND U2990 ( .A(n3141), .B(n3380), .Z(n3378) );
  XNOR U2991 ( .A(n3381), .B(n2961), .Z(out[451]) );
  XNOR U2992 ( .A(n3382), .B(n2265), .Z(n2961) );
  AND U2993 ( .A(n3383), .B(n3384), .Z(n3381) );
  XNOR U2994 ( .A(n3385), .B(n2965), .Z(out[450]) );
  XNOR U2995 ( .A(n3386), .B(n2272), .Z(n2965) );
  AND U2996 ( .A(n3387), .B(n3388), .Z(n3385) );
  XNOR U2997 ( .A(n3389), .B(n3390), .Z(out[44]) );
  AND U2998 ( .A(n3391), .B(n3392), .Z(n3389) );
  XNOR U2999 ( .A(n3393), .B(n2969), .Z(out[449]) );
  XNOR U3000 ( .A(n3394), .B(n2279), .Z(n2969) );
  AND U3001 ( .A(n3395), .B(n3396), .Z(n3393) );
  XNOR U3002 ( .A(n3397), .B(n2973), .Z(out[448]) );
  XNOR U3003 ( .A(n3398), .B(n2286), .Z(n2973) );
  AND U3004 ( .A(n3399), .B(n3400), .Z(n3397) );
  XOR U3005 ( .A(n3401), .B(n2975), .Z(out[447]) );
  IV U3006 ( .A(n3153), .Z(n2975) );
  XNOR U3007 ( .A(n3402), .B(n2291), .Z(n3153) );
  NOR U3008 ( .A(n2698), .B(n3152), .Z(n3401) );
  XOR U3009 ( .A(n3403), .B(n2977), .Z(out[446]) );
  IV U3010 ( .A(n3157), .Z(n2977) );
  XNOR U3011 ( .A(n3404), .B(n2298), .Z(n3157) );
  NOR U3012 ( .A(n2702), .B(n3156), .Z(n3403) );
  XOR U3013 ( .A(n3405), .B(n2979), .Z(out[445]) );
  IV U3014 ( .A(n3165), .Z(n2979) );
  XNOR U3015 ( .A(n3406), .B(n2305), .Z(n3165) );
  NOR U3016 ( .A(n2706), .B(n3164), .Z(n3405) );
  XOR U3017 ( .A(n3407), .B(n2981), .Z(out[444]) );
  IV U3018 ( .A(n3169), .Z(n2981) );
  XNOR U3019 ( .A(n3408), .B(n2312), .Z(n3169) );
  NOR U3020 ( .A(n2710), .B(n3168), .Z(n3407) );
  XOR U3021 ( .A(n3409), .B(n2983), .Z(out[443]) );
  IV U3022 ( .A(n3173), .Z(n2983) );
  XNOR U3023 ( .A(n3410), .B(n2319), .Z(n3173) );
  ANDN U3024 ( .B(n2714), .A(n3172), .Z(n3409) );
  XOR U3025 ( .A(n3411), .B(n2985), .Z(out[442]) );
  IV U3026 ( .A(n3177), .Z(n2985) );
  XNOR U3027 ( .A(n3412), .B(n2330), .Z(n3177) );
  NOR U3028 ( .A(n2718), .B(n3176), .Z(n3411) );
  XOR U3029 ( .A(n3413), .B(n2991), .Z(out[441]) );
  XOR U3030 ( .A(n2338), .B(n3414), .Z(n2991) );
  NOR U3031 ( .A(n2722), .B(n3180), .Z(n3413) );
  XOR U3032 ( .A(n3415), .B(n2993), .Z(out[440]) );
  XOR U3033 ( .A(n2345), .B(n3416), .Z(n2993) );
  NOR U3034 ( .A(n2726), .B(n3183), .Z(n3415) );
  XNOR U3035 ( .A(n3417), .B(n3418), .Z(out[43]) );
  AND U3036 ( .A(n3419), .B(n3420), .Z(n3417) );
  XOR U3037 ( .A(n3421), .B(n2995), .Z(out[439]) );
  XOR U3038 ( .A(n2352), .B(n3422), .Z(n2995) );
  NOR U3039 ( .A(n2730), .B(n3186), .Z(n3421) );
  XOR U3040 ( .A(n3423), .B(n2998), .Z(out[438]) );
  XOR U3041 ( .A(n2359), .B(n3424), .Z(n2998) );
  NOR U3042 ( .A(n2734), .B(n3189), .Z(n3423) );
  XOR U3043 ( .A(n3425), .B(n3001), .Z(out[437]) );
  XOR U3044 ( .A(n2366), .B(n3426), .Z(n3001) );
  NOR U3045 ( .A(n2742), .B(n3192), .Z(n3425) );
  XOR U3046 ( .A(n3427), .B(n3004), .Z(out[436]) );
  XOR U3047 ( .A(n2371), .B(n3428), .Z(n3004) );
  NOR U3048 ( .A(n2746), .B(n3195), .Z(n3427) );
  XOR U3049 ( .A(n3429), .B(n3007), .Z(out[435]) );
  XOR U3050 ( .A(n2380), .B(n3430), .Z(n3007) );
  NOR U3051 ( .A(n2750), .B(n3205), .Z(n3429) );
  XOR U3052 ( .A(n3431), .B(n3010), .Z(out[434]) );
  XOR U3053 ( .A(n2387), .B(n3432), .Z(n3010) );
  NOR U3054 ( .A(n2754), .B(n3208), .Z(n3431) );
  XOR U3055 ( .A(n3433), .B(n3013), .Z(out[433]) );
  XOR U3056 ( .A(n2392), .B(n3434), .Z(n3013) );
  NOR U3057 ( .A(n2758), .B(n3211), .Z(n3433) );
  XOR U3058 ( .A(n3435), .B(n3016), .Z(out[432]) );
  XNOR U3059 ( .A(n2405), .B(n3436), .Z(n3016) );
  NOR U3060 ( .A(n2762), .B(n3214), .Z(n3435) );
  XOR U3061 ( .A(n3437), .B(n3023), .Z(out[431]) );
  XOR U3062 ( .A(n3438), .B(n2411), .Z(n3023) );
  NOR U3063 ( .A(n2766), .B(n3217), .Z(n3437) );
  XOR U3064 ( .A(n3439), .B(n3026), .Z(out[430]) );
  XOR U3065 ( .A(n3440), .B(n2418), .Z(n3026) );
  NOR U3066 ( .A(n2770), .B(n3220), .Z(n3439) );
  XNOR U3067 ( .A(n3441), .B(n3442), .Z(out[42]) );
  AND U3068 ( .A(n3443), .B(n3444), .Z(n3441) );
  XOR U3069 ( .A(n3445), .B(n3029), .Z(out[429]) );
  XOR U3070 ( .A(n2424), .B(n3446), .Z(n3029) );
  NOR U3071 ( .A(n2774), .B(n3223), .Z(n3445) );
  XOR U3072 ( .A(n3447), .B(n3032), .Z(out[428]) );
  XOR U3073 ( .A(n2431), .B(n3448), .Z(n3032) );
  NOR U3074 ( .A(n2778), .B(n3226), .Z(n3447) );
  XOR U3075 ( .A(n3449), .B(n3035), .Z(out[427]) );
  XOR U3076 ( .A(n2440), .B(n3450), .Z(n3035) );
  NOR U3077 ( .A(n3229), .B(n2786), .Z(n3449) );
  XOR U3078 ( .A(n3451), .B(n3037), .Z(out[426]) );
  XOR U3079 ( .A(n2447), .B(n3452), .Z(n3037) );
  NOR U3080 ( .A(n2790), .B(n3232), .Z(n3451) );
  XOR U3081 ( .A(n3453), .B(n3040), .Z(out[425]) );
  XOR U3082 ( .A(n2452), .B(n3454), .Z(n3040) );
  NOR U3083 ( .A(n2794), .B(n3240), .Z(n3453) );
  XOR U3084 ( .A(n3455), .B(n3042), .Z(out[424]) );
  XOR U3085 ( .A(n2459), .B(n3456), .Z(n3042) );
  NOR U3086 ( .A(n2798), .B(n3243), .Z(n3455) );
  XOR U3087 ( .A(n3457), .B(n3044), .Z(out[423]) );
  XOR U3088 ( .A(n2466), .B(n3458), .Z(n3044) );
  NOR U3089 ( .A(n2802), .B(n3246), .Z(n3457) );
  XOR U3090 ( .A(n3459), .B(n3046), .Z(out[422]) );
  XOR U3091 ( .A(n2477), .B(n3460), .Z(n3046) );
  ANDN U3092 ( .B(n2806), .A(n3249), .Z(n3459) );
  XOR U3093 ( .A(n3461), .B(n3052), .Z(out[421]) );
  XOR U3094 ( .A(n2484), .B(n3462), .Z(n3052) );
  NOR U3095 ( .A(n2810), .B(n3252), .Z(n3461) );
  XOR U3096 ( .A(n3463), .B(n3055), .Z(out[420]) );
  XOR U3097 ( .A(n2493), .B(n3464), .Z(n3055) );
  NOR U3098 ( .A(n2814), .B(n3255), .Z(n3463) );
  XNOR U3099 ( .A(n3465), .B(n3466), .Z(out[41]) );
  AND U3100 ( .A(n3467), .B(n3468), .Z(n3465) );
  XOR U3101 ( .A(n3469), .B(n3058), .Z(out[419]) );
  XOR U3102 ( .A(n2500), .B(n3470), .Z(n3058) );
  NOR U3103 ( .A(n3258), .B(n2818), .Z(n3469) );
  XOR U3104 ( .A(n3471), .B(n3061), .Z(out[418]) );
  XOR U3105 ( .A(n2505), .B(n3472), .Z(n3061) );
  NOR U3106 ( .A(n2822), .B(n3261), .Z(n3471) );
  XOR U3107 ( .A(n3473), .B(n3064), .Z(out[417]) );
  XOR U3108 ( .A(n3474), .B(n2513), .Z(n3064) );
  AND U3109 ( .A(n3264), .B(n2830), .Z(n3473) );
  IV U3110 ( .A(n3475), .Z(n2830) );
  XOR U3111 ( .A(n3476), .B(n3067), .Z(out[416]) );
  XNOR U3112 ( .A(n2519), .B(n3477), .Z(n3067) );
  AND U3113 ( .A(n3267), .B(n2834), .Z(n3476) );
  IV U3114 ( .A(n3478), .Z(n2834) );
  XOR U3115 ( .A(n3479), .B(n3070), .Z(out[415]) );
  IV U3116 ( .A(n3275), .Z(n3070) );
  XOR U3117 ( .A(n2526), .B(n3480), .Z(n3275) );
  XOR U3118 ( .A(n3481), .B(n3072), .Z(out[414]) );
  XNOR U3119 ( .A(n2533), .B(n3482), .Z(n3072) );
  AND U3120 ( .A(n3278), .B(n2842), .Z(n3481) );
  IV U3121 ( .A(n3483), .Z(n2842) );
  XOR U3122 ( .A(n3484), .B(n3075), .Z(out[413]) );
  XOR U3123 ( .A(n3485), .B(n3486), .Z(n3075) );
  XOR U3124 ( .A(n3487), .B(n3077), .Z(out[412]) );
  XOR U3125 ( .A(n3488), .B(n3489), .Z(n3077) );
  XOR U3126 ( .A(n3490), .B(n3083), .Z(out[411]) );
  XOR U3127 ( .A(n3491), .B(n3492), .Z(n3083) );
  XOR U3128 ( .A(n3493), .B(n3085), .Z(out[410]) );
  XOR U3129 ( .A(n2565), .B(n3494), .Z(n3085) );
  ANDN U3130 ( .B(n3291), .A(n2858), .Z(n3493) );
  XNOR U3131 ( .A(n3495), .B(n3496), .Z(out[40]) );
  XOR U3132 ( .A(n3499), .B(n3088), .Z(out[409]) );
  IV U3133 ( .A(n3295), .Z(n3088) );
  XNOR U3134 ( .A(n3500), .B(n2573), .Z(n3295) );
  NOR U3135 ( .A(n2862), .B(n3294), .Z(n3499) );
  XOR U3136 ( .A(n3501), .B(n3090), .Z(out[408]) );
  XOR U3137 ( .A(n3502), .B(n2580), .Z(n3090) );
  AND U3138 ( .A(n3298), .B(n2866), .Z(n3501) );
  IV U3139 ( .A(n3503), .Z(n2866) );
  XOR U3140 ( .A(n3504), .B(n3093), .Z(out[407]) );
  XOR U3141 ( .A(n3505), .B(n2587), .Z(n3093) );
  AND U3142 ( .A(n3301), .B(n2877), .Z(n3504) );
  IV U3143 ( .A(n3506), .Z(n2877) );
  XOR U3144 ( .A(n3507), .B(n3096), .Z(out[406]) );
  XOR U3145 ( .A(n3508), .B(n2594), .Z(n3096) );
  AND U3146 ( .A(n3304), .B(n2881), .Z(n3507) );
  IV U3147 ( .A(n3509), .Z(n2881) );
  XOR U3148 ( .A(n3510), .B(n3099), .Z(out[405]) );
  XOR U3149 ( .A(n3511), .B(n2601), .Z(n3099) );
  AND U3150 ( .A(n3311), .B(n2885), .Z(n3510) );
  IV U3151 ( .A(n3512), .Z(n2885) );
  XOR U3152 ( .A(n3513), .B(n3101), .Z(out[404]) );
  XOR U3153 ( .A(n3514), .B(n2608), .Z(n3101) );
  AND U3154 ( .A(n3314), .B(n2889), .Z(n3513) );
  IV U3155 ( .A(n3515), .Z(n2889) );
  XOR U3156 ( .A(n3516), .B(n3103), .Z(out[403]) );
  XOR U3157 ( .A(n3517), .B(n2615), .Z(n3103) );
  ANDN U3158 ( .B(n3317), .A(n2893), .Z(n3516) );
  XOR U3159 ( .A(n3518), .B(n3105), .Z(out[402]) );
  XOR U3160 ( .A(n3519), .B(n2627), .Z(n3105) );
  ANDN U3161 ( .B(n3320), .A(n2897), .Z(n3518) );
  XOR U3162 ( .A(n3520), .B(n3111), .Z(out[401]) );
  IV U3163 ( .A(n3324), .Z(n3111) );
  XNOR U3164 ( .A(n3521), .B(n2634), .Z(n3324) );
  NOR U3165 ( .A(n3323), .B(n2901), .Z(n3520) );
  XOR U3166 ( .A(n3522), .B(n3113), .Z(out[400]) );
  IV U3167 ( .A(n3328), .Z(n3113) );
  XNOR U3168 ( .A(n3523), .B(n2641), .Z(n3328) );
  NOR U3169 ( .A(n3327), .B(n2905), .Z(n3522) );
  XOR U3170 ( .A(n3524), .B(n2399), .Z(out[3]) );
  AND U3171 ( .A(n3525), .B(n3526), .Z(n3524) );
  XNOR U3172 ( .A(n3527), .B(n3528), .Z(out[39]) );
  XOR U3173 ( .A(n3531), .B(n3115), .Z(out[399]) );
  IV U3174 ( .A(n3332), .Z(n3115) );
  XNOR U3175 ( .A(n3532), .B(n2648), .Z(n3332) );
  XOR U3176 ( .A(n3534), .B(n3117), .Z(out[398]) );
  IV U3177 ( .A(n3336), .Z(n3117) );
  XNOR U3178 ( .A(n3535), .B(n2655), .Z(n3336) );
  XOR U3179 ( .A(n3537), .B(n3119), .Z(out[397]) );
  IV U3180 ( .A(n3341), .Z(n3119) );
  XNOR U3181 ( .A(n3538), .B(n2662), .Z(n3341) );
  XOR U3182 ( .A(n3540), .B(n3121), .Z(out[396]) );
  IV U3183 ( .A(n3346), .Z(n3121) );
  XNOR U3184 ( .A(n3541), .B(n2669), .Z(n3346) );
  XOR U3185 ( .A(n3543), .B(n3123), .Z(out[395]) );
  IV U3186 ( .A(n3355), .Z(n3123) );
  XNOR U3187 ( .A(n3544), .B(n2676), .Z(n3355) );
  XOR U3188 ( .A(n3546), .B(n3125), .Z(out[394]) );
  IV U3189 ( .A(n3360), .Z(n3125) );
  XNOR U3190 ( .A(n3547), .B(n2683), .Z(n3360) );
  NOR U3191 ( .A(n2928), .B(n3359), .Z(n3546) );
  XOR U3192 ( .A(n3548), .B(n3127), .Z(out[393]) );
  IV U3193 ( .A(n3365), .Z(n3127) );
  XNOR U3194 ( .A(n3549), .B(n2690), .Z(n3365) );
  XNOR U3195 ( .A(n3551), .B(n3129), .Z(out[392]) );
  XNOR U3196 ( .A(n3552), .B(n2221), .Z(n3129) );
  XNOR U3197 ( .A(n3553), .B(n3135), .Z(out[391]) );
  XNOR U3198 ( .A(n3554), .B(n3555), .Z(n3135) );
  XNOR U3199 ( .A(n3556), .B(n3137), .Z(out[390]) );
  XNOR U3200 ( .A(n3557), .B(n3558), .Z(n3137) );
  XNOR U3201 ( .A(n3559), .B(n3560), .Z(out[38]) );
  XNOR U3202 ( .A(n3563), .B(n3139), .Z(out[389]) );
  XNOR U3203 ( .A(n3564), .B(n2242), .Z(n3139) );
  XNOR U3204 ( .A(n3565), .B(n3141), .Z(out[388]) );
  XNOR U3205 ( .A(n3566), .B(n2256), .Z(n3141) );
  XOR U3206 ( .A(n3567), .B(n3143), .Z(out[387]) );
  IV U3207 ( .A(n3384), .Z(n3143) );
  XNOR U3208 ( .A(n3568), .B(n2263), .Z(n3384) );
  NOR U3209 ( .A(n2959), .B(n3383), .Z(n3567) );
  XOR U3210 ( .A(n3569), .B(n3145), .Z(out[386]) );
  IV U3211 ( .A(n3388), .Z(n3145) );
  XNOR U3212 ( .A(n3570), .B(n2270), .Z(n3388) );
  NOR U3213 ( .A(n3387), .B(n2963), .Z(n3569) );
  XOR U3214 ( .A(n3571), .B(n3147), .Z(out[385]) );
  IV U3215 ( .A(n3396), .Z(n3147) );
  XNOR U3216 ( .A(n3572), .B(n2277), .Z(n3396) );
  NOR U3217 ( .A(n2967), .B(n3395), .Z(n3571) );
  XOR U3218 ( .A(n3573), .B(n3149), .Z(out[384]) );
  IV U3219 ( .A(n3400), .Z(n3149) );
  XNOR U3220 ( .A(n3574), .B(n2284), .Z(n3400) );
  NOR U3221 ( .A(n2971), .B(n3399), .Z(n3573) );
  XOR U3222 ( .A(n3575), .B(n3152), .Z(out[383]) );
  XNOR U3223 ( .A(n1811), .B(n3576), .Z(n3152) );
  ANDN U3224 ( .B(n2698), .A(n2699), .Z(n3575) );
  XOR U3225 ( .A(n3577), .B(n2356), .Z(n2699) );
  XOR U3226 ( .A(n3578), .B(n2052), .Z(n2698) );
  XOR U3227 ( .A(n3579), .B(n3156), .Z(out[382]) );
  XOR U3228 ( .A(n1823), .B(n3580), .Z(n3156) );
  ANDN U3229 ( .B(n2702), .A(n2703), .Z(n3579) );
  XOR U3230 ( .A(n3581), .B(n2363), .Z(n2703) );
  XOR U3231 ( .A(n3582), .B(n2056), .Z(n2702) );
  XOR U3232 ( .A(n3583), .B(n3164), .Z(out[381]) );
  XOR U3233 ( .A(n1827), .B(n3584), .Z(n3164) );
  ANDN U3234 ( .B(n2706), .A(n2707), .Z(n3583) );
  XOR U3235 ( .A(n3585), .B(n2370), .Z(n2707) );
  IV U3236 ( .A(n3586), .Z(n2370) );
  XOR U3237 ( .A(n3587), .B(n2060), .Z(n2706) );
  XOR U3238 ( .A(n3588), .B(n3168), .Z(out[380]) );
  XOR U3239 ( .A(n1831), .B(n3589), .Z(n3168) );
  ANDN U3240 ( .B(n2710), .A(n2711), .Z(n3588) );
  XOR U3241 ( .A(n3590), .B(n2377), .Z(n2711) );
  IV U3242 ( .A(n3591), .Z(n2377) );
  XOR U3243 ( .A(n3592), .B(n2063), .Z(n2710) );
  XNOR U3244 ( .A(n3593), .B(n3594), .Z(out[37]) );
  XOR U3245 ( .A(n3597), .B(n3172), .Z(out[379]) );
  XOR U3246 ( .A(n1835), .B(n3598), .Z(n3172) );
  NOR U3247 ( .A(n2715), .B(n2714), .Z(n3597) );
  XOR U3248 ( .A(n3599), .B(n2066), .Z(n2714) );
  XOR U3249 ( .A(n3600), .B(n2384), .Z(n2715) );
  XOR U3250 ( .A(n3601), .B(n3176), .Z(out[378]) );
  XOR U3251 ( .A(n1839), .B(n3602), .Z(n3176) );
  ANDN U3252 ( .B(n2718), .A(n2719), .Z(n3601) );
  XOR U3253 ( .A(n3603), .B(n2391), .Z(n2719) );
  XOR U3254 ( .A(n3604), .B(n2070), .Z(n2718) );
  XOR U3255 ( .A(n3605), .B(n3180), .Z(out[377]) );
  XOR U3256 ( .A(n1843), .B(n3606), .Z(n3180) );
  ANDN U3257 ( .B(n2722), .A(n2723), .Z(n3605) );
  XOR U3258 ( .A(n3607), .B(n2402), .Z(n2723) );
  XOR U3259 ( .A(n3608), .B(n2073), .Z(n2722) );
  XOR U3260 ( .A(n3609), .B(n3183), .Z(out[376]) );
  XOR U3261 ( .A(n1847), .B(n3610), .Z(n3183) );
  ANDN U3262 ( .B(n2726), .A(n2727), .Z(n3609) );
  XOR U3263 ( .A(n3611), .B(n2409), .Z(n2727) );
  XOR U3264 ( .A(n3612), .B(n2076), .Z(n2726) );
  XOR U3265 ( .A(n3613), .B(n3186), .Z(out[375]) );
  XOR U3266 ( .A(n1852), .B(n3614), .Z(n3186) );
  ANDN U3267 ( .B(n2730), .A(n2731), .Z(n3613) );
  XOR U3268 ( .A(n3615), .B(n2416), .Z(n2731) );
  XOR U3269 ( .A(n3616), .B(n2080), .Z(n2730) );
  XOR U3270 ( .A(n3617), .B(n3189), .Z(out[374]) );
  XOR U3271 ( .A(n1856), .B(n3618), .Z(n3189) );
  ANDN U3272 ( .B(n2734), .A(n2735), .Z(n3617) );
  XNOR U3273 ( .A(n3619), .B(n2423), .Z(n2735) );
  XOR U3274 ( .A(n3620), .B(n2087), .Z(n2734) );
  XOR U3275 ( .A(n3621), .B(n3192), .Z(out[373]) );
  XOR U3276 ( .A(n1860), .B(n3622), .Z(n3192) );
  ANDN U3277 ( .B(n2742), .A(n2743), .Z(n3621) );
  XOR U3278 ( .A(n3623), .B(n2430), .Z(n2743) );
  XOR U3279 ( .A(n3624), .B(n2090), .Z(n2742) );
  XOR U3280 ( .A(n3625), .B(n3195), .Z(out[372]) );
  XOR U3281 ( .A(n1868), .B(n3626), .Z(n3195) );
  ANDN U3282 ( .B(n2746), .A(n2747), .Z(n3625) );
  XNOR U3283 ( .A(n3627), .B(n2437), .Z(n2747) );
  XOR U3284 ( .A(n3628), .B(n2094), .Z(n2746) );
  XOR U3285 ( .A(n3629), .B(n3205), .Z(out[371]) );
  XOR U3286 ( .A(n1872), .B(n3630), .Z(n3205) );
  ANDN U3287 ( .B(n2750), .A(n2751), .Z(n3629) );
  XNOR U3288 ( .A(n3631), .B(n2444), .Z(n2751) );
  XOR U3289 ( .A(n3632), .B(n2098), .Z(n2750) );
  XOR U3290 ( .A(n3633), .B(n3208), .Z(out[370]) );
  XOR U3291 ( .A(n1876), .B(n3634), .Z(n3208) );
  ANDN U3292 ( .B(n2754), .A(n2755), .Z(n3633) );
  XNOR U3293 ( .A(n3635), .B(n2451), .Z(n2755) );
  XOR U3294 ( .A(n3636), .B(n2101), .Z(n2754) );
  XNOR U3295 ( .A(n3637), .B(n3638), .Z(out[36]) );
  XOR U3296 ( .A(n3641), .B(n3211), .Z(out[369]) );
  XNOR U3297 ( .A(n3642), .B(n3643), .Z(n3211) );
  ANDN U3298 ( .B(n2758), .A(n2759), .Z(n3641) );
  XNOR U3299 ( .A(n3644), .B(n2458), .Z(n2759) );
  XOR U3300 ( .A(n3645), .B(n2105), .Z(n2758) );
  XOR U3301 ( .A(n3646), .B(n3214), .Z(out[368]) );
  XNOR U3302 ( .A(n1885), .B(n3647), .Z(n3214) );
  ANDN U3303 ( .B(n2762), .A(n2763), .Z(n3646) );
  XNOR U3304 ( .A(n3648), .B(n2465), .Z(n2763) );
  XOR U3305 ( .A(n3649), .B(n2108), .Z(n2762) );
  XOR U3306 ( .A(n3650), .B(n3217), .Z(out[367]) );
  XNOR U3307 ( .A(n1889), .B(n3651), .Z(n3217) );
  ANDN U3308 ( .B(n2766), .A(n2767), .Z(n3650) );
  XNOR U3309 ( .A(n3652), .B(n2476), .Z(n2767) );
  XOR U3310 ( .A(n3653), .B(n2111), .Z(n2766) );
  XOR U3311 ( .A(n3654), .B(n3220), .Z(out[366]) );
  XOR U3312 ( .A(n1893), .B(n3655), .Z(n3220) );
  ANDN U3313 ( .B(n2770), .A(n2771), .Z(n3654) );
  XOR U3314 ( .A(n3656), .B(n2483), .Z(n2771) );
  XNOR U3315 ( .A(n2114), .B(n3657), .Z(n2770) );
  XOR U3316 ( .A(n3658), .B(n3223), .Z(out[365]) );
  XOR U3317 ( .A(n1897), .B(n3659), .Z(n3223) );
  ANDN U3318 ( .B(n2774), .A(n2775), .Z(n3658) );
  XOR U3319 ( .A(n3660), .B(n2490), .Z(n2775) );
  XOR U3320 ( .A(n2118), .B(n3661), .Z(n2774) );
  XOR U3321 ( .A(n3662), .B(n3226), .Z(out[364]) );
  XOR U3322 ( .A(n1901), .B(n3663), .Z(n3226) );
  ANDN U3323 ( .B(n2778), .A(n2779), .Z(n3662) );
  XOR U3324 ( .A(n3664), .B(n2497), .Z(n2779) );
  XNOR U3325 ( .A(n3665), .B(n2125), .Z(n2778) );
  XOR U3326 ( .A(n3666), .B(n3229), .Z(out[363]) );
  XOR U3327 ( .A(n1906), .B(n3667), .Z(n3229) );
  ANDN U3328 ( .B(n2786), .A(n2787), .Z(n3666) );
  XNOR U3329 ( .A(n3668), .B(n2504), .Z(n2787) );
  XNOR U3330 ( .A(n2127), .B(n3669), .Z(n2786) );
  XOR U3331 ( .A(n3670), .B(n3232), .Z(out[362]) );
  XOR U3332 ( .A(n1914), .B(n3671), .Z(n3232) );
  ANDN U3333 ( .B(n2790), .A(n2791), .Z(n3670) );
  XOR U3334 ( .A(n3672), .B(n2511), .Z(n2791) );
  XNOR U3335 ( .A(n2131), .B(n3673), .Z(n2790) );
  XOR U3336 ( .A(n3674), .B(n3240), .Z(out[361]) );
  XOR U3337 ( .A(n1919), .B(n3675), .Z(n3240) );
  ANDN U3338 ( .B(n2794), .A(n2796), .Z(n3674) );
  XOR U3339 ( .A(n3676), .B(n2518), .Z(n2796) );
  XNOR U3340 ( .A(n2135), .B(n3677), .Z(n2794) );
  XOR U3341 ( .A(n3678), .B(n3243), .Z(out[360]) );
  XOR U3342 ( .A(n1923), .B(n3679), .Z(n3243) );
  ANDN U3343 ( .B(n2798), .A(n2799), .Z(n3678) );
  XOR U3344 ( .A(n3680), .B(n2525), .Z(n2799) );
  XNOR U3345 ( .A(n2139), .B(n3681), .Z(n2798) );
  XNOR U3346 ( .A(n3682), .B(n1045), .Z(out[35]) );
  XOR U3347 ( .A(n3684), .B(n3246), .Z(out[359]) );
  XOR U3348 ( .A(n1927), .B(n3685), .Z(n3246) );
  ANDN U3349 ( .B(n2802), .A(n2803), .Z(n3684) );
  XOR U3350 ( .A(n3686), .B(n2532), .Z(n2803) );
  XNOR U3351 ( .A(n2143), .B(n3687), .Z(n2802) );
  XOR U3352 ( .A(n3688), .B(n3249), .Z(out[358]) );
  XOR U3353 ( .A(n1931), .B(n3689), .Z(n3249) );
  NOR U3354 ( .A(n2807), .B(n2806), .Z(n3688) );
  XNOR U3355 ( .A(n2147), .B(n3690), .Z(n2806) );
  XOR U3356 ( .A(n3691), .B(n2539), .Z(n2807) );
  XOR U3357 ( .A(n3692), .B(n3252), .Z(out[357]) );
  XOR U3358 ( .A(n1936), .B(n3693), .Z(n3252) );
  ANDN U3359 ( .B(n2810), .A(n2811), .Z(n3692) );
  XOR U3360 ( .A(n3694), .B(n2550), .Z(n2811) );
  XOR U3361 ( .A(n3695), .B(n2152), .Z(n2810) );
  XOR U3362 ( .A(n3696), .B(n3255), .Z(out[356]) );
  XOR U3363 ( .A(n1941), .B(n3697), .Z(n3255) );
  ANDN U3364 ( .B(n2814), .A(n2815), .Z(n3696) );
  XOR U3365 ( .A(n3698), .B(n2557), .Z(n2815) );
  XNOR U3366 ( .A(n3699), .B(n2155), .Z(n2814) );
  XOR U3367 ( .A(n3700), .B(n3258), .Z(out[355]) );
  XOR U3368 ( .A(n1946), .B(n3701), .Z(n3258) );
  ANDN U3369 ( .B(n2818), .A(n2819), .Z(n3700) );
  XOR U3370 ( .A(n3702), .B(n2564), .Z(n2819) );
  XNOR U3371 ( .A(n3703), .B(n2159), .Z(n2818) );
  XOR U3372 ( .A(n3704), .B(n3261), .Z(out[354]) );
  XNOR U3373 ( .A(n1951), .B(n3705), .Z(n3261) );
  ANDN U3374 ( .B(n2822), .A(n2823), .Z(n3704) );
  XOR U3375 ( .A(n3706), .B(n3707), .Z(n2823) );
  XNOR U3376 ( .A(n3708), .B(n2164), .Z(n2822) );
  XNOR U3377 ( .A(n3709), .B(n3264), .Z(out[353]) );
  XOR U3378 ( .A(n3710), .B(n1957), .Z(n3264) );
  ANDN U3379 ( .B(n3475), .A(n2831), .Z(n3709) );
  XOR U3380 ( .A(n3711), .B(n2578), .Z(n2831) );
  XNOR U3381 ( .A(n3712), .B(n2168), .Z(n3475) );
  XNOR U3382 ( .A(n3713), .B(n3267), .Z(out[352]) );
  XOR U3383 ( .A(n3714), .B(n1966), .Z(n3267) );
  ANDN U3384 ( .B(n3478), .A(n2835), .Z(n3713) );
  XOR U3385 ( .A(n3715), .B(n2585), .Z(n2835) );
  XNOR U3386 ( .A(n3716), .B(n2172), .Z(n3478) );
  XOR U3387 ( .A(n3717), .B(n3274), .Z(out[351]) );
  XNOR U3388 ( .A(n3718), .B(n1971), .Z(n3274) );
  ANDN U3389 ( .B(n2838), .A(n2839), .Z(n3717) );
  XOR U3390 ( .A(n3719), .B(n2592), .Z(n2839) );
  XOR U3391 ( .A(n3720), .B(n2175), .Z(n2838) );
  XNOR U3392 ( .A(n3721), .B(n3278), .Z(out[350]) );
  XOR U3393 ( .A(n3722), .B(n1658), .Z(n3278) );
  ANDN U3394 ( .B(n3483), .A(n2843), .Z(n3721) );
  XNOR U3395 ( .A(n2598), .B(n3723), .Z(n2843) );
  XNOR U3396 ( .A(n3724), .B(n2178), .Z(n3483) );
  XNOR U3397 ( .A(n3725), .B(n1089), .Z(out[34]) );
  XOR U3398 ( .A(n3727), .B(n3281), .Z(out[349]) );
  XNOR U3399 ( .A(n3728), .B(n1663), .Z(n3281) );
  ANDN U3400 ( .B(n2846), .A(n2847), .Z(n3727) );
  XNOR U3401 ( .A(n2605), .B(n3729), .Z(n2847) );
  XNOR U3402 ( .A(n3730), .B(n2181), .Z(n2846) );
  XOR U3403 ( .A(n3731), .B(n3285), .Z(out[348]) );
  XNOR U3404 ( .A(n3732), .B(n1671), .Z(n3285) );
  ANDN U3405 ( .B(n2850), .A(n2851), .Z(n3731) );
  XNOR U3406 ( .A(n2612), .B(n3733), .Z(n2851) );
  XNOR U3407 ( .A(n3734), .B(n2184), .Z(n2850) );
  XOR U3408 ( .A(n3735), .B(n3288), .Z(out[347]) );
  XNOR U3409 ( .A(n3736), .B(n1675), .Z(n3288) );
  ANDN U3410 ( .B(n2854), .A(n2855), .Z(n3735) );
  XOR U3411 ( .A(n3737), .B(n2625), .Z(n2855) );
  XNOR U3412 ( .A(n3738), .B(n2188), .Z(n2854) );
  XNOR U3413 ( .A(n3739), .B(n3291), .Z(out[346]) );
  XNOR U3414 ( .A(n3740), .B(n1680), .Z(n3291) );
  ANDN U3415 ( .B(n2858), .A(n2859), .Z(n3739) );
  XOR U3416 ( .A(n3741), .B(n3742), .Z(n2859) );
  XOR U3417 ( .A(n3743), .B(n2191), .Z(n2858) );
  XOR U3418 ( .A(n3744), .B(n3294), .Z(out[345]) );
  XOR U3419 ( .A(n3745), .B(n1685), .Z(n3294) );
  ANDN U3420 ( .B(n2862), .A(n2864), .Z(n3744) );
  XOR U3421 ( .A(n3746), .B(n2639), .Z(n2864) );
  XNOR U3422 ( .A(n3747), .B(n2194), .Z(n2862) );
  XNOR U3423 ( .A(n3748), .B(n3298), .Z(out[344]) );
  XOR U3424 ( .A(n3749), .B(n1690), .Z(n3298) );
  ANDN U3425 ( .B(n3503), .A(n2867), .Z(n3748) );
  XOR U3426 ( .A(n3750), .B(n2646), .Z(n2867) );
  XNOR U3427 ( .A(n3751), .B(n2201), .Z(n3503) );
  XNOR U3428 ( .A(n3752), .B(n3301), .Z(out[343]) );
  XOR U3429 ( .A(n3753), .B(n1695), .Z(n3301) );
  ANDN U3430 ( .B(n3506), .A(n2878), .Z(n3752) );
  XOR U3431 ( .A(n3754), .B(n2653), .Z(n2878) );
  XNOR U3432 ( .A(n3755), .B(n2204), .Z(n3506) );
  XNOR U3433 ( .A(n3756), .B(n3304), .Z(out[342]) );
  XNOR U3434 ( .A(n3757), .B(n1700), .Z(n3304) );
  ANDN U3435 ( .B(n3509), .A(n2882), .Z(n3756) );
  XOR U3436 ( .A(n3758), .B(n2660), .Z(n2882) );
  XNOR U3437 ( .A(n3759), .B(n2207), .Z(n3509) );
  XNOR U3438 ( .A(n3760), .B(n3311), .Z(out[341]) );
  XNOR U3439 ( .A(n3761), .B(n1705), .Z(n3311) );
  ANDN U3440 ( .B(n3512), .A(n2886), .Z(n3760) );
  XOR U3441 ( .A(n3762), .B(n2667), .Z(n2886) );
  XNOR U3442 ( .A(n3763), .B(n2210), .Z(n3512) );
  XNOR U3443 ( .A(n3764), .B(n3314), .Z(out[340]) );
  XNOR U3444 ( .A(n3765), .B(n1710), .Z(n3314) );
  ANDN U3445 ( .B(n3515), .A(n2890), .Z(n3764) );
  XOR U3446 ( .A(n3766), .B(n2674), .Z(n2890) );
  XNOR U3447 ( .A(n3767), .B(n2213), .Z(n3515) );
  XOR U3448 ( .A(n3768), .B(n1134), .Z(out[33]) );
  AND U3449 ( .A(n3769), .B(n3770), .Z(n3768) );
  XNOR U3450 ( .A(n3771), .B(n3317), .Z(out[339]) );
  XNOR U3451 ( .A(n3772), .B(n1715), .Z(n3317) );
  ANDN U3452 ( .B(n2893), .A(n2894), .Z(n3771) );
  XOR U3453 ( .A(n3773), .B(n2681), .Z(n2894) );
  XNOR U3454 ( .A(n3774), .B(n2216), .Z(n2893) );
  XNOR U3455 ( .A(n3775), .B(n3320), .Z(out[338]) );
  XOR U3456 ( .A(n3776), .B(n1724), .Z(n3320) );
  ANDN U3457 ( .B(n2897), .A(n2898), .Z(n3775) );
  XOR U3458 ( .A(n3777), .B(n2688), .Z(n2898) );
  XNOR U3459 ( .A(n3778), .B(n1976), .Z(n2897) );
  XOR U3460 ( .A(n3779), .B(n3323), .Z(out[337]) );
  XNOR U3461 ( .A(n3780), .B(n1728), .Z(n3323) );
  ANDN U3462 ( .B(n2901), .A(n2902), .Z(n3779) );
  XOR U3463 ( .A(n3781), .B(n2219), .Z(n2902) );
  XNOR U3464 ( .A(n3782), .B(n1979), .Z(n2901) );
  XOR U3465 ( .A(n3783), .B(n3327), .Z(out[336]) );
  XNOR U3466 ( .A(n3784), .B(n1732), .Z(n3327) );
  ANDN U3467 ( .B(n2905), .A(n2906), .Z(n3783) );
  XOR U3468 ( .A(n3785), .B(n2226), .Z(n2906) );
  XNOR U3469 ( .A(n3786), .B(n1982), .Z(n2905) );
  XOR U3470 ( .A(n3787), .B(n3331), .Z(out[335]) );
  XNOR U3471 ( .A(n3788), .B(n1737), .Z(n3331) );
  ANDN U3472 ( .B(n3533), .A(n2909), .Z(n3787) );
  XOR U3473 ( .A(n3789), .B(n2233), .Z(n2909) );
  XNOR U3474 ( .A(n3790), .B(n1985), .Z(n3533) );
  XOR U3475 ( .A(n3791), .B(n3335), .Z(out[334]) );
  XNOR U3476 ( .A(n3792), .B(n1742), .Z(n3335) );
  ANDN U3477 ( .B(n3536), .A(n2912), .Z(n3791) );
  XNOR U3478 ( .A(n3793), .B(n2240), .Z(n2912) );
  XNOR U3479 ( .A(n3794), .B(n1988), .Z(n3536) );
  XOR U3480 ( .A(n3795), .B(n3340), .Z(out[333]) );
  XNOR U3481 ( .A(n3796), .B(n1747), .Z(n3340) );
  ANDN U3482 ( .B(n3539), .A(n2920), .Z(n3795) );
  XOR U3483 ( .A(n3797), .B(n2254), .Z(n2920) );
  XNOR U3484 ( .A(n3798), .B(n1992), .Z(n3539) );
  XOR U3485 ( .A(n3799), .B(n3345), .Z(out[332]) );
  XNOR U3486 ( .A(n3800), .B(n1752), .Z(n3345) );
  ANDN U3487 ( .B(n3542), .A(n2922), .Z(n3799) );
  XOR U3488 ( .A(n3801), .B(n2261), .Z(n2922) );
  IV U3489 ( .A(n3802), .Z(n2261) );
  XNOR U3490 ( .A(n3803), .B(n1995), .Z(n3542) );
  XOR U3491 ( .A(n3804), .B(n3354), .Z(out[331]) );
  XNOR U3492 ( .A(n3805), .B(n1757), .Z(n3354) );
  ANDN U3493 ( .B(n3545), .A(n2926), .Z(n3804) );
  XOR U3494 ( .A(n3806), .B(n2268), .Z(n2926) );
  XNOR U3495 ( .A(n3807), .B(n1998), .Z(n3545) );
  XOR U3496 ( .A(n3808), .B(n3359), .Z(out[330]) );
  XOR U3497 ( .A(n1761), .B(n3809), .Z(n3359) );
  ANDN U3498 ( .B(n2928), .A(n2930), .Z(n3808) );
  XOR U3499 ( .A(n3810), .B(n2275), .Z(n2930) );
  XNOR U3500 ( .A(n3811), .B(n2005), .Z(n2928) );
  XNOR U3501 ( .A(n3812), .B(n1177), .Z(out[32]) );
  XOR U3502 ( .A(n3814), .B(n3364), .Z(out[329]) );
  XOR U3503 ( .A(n3815), .B(n1766), .Z(n3364) );
  ANDN U3504 ( .B(n3550), .A(n2933), .Z(n3814) );
  XOR U3505 ( .A(n3816), .B(n2282), .Z(n2933) );
  XNOR U3506 ( .A(n3817), .B(n2009), .Z(n3550) );
  XOR U3507 ( .A(n3818), .B(n3368), .Z(out[328]) );
  XOR U3508 ( .A(n3819), .B(n1775), .Z(n3368) );
  ANDN U3509 ( .B(n2935), .A(n2937), .Z(n3818) );
  XOR U3510 ( .A(n3820), .B(n2289), .Z(n2937) );
  XNOR U3511 ( .A(n3821), .B(n2013), .Z(n2935) );
  XOR U3512 ( .A(n3822), .B(n3371), .Z(out[327]) );
  XOR U3513 ( .A(n3823), .B(n1780), .Z(n3371) );
  ANDN U3514 ( .B(n2939), .A(n2941), .Z(n3822) );
  XOR U3515 ( .A(n3824), .B(n2296), .Z(n2941) );
  XOR U3516 ( .A(n3825), .B(n2017), .Z(n2939) );
  XOR U3517 ( .A(n3826), .B(n3374), .Z(out[326]) );
  XOR U3518 ( .A(n3827), .B(n1784), .Z(n3374) );
  ANDN U3519 ( .B(n2943), .A(n2945), .Z(n3826) );
  XOR U3520 ( .A(n3828), .B(n2303), .Z(n2945) );
  XOR U3521 ( .A(n3829), .B(n2021), .Z(n2943) );
  XOR U3522 ( .A(n3830), .B(n3377), .Z(out[325]) );
  XOR U3523 ( .A(n3831), .B(n1788), .Z(n3377) );
  ANDN U3524 ( .B(n2947), .A(n2949), .Z(n3830) );
  XNOR U3525 ( .A(n3832), .B(n2310), .Z(n2949) );
  XOR U3526 ( .A(n3833), .B(n2024), .Z(n2947) );
  XOR U3527 ( .A(n3834), .B(n3380), .Z(out[324]) );
  XOR U3528 ( .A(n3835), .B(n1792), .Z(n3380) );
  ANDN U3529 ( .B(n2951), .A(n2953), .Z(n3834) );
  XOR U3530 ( .A(n3836), .B(n2317), .Z(n2953) );
  XOR U3531 ( .A(n3837), .B(n2028), .Z(n2951) );
  XOR U3532 ( .A(n3838), .B(n3383), .Z(out[323]) );
  XNOR U3533 ( .A(n1795), .B(n3839), .Z(n3383) );
  ANDN U3534 ( .B(n2959), .A(n2960), .Z(n3838) );
  XOR U3535 ( .A(n3840), .B(n2328), .Z(n2960) );
  XOR U3536 ( .A(n3841), .B(n2032), .Z(n2959) );
  XOR U3537 ( .A(n3842), .B(n3387), .Z(out[322]) );
  XOR U3538 ( .A(n3843), .B(n1800), .Z(n3387) );
  ANDN U3539 ( .B(n2963), .A(n2964), .Z(n3842) );
  XOR U3540 ( .A(n3844), .B(n2335), .Z(n2964) );
  XOR U3541 ( .A(n3845), .B(n2036), .Z(n2963) );
  XOR U3542 ( .A(n3846), .B(n3395), .Z(out[321]) );
  XOR U3543 ( .A(n1803), .B(n3847), .Z(n3395) );
  ANDN U3544 ( .B(n2967), .A(n2968), .Z(n3846) );
  XOR U3545 ( .A(n3848), .B(n2342), .Z(n2968) );
  XOR U3546 ( .A(n3849), .B(n2040), .Z(n2967) );
  XOR U3547 ( .A(n3850), .B(n3399), .Z(out[320]) );
  XOR U3548 ( .A(n1807), .B(n3851), .Z(n3399) );
  ANDN U3549 ( .B(n2971), .A(n2972), .Z(n3850) );
  XOR U3550 ( .A(n3852), .B(n2349), .Z(n2972) );
  XOR U3551 ( .A(n3853), .B(n2048), .Z(n2971) );
  XNOR U3552 ( .A(n3854), .B(n1221), .Z(out[31]) );
  XNOR U3553 ( .A(n3856), .B(n2696), .Z(out[319]) );
  NOR U3554 ( .A(n3857), .B(n2695), .Z(n3856) );
  XNOR U3555 ( .A(n3858), .B(n2740), .Z(out[318]) );
  NOR U3556 ( .A(n3859), .B(n2739), .Z(n3858) );
  XNOR U3557 ( .A(n3860), .B(n2784), .Z(out[317]) );
  NOR U3558 ( .A(n3861), .B(n2783), .Z(n3860) );
  XNOR U3559 ( .A(n3862), .B(n2828), .Z(out[316]) );
  NOR U3560 ( .A(n3863), .B(n2827), .Z(n3862) );
  XNOR U3561 ( .A(n3864), .B(n2875), .Z(out[315]) );
  NOR U3562 ( .A(n3865), .B(n2874), .Z(n3864) );
  XNOR U3563 ( .A(n3866), .B(n2917), .Z(out[314]) );
  ANDN U3564 ( .B(n3867), .A(n2916), .Z(n3866) );
  XNOR U3565 ( .A(n3868), .B(n2957), .Z(out[313]) );
  ANDN U3566 ( .B(n3869), .A(n2956), .Z(n3868) );
  XNOR U3567 ( .A(n3870), .B(n2989), .Z(out[312]) );
  ANDN U3568 ( .B(n3871), .A(n2988), .Z(n3870) );
  XNOR U3569 ( .A(n3872), .B(n3021), .Z(out[311]) );
  NOR U3570 ( .A(n3873), .B(n3020), .Z(n3872) );
  XNOR U3571 ( .A(n3874), .B(n3050), .Z(out[310]) );
  ANDN U3572 ( .B(n3875), .A(n3049), .Z(n3874) );
  XNOR U3573 ( .A(n3876), .B(n1263), .Z(out[30]) );
  AND U3574 ( .A(n3877), .B(n3878), .Z(n3876) );
  XNOR U3575 ( .A(n3879), .B(n3081), .Z(out[309]) );
  ANDN U3576 ( .B(n3880), .A(n3080), .Z(n3879) );
  XNOR U3577 ( .A(n3881), .B(n3109), .Z(out[308]) );
  ANDN U3578 ( .B(n3882), .A(n3108), .Z(n3881) );
  XNOR U3579 ( .A(n3883), .B(n3133), .Z(out[307]) );
  ANDN U3580 ( .B(n3884), .A(n3132), .Z(n3883) );
  XNOR U3581 ( .A(n3885), .B(n3161), .Z(out[306]) );
  ANDN U3582 ( .B(n3886), .A(n3160), .Z(n3885) );
  XNOR U3583 ( .A(n3887), .B(n3202), .Z(out[305]) );
  ANDN U3584 ( .B(n3888), .A(n3201), .Z(n3887) );
  XNOR U3585 ( .A(n3889), .B(n3236), .Z(out[304]) );
  ANDN U3586 ( .B(n3890), .A(n3235), .Z(n3889) );
  XNOR U3587 ( .A(n3891), .B(n3270), .Z(out[303]) );
  AND U3588 ( .A(n3892), .B(n3893), .Z(n3891) );
  XNOR U3589 ( .A(n3894), .B(n3307), .Z(out[302]) );
  AND U3590 ( .A(n3895), .B(n3896), .Z(n3894) );
  XNOR U3591 ( .A(n3897), .B(n3349), .Z(out[301]) );
  XNOR U3592 ( .A(n3899), .B(n3391), .Z(out[300]) );
  XOR U3593 ( .A(n3901), .B(n2473), .Z(out[2]) );
  AND U3594 ( .A(n3902), .B(n3903), .Z(n3901) );
  XNOR U3595 ( .A(n3904), .B(n1304), .Z(out[29]) );
  AND U3596 ( .A(n3905), .B(n3906), .Z(n3904) );
  XNOR U3597 ( .A(n3907), .B(n3420), .Z(out[299]) );
  NOR U3598 ( .A(n3908), .B(n3419), .Z(n3907) );
  XNOR U3599 ( .A(n3909), .B(n3444), .Z(out[298]) );
  ANDN U3600 ( .B(n3910), .A(n3443), .Z(n3909) );
  XNOR U3601 ( .A(n3911), .B(n3468), .Z(out[297]) );
  NOR U3602 ( .A(n3912), .B(n3467), .Z(n3911) );
  XOR U3603 ( .A(n3913), .B(n3498), .Z(out[296]) );
  NOR U3604 ( .A(n3914), .B(n3497), .Z(n3913) );
  XOR U3605 ( .A(n3915), .B(n3530), .Z(out[295]) );
  NOR U3606 ( .A(n3916), .B(n3529), .Z(n3915) );
  XOR U3607 ( .A(n3917), .B(n3562), .Z(out[294]) );
  ANDN U3608 ( .B(n3918), .A(n3561), .Z(n3917) );
  XOR U3609 ( .A(n3919), .B(n3596), .Z(out[293]) );
  ANDN U3610 ( .B(n3920), .A(n3595), .Z(n3919) );
  XOR U3611 ( .A(n3921), .B(n3640), .Z(out[292]) );
  ANDN U3612 ( .B(n3922), .A(n3639), .Z(n3921) );
  XOR U3613 ( .A(n3923), .B(n1046), .Z(out[291]) );
  XOR U3614 ( .A(n2371), .B(n3924), .Z(n1046) );
  ANDN U3615 ( .B(n3925), .A(n3683), .Z(n3923) );
  XOR U3616 ( .A(n3926), .B(n1090), .Z(out[290]) );
  XOR U3617 ( .A(n2380), .B(n3927), .Z(n1090) );
  ANDN U3618 ( .B(n3928), .A(n3726), .Z(n3926) );
  XNOR U3619 ( .A(n3929), .B(n1350), .Z(out[28]) );
  ANDN U3620 ( .B(n3930), .A(n1349), .Z(n3929) );
  XOR U3621 ( .A(n3931), .B(n1133), .Z(out[289]) );
  IV U3622 ( .A(n3770), .Z(n1133) );
  XNOR U3623 ( .A(n2387), .B(n3932), .Z(n3770) );
  ANDN U3624 ( .B(n3933), .A(n3769), .Z(n3931) );
  XOR U3625 ( .A(n3934), .B(n1178), .Z(out[288]) );
  XOR U3626 ( .A(n2392), .B(n3935), .Z(n1178) );
  ANDN U3627 ( .B(n3936), .A(n3813), .Z(n3934) );
  XOR U3628 ( .A(n3937), .B(n1222), .Z(out[287]) );
  XOR U3629 ( .A(n2405), .B(n3938), .Z(n1222) );
  NOR U3630 ( .A(n3939), .B(n3855), .Z(n3937) );
  XOR U3631 ( .A(n3940), .B(n1264), .Z(out[286]) );
  IV U3632 ( .A(n3878), .Z(n1264) );
  XNOR U3633 ( .A(n3941), .B(n2411), .Z(n3878) );
  NOR U3634 ( .A(n3942), .B(n3877), .Z(n3940) );
  XOR U3635 ( .A(n3943), .B(n1305), .Z(out[285]) );
  IV U3636 ( .A(n3906), .Z(n1305) );
  XNOR U3637 ( .A(n3944), .B(n2418), .Z(n3906) );
  NOR U3638 ( .A(n3945), .B(n3905), .Z(n3943) );
  XOR U3639 ( .A(n3946), .B(n1349), .Z(out[284]) );
  XOR U3640 ( .A(n2424), .B(n3947), .Z(n1349) );
  ANDN U3641 ( .B(n3948), .A(n3930), .Z(n3946) );
  XOR U3642 ( .A(n3949), .B(n1393), .Z(out[283]) );
  XOR U3643 ( .A(n3952), .B(n1437), .Z(out[282]) );
  XOR U3644 ( .A(n3955), .B(n1485), .Z(out[281]) );
  ANDN U3645 ( .B(n3956), .A(n3957), .Z(n3955) );
  XOR U3646 ( .A(n3958), .B(n1517), .Z(out[280]) );
  ANDN U3647 ( .B(n3959), .A(n3960), .Z(n3958) );
  XNOR U3648 ( .A(n3961), .B(n1394), .Z(out[27]) );
  ANDN U3649 ( .B(n3951), .A(n1393), .Z(n3961) );
  XOR U3650 ( .A(n2431), .B(n3962), .Z(n1393) );
  XOR U3651 ( .A(n3963), .B(n1541), .Z(out[279]) );
  ANDN U3652 ( .B(n3964), .A(n3965), .Z(n3963) );
  XOR U3653 ( .A(n3966), .B(n1566), .Z(out[278]) );
  ANDN U3654 ( .B(n3967), .A(n3968), .Z(n3966) );
  XOR U3655 ( .A(n3969), .B(n1590), .Z(out[277]) );
  ANDN U3656 ( .B(n3970), .A(n3971), .Z(n3969) );
  XOR U3657 ( .A(n3972), .B(n1614), .Z(out[276]) );
  AND U3658 ( .A(n3973), .B(n3974), .Z(n3972) );
  XOR U3659 ( .A(n3975), .B(n1638), .Z(out[275]) );
  AND U3660 ( .A(n3976), .B(n3977), .Z(n3975) );
  XOR U3661 ( .A(n3978), .B(n1667), .Z(out[274]) );
  ANDN U3662 ( .B(n3979), .A(n3980), .Z(n3978) );
  XNOR U3663 ( .A(n3981), .B(n1720), .Z(out[273]) );
  AND U3664 ( .A(n3982), .B(n3983), .Z(n3981) );
  XOR U3665 ( .A(n3984), .B(n1772), .Z(out[272]) );
  IV U3666 ( .A(n3985), .Z(n1772) );
  ANDN U3667 ( .B(n3986), .A(n3987), .Z(n3984) );
  XOR U3668 ( .A(n3988), .B(n1820), .Z(out[271]) );
  ANDN U3669 ( .B(n3989), .A(n3990), .Z(n3988) );
  XOR U3670 ( .A(n3991), .B(n1865), .Z(out[270]) );
  ANDN U3671 ( .B(n3992), .A(n3993), .Z(n3991) );
  XNOR U3672 ( .A(n3994), .B(n1438), .Z(out[26]) );
  ANDN U3673 ( .B(n3954), .A(n1437), .Z(n3994) );
  XOR U3674 ( .A(n2440), .B(n3995), .Z(n1437) );
  XOR U3675 ( .A(n3996), .B(n1911), .Z(out[269]) );
  ANDN U3676 ( .B(n3997), .A(n3998), .Z(n3996) );
  XOR U3677 ( .A(n3999), .B(n1962), .Z(out[268]) );
  ANDN U3678 ( .B(n4000), .A(n4001), .Z(n3999) );
  XOR U3679 ( .A(n4002), .B(n2001), .Z(out[267]) );
  ANDN U3680 ( .B(n4003), .A(n4004), .Z(n4002) );
  XOR U3681 ( .A(n4005), .B(n2044), .Z(out[266]) );
  ANDN U3682 ( .B(n4006), .A(n4007), .Z(n4005) );
  XOR U3683 ( .A(n4008), .B(n1042), .Z(out[265]) );
  XOR U3684 ( .A(n2565), .B(n4009), .Z(n1042) );
  XOR U3685 ( .A(n4011), .B(n1482), .Z(out[264]) );
  XNOR U3686 ( .A(n4012), .B(n2573), .Z(n1482) );
  AND U3687 ( .A(n1481), .B(n4013), .Z(n4011) );
  IV U3688 ( .A(n4014), .Z(n1481) );
  XOR U3689 ( .A(n4015), .B(n1817), .Z(out[263]) );
  XNOR U3690 ( .A(n4016), .B(n2580), .Z(n1817) );
  AND U3691 ( .A(n4017), .B(n1816), .Z(n4015) );
  IV U3692 ( .A(n4018), .Z(n1816) );
  XOR U3693 ( .A(n4019), .B(n2198), .Z(out[262]) );
  IV U3694 ( .A(n2247), .Z(n2198) );
  XOR U3695 ( .A(n4020), .B(n2587), .Z(n2247) );
  XOR U3696 ( .A(n4022), .B(n2250), .Z(out[261]) );
  IV U3697 ( .A(n2871), .Z(n2250) );
  XOR U3698 ( .A(n4023), .B(n2594), .Z(n2871) );
  XOR U3699 ( .A(n4025), .B(n2325), .Z(out[260]) );
  IV U3700 ( .A(n3198), .Z(n2325) );
  XOR U3701 ( .A(n4026), .B(n2601), .Z(n3198) );
  XNOR U3702 ( .A(n4028), .B(n1486), .Z(out[25]) );
  ANDN U3703 ( .B(n3957), .A(n1485), .Z(n4028) );
  XOR U3704 ( .A(n2447), .B(n4029), .Z(n1485) );
  XOR U3705 ( .A(n4030), .B(n2398), .Z(out[259]) );
  IV U3706 ( .A(n3526), .Z(n2398) );
  XOR U3707 ( .A(n4031), .B(n2608), .Z(n3526) );
  XOR U3708 ( .A(n4033), .B(n2472), .Z(out[258]) );
  IV U3709 ( .A(n3903), .Z(n2472) );
  XOR U3710 ( .A(n4034), .B(n2615), .Z(n3903) );
  ANDN U3711 ( .B(n4035), .A(n3902), .Z(n4033) );
  XOR U3712 ( .A(n4036), .B(n2546), .Z(out[257]) );
  IV U3713 ( .A(n4037), .Z(n2546) );
  XOR U3714 ( .A(n4040), .B(n2620), .Z(out[256]) );
  IV U3715 ( .A(n4041), .Z(n2620) );
  XOR U3716 ( .A(n4044), .B(n2695), .Z(out[255]) );
  XOR U3717 ( .A(n1807), .B(n4045), .Z(n2695) );
  AND U3718 ( .A(n3857), .B(n4046), .Z(n4044) );
  XOR U3719 ( .A(n4047), .B(n2739), .Z(out[254]) );
  XOR U3720 ( .A(n1811), .B(n4048), .Z(n2739) );
  AND U3721 ( .A(n3859), .B(n4049), .Z(n4047) );
  XOR U3722 ( .A(n4050), .B(n2783), .Z(out[253]) );
  XOR U3723 ( .A(n1823), .B(n4051), .Z(n2783) );
  AND U3724 ( .A(n3861), .B(n4052), .Z(n4050) );
  XOR U3725 ( .A(n4053), .B(n2827), .Z(out[252]) );
  XOR U3726 ( .A(n1827), .B(n4054), .Z(n2827) );
  AND U3727 ( .A(n3863), .B(n4055), .Z(n4053) );
  XOR U3728 ( .A(n4056), .B(n2874), .Z(out[251]) );
  XOR U3729 ( .A(n1831), .B(n4057), .Z(n2874) );
  AND U3730 ( .A(n3865), .B(n4058), .Z(n4056) );
  XOR U3731 ( .A(n4059), .B(n2916), .Z(out[250]) );
  XOR U3732 ( .A(n1835), .B(n4060), .Z(n2916) );
  ANDN U3733 ( .B(n4061), .A(n3867), .Z(n4059) );
  XNOR U3734 ( .A(n4062), .B(n1518), .Z(out[24]) );
  ANDN U3735 ( .B(n3960), .A(n1517), .Z(n4062) );
  XOR U3736 ( .A(n2452), .B(n4063), .Z(n1517) );
  XOR U3737 ( .A(n4064), .B(n2956), .Z(out[249]) );
  XOR U3738 ( .A(n1839), .B(n4065), .Z(n2956) );
  ANDN U3739 ( .B(n4066), .A(n3869), .Z(n4064) );
  XOR U3740 ( .A(n4067), .B(n2988), .Z(out[248]) );
  XOR U3741 ( .A(n1843), .B(n4068), .Z(n2988) );
  ANDN U3742 ( .B(n4069), .A(n3871), .Z(n4067) );
  XOR U3743 ( .A(n4070), .B(n3020), .Z(out[247]) );
  XOR U3744 ( .A(n1847), .B(n4071), .Z(n3020) );
  AND U3745 ( .A(n3873), .B(n4072), .Z(n4070) );
  XOR U3746 ( .A(n4073), .B(n3049), .Z(out[246]) );
  XOR U3747 ( .A(n1852), .B(n4074), .Z(n3049) );
  NOR U3748 ( .A(n4075), .B(n3875), .Z(n4073) );
  XOR U3749 ( .A(n4076), .B(n3080), .Z(out[245]) );
  XOR U3750 ( .A(n1856), .B(n4077), .Z(n3080) );
  NOR U3751 ( .A(n4078), .B(n3880), .Z(n4076) );
  XOR U3752 ( .A(n4079), .B(n3108), .Z(out[244]) );
  XOR U3753 ( .A(n1860), .B(n4080), .Z(n3108) );
  AND U3754 ( .A(n4081), .B(n4082), .Z(n4079) );
  XOR U3755 ( .A(n4083), .B(n3132), .Z(out[243]) );
  XOR U3756 ( .A(n1868), .B(n4084), .Z(n3132) );
  AND U3757 ( .A(n4085), .B(n4086), .Z(n4083) );
  XOR U3758 ( .A(n4087), .B(n3160), .Z(out[242]) );
  XOR U3759 ( .A(n1872), .B(n4088), .Z(n3160) );
  AND U3760 ( .A(n4089), .B(n4090), .Z(n4087) );
  XOR U3761 ( .A(n4091), .B(n3201), .Z(out[241]) );
  XOR U3762 ( .A(n1876), .B(n4092), .Z(n3201) );
  ANDN U3763 ( .B(n4093), .A(n3888), .Z(n4091) );
  XOR U3764 ( .A(n4094), .B(n3235), .Z(out[240]) );
  XNOR U3765 ( .A(n3642), .B(n4095), .Z(n3235) );
  ANDN U3766 ( .B(n4096), .A(n3890), .Z(n4094) );
  XNOR U3767 ( .A(n4097), .B(n1542), .Z(out[23]) );
  ANDN U3768 ( .B(n3965), .A(n1541), .Z(n4097) );
  XOR U3769 ( .A(n2459), .B(n4098), .Z(n1541) );
  XOR U3770 ( .A(n4099), .B(n3271), .Z(out[239]) );
  IV U3771 ( .A(n3893), .Z(n3271) );
  XOR U3772 ( .A(n1885), .B(n4100), .Z(n3893) );
  ANDN U3773 ( .B(n4101), .A(n3892), .Z(n4099) );
  XOR U3774 ( .A(n4102), .B(n3308), .Z(out[238]) );
  IV U3775 ( .A(n3896), .Z(n3308) );
  XOR U3776 ( .A(n1889), .B(n4103), .Z(n3896) );
  NOR U3777 ( .A(n4104), .B(n3895), .Z(n4102) );
  XOR U3778 ( .A(n4105), .B(n3350), .Z(out[237]) );
  XOR U3779 ( .A(n1893), .B(n4106), .Z(n3350) );
  NOR U3780 ( .A(n4107), .B(n3898), .Z(n4105) );
  XOR U3781 ( .A(n4108), .B(n3392), .Z(out[236]) );
  XOR U3782 ( .A(n1897), .B(n4109), .Z(n3392) );
  ANDN U3783 ( .B(n4110), .A(n3900), .Z(n4108) );
  XOR U3784 ( .A(n4111), .B(n3419), .Z(out[235]) );
  XOR U3785 ( .A(n1901), .B(n4112), .Z(n3419) );
  AND U3786 ( .A(n3908), .B(n4113), .Z(n4111) );
  XOR U3787 ( .A(n4114), .B(n3443), .Z(out[234]) );
  XOR U3788 ( .A(n1906), .B(n4115), .Z(n3443) );
  ANDN U3789 ( .B(n4116), .A(n3910), .Z(n4114) );
  XOR U3790 ( .A(n4117), .B(n3467), .Z(out[233]) );
  XOR U3791 ( .A(n1914), .B(n4118), .Z(n3467) );
  AND U3792 ( .A(n3912), .B(n4119), .Z(n4117) );
  XOR U3793 ( .A(n4120), .B(n3497), .Z(out[232]) );
  XOR U3794 ( .A(n1919), .B(n4121), .Z(n3497) );
  AND U3795 ( .A(n3914), .B(n4122), .Z(n4120) );
  XOR U3796 ( .A(n4123), .B(n3529), .Z(out[231]) );
  XOR U3797 ( .A(n1923), .B(n4124), .Z(n3529) );
  AND U3798 ( .A(n3916), .B(n4125), .Z(n4123) );
  XOR U3799 ( .A(n4126), .B(n3561), .Z(out[230]) );
  XOR U3800 ( .A(n1927), .B(n4127), .Z(n3561) );
  ANDN U3801 ( .B(n4128), .A(n3918), .Z(n4126) );
  XNOR U3802 ( .A(n4129), .B(n1567), .Z(out[22]) );
  ANDN U3803 ( .B(n3968), .A(n1566), .Z(n4129) );
  XOR U3804 ( .A(n2466), .B(n4130), .Z(n1566) );
  XOR U3805 ( .A(n4131), .B(n3595), .Z(out[229]) );
  XOR U3806 ( .A(n1931), .B(n4132), .Z(n3595) );
  ANDN U3807 ( .B(n4133), .A(n3920), .Z(n4131) );
  XOR U3808 ( .A(n4134), .B(n3639), .Z(out[228]) );
  XOR U3809 ( .A(n1936), .B(n4135), .Z(n3639) );
  ANDN U3810 ( .B(n4136), .A(n3922), .Z(n4134) );
  XOR U3811 ( .A(n4137), .B(n3683), .Z(out[227]) );
  XOR U3812 ( .A(n1941), .B(n4138), .Z(n3683) );
  NOR U3813 ( .A(n1044), .B(n3925), .Z(n4137) );
  XOR U3814 ( .A(n4139), .B(n3726), .Z(out[226]) );
  XOR U3815 ( .A(n1946), .B(n4140), .Z(n3726) );
  NOR U3816 ( .A(n1088), .B(n3928), .Z(n4139) );
  XOR U3817 ( .A(n4141), .B(n3769), .Z(out[225]) );
  XNOR U3818 ( .A(n1951), .B(n4142), .Z(n3769) );
  ANDN U3819 ( .B(n1132), .A(n3933), .Z(n4141) );
  XOR U3820 ( .A(n4143), .B(n3813), .Z(out[224]) );
  XNOR U3821 ( .A(n4144), .B(n1957), .Z(n3813) );
  ANDN U3822 ( .B(n1176), .A(n3936), .Z(n4143) );
  IV U3823 ( .A(n4145), .Z(n1176) );
  XOR U3824 ( .A(n4146), .B(n3855), .Z(out[223]) );
  XNOR U3825 ( .A(n4147), .B(n1966), .Z(n3855) );
  AND U3826 ( .A(n3939), .B(n1220), .Z(n4146) );
  IV U3827 ( .A(n4148), .Z(n1220) );
  XOR U3828 ( .A(n4149), .B(n3877), .Z(out[222]) );
  XNOR U3829 ( .A(n4150), .B(n1971), .Z(n3877) );
  AND U3830 ( .A(n3942), .B(n1262), .Z(n4149) );
  IV U3831 ( .A(n4151), .Z(n1262) );
  XOR U3832 ( .A(n4152), .B(n3905), .Z(out[221]) );
  XNOR U3833 ( .A(n4153), .B(n1658), .Z(n3905) );
  AND U3834 ( .A(n3945), .B(n1303), .Z(n4152) );
  IV U3835 ( .A(n4154), .Z(n1303) );
  XOR U3836 ( .A(n4155), .B(n3930), .Z(out[220]) );
  XNOR U3837 ( .A(n4156), .B(n1663), .Z(n3930) );
  XNOR U3838 ( .A(n4157), .B(n1591), .Z(out[21]) );
  ANDN U3839 ( .B(n3971), .A(n1590), .Z(n4157) );
  XOR U3840 ( .A(n2477), .B(n4158), .Z(n1590) );
  XOR U3841 ( .A(n4159), .B(n3951), .Z(out[219]) );
  XNOR U3842 ( .A(n4160), .B(n1671), .Z(n3951) );
  ANDN U3843 ( .B(n1392), .A(n3950), .Z(n4159) );
  IV U3844 ( .A(n4161), .Z(n1392) );
  XOR U3845 ( .A(n4162), .B(n3954), .Z(out[218]) );
  XNOR U3846 ( .A(n4163), .B(n1675), .Z(n3954) );
  ANDN U3847 ( .B(n1436), .A(n3953), .Z(n4162) );
  IV U3848 ( .A(n4164), .Z(n1436) );
  XOR U3849 ( .A(n4165), .B(n3957), .Z(out[217]) );
  XNOR U3850 ( .A(n4166), .B(n1680), .Z(n3957) );
  ANDN U3851 ( .B(n1484), .A(n3956), .Z(n4165) );
  IV U3852 ( .A(n4167), .Z(n1484) );
  XOR U3853 ( .A(n4168), .B(n3960), .Z(out[216]) );
  XOR U3854 ( .A(n4169), .B(n1685), .Z(n3960) );
  ANDN U3855 ( .B(n1516), .A(n3959), .Z(n4168) );
  IV U3856 ( .A(n4170), .Z(n1516) );
  XOR U3857 ( .A(n4171), .B(n3965), .Z(out[215]) );
  XNOR U3858 ( .A(n4172), .B(n1690), .Z(n3965) );
  ANDN U3859 ( .B(n1540), .A(n3964), .Z(n4171) );
  IV U3860 ( .A(n4173), .Z(n1540) );
  XOR U3861 ( .A(n4174), .B(n3968), .Z(out[214]) );
  XNOR U3862 ( .A(n4175), .B(n1695), .Z(n3968) );
  ANDN U3863 ( .B(n1565), .A(n3967), .Z(n4174) );
  IV U3864 ( .A(n4176), .Z(n1565) );
  XOR U3865 ( .A(n4177), .B(n3971), .Z(out[213]) );
  XOR U3866 ( .A(n4178), .B(n1700), .Z(n3971) );
  ANDN U3867 ( .B(n1589), .A(n3970), .Z(n4177) );
  IV U3868 ( .A(n4179), .Z(n1589) );
  XNOR U3869 ( .A(n4180), .B(n3974), .Z(out[212]) );
  ANDN U3870 ( .B(n1613), .A(n3973), .Z(n4180) );
  IV U3871 ( .A(n4181), .Z(n1613) );
  XNOR U3872 ( .A(n4182), .B(n3977), .Z(out[211]) );
  NOR U3873 ( .A(n1637), .B(n3976), .Z(n4182) );
  XNOR U3874 ( .A(n4183), .B(n3979), .Z(out[210]) );
  ANDN U3875 ( .B(n3980), .A(n1666), .Z(n4183) );
  XNOR U3876 ( .A(n4184), .B(n1615), .Z(out[20]) );
  NOR U3877 ( .A(n3974), .B(n1614), .Z(n4184) );
  XOR U3878 ( .A(n2484), .B(n4185), .Z(n1614) );
  XNOR U3879 ( .A(n4186), .B(n1705), .Z(n3974) );
  XNOR U3880 ( .A(n4187), .B(n3982), .Z(out[209]) );
  XNOR U3881 ( .A(n4188), .B(n3986), .Z(out[208]) );
  ANDN U3882 ( .B(n3987), .A(n1770), .Z(n4188) );
  XNOR U3883 ( .A(n4189), .B(n3989), .Z(out[207]) );
  ANDN U3884 ( .B(n3990), .A(n1819), .Z(n4189) );
  XNOR U3885 ( .A(n4190), .B(n3992), .Z(out[206]) );
  ANDN U3886 ( .B(n3993), .A(n1864), .Z(n4190) );
  XNOR U3887 ( .A(n4191), .B(n3997), .Z(out[205]) );
  ANDN U3888 ( .B(n3998), .A(n1910), .Z(n4191) );
  XNOR U3889 ( .A(n4192), .B(n4000), .Z(out[204]) );
  ANDN U3890 ( .B(n4001), .A(n1961), .Z(n4192) );
  XNOR U3891 ( .A(n4193), .B(n4003), .Z(out[203]) );
  ANDN U3892 ( .B(n4004), .A(n2000), .Z(n4193) );
  XNOR U3893 ( .A(n4194), .B(n4006), .Z(out[202]) );
  ANDN U3894 ( .B(n4007), .A(n2043), .Z(n4194) );
  XOR U3895 ( .A(n4195), .B(n1041), .Z(out[201]) );
  XOR U3896 ( .A(n1761), .B(n4196), .Z(n1041) );
  ANDN U3897 ( .B(n4197), .A(n2083), .Z(n4195) );
  XOR U3898 ( .A(n4198), .B(n4014), .Z(out[200]) );
  XOR U3899 ( .A(n4199), .B(n1766), .Z(n4014) );
  ANDN U3900 ( .B(n4200), .A(n2122), .Z(n4198) );
  XOR U3901 ( .A(n4201), .B(n2547), .Z(out[1]) );
  AND U3902 ( .A(n4039), .B(n4037), .Z(n4201) );
  XOR U3903 ( .A(n4202), .B(n2627), .Z(n4037) );
  XNOR U3904 ( .A(n4203), .B(n1639), .Z(out[19]) );
  NOR U3905 ( .A(n3977), .B(n1638), .Z(n4203) );
  XOR U3906 ( .A(n2493), .B(n4204), .Z(n1638) );
  XNOR U3907 ( .A(n4205), .B(n1710), .Z(n3977) );
  XOR U3908 ( .A(n4206), .B(n4018), .Z(out[199]) );
  XOR U3909 ( .A(n4207), .B(n1775), .Z(n4018) );
  NOR U3910 ( .A(n2161), .B(n4017), .Z(n4206) );
  XOR U3911 ( .A(n4208), .B(n2246), .Z(out[198]) );
  XOR U3912 ( .A(n4209), .B(n1780), .Z(n2246) );
  XOR U3913 ( .A(n4210), .B(n2870), .Z(out[197]) );
  XOR U3914 ( .A(n4211), .B(n1784), .Z(n2870) );
  IV U3915 ( .A(n4212), .Z(n2249) );
  XOR U3916 ( .A(n4213), .B(n3197), .Z(out[196]) );
  XOR U3917 ( .A(n4214), .B(n1788), .Z(n3197) );
  XOR U3918 ( .A(n4215), .B(n3525), .Z(out[195]) );
  XOR U3919 ( .A(n4216), .B(n1792), .Z(n3525) );
  AND U3920 ( .A(n2397), .B(n4217), .Z(n4215) );
  IV U3921 ( .A(n4218), .Z(n2397) );
  XOR U3922 ( .A(n4219), .B(n3902), .Z(out[194]) );
  XNOR U3923 ( .A(n1795), .B(n4220), .Z(n3902) );
  AND U3924 ( .A(n2471), .B(n4221), .Z(n4219) );
  XOR U3925 ( .A(n4222), .B(n4039), .Z(out[193]) );
  XOR U3926 ( .A(n4223), .B(n1800), .Z(n4039) );
  ANDN U3927 ( .B(n2545), .A(n4038), .Z(n4222) );
  XOR U3928 ( .A(n4224), .B(n4043), .Z(out[192]) );
  NOR U3929 ( .A(n2619), .B(n4042), .Z(n4224) );
  XNOR U3930 ( .A(n4225), .B(n3857), .Z(out[191]) );
  XOR U3931 ( .A(n4226), .B(n2098), .Z(n3857) );
  AND U3932 ( .A(n2694), .B(n4227), .Z(n4225) );
  XNOR U3933 ( .A(n4228), .B(n3859), .Z(out[190]) );
  XOR U3934 ( .A(n4229), .B(n2101), .Z(n3859) );
  AND U3935 ( .A(n2738), .B(n4230), .Z(n4228) );
  XNOR U3936 ( .A(n4231), .B(n1668), .Z(out[18]) );
  NOR U3937 ( .A(n3979), .B(n1667), .Z(n4231) );
  XOR U3938 ( .A(n2500), .B(n4232), .Z(n1667) );
  XNOR U3939 ( .A(n4233), .B(n1715), .Z(n3979) );
  XNOR U3940 ( .A(n4234), .B(n3861), .Z(out[189]) );
  XOR U3941 ( .A(n4235), .B(n2105), .Z(n3861) );
  AND U3942 ( .A(n2782), .B(n4236), .Z(n4234) );
  XNOR U3943 ( .A(n4237), .B(n3863), .Z(out[188]) );
  XOR U3944 ( .A(n4238), .B(n2108), .Z(n3863) );
  XNOR U3945 ( .A(n4239), .B(n3865), .Z(out[187]) );
  XOR U3946 ( .A(n4240), .B(n2111), .Z(n3865) );
  XOR U3947 ( .A(n4241), .B(n3867), .Z(out[186]) );
  XOR U3948 ( .A(n2114), .B(n4242), .Z(n3867) );
  ANDN U3949 ( .B(n4243), .A(n2915), .Z(n4241) );
  XOR U3950 ( .A(n4244), .B(n3869), .Z(out[185]) );
  XNOR U3951 ( .A(n2118), .B(n4245), .Z(n3869) );
  XOR U3952 ( .A(n4246), .B(n3871), .Z(out[184]) );
  XOR U3953 ( .A(n4247), .B(n2125), .Z(n3871) );
  XNOR U3954 ( .A(n4248), .B(n3873), .Z(out[183]) );
  XNOR U3955 ( .A(n2127), .B(n4249), .Z(n3873) );
  XOR U3956 ( .A(n4250), .B(n3875), .Z(out[182]) );
  XOR U3957 ( .A(n2131), .B(n4251), .Z(n3875) );
  ANDN U3958 ( .B(n4075), .A(n3048), .Z(n4250) );
  XOR U3959 ( .A(n4252), .B(n3880), .Z(out[181]) );
  XOR U3960 ( .A(n2135), .B(n4253), .Z(n3880) );
  ANDN U3961 ( .B(n4078), .A(n3079), .Z(n4252) );
  XOR U3962 ( .A(n4254), .B(n3882), .Z(out[180]) );
  IV U3963 ( .A(n4082), .Z(n3882) );
  XNOR U3964 ( .A(n2139), .B(n4255), .Z(n4082) );
  NOR U3965 ( .A(n4081), .B(n3107), .Z(n4254) );
  XOR U3966 ( .A(n4256), .B(n1721), .Z(out[17]) );
  ANDN U3967 ( .B(n1720), .A(n3982), .Z(n4256) );
  XOR U3968 ( .A(n4257), .B(n1724), .Z(n3982) );
  XNOR U3969 ( .A(n2505), .B(n4258), .Z(n1720) );
  XOR U3970 ( .A(n4259), .B(n3884), .Z(out[179]) );
  IV U3971 ( .A(n4086), .Z(n3884) );
  XNOR U3972 ( .A(n2143), .B(n4260), .Z(n4086) );
  NOR U3973 ( .A(n3131), .B(n4085), .Z(n4259) );
  XOR U3974 ( .A(n4261), .B(n3886), .Z(out[178]) );
  IV U3975 ( .A(n4090), .Z(n3886) );
  XOR U3976 ( .A(n2147), .B(n4262), .Z(n4090) );
  NOR U3977 ( .A(n3159), .B(n4089), .Z(n4261) );
  XOR U3978 ( .A(n4263), .B(n3888), .Z(out[177]) );
  XNOR U3979 ( .A(n4264), .B(n2152), .Z(n3888) );
  ANDN U3980 ( .B(n4265), .A(n3200), .Z(n4263) );
  XOR U3981 ( .A(n4266), .B(n3890), .Z(out[176]) );
  XNOR U3982 ( .A(n4267), .B(n2155), .Z(n3890) );
  ANDN U3983 ( .B(n4268), .A(n3234), .Z(n4266) );
  XOR U3984 ( .A(n4269), .B(n3892), .Z(out[175]) );
  XNOR U3985 ( .A(n4270), .B(n2159), .Z(n3892) );
  ANDN U3986 ( .B(n4271), .A(n3269), .Z(n4269) );
  XOR U3987 ( .A(n4272), .B(n3895), .Z(out[174]) );
  XNOR U3988 ( .A(n4273), .B(n2164), .Z(n3895) );
  AND U3989 ( .A(n4104), .B(n3306), .Z(n4272) );
  IV U3990 ( .A(n4274), .Z(n3306) );
  XOR U3991 ( .A(n4275), .B(n3898), .Z(out[173]) );
  XNOR U3992 ( .A(n4276), .B(n2168), .Z(n3898) );
  AND U3993 ( .A(n4107), .B(n3348), .Z(n4275) );
  IV U3994 ( .A(n4277), .Z(n3348) );
  XOR U3995 ( .A(n4278), .B(n3900), .Z(out[172]) );
  XOR U3996 ( .A(n4279), .B(n2172), .Z(n3900) );
  ANDN U3997 ( .B(n4280), .A(n3390), .Z(n4278) );
  XNOR U3998 ( .A(n4281), .B(n3908), .Z(out[171]) );
  XOR U3999 ( .A(n4282), .B(n2175), .Z(n3908) );
  ANDN U4000 ( .B(n4283), .A(n3418), .Z(n4281) );
  XOR U4001 ( .A(n4284), .B(n3910), .Z(out[170]) );
  XOR U4002 ( .A(n4285), .B(n2178), .Z(n3910) );
  ANDN U4003 ( .B(n4286), .A(n3442), .Z(n4284) );
  XNOR U4004 ( .A(n4287), .B(n1771), .Z(out[16]) );
  ANDN U4005 ( .B(n3985), .A(n3986), .Z(n4287) );
  XOR U4006 ( .A(n4288), .B(n1728), .Z(n3986) );
  XNOR U4007 ( .A(n4289), .B(n2513), .Z(n3985) );
  XNOR U4008 ( .A(n4290), .B(n3912), .Z(out[169]) );
  XNOR U4009 ( .A(n4291), .B(n2181), .Z(n3912) );
  ANDN U4010 ( .B(n4292), .A(n3466), .Z(n4290) );
  XNOR U4011 ( .A(n4293), .B(n3914), .Z(out[168]) );
  XNOR U4012 ( .A(n4294), .B(n2184), .Z(n3914) );
  IV U4013 ( .A(n4295), .Z(n2184) );
  ANDN U4014 ( .B(n4296), .A(n3496), .Z(n4293) );
  XNOR U4015 ( .A(n4297), .B(n3916), .Z(out[167]) );
  XNOR U4016 ( .A(n4298), .B(n2188), .Z(n3916) );
  ANDN U4017 ( .B(n4299), .A(n3528), .Z(n4297) );
  XOR U4018 ( .A(n4300), .B(n3918), .Z(out[166]) );
  XNOR U4019 ( .A(n4301), .B(n2191), .Z(n3918) );
  ANDN U4020 ( .B(n4302), .A(n3560), .Z(n4300) );
  XOR U4021 ( .A(n4303), .B(n3920), .Z(out[165]) );
  XOR U4022 ( .A(n4304), .B(n2194), .Z(n3920) );
  ANDN U4023 ( .B(n4305), .A(n3594), .Z(n4303) );
  XOR U4024 ( .A(n4306), .B(n3922), .Z(out[164]) );
  XOR U4025 ( .A(n4307), .B(n2201), .Z(n3922) );
  ANDN U4026 ( .B(n4308), .A(n3638), .Z(n4306) );
  XOR U4027 ( .A(n4309), .B(n3925), .Z(out[163]) );
  XOR U4028 ( .A(n4310), .B(n2204), .Z(n3925) );
  ANDN U4029 ( .B(n1044), .A(n1045), .Z(n4309) );
  XNOR U4030 ( .A(n2438), .B(n4311), .Z(n1045) );
  XNOR U4031 ( .A(n2598), .B(n4312), .Z(n1044) );
  XOR U4032 ( .A(n4313), .B(n3928), .Z(out[162]) );
  XOR U4033 ( .A(n4314), .B(n2207), .Z(n3928) );
  ANDN U4034 ( .B(n1088), .A(n1089), .Z(n4313) );
  XNOR U4035 ( .A(n2445), .B(n4315), .Z(n1089) );
  XNOR U4036 ( .A(n2605), .B(n4316), .Z(n1088) );
  XOR U4037 ( .A(n4317), .B(n3933), .Z(out[161]) );
  XOR U4038 ( .A(n4318), .B(n2210), .Z(n3933) );
  ANDN U4039 ( .B(n1134), .A(n1132), .Z(n4317) );
  XNOR U4040 ( .A(n4319), .B(n4320), .Z(n1132) );
  XOR U4041 ( .A(n4321), .B(n2455), .Z(n1134) );
  XOR U4042 ( .A(n4322), .B(n3936), .Z(out[160]) );
  XOR U4043 ( .A(n4323), .B(n2213), .Z(n3936) );
  ANDN U4044 ( .B(n4145), .A(n1177), .Z(n4322) );
  XNOR U4045 ( .A(n4324), .B(n2462), .Z(n1177) );
  XOR U4046 ( .A(n4325), .B(n2625), .Z(n4145) );
  XNOR U4047 ( .A(n4326), .B(n1821), .Z(out[15]) );
  NOR U4048 ( .A(n3989), .B(n1820), .Z(n4326) );
  XNOR U4049 ( .A(n2519), .B(n4327), .Z(n1820) );
  XOR U4050 ( .A(n4328), .B(n1732), .Z(n3989) );
  XNOR U4051 ( .A(n4329), .B(n3939), .Z(out[159]) );
  XNOR U4052 ( .A(n4330), .B(n2216), .Z(n3939) );
  ANDN U4053 ( .B(n4148), .A(n1221), .Z(n4329) );
  XOR U4054 ( .A(n4331), .B(n2469), .Z(n1221) );
  XOR U4055 ( .A(n4332), .B(n3742), .Z(n4148) );
  XOR U4056 ( .A(n4333), .B(n4334), .Z(out[1599]) );
  XOR U4057 ( .A(n4335), .B(n4336), .Z(n4334) );
  AND U4058 ( .A(n4337), .B(n4338), .Z(n4336) );
  AND U4059 ( .A(n4339), .B(n4340), .Z(n4338) );
  ANDN U4060 ( .B(n4341), .A(n4342), .Z(n4337) );
  ANDN U4061 ( .B(n4343), .A(n4344), .Z(n4341) );
  XOR U4062 ( .A(n4347), .B(n4348), .Z(out[1598]) );
  AND U4063 ( .A(n4349), .B(n4350), .Z(n4347) );
  XOR U4064 ( .A(n4351), .B(n4352), .Z(out[1597]) );
  AND U4065 ( .A(n4353), .B(n4354), .Z(n4351) );
  XOR U4066 ( .A(n4355), .B(n4356), .Z(out[1596]) );
  AND U4067 ( .A(n4357), .B(n4358), .Z(n4355) );
  XOR U4068 ( .A(n4359), .B(n4360), .Z(out[1595]) );
  AND U4069 ( .A(n4361), .B(n4362), .Z(n4359) );
  XOR U4070 ( .A(n4363), .B(n4364), .Z(out[1594]) );
  AND U4071 ( .A(n4365), .B(n4366), .Z(n4363) );
  XOR U4072 ( .A(n4367), .B(n4368), .Z(out[1593]) );
  AND U4073 ( .A(n4369), .B(n4370), .Z(n4367) );
  XOR U4074 ( .A(n4371), .B(n4372), .Z(out[1592]) );
  AND U4075 ( .A(n4373), .B(n4374), .Z(n4371) );
  XOR U4076 ( .A(n4375), .B(n4376), .Z(out[1591]) );
  AND U4077 ( .A(n4377), .B(n4378), .Z(n4375) );
  XOR U4078 ( .A(n4379), .B(n4380), .Z(out[1590]) );
  AND U4079 ( .A(n4381), .B(n4382), .Z(n4379) );
  XNOR U4080 ( .A(n4383), .B(n3942), .Z(out[158]) );
  XNOR U4081 ( .A(n4384), .B(n1976), .Z(n3942) );
  ANDN U4082 ( .B(n4151), .A(n1263), .Z(n4383) );
  XNOR U4083 ( .A(n4385), .B(n2480), .Z(n1263) );
  XOR U4084 ( .A(n4386), .B(n2639), .Z(n4151) );
  XOR U4085 ( .A(n4387), .B(n4388), .Z(out[1589]) );
  AND U4086 ( .A(n4389), .B(n4390), .Z(n4387) );
  XOR U4087 ( .A(n4391), .B(n4392), .Z(out[1588]) );
  AND U4088 ( .A(n4393), .B(n4394), .Z(n4391) );
  XOR U4089 ( .A(n4395), .B(n4396), .Z(out[1587]) );
  XOR U4090 ( .A(n4399), .B(n4400), .Z(out[1586]) );
  AND U4091 ( .A(n4401), .B(n4402), .Z(n4399) );
  XOR U4092 ( .A(n4403), .B(n4404), .Z(out[1585]) );
  AND U4093 ( .A(n4405), .B(n4406), .Z(n4403) );
  XOR U4094 ( .A(n4407), .B(n4408), .Z(out[1584]) );
  AND U4095 ( .A(n4409), .B(n4410), .Z(n4407) );
  XOR U4096 ( .A(n4411), .B(n4412), .Z(out[1583]) );
  ANDN U4097 ( .B(n4413), .A(n4414), .Z(n4411) );
  XOR U4098 ( .A(n4415), .B(n4416), .Z(out[1582]) );
  AND U4099 ( .A(n4417), .B(n4418), .Z(n4415) );
  XOR U4100 ( .A(n4419), .B(n4420), .Z(out[1581]) );
  ANDN U4101 ( .B(n4421), .A(n4422), .Z(n4419) );
  XOR U4102 ( .A(n4423), .B(n4424), .Z(out[1580]) );
  ANDN U4103 ( .B(n4425), .A(n4426), .Z(n4423) );
  XNOR U4104 ( .A(n4427), .B(n3945), .Z(out[157]) );
  XNOR U4105 ( .A(n4428), .B(n1979), .Z(n3945) );
  ANDN U4106 ( .B(n4154), .A(n1304), .Z(n4427) );
  XNOR U4107 ( .A(n4429), .B(n2487), .Z(n1304) );
  XOR U4108 ( .A(n4430), .B(n2646), .Z(n4154) );
  XOR U4109 ( .A(n4431), .B(n4432), .Z(out[1579]) );
  ANDN U4110 ( .B(n4433), .A(n4434), .Z(n4431) );
  XOR U4111 ( .A(n4435), .B(n4436), .Z(out[1578]) );
  AND U4112 ( .A(n4437), .B(n4438), .Z(n4435) );
  XOR U4113 ( .A(n4439), .B(n4440), .Z(out[1577]) );
  AND U4114 ( .A(n4441), .B(n4442), .Z(n4439) );
  XOR U4115 ( .A(n4443), .B(n4444), .Z(out[1576]) );
  AND U4116 ( .A(n4445), .B(n4446), .Z(n4443) );
  XOR U4117 ( .A(n4447), .B(n4448), .Z(out[1575]) );
  AND U4118 ( .A(n4449), .B(n4450), .Z(n4447) );
  XOR U4119 ( .A(n4451), .B(n4452), .Z(out[1574]) );
  AND U4120 ( .A(n4453), .B(n4454), .Z(n4451) );
  XOR U4121 ( .A(n4455), .B(n4456), .Z(out[1573]) );
  AND U4122 ( .A(n4457), .B(n4458), .Z(n4455) );
  XNOR U4123 ( .A(n4459), .B(n4460), .Z(out[1572]) );
  AND U4124 ( .A(n4461), .B(n4462), .Z(n4459) );
  XOR U4125 ( .A(n4463), .B(n4464), .Z(out[1571]) );
  AND U4126 ( .A(n4465), .B(n4466), .Z(n4463) );
  XOR U4127 ( .A(n4467), .B(n4468), .Z(out[1570]) );
  ANDN U4128 ( .B(n4469), .A(n4470), .Z(n4467) );
  XOR U4129 ( .A(n4471), .B(n3948), .Z(out[156]) );
  XOR U4130 ( .A(n4472), .B(n1982), .Z(n3948) );
  ANDN U4131 ( .B(n1348), .A(n1350), .Z(n4471) );
  XNOR U4132 ( .A(n4473), .B(n2492), .Z(n1350) );
  XOR U4133 ( .A(n4474), .B(n2653), .Z(n1348) );
  XNOR U4134 ( .A(n4475), .B(n4476), .Z(out[1569]) );
  ANDN U4135 ( .B(n4477), .A(n4478), .Z(n4475) );
  XNOR U4136 ( .A(n4479), .B(n4480), .Z(out[1568]) );
  AND U4137 ( .A(n4481), .B(n4482), .Z(n4479) );
  XOR U4138 ( .A(n4483), .B(n4484), .Z(out[1567]) );
  XOR U4139 ( .A(n4485), .B(n4486), .Z(n4484) );
  AND U4140 ( .A(n4487), .B(n4488), .Z(n4486) );
  AND U4141 ( .A(n4489), .B(n4490), .Z(n4488) );
  NOR U4142 ( .A(rc_i[5]), .B(rc_i[9]), .Z(n4489) );
  AND U4143 ( .A(n4491), .B(n4343), .Z(n4487) );
  AND U4144 ( .A(n4492), .B(n4493), .Z(n4485) );
  XNOR U4145 ( .A(n4494), .B(n4495), .Z(out[1566]) );
  AND U4146 ( .A(n4496), .B(n4497), .Z(n4494) );
  XNOR U4147 ( .A(n4498), .B(n4499), .Z(out[1565]) );
  AND U4148 ( .A(n4500), .B(n4501), .Z(n4498) );
  XOR U4149 ( .A(n4502), .B(n4503), .Z(out[1564]) );
  AND U4150 ( .A(n4504), .B(n4505), .Z(n4502) );
  XOR U4151 ( .A(n4506), .B(n4507), .Z(out[1563]) );
  AND U4152 ( .A(n4508), .B(n4509), .Z(n4506) );
  XOR U4153 ( .A(n4510), .B(n4511), .Z(out[1562]) );
  AND U4154 ( .A(n4512), .B(n4513), .Z(n4510) );
  XOR U4155 ( .A(n4514), .B(n4515), .Z(out[1561]) );
  XOR U4156 ( .A(n4518), .B(n4519), .Z(out[1560]) );
  XOR U4157 ( .A(n4522), .B(n3950), .Z(out[155]) );
  XOR U4158 ( .A(n4523), .B(n1985), .Z(n3950) );
  ANDN U4159 ( .B(n4161), .A(n1394), .Z(n4522) );
  XNOR U4160 ( .A(n4524), .B(n2499), .Z(n1394) );
  XOR U4161 ( .A(n4525), .B(n2660), .Z(n4161) );
  XOR U4162 ( .A(n4526), .B(n4527), .Z(out[1559]) );
  XOR U4163 ( .A(n4530), .B(n4531), .Z(out[1558]) );
  XNOR U4164 ( .A(n4534), .B(n4535), .Z(out[1557]) );
  XNOR U4165 ( .A(n4538), .B(n4539), .Z(out[1556]) );
  XNOR U4166 ( .A(n4542), .B(n4543), .Z(out[1555]) );
  XNOR U4167 ( .A(n4546), .B(n4547), .Z(out[1554]) );
  XOR U4168 ( .A(n4550), .B(n4551), .Z(out[1553]) );
  XNOR U4169 ( .A(n4554), .B(n4555), .Z(out[1552]) );
  XOR U4170 ( .A(n4558), .B(n4559), .Z(out[1551]) );
  XOR U4171 ( .A(n4560), .B(n4561), .Z(n4559) );
  AND U4172 ( .A(n4562), .B(n4563), .Z(n4561) );
  AND U4173 ( .A(n4564), .B(n4343), .Z(n4563) );
  ANDN U4174 ( .B(n4565), .A(n4344), .Z(n4562) );
  NAND U4175 ( .A(n4566), .B(n4491), .Z(n4344) );
  XNOR U4176 ( .A(n4569), .B(n4570), .Z(out[1550]) );
  XOR U4177 ( .A(n4573), .B(n3953), .Z(out[154]) );
  XOR U4178 ( .A(n4574), .B(n1988), .Z(n3953) );
  ANDN U4179 ( .B(n4164), .A(n1438), .Z(n4573) );
  XNOR U4180 ( .A(n4575), .B(n2508), .Z(n1438) );
  XOR U4181 ( .A(n4576), .B(n2667), .Z(n4164) );
  XNOR U4182 ( .A(n4577), .B(n4578), .Z(out[1549]) );
  XOR U4183 ( .A(n4581), .B(n4582), .Z(out[1548]) );
  XNOR U4184 ( .A(n4585), .B(n4586), .Z(out[1547]) );
  AND U4185 ( .A(n4587), .B(n4588), .Z(n4585) );
  XOR U4186 ( .A(n4589), .B(n4590), .Z(out[1546]) );
  XOR U4187 ( .A(n4593), .B(n4594), .Z(out[1545]) );
  XOR U4188 ( .A(n4597), .B(n4598), .Z(out[1544]) );
  XOR U4189 ( .A(n4601), .B(n4602), .Z(out[1543]) );
  XOR U4190 ( .A(n4603), .B(n4604), .Z(n4602) );
  AND U4191 ( .A(n4605), .B(n4606), .Z(n4604) );
  ANDN U4192 ( .B(n4607), .A(rc_i[4]), .Z(n4606) );
  AND U4193 ( .A(n4608), .B(n4609), .Z(n4607) );
  XOR U4194 ( .A(n4612), .B(n4613), .Z(out[1542]) );
  XOR U4195 ( .A(n4616), .B(n4617), .Z(out[1541]) );
  XOR U4196 ( .A(n4620), .B(n4621), .Z(out[1540]) );
  XOR U4197 ( .A(n4624), .B(n3956), .Z(out[153]) );
  XOR U4198 ( .A(n4625), .B(n1992), .Z(n3956) );
  ANDN U4199 ( .B(n4167), .A(n1486), .Z(n4624) );
  XNOR U4200 ( .A(n4626), .B(n2515), .Z(n1486) );
  XOR U4201 ( .A(n4627), .B(n2674), .Z(n4167) );
  XOR U4202 ( .A(n4628), .B(n4629), .Z(out[1539]) );
  XOR U4203 ( .A(n4630), .B(n4631), .Z(n4629) );
  AND U4204 ( .A(n4632), .B(n4633), .Z(n4631) );
  AND U4205 ( .A(n4634), .B(n4635), .Z(n4633) );
  NOR U4206 ( .A(rc_i[6]), .B(rc_i[9]), .Z(n4634) );
  AND U4207 ( .A(n4636), .B(n4491), .Z(n4632) );
  NOR U4208 ( .A(rc_i[3]), .B(rc_i[4]), .Z(n4636) );
  XOR U4209 ( .A(n4639), .B(n4640), .Z(out[1538]) );
  XOR U4210 ( .A(n4643), .B(n4644), .Z(out[1537]) );
  XOR U4211 ( .A(n4645), .B(n4646), .Z(n4644) );
  AND U4212 ( .A(n4647), .B(n4648), .Z(n4646) );
  AND U4213 ( .A(n4649), .B(n4608), .Z(n4648) );
  AND U4214 ( .A(n4565), .B(n4635), .Z(n4647) );
  XOR U4215 ( .A(n4652), .B(n4653), .Z(out[1536]) );
  XOR U4216 ( .A(n4654), .B(n4655), .Z(n4653) );
  ANDN U4217 ( .B(n4656), .A(n4342), .Z(n4655) );
  NAND U4218 ( .A(n4608), .B(n4657), .Z(n4342) );
  AND U4219 ( .A(n4490), .B(n4340), .Z(n4656) );
  XOR U4220 ( .A(n4660), .B(n4346), .Z(out[1535]) );
  ANDN U4221 ( .B(n4661), .A(n4345), .Z(n4660) );
  XNOR U4222 ( .A(n4662), .B(n4350), .Z(out[1534]) );
  ANDN U4223 ( .B(n4663), .A(n4349), .Z(n4662) );
  XNOR U4224 ( .A(n4664), .B(n4354), .Z(out[1533]) );
  ANDN U4225 ( .B(n4665), .A(n4353), .Z(n4664) );
  XNOR U4226 ( .A(n4666), .B(n4357), .Z(out[1532]) );
  XNOR U4227 ( .A(n4668), .B(n4361), .Z(out[1531]) );
  AND U4228 ( .A(n4669), .B(n4670), .Z(n4668) );
  XNOR U4229 ( .A(n4671), .B(n4365), .Z(out[1530]) );
  AND U4230 ( .A(n4672), .B(n4673), .Z(n4671) );
  IV U4231 ( .A(n4366), .Z(n4673) );
  XOR U4232 ( .A(n4674), .B(n3959), .Z(out[152]) );
  XOR U4233 ( .A(n4675), .B(n1995), .Z(n3959) );
  ANDN U4234 ( .B(n4170), .A(n1518), .Z(n4674) );
  XOR U4235 ( .A(n4676), .B(n2522), .Z(n1518) );
  XOR U4236 ( .A(n4677), .B(n2681), .Z(n4170) );
  XNOR U4237 ( .A(n4678), .B(n4369), .Z(out[1529]) );
  AND U4238 ( .A(n4679), .B(n4680), .Z(n4678) );
  IV U4239 ( .A(n4370), .Z(n4680) );
  XNOR U4240 ( .A(n4681), .B(n4373), .Z(out[1528]) );
  XNOR U4241 ( .A(n4683), .B(n4377), .Z(out[1527]) );
  XNOR U4242 ( .A(n4685), .B(n4382), .Z(out[1526]) );
  ANDN U4243 ( .B(n4686), .A(n4381), .Z(n4685) );
  XNOR U4244 ( .A(n4687), .B(n4390), .Z(out[1525]) );
  ANDN U4245 ( .B(n4688), .A(n4389), .Z(n4687) );
  XNOR U4246 ( .A(n4689), .B(n4394), .Z(out[1524]) );
  ANDN U4247 ( .B(n4690), .A(n4393), .Z(n4689) );
  XOR U4248 ( .A(n4691), .B(n4398), .Z(out[1523]) );
  ANDN U4249 ( .B(n4692), .A(n4397), .Z(n4691) );
  XNOR U4250 ( .A(n4693), .B(n4402), .Z(out[1522]) );
  ANDN U4251 ( .B(n4694), .A(n4401), .Z(n4693) );
  XNOR U4252 ( .A(n4695), .B(n4406), .Z(out[1521]) );
  ANDN U4253 ( .B(n4696), .A(n4405), .Z(n4695) );
  XNOR U4254 ( .A(n4697), .B(n4410), .Z(out[1520]) );
  ANDN U4255 ( .B(n4698), .A(n4409), .Z(n4697) );
  XOR U4256 ( .A(n4699), .B(n3964), .Z(out[151]) );
  XOR U4257 ( .A(n4700), .B(n1998), .Z(n3964) );
  ANDN U4258 ( .B(n4173), .A(n1542), .Z(n4699) );
  XNOR U4259 ( .A(n4701), .B(n2529), .Z(n1542) );
  XOR U4260 ( .A(n4702), .B(n2688), .Z(n4173) );
  XOR U4261 ( .A(n4703), .B(n4414), .Z(out[1519]) );
  ANDN U4262 ( .B(n4704), .A(n4413), .Z(n4703) );
  XNOR U4263 ( .A(n4705), .B(n4418), .Z(out[1518]) );
  ANDN U4264 ( .B(n4706), .A(n4417), .Z(n4705) );
  XOR U4265 ( .A(n4707), .B(n4422), .Z(out[1517]) );
  ANDN U4266 ( .B(n4708), .A(n4421), .Z(n4707) );
  XOR U4267 ( .A(n4709), .B(n4426), .Z(out[1516]) );
  ANDN U4268 ( .B(n4710), .A(n4425), .Z(n4709) );
  XOR U4269 ( .A(n4711), .B(n4434), .Z(out[1515]) );
  ANDN U4270 ( .B(n4712), .A(n4433), .Z(n4711) );
  XNOR U4271 ( .A(n4713), .B(n4438), .Z(out[1514]) );
  ANDN U4272 ( .B(n4714), .A(n4437), .Z(n4713) );
  XNOR U4273 ( .A(n4715), .B(n4442), .Z(out[1513]) );
  ANDN U4274 ( .B(n4716), .A(n4441), .Z(n4715) );
  XNOR U4275 ( .A(n4717), .B(n4446), .Z(out[1512]) );
  ANDN U4276 ( .B(n4718), .A(n4445), .Z(n4717) );
  XNOR U4277 ( .A(n4719), .B(n4450), .Z(out[1511]) );
  ANDN U4278 ( .B(n4720), .A(n4449), .Z(n4719) );
  XNOR U4279 ( .A(n4721), .B(n4454), .Z(out[1510]) );
  ANDN U4280 ( .B(n4722), .A(n4453), .Z(n4721) );
  XOR U4281 ( .A(n4723), .B(n3967), .Z(out[150]) );
  XOR U4282 ( .A(n4724), .B(n2005), .Z(n3967) );
  ANDN U4283 ( .B(n4176), .A(n1567), .Z(n4723) );
  XNOR U4284 ( .A(n4725), .B(n2536), .Z(n1567) );
  XOR U4285 ( .A(n4726), .B(n2219), .Z(n4176) );
  XNOR U4286 ( .A(n4727), .B(n4458), .Z(out[1509]) );
  ANDN U4287 ( .B(n4728), .A(n4457), .Z(n4727) );
  XNOR U4288 ( .A(n4729), .B(n4462), .Z(out[1508]) );
  ANDN U4289 ( .B(n4730), .A(n4461), .Z(n4729) );
  XNOR U4290 ( .A(n4731), .B(n4466), .Z(out[1507]) );
  ANDN U4291 ( .B(n4732), .A(n4465), .Z(n4731) );
  XNOR U4292 ( .A(n4733), .B(n4469), .Z(out[1506]) );
  AND U4293 ( .A(n4470), .B(n4734), .Z(n4733) );
  XNOR U4294 ( .A(n4735), .B(n4477), .Z(out[1505]) );
  AND U4295 ( .A(n4478), .B(n4736), .Z(n4735) );
  XNOR U4296 ( .A(n4737), .B(n4481), .Z(out[1504]) );
  XNOR U4297 ( .A(n4739), .B(n4493), .Z(out[1503]) );
  ANDN U4298 ( .B(n4740), .A(n4492), .Z(n4739) );
  XNOR U4299 ( .A(n4741), .B(n4497), .Z(out[1502]) );
  ANDN U4300 ( .B(n4742), .A(n4496), .Z(n4741) );
  XNOR U4301 ( .A(n4743), .B(n4501), .Z(out[1501]) );
  ANDN U4302 ( .B(n4744), .A(n4500), .Z(n4743) );
  XNOR U4303 ( .A(n4745), .B(n4505), .Z(out[1500]) );
  ANDN U4304 ( .B(n4746), .A(n4504), .Z(n4745) );
  XNOR U4305 ( .A(n4747), .B(n1866), .Z(out[14]) );
  NOR U4306 ( .A(n3992), .B(n1865), .Z(n4747) );
  XNOR U4307 ( .A(n2526), .B(n4748), .Z(n1865) );
  XOR U4308 ( .A(n4749), .B(n1737), .Z(n3992) );
  XOR U4309 ( .A(n4750), .B(n3970), .Z(out[149]) );
  XOR U4310 ( .A(n4751), .B(n2009), .Z(n3970) );
  ANDN U4311 ( .B(n4179), .A(n1591), .Z(n4750) );
  XOR U4312 ( .A(n4752), .B(n2543), .Z(n1591) );
  XOR U4313 ( .A(n4753), .B(n2226), .Z(n4179) );
  XNOR U4314 ( .A(n4754), .B(n4509), .Z(out[1499]) );
  ANDN U4315 ( .B(n4755), .A(n4508), .Z(n4754) );
  XNOR U4316 ( .A(n4756), .B(n4513), .Z(out[1498]) );
  ANDN U4317 ( .B(n4757), .A(n4512), .Z(n4756) );
  XOR U4318 ( .A(n4758), .B(n4517), .Z(out[1497]) );
  ANDN U4319 ( .B(n4759), .A(n4516), .Z(n4758) );
  XOR U4320 ( .A(n4760), .B(n4521), .Z(out[1496]) );
  ANDN U4321 ( .B(n4761), .A(n4520), .Z(n4760) );
  XOR U4322 ( .A(n4762), .B(n4529), .Z(out[1495]) );
  ANDN U4323 ( .B(n4763), .A(n4528), .Z(n4762) );
  XOR U4324 ( .A(n4764), .B(n4533), .Z(out[1494]) );
  ANDN U4325 ( .B(n4765), .A(n4532), .Z(n4764) );
  XOR U4326 ( .A(n4766), .B(n4537), .Z(out[1493]) );
  ANDN U4327 ( .B(n4767), .A(n4536), .Z(n4766) );
  XOR U4328 ( .A(n4768), .B(n4541), .Z(out[1492]) );
  ANDN U4329 ( .B(n4769), .A(n4540), .Z(n4768) );
  XOR U4330 ( .A(n4770), .B(n4545), .Z(out[1491]) );
  ANDN U4331 ( .B(n4771), .A(n4544), .Z(n4770) );
  XOR U4332 ( .A(n4772), .B(n4549), .Z(out[1490]) );
  NOR U4333 ( .A(n4773), .B(n4548), .Z(n4772) );
  XOR U4334 ( .A(n4774), .B(n3973), .Z(out[148]) );
  XOR U4335 ( .A(n4775), .B(n2013), .Z(n3973) );
  ANDN U4336 ( .B(n4181), .A(n1615), .Z(n4774) );
  XOR U4337 ( .A(n4776), .B(n2554), .Z(n1615) );
  XOR U4338 ( .A(n4777), .B(n2233), .Z(n4181) );
  IV U4339 ( .A(n4778), .Z(n2233) );
  XOR U4340 ( .A(n4779), .B(n4553), .Z(out[1489]) );
  ANDN U4341 ( .B(n4780), .A(n4552), .Z(n4779) );
  XOR U4342 ( .A(n4781), .B(n4557), .Z(out[1488]) );
  NOR U4343 ( .A(n4782), .B(n4556), .Z(n4781) );
  XOR U4344 ( .A(n4783), .B(n4568), .Z(out[1487]) );
  ANDN U4345 ( .B(n4784), .A(n4567), .Z(n4783) );
  XOR U4346 ( .A(n4785), .B(n4572), .Z(out[1486]) );
  ANDN U4347 ( .B(n4786), .A(n4571), .Z(n4785) );
  XOR U4348 ( .A(n4787), .B(n4580), .Z(out[1485]) );
  ANDN U4349 ( .B(n4788), .A(n4579), .Z(n4787) );
  XOR U4350 ( .A(n4789), .B(n4584), .Z(out[1484]) );
  ANDN U4351 ( .B(n4790), .A(n4583), .Z(n4789) );
  XNOR U4352 ( .A(n4791), .B(n4587), .Z(out[1483]) );
  ANDN U4353 ( .B(n4792), .A(n4588), .Z(n4791) );
  XOR U4354 ( .A(n4793), .B(n4592), .Z(out[1482]) );
  ANDN U4355 ( .B(n4794), .A(n4591), .Z(n4793) );
  XOR U4356 ( .A(n4795), .B(n4596), .Z(out[1481]) );
  ANDN U4357 ( .B(n4796), .A(n4595), .Z(n4795) );
  XOR U4358 ( .A(n4797), .B(n4600), .Z(out[1480]) );
  ANDN U4359 ( .B(n4798), .A(n4599), .Z(n4797) );
  XOR U4360 ( .A(n4799), .B(n3976), .Z(out[147]) );
  XOR U4361 ( .A(n4800), .B(n2017), .Z(n3976) );
  ANDN U4362 ( .B(n1637), .A(n1639), .Z(n4799) );
  XOR U4363 ( .A(n4801), .B(n2561), .Z(n1639) );
  XNOR U4364 ( .A(n4802), .B(n2240), .Z(n1637) );
  IV U4365 ( .A(n4803), .Z(n2240) );
  XOR U4366 ( .A(n4804), .B(n4611), .Z(out[1479]) );
  ANDN U4367 ( .B(n4805), .A(n4610), .Z(n4804) );
  XOR U4368 ( .A(n4806), .B(n4615), .Z(out[1478]) );
  ANDN U4369 ( .B(n4807), .A(n4614), .Z(n4806) );
  XOR U4370 ( .A(n4808), .B(n4619), .Z(out[1477]) );
  ANDN U4371 ( .B(n4809), .A(n4618), .Z(n4808) );
  XOR U4372 ( .A(n4810), .B(n4623), .Z(out[1476]) );
  ANDN U4373 ( .B(n4811), .A(n4622), .Z(n4810) );
  XOR U4374 ( .A(n4812), .B(n4638), .Z(out[1475]) );
  ANDN U4375 ( .B(n4813), .A(n4637), .Z(n4812) );
  XOR U4376 ( .A(n4814), .B(n4642), .Z(out[1474]) );
  ANDN U4377 ( .B(n4815), .A(n4641), .Z(n4814) );
  XOR U4378 ( .A(n4816), .B(n4651), .Z(out[1473]) );
  ANDN U4379 ( .B(n4817), .A(n4650), .Z(n4816) );
  XOR U4380 ( .A(n4818), .B(n4659), .Z(out[1472]) );
  ANDN U4381 ( .B(n4819), .A(n4658), .Z(n4818) );
  XOR U4382 ( .A(n4820), .B(n4345), .Z(out[1471]) );
  XNOR U4383 ( .A(n4821), .B(n4822), .Z(n4345) );
  AND U4384 ( .A(n4823), .B(n4824), .Z(n4820) );
  XOR U4385 ( .A(n4825), .B(n4349), .Z(out[1470]) );
  XNOR U4386 ( .A(n4826), .B(n4827), .Z(n4349) );
  ANDN U4387 ( .B(n4828), .A(n4663), .Z(n4825) );
  XNOR U4388 ( .A(n4829), .B(n3980), .Z(out[146]) );
  XNOR U4389 ( .A(n4830), .B(n2021), .Z(n3980) );
  ANDN U4390 ( .B(n1666), .A(n1668), .Z(n4829) );
  XOR U4391 ( .A(n4831), .B(n2568), .Z(n1668) );
  XNOR U4392 ( .A(n4832), .B(n2254), .Z(n1666) );
  IV U4393 ( .A(n4833), .Z(n2254) );
  XOR U4394 ( .A(n4834), .B(n4353), .Z(out[1469]) );
  XOR U4395 ( .A(n4835), .B(n2513), .Z(n4353) );
  ANDN U4396 ( .B(n4836), .A(n4665), .Z(n4834) );
  XOR U4397 ( .A(n4837), .B(n4358), .Z(out[1468]) );
  XOR U4398 ( .A(n4838), .B(n4839), .Z(n4358) );
  ANDN U4399 ( .B(n4840), .A(n4667), .Z(n4837) );
  XOR U4400 ( .A(n4841), .B(n4362), .Z(out[1467]) );
  IV U4401 ( .A(n4670), .Z(n4362) );
  XOR U4402 ( .A(n2526), .B(n4842), .Z(n4670) );
  ANDN U4403 ( .B(n4843), .A(n4669), .Z(n4841) );
  XOR U4404 ( .A(n4844), .B(n4366), .Z(out[1466]) );
  XOR U4405 ( .A(n4845), .B(n4846), .Z(n4366) );
  ANDN U4406 ( .B(n4847), .A(n4672), .Z(n4844) );
  XOR U4407 ( .A(n4848), .B(n4370), .Z(out[1465]) );
  XOR U4408 ( .A(n3485), .B(n4849), .Z(n4370) );
  ANDN U4409 ( .B(n4850), .A(n4679), .Z(n4848) );
  XOR U4410 ( .A(n4851), .B(n4374), .Z(out[1464]) );
  XOR U4411 ( .A(n3488), .B(n4852), .Z(n4374) );
  ANDN U4412 ( .B(n4853), .A(n4682), .Z(n4851) );
  XOR U4413 ( .A(n4854), .B(n4378), .Z(out[1463]) );
  XOR U4414 ( .A(n3491), .B(n4855), .Z(n4378) );
  ANDN U4415 ( .B(n4856), .A(n4684), .Z(n4854) );
  XOR U4416 ( .A(n4857), .B(n4381), .Z(out[1462]) );
  XNOR U4417 ( .A(n4858), .B(n4859), .Z(n4381) );
  ANDN U4418 ( .B(n4860), .A(n4686), .Z(n4857) );
  XOR U4419 ( .A(n4861), .B(n4389), .Z(out[1461]) );
  XOR U4420 ( .A(n4862), .B(n2573), .Z(n4389) );
  ANDN U4421 ( .B(n4863), .A(n4688), .Z(n4861) );
  XOR U4422 ( .A(n4864), .B(n4393), .Z(out[1460]) );
  XOR U4423 ( .A(n4865), .B(n2580), .Z(n4393) );
  ANDN U4424 ( .B(n4866), .A(n4690), .Z(n4864) );
  XOR U4425 ( .A(n4867), .B(n3983), .Z(out[145]) );
  XOR U4426 ( .A(n4868), .B(n2024), .Z(n3983) );
  ANDN U4427 ( .B(n1721), .A(n1719), .Z(n4867) );
  XNOR U4428 ( .A(n4869), .B(n3802), .Z(n1719) );
  XOR U4429 ( .A(n4870), .B(n2575), .Z(n1721) );
  XOR U4430 ( .A(n4871), .B(n4397), .Z(out[1459]) );
  XOR U4431 ( .A(n4872), .B(n2587), .Z(n4397) );
  ANDN U4432 ( .B(n4873), .A(n4692), .Z(n4871) );
  XOR U4433 ( .A(n4874), .B(n4401), .Z(out[1458]) );
  XOR U4434 ( .A(n4875), .B(n2594), .Z(n4401) );
  ANDN U4435 ( .B(n4876), .A(n4694), .Z(n4874) );
  XOR U4436 ( .A(n4877), .B(n4405), .Z(out[1457]) );
  XOR U4437 ( .A(n4878), .B(n2601), .Z(n4405) );
  ANDN U4438 ( .B(n4879), .A(n4696), .Z(n4877) );
  XOR U4439 ( .A(n4880), .B(n4409), .Z(out[1456]) );
  XOR U4440 ( .A(n4881), .B(n2608), .Z(n4409) );
  ANDN U4441 ( .B(n4882), .A(n4698), .Z(n4880) );
  XOR U4442 ( .A(n4883), .B(n4413), .Z(out[1455]) );
  XOR U4443 ( .A(n4884), .B(n2615), .Z(n4413) );
  ANDN U4444 ( .B(n4885), .A(n4704), .Z(n4883) );
  XOR U4445 ( .A(n4886), .B(n4417), .Z(out[1454]) );
  XOR U4446 ( .A(n4887), .B(n2627), .Z(n4417) );
  ANDN U4447 ( .B(n4888), .A(n4706), .Z(n4886) );
  XOR U4448 ( .A(n4889), .B(n4421), .Z(out[1453]) );
  XOR U4449 ( .A(n4890), .B(n2634), .Z(n4421) );
  ANDN U4450 ( .B(n4891), .A(n4708), .Z(n4889) );
  XOR U4451 ( .A(n4892), .B(n4425), .Z(out[1452]) );
  XOR U4452 ( .A(n4893), .B(n2641), .Z(n4425) );
  ANDN U4453 ( .B(n4894), .A(n4710), .Z(n4892) );
  XOR U4454 ( .A(n4895), .B(n4433), .Z(out[1451]) );
  XOR U4455 ( .A(n4896), .B(n2648), .Z(n4433) );
  ANDN U4456 ( .B(n4897), .A(n4712), .Z(n4895) );
  XOR U4457 ( .A(n4898), .B(n4437), .Z(out[1450]) );
  XOR U4458 ( .A(n4899), .B(n2655), .Z(n4437) );
  ANDN U4459 ( .B(n4900), .A(n4714), .Z(n4898) );
  XNOR U4460 ( .A(n4901), .B(n3987), .Z(out[144]) );
  XOR U4461 ( .A(n4902), .B(n2028), .Z(n3987) );
  ANDN U4462 ( .B(n1770), .A(n1771), .Z(n4901) );
  XOR U4463 ( .A(n4903), .B(n2582), .Z(n1771) );
  XNOR U4464 ( .A(n4904), .B(n2268), .Z(n1770) );
  IV U4465 ( .A(n4905), .Z(n2268) );
  XOR U4466 ( .A(n4906), .B(n4441), .Z(out[1449]) );
  XOR U4467 ( .A(n4907), .B(n2662), .Z(n4441) );
  ANDN U4468 ( .B(n4908), .A(n4716), .Z(n4906) );
  XOR U4469 ( .A(n4909), .B(n4445), .Z(out[1448]) );
  XOR U4470 ( .A(n4910), .B(n2669), .Z(n4445) );
  ANDN U4471 ( .B(n4911), .A(n4718), .Z(n4909) );
  XOR U4472 ( .A(n4912), .B(n4449), .Z(out[1447]) );
  XOR U4473 ( .A(n4913), .B(n2676), .Z(n4449) );
  XOR U4474 ( .A(n4915), .B(n4453), .Z(out[1446]) );
  XOR U4475 ( .A(n4916), .B(n2683), .Z(n4453) );
  AND U4476 ( .A(n4917), .B(n4918), .Z(n4915) );
  XOR U4477 ( .A(n4919), .B(n4457), .Z(out[1445]) );
  XOR U4478 ( .A(n4920), .B(n2690), .Z(n4457) );
  AND U4479 ( .A(n4921), .B(n4922), .Z(n4919) );
  XOR U4480 ( .A(n4923), .B(n4461), .Z(out[1444]) );
  XOR U4481 ( .A(n4924), .B(n4925), .Z(n4461) );
  AND U4482 ( .A(n4926), .B(n4927), .Z(n4923) );
  XOR U4483 ( .A(n4928), .B(n4465), .Z(out[1443]) );
  XOR U4484 ( .A(n4929), .B(n3555), .Z(n4465) );
  AND U4485 ( .A(n4930), .B(n4931), .Z(n4928) );
  XNOR U4486 ( .A(n4932), .B(n4470), .Z(out[1442]) );
  XNOR U4487 ( .A(n4933), .B(n3558), .Z(n4470) );
  AND U4488 ( .A(n4934), .B(n4935), .Z(n4932) );
  XNOR U4489 ( .A(n4936), .B(n4478), .Z(out[1441]) );
  XNOR U4490 ( .A(n4937), .B(n2242), .Z(n4478) );
  AND U4491 ( .A(n4938), .B(n4939), .Z(n4936) );
  IV U4492 ( .A(n4736), .Z(n4939) );
  XOR U4493 ( .A(n4940), .B(n4482), .Z(out[1440]) );
  XOR U4494 ( .A(n4941), .B(n2256), .Z(n4482) );
  NOR U4495 ( .A(n4942), .B(n4738), .Z(n4940) );
  XNOR U4496 ( .A(n4943), .B(n3990), .Z(out[143]) );
  XOR U4497 ( .A(n4944), .B(n2032), .Z(n3990) );
  ANDN U4498 ( .B(n1819), .A(n1821), .Z(n4943) );
  XOR U4499 ( .A(n4945), .B(n2589), .Z(n1821) );
  XNOR U4500 ( .A(n4946), .B(n2275), .Z(n1819) );
  IV U4501 ( .A(n4947), .Z(n2275) );
  XOR U4502 ( .A(n4948), .B(n4492), .Z(out[1439]) );
  XOR U4503 ( .A(n4949), .B(n2263), .Z(n4492) );
  ANDN U4504 ( .B(n4950), .A(n4740), .Z(n4948) );
  XOR U4505 ( .A(n4951), .B(n4496), .Z(out[1438]) );
  XOR U4506 ( .A(n4952), .B(n2270), .Z(n4496) );
  ANDN U4507 ( .B(n4953), .A(n4742), .Z(n4951) );
  XOR U4508 ( .A(n4954), .B(n4500), .Z(out[1437]) );
  XOR U4509 ( .A(n4955), .B(n2277), .Z(n4500) );
  NOR U4510 ( .A(n4956), .B(n4744), .Z(n4954) );
  XOR U4511 ( .A(n4957), .B(n4504), .Z(out[1436]) );
  XOR U4512 ( .A(n4958), .B(n2284), .Z(n4504) );
  NOR U4513 ( .A(n4959), .B(n4746), .Z(n4957) );
  XOR U4514 ( .A(n4960), .B(n4508), .Z(out[1435]) );
  XOR U4515 ( .A(n4961), .B(n2291), .Z(n4508) );
  NOR U4516 ( .A(n4962), .B(n4755), .Z(n4960) );
  XOR U4517 ( .A(n4963), .B(n4512), .Z(out[1434]) );
  XOR U4518 ( .A(n4964), .B(n2298), .Z(n4512) );
  NOR U4519 ( .A(n4965), .B(n4757), .Z(n4963) );
  XOR U4520 ( .A(n4966), .B(n4516), .Z(out[1433]) );
  XOR U4521 ( .A(n4967), .B(n2305), .Z(n4516) );
  ANDN U4522 ( .B(n4968), .A(n4759), .Z(n4966) );
  XOR U4523 ( .A(n4969), .B(n4520), .Z(out[1432]) );
  XOR U4524 ( .A(n4970), .B(n2312), .Z(n4520) );
  ANDN U4525 ( .B(n4971), .A(n4761), .Z(n4969) );
  XOR U4526 ( .A(n4972), .B(n4528), .Z(out[1431]) );
  XOR U4527 ( .A(n4973), .B(n2319), .Z(n4528) );
  ANDN U4528 ( .B(n4974), .A(n4763), .Z(n4972) );
  XOR U4529 ( .A(n4975), .B(n4532), .Z(out[1430]) );
  XOR U4530 ( .A(n4976), .B(n2330), .Z(n4532) );
  ANDN U4531 ( .B(n4977), .A(n4765), .Z(n4975) );
  XNOR U4532 ( .A(n4978), .B(n3993), .Z(out[142]) );
  XOR U4533 ( .A(n4979), .B(n2036), .Z(n3993) );
  ANDN U4534 ( .B(n1864), .A(n1866), .Z(n4978) );
  XOR U4535 ( .A(n4980), .B(n2596), .Z(n1866) );
  XNOR U4536 ( .A(n4981), .B(n2282), .Z(n1864) );
  IV U4537 ( .A(n4982), .Z(n2282) );
  XOR U4538 ( .A(n4983), .B(n4536), .Z(out[1429]) );
  XNOR U4539 ( .A(n4984), .B(n4985), .Z(n4536) );
  ANDN U4540 ( .B(n4986), .A(n4767), .Z(n4983) );
  XOR U4541 ( .A(n4987), .B(n4540), .Z(out[1428]) );
  XNOR U4542 ( .A(n4988), .B(n4989), .Z(n4540) );
  AND U4543 ( .A(n4990), .B(n4991), .Z(n4987) );
  XOR U4544 ( .A(n4992), .B(n4544), .Z(out[1427]) );
  XNOR U4545 ( .A(n4993), .B(n4994), .Z(n4544) );
  AND U4546 ( .A(n4995), .B(n4996), .Z(n4992) );
  XOR U4547 ( .A(n4997), .B(n4548), .Z(out[1426]) );
  XNOR U4548 ( .A(n4998), .B(n4999), .Z(n4548) );
  AND U4549 ( .A(n4773), .B(n5000), .Z(n4997) );
  XOR U4550 ( .A(n5001), .B(n4552), .Z(out[1425]) );
  XNOR U4551 ( .A(n5002), .B(n5003), .Z(n4552) );
  AND U4552 ( .A(n5004), .B(n5005), .Z(n5001) );
  XOR U4553 ( .A(n5006), .B(n4556), .Z(out[1424]) );
  XNOR U4554 ( .A(n5007), .B(n5008), .Z(n4556) );
  AND U4555 ( .A(n4782), .B(n5009), .Z(n5006) );
  XOR U4556 ( .A(n5010), .B(n4567), .Z(out[1423]) );
  XNOR U4557 ( .A(n5011), .B(n5012), .Z(n4567) );
  AND U4558 ( .A(n5013), .B(n5014), .Z(n5010) );
  XOR U4559 ( .A(n5015), .B(n4571), .Z(out[1422]) );
  XOR U4560 ( .A(n2387), .B(n5016), .Z(n4571) );
  XOR U4561 ( .A(n5018), .B(n4579), .Z(out[1421]) );
  XNOR U4562 ( .A(n5019), .B(n5020), .Z(n4579) );
  XOR U4563 ( .A(n5022), .B(n4583), .Z(out[1420]) );
  XOR U4564 ( .A(n5023), .B(n5024), .Z(n4583) );
  XNOR U4565 ( .A(n5026), .B(n3998), .Z(out[141]) );
  XOR U4566 ( .A(n5027), .B(n2040), .Z(n3998) );
  AND U4567 ( .A(n1910), .B(n1912), .Z(n5026) );
  XNOR U4568 ( .A(n5028), .B(n2289), .Z(n1910) );
  XOR U4569 ( .A(n5029), .B(n4588), .Z(out[1419]) );
  XOR U4570 ( .A(n5030), .B(n2411), .Z(n4588) );
  AND U4571 ( .A(n5031), .B(n5032), .Z(n5029) );
  XOR U4572 ( .A(n5033), .B(n4591), .Z(out[1418]) );
  XOR U4573 ( .A(n5034), .B(n2418), .Z(n4591) );
  AND U4574 ( .A(n5035), .B(n5036), .Z(n5033) );
  XOR U4575 ( .A(n5037), .B(n4595), .Z(out[1417]) );
  XNOR U4576 ( .A(n5038), .B(n5039), .Z(n4595) );
  AND U4577 ( .A(n5040), .B(n5041), .Z(n5037) );
  XOR U4578 ( .A(n5042), .B(n4599), .Z(out[1416]) );
  XNOR U4579 ( .A(n5043), .B(n5044), .Z(n4599) );
  AND U4580 ( .A(n5045), .B(n5046), .Z(n5042) );
  XOR U4581 ( .A(n5047), .B(n4610), .Z(out[1415]) );
  XNOR U4582 ( .A(n5048), .B(n5049), .Z(n4610) );
  AND U4583 ( .A(n5050), .B(n5051), .Z(n5047) );
  XOR U4584 ( .A(n5052), .B(n4614), .Z(out[1414]) );
  XNOR U4585 ( .A(n5053), .B(n5054), .Z(n4614) );
  AND U4586 ( .A(n5055), .B(n5056), .Z(n5052) );
  XOR U4587 ( .A(n5057), .B(n4618), .Z(out[1413]) );
  XNOR U4588 ( .A(n5058), .B(n5059), .Z(n4618) );
  AND U4589 ( .A(n5060), .B(n5061), .Z(n5057) );
  XOR U4590 ( .A(n5062), .B(n4622), .Z(out[1412]) );
  XNOR U4591 ( .A(n5063), .B(n5064), .Z(n4622) );
  AND U4592 ( .A(n5065), .B(n5066), .Z(n5062) );
  XOR U4593 ( .A(n5067), .B(n4637), .Z(out[1411]) );
  XNOR U4594 ( .A(n5068), .B(n5069), .Z(n4637) );
  AND U4595 ( .A(n5070), .B(n5071), .Z(n5067) );
  XOR U4596 ( .A(n5072), .B(n4641), .Z(out[1410]) );
  XNOR U4597 ( .A(n5073), .B(n5074), .Z(n4641) );
  AND U4598 ( .A(n5075), .B(n5076), .Z(n5072) );
  XNOR U4599 ( .A(n5077), .B(n4001), .Z(out[140]) );
  XOR U4600 ( .A(n5078), .B(n2048), .Z(n4001) );
  AND U4601 ( .A(n1963), .B(n1961), .Z(n5077) );
  XNOR U4602 ( .A(n5079), .B(n2296), .Z(n1961) );
  IV U4603 ( .A(n5080), .Z(n2296) );
  XOR U4604 ( .A(n5081), .B(n4650), .Z(out[1409]) );
  XNOR U4605 ( .A(n5082), .B(n5083), .Z(n4650) );
  AND U4606 ( .A(n5084), .B(n5085), .Z(n5081) );
  XOR U4607 ( .A(n5086), .B(n4658), .Z(out[1408]) );
  XNOR U4608 ( .A(n5087), .B(n5088), .Z(n4658) );
  AND U4609 ( .A(n5089), .B(n5090), .Z(n5086) );
  XOR U4610 ( .A(n5091), .B(n4661), .Z(out[1407]) );
  IV U4611 ( .A(n4824), .Z(n4661) );
  XOR U4612 ( .A(n1951), .B(n5092), .Z(n4824) );
  NOR U4613 ( .A(n4333), .B(n4823), .Z(n5091) );
  XOR U4614 ( .A(n5093), .B(n4663), .Z(out[1406]) );
  XNOR U4615 ( .A(n5094), .B(n1957), .Z(n4663) );
  ANDN U4616 ( .B(n4348), .A(n4828), .Z(n5093) );
  XOR U4617 ( .A(n5095), .B(n4665), .Z(out[1405]) );
  XNOR U4618 ( .A(n5096), .B(n1966), .Z(n4665) );
  ANDN U4619 ( .B(n4352), .A(n4836), .Z(n5095) );
  XOR U4620 ( .A(n5097), .B(n4667), .Z(out[1404]) );
  XNOR U4621 ( .A(n5098), .B(n1971), .Z(n4667) );
  ANDN U4622 ( .B(n4356), .A(n4840), .Z(n5097) );
  XOR U4623 ( .A(n5099), .B(n4669), .Z(out[1403]) );
  XNOR U4624 ( .A(n5100), .B(n1658), .Z(n4669) );
  ANDN U4625 ( .B(n4360), .A(n4843), .Z(n5099) );
  XOR U4626 ( .A(n5101), .B(n4672), .Z(out[1402]) );
  XNOR U4627 ( .A(n5102), .B(n1663), .Z(n4672) );
  ANDN U4628 ( .B(n4364), .A(n4847), .Z(n5101) );
  XOR U4629 ( .A(n5103), .B(n4679), .Z(out[1401]) );
  XNOR U4630 ( .A(n5104), .B(n1671), .Z(n4679) );
  XOR U4631 ( .A(n5105), .B(n4682), .Z(out[1400]) );
  XOR U4632 ( .A(n5106), .B(n1675), .Z(n4682) );
  XOR U4633 ( .A(n5107), .B(n1912), .Z(out[13]) );
  XOR U4634 ( .A(n5108), .B(n2603), .Z(n1912) );
  NOR U4635 ( .A(n3997), .B(n1911), .Z(n5107) );
  XNOR U4636 ( .A(n2533), .B(n5109), .Z(n1911) );
  XOR U4637 ( .A(n5110), .B(n1742), .Z(n3997) );
  XNOR U4638 ( .A(n5111), .B(n4004), .Z(out[139]) );
  XOR U4639 ( .A(n5112), .B(n2052), .Z(n4004) );
  AND U4640 ( .A(n2000), .B(n2002), .Z(n5111) );
  XNOR U4641 ( .A(n5113), .B(n2303), .Z(n2000) );
  IV U4642 ( .A(n5114), .Z(n2303) );
  XOR U4643 ( .A(n5115), .B(n4684), .Z(out[1399]) );
  XOR U4644 ( .A(n5116), .B(n1680), .Z(n4684) );
  ANDN U4645 ( .B(n4376), .A(n4856), .Z(n5115) );
  XOR U4646 ( .A(n5117), .B(n4686), .Z(out[1398]) );
  XNOR U4647 ( .A(n5118), .B(n1685), .Z(n4686) );
  ANDN U4648 ( .B(n4380), .A(n4860), .Z(n5117) );
  XOR U4649 ( .A(n5119), .B(n4688), .Z(out[1397]) );
  XNOR U4650 ( .A(n5120), .B(n1690), .Z(n4688) );
  ANDN U4651 ( .B(n4388), .A(n4863), .Z(n5119) );
  XOR U4652 ( .A(n5121), .B(n4690), .Z(out[1396]) );
  XNOR U4653 ( .A(n5122), .B(n1695), .Z(n4690) );
  ANDN U4654 ( .B(n4392), .A(n4866), .Z(n5121) );
  XOR U4655 ( .A(n5123), .B(n4692), .Z(out[1395]) );
  XNOR U4656 ( .A(n5124), .B(n1700), .Z(n4692) );
  ANDN U4657 ( .B(n4396), .A(n4873), .Z(n5123) );
  XOR U4658 ( .A(n5125), .B(n4694), .Z(out[1394]) );
  XNOR U4659 ( .A(n5126), .B(n1705), .Z(n4694) );
  ANDN U4660 ( .B(n4400), .A(n4876), .Z(n5125) );
  XOR U4661 ( .A(n5127), .B(n4696), .Z(out[1393]) );
  XOR U4662 ( .A(n5128), .B(n1710), .Z(n4696) );
  ANDN U4663 ( .B(n4404), .A(n4879), .Z(n5127) );
  XOR U4664 ( .A(n5129), .B(n4698), .Z(out[1392]) );
  XOR U4665 ( .A(n5130), .B(n1715), .Z(n4698) );
  ANDN U4666 ( .B(n4408), .A(n4882), .Z(n5129) );
  XOR U4667 ( .A(n5131), .B(n4704), .Z(out[1391]) );
  XNOR U4668 ( .A(n5132), .B(n1724), .Z(n4704) );
  AND U4669 ( .A(n4412), .B(n5133), .Z(n5131) );
  XOR U4670 ( .A(n5134), .B(n4706), .Z(out[1390]) );
  XNOR U4671 ( .A(n5135), .B(n1728), .Z(n4706) );
  ANDN U4672 ( .B(n4416), .A(n4888), .Z(n5134) );
  XNOR U4673 ( .A(n5136), .B(n4007), .Z(out[138]) );
  XOR U4674 ( .A(n5137), .B(n2056), .Z(n4007) );
  AND U4675 ( .A(n2043), .B(n2045), .Z(n5136) );
  XNOR U4676 ( .A(n5138), .B(n2310), .Z(n2043) );
  XOR U4677 ( .A(n5139), .B(n4708), .Z(out[1389]) );
  XNOR U4678 ( .A(n5140), .B(n1732), .Z(n4708) );
  AND U4679 ( .A(n4420), .B(n5141), .Z(n5139) );
  XOR U4680 ( .A(n5142), .B(n4710), .Z(out[1388]) );
  XNOR U4681 ( .A(n5143), .B(n1737), .Z(n4710) );
  AND U4682 ( .A(n4424), .B(n5144), .Z(n5142) );
  XOR U4683 ( .A(n5145), .B(n4712), .Z(out[1387]) );
  XNOR U4684 ( .A(n5146), .B(n1742), .Z(n4712) );
  AND U4685 ( .A(n4432), .B(n5147), .Z(n5145) );
  IV U4686 ( .A(n4897), .Z(n5147) );
  XOR U4687 ( .A(n5148), .B(n4714), .Z(out[1386]) );
  XNOR U4688 ( .A(n5149), .B(n1747), .Z(n4714) );
  ANDN U4689 ( .B(n4436), .A(n4900), .Z(n5148) );
  XOR U4690 ( .A(n5150), .B(n4716), .Z(out[1385]) );
  XNOR U4691 ( .A(n5151), .B(n1752), .Z(n4716) );
  ANDN U4692 ( .B(n4440), .A(n4908), .Z(n5150) );
  XOR U4693 ( .A(n5152), .B(n4718), .Z(out[1384]) );
  XNOR U4694 ( .A(n5153), .B(n1757), .Z(n4718) );
  ANDN U4695 ( .B(n4444), .A(n4911), .Z(n5152) );
  XOR U4696 ( .A(n5154), .B(n4720), .Z(out[1383]) );
  XOR U4697 ( .A(n1761), .B(n5155), .Z(n4720) );
  IV U4698 ( .A(n5156), .Z(n1761) );
  ANDN U4699 ( .B(n4448), .A(n4914), .Z(n5154) );
  XOR U4700 ( .A(n5157), .B(n4722), .Z(out[1382]) );
  IV U4701 ( .A(n4918), .Z(n4722) );
  XOR U4702 ( .A(n5158), .B(n1766), .Z(n4918) );
  IV U4703 ( .A(n5159), .Z(n1766) );
  ANDN U4704 ( .B(n4452), .A(n4917), .Z(n5157) );
  XOR U4705 ( .A(n5160), .B(n4728), .Z(out[1381]) );
  IV U4706 ( .A(n4922), .Z(n4728) );
  XOR U4707 ( .A(n5161), .B(n1775), .Z(n4922) );
  IV U4708 ( .A(n5162), .Z(n1775) );
  ANDN U4709 ( .B(n4456), .A(n4921), .Z(n5160) );
  XOR U4710 ( .A(n5163), .B(n4730), .Z(out[1380]) );
  IV U4711 ( .A(n4927), .Z(n4730) );
  XOR U4712 ( .A(n5164), .B(n1780), .Z(n4927) );
  IV U4713 ( .A(n5165), .Z(n1780) );
  NOR U4714 ( .A(n4460), .B(n4926), .Z(n5163) );
  XOR U4715 ( .A(n5166), .B(n4010), .Z(out[137]) );
  IV U4716 ( .A(n4197), .Z(n4010) );
  XOR U4717 ( .A(n5167), .B(n2060), .Z(n4197) );
  IV U4718 ( .A(n5168), .Z(n2060) );
  AND U4719 ( .A(n2083), .B(n1040), .Z(n5166) );
  IV U4720 ( .A(n2084), .Z(n1040) );
  XOR U4721 ( .A(n5169), .B(n2635), .Z(n2084) );
  XNOR U4722 ( .A(n5170), .B(n2317), .Z(n2083) );
  XOR U4723 ( .A(n5171), .B(n4732), .Z(out[1379]) );
  IV U4724 ( .A(n4931), .Z(n4732) );
  XOR U4725 ( .A(n5172), .B(n1784), .Z(n4931) );
  IV U4726 ( .A(n5173), .Z(n1784) );
  ANDN U4727 ( .B(n4464), .A(n4930), .Z(n5171) );
  XOR U4728 ( .A(n5174), .B(n4734), .Z(out[1378]) );
  IV U4729 ( .A(n4935), .Z(n4734) );
  XOR U4730 ( .A(n5175), .B(n1788), .Z(n4935) );
  IV U4731 ( .A(n5176), .Z(n1788) );
  ANDN U4732 ( .B(n4468), .A(n4934), .Z(n5174) );
  XOR U4733 ( .A(n5177), .B(n4736), .Z(out[1377]) );
  XOR U4734 ( .A(n5178), .B(n1792), .Z(n4736) );
  IV U4735 ( .A(n5179), .Z(n1792) );
  NOR U4736 ( .A(n4938), .B(n4476), .Z(n5177) );
  XOR U4737 ( .A(n5180), .B(n4738), .Z(out[1376]) );
  XOR U4738 ( .A(n5181), .B(n5182), .Z(n4738) );
  ANDN U4739 ( .B(n4942), .A(n4480), .Z(n5180) );
  XOR U4740 ( .A(n5183), .B(n4740), .Z(out[1375]) );
  XOR U4741 ( .A(n5184), .B(n1800), .Z(n4740) );
  NOR U4742 ( .A(n4483), .B(n4950), .Z(n5183) );
  XOR U4743 ( .A(n5185), .B(n4742), .Z(out[1374]) );
  XNOR U4744 ( .A(n5186), .B(n5187), .Z(n4742) );
  NOR U4745 ( .A(n4495), .B(n4953), .Z(n5185) );
  XOR U4746 ( .A(n5188), .B(n4744), .Z(out[1373]) );
  XNOR U4747 ( .A(n5189), .B(n5190), .Z(n4744) );
  ANDN U4748 ( .B(n4956), .A(n4499), .Z(n5188) );
  XOR U4749 ( .A(n5191), .B(n4746), .Z(out[1372]) );
  XNOR U4750 ( .A(n5192), .B(n5193), .Z(n4746) );
  AND U4751 ( .A(n4959), .B(n4503), .Z(n5191) );
  IV U4752 ( .A(n5194), .Z(n4503) );
  XOR U4753 ( .A(n5195), .B(n4755), .Z(out[1371]) );
  XNOR U4754 ( .A(n5196), .B(n5197), .Z(n4755) );
  AND U4755 ( .A(n4962), .B(n4507), .Z(n5195) );
  IV U4756 ( .A(n5198), .Z(n4507) );
  XOR U4757 ( .A(n5199), .B(n4757), .Z(out[1370]) );
  XNOR U4758 ( .A(n5200), .B(n5201), .Z(n4757) );
  AND U4759 ( .A(n4965), .B(n4511), .Z(n5199) );
  IV U4760 ( .A(n5202), .Z(n4511) );
  XOR U4761 ( .A(n5203), .B(n4013), .Z(out[136]) );
  IV U4762 ( .A(n4200), .Z(n4013) );
  XOR U4763 ( .A(n5204), .B(n2063), .Z(n4200) );
  ANDN U4764 ( .B(n2122), .A(n1480), .Z(n5203) );
  XOR U4765 ( .A(n5205), .B(n2643), .Z(n1480) );
  XNOR U4766 ( .A(n5206), .B(n2328), .Z(n2122) );
  IV U4767 ( .A(n5207), .Z(n2328) );
  XOR U4768 ( .A(n5208), .B(n4759), .Z(out[1369]) );
  XNOR U4769 ( .A(n5209), .B(n5210), .Z(n4759) );
  AND U4770 ( .A(n4515), .B(n5211), .Z(n5208) );
  XOR U4771 ( .A(n5212), .B(n4761), .Z(out[1368]) );
  XNOR U4772 ( .A(n5213), .B(n5214), .Z(n4761) );
  AND U4773 ( .A(n4519), .B(n5215), .Z(n5212) );
  XOR U4774 ( .A(n5216), .B(n4763), .Z(out[1367]) );
  XNOR U4775 ( .A(n5217), .B(n5218), .Z(n4763) );
  ANDN U4776 ( .B(n4527), .A(n4974), .Z(n5216) );
  XOR U4777 ( .A(n5219), .B(n4765), .Z(out[1366]) );
  XNOR U4778 ( .A(n5220), .B(n5221), .Z(n4765) );
  AND U4779 ( .A(n4531), .B(n5222), .Z(n5219) );
  XOR U4780 ( .A(n5223), .B(n4767), .Z(out[1365]) );
  XNOR U4781 ( .A(n5224), .B(n5225), .Z(n4767) );
  NOR U4782 ( .A(n4535), .B(n4986), .Z(n5223) );
  XOR U4783 ( .A(n5226), .B(n4769), .Z(out[1364]) );
  IV U4784 ( .A(n4991), .Z(n4769) );
  XOR U4785 ( .A(n5227), .B(n5228), .Z(n4991) );
  NOR U4786 ( .A(n4539), .B(n4990), .Z(n5226) );
  XOR U4787 ( .A(n5229), .B(n4771), .Z(out[1363]) );
  IV U4788 ( .A(n4996), .Z(n4771) );
  XOR U4789 ( .A(n5230), .B(n5231), .Z(n4996) );
  NOR U4790 ( .A(n4543), .B(n4995), .Z(n5229) );
  XNOR U4791 ( .A(n5232), .B(n4773), .Z(out[1362]) );
  XNOR U4792 ( .A(n1860), .B(n5233), .Z(n4773) );
  ANDN U4793 ( .B(n5234), .A(n4547), .Z(n5232) );
  XOR U4794 ( .A(n5235), .B(n4780), .Z(out[1361]) );
  IV U4795 ( .A(n5005), .Z(n4780) );
  XOR U4796 ( .A(n5236), .B(n5237), .Z(n5005) );
  ANDN U4797 ( .B(n4551), .A(n5004), .Z(n5235) );
  XNOR U4798 ( .A(n5238), .B(n4782), .Z(out[1360]) );
  XNOR U4799 ( .A(n1872), .B(n5239), .Z(n4782) );
  ANDN U4800 ( .B(n5240), .A(n4555), .Z(n5238) );
  XOR U4801 ( .A(n5241), .B(n4017), .Z(out[135]) );
  XNOR U4802 ( .A(n5242), .B(n2066), .Z(n4017) );
  ANDN U4803 ( .B(n2161), .A(n1815), .Z(n5241) );
  XNOR U4804 ( .A(n5243), .B(n2650), .Z(n1815) );
  XNOR U4805 ( .A(n5244), .B(n2335), .Z(n2161) );
  XOR U4806 ( .A(n5245), .B(n4784), .Z(out[1359]) );
  IV U4807 ( .A(n5014), .Z(n4784) );
  XOR U4808 ( .A(n5246), .B(n5247), .Z(n5014) );
  XOR U4809 ( .A(n5248), .B(n4786), .Z(out[1358]) );
  XOR U4810 ( .A(n1880), .B(n5249), .Z(n4786) );
  NOR U4811 ( .A(n5017), .B(n4570), .Z(n5248) );
  XOR U4812 ( .A(n5250), .B(n4788), .Z(out[1357]) );
  XOR U4813 ( .A(n5251), .B(n5252), .Z(n4788) );
  NOR U4814 ( .A(n4578), .B(n5021), .Z(n5250) );
  XOR U4815 ( .A(n5253), .B(n4790), .Z(out[1356]) );
  XOR U4816 ( .A(n5254), .B(n5255), .Z(n4790) );
  ANDN U4817 ( .B(n4582), .A(n5025), .Z(n5253) );
  XOR U4818 ( .A(n5256), .B(n4792), .Z(out[1355]) );
  IV U4819 ( .A(n5032), .Z(n4792) );
  XOR U4820 ( .A(n5257), .B(n5258), .Z(n5032) );
  NOR U4821 ( .A(n4586), .B(n5031), .Z(n5256) );
  XOR U4822 ( .A(n5259), .B(n4794), .Z(out[1354]) );
  IV U4823 ( .A(n5036), .Z(n4794) );
  XOR U4824 ( .A(n5260), .B(n5261), .Z(n5036) );
  ANDN U4825 ( .B(n4590), .A(n5035), .Z(n5259) );
  XOR U4826 ( .A(n5262), .B(n4796), .Z(out[1353]) );
  IV U4827 ( .A(n5041), .Z(n4796) );
  XOR U4828 ( .A(n5263), .B(n5264), .Z(n5041) );
  ANDN U4829 ( .B(n4594), .A(n5040), .Z(n5262) );
  XOR U4830 ( .A(n5265), .B(n4798), .Z(out[1352]) );
  IV U4831 ( .A(n5046), .Z(n4798) );
  XOR U4832 ( .A(n5266), .B(n5267), .Z(n5046) );
  ANDN U4833 ( .B(n4598), .A(n5045), .Z(n5265) );
  XOR U4834 ( .A(n5268), .B(n4805), .Z(out[1351]) );
  IV U4835 ( .A(n5051), .Z(n4805) );
  XOR U4836 ( .A(n5269), .B(n5270), .Z(n5051) );
  NOR U4837 ( .A(n4601), .B(n5050), .Z(n5268) );
  XOR U4838 ( .A(n5271), .B(n4807), .Z(out[1350]) );
  IV U4839 ( .A(n5056), .Z(n4807) );
  XOR U4840 ( .A(n5272), .B(n5273), .Z(n5056) );
  ANDN U4841 ( .B(n4613), .A(n5055), .Z(n5271) );
  XOR U4842 ( .A(n5274), .B(n4021), .Z(out[134]) );
  XOR U4843 ( .A(n5275), .B(n2070), .Z(n4021) );
  ANDN U4844 ( .B(n2196), .A(n2197), .Z(n5274) );
  XOR U4845 ( .A(n5276), .B(n2657), .Z(n2197) );
  XNOR U4846 ( .A(n5277), .B(n2342), .Z(n2196) );
  XOR U4847 ( .A(n5278), .B(n4809), .Z(out[1349]) );
  IV U4848 ( .A(n5061), .Z(n4809) );
  XOR U4849 ( .A(n5279), .B(n5280), .Z(n5061) );
  ANDN U4850 ( .B(n4617), .A(n5060), .Z(n5278) );
  XOR U4851 ( .A(n5281), .B(n4811), .Z(out[1348]) );
  IV U4852 ( .A(n5066), .Z(n4811) );
  XOR U4853 ( .A(n5282), .B(n5283), .Z(n5066) );
  ANDN U4854 ( .B(n4621), .A(n5065), .Z(n5281) );
  XOR U4855 ( .A(n5284), .B(n4813), .Z(out[1347]) );
  IV U4856 ( .A(n5071), .Z(n4813) );
  XOR U4857 ( .A(n5285), .B(n5286), .Z(n5071) );
  NOR U4858 ( .A(n4628), .B(n5070), .Z(n5284) );
  XOR U4859 ( .A(n5287), .B(n4815), .Z(out[1346]) );
  IV U4860 ( .A(n5076), .Z(n4815) );
  XOR U4861 ( .A(n5288), .B(n5289), .Z(n5076) );
  ANDN U4862 ( .B(n4640), .A(n5075), .Z(n5287) );
  XOR U4863 ( .A(n5290), .B(n4817), .Z(out[1345]) );
  IV U4864 ( .A(n5085), .Z(n4817) );
  XNOR U4865 ( .A(n1941), .B(n5291), .Z(n5085) );
  NOR U4866 ( .A(n4643), .B(n5084), .Z(n5290) );
  XOR U4867 ( .A(n5292), .B(n4819), .Z(out[1344]) );
  IV U4868 ( .A(n5090), .Z(n4819) );
  XNOR U4869 ( .A(n1946), .B(n5293), .Z(n5090) );
  NOR U4870 ( .A(n4652), .B(n5089), .Z(n5292) );
  XOR U4871 ( .A(n5294), .B(n4823), .Z(out[1343]) );
  XOR U4872 ( .A(n5295), .B(n1995), .Z(n4823) );
  AND U4873 ( .A(n4333), .B(n4346), .Z(n5294) );
  XOR U4874 ( .A(n5296), .B(n2543), .Z(n4346) );
  XOR U4875 ( .A(n5297), .B(n2564), .Z(n4333) );
  XOR U4876 ( .A(n5298), .B(n4828), .Z(out[1342]) );
  XOR U4877 ( .A(n5299), .B(n1998), .Z(n4828) );
  NOR U4878 ( .A(n4350), .B(n4348), .Z(n5298) );
  XOR U4879 ( .A(n5300), .B(n2571), .Z(n4348) );
  XNOR U4880 ( .A(n5301), .B(n2554), .Z(n4350) );
  IV U4881 ( .A(n3284), .Z(n2554) );
  XOR U4882 ( .A(n5302), .B(n4836), .Z(out[1341]) );
  XOR U4883 ( .A(n5303), .B(n2005), .Z(n4836) );
  NOR U4884 ( .A(n4354), .B(n4352), .Z(n5302) );
  XNOR U4885 ( .A(n5304), .B(n2578), .Z(n4352) );
  XNOR U4886 ( .A(n5305), .B(n2561), .Z(n4354) );
  IV U4887 ( .A(n5306), .Z(n2561) );
  XOR U4888 ( .A(n5307), .B(n4840), .Z(out[1340]) );
  XOR U4889 ( .A(n5308), .B(n2009), .Z(n4840) );
  NOR U4890 ( .A(n4357), .B(n4356), .Z(n5307) );
  XNOR U4891 ( .A(n5309), .B(n2585), .Z(n4356) );
  XOR U4892 ( .A(n5310), .B(n2568), .Z(n4357) );
  IV U4893 ( .A(n5311), .Z(n2568) );
  XOR U4894 ( .A(n5312), .B(n4024), .Z(out[133]) );
  XOR U4895 ( .A(n5313), .B(n2073), .Z(n4024) );
  AND U4896 ( .A(n2251), .B(n4212), .Z(n5312) );
  XOR U4897 ( .A(n5314), .B(n2349), .Z(n4212) );
  XOR U4898 ( .A(n5315), .B(n3339), .Z(n2251) );
  IV U4899 ( .A(n2664), .Z(n3339) );
  XOR U4900 ( .A(n5316), .B(n4843), .Z(out[1339]) );
  XOR U4901 ( .A(n5317), .B(n2013), .Z(n4843) );
  NOR U4902 ( .A(n4361), .B(n4360), .Z(n5316) );
  XNOR U4903 ( .A(n5318), .B(n2592), .Z(n4360) );
  XOR U4904 ( .A(n5319), .B(n2575), .Z(n4361) );
  XOR U4905 ( .A(n5320), .B(n4847), .Z(out[1338]) );
  XOR U4906 ( .A(n5321), .B(n2017), .Z(n4847) );
  NOR U4907 ( .A(n4365), .B(n4364), .Z(n5320) );
  XNOR U4908 ( .A(n2598), .B(n5322), .Z(n4364) );
  IV U4909 ( .A(n5323), .Z(n2598) );
  XNOR U4910 ( .A(n5324), .B(n2582), .Z(n4365) );
  IV U4911 ( .A(n5325), .Z(n2582) );
  XOR U4912 ( .A(n5326), .B(n4850), .Z(out[1337]) );
  XOR U4913 ( .A(n5327), .B(n2021), .Z(n4850) );
  IV U4914 ( .A(n5328), .Z(n2021) );
  NOR U4915 ( .A(n4369), .B(n4368), .Z(n5326) );
  XNOR U4916 ( .A(n2605), .B(n5329), .Z(n4368) );
  IV U4917 ( .A(n5330), .Z(n2605) );
  XNOR U4918 ( .A(n5331), .B(n2589), .Z(n4369) );
  IV U4919 ( .A(n5332), .Z(n2589) );
  XOR U4920 ( .A(n5333), .B(n4853), .Z(out[1336]) );
  XOR U4921 ( .A(n5334), .B(n2024), .Z(n4853) );
  IV U4922 ( .A(n5335), .Z(n2024) );
  NOR U4923 ( .A(n4373), .B(n4372), .Z(n5333) );
  XNOR U4924 ( .A(n2612), .B(n5336), .Z(n4372) );
  IV U4925 ( .A(n4319), .Z(n2612) );
  XNOR U4926 ( .A(n5337), .B(n2596), .Z(n4373) );
  IV U4927 ( .A(n5338), .Z(n2596) );
  XOR U4928 ( .A(n5339), .B(n4856), .Z(out[1335]) );
  XOR U4929 ( .A(n5340), .B(n2028), .Z(n4856) );
  NOR U4930 ( .A(n4377), .B(n4376), .Z(n5339) );
  XOR U4931 ( .A(n5341), .B(n2625), .Z(n4376) );
  XNOR U4932 ( .A(n5342), .B(n2603), .Z(n4377) );
  IV U4933 ( .A(n5343), .Z(n2603) );
  XOR U4934 ( .A(n5344), .B(n4860), .Z(out[1334]) );
  XOR U4935 ( .A(n5345), .B(n2032), .Z(n4860) );
  NOR U4936 ( .A(n4382), .B(n4380), .Z(n5344) );
  XOR U4937 ( .A(n5346), .B(n2632), .Z(n4380) );
  XNOR U4938 ( .A(n5347), .B(n2610), .Z(n4382) );
  XOR U4939 ( .A(n5348), .B(n4863), .Z(out[1333]) );
  XOR U4940 ( .A(n5349), .B(n2036), .Z(n4863) );
  NOR U4941 ( .A(n4390), .B(n4388), .Z(n5348) );
  XNOR U4942 ( .A(n5350), .B(n2639), .Z(n4388) );
  XOR U4943 ( .A(n5351), .B(n2617), .Z(n4390) );
  XOR U4944 ( .A(n5352), .B(n4866), .Z(out[1332]) );
  XOR U4945 ( .A(n5353), .B(n2040), .Z(n4866) );
  NOR U4946 ( .A(n4394), .B(n4392), .Z(n5352) );
  XNOR U4947 ( .A(n5354), .B(n2646), .Z(n4392) );
  XOR U4948 ( .A(n5355), .B(n2629), .Z(n4394) );
  XOR U4949 ( .A(n5356), .B(n4873), .Z(out[1331]) );
  XNOR U4950 ( .A(n5357), .B(n2048), .Z(n4873) );
  ANDN U4951 ( .B(n4398), .A(n4396), .Z(n5356) );
  XNOR U4952 ( .A(n5358), .B(n2653), .Z(n4396) );
  XOR U4953 ( .A(n2635), .B(n5359), .Z(n4398) );
  IV U4954 ( .A(n5360), .Z(n2635) );
  XOR U4955 ( .A(n5361), .B(n4876), .Z(out[1330]) );
  XOR U4956 ( .A(n5362), .B(n2052), .Z(n4876) );
  NOR U4957 ( .A(n4402), .B(n4400), .Z(n5361) );
  XNOR U4958 ( .A(n5363), .B(n2660), .Z(n4400) );
  XOR U4959 ( .A(n5364), .B(n2643), .Z(n4402) );
  IV U4960 ( .A(n5365), .Z(n2643) );
  XOR U4961 ( .A(n5366), .B(n4027), .Z(out[132]) );
  XOR U4962 ( .A(n5367), .B(n2076), .Z(n4027) );
  ANDN U4963 ( .B(n2323), .A(n2324), .Z(n5366) );
  XOR U4964 ( .A(n5368), .B(n2671), .Z(n2324) );
  XNOR U4965 ( .A(n5369), .B(n2356), .Z(n2323) );
  XOR U4966 ( .A(n5370), .B(n4879), .Z(out[1329]) );
  XOR U4967 ( .A(n5371), .B(n2056), .Z(n4879) );
  NOR U4968 ( .A(n4406), .B(n4404), .Z(n5370) );
  XNOR U4969 ( .A(n5372), .B(n2667), .Z(n4404) );
  XOR U4970 ( .A(n5373), .B(n2650), .Z(n4406) );
  IV U4971 ( .A(n5374), .Z(n2650) );
  XOR U4972 ( .A(n5375), .B(n4882), .Z(out[1328]) );
  XOR U4973 ( .A(n5376), .B(n5168), .Z(n4882) );
  NOR U4974 ( .A(n4410), .B(n4408), .Z(n5375) );
  XNOR U4975 ( .A(n5377), .B(n2674), .Z(n4408) );
  XOR U4976 ( .A(n5378), .B(n2657), .Z(n4410) );
  IV U4977 ( .A(n5379), .Z(n2657) );
  XOR U4978 ( .A(n5380), .B(n4885), .Z(out[1327]) );
  IV U4979 ( .A(n5133), .Z(n4885) );
  XOR U4980 ( .A(n5381), .B(n2063), .Z(n5133) );
  IV U4981 ( .A(n5382), .Z(n2063) );
  ANDN U4982 ( .B(n4414), .A(n4412), .Z(n5380) );
  XNOR U4983 ( .A(n5383), .B(n2681), .Z(n4412) );
  XNOR U4984 ( .A(n5384), .B(n2664), .Z(n4414) );
  XOR U4985 ( .A(n5385), .B(n4888), .Z(out[1326]) );
  XNOR U4986 ( .A(n5386), .B(n2066), .Z(n4888) );
  NOR U4987 ( .A(n4418), .B(n4416), .Z(n5385) );
  XNOR U4988 ( .A(n5387), .B(n2688), .Z(n4416) );
  XOR U4989 ( .A(n5388), .B(n2671), .Z(n4418) );
  IV U4990 ( .A(n3344), .Z(n2671) );
  XOR U4991 ( .A(n5389), .B(n4891), .Z(out[1325]) );
  IV U4992 ( .A(n5141), .Z(n4891) );
  XOR U4993 ( .A(n5390), .B(n2070), .Z(n5141) );
  IV U4994 ( .A(n5391), .Z(n2070) );
  ANDN U4995 ( .B(n4422), .A(n4420), .Z(n5389) );
  XNOR U4996 ( .A(n5392), .B(n2219), .Z(n4420) );
  XNOR U4997 ( .A(n5393), .B(n2678), .Z(n4422) );
  XOR U4998 ( .A(n5394), .B(n4894), .Z(out[1324]) );
  IV U4999 ( .A(n5144), .Z(n4894) );
  XOR U5000 ( .A(n5395), .B(n2073), .Z(n5144) );
  IV U5001 ( .A(n5396), .Z(n2073) );
  ANDN U5002 ( .B(n4426), .A(n4424), .Z(n5394) );
  XNOR U5003 ( .A(n5397), .B(n2226), .Z(n4424) );
  XNOR U5004 ( .A(n5398), .B(n2685), .Z(n4426) );
  XOR U5005 ( .A(n5399), .B(n4897), .Z(out[1323]) );
  XOR U5006 ( .A(n5400), .B(n2076), .Z(n4897) );
  IV U5007 ( .A(n5401), .Z(n2076) );
  ANDN U5008 ( .B(n4434), .A(n4432), .Z(n5399) );
  XOR U5009 ( .A(n5402), .B(n4778), .Z(n4432) );
  XNOR U5010 ( .A(n5403), .B(n2692), .Z(n4434) );
  XOR U5011 ( .A(n5404), .B(n4900), .Z(out[1322]) );
  XNOR U5012 ( .A(n5405), .B(n2080), .Z(n4900) );
  NOR U5013 ( .A(n4438), .B(n4436), .Z(n5404) );
  XOR U5014 ( .A(n5406), .B(n4803), .Z(n4436) );
  XOR U5015 ( .A(n2222), .B(n5407), .Z(n4438) );
  XOR U5016 ( .A(n5408), .B(n4908), .Z(out[1321]) );
  XNOR U5017 ( .A(n5409), .B(n2087), .Z(n4908) );
  NOR U5018 ( .A(n4442), .B(n4440), .Z(n5408) );
  XNOR U5019 ( .A(n5410), .B(n4833), .Z(n4440) );
  XOR U5020 ( .A(n2229), .B(n5411), .Z(n4442) );
  XOR U5021 ( .A(n5412), .B(n4911), .Z(out[1320]) );
  XNOR U5022 ( .A(n5413), .B(n2090), .Z(n4911) );
  NOR U5023 ( .A(n4446), .B(n4444), .Z(n5412) );
  XNOR U5024 ( .A(n5414), .B(n3802), .Z(n4444) );
  XOR U5025 ( .A(n2236), .B(n5415), .Z(n4446) );
  XOR U5026 ( .A(n5416), .B(n4032), .Z(out[131]) );
  IV U5027 ( .A(n4217), .Z(n4032) );
  XNOR U5028 ( .A(n5417), .B(n2080), .Z(n4217) );
  AND U5029 ( .A(n2399), .B(n4218), .Z(n5416) );
  XOR U5030 ( .A(n5418), .B(n2363), .Z(n4218) );
  XOR U5031 ( .A(n5419), .B(n3353), .Z(n2399) );
  IV U5032 ( .A(n2678), .Z(n3353) );
  XOR U5033 ( .A(n5420), .B(n4914), .Z(out[1319]) );
  XNOR U5034 ( .A(n5421), .B(n2094), .Z(n4914) );
  NOR U5035 ( .A(n4450), .B(n4448), .Z(n5420) );
  XNOR U5036 ( .A(n5422), .B(n4905), .Z(n4448) );
  XOR U5037 ( .A(n2243), .B(n5423), .Z(n4450) );
  XOR U5038 ( .A(n5424), .B(n4917), .Z(out[1318]) );
  XNOR U5039 ( .A(n5425), .B(n2098), .Z(n4917) );
  NOR U5040 ( .A(n4454), .B(n4452), .Z(n5424) );
  XNOR U5041 ( .A(n5426), .B(n4947), .Z(n4452) );
  XOR U5042 ( .A(n2257), .B(n5427), .Z(n4454) );
  XOR U5043 ( .A(n5428), .B(n4921), .Z(out[1317]) );
  XNOR U5044 ( .A(n5429), .B(n2101), .Z(n4921) );
  NOR U5045 ( .A(n4458), .B(n4456), .Z(n5428) );
  XNOR U5046 ( .A(n5430), .B(n4982), .Z(n4456) );
  XNOR U5047 ( .A(n5431), .B(n2265), .Z(n4458) );
  XOR U5048 ( .A(n5432), .B(n4926), .Z(out[1316]) );
  XNOR U5049 ( .A(n5433), .B(n2105), .Z(n4926) );
  ANDN U5050 ( .B(n4460), .A(n4462), .Z(n5432) );
  XNOR U5051 ( .A(n5434), .B(n2272), .Z(n4462) );
  XNOR U5052 ( .A(n5435), .B(n2289), .Z(n4460) );
  IV U5053 ( .A(n5436), .Z(n2289) );
  XOR U5054 ( .A(n5437), .B(n4930), .Z(out[1315]) );
  XNOR U5055 ( .A(n5438), .B(n2108), .Z(n4930) );
  NOR U5056 ( .A(n4466), .B(n4464), .Z(n5437) );
  XNOR U5057 ( .A(n5439), .B(n5080), .Z(n4464) );
  XNOR U5058 ( .A(n5440), .B(n2279), .Z(n4466) );
  XOR U5059 ( .A(n5441), .B(n4934), .Z(out[1314]) );
  XNOR U5060 ( .A(n5442), .B(n2111), .Z(n4934) );
  NOR U5061 ( .A(n4469), .B(n4468), .Z(n5441) );
  XOR U5062 ( .A(n5443), .B(n5114), .Z(n4468) );
  XOR U5063 ( .A(n5444), .B(n2286), .Z(n4469) );
  XOR U5064 ( .A(n5445), .B(n4938), .Z(out[1313]) );
  XOR U5065 ( .A(n5446), .B(n5447), .Z(n4938) );
  ANDN U5066 ( .B(n4476), .A(n4477), .Z(n5445) );
  XOR U5067 ( .A(n5448), .B(n2293), .Z(n4477) );
  XNOR U5068 ( .A(n5449), .B(n2310), .Z(n4476) );
  IV U5069 ( .A(n5450), .Z(n2310) );
  XNOR U5070 ( .A(n5451), .B(n4942), .Z(out[1312]) );
  XNOR U5071 ( .A(n5452), .B(n5453), .Z(n4942) );
  ANDN U5072 ( .B(n4480), .A(n4481), .Z(n5451) );
  XOR U5073 ( .A(n5454), .B(n2300), .Z(n4481) );
  XNOR U5074 ( .A(n5455), .B(n2317), .Z(n4480) );
  IV U5075 ( .A(n5456), .Z(n2317) );
  XOR U5076 ( .A(n5457), .B(n4950), .Z(out[1311]) );
  XOR U5077 ( .A(n5458), .B(n2125), .Z(n4950) );
  ANDN U5078 ( .B(n4483), .A(n4493), .Z(n5457) );
  XOR U5079 ( .A(n5459), .B(n2307), .Z(n4493) );
  XNOR U5080 ( .A(n5460), .B(n5207), .Z(n4483) );
  XOR U5081 ( .A(n5461), .B(n4953), .Z(out[1310]) );
  XNOR U5082 ( .A(n2127), .B(n5462), .Z(n4953) );
  ANDN U5083 ( .B(n4495), .A(n4497), .Z(n5461) );
  XOR U5084 ( .A(n5463), .B(n2314), .Z(n4497) );
  XNOR U5085 ( .A(n5464), .B(n2335), .Z(n4495) );
  IV U5086 ( .A(n5465), .Z(n2335) );
  XOR U5087 ( .A(n5466), .B(n4035), .Z(out[130]) );
  IV U5088 ( .A(n4221), .Z(n4035) );
  XNOR U5089 ( .A(n5467), .B(n2087), .Z(n4221) );
  ANDN U5090 ( .B(n2473), .A(n2471), .Z(n5466) );
  XOR U5091 ( .A(n5468), .B(n3586), .Z(n2471) );
  XOR U5092 ( .A(n5469), .B(n3358), .Z(n2473) );
  IV U5093 ( .A(n2685), .Z(n3358) );
  XNOR U5094 ( .A(n5470), .B(n4956), .Z(out[1309]) );
  XNOR U5095 ( .A(n5471), .B(n5472), .Z(n4956) );
  ANDN U5096 ( .B(n4499), .A(n4501), .Z(n5470) );
  XNOR U5097 ( .A(n5473), .B(n2321), .Z(n4501) );
  XNOR U5098 ( .A(n5474), .B(n2342), .Z(n4499) );
  IV U5099 ( .A(n5475), .Z(n2342) );
  XNOR U5100 ( .A(n5476), .B(n4959), .Z(out[1308]) );
  XNOR U5101 ( .A(n5477), .B(n5478), .Z(n4959) );
  ANDN U5102 ( .B(n5194), .A(n4505), .Z(n5476) );
  XNOR U5103 ( .A(n5479), .B(n2332), .Z(n4505) );
  XOR U5104 ( .A(n5480), .B(n2349), .Z(n5194) );
  IV U5105 ( .A(n5481), .Z(n2349) );
  XNOR U5106 ( .A(n5482), .B(n4962), .Z(out[1307]) );
  XOR U5107 ( .A(n2139), .B(n5483), .Z(n4962) );
  ANDN U5108 ( .B(n5198), .A(n4509), .Z(n5482) );
  XNOR U5109 ( .A(n5484), .B(n2337), .Z(n4509) );
  XOR U5110 ( .A(n5485), .B(n2356), .Z(n5198) );
  IV U5111 ( .A(n5486), .Z(n2356) );
  XNOR U5112 ( .A(n5487), .B(n4965), .Z(out[1306]) );
  XOR U5113 ( .A(n2143), .B(n5488), .Z(n4965) );
  ANDN U5114 ( .B(n5202), .A(n4513), .Z(n5487) );
  XNOR U5115 ( .A(n5489), .B(n2344), .Z(n4513) );
  XOR U5116 ( .A(n5490), .B(n2363), .Z(n5202) );
  IV U5117 ( .A(n5491), .Z(n2363) );
  XOR U5118 ( .A(n5492), .B(n4968), .Z(out[1305]) );
  IV U5119 ( .A(n5211), .Z(n4968) );
  XOR U5120 ( .A(n2147), .B(n5493), .Z(n5211) );
  ANDN U5121 ( .B(n4517), .A(n4515), .Z(n5492) );
  XNOR U5122 ( .A(n5494), .B(n3586), .Z(n4515) );
  XOR U5123 ( .A(n5495), .B(n2351), .Z(n4517) );
  XOR U5124 ( .A(n5496), .B(n4971), .Z(out[1304]) );
  IV U5125 ( .A(n5215), .Z(n4971) );
  XOR U5126 ( .A(n5497), .B(n2152), .Z(n5215) );
  ANDN U5127 ( .B(n4521), .A(n4519), .Z(n5496) );
  XNOR U5128 ( .A(n5498), .B(n3591), .Z(n4519) );
  XOR U5129 ( .A(n5499), .B(n2358), .Z(n4521) );
  XOR U5130 ( .A(n5500), .B(n4974), .Z(out[1303]) );
  XOR U5131 ( .A(n5501), .B(n2155), .Z(n4974) );
  ANDN U5132 ( .B(n4529), .A(n4527), .Z(n5500) );
  XNOR U5133 ( .A(n5502), .B(n5503), .Z(n4527) );
  XOR U5134 ( .A(n5504), .B(n2365), .Z(n4529) );
  XOR U5135 ( .A(n5505), .B(n4977), .Z(out[1302]) );
  IV U5136 ( .A(n5222), .Z(n4977) );
  XNOR U5137 ( .A(n5506), .B(n2159), .Z(n5222) );
  ANDN U5138 ( .B(n4533), .A(n4531), .Z(n5505) );
  XOR U5139 ( .A(n5507), .B(n5508), .Z(n4531) );
  XOR U5140 ( .A(n5509), .B(n2374), .Z(n4533) );
  XOR U5141 ( .A(n5510), .B(n4986), .Z(out[1301]) );
  XOR U5142 ( .A(n5511), .B(n2164), .Z(n4986) );
  AND U5143 ( .A(n4535), .B(n4537), .Z(n5510) );
  XOR U5144 ( .A(n5512), .B(n2379), .Z(n4537) );
  XNOR U5145 ( .A(n5513), .B(n2402), .Z(n4535) );
  XOR U5146 ( .A(n5514), .B(n4990), .Z(out[1300]) );
  XOR U5147 ( .A(n5515), .B(n2168), .Z(n4990) );
  AND U5148 ( .A(n4539), .B(n4541), .Z(n5514) );
  XOR U5149 ( .A(n5516), .B(n2386), .Z(n4541) );
  XNOR U5150 ( .A(n5517), .B(n2409), .Z(n4539) );
  XOR U5151 ( .A(n5518), .B(n1963), .Z(out[12]) );
  XNOR U5152 ( .A(n5519), .B(n2610), .Z(n1963) );
  IV U5153 ( .A(n5520), .Z(n2610) );
  NOR U5154 ( .A(n4000), .B(n1962), .Z(n5518) );
  XNOR U5155 ( .A(n2540), .B(n5521), .Z(n1962) );
  XOR U5156 ( .A(n5522), .B(n1747), .Z(n4000) );
  XOR U5157 ( .A(n5523), .B(n4038), .Z(out[129]) );
  XNOR U5158 ( .A(n5524), .B(n2090), .Z(n4038) );
  ANDN U5159 ( .B(n2547), .A(n2545), .Z(n5523) );
  XOR U5160 ( .A(n5525), .B(n3591), .Z(n2545) );
  XOR U5161 ( .A(n5526), .B(n3363), .Z(n2547) );
  IV U5162 ( .A(n2692), .Z(n3363) );
  XOR U5163 ( .A(n5527), .B(n4995), .Z(out[1299]) );
  XNOR U5164 ( .A(n5528), .B(n2172), .Z(n4995) );
  AND U5165 ( .A(n4543), .B(n4545), .Z(n5527) );
  XOR U5166 ( .A(n5529), .B(n2395), .Z(n4545) );
  XNOR U5167 ( .A(n5530), .B(n2416), .Z(n4543) );
  XOR U5168 ( .A(n5531), .B(n5000), .Z(out[1298]) );
  IV U5169 ( .A(n5234), .Z(n5000) );
  XNOR U5170 ( .A(n5532), .B(n2175), .Z(n5234) );
  AND U5171 ( .A(n4547), .B(n4549), .Z(n5531) );
  XOR U5172 ( .A(n5533), .B(n2404), .Z(n4549) );
  XNOR U5173 ( .A(n5534), .B(n2423), .Z(n4547) );
  XOR U5174 ( .A(n5535), .B(n5004), .Z(out[1297]) );
  XNOR U5175 ( .A(n5536), .B(n2178), .Z(n5004) );
  ANDN U5176 ( .B(n4553), .A(n4551), .Z(n5535) );
  XNOR U5177 ( .A(n5537), .B(n2430), .Z(n4551) );
  XOR U5178 ( .A(n5538), .B(n2413), .Z(n4553) );
  XOR U5179 ( .A(n5539), .B(n5009), .Z(out[1296]) );
  IV U5180 ( .A(n5240), .Z(n5009) );
  XNOR U5181 ( .A(n5540), .B(n2181), .Z(n5240) );
  AND U5182 ( .A(n4555), .B(n4557), .Z(n5539) );
  XOR U5183 ( .A(n5541), .B(n2420), .Z(n4557) );
  XNOR U5184 ( .A(n5542), .B(n2437), .Z(n4555) );
  XOR U5185 ( .A(n5543), .B(n5013), .Z(out[1295]) );
  XNOR U5186 ( .A(n5544), .B(n4295), .Z(n5013) );
  AND U5187 ( .A(n4568), .B(n4558), .Z(n5543) );
  XOR U5188 ( .A(n5545), .B(n2444), .Z(n4558) );
  XOR U5189 ( .A(n5546), .B(n2427), .Z(n4568) );
  XOR U5190 ( .A(n5547), .B(n5017), .Z(out[1294]) );
  XOR U5191 ( .A(n5548), .B(n2188), .Z(n5017) );
  AND U5192 ( .A(n4570), .B(n4572), .Z(n5547) );
  XOR U5193 ( .A(n5549), .B(n2434), .Z(n4572) );
  XNOR U5194 ( .A(n5550), .B(n2451), .Z(n4570) );
  XOR U5195 ( .A(n5551), .B(n5021), .Z(out[1293]) );
  XNOR U5196 ( .A(n5552), .B(n2191), .Z(n5021) );
  AND U5197 ( .A(n4578), .B(n4580), .Z(n5551) );
  XOR U5198 ( .A(n2438), .B(n5553), .Z(n4580) );
  XNOR U5199 ( .A(n5554), .B(n2458), .Z(n4578) );
  XOR U5200 ( .A(n5555), .B(n5025), .Z(out[1292]) );
  XOR U5201 ( .A(n5556), .B(n2194), .Z(n5025) );
  ANDN U5202 ( .B(n4584), .A(n4582), .Z(n5555) );
  XNOR U5203 ( .A(n5557), .B(n5558), .Z(n4582) );
  XOR U5204 ( .A(n2445), .B(n5559), .Z(n4584) );
  XOR U5205 ( .A(n5560), .B(n5031), .Z(out[1291]) );
  XOR U5206 ( .A(n5561), .B(n2201), .Z(n5031) );
  ANDN U5207 ( .B(n4586), .A(n4587), .Z(n5560) );
  XNOR U5208 ( .A(n5562), .B(n2455), .Z(n4587) );
  XNOR U5209 ( .A(n5563), .B(n2476), .Z(n4586) );
  XOR U5210 ( .A(n5564), .B(n5035), .Z(out[1290]) );
  XOR U5211 ( .A(n5565), .B(n2204), .Z(n5035) );
  ANDN U5212 ( .B(n4592), .A(n4590), .Z(n5564) );
  XOR U5213 ( .A(n5566), .B(n2483), .Z(n4590) );
  XNOR U5214 ( .A(n5567), .B(n2462), .Z(n4592) );
  XOR U5215 ( .A(n5568), .B(n4042), .Z(out[128]) );
  XNOR U5216 ( .A(n5569), .B(n2094), .Z(n4042) );
  AND U5217 ( .A(n2622), .B(n2619), .Z(n5568) );
  XOR U5218 ( .A(n5570), .B(n2384), .Z(n2619) );
  IV U5219 ( .A(n5503), .Z(n2384) );
  XOR U5220 ( .A(n5571), .B(n5040), .Z(out[1289]) );
  XOR U5221 ( .A(n5572), .B(n2207), .Z(n5040) );
  ANDN U5222 ( .B(n4596), .A(n4594), .Z(n5571) );
  XOR U5223 ( .A(n5573), .B(n2490), .Z(n4594) );
  XNOR U5224 ( .A(n5574), .B(n2469), .Z(n4596) );
  XOR U5225 ( .A(n5575), .B(n5045), .Z(out[1288]) );
  XOR U5226 ( .A(n5576), .B(n2210), .Z(n5045) );
  ANDN U5227 ( .B(n4600), .A(n4598), .Z(n5575) );
  XOR U5228 ( .A(n5577), .B(n2497), .Z(n4598) );
  XNOR U5229 ( .A(n5578), .B(n2480), .Z(n4600) );
  XOR U5230 ( .A(n5579), .B(n5050), .Z(out[1287]) );
  XOR U5231 ( .A(n5580), .B(n2213), .Z(n5050) );
  AND U5232 ( .A(n4601), .B(n4611), .Z(n5579) );
  XOR U5233 ( .A(n5581), .B(n2487), .Z(n4611) );
  XOR U5234 ( .A(n5582), .B(n2504), .Z(n4601) );
  XOR U5235 ( .A(n5583), .B(n5055), .Z(out[1286]) );
  XNOR U5236 ( .A(n5584), .B(n5585), .Z(n5055) );
  ANDN U5237 ( .B(n4615), .A(n4613), .Z(n5583) );
  XOR U5238 ( .A(n5586), .B(n2511), .Z(n4613) );
  XOR U5239 ( .A(n5587), .B(n2492), .Z(n4615) );
  XOR U5240 ( .A(n5588), .B(n5060), .Z(out[1285]) );
  XNOR U5241 ( .A(n5589), .B(n5590), .Z(n5060) );
  ANDN U5242 ( .B(n4619), .A(n4617), .Z(n5588) );
  XOR U5243 ( .A(n5591), .B(n2518), .Z(n4617) );
  XOR U5244 ( .A(n5592), .B(n2499), .Z(n4619) );
  XOR U5245 ( .A(n5593), .B(n5065), .Z(out[1284]) );
  XNOR U5246 ( .A(n5594), .B(n5595), .Z(n5065) );
  ANDN U5247 ( .B(n4623), .A(n4621), .Z(n5593) );
  XOR U5248 ( .A(n5596), .B(n2525), .Z(n4621) );
  XOR U5249 ( .A(n5597), .B(n2508), .Z(n4623) );
  XOR U5250 ( .A(n5598), .B(n5070), .Z(out[1283]) );
  XNOR U5251 ( .A(n5599), .B(n5600), .Z(n5070) );
  AND U5252 ( .A(n4628), .B(n4638), .Z(n5598) );
  XOR U5253 ( .A(n5601), .B(n2515), .Z(n4638) );
  XOR U5254 ( .A(n5602), .B(n2532), .Z(n4628) );
  XOR U5255 ( .A(n5603), .B(n5075), .Z(out[1282]) );
  XOR U5256 ( .A(n5604), .B(n1985), .Z(n5075) );
  ANDN U5257 ( .B(n4642), .A(n4640), .Z(n5603) );
  XOR U5258 ( .A(n5605), .B(n2539), .Z(n4640) );
  XOR U5259 ( .A(n5606), .B(n2522), .Z(n4642) );
  XOR U5260 ( .A(n5607), .B(n5084), .Z(out[1281]) );
  XOR U5261 ( .A(n5608), .B(n1988), .Z(n5084) );
  AND U5262 ( .A(n4643), .B(n4651), .Z(n5607) );
  XOR U5263 ( .A(n5609), .B(n2529), .Z(n4651) );
  XOR U5264 ( .A(n5610), .B(n2550), .Z(n4643) );
  XOR U5265 ( .A(n5611), .B(n5089), .Z(out[1280]) );
  XOR U5266 ( .A(n5612), .B(n1992), .Z(n5089) );
  AND U5267 ( .A(n4652), .B(n4659), .Z(n5611) );
  XOR U5268 ( .A(n5613), .B(n2536), .Z(n4659) );
  XOR U5269 ( .A(n5614), .B(n2557), .Z(n4652) );
  XOR U5270 ( .A(n5615), .B(n4046), .Z(out[127]) );
  IV U5271 ( .A(n4227), .Z(n4046) );
  XOR U5272 ( .A(n5616), .B(n2391), .Z(n4227) );
  IV U5273 ( .A(n5508), .Z(n2391) );
  NOR U5274 ( .A(n2696), .B(n2694), .Z(n5615) );
  XNOR U5275 ( .A(n2229), .B(n5617), .Z(n2694) );
  XOR U5276 ( .A(n5618), .B(n2641), .Z(n2696) );
  XOR U5277 ( .A(n5619), .B(n5620), .Z(out[1279]) );
  ANDN U5278 ( .B(n5621), .A(n5622), .Z(n5619) );
  XOR U5279 ( .A(n5623), .B(n5624), .Z(out[1278]) );
  ANDN U5280 ( .B(n5625), .A(n5626), .Z(n5623) );
  XOR U5281 ( .A(n5627), .B(n5628), .Z(out[1277]) );
  AND U5282 ( .A(n5629), .B(n5630), .Z(n5627) );
  XNOR U5283 ( .A(n5631), .B(n5632), .Z(out[1276]) );
  AND U5284 ( .A(n5633), .B(n5634), .Z(n5631) );
  XNOR U5285 ( .A(n5635), .B(n5636), .Z(out[1275]) );
  AND U5286 ( .A(n5637), .B(n5638), .Z(n5635) );
  XOR U5287 ( .A(n5639), .B(n5640), .Z(out[1274]) );
  AND U5288 ( .A(n5641), .B(n5642), .Z(n5639) );
  XOR U5289 ( .A(n5643), .B(n5644), .Z(out[1273]) );
  AND U5290 ( .A(n5645), .B(n5646), .Z(n5643) );
  XOR U5291 ( .A(n5647), .B(n5648), .Z(out[1272]) );
  AND U5292 ( .A(n5649), .B(n5650), .Z(n5647) );
  XOR U5293 ( .A(n5651), .B(n5652), .Z(out[1271]) );
  AND U5294 ( .A(n5653), .B(n5654), .Z(n5651) );
  XOR U5295 ( .A(n5655), .B(n5656), .Z(out[1270]) );
  XOR U5296 ( .A(n5659), .B(n4049), .Z(out[126]) );
  IV U5297 ( .A(n4230), .Z(n4049) );
  XOR U5298 ( .A(n5660), .B(n2402), .Z(n4230) );
  IV U5299 ( .A(n5661), .Z(n2402) );
  NOR U5300 ( .A(n2740), .B(n2738), .Z(n5659) );
  XNOR U5301 ( .A(n2236), .B(n5662), .Z(n2738) );
  IV U5302 ( .A(n5663), .Z(n2236) );
  XNOR U5303 ( .A(n5664), .B(n2648), .Z(n2740) );
  XOR U5304 ( .A(n5665), .B(n5666), .Z(out[1269]) );
  XOR U5305 ( .A(n5669), .B(n5670), .Z(out[1268]) );
  ANDN U5306 ( .B(n5671), .A(n5672), .Z(n5669) );
  XOR U5307 ( .A(n5673), .B(n5674), .Z(out[1267]) );
  XOR U5308 ( .A(n5677), .B(n5678), .Z(out[1266]) );
  XOR U5309 ( .A(n5681), .B(n5682), .Z(out[1265]) );
  XOR U5310 ( .A(n5685), .B(n5686), .Z(out[1264]) );
  AND U5311 ( .A(n5687), .B(n5688), .Z(n5685) );
  XOR U5312 ( .A(n5689), .B(n5690), .Z(out[1263]) );
  AND U5313 ( .A(n5691), .B(n5692), .Z(n5689) );
  XNOR U5314 ( .A(n5693), .B(n5694), .Z(out[1262]) );
  AND U5315 ( .A(n5695), .B(n5696), .Z(n5693) );
  XOR U5316 ( .A(n5697), .B(n5698), .Z(out[1261]) );
  AND U5317 ( .A(n5699), .B(n5700), .Z(n5697) );
  XOR U5318 ( .A(n5701), .B(n5702), .Z(out[1260]) );
  AND U5319 ( .A(n5703), .B(n5704), .Z(n5701) );
  XOR U5320 ( .A(n5705), .B(n4052), .Z(out[125]) );
  IV U5321 ( .A(n4236), .Z(n4052) );
  XOR U5322 ( .A(n5706), .B(n2409), .Z(n4236) );
  IV U5323 ( .A(n5707), .Z(n2409) );
  NOR U5324 ( .A(n2784), .B(n2782), .Z(n5705) );
  XNOR U5325 ( .A(n2243), .B(n5708), .Z(n2782) );
  IV U5326 ( .A(n5709), .Z(n2243) );
  XNOR U5327 ( .A(n5710), .B(n2655), .Z(n2784) );
  XOR U5328 ( .A(n5711), .B(n5712), .Z(out[1259]) );
  AND U5329 ( .A(n5713), .B(n5714), .Z(n5711) );
  XOR U5330 ( .A(n5715), .B(n5716), .Z(out[1258]) );
  AND U5331 ( .A(n5717), .B(n5718), .Z(n5715) );
  XOR U5332 ( .A(n5719), .B(n5720), .Z(out[1257]) );
  AND U5333 ( .A(n5721), .B(n5722), .Z(n5719) );
  XOR U5334 ( .A(n5723), .B(n5724), .Z(out[1256]) );
  AND U5335 ( .A(n5725), .B(n5726), .Z(n5723) );
  XNOR U5336 ( .A(n5727), .B(n1049), .Z(out[1255]) );
  XNOR U5337 ( .A(n5729), .B(n1053), .Z(out[1254]) );
  XNOR U5338 ( .A(n5731), .B(n1057), .Z(out[1253]) );
  AND U5339 ( .A(n5732), .B(n5733), .Z(n5731) );
  XNOR U5340 ( .A(n5734), .B(n1062), .Z(out[1252]) );
  ANDN U5341 ( .B(n5735), .A(n1061), .Z(n5734) );
  XNOR U5342 ( .A(n5736), .B(n1065), .Z(out[1251]) );
  XNOR U5343 ( .A(n5738), .B(n1069), .Z(out[1250]) );
  XOR U5344 ( .A(n5740), .B(n4055), .Z(out[124]) );
  XOR U5345 ( .A(n5741), .B(n2416), .Z(n4055) );
  IV U5346 ( .A(n5742), .Z(n2416) );
  NOR U5347 ( .A(n2828), .B(n2826), .Z(n5740) );
  XNOR U5348 ( .A(n2257), .B(n5743), .Z(n2826) );
  XNOR U5349 ( .A(n5744), .B(n2662), .Z(n2828) );
  XNOR U5350 ( .A(n5745), .B(n1073), .Z(out[1249]) );
  AND U5351 ( .A(n5746), .B(n5747), .Z(n5745) );
  XNOR U5352 ( .A(n5748), .B(n1077), .Z(out[1248]) );
  AND U5353 ( .A(n5749), .B(n5750), .Z(n5748) );
  XNOR U5354 ( .A(n5751), .B(n1081), .Z(out[1247]) );
  AND U5355 ( .A(n5752), .B(n5753), .Z(n5751) );
  XNOR U5356 ( .A(n5754), .B(n1085), .Z(out[1246]) );
  AND U5357 ( .A(n5755), .B(n5756), .Z(n5754) );
  XNOR U5358 ( .A(n5757), .B(n1093), .Z(out[1245]) );
  AND U5359 ( .A(n5758), .B(n5759), .Z(n5757) );
  XNOR U5360 ( .A(n5760), .B(n1098), .Z(out[1244]) );
  ANDN U5361 ( .B(n5761), .A(n1097), .Z(n5760) );
  XNOR U5362 ( .A(n5762), .B(n1101), .Z(out[1243]) );
  AND U5363 ( .A(n5763), .B(n5764), .Z(n5762) );
  XNOR U5364 ( .A(n5765), .B(n1105), .Z(out[1242]) );
  AND U5365 ( .A(n5766), .B(n5767), .Z(n5765) );
  XNOR U5366 ( .A(n5768), .B(n1109), .Z(out[1241]) );
  AND U5367 ( .A(n5769), .B(n5770), .Z(n5768) );
  XNOR U5368 ( .A(n5771), .B(n1114), .Z(out[1240]) );
  ANDN U5369 ( .B(n5772), .A(n1113), .Z(n5771) );
  XOR U5370 ( .A(n5773), .B(n4058), .Z(out[123]) );
  XOR U5371 ( .A(n5774), .B(n2423), .Z(n4058) );
  IV U5372 ( .A(n5775), .Z(n2423) );
  ANDN U5373 ( .B(n2873), .A(n2875), .Z(n5773) );
  XNOR U5374 ( .A(n5776), .B(n2669), .Z(n2875) );
  XNOR U5375 ( .A(n5777), .B(n2265), .Z(n2873) );
  IV U5376 ( .A(n5778), .Z(n2265) );
  XNOR U5377 ( .A(n5779), .B(n1117), .Z(out[1239]) );
  AND U5378 ( .A(n5780), .B(n5781), .Z(n5779) );
  XNOR U5379 ( .A(n5782), .B(n1122), .Z(out[1238]) );
  ANDN U5380 ( .B(n5783), .A(n1121), .Z(n5782) );
  XNOR U5381 ( .A(n5784), .B(n1126), .Z(out[1237]) );
  ANDN U5382 ( .B(n5785), .A(n1125), .Z(n5784) );
  XNOR U5383 ( .A(n5786), .B(n1130), .Z(out[1236]) );
  ANDN U5384 ( .B(n5787), .A(n1129), .Z(n5786) );
  XNOR U5385 ( .A(n5788), .B(n1137), .Z(out[1235]) );
  XNOR U5386 ( .A(n5790), .B(n1141), .Z(out[1234]) );
  AND U5387 ( .A(n5791), .B(n5792), .Z(n5790) );
  XNOR U5388 ( .A(n5793), .B(n1145), .Z(out[1233]) );
  AND U5389 ( .A(n5794), .B(n5795), .Z(n5793) );
  XNOR U5390 ( .A(n5796), .B(n1149), .Z(out[1232]) );
  AND U5391 ( .A(n5797), .B(n5798), .Z(n5796) );
  XNOR U5392 ( .A(n5799), .B(n1153), .Z(out[1231]) );
  AND U5393 ( .A(n5800), .B(n5801), .Z(n5799) );
  XNOR U5394 ( .A(n5802), .B(n1157), .Z(out[1230]) );
  AND U5395 ( .A(n5803), .B(n5804), .Z(n5802) );
  XOR U5396 ( .A(n5805), .B(n4061), .Z(out[122]) );
  IV U5397 ( .A(n4243), .Z(n4061) );
  XOR U5398 ( .A(n5806), .B(n2430), .Z(n4243) );
  ANDN U5399 ( .B(n2915), .A(n2917), .Z(n5805) );
  XNOR U5400 ( .A(n5807), .B(n2676), .Z(n2917) );
  XNOR U5401 ( .A(n5808), .B(n2272), .Z(n2915) );
  IV U5402 ( .A(n5809), .Z(n2272) );
  XNOR U5403 ( .A(n5810), .B(n1161), .Z(out[1229]) );
  AND U5404 ( .A(n5811), .B(n5812), .Z(n5810) );
  XNOR U5405 ( .A(n5813), .B(n1165), .Z(out[1228]) );
  AND U5406 ( .A(n1166), .B(n5814), .Z(n5813) );
  XNOR U5407 ( .A(n5815), .B(n1169), .Z(out[1227]) );
  AND U5408 ( .A(n1170), .B(n5816), .Z(n5815) );
  XNOR U5409 ( .A(n5817), .B(n1173), .Z(out[1226]) );
  XNOR U5410 ( .A(n5819), .B(n1181), .Z(out[1225]) );
  AND U5411 ( .A(n1182), .B(n5820), .Z(n5819) );
  XOR U5412 ( .A(n5821), .B(n1186), .Z(out[1224]) );
  ANDN U5413 ( .B(n5822), .A(n1185), .Z(n5821) );
  XOR U5414 ( .A(n5823), .B(n1190), .Z(out[1223]) );
  ANDN U5415 ( .B(n5824), .A(n1189), .Z(n5823) );
  XNOR U5416 ( .A(n5825), .B(n1193), .Z(out[1222]) );
  AND U5417 ( .A(n1194), .B(n5826), .Z(n5825) );
  XNOR U5418 ( .A(n5827), .B(n1197), .Z(out[1221]) );
  AND U5419 ( .A(n1198), .B(n5828), .Z(n5827) );
  XNOR U5420 ( .A(n5829), .B(n1201), .Z(out[1220]) );
  AND U5421 ( .A(n1202), .B(n5830), .Z(n5829) );
  XOR U5422 ( .A(n5831), .B(n4066), .Z(out[121]) );
  XOR U5423 ( .A(n5832), .B(n2437), .Z(n4066) );
  IV U5424 ( .A(n5833), .Z(n2437) );
  ANDN U5425 ( .B(n2955), .A(n2957), .Z(n5831) );
  XNOR U5426 ( .A(n5834), .B(n2683), .Z(n2957) );
  XOR U5427 ( .A(n5835), .B(n2279), .Z(n2955) );
  IV U5428 ( .A(n5836), .Z(n2279) );
  XNOR U5429 ( .A(n5837), .B(n1205), .Z(out[1219]) );
  AND U5430 ( .A(n1206), .B(n5838), .Z(n5837) );
  XNOR U5431 ( .A(n5839), .B(n1209), .Z(out[1218]) );
  AND U5432 ( .A(n1210), .B(n5840), .Z(n5839) );
  XNOR U5433 ( .A(n5841), .B(n1213), .Z(out[1217]) );
  AND U5434 ( .A(n5842), .B(n5843), .Z(n5841) );
  XNOR U5435 ( .A(n5844), .B(n1217), .Z(out[1216]) );
  AND U5436 ( .A(n1218), .B(n5845), .Z(n5844) );
  XOR U5437 ( .A(n5846), .B(n5622), .Z(out[1215]) );
  ANDN U5438 ( .B(n5847), .A(n5621), .Z(n5846) );
  XOR U5439 ( .A(n5848), .B(n5626), .Z(out[1214]) );
  ANDN U5440 ( .B(n5849), .A(n5625), .Z(n5848) );
  XNOR U5441 ( .A(n5850), .B(n5629), .Z(out[1213]) );
  AND U5442 ( .A(n5851), .B(n5852), .Z(n5850) );
  XNOR U5443 ( .A(n5853), .B(n5633), .Z(out[1212]) );
  AND U5444 ( .A(n5854), .B(n5855), .Z(n5853) );
  XNOR U5445 ( .A(n5856), .B(n5637), .Z(out[1211]) );
  AND U5446 ( .A(n5857), .B(n5858), .Z(n5856) );
  XNOR U5447 ( .A(n5859), .B(n5641), .Z(out[1210]) );
  AND U5448 ( .A(n5860), .B(n5861), .Z(n5859) );
  XOR U5449 ( .A(n5862), .B(n4069), .Z(out[120]) );
  XOR U5450 ( .A(n5863), .B(n2444), .Z(n4069) );
  IV U5451 ( .A(n5864), .Z(n2444) );
  ANDN U5452 ( .B(n2987), .A(n2989), .Z(n5862) );
  XNOR U5453 ( .A(n5865), .B(n2690), .Z(n2989) );
  XNOR U5454 ( .A(n5866), .B(n2286), .Z(n2987) );
  IV U5455 ( .A(n5867), .Z(n2286) );
  XNOR U5456 ( .A(n5868), .B(n5646), .Z(out[1209]) );
  ANDN U5457 ( .B(n5869), .A(n5645), .Z(n5868) );
  XNOR U5458 ( .A(n5870), .B(n5649), .Z(out[1208]) );
  AND U5459 ( .A(n5871), .B(n5872), .Z(n5870) );
  XNOR U5460 ( .A(n5873), .B(n5653), .Z(out[1207]) );
  AND U5461 ( .A(n5874), .B(n5875), .Z(n5873) );
  XOR U5462 ( .A(n5876), .B(n5658), .Z(out[1206]) );
  ANDN U5463 ( .B(n5877), .A(n5657), .Z(n5876) );
  XOR U5464 ( .A(n5878), .B(n5668), .Z(out[1205]) );
  ANDN U5465 ( .B(n5879), .A(n5667), .Z(n5878) );
  XOR U5466 ( .A(n5880), .B(n5672), .Z(out[1204]) );
  AND U5467 ( .A(n5881), .B(n5882), .Z(n5880) );
  XOR U5468 ( .A(n5883), .B(n5676), .Z(out[1203]) );
  ANDN U5469 ( .B(n5884), .A(n5675), .Z(n5883) );
  XOR U5470 ( .A(n5885), .B(n5680), .Z(out[1202]) );
  ANDN U5471 ( .B(n5886), .A(n5679), .Z(n5885) );
  XOR U5472 ( .A(n5887), .B(n5684), .Z(out[1201]) );
  ANDN U5473 ( .B(n5888), .A(n5683), .Z(n5887) );
  XNOR U5474 ( .A(n5889), .B(n5687), .Z(out[1200]) );
  AND U5475 ( .A(n5890), .B(n5891), .Z(n5889) );
  XOR U5476 ( .A(n5892), .B(n2002), .Z(out[11]) );
  XOR U5477 ( .A(n5893), .B(n2617), .Z(n2002) );
  IV U5478 ( .A(n5894), .Z(n2617) );
  NOR U5479 ( .A(n4003), .B(n2001), .Z(n5892) );
  XNOR U5480 ( .A(n2551), .B(n5895), .Z(n2001) );
  XOR U5481 ( .A(n5896), .B(n1752), .Z(n4003) );
  XOR U5482 ( .A(n5897), .B(n4072), .Z(out[119]) );
  XOR U5483 ( .A(n5898), .B(n2451), .Z(n4072) );
  IV U5484 ( .A(n5899), .Z(n2451) );
  ANDN U5485 ( .B(n3019), .A(n3021), .Z(n5897) );
  XOR U5486 ( .A(n5900), .B(n2221), .Z(n3021) );
  IV U5487 ( .A(n4925), .Z(n2221) );
  XNOR U5488 ( .A(n5901), .B(n2293), .Z(n3019) );
  IV U5489 ( .A(n5902), .Z(n2293) );
  XNOR U5490 ( .A(n5903), .B(n5691), .Z(out[1199]) );
  AND U5491 ( .A(n5904), .B(n5905), .Z(n5903) );
  XNOR U5492 ( .A(n5906), .B(n5696), .Z(out[1198]) );
  ANDN U5493 ( .B(n5907), .A(n5695), .Z(n5906) );
  XNOR U5494 ( .A(n5908), .B(n5700), .Z(out[1197]) );
  ANDN U5495 ( .B(n5909), .A(n5699), .Z(n5908) );
  XNOR U5496 ( .A(n5910), .B(n5704), .Z(out[1196]) );
  ANDN U5497 ( .B(n5911), .A(n5703), .Z(n5910) );
  XNOR U5498 ( .A(n5912), .B(n5714), .Z(out[1195]) );
  ANDN U5499 ( .B(n5913), .A(n5713), .Z(n5912) );
  XNOR U5500 ( .A(n5914), .B(n5718), .Z(out[1194]) );
  ANDN U5501 ( .B(n5915), .A(n5717), .Z(n5914) );
  XNOR U5502 ( .A(n5916), .B(n5722), .Z(out[1193]) );
  ANDN U5503 ( .B(n5917), .A(n5721), .Z(n5916) );
  XNOR U5504 ( .A(n5918), .B(n5726), .Z(out[1192]) );
  ANDN U5505 ( .B(n5919), .A(n5725), .Z(n5918) );
  XOR U5506 ( .A(n5920), .B(n1050), .Z(out[1191]) );
  XOR U5507 ( .A(n2114), .B(n5921), .Z(n1050) );
  IV U5508 ( .A(n5446), .Z(n2114) );
  XOR U5509 ( .A(n5922), .B(n5923), .Z(n5446) );
  NOR U5510 ( .A(n5924), .B(n5728), .Z(n5920) );
  XOR U5511 ( .A(n5925), .B(n1054), .Z(out[1190]) );
  XOR U5512 ( .A(n2118), .B(n5926), .Z(n1054) );
  IV U5513 ( .A(n5452), .Z(n2118) );
  XOR U5514 ( .A(n5927), .B(n5928), .Z(n5452) );
  ANDN U5515 ( .B(n5929), .A(n5730), .Z(n5925) );
  XNOR U5516 ( .A(n5930), .B(n4075), .Z(out[118]) );
  XNOR U5517 ( .A(n5931), .B(n2458), .Z(n4075) );
  IV U5518 ( .A(n5932), .Z(n2458) );
  ANDN U5519 ( .B(n3048), .A(n3050), .Z(n5930) );
  XOR U5520 ( .A(n5933), .B(n2228), .Z(n3050) );
  IV U5521 ( .A(n3555), .Z(n2228) );
  XNOR U5522 ( .A(n5934), .B(n2300), .Z(n3048) );
  IV U5523 ( .A(n5935), .Z(n2300) );
  XOR U5524 ( .A(n5936), .B(n1058), .Z(out[1189]) );
  IV U5525 ( .A(n5733), .Z(n1058) );
  XNOR U5526 ( .A(n5937), .B(n2125), .Z(n5733) );
  XOR U5527 ( .A(n5938), .B(n5939), .Z(n2125) );
  ANDN U5528 ( .B(n5940), .A(n5732), .Z(n5936) );
  XOR U5529 ( .A(n5941), .B(n1061), .Z(out[1188]) );
  XOR U5530 ( .A(n5943), .B(n5944), .Z(n2127) );
  ANDN U5531 ( .B(n5945), .A(n5735), .Z(n5941) );
  XOR U5532 ( .A(n5946), .B(n1066), .Z(out[1187]) );
  XOR U5533 ( .A(n2131), .B(n5947), .Z(n1066) );
  IV U5534 ( .A(n5471), .Z(n2131) );
  XOR U5535 ( .A(n5948), .B(n5949), .Z(n5471) );
  ANDN U5536 ( .B(n5950), .A(n5737), .Z(n5946) );
  XOR U5537 ( .A(n5951), .B(n1070), .Z(out[1186]) );
  XOR U5538 ( .A(n2135), .B(n5952), .Z(n1070) );
  IV U5539 ( .A(n5477), .Z(n2135) );
  XOR U5540 ( .A(n5953), .B(n5954), .Z(n5477) );
  ANDN U5541 ( .B(n5955), .A(n5739), .Z(n5951) );
  XOR U5542 ( .A(n5956), .B(n1074), .Z(out[1185]) );
  IV U5543 ( .A(n5747), .Z(n1074) );
  XNOR U5544 ( .A(n2139), .B(n5957), .Z(n5747) );
  XOR U5545 ( .A(n5958), .B(n5959), .Z(n2139) );
  ANDN U5546 ( .B(n5960), .A(n5746), .Z(n5956) );
  XOR U5547 ( .A(n5961), .B(n1078), .Z(out[1184]) );
  IV U5548 ( .A(n5750), .Z(n1078) );
  XNOR U5549 ( .A(n2143), .B(n5962), .Z(n5750) );
  XOR U5550 ( .A(n5963), .B(n5964), .Z(n2143) );
  ANDN U5551 ( .B(n5965), .A(n5749), .Z(n5961) );
  XOR U5552 ( .A(n5966), .B(n1082), .Z(out[1183]) );
  IV U5553 ( .A(n5753), .Z(n1082) );
  XNOR U5554 ( .A(n2147), .B(n5967), .Z(n5753) );
  XOR U5555 ( .A(n5968), .B(n5969), .Z(n2147) );
  ANDN U5556 ( .B(n5970), .A(n5752), .Z(n5966) );
  XOR U5557 ( .A(n5971), .B(n1086), .Z(out[1182]) );
  IV U5558 ( .A(n5756), .Z(n1086) );
  XOR U5559 ( .A(n5972), .B(n2152), .Z(n5756) );
  XNOR U5560 ( .A(n5973), .B(n5974), .Z(n2152) );
  ANDN U5561 ( .B(n5975), .A(n5755), .Z(n5971) );
  XOR U5562 ( .A(n5976), .B(n1094), .Z(out[1181]) );
  IV U5563 ( .A(n5759), .Z(n1094) );
  XNOR U5564 ( .A(n5977), .B(n2155), .Z(n5759) );
  XNOR U5565 ( .A(n5978), .B(n5979), .Z(n2155) );
  ANDN U5566 ( .B(n5980), .A(n5758), .Z(n5976) );
  XOR U5567 ( .A(n5981), .B(n1097), .Z(out[1180]) );
  XOR U5568 ( .A(n5982), .B(n2159), .Z(n1097) );
  XNOR U5569 ( .A(n5983), .B(n5984), .Z(n2159) );
  ANDN U5570 ( .B(n5985), .A(n5761), .Z(n5981) );
  XNOR U5571 ( .A(n5986), .B(n4078), .Z(out[117]) );
  XNOR U5572 ( .A(n5987), .B(n2465), .Z(n4078) );
  IV U5573 ( .A(n5558), .Z(n2465) );
  ANDN U5574 ( .B(n3079), .A(n3081), .Z(n5986) );
  XOR U5575 ( .A(n5988), .B(n2235), .Z(n3081) );
  IV U5576 ( .A(n3558), .Z(n2235) );
  XNOR U5577 ( .A(n5989), .B(n2307), .Z(n3079) );
  IV U5578 ( .A(n5990), .Z(n2307) );
  XOR U5579 ( .A(n5991), .B(n1102), .Z(out[1179]) );
  IV U5580 ( .A(n5764), .Z(n1102) );
  XNOR U5581 ( .A(n5992), .B(n2164), .Z(n5764) );
  XNOR U5582 ( .A(n5993), .B(n5994), .Z(n2164) );
  ANDN U5583 ( .B(n5995), .A(n5763), .Z(n5991) );
  XOR U5584 ( .A(n5996), .B(n1106), .Z(out[1178]) );
  IV U5585 ( .A(n5767), .Z(n1106) );
  XNOR U5586 ( .A(n5997), .B(n2168), .Z(n5767) );
  XNOR U5587 ( .A(n5998), .B(n5999), .Z(n2168) );
  ANDN U5588 ( .B(n6000), .A(n5766), .Z(n5996) );
  XOR U5589 ( .A(n6001), .B(n1110), .Z(out[1177]) );
  IV U5590 ( .A(n5770), .Z(n1110) );
  XNOR U5591 ( .A(n6002), .B(n2172), .Z(n5770) );
  XNOR U5592 ( .A(n6003), .B(n6004), .Z(n2172) );
  ANDN U5593 ( .B(n6005), .A(n5769), .Z(n6001) );
  XOR U5594 ( .A(n6006), .B(n1113), .Z(out[1176]) );
  XNOR U5595 ( .A(n6007), .B(n2175), .Z(n1113) );
  XNOR U5596 ( .A(n6008), .B(n6009), .Z(n2175) );
  ANDN U5597 ( .B(n6010), .A(n5772), .Z(n6006) );
  XOR U5598 ( .A(n6011), .B(n1118), .Z(out[1175]) );
  IV U5599 ( .A(n5781), .Z(n1118) );
  XNOR U5600 ( .A(n6012), .B(n2178), .Z(n5781) );
  XNOR U5601 ( .A(n6013), .B(n6014), .Z(n2178) );
  ANDN U5602 ( .B(n6015), .A(n5780), .Z(n6011) );
  XOR U5603 ( .A(n6016), .B(n1121), .Z(out[1174]) );
  XOR U5604 ( .A(n6017), .B(n2181), .Z(n1121) );
  XOR U5605 ( .A(n6018), .B(n6019), .Z(n2181) );
  ANDN U5606 ( .B(n6020), .A(n5783), .Z(n6016) );
  XOR U5607 ( .A(n6021), .B(n1125), .Z(out[1173]) );
  XNOR U5608 ( .A(n6022), .B(n4295), .Z(n1125) );
  XNOR U5609 ( .A(n6023), .B(n6024), .Z(n4295) );
  ANDN U5610 ( .B(n6025), .A(n5785), .Z(n6021) );
  XOR U5611 ( .A(n6026), .B(n1129), .Z(out[1172]) );
  XOR U5612 ( .A(n6027), .B(n2188), .Z(n1129) );
  XOR U5613 ( .A(n6028), .B(n6029), .Z(n2188) );
  AND U5614 ( .A(n6030), .B(n6031), .Z(n6026) );
  XOR U5615 ( .A(n6032), .B(n1138), .Z(out[1171]) );
  XNOR U5616 ( .A(n6033), .B(n2191), .Z(n1138) );
  ANDN U5617 ( .B(n6036), .A(n5789), .Z(n6032) );
  XOR U5618 ( .A(n6037), .B(n1142), .Z(out[1170]) );
  IV U5619 ( .A(n5792), .Z(n1142) );
  XNOR U5620 ( .A(n6038), .B(n2194), .Z(n5792) );
  XNOR U5621 ( .A(n6039), .B(n6040), .Z(n2194) );
  ANDN U5622 ( .B(n6041), .A(n5791), .Z(n6037) );
  XOR U5623 ( .A(n6042), .B(n4081), .Z(out[116]) );
  XOR U5624 ( .A(n6043), .B(n2476), .Z(n4081) );
  IV U5625 ( .A(n6044), .Z(n2476) );
  ANDN U5626 ( .B(n3107), .A(n3109), .Z(n6042) );
  XNOR U5627 ( .A(n6045), .B(n2242), .Z(n3109) );
  IV U5628 ( .A(n6046), .Z(n2242) );
  XNOR U5629 ( .A(n6047), .B(n2314), .Z(n3107) );
  IV U5630 ( .A(n6048), .Z(n2314) );
  XOR U5631 ( .A(n6049), .B(n1146), .Z(out[1169]) );
  IV U5632 ( .A(n5795), .Z(n1146) );
  XNOR U5633 ( .A(n6050), .B(n2201), .Z(n5795) );
  XNOR U5634 ( .A(n6051), .B(n6052), .Z(n2201) );
  ANDN U5635 ( .B(n6053), .A(n5794), .Z(n6049) );
  XOR U5636 ( .A(n6054), .B(n1150), .Z(out[1168]) );
  IV U5637 ( .A(n5798), .Z(n1150) );
  XNOR U5638 ( .A(n6055), .B(n2204), .Z(n5798) );
  XNOR U5639 ( .A(n6056), .B(n6057), .Z(n2204) );
  ANDN U5640 ( .B(n6058), .A(n5797), .Z(n6054) );
  XOR U5641 ( .A(n6059), .B(n1154), .Z(out[1167]) );
  IV U5642 ( .A(n5801), .Z(n1154) );
  XNOR U5643 ( .A(n6060), .B(n2207), .Z(n5801) );
  XNOR U5644 ( .A(n6061), .B(n6062), .Z(n2207) );
  ANDN U5645 ( .B(n6063), .A(n5800), .Z(n6059) );
  XOR U5646 ( .A(n6064), .B(n1158), .Z(out[1166]) );
  IV U5647 ( .A(n5804), .Z(n1158) );
  XNOR U5648 ( .A(n6065), .B(n2210), .Z(n5804) );
  XNOR U5649 ( .A(n6066), .B(n6067), .Z(n2210) );
  NOR U5650 ( .A(n6068), .B(n5803), .Z(n6064) );
  XOR U5651 ( .A(n6069), .B(n1162), .Z(out[1165]) );
  IV U5652 ( .A(n5812), .Z(n1162) );
  XNOR U5653 ( .A(n6070), .B(n2213), .Z(n5812) );
  XNOR U5654 ( .A(n6071), .B(n6072), .Z(n2213) );
  ANDN U5655 ( .B(n6073), .A(n5811), .Z(n6069) );
  XNOR U5656 ( .A(n6074), .B(n1166), .Z(out[1164]) );
  XNOR U5657 ( .A(n6075), .B(n2216), .Z(n1166) );
  IV U5658 ( .A(n5585), .Z(n2216) );
  AND U5659 ( .A(n6078), .B(n6079), .Z(n6074) );
  XNOR U5660 ( .A(n6080), .B(n1170), .Z(out[1163]) );
  XNOR U5661 ( .A(n6081), .B(n1976), .Z(n1170) );
  IV U5662 ( .A(n5590), .Z(n1976) );
  AND U5663 ( .A(n6084), .B(n6085), .Z(n6080) );
  XOR U5664 ( .A(n6086), .B(n1174), .Z(out[1162]) );
  XOR U5665 ( .A(n6087), .B(n1979), .Z(n1174) );
  IV U5666 ( .A(n5595), .Z(n1979) );
  ANDN U5667 ( .B(n6090), .A(n5818), .Z(n6086) );
  XNOR U5668 ( .A(n6091), .B(n1182), .Z(out[1161]) );
  XNOR U5669 ( .A(n6092), .B(n1982), .Z(n1182) );
  IV U5670 ( .A(n5600), .Z(n1982) );
  AND U5671 ( .A(n6095), .B(n6096), .Z(n6091) );
  XOR U5672 ( .A(n6097), .B(n1185), .Z(out[1160]) );
  XOR U5673 ( .A(n6098), .B(n1985), .Z(n1185) );
  XNOR U5674 ( .A(n6099), .B(n6100), .Z(n1985) );
  ANDN U5675 ( .B(n6101), .A(n5822), .Z(n6097) );
  XOR U5676 ( .A(n6102), .B(n4085), .Z(out[115]) );
  XOR U5677 ( .A(n6103), .B(n2483), .Z(n4085) );
  ANDN U5678 ( .B(n3131), .A(n3133), .Z(n6102) );
  XNOR U5679 ( .A(n6104), .B(n2256), .Z(n3133) );
  IV U5680 ( .A(n6105), .Z(n2256) );
  XOR U5681 ( .A(n6106), .B(n2321), .Z(n3131) );
  IV U5682 ( .A(n6107), .Z(n2321) );
  XOR U5683 ( .A(n6108), .B(n1189), .Z(out[1159]) );
  XOR U5684 ( .A(n6109), .B(n1988), .Z(n1189) );
  XNOR U5685 ( .A(n6110), .B(n6111), .Z(n1988) );
  ANDN U5686 ( .B(n6112), .A(n5824), .Z(n6108) );
  XNOR U5687 ( .A(n6113), .B(n1194), .Z(out[1158]) );
  XNOR U5688 ( .A(n6114), .B(n1992), .Z(n1194) );
  XNOR U5689 ( .A(n6115), .B(n6116), .Z(n1992) );
  AND U5690 ( .A(n6117), .B(n6118), .Z(n6113) );
  XNOR U5691 ( .A(n6119), .B(n1198), .Z(out[1157]) );
  XNOR U5692 ( .A(n6120), .B(n1995), .Z(n1198) );
  XNOR U5693 ( .A(n6121), .B(n6122), .Z(n1995) );
  AND U5694 ( .A(n6123), .B(n6124), .Z(n6119) );
  XNOR U5695 ( .A(n6125), .B(n1202), .Z(out[1156]) );
  XNOR U5696 ( .A(n6126), .B(n1998), .Z(n1202) );
  XNOR U5697 ( .A(n6127), .B(n6128), .Z(n1998) );
  AND U5698 ( .A(n6129), .B(n6130), .Z(n6125) );
  XNOR U5699 ( .A(n6131), .B(n1206), .Z(out[1155]) );
  XNOR U5700 ( .A(n6132), .B(n2005), .Z(n1206) );
  XNOR U5701 ( .A(n6133), .B(n6134), .Z(n2005) );
  AND U5702 ( .A(n6135), .B(n6136), .Z(n6131) );
  XNOR U5703 ( .A(n6137), .B(n1210), .Z(out[1154]) );
  XNOR U5704 ( .A(n6138), .B(n2009), .Z(n1210) );
  XNOR U5705 ( .A(n6139), .B(n6140), .Z(n2009) );
  AND U5706 ( .A(n6141), .B(n6142), .Z(n6137) );
  XOR U5707 ( .A(n6143), .B(n1214), .Z(out[1153]) );
  IV U5708 ( .A(n5843), .Z(n1214) );
  XNOR U5709 ( .A(n6144), .B(n2013), .Z(n5843) );
  XNOR U5710 ( .A(n6145), .B(n6146), .Z(n2013) );
  ANDN U5711 ( .B(n6147), .A(n5842), .Z(n6143) );
  XNOR U5712 ( .A(n6148), .B(n1218), .Z(out[1152]) );
  XNOR U5713 ( .A(n6149), .B(n2017), .Z(n1218) );
  XNOR U5714 ( .A(n6150), .B(n6151), .Z(n2017) );
  AND U5715 ( .A(n6152), .B(n6153), .Z(n6148) );
  XOR U5716 ( .A(n6154), .B(n5621), .Z(out[1151]) );
  XNOR U5717 ( .A(n6155), .B(n2585), .Z(n5621) );
  ANDN U5718 ( .B(n6156), .A(n5847), .Z(n6154) );
  XOR U5719 ( .A(n6157), .B(n5625), .Z(out[1150]) );
  XNOR U5720 ( .A(n6158), .B(n2592), .Z(n5625) );
  ANDN U5721 ( .B(n6159), .A(n5849), .Z(n6157) );
  XOR U5722 ( .A(n6160), .B(n4089), .Z(out[114]) );
  XNOR U5723 ( .A(n6161), .B(n2490), .Z(n4089) );
  ANDN U5724 ( .B(n3159), .A(n3161), .Z(n6160) );
  XNOR U5725 ( .A(n6162), .B(n2263), .Z(n3161) );
  XOR U5726 ( .A(n6163), .B(n2332), .Z(n3159) );
  IV U5727 ( .A(n6164), .Z(n2332) );
  XOR U5728 ( .A(n6165), .B(n5630), .Z(out[1149]) );
  IV U5729 ( .A(n5852), .Z(n5630) );
  XOR U5730 ( .A(n5323), .B(n6166), .Z(n5852) );
  XOR U5731 ( .A(n6167), .B(n6168), .Z(n5323) );
  ANDN U5732 ( .B(n6169), .A(n5851), .Z(n6165) );
  XOR U5733 ( .A(n6170), .B(n5634), .Z(out[1148]) );
  IV U5734 ( .A(n5855), .Z(n5634) );
  XOR U5735 ( .A(n5330), .B(n6171), .Z(n5855) );
  XOR U5736 ( .A(n6172), .B(n6173), .Z(n5330) );
  ANDN U5737 ( .B(n6174), .A(n5854), .Z(n6170) );
  XOR U5738 ( .A(n6175), .B(n5638), .Z(out[1147]) );
  IV U5739 ( .A(n5858), .Z(n5638) );
  XOR U5740 ( .A(n4319), .B(n6176), .Z(n5858) );
  XOR U5741 ( .A(n6177), .B(n6178), .Z(n4319) );
  ANDN U5742 ( .B(n6179), .A(n5857), .Z(n6175) );
  XOR U5743 ( .A(n6180), .B(n5642), .Z(out[1146]) );
  IV U5744 ( .A(n5861), .Z(n5642) );
  XOR U5745 ( .A(n6181), .B(n2625), .Z(n5861) );
  XOR U5746 ( .A(n6182), .B(n6183), .Z(n2625) );
  ANDN U5747 ( .B(n6184), .A(n5860), .Z(n6180) );
  XOR U5748 ( .A(n6185), .B(n5645), .Z(out[1145]) );
  XOR U5749 ( .A(n6186), .B(n2632), .Z(n5645) );
  IV U5750 ( .A(n3742), .Z(n2632) );
  XNOR U5751 ( .A(n6187), .B(n6188), .Z(n3742) );
  ANDN U5752 ( .B(n6189), .A(n5869), .Z(n6185) );
  XOR U5753 ( .A(n6190), .B(n5650), .Z(out[1144]) );
  IV U5754 ( .A(n5872), .Z(n5650) );
  XOR U5755 ( .A(n6191), .B(n2639), .Z(n5872) );
  XNOR U5756 ( .A(n6192), .B(n6193), .Z(n2639) );
  ANDN U5757 ( .B(n6194), .A(n5871), .Z(n6190) );
  XOR U5758 ( .A(n6195), .B(n5654), .Z(out[1143]) );
  IV U5759 ( .A(n5875), .Z(n5654) );
  XOR U5760 ( .A(n6196), .B(n2646), .Z(n5875) );
  XNOR U5761 ( .A(n6197), .B(n6198), .Z(n2646) );
  ANDN U5762 ( .B(n6199), .A(n5874), .Z(n6195) );
  XOR U5763 ( .A(n6200), .B(n5657), .Z(out[1142]) );
  XNOR U5764 ( .A(n6201), .B(n2653), .Z(n5657) );
  XNOR U5765 ( .A(n6202), .B(n6203), .Z(n2653) );
  ANDN U5766 ( .B(n6204), .A(n5877), .Z(n6200) );
  XOR U5767 ( .A(n6205), .B(n5667), .Z(out[1141]) );
  XNOR U5768 ( .A(n6206), .B(n2660), .Z(n5667) );
  XNOR U5769 ( .A(n6207), .B(n6208), .Z(n2660) );
  ANDN U5770 ( .B(n6209), .A(n5879), .Z(n6205) );
  XOR U5771 ( .A(n6210), .B(n5671), .Z(out[1140]) );
  IV U5772 ( .A(n5882), .Z(n5671) );
  XOR U5773 ( .A(n6211), .B(n2667), .Z(n5882) );
  XNOR U5774 ( .A(n6212), .B(n6213), .Z(n2667) );
  ANDN U5775 ( .B(n6214), .A(n5881), .Z(n6210) );
  XOR U5776 ( .A(n6215), .B(n4093), .Z(out[113]) );
  IV U5777 ( .A(n4265), .Z(n4093) );
  XOR U5778 ( .A(n6216), .B(n2497), .Z(n4265) );
  ANDN U5779 ( .B(n3200), .A(n3202), .Z(n6215) );
  XNOR U5780 ( .A(n6217), .B(n2270), .Z(n3202) );
  XNOR U5781 ( .A(n6218), .B(n2337), .Z(n3200) );
  IV U5782 ( .A(n6219), .Z(n2337) );
  XOR U5783 ( .A(n6220), .B(n5675), .Z(out[1139]) );
  XNOR U5784 ( .A(n6221), .B(n2674), .Z(n5675) );
  XNOR U5785 ( .A(n6222), .B(n6223), .Z(n2674) );
  ANDN U5786 ( .B(n6224), .A(n5884), .Z(n6220) );
  XOR U5787 ( .A(n6225), .B(n5679), .Z(out[1138]) );
  XNOR U5788 ( .A(n6226), .B(n2681), .Z(n5679) );
  XNOR U5789 ( .A(n6227), .B(n6228), .Z(n2681) );
  ANDN U5790 ( .B(n6229), .A(n5886), .Z(n6225) );
  XOR U5791 ( .A(n6230), .B(n5683), .Z(out[1137]) );
  XNOR U5792 ( .A(n6231), .B(n2688), .Z(n5683) );
  XNOR U5793 ( .A(n6232), .B(n6233), .Z(n2688) );
  ANDN U5794 ( .B(n6234), .A(n5888), .Z(n6230) );
  XOR U5795 ( .A(n6235), .B(n5688), .Z(out[1136]) );
  IV U5796 ( .A(n5891), .Z(n5688) );
  XOR U5797 ( .A(n6236), .B(n2219), .Z(n5891) );
  XNOR U5798 ( .A(n6237), .B(n6238), .Z(n2219) );
  XOR U5799 ( .A(n6240), .B(n5692), .Z(out[1135]) );
  IV U5800 ( .A(n5905), .Z(n5692) );
  XOR U5801 ( .A(n6241), .B(n2226), .Z(n5905) );
  XNOR U5802 ( .A(n6242), .B(n6243), .Z(n2226) );
  ANDN U5803 ( .B(n6244), .A(n5904), .Z(n6240) );
  XOR U5804 ( .A(n6245), .B(n5695), .Z(out[1134]) );
  XOR U5805 ( .A(n6246), .B(n4778), .Z(n5695) );
  XOR U5806 ( .A(n6247), .B(n6248), .Z(n4778) );
  XOR U5807 ( .A(n6250), .B(n5699), .Z(out[1133]) );
  XNOR U5808 ( .A(n6251), .B(n4803), .Z(n5699) );
  XOR U5809 ( .A(n6252), .B(n6253), .Z(n4803) );
  XOR U5810 ( .A(n6255), .B(n5703), .Z(out[1132]) );
  XNOR U5811 ( .A(n6256), .B(n4833), .Z(n5703) );
  XOR U5812 ( .A(n6257), .B(n6258), .Z(n4833) );
  XOR U5813 ( .A(n6260), .B(n5713), .Z(out[1131]) );
  XNOR U5814 ( .A(n6261), .B(n3802), .Z(n5713) );
  XOR U5815 ( .A(n6262), .B(n6263), .Z(n3802) );
  AND U5816 ( .A(n6264), .B(n6265), .Z(n6260) );
  XOR U5817 ( .A(n6266), .B(n5717), .Z(out[1130]) );
  XOR U5818 ( .A(n6267), .B(n4905), .Z(n5717) );
  XOR U5819 ( .A(n6268), .B(n6269), .Z(n4905) );
  AND U5820 ( .A(n6270), .B(n6271), .Z(n6266) );
  XOR U5821 ( .A(n6272), .B(n4096), .Z(out[112]) );
  IV U5822 ( .A(n4268), .Z(n4096) );
  XNOR U5823 ( .A(n6273), .B(n2504), .Z(n4268) );
  ANDN U5824 ( .B(n3234), .A(n3236), .Z(n6272) );
  XNOR U5825 ( .A(n6274), .B(n2277), .Z(n3236) );
  XOR U5826 ( .A(n6275), .B(n2344), .Z(n3234) );
  IV U5827 ( .A(n6276), .Z(n2344) );
  XOR U5828 ( .A(n6277), .B(n5721), .Z(out[1129]) );
  XNOR U5829 ( .A(n6278), .B(n4947), .Z(n5721) );
  XOR U5830 ( .A(n6279), .B(n6280), .Z(n4947) );
  XOR U5831 ( .A(n6282), .B(n5725), .Z(out[1128]) );
  XOR U5832 ( .A(n6283), .B(n4982), .Z(n5725) );
  XOR U5833 ( .A(n6284), .B(n6285), .Z(n4982) );
  XOR U5834 ( .A(n6287), .B(n5728), .Z(out[1127]) );
  XNOR U5835 ( .A(n6288), .B(n5436), .Z(n5728) );
  XOR U5836 ( .A(n6289), .B(n6290), .Z(n5436) );
  ANDN U5837 ( .B(n5924), .A(n1048), .Z(n6287) );
  XOR U5838 ( .A(n6291), .B(n5730), .Z(out[1126]) );
  XOR U5839 ( .A(n6292), .B(n5080), .Z(n5730) );
  XOR U5840 ( .A(n6293), .B(n6294), .Z(n5080) );
  NOR U5841 ( .A(n1052), .B(n5929), .Z(n6291) );
  XOR U5842 ( .A(n6295), .B(n5732), .Z(out[1125]) );
  XNOR U5843 ( .A(n6296), .B(n5114), .Z(n5732) );
  XOR U5844 ( .A(n6297), .B(n6298), .Z(n5114) );
  NOR U5845 ( .A(n1056), .B(n5940), .Z(n6295) );
  XOR U5846 ( .A(n6299), .B(n5735), .Z(out[1124]) );
  XNOR U5847 ( .A(n6300), .B(n5450), .Z(n5735) );
  XOR U5848 ( .A(n6301), .B(n6302), .Z(n5450) );
  NOR U5849 ( .A(n1060), .B(n5945), .Z(n6299) );
  XOR U5850 ( .A(n6303), .B(n5737), .Z(out[1123]) );
  XNOR U5851 ( .A(n6304), .B(n5456), .Z(n5737) );
  XOR U5852 ( .A(n6305), .B(n6306), .Z(n5456) );
  NOR U5853 ( .A(n1064), .B(n5950), .Z(n6303) );
  XOR U5854 ( .A(n6307), .B(n5739), .Z(out[1122]) );
  XNOR U5855 ( .A(n6308), .B(n5207), .Z(n5739) );
  XOR U5856 ( .A(n6309), .B(n6310), .Z(n5207) );
  NOR U5857 ( .A(n1068), .B(n5955), .Z(n6307) );
  XOR U5858 ( .A(n6311), .B(n5746), .Z(out[1121]) );
  XNOR U5859 ( .A(n6312), .B(n5465), .Z(n5746) );
  XOR U5860 ( .A(n6313), .B(n6314), .Z(n5465) );
  NOR U5861 ( .A(n1072), .B(n5960), .Z(n6311) );
  XOR U5862 ( .A(n6315), .B(n5749), .Z(out[1120]) );
  XNOR U5863 ( .A(n6316), .B(n5475), .Z(n5749) );
  XOR U5864 ( .A(n6317), .B(n6318), .Z(n5475) );
  ANDN U5865 ( .B(n1076), .A(n5965), .Z(n6315) );
  XOR U5866 ( .A(n6319), .B(n4101), .Z(out[111]) );
  IV U5867 ( .A(n4271), .Z(n4101) );
  XOR U5868 ( .A(n6320), .B(n2511), .Z(n4271) );
  ANDN U5869 ( .B(n3269), .A(n3270), .Z(n6319) );
  XNOR U5870 ( .A(n6321), .B(n2284), .Z(n3270) );
  XOR U5871 ( .A(n6322), .B(n2351), .Z(n3269) );
  XOR U5872 ( .A(n6323), .B(n5752), .Z(out[1119]) );
  XOR U5873 ( .A(n6324), .B(n5481), .Z(n5752) );
  XOR U5874 ( .A(n6325), .B(n6326), .Z(n5481) );
  NOR U5875 ( .A(n1080), .B(n5970), .Z(n6323) );
  XOR U5876 ( .A(n6327), .B(n5755), .Z(out[1118]) );
  XOR U5877 ( .A(n6328), .B(n5486), .Z(n5755) );
  XOR U5878 ( .A(n6329), .B(n6330), .Z(n5486) );
  NOR U5879 ( .A(n1084), .B(n5975), .Z(n6327) );
  XOR U5880 ( .A(n6331), .B(n5758), .Z(out[1117]) );
  XOR U5881 ( .A(n6332), .B(n5491), .Z(n5758) );
  XOR U5882 ( .A(n6333), .B(n6334), .Z(n5491) );
  NOR U5883 ( .A(n1092), .B(n5980), .Z(n6331) );
  XOR U5884 ( .A(n6335), .B(n5761), .Z(out[1116]) );
  XOR U5885 ( .A(n6336), .B(n3586), .Z(n5761) );
  XOR U5886 ( .A(n6337), .B(n6338), .Z(n3586) );
  NOR U5887 ( .A(n1096), .B(n5985), .Z(n6335) );
  XOR U5888 ( .A(n6339), .B(n5763), .Z(out[1115]) );
  XNOR U5889 ( .A(n6340), .B(n3591), .Z(n5763) );
  XOR U5890 ( .A(n6341), .B(n6342), .Z(n3591) );
  NOR U5891 ( .A(n1100), .B(n5995), .Z(n6339) );
  XOR U5892 ( .A(n6343), .B(n5766), .Z(out[1114]) );
  XNOR U5893 ( .A(n6344), .B(n5503), .Z(n5766) );
  XOR U5894 ( .A(n6345), .B(n6346), .Z(n5503) );
  NOR U5895 ( .A(n1104), .B(n6000), .Z(n6343) );
  XOR U5896 ( .A(n6347), .B(n5769), .Z(out[1113]) );
  XOR U5897 ( .A(n6348), .B(n5508), .Z(n5769) );
  XOR U5898 ( .A(n6349), .B(n6350), .Z(n5508) );
  NOR U5899 ( .A(n1108), .B(n6005), .Z(n6347) );
  XOR U5900 ( .A(n6351), .B(n5772), .Z(out[1112]) );
  XNOR U5901 ( .A(n6352), .B(n5661), .Z(n5772) );
  XOR U5902 ( .A(n6353), .B(n6354), .Z(n5661) );
  NOR U5903 ( .A(n1112), .B(n6010), .Z(n6351) );
  XOR U5904 ( .A(n6355), .B(n5780), .Z(out[1111]) );
  XNOR U5905 ( .A(n6356), .B(n5707), .Z(n5780) );
  XOR U5906 ( .A(n6357), .B(n6358), .Z(n5707) );
  NOR U5907 ( .A(n1116), .B(n6015), .Z(n6355) );
  XOR U5908 ( .A(n6359), .B(n5783), .Z(out[1110]) );
  XNOR U5909 ( .A(n6360), .B(n5742), .Z(n5783) );
  XOR U5910 ( .A(n6361), .B(n6362), .Z(n5742) );
  NOR U5911 ( .A(n1120), .B(n6020), .Z(n6359) );
  XNOR U5912 ( .A(n6363), .B(n4104), .Z(out[110]) );
  XOR U5913 ( .A(n6364), .B(n2518), .Z(n4104) );
  ANDN U5914 ( .B(n4274), .A(n3307), .Z(n6363) );
  XNOR U5915 ( .A(n6365), .B(n2291), .Z(n3307) );
  XOR U5916 ( .A(n6366), .B(n2358), .Z(n4274) );
  XOR U5917 ( .A(n6367), .B(n5785), .Z(out[1109]) );
  XNOR U5918 ( .A(n6368), .B(n5775), .Z(n5785) );
  XOR U5919 ( .A(n6369), .B(n6370), .Z(n5775) );
  NOR U5920 ( .A(n1124), .B(n6025), .Z(n6367) );
  XOR U5921 ( .A(n6371), .B(n5787), .Z(out[1108]) );
  IV U5922 ( .A(n6031), .Z(n5787) );
  XOR U5923 ( .A(n6372), .B(n2430), .Z(n6031) );
  XNOR U5924 ( .A(n6373), .B(n6374), .Z(n2430) );
  NOR U5925 ( .A(n1128), .B(n6030), .Z(n6371) );
  XOR U5926 ( .A(n6375), .B(n5789), .Z(out[1107]) );
  XNOR U5927 ( .A(n6376), .B(n5833), .Z(n5789) );
  XOR U5928 ( .A(n6377), .B(n6378), .Z(n5833) );
  NOR U5929 ( .A(n1136), .B(n6036), .Z(n6375) );
  XOR U5930 ( .A(n6379), .B(n5791), .Z(out[1106]) );
  XNOR U5931 ( .A(n6380), .B(n5864), .Z(n5791) );
  XOR U5932 ( .A(n6381), .B(n6382), .Z(n5864) );
  NOR U5933 ( .A(n1140), .B(n6041), .Z(n6379) );
  XOR U5934 ( .A(n6383), .B(n5794), .Z(out[1105]) );
  XNOR U5935 ( .A(n6384), .B(n5899), .Z(n5794) );
  XOR U5936 ( .A(n6385), .B(n6386), .Z(n5899) );
  NOR U5937 ( .A(n1144), .B(n6053), .Z(n6383) );
  XOR U5938 ( .A(n6387), .B(n5797), .Z(out[1104]) );
  XNOR U5939 ( .A(n6388), .B(n5932), .Z(n5797) );
  XOR U5940 ( .A(n6389), .B(n6390), .Z(n5932) );
  NOR U5941 ( .A(n1148), .B(n6058), .Z(n6387) );
  XOR U5942 ( .A(n6391), .B(n5800), .Z(out[1103]) );
  XNOR U5943 ( .A(n6392), .B(n5558), .Z(n5800) );
  XOR U5944 ( .A(n6393), .B(n6394), .Z(n5558) );
  NOR U5945 ( .A(n1152), .B(n6063), .Z(n6391) );
  XOR U5946 ( .A(n6395), .B(n5803), .Z(out[1102]) );
  XNOR U5947 ( .A(n6396), .B(n6044), .Z(n5803) );
  XOR U5948 ( .A(n6397), .B(n6398), .Z(n6044) );
  ANDN U5949 ( .B(n6068), .A(n1156), .Z(n6395) );
  XOR U5950 ( .A(n6399), .B(n5811), .Z(out[1101]) );
  XOR U5951 ( .A(n6400), .B(n2483), .Z(n5811) );
  XNOR U5952 ( .A(n6401), .B(n6402), .Z(n2483) );
  ANDN U5953 ( .B(n1160), .A(n6073), .Z(n6399) );
  IV U5954 ( .A(n6403), .Z(n1160) );
  XOR U5955 ( .A(n6404), .B(n5814), .Z(out[1100]) );
  IV U5956 ( .A(n6079), .Z(n5814) );
  XOR U5957 ( .A(n6405), .B(n2490), .Z(n6079) );
  XNOR U5958 ( .A(n6406), .B(n6407), .Z(n2490) );
  NOR U5959 ( .A(n6078), .B(n1164), .Z(n6404) );
  XOR U5960 ( .A(n6408), .B(n2045), .Z(out[10]) );
  XOR U5961 ( .A(n6409), .B(n2629), .Z(n2045) );
  IV U5962 ( .A(n6410), .Z(n2629) );
  NOR U5963 ( .A(n4006), .B(n2044), .Z(n6408) );
  XNOR U5964 ( .A(n2558), .B(n6411), .Z(n2044) );
  XOR U5965 ( .A(n6412), .B(n1757), .Z(n4006) );
  XNOR U5966 ( .A(n6413), .B(n4107), .Z(out[109]) );
  XOR U5967 ( .A(n6414), .B(n2525), .Z(n4107) );
  ANDN U5968 ( .B(n4277), .A(n3349), .Z(n6413) );
  XNOR U5969 ( .A(n6415), .B(n2298), .Z(n3349) );
  XNOR U5970 ( .A(n6416), .B(n2365), .Z(n4277) );
  XOR U5971 ( .A(n6417), .B(n5816), .Z(out[1099]) );
  IV U5972 ( .A(n6085), .Z(n5816) );
  XOR U5973 ( .A(n6418), .B(n2497), .Z(n6085) );
  XNOR U5974 ( .A(n6419), .B(n6420), .Z(n2497) );
  NOR U5975 ( .A(n1168), .B(n6084), .Z(n6417) );
  XOR U5976 ( .A(n6421), .B(n5818), .Z(out[1098]) );
  XOR U5977 ( .A(n6422), .B(n2504), .Z(n5818) );
  XNOR U5978 ( .A(n6423), .B(n6424), .Z(n2504) );
  NOR U5979 ( .A(n1172), .B(n6090), .Z(n6421) );
  XOR U5980 ( .A(n6425), .B(n5820), .Z(out[1097]) );
  IV U5981 ( .A(n6096), .Z(n5820) );
  XOR U5982 ( .A(n6426), .B(n2511), .Z(n6096) );
  XNOR U5983 ( .A(n6427), .B(n6428), .Z(n2511) );
  NOR U5984 ( .A(n1180), .B(n6095), .Z(n6425) );
  XOR U5985 ( .A(n6429), .B(n5822), .Z(out[1096]) );
  XNOR U5986 ( .A(n6430), .B(n2518), .Z(n5822) );
  XNOR U5987 ( .A(n6431), .B(n6432), .Z(n2518) );
  ANDN U5988 ( .B(n1184), .A(n6101), .Z(n6429) );
  XOR U5989 ( .A(n6433), .B(n5824), .Z(out[1095]) );
  XNOR U5990 ( .A(n6434), .B(n2525), .Z(n5824) );
  XNOR U5991 ( .A(n6435), .B(n6436), .Z(n2525) );
  NOR U5992 ( .A(n1188), .B(n6112), .Z(n6433) );
  XOR U5993 ( .A(n6437), .B(n5826), .Z(out[1094]) );
  IV U5994 ( .A(n6118), .Z(n5826) );
  XOR U5995 ( .A(n6438), .B(n2532), .Z(n6118) );
  NOR U5996 ( .A(n1192), .B(n6117), .Z(n6437) );
  XOR U5997 ( .A(n6439), .B(n5828), .Z(out[1093]) );
  IV U5998 ( .A(n6124), .Z(n5828) );
  XOR U5999 ( .A(n6440), .B(n2539), .Z(n6124) );
  NOR U6000 ( .A(n1196), .B(n6123), .Z(n6439) );
  XOR U6001 ( .A(n6441), .B(n5830), .Z(out[1092]) );
  IV U6002 ( .A(n6130), .Z(n5830) );
  XOR U6003 ( .A(n6442), .B(n2550), .Z(n6130) );
  NOR U6004 ( .A(n1200), .B(n6129), .Z(n6441) );
  XOR U6005 ( .A(n6443), .B(n5838), .Z(out[1091]) );
  IV U6006 ( .A(n6136), .Z(n5838) );
  XOR U6007 ( .A(n6444), .B(n2557), .Z(n6136) );
  NOR U6008 ( .A(n1204), .B(n6135), .Z(n6443) );
  XOR U6009 ( .A(n6445), .B(n5840), .Z(out[1090]) );
  IV U6010 ( .A(n6142), .Z(n5840) );
  XOR U6011 ( .A(n6446), .B(n2564), .Z(n6142) );
  NOR U6012 ( .A(n1208), .B(n6141), .Z(n6445) );
  XOR U6013 ( .A(n6447), .B(n4110), .Z(out[108]) );
  IV U6014 ( .A(n4280), .Z(n4110) );
  XOR U6015 ( .A(n6448), .B(n2532), .Z(n4280) );
  XNOR U6016 ( .A(n6449), .B(n6450), .Z(n2532) );
  ANDN U6017 ( .B(n3390), .A(n3391), .Z(n6447) );
  XNOR U6018 ( .A(n6451), .B(n2305), .Z(n3391) );
  XOR U6019 ( .A(n6452), .B(n2374), .Z(n3390) );
  XOR U6020 ( .A(n6453), .B(n5842), .Z(out[1089]) );
  XOR U6021 ( .A(n6454), .B(n2571), .Z(n5842) );
  IV U6022 ( .A(n3707), .Z(n2571) );
  NOR U6023 ( .A(n1212), .B(n6147), .Z(n6453) );
  XOR U6024 ( .A(n6455), .B(n5845), .Z(out[1088]) );
  IV U6025 ( .A(n6153), .Z(n5845) );
  XOR U6026 ( .A(n6456), .B(n2578), .Z(n6153) );
  NOR U6027 ( .A(n1216), .B(n6152), .Z(n6455) );
  XOR U6028 ( .A(n6457), .B(n5847), .Z(out[1087]) );
  XOR U6029 ( .A(n6458), .B(n3284), .Z(n5847) );
  XOR U6030 ( .A(n5922), .B(n6459), .Z(n3284) );
  XOR U6031 ( .A(n6460), .B(n6461), .Z(n5922) );
  XOR U6032 ( .A(n6368), .B(n2422), .Z(n6461) );
  XOR U6033 ( .A(n6462), .B(n6463), .Z(n2422) );
  ANDN U6034 ( .B(n6464), .A(n6465), .Z(n6462) );
  XNOR U6035 ( .A(n6466), .B(n6467), .Z(n6368) );
  ANDN U6036 ( .B(n6468), .A(n6469), .Z(n6466) );
  XOR U6037 ( .A(n3619), .B(n6470), .Z(n6460) );
  XOR U6038 ( .A(n5774), .B(n5534), .Z(n6470) );
  XNOR U6039 ( .A(n6471), .B(n6472), .Z(n5534) );
  ANDN U6040 ( .B(n6473), .A(n6474), .Z(n6471) );
  XNOR U6041 ( .A(n6475), .B(n6476), .Z(n5774) );
  ANDN U6042 ( .B(n6477), .A(n6478), .Z(n6475) );
  XNOR U6043 ( .A(n6479), .B(n6480), .Z(n3619) );
  ANDN U6044 ( .B(n6481), .A(n6482), .Z(n6479) );
  ANDN U6045 ( .B(n5620), .A(n6156), .Z(n6457) );
  XOR U6046 ( .A(n6483), .B(n5849), .Z(out[1086]) );
  XNOR U6047 ( .A(n6484), .B(n5306), .Z(n5849) );
  XOR U6048 ( .A(n5927), .B(n6485), .Z(n5306) );
  XOR U6049 ( .A(n6486), .B(n6487), .Z(n5927) );
  XNOR U6050 ( .A(n6372), .B(n2429), .Z(n6487) );
  XNOR U6051 ( .A(n6488), .B(n6489), .Z(n2429) );
  ANDN U6052 ( .B(n6490), .A(n6491), .Z(n6488) );
  XOR U6053 ( .A(n6492), .B(n6493), .Z(n6372) );
  ANDN U6054 ( .B(n6494), .A(n6495), .Z(n6492) );
  XNOR U6055 ( .A(n3623), .B(n6496), .Z(n6486) );
  XOR U6056 ( .A(n5806), .B(n5537), .Z(n6496) );
  XNOR U6057 ( .A(n6497), .B(n6498), .Z(n5537) );
  ANDN U6058 ( .B(n6499), .A(n6500), .Z(n6497) );
  XNOR U6059 ( .A(n6501), .B(n6502), .Z(n5806) );
  ANDN U6060 ( .B(n6503), .A(n6504), .Z(n6501) );
  XNOR U6061 ( .A(n6505), .B(n6506), .Z(n3623) );
  ANDN U6062 ( .B(n6507), .A(n6508), .Z(n6505) );
  ANDN U6063 ( .B(n5624), .A(n6159), .Z(n6483) );
  XOR U6064 ( .A(n6509), .B(n5851), .Z(out[1085]) );
  XOR U6065 ( .A(n6510), .B(n5311), .Z(n5851) );
  XOR U6066 ( .A(n5938), .B(n6511), .Z(n5311) );
  XOR U6067 ( .A(n6512), .B(n6513), .Z(n5938) );
  XOR U6068 ( .A(n6376), .B(n2436), .Z(n6513) );
  XOR U6069 ( .A(n6514), .B(n6515), .Z(n2436) );
  ANDN U6070 ( .B(n6516), .A(n6517), .Z(n6514) );
  XNOR U6071 ( .A(n6518), .B(n6519), .Z(n6376) );
  ANDN U6072 ( .B(n6520), .A(n6521), .Z(n6518) );
  XOR U6073 ( .A(n3627), .B(n6522), .Z(n6512) );
  XOR U6074 ( .A(n5832), .B(n5542), .Z(n6522) );
  XNOR U6075 ( .A(n6523), .B(n6524), .Z(n5542) );
  ANDN U6076 ( .B(n6525), .A(n6526), .Z(n6523) );
  XNOR U6077 ( .A(n6527), .B(n6528), .Z(n5832) );
  ANDN U6078 ( .B(n6529), .A(n6530), .Z(n6527) );
  XNOR U6079 ( .A(n6531), .B(n6532), .Z(n3627) );
  ANDN U6080 ( .B(n6533), .A(n6534), .Z(n6531) );
  ANDN U6081 ( .B(n5628), .A(n6169), .Z(n6509) );
  XOR U6082 ( .A(n6535), .B(n5854), .Z(out[1084]) );
  XOR U6083 ( .A(n6536), .B(n2575), .Z(n5854) );
  XNOR U6084 ( .A(n5943), .B(n6537), .Z(n2575) );
  XOR U6085 ( .A(n6538), .B(n6539), .Z(n5943) );
  XOR U6086 ( .A(n6380), .B(n2443), .Z(n6539) );
  XOR U6087 ( .A(n6540), .B(n6541), .Z(n2443) );
  ANDN U6088 ( .B(n6542), .A(n6543), .Z(n6540) );
  XNOR U6089 ( .A(n6544), .B(n6545), .Z(n6380) );
  ANDN U6090 ( .B(n6546), .A(n6547), .Z(n6544) );
  XOR U6091 ( .A(n3631), .B(n6548), .Z(n6538) );
  XOR U6092 ( .A(n5863), .B(n5545), .Z(n6548) );
  XOR U6093 ( .A(n6549), .B(n6550), .Z(n5545) );
  XOR U6094 ( .A(n6551), .B(n6552), .Z(n6550) );
  NAND U6095 ( .A(n6553), .B(n6554), .Z(n6552) );
  AND U6096 ( .A(n4564), .B(n6555), .Z(n6554) );
  ANDN U6097 ( .B(n4609), .A(rc_i[9]), .Z(n6555) );
  AND U6098 ( .A(n6556), .B(n6557), .Z(n6553) );
  AND U6099 ( .A(n4343), .B(n4490), .Z(n6557) );
  ANDN U6100 ( .B(n4566), .A(n6558), .Z(n6556) );
  ANDN U6101 ( .B(n6559), .A(n6560), .Z(n6551) );
  XNOR U6102 ( .A(n6561), .B(n6562), .Z(n5863) );
  ANDN U6103 ( .B(n6563), .A(n6564), .Z(n6561) );
  XNOR U6104 ( .A(n6565), .B(n6566), .Z(n3631) );
  ANDN U6105 ( .B(n6567), .A(n6568), .Z(n6565) );
  NOR U6106 ( .A(n5632), .B(n6174), .Z(n6535) );
  XOR U6107 ( .A(n6569), .B(n5857), .Z(out[1083]) );
  XOR U6108 ( .A(n6570), .B(n5325), .Z(n5857) );
  XOR U6109 ( .A(n5948), .B(n6571), .Z(n5325) );
  XOR U6110 ( .A(n6572), .B(n6573), .Z(n5948) );
  XOR U6111 ( .A(n6384), .B(n2450), .Z(n6573) );
  XOR U6112 ( .A(n6574), .B(n6575), .Z(n2450) );
  ANDN U6113 ( .B(n6576), .A(n6577), .Z(n6574) );
  XNOR U6114 ( .A(n6578), .B(n6579), .Z(n6384) );
  ANDN U6115 ( .B(n6580), .A(n6581), .Z(n6578) );
  XOR U6116 ( .A(n3635), .B(n6582), .Z(n6572) );
  XOR U6117 ( .A(n5898), .B(n5550), .Z(n6582) );
  XNOR U6118 ( .A(n6583), .B(n6584), .Z(n5550) );
  AND U6119 ( .A(n6585), .B(n6586), .Z(n6583) );
  XNOR U6120 ( .A(n6587), .B(n6588), .Z(n5898) );
  ANDN U6121 ( .B(n6589), .A(n6590), .Z(n6587) );
  XOR U6122 ( .A(n6591), .B(n6592), .Z(n3635) );
  ANDN U6123 ( .B(n6593), .A(n6594), .Z(n6591) );
  NOR U6124 ( .A(n6179), .B(n5636), .Z(n6569) );
  XOR U6125 ( .A(n6595), .B(n5860), .Z(out[1082]) );
  XOR U6126 ( .A(n6596), .B(n5332), .Z(n5860) );
  XOR U6127 ( .A(n5953), .B(n6597), .Z(n5332) );
  XOR U6128 ( .A(n6598), .B(n6599), .Z(n5953) );
  XOR U6129 ( .A(n6388), .B(n2457), .Z(n6599) );
  XOR U6130 ( .A(n6600), .B(n6601), .Z(n2457) );
  ANDN U6131 ( .B(n6602), .A(n6603), .Z(n6600) );
  XNOR U6132 ( .A(n6604), .B(n6605), .Z(n6388) );
  ANDN U6133 ( .B(n6606), .A(n6607), .Z(n6604) );
  XOR U6134 ( .A(n3644), .B(n6608), .Z(n6598) );
  XOR U6135 ( .A(n5931), .B(n5554), .Z(n6608) );
  XNOR U6136 ( .A(n6609), .B(n6610), .Z(n5554) );
  ANDN U6137 ( .B(n6611), .A(n6612), .Z(n6609) );
  XNOR U6138 ( .A(n6613), .B(n6614), .Z(n5931) );
  ANDN U6139 ( .B(n6615), .A(n6616), .Z(n6613) );
  XOR U6140 ( .A(n6617), .B(n6618), .Z(n3644) );
  ANDN U6141 ( .B(n6619), .A(n6620), .Z(n6617) );
  ANDN U6142 ( .B(n5640), .A(n6184), .Z(n6595) );
  XOR U6143 ( .A(n6621), .B(n5869), .Z(out[1081]) );
  XOR U6144 ( .A(n6622), .B(n5338), .Z(n5869) );
  XOR U6145 ( .A(n6623), .B(n5959), .Z(n5338) );
  XNOR U6146 ( .A(n6624), .B(n6625), .Z(n5959) );
  XNOR U6147 ( .A(n5557), .B(n3648), .Z(n6625) );
  XOR U6148 ( .A(n6626), .B(n6627), .Z(n3648) );
  ANDN U6149 ( .B(n6628), .A(n6629), .Z(n6626) );
  XNOR U6150 ( .A(n6630), .B(n6631), .Z(n5557) );
  NOR U6151 ( .A(n6632), .B(n6633), .Z(n6630) );
  XOR U6152 ( .A(n6392), .B(n6634), .Z(n6624) );
  XOR U6153 ( .A(n2464), .B(n5987), .Z(n6634) );
  XNOR U6154 ( .A(n6635), .B(n6636), .Z(n5987) );
  ANDN U6155 ( .B(n6637), .A(n6638), .Z(n6635) );
  XNOR U6156 ( .A(n6639), .B(n6640), .Z(n2464) );
  ANDN U6157 ( .B(n6641), .A(n6642), .Z(n6639) );
  XNOR U6158 ( .A(n6643), .B(n6644), .Z(n6392) );
  AND U6159 ( .A(n6645), .B(n6646), .Z(n6643) );
  ANDN U6160 ( .B(n5644), .A(n6189), .Z(n6621) );
  XOR U6161 ( .A(n6647), .B(n5871), .Z(out[1080]) );
  XNOR U6162 ( .A(n6648), .B(n5343), .Z(n5871) );
  XOR U6163 ( .A(n6649), .B(n5964), .Z(n5343) );
  XNOR U6164 ( .A(n6650), .B(n6651), .Z(n5964) );
  XNOR U6165 ( .A(n5563), .B(n3652), .Z(n6651) );
  XOR U6166 ( .A(n6652), .B(n6653), .Z(n3652) );
  XNOR U6167 ( .A(n6656), .B(n6657), .Z(n5563) );
  AND U6168 ( .A(n6658), .B(n6659), .Z(n6656) );
  XOR U6169 ( .A(n6396), .B(n6660), .Z(n6650) );
  XOR U6170 ( .A(n2475), .B(n6043), .Z(n6660) );
  XNOR U6171 ( .A(n6661), .B(n6662), .Z(n6043) );
  AND U6172 ( .A(n6663), .B(n6664), .Z(n6661) );
  XNOR U6173 ( .A(n6665), .B(n6666), .Z(n2475) );
  XNOR U6174 ( .A(n6669), .B(n6670), .Z(n6396) );
  AND U6175 ( .A(n6671), .B(n6672), .Z(n6669) );
  ANDN U6176 ( .B(n5648), .A(n6194), .Z(n6647) );
  XOR U6177 ( .A(n6673), .B(n4113), .Z(out[107]) );
  IV U6178 ( .A(n4283), .Z(n4113) );
  XOR U6179 ( .A(n6674), .B(n2539), .Z(n4283) );
  XNOR U6180 ( .A(n6675), .B(n6676), .Z(n2539) );
  ANDN U6181 ( .B(n3418), .A(n3420), .Z(n6673) );
  XNOR U6182 ( .A(n6677), .B(n2312), .Z(n3420) );
  XOR U6183 ( .A(n6678), .B(n2379), .Z(n3418) );
  XOR U6184 ( .A(n6679), .B(n5874), .Z(out[1079]) );
  XNOR U6185 ( .A(n6680), .B(n5520), .Z(n5874) );
  XOR U6186 ( .A(n6681), .B(n5969), .Z(n5520) );
  XNOR U6187 ( .A(n6682), .B(n6683), .Z(n5969) );
  XOR U6188 ( .A(n5566), .B(n3656), .Z(n6683) );
  XOR U6189 ( .A(n6684), .B(n6685), .Z(n3656) );
  ANDN U6190 ( .B(n6686), .A(n6687), .Z(n6684) );
  XNOR U6191 ( .A(n6688), .B(n6689), .Z(n5566) );
  ANDN U6192 ( .B(n6690), .A(n6691), .Z(n6688) );
  XOR U6193 ( .A(n6400), .B(n6692), .Z(n6682) );
  XOR U6194 ( .A(n2482), .B(n6103), .Z(n6692) );
  XNOR U6195 ( .A(n6693), .B(n6694), .Z(n6103) );
  ANDN U6196 ( .B(n6695), .A(n6696), .Z(n6693) );
  XNOR U6197 ( .A(n6697), .B(n6698), .Z(n2482) );
  ANDN U6198 ( .B(n6699), .A(n6700), .Z(n6697) );
  XNOR U6199 ( .A(n6701), .B(n6702), .Z(n6400) );
  ANDN U6200 ( .B(n6703), .A(n6704), .Z(n6701) );
  ANDN U6201 ( .B(n5652), .A(n6199), .Z(n6679) );
  XOR U6202 ( .A(n6705), .B(n5877), .Z(out[1078]) );
  XNOR U6203 ( .A(n6706), .B(n5894), .Z(n5877) );
  XOR U6204 ( .A(n6707), .B(n5974), .Z(n5894) );
  XNOR U6205 ( .A(n6708), .B(n6709), .Z(n5974) );
  XOR U6206 ( .A(n5573), .B(n3660), .Z(n6709) );
  XNOR U6207 ( .A(n6710), .B(n6711), .Z(n3660) );
  ANDN U6208 ( .B(n6712), .A(n6713), .Z(n6710) );
  XNOR U6209 ( .A(n6714), .B(n6715), .Z(n5573) );
  ANDN U6210 ( .B(n6716), .A(n6717), .Z(n6714) );
  XNOR U6211 ( .A(n6405), .B(n6718), .Z(n6708) );
  XOR U6212 ( .A(n2489), .B(n6161), .Z(n6718) );
  XOR U6213 ( .A(n6719), .B(n6720), .Z(n6161) );
  ANDN U6214 ( .B(n6721), .A(n6722), .Z(n6719) );
  XOR U6215 ( .A(n6723), .B(n6724), .Z(n2489) );
  ANDN U6216 ( .B(n6725), .A(n6726), .Z(n6723) );
  XOR U6217 ( .A(n6727), .B(n6728), .Z(n6405) );
  ANDN U6218 ( .B(n6729), .A(n6730), .Z(n6727) );
  ANDN U6219 ( .B(n5656), .A(n6204), .Z(n6705) );
  XOR U6220 ( .A(n6731), .B(n5879), .Z(out[1077]) );
  XNOR U6221 ( .A(n6732), .B(n6410), .Z(n5879) );
  XOR U6222 ( .A(n6733), .B(n5979), .Z(n6410) );
  XNOR U6223 ( .A(n6734), .B(n6735), .Z(n5979) );
  XOR U6224 ( .A(n5577), .B(n3664), .Z(n6735) );
  XOR U6225 ( .A(n6736), .B(n6737), .Z(n3664) );
  ANDN U6226 ( .B(n6738), .A(n6739), .Z(n6736) );
  XNOR U6227 ( .A(n6740), .B(n6741), .Z(n5577) );
  ANDN U6228 ( .B(n6742), .A(n6743), .Z(n6740) );
  XNOR U6229 ( .A(n6418), .B(n6744), .Z(n6734) );
  XOR U6230 ( .A(n2496), .B(n6216), .Z(n6744) );
  XOR U6231 ( .A(n6745), .B(n6746), .Z(n6216) );
  ANDN U6232 ( .B(n6747), .A(n6748), .Z(n6745) );
  XNOR U6233 ( .A(n6749), .B(n6750), .Z(n2496) );
  ANDN U6234 ( .B(n6751), .A(n6752), .Z(n6749) );
  XOR U6235 ( .A(n6753), .B(n6754), .Z(n6418) );
  ANDN U6236 ( .B(n6755), .A(n6756), .Z(n6753) );
  ANDN U6237 ( .B(n5666), .A(n6209), .Z(n6731) );
  XOR U6238 ( .A(n6757), .B(n5881), .Z(out[1076]) );
  XNOR U6239 ( .A(n5360), .B(n6758), .Z(n5881) );
  XOR U6240 ( .A(n5983), .B(n6759), .Z(n5360) );
  XOR U6241 ( .A(n6760), .B(n6761), .Z(n5983) );
  XNOR U6242 ( .A(n6422), .B(n2503), .Z(n6761) );
  XOR U6243 ( .A(n6762), .B(n6763), .Z(n2503) );
  NOR U6244 ( .A(n6764), .B(n6765), .Z(n6762) );
  XOR U6245 ( .A(n6766), .B(n6767), .Z(n6422) );
  ANDN U6246 ( .B(n6768), .A(n6769), .Z(n6766) );
  XOR U6247 ( .A(n3668), .B(n6770), .Z(n6760) );
  XOR U6248 ( .A(n6273), .B(n5582), .Z(n6770) );
  XNOR U6249 ( .A(n6771), .B(n6772), .Z(n5582) );
  XOR U6250 ( .A(n6773), .B(n6774), .Z(n6772) );
  NAND U6251 ( .A(n6775), .B(n6776), .Z(n6774) );
  ANDN U6252 ( .B(n6777), .A(rc_i[4]), .Z(n6776) );
  AND U6253 ( .A(n4608), .B(n4657), .Z(n6777) );
  ANDN U6254 ( .B(n6778), .A(n6779), .Z(n6775) );
  AND U6255 ( .A(n4566), .B(n4340), .Z(n6778) );
  ANDN U6256 ( .B(n6780), .A(n6781), .Z(n6773) );
  XOR U6257 ( .A(n6782), .B(n6783), .Z(n6273) );
  ANDN U6258 ( .B(n6784), .A(n6785), .Z(n6782) );
  XOR U6259 ( .A(n6786), .B(n6787), .Z(n3668) );
  ANDN U6260 ( .B(n6788), .A(n6789), .Z(n6786) );
  ANDN U6261 ( .B(n5670), .A(n6214), .Z(n6757) );
  XOR U6262 ( .A(n6790), .B(n5884), .Z(out[1075]) );
  XNOR U6263 ( .A(n6791), .B(n5365), .Z(n5884) );
  XOR U6264 ( .A(n6792), .B(n5994), .Z(n5365) );
  XNOR U6265 ( .A(n6793), .B(n6794), .Z(n5994) );
  XOR U6266 ( .A(n5586), .B(n3672), .Z(n6794) );
  XOR U6267 ( .A(n6795), .B(n6796), .Z(n3672) );
  ANDN U6268 ( .B(n6797), .A(n6798), .Z(n6795) );
  XNOR U6269 ( .A(n6799), .B(n6800), .Z(n5586) );
  ANDN U6270 ( .B(n6801), .A(n6802), .Z(n6799) );
  XNOR U6271 ( .A(n6426), .B(n6803), .Z(n6793) );
  XOR U6272 ( .A(n2510), .B(n6320), .Z(n6803) );
  XOR U6273 ( .A(n6804), .B(n6805), .Z(n6320) );
  ANDN U6274 ( .B(n6806), .A(n6807), .Z(n6804) );
  XOR U6275 ( .A(n6808), .B(n6809), .Z(n2510) );
  NOR U6276 ( .A(n6810), .B(n6811), .Z(n6808) );
  XOR U6277 ( .A(n6812), .B(n6813), .Z(n6426) );
  ANDN U6278 ( .B(n6814), .A(n6815), .Z(n6812) );
  ANDN U6279 ( .B(n5674), .A(n6224), .Z(n6790) );
  XOR U6280 ( .A(n6816), .B(n5886), .Z(out[1074]) );
  XNOR U6281 ( .A(n6817), .B(n5374), .Z(n5886) );
  XOR U6282 ( .A(n6818), .B(n5999), .Z(n5374) );
  XNOR U6283 ( .A(n6819), .B(n6820), .Z(n5999) );
  XOR U6284 ( .A(n5591), .B(n3676), .Z(n6820) );
  XOR U6285 ( .A(n6821), .B(n6822), .Z(n3676) );
  ANDN U6286 ( .B(n6823), .A(n6824), .Z(n6821) );
  XNOR U6287 ( .A(n6825), .B(n6826), .Z(n5591) );
  ANDN U6288 ( .B(n6827), .A(n6828), .Z(n6825) );
  XNOR U6289 ( .A(n6430), .B(n6829), .Z(n6819) );
  XOR U6290 ( .A(n2517), .B(n6364), .Z(n6829) );
  XOR U6291 ( .A(n6830), .B(n6831), .Z(n6364) );
  ANDN U6292 ( .B(n6832), .A(n6833), .Z(n6830) );
  XOR U6293 ( .A(n6834), .B(n6835), .Z(n2517) );
  ANDN U6294 ( .B(n6836), .A(n6837), .Z(n6834) );
  XOR U6295 ( .A(n6838), .B(n6839), .Z(n6430) );
  ANDN U6296 ( .B(n6840), .A(n6841), .Z(n6838) );
  ANDN U6297 ( .B(n5678), .A(n6229), .Z(n6816) );
  XOR U6298 ( .A(n6842), .B(n5888), .Z(out[1073]) );
  XNOR U6299 ( .A(n6843), .B(n5379), .Z(n5888) );
  XOR U6300 ( .A(n6844), .B(n6004), .Z(n5379) );
  XNOR U6301 ( .A(n6845), .B(n6846), .Z(n6004) );
  XOR U6302 ( .A(n5596), .B(n3680), .Z(n6846) );
  XOR U6303 ( .A(n6847), .B(n6848), .Z(n3680) );
  AND U6304 ( .A(n6849), .B(n6850), .Z(n6847) );
  XNOR U6305 ( .A(n6851), .B(n6852), .Z(n5596) );
  ANDN U6306 ( .B(n6853), .A(n6854), .Z(n6851) );
  XNOR U6307 ( .A(n6434), .B(n6855), .Z(n6845) );
  XOR U6308 ( .A(n2524), .B(n6414), .Z(n6855) );
  XOR U6309 ( .A(n6856), .B(n6857), .Z(n6414) );
  ANDN U6310 ( .B(n6858), .A(n6859), .Z(n6856) );
  XOR U6311 ( .A(n6860), .B(n6861), .Z(n2524) );
  NOR U6312 ( .A(n6862), .B(n6863), .Z(n6860) );
  XOR U6313 ( .A(n6864), .B(n6865), .Z(n6434) );
  ANDN U6314 ( .B(n6866), .A(n6867), .Z(n6864) );
  ANDN U6315 ( .B(n5682), .A(n6234), .Z(n6842) );
  XOR U6316 ( .A(n6868), .B(n5890), .Z(out[1072]) );
  XOR U6317 ( .A(n6869), .B(n2664), .Z(n5890) );
  XOR U6318 ( .A(n6870), .B(n6009), .Z(n2664) );
  XNOR U6319 ( .A(n6871), .B(n6872), .Z(n6009) );
  XOR U6320 ( .A(n5602), .B(n3686), .Z(n6872) );
  XOR U6321 ( .A(n6873), .B(n6874), .Z(n3686) );
  AND U6322 ( .A(n6875), .B(n6876), .Z(n6873) );
  XOR U6323 ( .A(n6877), .B(n6878), .Z(n5602) );
  XOR U6324 ( .A(n6879), .B(n6880), .Z(n6878) );
  NAND U6325 ( .A(n6881), .B(n6882), .Z(n6880) );
  AND U6326 ( .A(n6883), .B(n4649), .Z(n6882) );
  NOR U6327 ( .A(rc_i[7]), .B(rc_i[9]), .Z(n4649) );
  AND U6328 ( .A(n6884), .B(n4343), .Z(n6881) );
  NOR U6329 ( .A(rc_i[2]), .B(rc_i[4]), .Z(n6884) );
  ANDN U6330 ( .B(n6885), .A(n6886), .Z(n6879) );
  XNOR U6331 ( .A(n6438), .B(n6887), .Z(n6871) );
  XOR U6332 ( .A(n2531), .B(n6448), .Z(n6887) );
  XNOR U6333 ( .A(n6888), .B(n6889), .Z(n6448) );
  AND U6334 ( .A(n6890), .B(n6891), .Z(n6888) );
  XOR U6335 ( .A(n6892), .B(n6893), .Z(n2531) );
  NOR U6336 ( .A(n6894), .B(n6895), .Z(n6892) );
  XOR U6337 ( .A(n6896), .B(n6897), .Z(n6438) );
  AND U6338 ( .A(n6898), .B(n6899), .Z(n6896) );
  ANDN U6339 ( .B(n5686), .A(n6239), .Z(n6868) );
  XOR U6340 ( .A(n6900), .B(n5904), .Z(out[1071]) );
  XNOR U6341 ( .A(n6901), .B(n3344), .Z(n5904) );
  XOR U6342 ( .A(n6902), .B(n6014), .Z(n3344) );
  XNOR U6343 ( .A(n6903), .B(n6904), .Z(n6014) );
  XOR U6344 ( .A(n5605), .B(n3691), .Z(n6904) );
  XOR U6345 ( .A(n6905), .B(n6906), .Z(n3691) );
  AND U6346 ( .A(n6907), .B(n6908), .Z(n6905) );
  XNOR U6347 ( .A(n6909), .B(n6910), .Z(n5605) );
  ANDN U6348 ( .B(n6911), .A(n6912), .Z(n6909) );
  XNOR U6349 ( .A(n6440), .B(n6913), .Z(n6903) );
  XOR U6350 ( .A(n2538), .B(n6674), .Z(n6913) );
  XOR U6351 ( .A(n6914), .B(n6915), .Z(n6674) );
  AND U6352 ( .A(n6916), .B(n6917), .Z(n6914) );
  XOR U6353 ( .A(n6918), .B(n6919), .Z(n2538) );
  NOR U6354 ( .A(n6920), .B(n6921), .Z(n6918) );
  XOR U6355 ( .A(n6922), .B(n6923), .Z(n6440) );
  NOR U6356 ( .A(n6924), .B(n6925), .Z(n6922) );
  ANDN U6357 ( .B(n5690), .A(n6244), .Z(n6900) );
  XOR U6358 ( .A(n6926), .B(n5907), .Z(out[1070]) );
  XOR U6359 ( .A(n6927), .B(n2678), .Z(n5907) );
  XOR U6360 ( .A(n6928), .B(n6019), .Z(n2678) );
  XNOR U6361 ( .A(n6929), .B(n6930), .Z(n6019) );
  XOR U6362 ( .A(n5610), .B(n3694), .Z(n6930) );
  XOR U6363 ( .A(n6931), .B(n6932), .Z(n3694) );
  AND U6364 ( .A(n6933), .B(n6934), .Z(n6931) );
  XOR U6365 ( .A(n6935), .B(n6936), .Z(n5610) );
  XOR U6366 ( .A(n6937), .B(n6938), .Z(n6936) );
  NAND U6367 ( .A(n6939), .B(n6940), .Z(n6938) );
  AND U6368 ( .A(n4339), .B(n4608), .Z(n6940) );
  NOR U6369 ( .A(rc_i[8]), .B(rc_i[9]), .Z(n4339) );
  NOR U6370 ( .A(rc_i[4]), .B(n6779), .Z(n6939) );
  NAND U6371 ( .A(n4490), .B(n4343), .Z(n6779) );
  ANDN U6372 ( .B(n6941), .A(n6942), .Z(n6937) );
  XNOR U6373 ( .A(n6442), .B(n6943), .Z(n6929) );
  XOR U6374 ( .A(n2549), .B(n6944), .Z(n6943) );
  XOR U6375 ( .A(n6945), .B(n6946), .Z(n2549) );
  NOR U6376 ( .A(n6947), .B(n6948), .Z(n6945) );
  XOR U6377 ( .A(n6949), .B(n6950), .Z(n6442) );
  ANDN U6378 ( .B(n6951), .A(n6952), .Z(n6949) );
  NOR U6379 ( .A(n5694), .B(n6249), .Z(n6926) );
  XOR U6380 ( .A(n6953), .B(n4116), .Z(out[106]) );
  IV U6381 ( .A(n4286), .Z(n4116) );
  XOR U6382 ( .A(n6944), .B(n2550), .Z(n4286) );
  XNOR U6383 ( .A(n6954), .B(n6955), .Z(n2550) );
  XOR U6384 ( .A(n6956), .B(n6957), .Z(n6944) );
  ANDN U6385 ( .B(n6958), .A(n6959), .Z(n6956) );
  ANDN U6386 ( .B(n3442), .A(n3444), .Z(n6953) );
  XNOR U6387 ( .A(n6960), .B(n2319), .Z(n3444) );
  XNOR U6388 ( .A(n6961), .B(n2386), .Z(n3442) );
  XOR U6389 ( .A(n6962), .B(n5909), .Z(out[1069]) );
  XOR U6390 ( .A(n6963), .B(n2685), .Z(n5909) );
  XOR U6391 ( .A(n6964), .B(n6024), .Z(n2685) );
  XNOR U6392 ( .A(n6965), .B(n6966), .Z(n6024) );
  XOR U6393 ( .A(n5614), .B(n3698), .Z(n6966) );
  XOR U6394 ( .A(n6967), .B(n6968), .Z(n3698) );
  AND U6395 ( .A(n6969), .B(n6970), .Z(n6967) );
  XOR U6396 ( .A(n6971), .B(n6972), .Z(n5614) );
  XOR U6397 ( .A(n6973), .B(n6974), .Z(n6972) );
  NAND U6398 ( .A(n6975), .B(n6976), .Z(n6974) );
  AND U6399 ( .A(n6977), .B(n4564), .Z(n6976) );
  AND U6400 ( .A(n4340), .B(n4657), .Z(n4564) );
  AND U6401 ( .A(n4491), .B(n4490), .Z(n6977) );
  IV U6402 ( .A(rc_i[2]), .Z(n4490) );
  ANDN U6403 ( .B(n4605), .A(n6558), .Z(n6975) );
  NAND U6404 ( .A(n4608), .B(n4635), .Z(n6558) );
  AND U6405 ( .A(n4565), .B(n4566), .Z(n4605) );
  IV U6406 ( .A(rc_i[0]), .Z(n4565) );
  AND U6407 ( .A(n6978), .B(n6979), .Z(n6973) );
  XNOR U6408 ( .A(n6444), .B(n6980), .Z(n6965) );
  XOR U6409 ( .A(n2556), .B(n6981), .Z(n6980) );
  XOR U6410 ( .A(n6982), .B(n6983), .Z(n2556) );
  NOR U6411 ( .A(n6984), .B(n6985), .Z(n6982) );
  XOR U6412 ( .A(n6986), .B(n6987), .Z(n6444) );
  ANDN U6413 ( .B(n6988), .A(n6989), .Z(n6986) );
  ANDN U6414 ( .B(n5698), .A(n6254), .Z(n6962) );
  XOR U6415 ( .A(n6990), .B(n5911), .Z(out[1068]) );
  XOR U6416 ( .A(n6991), .B(n2692), .Z(n5911) );
  XOR U6417 ( .A(n6992), .B(n6029), .Z(n2692) );
  XNOR U6418 ( .A(n6993), .B(n6994), .Z(n6029) );
  XOR U6419 ( .A(n5297), .B(n3702), .Z(n6994) );
  XOR U6420 ( .A(n6995), .B(n6996), .Z(n3702) );
  ANDN U6421 ( .B(n6997), .A(n6998), .Z(n6995) );
  XOR U6422 ( .A(n6999), .B(n7000), .Z(n5297) );
  XOR U6423 ( .A(n7001), .B(n7002), .Z(n7000) );
  NAND U6424 ( .A(n7003), .B(n7004), .Z(n7002) );
  AND U6425 ( .A(n7005), .B(n4340), .Z(n7004) );
  AND U6426 ( .A(n4657), .B(n4609), .Z(n7005) );
  IV U6427 ( .A(rc_i[8]), .Z(n4609) );
  IV U6428 ( .A(rc_i[7]), .Z(n4657) );
  AND U6429 ( .A(n4566), .B(n4343), .Z(n7003) );
  IV U6430 ( .A(rc_i[1]), .Z(n4343) );
  AND U6431 ( .A(n7006), .B(n7007), .Z(n7001) );
  XNOR U6432 ( .A(n6446), .B(n7008), .Z(n6993) );
  XOR U6433 ( .A(n2563), .B(n7009), .Z(n7008) );
  XNOR U6434 ( .A(n7010), .B(n7011), .Z(n2563) );
  NOR U6435 ( .A(n7012), .B(n7013), .Z(n7010) );
  XNOR U6436 ( .A(n7014), .B(n7015), .Z(n6446) );
  ANDN U6437 ( .B(n7016), .A(n7017), .Z(n7014) );
  ANDN U6438 ( .B(n5702), .A(n6259), .Z(n6990) );
  XOR U6439 ( .A(n7018), .B(n5913), .Z(out[1067]) );
  IV U6440 ( .A(n6265), .Z(n5913) );
  XOR U6441 ( .A(n2222), .B(n7019), .Z(n6265) );
  ANDN U6442 ( .B(n5712), .A(n6264), .Z(n7018) );
  XOR U6443 ( .A(n7020), .B(n5915), .Z(out[1066]) );
  IV U6444 ( .A(n6271), .Z(n5915) );
  XOR U6445 ( .A(n2229), .B(n7021), .Z(n6271) );
  XOR U6446 ( .A(n7022), .B(n6040), .Z(n2229) );
  XNOR U6447 ( .A(n7023), .B(n7024), .Z(n6040) );
  XNOR U6448 ( .A(n5304), .B(n3711), .Z(n7024) );
  XOR U6449 ( .A(n7025), .B(n7026), .Z(n3711) );
  AND U6450 ( .A(n7027), .B(n7028), .Z(n7025) );
  XNOR U6451 ( .A(n7029), .B(n7030), .Z(n5304) );
  ANDN U6452 ( .B(n7031), .A(n7032), .Z(n7029) );
  XNOR U6453 ( .A(n6456), .B(n7033), .Z(n7023) );
  XOR U6454 ( .A(n2577), .B(n7034), .Z(n7033) );
  XNOR U6455 ( .A(n7035), .B(n7036), .Z(n2577) );
  ANDN U6456 ( .B(n7037), .A(n7038), .Z(n7035) );
  XNOR U6457 ( .A(n7039), .B(n7040), .Z(n6456) );
  ANDN U6458 ( .B(n7041), .A(n7042), .Z(n7039) );
  ANDN U6459 ( .B(n5716), .A(n6270), .Z(n7020) );
  XOR U6460 ( .A(n7043), .B(n5917), .Z(out[1065]) );
  XOR U6461 ( .A(n5663), .B(n7044), .Z(n5917) );
  XNOR U6462 ( .A(n7045), .B(n6052), .Z(n5663) );
  XNOR U6463 ( .A(n7046), .B(n7047), .Z(n6052) );
  XNOR U6464 ( .A(n5309), .B(n3715), .Z(n7047) );
  XOR U6465 ( .A(n7048), .B(n7049), .Z(n3715) );
  AND U6466 ( .A(n7050), .B(n7051), .Z(n7048) );
  XNOR U6467 ( .A(n7052), .B(n7053), .Z(n5309) );
  ANDN U6468 ( .B(n7054), .A(n7055), .Z(n7052) );
  XNOR U6469 ( .A(n6155), .B(n7056), .Z(n7046) );
  XOR U6470 ( .A(n2584), .B(n7057), .Z(n7056) );
  XNOR U6471 ( .A(n7058), .B(n7059), .Z(n2584) );
  AND U6472 ( .A(n7060), .B(n7061), .Z(n7058) );
  XNOR U6473 ( .A(n7062), .B(n7063), .Z(n6155) );
  ANDN U6474 ( .B(n7064), .A(n7065), .Z(n7062) );
  ANDN U6475 ( .B(n5720), .A(n6281), .Z(n7043) );
  XOR U6476 ( .A(n7066), .B(n5919), .Z(out[1064]) );
  XOR U6477 ( .A(n5709), .B(n7067), .Z(n5919) );
  XNOR U6478 ( .A(n7068), .B(n6057), .Z(n5709) );
  XNOR U6479 ( .A(n7069), .B(n7070), .Z(n6057) );
  XNOR U6480 ( .A(n5318), .B(n3719), .Z(n7070) );
  XOR U6481 ( .A(n7071), .B(n7072), .Z(n3719) );
  AND U6482 ( .A(n7073), .B(n7074), .Z(n7071) );
  XNOR U6483 ( .A(n7075), .B(n7076), .Z(n5318) );
  ANDN U6484 ( .B(n7077), .A(n7078), .Z(n7075) );
  XNOR U6485 ( .A(n6158), .B(n7079), .Z(n7069) );
  XOR U6486 ( .A(n2591), .B(n7080), .Z(n7079) );
  XNOR U6487 ( .A(n7081), .B(n7082), .Z(n2591) );
  AND U6488 ( .A(n7083), .B(n7084), .Z(n7081) );
  XNOR U6489 ( .A(n7085), .B(n7086), .Z(n6158) );
  ANDN U6490 ( .B(n7087), .A(n7088), .Z(n7085) );
  ANDN U6491 ( .B(n5724), .A(n6286), .Z(n7066) );
  XNOR U6492 ( .A(n7089), .B(n5924), .Z(out[1063]) );
  XOR U6493 ( .A(n2257), .B(n7090), .Z(n5924) );
  XOR U6494 ( .A(n7091), .B(n6062), .Z(n2257) );
  XNOR U6495 ( .A(n7092), .B(n7093), .Z(n6062) );
  XOR U6496 ( .A(n5322), .B(n3723), .Z(n7093) );
  XOR U6497 ( .A(n7094), .B(n7095), .Z(n3723) );
  AND U6498 ( .A(n7096), .B(n7097), .Z(n7094) );
  XNOR U6499 ( .A(n7098), .B(n7099), .Z(n5322) );
  AND U6500 ( .A(n7100), .B(n7101), .Z(n7098) );
  XNOR U6501 ( .A(n6166), .B(n7102), .Z(n7092) );
  XOR U6502 ( .A(n4312), .B(n2599), .Z(n7102) );
  XOR U6503 ( .A(n7103), .B(n7104), .Z(n2599) );
  AND U6504 ( .A(n7105), .B(n7106), .Z(n7103) );
  XOR U6505 ( .A(n7107), .B(n7108), .Z(n4312) );
  ANDN U6506 ( .B(n7109), .A(n7110), .Z(n7107) );
  XOR U6507 ( .A(n7111), .B(n7112), .Z(n6166) );
  ANDN U6508 ( .B(n7113), .A(n7114), .Z(n7111) );
  ANDN U6509 ( .B(n1048), .A(n1049), .Z(n7089) );
  XNOR U6510 ( .A(n1795), .B(n7115), .Z(n1049) );
  IV U6511 ( .A(n5181), .Z(n1795) );
  XOR U6512 ( .A(n6623), .B(n6401), .Z(n5181) );
  XOR U6513 ( .A(n7116), .B(n7117), .Z(n6401) );
  XNOR U6514 ( .A(n5972), .B(n2151), .Z(n7117) );
  XNOR U6515 ( .A(n7118), .B(n7119), .Z(n2151) );
  ANDN U6516 ( .B(n6694), .A(n6695), .Z(n7118) );
  XNOR U6517 ( .A(n7120), .B(n7121), .Z(n5972) );
  ANDN U6518 ( .B(n6685), .A(n6686), .Z(n7120) );
  XNOR U6519 ( .A(n5497), .B(n7122), .Z(n7116) );
  XOR U6520 ( .A(n4264), .B(n3695), .Z(n7122) );
  XNOR U6521 ( .A(n7123), .B(n7124), .Z(n3695) );
  ANDN U6522 ( .B(n6689), .A(n6690), .Z(n7123) );
  XNOR U6523 ( .A(n7125), .B(n7126), .Z(n4264) );
  ANDN U6524 ( .B(n6702), .A(n6703), .Z(n7125) );
  XNOR U6525 ( .A(n7127), .B(n7128), .Z(n5497) );
  ANDN U6526 ( .B(n6698), .A(n6699), .Z(n7127) );
  XOR U6527 ( .A(n7129), .B(n7130), .Z(n6623) );
  XNOR U6528 ( .A(n3494), .B(n4859), .Z(n7130) );
  XNOR U6529 ( .A(n7131), .B(n6671), .Z(n4859) );
  ANDN U6530 ( .B(n7132), .A(n7133), .Z(n7131) );
  XNOR U6531 ( .A(n7134), .B(n6663), .Z(n3494) );
  ANDN U6532 ( .B(n7135), .A(n7136), .Z(n7134) );
  XNOR U6533 ( .A(n7137), .B(n7138), .Z(n7129) );
  XOR U6534 ( .A(n4009), .B(n2566), .Z(n7138) );
  XNOR U6535 ( .A(n7139), .B(n6654), .Z(n2566) );
  ANDN U6536 ( .B(n7140), .A(n7141), .Z(n7139) );
  XNOR U6537 ( .A(n7142), .B(n6658), .Z(n4009) );
  ANDN U6538 ( .B(n7143), .A(n7144), .Z(n7142) );
  XNOR U6539 ( .A(n2338), .B(n7145), .Z(n1048) );
  XOR U6540 ( .A(n7146), .B(n5929), .Z(out[1062]) );
  XNOR U6541 ( .A(n7147), .B(n5778), .Z(n5929) );
  XOR U6542 ( .A(n7148), .B(n6067), .Z(n5778) );
  XNOR U6543 ( .A(n7149), .B(n7150), .Z(n6067) );
  XOR U6544 ( .A(n5329), .B(n3729), .Z(n7150) );
  XOR U6545 ( .A(n7151), .B(n7152), .Z(n3729) );
  ANDN U6546 ( .B(n7153), .A(n7154), .Z(n7151) );
  XNOR U6547 ( .A(n7155), .B(n7156), .Z(n5329) );
  ANDN U6548 ( .B(n7157), .A(n7158), .Z(n7155) );
  XNOR U6549 ( .A(n6171), .B(n7159), .Z(n7149) );
  XOR U6550 ( .A(n4316), .B(n2606), .Z(n7159) );
  XOR U6551 ( .A(n7160), .B(n7161), .Z(n2606) );
  ANDN U6552 ( .B(n7162), .A(n7163), .Z(n7160) );
  XOR U6553 ( .A(n7164), .B(n7165), .Z(n4316) );
  ANDN U6554 ( .B(n7166), .A(n7167), .Z(n7164) );
  XNOR U6555 ( .A(n7168), .B(n7169), .Z(n6171) );
  ANDN U6556 ( .B(n7170), .A(n7171), .Z(n7168) );
  ANDN U6557 ( .B(n1052), .A(n1053), .Z(n7146) );
  XNOR U6558 ( .A(n7172), .B(n1800), .Z(n1053) );
  XOR U6559 ( .A(n6649), .B(n6406), .Z(n1800) );
  XOR U6560 ( .A(n7173), .B(n7174), .Z(n6406) );
  XOR U6561 ( .A(n5501), .B(n4267), .Z(n7174) );
  XOR U6562 ( .A(n7175), .B(n7176), .Z(n4267) );
  ANDN U6563 ( .B(n6728), .A(n6729), .Z(n7175) );
  XNOR U6564 ( .A(n7177), .B(n7178), .Z(n5501) );
  ANDN U6565 ( .B(n6724), .A(n6725), .Z(n7177) );
  XOR U6566 ( .A(n3699), .B(n7179), .Z(n7173) );
  XOR U6567 ( .A(n5977), .B(n2154), .Z(n7179) );
  XNOR U6568 ( .A(n7180), .B(n7181), .Z(n2154) );
  ANDN U6569 ( .B(n6720), .A(n6721), .Z(n7180) );
  XNOR U6570 ( .A(n7182), .B(n7183), .Z(n5977) );
  NOR U6571 ( .A(n6711), .B(n6712), .Z(n7182) );
  XNOR U6572 ( .A(n7184), .B(n7185), .Z(n3699) );
  ANDN U6573 ( .B(n6715), .A(n6716), .Z(n7184) );
  XOR U6574 ( .A(n7186), .B(n7187), .Z(n6649) );
  XOR U6575 ( .A(n4862), .B(n4012), .Z(n7187) );
  XOR U6576 ( .A(n7188), .B(n6691), .Z(n4012) );
  AND U6577 ( .A(n7124), .B(n7189), .Z(n7188) );
  XNOR U6578 ( .A(n7190), .B(n6704), .Z(n4862) );
  AND U6579 ( .A(n7126), .B(n7191), .Z(n7190) );
  XOR U6580 ( .A(n2572), .B(n7192), .Z(n7186) );
  XOR U6581 ( .A(n3500), .B(n7193), .Z(n7192) );
  XNOR U6582 ( .A(n7194), .B(n6696), .Z(n3500) );
  AND U6583 ( .A(n7119), .B(n7195), .Z(n7194) );
  XNOR U6584 ( .A(n7196), .B(n6687), .Z(n2572) );
  XNOR U6585 ( .A(n2345), .B(n7198), .Z(n1052) );
  XOR U6586 ( .A(n7199), .B(n5940), .Z(out[1061]) );
  XNOR U6587 ( .A(n7200), .B(n5809), .Z(n5940) );
  XOR U6588 ( .A(n7201), .B(n6072), .Z(n5809) );
  XNOR U6589 ( .A(n7202), .B(n7203), .Z(n6072) );
  XOR U6590 ( .A(n5336), .B(n3733), .Z(n7203) );
  XOR U6591 ( .A(n7204), .B(n7205), .Z(n3733) );
  ANDN U6592 ( .B(n7206), .A(n7207), .Z(n7204) );
  XOR U6593 ( .A(n7208), .B(n7209), .Z(n5336) );
  ANDN U6594 ( .B(n7210), .A(n7211), .Z(n7208) );
  XNOR U6595 ( .A(n6176), .B(n7212), .Z(n7202) );
  XOR U6596 ( .A(n4320), .B(n2613), .Z(n7212) );
  XNOR U6597 ( .A(n7213), .B(n7214), .Z(n2613) );
  ANDN U6598 ( .B(n7215), .A(n7216), .Z(n7213) );
  XOR U6599 ( .A(n7217), .B(n7218), .Z(n4320) );
  ANDN U6600 ( .B(n7219), .A(n7220), .Z(n7217) );
  XNOR U6601 ( .A(n7221), .B(n7222), .Z(n6176) );
  ANDN U6602 ( .B(n7223), .A(n7224), .Z(n7221) );
  ANDN U6603 ( .B(n1056), .A(n1057), .Z(n7199) );
  XNOR U6604 ( .A(n1803), .B(n7225), .Z(n1057) );
  XNOR U6605 ( .A(n2352), .B(n7226), .Z(n1056) );
  XOR U6606 ( .A(n7227), .B(n5945), .Z(out[1060]) );
  XNOR U6607 ( .A(n7228), .B(n5836), .Z(n5945) );
  XOR U6608 ( .A(n7229), .B(n6076), .Z(n5836) );
  XNOR U6609 ( .A(n7230), .B(n7231), .Z(n6076) );
  XOR U6610 ( .A(n5341), .B(n3737), .Z(n7231) );
  XOR U6611 ( .A(n7232), .B(n7233), .Z(n3737) );
  ANDN U6612 ( .B(n7234), .A(n7235), .Z(n7232) );
  XOR U6613 ( .A(n7236), .B(n7237), .Z(n5341) );
  ANDN U6614 ( .B(n7238), .A(n7239), .Z(n7236) );
  XNOR U6615 ( .A(n6181), .B(n7240), .Z(n7230) );
  XOR U6616 ( .A(n2624), .B(n4325), .Z(n7240) );
  XOR U6617 ( .A(n7241), .B(n7242), .Z(n4325) );
  ANDN U6618 ( .B(n7243), .A(n7244), .Z(n7241) );
  XNOR U6619 ( .A(n7245), .B(n7246), .Z(n2624) );
  ANDN U6620 ( .B(n7247), .A(n7248), .Z(n7245) );
  XNOR U6621 ( .A(n7249), .B(n7250), .Z(n6181) );
  ANDN U6622 ( .B(n7251), .A(n7252), .Z(n7249) );
  ANDN U6623 ( .B(n1060), .A(n1062), .Z(n7227) );
  XNOR U6624 ( .A(n1807), .B(n7253), .Z(n1062) );
  IV U6625 ( .A(n5189), .Z(n1807) );
  XOR U6626 ( .A(n6707), .B(n6423), .Z(n5189) );
  XOR U6627 ( .A(n7254), .B(n7255), .Z(n6423) );
  XOR U6628 ( .A(n5992), .B(n4273), .Z(n7255) );
  XOR U6629 ( .A(n7256), .B(n7257), .Z(n4273) );
  XNOR U6630 ( .A(n7258), .B(n7259), .Z(n5992) );
  ANDN U6631 ( .B(n7260), .A(n6788), .Z(n7258) );
  XOR U6632 ( .A(n3708), .B(n7261), .Z(n7254) );
  XOR U6633 ( .A(n5511), .B(n2163), .Z(n7261) );
  XNOR U6634 ( .A(n7262), .B(n7263), .Z(n2163) );
  ANDN U6635 ( .B(n7264), .A(n6784), .Z(n7262) );
  XNOR U6636 ( .A(n7265), .B(n7266), .Z(n5511) );
  XNOR U6637 ( .A(n7267), .B(n7268), .Z(n3708) );
  NOR U6638 ( .A(n6771), .B(n6780), .Z(n7267) );
  XOR U6639 ( .A(n7269), .B(n7270), .Z(n6707) );
  XOR U6640 ( .A(n4872), .B(n4020), .Z(n7270) );
  XOR U6641 ( .A(n7271), .B(n6743), .Z(n4020) );
  ANDN U6642 ( .B(n7272), .A(n7273), .Z(n7271) );
  XNOR U6643 ( .A(n7274), .B(n6756), .Z(n4872) );
  ANDN U6644 ( .B(n7275), .A(n7276), .Z(n7274) );
  XOR U6645 ( .A(n2586), .B(n7277), .Z(n7269) );
  XOR U6646 ( .A(n3505), .B(n7278), .Z(n7277) );
  XNOR U6647 ( .A(n7279), .B(n6748), .Z(n3505) );
  ANDN U6648 ( .B(n7280), .A(n7281), .Z(n7279) );
  XNOR U6649 ( .A(n7282), .B(n6739), .Z(n2586) );
  ANDN U6650 ( .B(n7283), .A(n7284), .Z(n7282) );
  XNOR U6651 ( .A(n2359), .B(n7285), .Z(n1060) );
  XOR U6652 ( .A(n7286), .B(n4119), .Z(out[105]) );
  IV U6653 ( .A(n4292), .Z(n4119) );
  XOR U6654 ( .A(n6981), .B(n2557), .Z(n4292) );
  XNOR U6655 ( .A(n7287), .B(n7288), .Z(n2557) );
  XOR U6656 ( .A(n7289), .B(n7290), .Z(n6981) );
  ANDN U6657 ( .B(n7291), .A(n7292), .Z(n7289) );
  ANDN U6658 ( .B(n3466), .A(n3468), .Z(n7286) );
  XNOR U6659 ( .A(n7293), .B(n2330), .Z(n3468) );
  XOR U6660 ( .A(n7294), .B(n2395), .Z(n3466) );
  XOR U6661 ( .A(n7295), .B(n5950), .Z(out[1059]) );
  XNOR U6662 ( .A(n7296), .B(n5867), .Z(n5950) );
  XOR U6663 ( .A(n7297), .B(n6082), .Z(n5867) );
  XNOR U6664 ( .A(n7298), .B(n7299), .Z(n6082) );
  XNOR U6665 ( .A(n5346), .B(n3741), .Z(n7299) );
  XOR U6666 ( .A(n7300), .B(n7301), .Z(n3741) );
  ANDN U6667 ( .B(n7302), .A(n7303), .Z(n7300) );
  XNOR U6668 ( .A(n7304), .B(n7305), .Z(n5346) );
  ANDN U6669 ( .B(n7306), .A(n7307), .Z(n7304) );
  XNOR U6670 ( .A(n6186), .B(n7308), .Z(n7298) );
  XOR U6671 ( .A(n2631), .B(n4332), .Z(n7308) );
  XNOR U6672 ( .A(n7309), .B(n7310), .Z(n4332) );
  ANDN U6673 ( .B(n7311), .A(n7312), .Z(n7309) );
  XNOR U6674 ( .A(n7313), .B(n7314), .Z(n2631) );
  NOR U6675 ( .A(n7315), .B(n7316), .Z(n7313) );
  XNOR U6676 ( .A(n7317), .B(n7318), .Z(n6186) );
  ANDN U6677 ( .B(n7319), .A(n7320), .Z(n7317) );
  ANDN U6678 ( .B(n1064), .A(n1065), .Z(n7295) );
  XNOR U6679 ( .A(n1811), .B(n7321), .Z(n1065) );
  IV U6680 ( .A(n5192), .Z(n1811) );
  XOR U6681 ( .A(n6733), .B(n6427), .Z(n5192) );
  XOR U6682 ( .A(n7322), .B(n7323), .Z(n6427) );
  XOR U6683 ( .A(n5997), .B(n4276), .Z(n7323) );
  XOR U6684 ( .A(n7324), .B(n7325), .Z(n4276) );
  ANDN U6685 ( .B(n6813), .A(n6814), .Z(n7324) );
  XNOR U6686 ( .A(n7326), .B(n7327), .Z(n5997) );
  ANDN U6687 ( .B(n6796), .A(n6797), .Z(n7326) );
  XOR U6688 ( .A(n3712), .B(n7328), .Z(n7322) );
  XOR U6689 ( .A(n5515), .B(n2167), .Z(n7328) );
  XNOR U6690 ( .A(n7329), .B(n7330), .Z(n2167) );
  ANDN U6691 ( .B(n6805), .A(n6806), .Z(n7329) );
  XNOR U6692 ( .A(n7331), .B(n7332), .Z(n5515) );
  AND U6693 ( .A(n6811), .B(n6809), .Z(n7331) );
  XNOR U6694 ( .A(n7333), .B(n7334), .Z(n3712) );
  ANDN U6695 ( .B(n6800), .A(n6801), .Z(n7333) );
  XOR U6696 ( .A(n7335), .B(n7336), .Z(n6733) );
  XOR U6697 ( .A(n4875), .B(n4023), .Z(n7336) );
  XOR U6698 ( .A(n7337), .B(n6781), .Z(n4023) );
  ANDN U6699 ( .B(n7338), .A(n7268), .Z(n7337) );
  XNOR U6700 ( .A(n7339), .B(n6769), .Z(n4875) );
  ANDN U6701 ( .B(n7340), .A(n7257), .Z(n7339) );
  XOR U6702 ( .A(n2593), .B(n7341), .Z(n7335) );
  XOR U6703 ( .A(n3508), .B(n7342), .Z(n7341) );
  XNOR U6704 ( .A(n7343), .B(n6785), .Z(n3508) );
  ANDN U6705 ( .B(n7344), .A(n7263), .Z(n7343) );
  XNOR U6706 ( .A(n7345), .B(n6789), .Z(n2593) );
  ANDN U6707 ( .B(n7346), .A(n7259), .Z(n7345) );
  XNOR U6708 ( .A(n2366), .B(n7347), .Z(n1064) );
  XOR U6709 ( .A(n7348), .B(n5955), .Z(out[1058]) );
  XNOR U6710 ( .A(n7349), .B(n5902), .Z(n5955) );
  XOR U6711 ( .A(n7350), .B(n6088), .Z(n5902) );
  XNOR U6712 ( .A(n7351), .B(n7352), .Z(n6088) );
  XNOR U6713 ( .A(n5350), .B(n3746), .Z(n7352) );
  XOR U6714 ( .A(n7353), .B(n7354), .Z(n3746) );
  ANDN U6715 ( .B(n7355), .A(n7356), .Z(n7353) );
  XNOR U6716 ( .A(n7357), .B(n7358), .Z(n5350) );
  ANDN U6717 ( .B(n7359), .A(n7360), .Z(n7357) );
  XNOR U6718 ( .A(n6191), .B(n7361), .Z(n7351) );
  XOR U6719 ( .A(n2638), .B(n4386), .Z(n7361) );
  XNOR U6720 ( .A(n7362), .B(n7363), .Z(n4386) );
  ANDN U6721 ( .B(n7364), .A(n7365), .Z(n7362) );
  XNOR U6722 ( .A(n7366), .B(n7367), .Z(n2638) );
  ANDN U6723 ( .B(n7368), .A(n7369), .Z(n7366) );
  XNOR U6724 ( .A(n7370), .B(n7371), .Z(n6191) );
  ANDN U6725 ( .B(n7372), .A(n7373), .Z(n7370) );
  ANDN U6726 ( .B(n1068), .A(n1069), .Z(n7348) );
  XNOR U6727 ( .A(n1823), .B(n7374), .Z(n1069) );
  IV U6728 ( .A(n5196), .Z(n1823) );
  XOR U6729 ( .A(n6759), .B(n6431), .Z(n5196) );
  XOR U6730 ( .A(n7375), .B(n7376), .Z(n6431) );
  XOR U6731 ( .A(n6002), .B(n5528), .Z(n7376) );
  XOR U6732 ( .A(n7377), .B(n7378), .Z(n5528) );
  ANDN U6733 ( .B(n6835), .A(n6836), .Z(n7377) );
  XNOR U6734 ( .A(n7379), .B(n7380), .Z(n6002) );
  ANDN U6735 ( .B(n6822), .A(n6823), .Z(n7379) );
  XOR U6736 ( .A(n3716), .B(n7381), .Z(n7375) );
  XOR U6737 ( .A(n4279), .B(n2171), .Z(n7381) );
  XNOR U6738 ( .A(n7382), .B(n7383), .Z(n2171) );
  ANDN U6739 ( .B(n6831), .A(n6832), .Z(n7382) );
  XNOR U6740 ( .A(n7384), .B(n7385), .Z(n4279) );
  ANDN U6741 ( .B(n6839), .A(n6840), .Z(n7384) );
  XNOR U6742 ( .A(n7386), .B(n7387), .Z(n3716) );
  ANDN U6743 ( .B(n6826), .A(n6827), .Z(n7386) );
  XOR U6744 ( .A(n7388), .B(n7389), .Z(n6759) );
  XOR U6745 ( .A(n4878), .B(n4026), .Z(n7389) );
  XOR U6746 ( .A(n7390), .B(n6802), .Z(n4026) );
  NOR U6747 ( .A(n7391), .B(n7334), .Z(n7390) );
  XNOR U6748 ( .A(n7392), .B(n6815), .Z(n4878) );
  NOR U6749 ( .A(n7393), .B(n7325), .Z(n7392) );
  XOR U6750 ( .A(n2600), .B(n7394), .Z(n7388) );
  XOR U6751 ( .A(n3511), .B(n7395), .Z(n7394) );
  XNOR U6752 ( .A(n7396), .B(n6807), .Z(n3511) );
  NOR U6753 ( .A(n7397), .B(n7330), .Z(n7396) );
  XNOR U6754 ( .A(n7398), .B(n6798), .Z(n2600) );
  NOR U6755 ( .A(n7399), .B(n7327), .Z(n7398) );
  XNOR U6756 ( .A(n2371), .B(n7400), .Z(n1068) );
  IV U6757 ( .A(n5007), .Z(n2371) );
  XOR U6758 ( .A(n6279), .B(n7401), .Z(n5007) );
  XOR U6759 ( .A(n7402), .B(n7403), .Z(n6279) );
  XOR U6760 ( .A(n3216), .B(n7404), .Z(n7403) );
  XNOR U6761 ( .A(n7405), .B(n7406), .Z(n3216) );
  ANDN U6762 ( .B(n7407), .A(n7408), .Z(n7405) );
  XOR U6763 ( .A(n5538), .B(n7409), .Z(n7402) );
  XOR U6764 ( .A(n7410), .B(n2412), .Z(n7409) );
  XNOR U6765 ( .A(n7411), .B(n7412), .Z(n2412) );
  NOR U6766 ( .A(n7413), .B(n7414), .Z(n7411) );
  XNOR U6767 ( .A(n7415), .B(n7416), .Z(n5538) );
  NOR U6768 ( .A(n7417), .B(n7418), .Z(n7415) );
  XOR U6769 ( .A(n7419), .B(n5960), .Z(out[1057]) );
  XNOR U6770 ( .A(n7420), .B(n5935), .Z(n5960) );
  XOR U6771 ( .A(n7421), .B(n6093), .Z(n5935) );
  XNOR U6772 ( .A(n7422), .B(n7423), .Z(n6093) );
  XNOR U6773 ( .A(n5354), .B(n3750), .Z(n7423) );
  XOR U6774 ( .A(n7424), .B(n7425), .Z(n3750) );
  AND U6775 ( .A(n7426), .B(n7427), .Z(n7424) );
  XNOR U6776 ( .A(n7428), .B(n7429), .Z(n5354) );
  ANDN U6777 ( .B(n7430), .A(n7431), .Z(n7428) );
  XNOR U6778 ( .A(n6196), .B(n7432), .Z(n7422) );
  XOR U6779 ( .A(n2645), .B(n4430), .Z(n7432) );
  XOR U6780 ( .A(n7433), .B(n7434), .Z(n4430) );
  ANDN U6781 ( .B(n7435), .A(n7436), .Z(n7433) );
  XNOR U6782 ( .A(n7437), .B(n7438), .Z(n2645) );
  ANDN U6783 ( .B(n7439), .A(n7440), .Z(n7437) );
  XNOR U6784 ( .A(n7441), .B(n7442), .Z(n6196) );
  AND U6785 ( .A(n7443), .B(n7444), .Z(n7441) );
  ANDN U6786 ( .B(n1072), .A(n1073), .Z(n7419) );
  XNOR U6787 ( .A(n1827), .B(n7445), .Z(n1073) );
  IV U6788 ( .A(n5200), .Z(n1827) );
  XOR U6789 ( .A(n6792), .B(n6435), .Z(n5200) );
  XOR U6790 ( .A(n7446), .B(n7447), .Z(n6435) );
  XOR U6791 ( .A(n6007), .B(n5532), .Z(n7447) );
  XOR U6792 ( .A(n7448), .B(n7449), .Z(n5532) );
  AND U6793 ( .A(n6863), .B(n6861), .Z(n7448) );
  XNOR U6794 ( .A(n7450), .B(n7451), .Z(n6007) );
  ANDN U6795 ( .B(n6848), .A(n6850), .Z(n7450) );
  XOR U6796 ( .A(n3720), .B(n7452), .Z(n7446) );
  XOR U6797 ( .A(n4282), .B(n2174), .Z(n7452) );
  XNOR U6798 ( .A(n7453), .B(n7454), .Z(n2174) );
  ANDN U6799 ( .B(n6857), .A(n6858), .Z(n7453) );
  XNOR U6800 ( .A(n7455), .B(n7456), .Z(n4282) );
  ANDN U6801 ( .B(n6865), .A(n6866), .Z(n7455) );
  XNOR U6802 ( .A(n7457), .B(n7458), .Z(n3720) );
  ANDN U6803 ( .B(n6852), .A(n6853), .Z(n7457) );
  XOR U6804 ( .A(n7459), .B(n7460), .Z(n6792) );
  XOR U6805 ( .A(n4881), .B(n4031), .Z(n7460) );
  XOR U6806 ( .A(n7461), .B(n6828), .Z(n4031) );
  ANDN U6807 ( .B(n7462), .A(n7387), .Z(n7461) );
  XNOR U6808 ( .A(n7463), .B(n6841), .Z(n4881) );
  ANDN U6809 ( .B(n7464), .A(n7385), .Z(n7463) );
  XOR U6810 ( .A(n2607), .B(n7465), .Z(n7459) );
  XOR U6811 ( .A(n3514), .B(n7466), .Z(n7465) );
  XNOR U6812 ( .A(n7467), .B(n6833), .Z(n3514) );
  ANDN U6813 ( .B(n7468), .A(n7383), .Z(n7467) );
  XNOR U6814 ( .A(n7469), .B(n6824), .Z(n2607) );
  ANDN U6815 ( .B(n7470), .A(n7380), .Z(n7469) );
  XNOR U6816 ( .A(n2380), .B(n7471), .Z(n1072) );
  IV U6817 ( .A(n5011), .Z(n2380) );
  XOR U6818 ( .A(n6284), .B(n7472), .Z(n5011) );
  XOR U6819 ( .A(n7473), .B(n7474), .Z(n6284) );
  XNOR U6820 ( .A(n3219), .B(n7475), .Z(n7474) );
  XNOR U6821 ( .A(n7476), .B(n7477), .Z(n3219) );
  ANDN U6822 ( .B(n7478), .A(n7479), .Z(n7476) );
  XOR U6823 ( .A(n5541), .B(n7480), .Z(n7473) );
  XOR U6824 ( .A(n7481), .B(n2419), .Z(n7480) );
  XNOR U6825 ( .A(n7482), .B(n7483), .Z(n2419) );
  ANDN U6826 ( .B(n7484), .A(n7485), .Z(n7482) );
  XNOR U6827 ( .A(n7486), .B(n7487), .Z(n5541) );
  ANDN U6828 ( .B(n7488), .A(n7489), .Z(n7486) );
  XOR U6829 ( .A(n7490), .B(n5965), .Z(out[1056]) );
  XNOR U6830 ( .A(n7491), .B(n5990), .Z(n5965) );
  XOR U6831 ( .A(n7492), .B(n6100), .Z(n5990) );
  XNOR U6832 ( .A(n7493), .B(n7494), .Z(n6100) );
  XNOR U6833 ( .A(n5358), .B(n3754), .Z(n7494) );
  XOR U6834 ( .A(n7495), .B(n7496), .Z(n3754) );
  ANDN U6835 ( .B(n7497), .A(n7498), .Z(n7495) );
  XNOR U6836 ( .A(n7499), .B(n7500), .Z(n5358) );
  ANDN U6837 ( .B(n7501), .A(n7502), .Z(n7499) );
  XNOR U6838 ( .A(n6201), .B(n7503), .Z(n7493) );
  XOR U6839 ( .A(n2652), .B(n4474), .Z(n7503) );
  XOR U6840 ( .A(n7504), .B(n7505), .Z(n4474) );
  ANDN U6841 ( .B(n7506), .A(n7507), .Z(n7504) );
  XNOR U6842 ( .A(n7508), .B(n7509), .Z(n2652) );
  ANDN U6843 ( .B(n7510), .A(n7511), .Z(n7508) );
  XNOR U6844 ( .A(n7512), .B(n7513), .Z(n6201) );
  AND U6845 ( .A(n7514), .B(n7515), .Z(n7512) );
  NOR U6846 ( .A(n1077), .B(n1076), .Z(n7490) );
  XOR U6847 ( .A(n7516), .B(n2387), .Z(n1076) );
  XOR U6848 ( .A(n7517), .B(n7518), .Z(n6289) );
  XNOR U6849 ( .A(n3222), .B(n7519), .Z(n7518) );
  XNOR U6850 ( .A(n7520), .B(n7521), .Z(n3222) );
  ANDN U6851 ( .B(n7522), .A(n7523), .Z(n7520) );
  XOR U6852 ( .A(n5546), .B(n7524), .Z(n7517) );
  XOR U6853 ( .A(n7525), .B(n2426), .Z(n7524) );
  XNOR U6854 ( .A(n7526), .B(n7527), .Z(n2426) );
  ANDN U6855 ( .B(n7528), .A(n7529), .Z(n7526) );
  XNOR U6856 ( .A(n7530), .B(n7531), .Z(n5546) );
  ANDN U6857 ( .B(n7532), .A(n7533), .Z(n7530) );
  XNOR U6858 ( .A(n1831), .B(n7535), .Z(n1077) );
  IV U6859 ( .A(n5209), .Z(n1831) );
  XOR U6860 ( .A(n6818), .B(n6449), .Z(n5209) );
  XOR U6861 ( .A(n7536), .B(n7537), .Z(n6449) );
  XOR U6862 ( .A(n6012), .B(n5536), .Z(n7537) );
  XOR U6863 ( .A(n7538), .B(n7539), .Z(n5536) );
  AND U6864 ( .A(n6895), .B(n6893), .Z(n7538) );
  XNOR U6865 ( .A(n7540), .B(n7541), .Z(n6012) );
  ANDN U6866 ( .B(n6874), .A(n6876), .Z(n7540) );
  XOR U6867 ( .A(n3724), .B(n7542), .Z(n7536) );
  XOR U6868 ( .A(n4285), .B(n2177), .Z(n7542) );
  XOR U6869 ( .A(n7543), .B(n7544), .Z(n2177) );
  XNOR U6870 ( .A(n7545), .B(n7546), .Z(n4285) );
  ANDN U6871 ( .B(n6897), .A(n6899), .Z(n7545) );
  XNOR U6872 ( .A(n7547), .B(n7548), .Z(n3724) );
  ANDN U6873 ( .B(n6877), .A(n6885), .Z(n7547) );
  IV U6874 ( .A(n7549), .Z(n6877) );
  XOR U6875 ( .A(n7550), .B(n7551), .Z(n6818) );
  XOR U6876 ( .A(n4884), .B(n4034), .Z(n7551) );
  XOR U6877 ( .A(n7552), .B(n6854), .Z(n4034) );
  NOR U6878 ( .A(n7553), .B(n7458), .Z(n7552) );
  XNOR U6879 ( .A(n7554), .B(n6867), .Z(n4884) );
  ANDN U6880 ( .B(n7555), .A(n7456), .Z(n7554) );
  XOR U6881 ( .A(n2614), .B(n7556), .Z(n7550) );
  XOR U6882 ( .A(n3517), .B(n7557), .Z(n7556) );
  XNOR U6883 ( .A(n7558), .B(n6859), .Z(n3517) );
  ANDN U6884 ( .B(n7559), .A(n7454), .Z(n7558) );
  XOR U6885 ( .A(n7560), .B(n6849), .Z(n2614) );
  XOR U6886 ( .A(n7562), .B(n5970), .Z(out[1055]) );
  XOR U6887 ( .A(n7563), .B(n6048), .Z(n5970) );
  XOR U6888 ( .A(n7564), .B(n6111), .Z(n6048) );
  XNOR U6889 ( .A(n7565), .B(n7566), .Z(n6111) );
  XNOR U6890 ( .A(n5363), .B(n3758), .Z(n7566) );
  XOR U6891 ( .A(n7567), .B(n7568), .Z(n3758) );
  ANDN U6892 ( .B(n7569), .A(n7570), .Z(n7567) );
  XNOR U6893 ( .A(n7571), .B(n7572), .Z(n5363) );
  ANDN U6894 ( .B(n7573), .A(n7574), .Z(n7571) );
  XNOR U6895 ( .A(n6206), .B(n7575), .Z(n7565) );
  XOR U6896 ( .A(n2659), .B(n4525), .Z(n7575) );
  XOR U6897 ( .A(n7576), .B(n7577), .Z(n4525) );
  ANDN U6898 ( .B(n7578), .A(n7579), .Z(n7576) );
  XNOR U6899 ( .A(n7580), .B(n7581), .Z(n2659) );
  ANDN U6900 ( .B(n7582), .A(n7583), .Z(n7580) );
  XNOR U6901 ( .A(n7584), .B(n7585), .Z(n6206) );
  AND U6902 ( .A(n7586), .B(n7587), .Z(n7584) );
  ANDN U6903 ( .B(n1080), .A(n1081), .Z(n7562) );
  XNOR U6904 ( .A(n1835), .B(n7588), .Z(n1081) );
  IV U6905 ( .A(n5213), .Z(n1835) );
  XOR U6906 ( .A(n6844), .B(n6675), .Z(n5213) );
  XOR U6907 ( .A(n7589), .B(n7590), .Z(n6675) );
  XOR U6908 ( .A(n6017), .B(n2180), .Z(n7590) );
  XOR U6909 ( .A(n7591), .B(n7592), .Z(n2180) );
  ANDN U6910 ( .B(n6915), .A(n6917), .Z(n7591) );
  XNOR U6911 ( .A(n7593), .B(n7594), .Z(n6017) );
  ANDN U6912 ( .B(n6906), .A(n6908), .Z(n7593) );
  XOR U6913 ( .A(n3730), .B(n7595), .Z(n7589) );
  XOR U6914 ( .A(n4291), .B(n5540), .Z(n7595) );
  XNOR U6915 ( .A(n7596), .B(n7597), .Z(n5540) );
  AND U6916 ( .A(n6921), .B(n6919), .Z(n7596) );
  XNOR U6917 ( .A(n7598), .B(n7599), .Z(n4291) );
  AND U6918 ( .A(n6925), .B(n6923), .Z(n7598) );
  XNOR U6919 ( .A(n7600), .B(n7601), .Z(n3730) );
  ANDN U6920 ( .B(n6910), .A(n6911), .Z(n7600) );
  XOR U6921 ( .A(n7602), .B(n7603), .Z(n6844) );
  XOR U6922 ( .A(n4887), .B(n4202), .Z(n7603) );
  XOR U6923 ( .A(n7604), .B(n6886), .Z(n4202) );
  NOR U6924 ( .A(n7605), .B(n7548), .Z(n7604) );
  XOR U6925 ( .A(n7606), .B(n6898), .Z(n4887) );
  XOR U6926 ( .A(n2626), .B(n7608), .Z(n7602) );
  XOR U6927 ( .A(n3519), .B(n7609), .Z(n7608) );
  XOR U6928 ( .A(n7610), .B(n6890), .Z(n3519) );
  AND U6929 ( .A(n7544), .B(n7611), .Z(n7610) );
  XOR U6930 ( .A(n7612), .B(n6875), .Z(n2626) );
  XNOR U6931 ( .A(n2392), .B(n7614), .Z(n1080) );
  IV U6932 ( .A(n5019), .Z(n2392) );
  XOR U6933 ( .A(n6293), .B(n7615), .Z(n5019) );
  XOR U6934 ( .A(n7616), .B(n7617), .Z(n6293) );
  XNOR U6935 ( .A(n3225), .B(n7618), .Z(n7617) );
  XNOR U6936 ( .A(n7619), .B(n7620), .Z(n3225) );
  ANDN U6937 ( .B(n7621), .A(n7622), .Z(n7619) );
  XOR U6938 ( .A(n5549), .B(n7623), .Z(n7616) );
  XOR U6939 ( .A(n7624), .B(n2433), .Z(n7623) );
  XNOR U6940 ( .A(n7625), .B(n7626), .Z(n2433) );
  AND U6941 ( .A(n7627), .B(n7628), .Z(n7625) );
  XNOR U6942 ( .A(n7629), .B(n7630), .Z(n5549) );
  ANDN U6943 ( .B(n7631), .A(n7632), .Z(n7629) );
  XOR U6944 ( .A(n7633), .B(n5975), .Z(out[1054]) );
  XNOR U6945 ( .A(n7634), .B(n6107), .Z(n5975) );
  XOR U6946 ( .A(n7635), .B(n6116), .Z(n6107) );
  XNOR U6947 ( .A(n7636), .B(n7637), .Z(n6116) );
  XNOR U6948 ( .A(n5372), .B(n3762), .Z(n7637) );
  XOR U6949 ( .A(n7638), .B(n7639), .Z(n3762) );
  ANDN U6950 ( .B(n7640), .A(n7641), .Z(n7638) );
  XNOR U6951 ( .A(n7642), .B(n7643), .Z(n5372) );
  ANDN U6952 ( .B(n7644), .A(n7645), .Z(n7642) );
  XNOR U6953 ( .A(n6211), .B(n7646), .Z(n7636) );
  XOR U6954 ( .A(n2666), .B(n4576), .Z(n7646) );
  XOR U6955 ( .A(n7647), .B(n7648), .Z(n4576) );
  XOR U6956 ( .A(n7651), .B(n7652), .Z(n2666) );
  ANDN U6957 ( .B(n7653), .A(n7654), .Z(n7651) );
  XOR U6958 ( .A(n7655), .B(n7656), .Z(n6211) );
  ANDN U6959 ( .B(n7657), .A(n7658), .Z(n7655) );
  ANDN U6960 ( .B(n1084), .A(n1085), .Z(n7633) );
  XNOR U6961 ( .A(n1839), .B(n7659), .Z(n1085) );
  IV U6962 ( .A(n5217), .Z(n1839) );
  XOR U6963 ( .A(n6870), .B(n6954), .Z(n5217) );
  XOR U6964 ( .A(n7660), .B(n7661), .Z(n6954) );
  XOR U6965 ( .A(n6022), .B(n2183), .Z(n7661) );
  XOR U6966 ( .A(n7662), .B(n7663), .Z(n2183) );
  ANDN U6967 ( .B(n6957), .A(n6958), .Z(n7662) );
  XNOR U6968 ( .A(n7664), .B(n7665), .Z(n6022) );
  ANDN U6969 ( .B(n6932), .A(n6934), .Z(n7664) );
  XOR U6970 ( .A(n3734), .B(n7666), .Z(n7660) );
  XOR U6971 ( .A(n4294), .B(n5544), .Z(n7666) );
  XNOR U6972 ( .A(n7667), .B(n7668), .Z(n5544) );
  AND U6973 ( .A(n6948), .B(n6946), .Z(n7667) );
  ANDN U6974 ( .B(n6950), .A(n6951), .Z(n7669) );
  XNOR U6975 ( .A(n7671), .B(n7672), .Z(n3734) );
  ANDN U6976 ( .B(n6935), .A(n6941), .Z(n7671) );
  XOR U6977 ( .A(n7673), .B(n7674), .Z(n6870) );
  XOR U6978 ( .A(n4890), .B(n7675), .Z(n7674) );
  XNOR U6979 ( .A(n7676), .B(n6924), .Z(n4890) );
  ANDN U6980 ( .B(n7677), .A(n7599), .Z(n7676) );
  XOR U6981 ( .A(n2633), .B(n7678), .Z(n7673) );
  XOR U6982 ( .A(n3521), .B(n7679), .Z(n7678) );
  XOR U6983 ( .A(n7680), .B(n6916), .Z(n3521) );
  ANDN U6984 ( .B(n7681), .A(n7592), .Z(n7680) );
  XOR U6985 ( .A(n7682), .B(n6907), .Z(n2633) );
  XNOR U6986 ( .A(n2405), .B(n7684), .Z(n1084) );
  IV U6987 ( .A(n5023), .Z(n2405) );
  XOR U6988 ( .A(n6297), .B(n7685), .Z(n5023) );
  XOR U6989 ( .A(n7686), .B(n7687), .Z(n6297) );
  XNOR U6990 ( .A(n7688), .B(n3228), .Z(n7687) );
  XOR U6991 ( .A(n7689), .B(n7690), .Z(n3228) );
  ANDN U6992 ( .B(n7691), .A(n7692), .Z(n7689) );
  XNOR U6993 ( .A(n2439), .B(n7693), .Z(n7686) );
  XOR U6994 ( .A(n4311), .B(n5553), .Z(n7693) );
  XOR U6995 ( .A(n7694), .B(n7695), .Z(n5553) );
  ANDN U6996 ( .B(n7696), .A(n7697), .Z(n7694) );
  XOR U6997 ( .A(n7698), .B(n7699), .Z(n4311) );
  ANDN U6998 ( .B(n7700), .A(n7701), .Z(n7698) );
  XOR U6999 ( .A(n7702), .B(n7703), .Z(n2439) );
  AND U7000 ( .A(n7704), .B(n7705), .Z(n7702) );
  XOR U7001 ( .A(n7706), .B(n5980), .Z(out[1053]) );
  XNOR U7002 ( .A(n7707), .B(n6164), .Z(n5980) );
  XOR U7003 ( .A(n7708), .B(n6122), .Z(n6164) );
  XNOR U7004 ( .A(n7709), .B(n7710), .Z(n6122) );
  XNOR U7005 ( .A(n5377), .B(n3766), .Z(n7710) );
  XNOR U7006 ( .A(n7711), .B(n7712), .Z(n3766) );
  AND U7007 ( .A(n7713), .B(n7714), .Z(n7711) );
  XNOR U7008 ( .A(n7715), .B(n7716), .Z(n5377) );
  ANDN U7009 ( .B(n7717), .A(n7718), .Z(n7715) );
  XNOR U7010 ( .A(n6221), .B(n7719), .Z(n7709) );
  XOR U7011 ( .A(n2673), .B(n4627), .Z(n7719) );
  XOR U7012 ( .A(n7720), .B(n7721), .Z(n4627) );
  AND U7013 ( .A(n7722), .B(n7723), .Z(n7720) );
  XOR U7014 ( .A(n7724), .B(n7725), .Z(n2673) );
  ANDN U7015 ( .B(n7726), .A(n7727), .Z(n7724) );
  XNOR U7016 ( .A(n7728), .B(n7729), .Z(n6221) );
  ANDN U7017 ( .B(n7730), .A(n7731), .Z(n7728) );
  ANDN U7018 ( .B(n1092), .A(n1093), .Z(n7706) );
  XNOR U7019 ( .A(n1843), .B(n7732), .Z(n1093) );
  IV U7020 ( .A(n5220), .Z(n1843) );
  XOR U7021 ( .A(n6902), .B(n7287), .Z(n5220) );
  XOR U7022 ( .A(n7733), .B(n7734), .Z(n7287) );
  XOR U7023 ( .A(n6027), .B(n2187), .Z(n7734) );
  XOR U7024 ( .A(n7735), .B(n7736), .Z(n2187) );
  ANDN U7025 ( .B(n7290), .A(n7291), .Z(n7735) );
  XNOR U7026 ( .A(n7737), .B(n7738), .Z(n6027) );
  ANDN U7027 ( .B(n6968), .A(n6970), .Z(n7737) );
  XOR U7028 ( .A(n5548), .B(n7739), .Z(n7733) );
  XOR U7029 ( .A(n4298), .B(n3738), .Z(n7739) );
  XNOR U7030 ( .A(n7740), .B(n7741), .Z(n3738) );
  ANDN U7031 ( .B(n6971), .A(n6979), .Z(n7740) );
  IV U7032 ( .A(n7742), .Z(n6971) );
  XNOR U7033 ( .A(n7743), .B(n7744), .Z(n4298) );
  ANDN U7034 ( .B(n6987), .A(n6988), .Z(n7743) );
  XNOR U7035 ( .A(n7745), .B(n7746), .Z(n5548) );
  AND U7036 ( .A(n6985), .B(n6983), .Z(n7745) );
  XOR U7037 ( .A(n7747), .B(n7748), .Z(n6902) );
  XOR U7038 ( .A(n4893), .B(n5618), .Z(n7748) );
  XOR U7039 ( .A(n7749), .B(n6942), .Z(n5618) );
  NOR U7040 ( .A(n7750), .B(n7672), .Z(n7749) );
  XNOR U7041 ( .A(n7751), .B(n6952), .Z(n4893) );
  NOR U7042 ( .A(n7670), .B(n7752), .Z(n7751) );
  XOR U7043 ( .A(n2640), .B(n7753), .Z(n7747) );
  XOR U7044 ( .A(n3523), .B(n7754), .Z(n7753) );
  XNOR U7045 ( .A(n7755), .B(n6959), .Z(n3523) );
  ANDN U7046 ( .B(n7756), .A(n7663), .Z(n7755) );
  XOR U7047 ( .A(n7757), .B(n6933), .Z(n2640) );
  XNOR U7048 ( .A(n7759), .B(n2411), .Z(n1092) );
  XOR U7049 ( .A(n6301), .B(n7760), .Z(n2411) );
  XOR U7050 ( .A(n7761), .B(n7762), .Z(n6301) );
  XNOR U7051 ( .A(n7763), .B(n3231), .Z(n7762) );
  XOR U7052 ( .A(n7764), .B(n7765), .Z(n3231) );
  ANDN U7053 ( .B(n7766), .A(n7767), .Z(n7764) );
  XNOR U7054 ( .A(n2446), .B(n7768), .Z(n7761) );
  XOR U7055 ( .A(n4315), .B(n5559), .Z(n7768) );
  XOR U7056 ( .A(n7769), .B(n7770), .Z(n5559) );
  ANDN U7057 ( .B(n7771), .A(n7772), .Z(n7769) );
  XOR U7058 ( .A(n7773), .B(n7774), .Z(n4315) );
  NOR U7059 ( .A(n7775), .B(n7776), .Z(n7773) );
  XNOR U7060 ( .A(n7777), .B(n7778), .Z(n2446) );
  ANDN U7061 ( .B(n7779), .A(n7780), .Z(n7777) );
  XOR U7062 ( .A(n7781), .B(n5985), .Z(out[1052]) );
  XNOR U7063 ( .A(n7782), .B(n6219), .Z(n5985) );
  XOR U7064 ( .A(n7783), .B(n6128), .Z(n6219) );
  XNOR U7065 ( .A(n7784), .B(n7785), .Z(n6128) );
  XNOR U7066 ( .A(n5383), .B(n3773), .Z(n7785) );
  XOR U7067 ( .A(n7786), .B(n7787), .Z(n3773) );
  XNOR U7068 ( .A(n7790), .B(n7791), .Z(n5383) );
  ANDN U7069 ( .B(n7792), .A(n7793), .Z(n7790) );
  XNOR U7070 ( .A(n6226), .B(n7794), .Z(n7784) );
  XOR U7071 ( .A(n2680), .B(n4677), .Z(n7794) );
  XNOR U7072 ( .A(n7795), .B(n7796), .Z(n4677) );
  ANDN U7073 ( .B(n7797), .A(n7798), .Z(n7795) );
  XOR U7074 ( .A(n7799), .B(n7800), .Z(n2680) );
  XNOR U7075 ( .A(n7803), .B(n7804), .Z(n6226) );
  NOR U7076 ( .A(n7805), .B(n7806), .Z(n7803) );
  ANDN U7077 ( .B(n1096), .A(n1098), .Z(n7781) );
  XNOR U7078 ( .A(n1847), .B(n7807), .Z(n1098) );
  IV U7079 ( .A(n5224), .Z(n1847) );
  XOR U7080 ( .A(n6928), .B(n7808), .Z(n5224) );
  XOR U7081 ( .A(n7809), .B(n7810), .Z(n6928) );
  XNOR U7082 ( .A(n4896), .B(n5664), .Z(n7810) );
  XOR U7083 ( .A(n7811), .B(n6978), .Z(n5664) );
  NOR U7084 ( .A(n7741), .B(n7812), .Z(n7811) );
  XNOR U7085 ( .A(n7813), .B(n6989), .Z(n4896) );
  NOR U7086 ( .A(n7814), .B(n7744), .Z(n7813) );
  XOR U7087 ( .A(n2647), .B(n7815), .Z(n7809) );
  XOR U7088 ( .A(n3532), .B(n7816), .Z(n7815) );
  XNOR U7089 ( .A(n7817), .B(n7292), .Z(n3532) );
  ANDN U7090 ( .B(n7818), .A(n7736), .Z(n7817) );
  XOR U7091 ( .A(n7819), .B(n6969), .Z(n2647) );
  XOR U7092 ( .A(n7821), .B(n2418), .Z(n1096) );
  XOR U7093 ( .A(n6305), .B(n7822), .Z(n2418) );
  XOR U7094 ( .A(n7823), .B(n7824), .Z(n6305) );
  XNOR U7095 ( .A(n3238), .B(n4321), .Z(n7824) );
  XOR U7096 ( .A(n7825), .B(n7826), .Z(n4321) );
  NOR U7097 ( .A(n7827), .B(n7828), .Z(n7825) );
  XOR U7098 ( .A(n7829), .B(n7830), .Z(n3238) );
  NOR U7099 ( .A(n7831), .B(n7832), .Z(n7829) );
  XOR U7100 ( .A(n5562), .B(n7833), .Z(n7823) );
  XOR U7101 ( .A(n7834), .B(n2454), .Z(n7833) );
  XOR U7102 ( .A(n7835), .B(n7836), .Z(n2454) );
  ANDN U7103 ( .B(n7837), .A(n7838), .Z(n7835) );
  XOR U7104 ( .A(n7839), .B(n7840), .Z(n5562) );
  ANDN U7105 ( .B(n7841), .A(n7842), .Z(n7839) );
  XOR U7106 ( .A(n7843), .B(n5995), .Z(out[1051]) );
  XNOR U7107 ( .A(n7844), .B(n6276), .Z(n5995) );
  XOR U7108 ( .A(n7845), .B(n6134), .Z(n6276) );
  XNOR U7109 ( .A(n7846), .B(n7847), .Z(n6134) );
  XNOR U7110 ( .A(n5387), .B(n3777), .Z(n7847) );
  XNOR U7111 ( .A(n7848), .B(n7849), .Z(n3777) );
  XNOR U7112 ( .A(n7852), .B(n7853), .Z(n5387) );
  ANDN U7113 ( .B(n7854), .A(n7855), .Z(n7852) );
  XNOR U7114 ( .A(n6231), .B(n7856), .Z(n7846) );
  XOR U7115 ( .A(n2687), .B(n4702), .Z(n7856) );
  XNOR U7116 ( .A(n7857), .B(n7858), .Z(n4702) );
  ANDN U7117 ( .B(n7859), .A(n7860), .Z(n7857) );
  XOR U7118 ( .A(n7861), .B(n7862), .Z(n2687) );
  ANDN U7119 ( .B(n7863), .A(n7864), .Z(n7861) );
  XNOR U7120 ( .A(n7865), .B(n7866), .Z(n6231) );
  ANDN U7121 ( .B(n7867), .A(n7868), .Z(n7865) );
  ANDN U7122 ( .B(n1100), .A(n1101), .Z(n7843) );
  XNOR U7123 ( .A(n1852), .B(n7869), .Z(n1101) );
  IV U7124 ( .A(n5227), .Z(n1852) );
  XOR U7125 ( .A(n6964), .B(n7870), .Z(n5227) );
  XOR U7126 ( .A(n7871), .B(n7872), .Z(n6964) );
  XOR U7127 ( .A(n4899), .B(n7873), .Z(n7872) );
  XNOR U7128 ( .A(n7874), .B(n7017), .Z(n4899) );
  NOR U7129 ( .A(n7875), .B(n7876), .Z(n7874) );
  XOR U7130 ( .A(n2654), .B(n7877), .Z(n7871) );
  XOR U7131 ( .A(n3535), .B(n5710), .Z(n7877) );
  XOR U7132 ( .A(n7878), .B(n7006), .Z(n5710) );
  ANDN U7133 ( .B(n7879), .A(n7880), .Z(n7878) );
  XNOR U7134 ( .A(n7881), .B(n7882), .Z(n3535) );
  ANDN U7135 ( .B(n7883), .A(n7884), .Z(n7881) );
  XOR U7136 ( .A(n7885), .B(n6997), .Z(n2654) );
  XNOR U7137 ( .A(n2424), .B(n7888), .Z(n1100) );
  IV U7138 ( .A(n5038), .Z(n2424) );
  XOR U7139 ( .A(n6309), .B(n7889), .Z(n5038) );
  XOR U7140 ( .A(n7890), .B(n7891), .Z(n6309) );
  XOR U7141 ( .A(n3242), .B(n4324), .Z(n7891) );
  XNOR U7142 ( .A(n7892), .B(n7893), .Z(n4324) );
  NOR U7143 ( .A(n7894), .B(n7895), .Z(n7892) );
  XOR U7144 ( .A(n7896), .B(n7897), .Z(n3242) );
  ANDN U7145 ( .B(n7898), .A(n7899), .Z(n7896) );
  XOR U7146 ( .A(n5567), .B(n7900), .Z(n7890) );
  XOR U7147 ( .A(n7901), .B(n2461), .Z(n7900) );
  XOR U7148 ( .A(n7902), .B(n7903), .Z(n2461) );
  AND U7149 ( .A(n7904), .B(n7905), .Z(n7902) );
  XOR U7150 ( .A(n7906), .B(n7907), .Z(n5567) );
  ANDN U7151 ( .B(n7908), .A(n7909), .Z(n7906) );
  XOR U7152 ( .A(n7910), .B(n6000), .Z(out[1050]) );
  XOR U7153 ( .A(n7911), .B(n2351), .Z(n6000) );
  XNOR U7154 ( .A(n7912), .B(n6140), .Z(n2351) );
  XNOR U7155 ( .A(n7913), .B(n7914), .Z(n6140) );
  XNOR U7156 ( .A(n5392), .B(n3781), .Z(n7914) );
  XOR U7157 ( .A(n7915), .B(n7916), .Z(n3781) );
  XNOR U7158 ( .A(n7919), .B(n7920), .Z(n5392) );
  ANDN U7159 ( .B(n7921), .A(n7922), .Z(n7919) );
  XNOR U7160 ( .A(n6236), .B(n7923), .Z(n7913) );
  XOR U7161 ( .A(n2218), .B(n4726), .Z(n7923) );
  XNOR U7162 ( .A(n7924), .B(n7925), .Z(n4726) );
  ANDN U7163 ( .B(n7926), .A(n7927), .Z(n7924) );
  XOR U7164 ( .A(n7928), .B(n7929), .Z(n2218) );
  ANDN U7165 ( .B(n7930), .A(n7931), .Z(n7928) );
  XNOR U7166 ( .A(n7932), .B(n7933), .Z(n6236) );
  ANDN U7167 ( .B(n7934), .A(n7935), .Z(n7932) );
  ANDN U7168 ( .B(n1104), .A(n1105), .Z(n7910) );
  XNOR U7169 ( .A(n1856), .B(n7936), .Z(n1105) );
  IV U7170 ( .A(n5230), .Z(n1856) );
  XOR U7171 ( .A(n6992), .B(n7937), .Z(n5230) );
  XOR U7172 ( .A(n7938), .B(n7939), .Z(n6992) );
  XOR U7173 ( .A(n4907), .B(n7940), .Z(n7939) );
  XNOR U7174 ( .A(n7941), .B(n7942), .Z(n4907) );
  AND U7175 ( .A(n7943), .B(n7944), .Z(n7941) );
  XOR U7176 ( .A(n2661), .B(n7945), .Z(n7938) );
  XOR U7177 ( .A(n3538), .B(n5744), .Z(n7945) );
  XOR U7178 ( .A(n7946), .B(n7947), .Z(n5744) );
  ANDN U7179 ( .B(n7948), .A(n7949), .Z(n7946) );
  XNOR U7180 ( .A(n7950), .B(n7951), .Z(n3538) );
  ANDN U7181 ( .B(n7952), .A(n7953), .Z(n7950) );
  XOR U7182 ( .A(n7954), .B(n7955), .Z(n2661) );
  XNOR U7183 ( .A(n2431), .B(n7958), .Z(n1104) );
  IV U7184 ( .A(n5043), .Z(n2431) );
  XOR U7185 ( .A(n6313), .B(n7959), .Z(n5043) );
  XOR U7186 ( .A(n7960), .B(n7961), .Z(n6313) );
  XNOR U7187 ( .A(n3245), .B(n4331), .Z(n7961) );
  XOR U7188 ( .A(n7962), .B(n7963), .Z(n4331) );
  NOR U7189 ( .A(n7964), .B(n7965), .Z(n7962) );
  XOR U7190 ( .A(n7966), .B(n7967), .Z(n3245) );
  ANDN U7191 ( .B(n7968), .A(n7969), .Z(n7966) );
  XOR U7192 ( .A(n5574), .B(n7970), .Z(n7960) );
  XNOR U7193 ( .A(n7971), .B(n2468), .Z(n7970) );
  XOR U7194 ( .A(n7972), .B(n7973), .Z(n2468) );
  AND U7195 ( .A(n7974), .B(n7975), .Z(n7972) );
  XOR U7196 ( .A(n7976), .B(n7977), .Z(n5574) );
  ANDN U7197 ( .B(n7978), .A(n7979), .Z(n7976) );
  XOR U7198 ( .A(n7980), .B(n4122), .Z(out[104]) );
  IV U7199 ( .A(n4296), .Z(n4122) );
  XOR U7200 ( .A(n7009), .B(n2564), .Z(n4296) );
  XNOR U7201 ( .A(n7808), .B(n7981), .Z(n2564) );
  XOR U7202 ( .A(n7982), .B(n7983), .Z(n7808) );
  XOR U7203 ( .A(n4301), .B(n2190), .Z(n7983) );
  XOR U7204 ( .A(n7984), .B(n7884), .Z(n2190) );
  ANDN U7205 ( .B(n7985), .A(n7986), .Z(n7984) );
  XNOR U7206 ( .A(n7987), .B(n7876), .Z(n4301) );
  XOR U7207 ( .A(n6033), .B(n7988), .Z(n7982) );
  XOR U7208 ( .A(n5552), .B(n3743), .Z(n7988) );
  XOR U7209 ( .A(n7989), .B(n7879), .Z(n3743) );
  ANDN U7210 ( .B(n6999), .A(n7007), .Z(n7989) );
  IV U7211 ( .A(n7990), .Z(n6999) );
  XOR U7212 ( .A(n7991), .B(n7992), .Z(n5552) );
  XNOR U7213 ( .A(n7993), .B(n7886), .Z(n6033) );
  AND U7214 ( .A(n6998), .B(n6996), .Z(n7993) );
  XOR U7215 ( .A(n7994), .B(n7985), .Z(n7009) );
  ANDN U7216 ( .B(n7986), .A(n7882), .Z(n7994) );
  AND U7217 ( .A(n3496), .B(n3498), .Z(n7980) );
  XOR U7218 ( .A(n2338), .B(n7995), .Z(n3498) );
  IV U7219 ( .A(n4984), .Z(n2338) );
  XOR U7220 ( .A(n6247), .B(n7996), .Z(n4984) );
  XOR U7221 ( .A(n7997), .B(n7998), .Z(n6247) );
  XOR U7222 ( .A(n3194), .B(n6452), .Z(n7998) );
  XOR U7223 ( .A(n7999), .B(n8000), .Z(n6452) );
  ANDN U7224 ( .B(n8001), .A(n8002), .Z(n7999) );
  XNOR U7225 ( .A(n8003), .B(n8004), .Z(n3194) );
  ANDN U7226 ( .B(n8005), .A(n8006), .Z(n8003) );
  XOR U7227 ( .A(n5509), .B(n8007), .Z(n7997) );
  XOR U7228 ( .A(n8008), .B(n2373), .Z(n8007) );
  XNOR U7229 ( .A(n8009), .B(n8010), .Z(n2373) );
  NOR U7230 ( .A(n8011), .B(n8012), .Z(n8009) );
  XNOR U7231 ( .A(n8013), .B(n8014), .Z(n5509) );
  NOR U7232 ( .A(n8015), .B(n8016), .Z(n8013) );
  XOR U7233 ( .A(n8017), .B(n2404), .Z(n3496) );
  XOR U7234 ( .A(n8018), .B(n6005), .Z(out[1049]) );
  XOR U7235 ( .A(n8019), .B(n2358), .Z(n6005) );
  XNOR U7236 ( .A(n8020), .B(n6146), .Z(n2358) );
  XNOR U7237 ( .A(n8021), .B(n8022), .Z(n6146) );
  XNOR U7238 ( .A(n5397), .B(n3785), .Z(n8022) );
  XOR U7239 ( .A(n8023), .B(n8024), .Z(n3785) );
  XNOR U7240 ( .A(n8027), .B(n8028), .Z(n5397) );
  ANDN U7241 ( .B(n8029), .A(n8030), .Z(n8027) );
  XNOR U7242 ( .A(n6241), .B(n8031), .Z(n8021) );
  XOR U7243 ( .A(n2225), .B(n4753), .Z(n8031) );
  XNOR U7244 ( .A(n8032), .B(n8033), .Z(n4753) );
  ANDN U7245 ( .B(n8034), .A(n8035), .Z(n8032) );
  XOR U7246 ( .A(n8036), .B(n8037), .Z(n2225) );
  ANDN U7247 ( .B(n8038), .A(n8039), .Z(n8036) );
  XOR U7248 ( .A(n8040), .B(n8041), .Z(n6241) );
  AND U7249 ( .A(n8042), .B(n8043), .Z(n8040) );
  ANDN U7250 ( .B(n1108), .A(n1109), .Z(n8018) );
  XNOR U7251 ( .A(n1860), .B(n8044), .Z(n1109) );
  XNOR U7252 ( .A(n8045), .B(n8046), .Z(n1860) );
  XNOR U7253 ( .A(n2440), .B(n8047), .Z(n1108) );
  IV U7254 ( .A(n5048), .Z(n2440) );
  XOR U7255 ( .A(n6317), .B(n8048), .Z(n5048) );
  XOR U7256 ( .A(n8049), .B(n8050), .Z(n6317) );
  XOR U7257 ( .A(n3248), .B(n4385), .Z(n8050) );
  XOR U7258 ( .A(n8051), .B(n8052), .Z(n4385) );
  NOR U7259 ( .A(n8053), .B(n8054), .Z(n8051) );
  XOR U7260 ( .A(n8055), .B(n8056), .Z(n3248) );
  ANDN U7261 ( .B(n8057), .A(n8058), .Z(n8055) );
  XOR U7262 ( .A(n5578), .B(n8059), .Z(n8049) );
  XOR U7263 ( .A(n8060), .B(n2479), .Z(n8059) );
  XNOR U7264 ( .A(n8061), .B(n8062), .Z(n2479) );
  AND U7265 ( .A(n8063), .B(n8064), .Z(n8061) );
  XNOR U7266 ( .A(n8065), .B(n8066), .Z(n5578) );
  ANDN U7267 ( .B(n8067), .A(n8068), .Z(n8065) );
  XOR U7268 ( .A(n8069), .B(n6010), .Z(out[1048]) );
  XOR U7269 ( .A(n8070), .B(n2365), .Z(n6010) );
  XNOR U7270 ( .A(n8071), .B(n6151), .Z(n2365) );
  XNOR U7271 ( .A(n8072), .B(n8073), .Z(n6151) );
  XNOR U7272 ( .A(n5402), .B(n3789), .Z(n8073) );
  XOR U7273 ( .A(n8074), .B(n8075), .Z(n3789) );
  AND U7274 ( .A(n8076), .B(n8077), .Z(n8074) );
  XNOR U7275 ( .A(n8078), .B(n8079), .Z(n5402) );
  ANDN U7276 ( .B(n8080), .A(n8081), .Z(n8078) );
  XNOR U7277 ( .A(n6246), .B(n8082), .Z(n8072) );
  XOR U7278 ( .A(n2232), .B(n4777), .Z(n8082) );
  XNOR U7279 ( .A(n8083), .B(n8084), .Z(n4777) );
  ANDN U7280 ( .B(n8085), .A(n8086), .Z(n8083) );
  XNOR U7281 ( .A(n8087), .B(n8088), .Z(n2232) );
  ANDN U7282 ( .B(n8089), .A(n8090), .Z(n8087) );
  XNOR U7283 ( .A(n8091), .B(n8092), .Z(n6246) );
  ANDN U7284 ( .B(n8093), .A(n8094), .Z(n8091) );
  ANDN U7285 ( .B(n1112), .A(n1114), .Z(n8069) );
  XNOR U7286 ( .A(n1868), .B(n8095), .Z(n1114) );
  IV U7287 ( .A(n5236), .Z(n1868) );
  XOR U7288 ( .A(n7022), .B(n8096), .Z(n5236) );
  XOR U7289 ( .A(n8097), .B(n8098), .Z(n7022) );
  XNOR U7290 ( .A(n4913), .B(n8099), .Z(n8098) );
  XNOR U7291 ( .A(n8100), .B(n7065), .Z(n4913) );
  AND U7292 ( .A(n8101), .B(n8102), .Z(n8100) );
  XOR U7293 ( .A(n2675), .B(n8103), .Z(n8097) );
  XOR U7294 ( .A(n3544), .B(n5807), .Z(n8103) );
  XOR U7295 ( .A(n8104), .B(n7054), .Z(n5807) );
  NOR U7296 ( .A(n8105), .B(n8106), .Z(n8104) );
  XNOR U7297 ( .A(n8107), .B(n8108), .Z(n3544) );
  ANDN U7298 ( .B(n8109), .A(n8110), .Z(n8107) );
  XOR U7299 ( .A(n8111), .B(n7050), .Z(n2675) );
  XNOR U7300 ( .A(n2447), .B(n8114), .Z(n1112) );
  IV U7301 ( .A(n5053), .Z(n2447) );
  XOR U7302 ( .A(n6325), .B(n8115), .Z(n5053) );
  XOR U7303 ( .A(n8116), .B(n8117), .Z(n6325) );
  XNOR U7304 ( .A(n3251), .B(n4429), .Z(n8117) );
  XOR U7305 ( .A(n8118), .B(n8119), .Z(n4429) );
  NOR U7306 ( .A(n8120), .B(n8121), .Z(n8118) );
  XOR U7307 ( .A(n8122), .B(n8123), .Z(n3251) );
  ANDN U7308 ( .B(n8124), .A(n8125), .Z(n8122) );
  XOR U7309 ( .A(n5581), .B(n8126), .Z(n8116) );
  XOR U7310 ( .A(n8127), .B(n2486), .Z(n8126) );
  XNOR U7311 ( .A(n8128), .B(n8129), .Z(n2486) );
  AND U7312 ( .A(n8130), .B(n8131), .Z(n8128) );
  XNOR U7313 ( .A(n8132), .B(n8133), .Z(n5581) );
  ANDN U7314 ( .B(n8134), .A(n8135), .Z(n8132) );
  XOR U7315 ( .A(n8136), .B(n6015), .Z(out[1047]) );
  XOR U7316 ( .A(n8008), .B(n2374), .Z(n6015) );
  XNOR U7317 ( .A(n8137), .B(n8138), .Z(n2374) );
  XNOR U7318 ( .A(n8139), .B(n8140), .Z(n8008) );
  ANDN U7319 ( .B(n8141), .A(n8142), .Z(n8139) );
  ANDN U7320 ( .B(n1116), .A(n1117), .Z(n8136) );
  XNOR U7321 ( .A(n1872), .B(n8143), .Z(n1117) );
  XNOR U7322 ( .A(n6168), .B(n7045), .Z(n1872) );
  XOR U7323 ( .A(n8144), .B(n8145), .Z(n7045) );
  XNOR U7324 ( .A(n4916), .B(n8146), .Z(n8145) );
  XNOR U7325 ( .A(n8147), .B(n7088), .Z(n4916) );
  ANDN U7326 ( .B(n8148), .A(n8149), .Z(n8147) );
  XOR U7327 ( .A(n2682), .B(n8150), .Z(n8144) );
  XOR U7328 ( .A(n3547), .B(n5834), .Z(n8150) );
  XOR U7329 ( .A(n8151), .B(n7077), .Z(n5834) );
  NOR U7330 ( .A(n8152), .B(n8153), .Z(n8151) );
  XNOR U7331 ( .A(n8154), .B(n8155), .Z(n3547) );
  AND U7332 ( .A(n8156), .B(n8157), .Z(n8154) );
  XOR U7333 ( .A(n8158), .B(n7073), .Z(n2682) );
  ANDN U7334 ( .B(n8159), .A(n8160), .Z(n8158) );
  XOR U7335 ( .A(n8161), .B(n8162), .Z(n6168) );
  XOR U7336 ( .A(n4318), .B(n2209), .Z(n8162) );
  XOR U7337 ( .A(n8163), .B(n8164), .Z(n2209) );
  ANDN U7338 ( .B(n7108), .A(n7109), .Z(n8163) );
  XOR U7339 ( .A(n8165), .B(n8166), .Z(n4318) );
  ANDN U7340 ( .B(n7112), .A(n7113), .Z(n8165) );
  XOR U7341 ( .A(n6065), .B(n8167), .Z(n8161) );
  XOR U7342 ( .A(n5576), .B(n3763), .Z(n8167) );
  XOR U7343 ( .A(n8168), .B(n8169), .Z(n3763) );
  ANDN U7344 ( .B(n7099), .A(n7101), .Z(n8168) );
  XNOR U7345 ( .A(n8170), .B(n8171), .Z(n5576) );
  ANDN U7346 ( .B(n7104), .A(n7106), .Z(n8170) );
  XNOR U7347 ( .A(n8172), .B(n8173), .Z(n6065) );
  ANDN U7348 ( .B(n7095), .A(n7097), .Z(n8172) );
  XNOR U7349 ( .A(n2452), .B(n8174), .Z(n1116) );
  IV U7350 ( .A(n5058), .Z(n2452) );
  XOR U7351 ( .A(n6329), .B(n8175), .Z(n5058) );
  XOR U7352 ( .A(n8176), .B(n8177), .Z(n6329) );
  XNOR U7353 ( .A(n3254), .B(n4473), .Z(n8177) );
  XOR U7354 ( .A(n8178), .B(n8179), .Z(n4473) );
  NOR U7355 ( .A(n8180), .B(n8181), .Z(n8178) );
  XOR U7356 ( .A(n8182), .B(n8183), .Z(n3254) );
  ANDN U7357 ( .B(n8184), .A(n8185), .Z(n8182) );
  XOR U7358 ( .A(n5587), .B(n8186), .Z(n8176) );
  XOR U7359 ( .A(n8187), .B(n2491), .Z(n8186) );
  XNOR U7360 ( .A(n8188), .B(n8189), .Z(n2491) );
  AND U7361 ( .A(n8190), .B(n8191), .Z(n8188) );
  XNOR U7362 ( .A(n8192), .B(n8193), .Z(n5587) );
  ANDN U7363 ( .B(n8194), .A(n8195), .Z(n8192) );
  XOR U7364 ( .A(n8196), .B(n6020), .Z(out[1046]) );
  XOR U7365 ( .A(n8197), .B(n2379), .Z(n6020) );
  XNOR U7366 ( .A(n8198), .B(n8199), .Z(n2379) );
  ANDN U7367 ( .B(n1120), .A(n1122), .Z(n8196) );
  XNOR U7368 ( .A(n1876), .B(n8200), .Z(n1122) );
  IV U7369 ( .A(n5246), .Z(n1876) );
  XOR U7370 ( .A(n6173), .B(n7068), .Z(n5246) );
  XOR U7371 ( .A(n8201), .B(n8202), .Z(n7068) );
  XNOR U7372 ( .A(n4920), .B(n8203), .Z(n8202) );
  XNOR U7373 ( .A(n8204), .B(n7114), .Z(n4920) );
  ANDN U7374 ( .B(n8166), .A(n8205), .Z(n8204) );
  XOR U7375 ( .A(n2689), .B(n8206), .Z(n8201) );
  XOR U7376 ( .A(n3549), .B(n5865), .Z(n8206) );
  XOR U7377 ( .A(n8207), .B(n7100), .Z(n5865) );
  ANDN U7378 ( .B(n8169), .A(n8208), .Z(n8207) );
  IV U7379 ( .A(n8209), .Z(n8169) );
  XNOR U7380 ( .A(n8210), .B(n7110), .Z(n3549) );
  ANDN U7381 ( .B(n8211), .A(n8164), .Z(n8210) );
  XOR U7382 ( .A(n8212), .B(n7096), .Z(n2689) );
  XOR U7383 ( .A(n8214), .B(n8215), .Z(n6173) );
  XOR U7384 ( .A(n4323), .B(n2212), .Z(n8215) );
  XOR U7385 ( .A(n8216), .B(n8217), .Z(n2212) );
  ANDN U7386 ( .B(n7165), .A(n7166), .Z(n8216) );
  XOR U7387 ( .A(n8218), .B(n8219), .Z(n4323) );
  ANDN U7388 ( .B(n8220), .A(n7169), .Z(n8218) );
  XOR U7389 ( .A(n6070), .B(n8221), .Z(n8214) );
  XOR U7390 ( .A(n5580), .B(n3767), .Z(n8221) );
  XNOR U7391 ( .A(n8222), .B(n8223), .Z(n3767) );
  ANDN U7392 ( .B(n7156), .A(n7157), .Z(n8222) );
  XNOR U7393 ( .A(n8224), .B(n8225), .Z(n5580) );
  ANDN U7394 ( .B(n7161), .A(n7162), .Z(n8224) );
  XOR U7395 ( .A(n8226), .B(n8227), .Z(n6070) );
  ANDN U7396 ( .B(n7152), .A(n7153), .Z(n8226) );
  XNOR U7397 ( .A(n2459), .B(n8228), .Z(n1120) );
  IV U7398 ( .A(n5063), .Z(n2459) );
  XOR U7399 ( .A(n6333), .B(n8229), .Z(n5063) );
  XOR U7400 ( .A(n8230), .B(n8231), .Z(n6333) );
  XNOR U7401 ( .A(n3257), .B(n4524), .Z(n8231) );
  XOR U7402 ( .A(n8232), .B(n8233), .Z(n4524) );
  NOR U7403 ( .A(n8234), .B(n8235), .Z(n8232) );
  XOR U7404 ( .A(n8236), .B(n8237), .Z(n3257) );
  ANDN U7405 ( .B(n8238), .A(n8239), .Z(n8236) );
  XOR U7406 ( .A(n5592), .B(n8240), .Z(n8230) );
  XOR U7407 ( .A(n8241), .B(n2498), .Z(n8240) );
  XNOR U7408 ( .A(n8242), .B(n8243), .Z(n2498) );
  AND U7409 ( .A(n8244), .B(n8245), .Z(n8242) );
  XOR U7410 ( .A(n8246), .B(n8247), .Z(n5592) );
  XOR U7411 ( .A(n8250), .B(n6025), .Z(out[1045]) );
  XOR U7412 ( .A(n8251), .B(n2386), .Z(n6025) );
  XNOR U7413 ( .A(n8252), .B(n8253), .Z(n2386) );
  ANDN U7414 ( .B(n1124), .A(n1126), .Z(n8250) );
  XNOR U7415 ( .A(n3642), .B(n8254), .Z(n1126) );
  IV U7416 ( .A(n1880), .Z(n3642) );
  XOR U7417 ( .A(n7091), .B(n6177), .Z(n1880) );
  XOR U7418 ( .A(n8255), .B(n8256), .Z(n6177) );
  XOR U7419 ( .A(n4330), .B(n2215), .Z(n8256) );
  XOR U7420 ( .A(n8257), .B(n8258), .Z(n2215) );
  ANDN U7421 ( .B(n7218), .A(n7219), .Z(n8257) );
  XOR U7422 ( .A(n8259), .B(n8260), .Z(n4330) );
  NOR U7423 ( .A(n7223), .B(n7222), .Z(n8259) );
  XOR U7424 ( .A(n6075), .B(n8261), .Z(n8255) );
  XOR U7425 ( .A(n5584), .B(n3774), .Z(n8261) );
  XOR U7426 ( .A(n8262), .B(n8263), .Z(n3774) );
  XOR U7427 ( .A(n8264), .B(n8265), .Z(n5584) );
  NOR U7428 ( .A(n7215), .B(n7214), .Z(n8264) );
  XOR U7429 ( .A(n8266), .B(n8267), .Z(n6075) );
  ANDN U7430 ( .B(n7205), .A(n7206), .Z(n8266) );
  XOR U7431 ( .A(n8268), .B(n8269), .Z(n7091) );
  XNOR U7432 ( .A(n4924), .B(n8270), .Z(n8269) );
  XOR U7433 ( .A(n8271), .B(n7171), .Z(n4924) );
  AND U7434 ( .A(n8219), .B(n8272), .Z(n8271) );
  XNOR U7435 ( .A(n2220), .B(n8273), .Z(n8268) );
  XNOR U7436 ( .A(n3552), .B(n5900), .Z(n8273) );
  XOR U7437 ( .A(n8274), .B(n7158), .Z(n5900) );
  ANDN U7438 ( .B(n8275), .A(n8223), .Z(n8274) );
  XNOR U7439 ( .A(n8276), .B(n7167), .Z(n3552) );
  ANDN U7440 ( .B(n8277), .A(n8217), .Z(n8276) );
  XOR U7441 ( .A(n8278), .B(n7154), .Z(n2220) );
  AND U7442 ( .A(n8227), .B(n8279), .Z(n8278) );
  XNOR U7443 ( .A(n2466), .B(n8280), .Z(n1124) );
  IV U7444 ( .A(n5068), .Z(n2466) );
  XOR U7445 ( .A(n6337), .B(n8281), .Z(n5068) );
  XOR U7446 ( .A(n8282), .B(n8283), .Z(n6337) );
  XNOR U7447 ( .A(n3260), .B(n4575), .Z(n8283) );
  XOR U7448 ( .A(n8284), .B(n8285), .Z(n4575) );
  ANDN U7449 ( .B(n8286), .A(n8287), .Z(n8284) );
  XOR U7450 ( .A(n8288), .B(n8289), .Z(n3260) );
  ANDN U7451 ( .B(n8290), .A(n8291), .Z(n8288) );
  XOR U7452 ( .A(n5597), .B(n8292), .Z(n8282) );
  XOR U7453 ( .A(n8293), .B(n2507), .Z(n8292) );
  XNOR U7454 ( .A(n8294), .B(n8295), .Z(n2507) );
  AND U7455 ( .A(n8296), .B(n8297), .Z(n8294) );
  XNOR U7456 ( .A(n8298), .B(n8299), .Z(n5597) );
  ANDN U7457 ( .B(n8300), .A(n8301), .Z(n8298) );
  XOR U7458 ( .A(n8302), .B(n6030), .Z(out[1044]) );
  XOR U7459 ( .A(n8303), .B(n2395), .Z(n6030) );
  XNOR U7460 ( .A(n8304), .B(n8305), .Z(n2395) );
  ANDN U7461 ( .B(n1128), .A(n1130), .Z(n8302) );
  XNOR U7462 ( .A(n1885), .B(n8306), .Z(n1130) );
  IV U7463 ( .A(n5251), .Z(n1885) );
  XOR U7464 ( .A(n7148), .B(n6182), .Z(n5251) );
  XOR U7465 ( .A(n8307), .B(n8308), .Z(n6182) );
  XOR U7466 ( .A(n4384), .B(n1975), .Z(n8308) );
  XOR U7467 ( .A(n8309), .B(n8310), .Z(n1975) );
  AND U7468 ( .A(n7244), .B(n7242), .Z(n8309) );
  XOR U7469 ( .A(n8311), .B(n8312), .Z(n4384) );
  NOR U7470 ( .A(n7250), .B(n7251), .Z(n8311) );
  XOR U7471 ( .A(n6081), .B(n8313), .Z(n8307) );
  XOR U7472 ( .A(n5589), .B(n3778), .Z(n8313) );
  XOR U7473 ( .A(n8314), .B(n8315), .Z(n3778) );
  XOR U7474 ( .A(n8316), .B(n8317), .Z(n5589) );
  NOR U7475 ( .A(n7246), .B(n7247), .Z(n8316) );
  XOR U7476 ( .A(n8318), .B(n8319), .Z(n6081) );
  ANDN U7477 ( .B(n7233), .A(n7234), .Z(n8318) );
  XOR U7478 ( .A(n8320), .B(n8321), .Z(n7148) );
  XNOR U7479 ( .A(n4929), .B(n8322), .Z(n8321) );
  XOR U7480 ( .A(n8323), .B(n7224), .Z(n4929) );
  AND U7481 ( .A(n8260), .B(n8324), .Z(n8323) );
  XNOR U7482 ( .A(n2227), .B(n8325), .Z(n8320) );
  XOR U7483 ( .A(n3554), .B(n5933), .Z(n8325) );
  XNOR U7484 ( .A(n8326), .B(n7210), .Z(n5933) );
  AND U7485 ( .A(n8263), .B(n8327), .Z(n8326) );
  XOR U7486 ( .A(n8328), .B(n7220), .Z(n3554) );
  ANDN U7487 ( .B(n8329), .A(n8258), .Z(n8328) );
  XOR U7488 ( .A(n8330), .B(n7207), .Z(n2227) );
  AND U7489 ( .A(n8267), .B(n8331), .Z(n8330) );
  XNOR U7490 ( .A(n2477), .B(n8332), .Z(n1128) );
  IV U7491 ( .A(n5073), .Z(n2477) );
  XOR U7492 ( .A(n6341), .B(n8333), .Z(n5073) );
  XOR U7493 ( .A(n8334), .B(n8335), .Z(n6341) );
  XNOR U7494 ( .A(n3263), .B(n4626), .Z(n8335) );
  XOR U7495 ( .A(n8336), .B(n8337), .Z(n4626) );
  NOR U7496 ( .A(n8338), .B(n8339), .Z(n8336) );
  XOR U7497 ( .A(n8340), .B(n8341), .Z(n3263) );
  ANDN U7498 ( .B(n8342), .A(n8343), .Z(n8340) );
  XOR U7499 ( .A(n5601), .B(n8344), .Z(n8334) );
  XOR U7500 ( .A(n8345), .B(n2514), .Z(n8344) );
  XNOR U7501 ( .A(n8346), .B(n8347), .Z(n2514) );
  AND U7502 ( .A(n8348), .B(n8349), .Z(n8346) );
  XOR U7503 ( .A(n8350), .B(n8351), .Z(n5601) );
  XOR U7504 ( .A(n8354), .B(n6036), .Z(out[1043]) );
  XOR U7505 ( .A(n8355), .B(n2404), .Z(n6036) );
  XNOR U7506 ( .A(n8356), .B(n8357), .Z(n2404) );
  ANDN U7507 ( .B(n1136), .A(n1137), .Z(n8354) );
  XNOR U7508 ( .A(n1889), .B(n8358), .Z(n1137) );
  IV U7509 ( .A(n5254), .Z(n1889) );
  XOR U7510 ( .A(n7201), .B(n6187), .Z(n5254) );
  XOR U7511 ( .A(n8359), .B(n8360), .Z(n6187) );
  XNOR U7512 ( .A(n4428), .B(n1978), .Z(n8360) );
  XOR U7513 ( .A(n8361), .B(n8362), .Z(n1978) );
  XOR U7514 ( .A(n8363), .B(n8364), .Z(n4428) );
  XOR U7515 ( .A(n6087), .B(n8365), .Z(n8359) );
  XOR U7516 ( .A(n5594), .B(n3782), .Z(n8365) );
  XOR U7517 ( .A(n8366), .B(n8367), .Z(n3782) );
  ANDN U7518 ( .B(n7307), .A(n7305), .Z(n8366) );
  XNOR U7519 ( .A(n8368), .B(n8369), .Z(n5594) );
  ANDN U7520 ( .B(n7315), .A(n7314), .Z(n8368) );
  XOR U7521 ( .A(n8370), .B(n8371), .Z(n6087) );
  AND U7522 ( .A(n7303), .B(n7301), .Z(n8370) );
  XOR U7523 ( .A(n8372), .B(n8373), .Z(n7201) );
  XNOR U7524 ( .A(n4933), .B(n8374), .Z(n8373) );
  XOR U7525 ( .A(n8375), .B(n7252), .Z(n4933) );
  ANDN U7526 ( .B(n8312), .A(n8376), .Z(n8375) );
  XNOR U7527 ( .A(n2234), .B(n8377), .Z(n8372) );
  XOR U7528 ( .A(n3557), .B(n5988), .Z(n8377) );
  XNOR U7529 ( .A(n8378), .B(n7238), .Z(n5988) );
  ANDN U7530 ( .B(n8315), .A(n8379), .Z(n8378) );
  XNOR U7531 ( .A(n8380), .B(n7243), .Z(n3557) );
  ANDN U7532 ( .B(n8381), .A(n8310), .Z(n8380) );
  XOR U7533 ( .A(n8382), .B(n7235), .Z(n2234) );
  AND U7534 ( .A(n8319), .B(n8383), .Z(n8382) );
  XNOR U7535 ( .A(n2484), .B(n8384), .Z(n1136) );
  IV U7536 ( .A(n5082), .Z(n2484) );
  XOR U7537 ( .A(n6345), .B(n8385), .Z(n5082) );
  XOR U7538 ( .A(n8386), .B(n8387), .Z(n6345) );
  XOR U7539 ( .A(n3266), .B(n4676), .Z(n8387) );
  XOR U7540 ( .A(n8388), .B(n8389), .Z(n4676) );
  NOR U7541 ( .A(n8390), .B(n8391), .Z(n8388) );
  XOR U7542 ( .A(n8392), .B(n8393), .Z(n3266) );
  AND U7543 ( .A(n8394), .B(n8395), .Z(n8392) );
  XOR U7544 ( .A(n5606), .B(n8396), .Z(n8386) );
  XOR U7545 ( .A(n8397), .B(n2521), .Z(n8396) );
  XNOR U7546 ( .A(n8398), .B(n8399), .Z(n2521) );
  ANDN U7547 ( .B(n8400), .A(n8401), .Z(n8398) );
  XOR U7548 ( .A(n8402), .B(n8403), .Z(n5606) );
  NOR U7549 ( .A(n8404), .B(n8405), .Z(n8402) );
  XOR U7550 ( .A(n8406), .B(n6041), .Z(out[1042]) );
  XOR U7551 ( .A(n7410), .B(n2413), .Z(n6041) );
  XNOR U7552 ( .A(n8407), .B(n8408), .Z(n7410) );
  ANDN U7553 ( .B(n8409), .A(n8410), .Z(n8407) );
  ANDN U7554 ( .B(n1140), .A(n1141), .Z(n8406) );
  XNOR U7555 ( .A(n1893), .B(n8411), .Z(n1141) );
  IV U7556 ( .A(n5257), .Z(n1893) );
  XOR U7557 ( .A(n7229), .B(n6192), .Z(n5257) );
  XOR U7558 ( .A(n8412), .B(n8413), .Z(n6192) );
  XNOR U7559 ( .A(n4472), .B(n1981), .Z(n8413) );
  XOR U7560 ( .A(n8414), .B(n8415), .Z(n1981) );
  XOR U7561 ( .A(n8416), .B(n8417), .Z(n4472) );
  NOR U7562 ( .A(n7371), .B(n7372), .Z(n8416) );
  XOR U7563 ( .A(n6092), .B(n8418), .Z(n8412) );
  XOR U7564 ( .A(n5599), .B(n3786), .Z(n8418) );
  XOR U7565 ( .A(n8419), .B(n8420), .Z(n3786) );
  ANDN U7566 ( .B(n7360), .A(n7358), .Z(n8419) );
  XOR U7567 ( .A(n8421), .B(n8422), .Z(n5599) );
  ANDN U7568 ( .B(n7369), .A(n7367), .Z(n8421) );
  XOR U7569 ( .A(n8423), .B(n8424), .Z(n6092) );
  AND U7570 ( .A(n7356), .B(n7354), .Z(n8423) );
  XOR U7571 ( .A(n8425), .B(n8426), .Z(n7229) );
  XOR U7572 ( .A(n4937), .B(n8427), .Z(n8426) );
  XNOR U7573 ( .A(n8428), .B(n7320), .Z(n4937) );
  ANDN U7574 ( .B(n8364), .A(n8429), .Z(n8428) );
  XOR U7575 ( .A(n2241), .B(n8430), .Z(n8425) );
  XOR U7576 ( .A(n3564), .B(n6045), .Z(n8430) );
  XOR U7577 ( .A(n8431), .B(n7306), .Z(n6045) );
  ANDN U7578 ( .B(n8367), .A(n8432), .Z(n8431) );
  XNOR U7579 ( .A(n8433), .B(n7312), .Z(n3564) );
  ANDN U7580 ( .B(n8362), .A(n8434), .Z(n8433) );
  XOR U7581 ( .A(n8435), .B(n7302), .Z(n2241) );
  AND U7582 ( .A(n8371), .B(n8436), .Z(n8435) );
  XNOR U7583 ( .A(n2493), .B(n8437), .Z(n1140) );
  IV U7584 ( .A(n5087), .Z(n2493) );
  XOR U7585 ( .A(n6349), .B(n8438), .Z(n5087) );
  XOR U7586 ( .A(n8439), .B(n8440), .Z(n6349) );
  XNOR U7587 ( .A(n3273), .B(n4701), .Z(n8440) );
  XOR U7588 ( .A(n8441), .B(n8442), .Z(n4701) );
  ANDN U7589 ( .B(n8443), .A(n8444), .Z(n8441) );
  XOR U7590 ( .A(n8445), .B(n8446), .Z(n3273) );
  ANDN U7591 ( .B(n8447), .A(n8448), .Z(n8445) );
  XOR U7592 ( .A(n5609), .B(n8449), .Z(n8439) );
  XOR U7593 ( .A(n8450), .B(n2528), .Z(n8449) );
  XNOR U7594 ( .A(n8451), .B(n8452), .Z(n2528) );
  ANDN U7595 ( .B(n8453), .A(n8454), .Z(n8451) );
  XOR U7596 ( .A(n8455), .B(n8456), .Z(n5609) );
  NOR U7597 ( .A(n8457), .B(n8458), .Z(n8455) );
  XOR U7598 ( .A(n8459), .B(n6053), .Z(out[1041]) );
  XOR U7599 ( .A(n7481), .B(n2420), .Z(n6053) );
  XNOR U7600 ( .A(n8460), .B(n8461), .Z(n7481) );
  ANDN U7601 ( .B(n8462), .A(n8463), .Z(n8460) );
  ANDN U7602 ( .B(n1144), .A(n1145), .Z(n8459) );
  XNOR U7603 ( .A(n1897), .B(n8464), .Z(n1145) );
  IV U7604 ( .A(n5260), .Z(n1897) );
  XOR U7605 ( .A(n7297), .B(n6197), .Z(n5260) );
  XOR U7606 ( .A(n8465), .B(n8466), .Z(n6197) );
  XNOR U7607 ( .A(n4523), .B(n1984), .Z(n8466) );
  XNOR U7608 ( .A(n8467), .B(n8468), .Z(n1984) );
  AND U7609 ( .A(n7434), .B(n8469), .Z(n8467) );
  XOR U7610 ( .A(n8470), .B(n8471), .Z(n4523) );
  XOR U7611 ( .A(n6098), .B(n8472), .Z(n8465) );
  XOR U7612 ( .A(n5604), .B(n3790), .Z(n8472) );
  XOR U7613 ( .A(n8473), .B(n8474), .Z(n3790) );
  ANDN U7614 ( .B(n7431), .A(n7429), .Z(n8473) );
  XNOR U7615 ( .A(n8475), .B(n8476), .Z(n5604) );
  ANDN U7616 ( .B(n7440), .A(n7438), .Z(n8475) );
  XOR U7617 ( .A(n8477), .B(n8478), .Z(n6098) );
  ANDN U7618 ( .B(n7425), .A(n7427), .Z(n8477) );
  XOR U7619 ( .A(n8479), .B(n8480), .Z(n7297) );
  XNOR U7620 ( .A(n4941), .B(n8481), .Z(n8480) );
  XNOR U7621 ( .A(n8482), .B(n7373), .Z(n4941) );
  ANDN U7622 ( .B(n8417), .A(n8483), .Z(n8482) );
  XOR U7623 ( .A(n2255), .B(n8484), .Z(n8479) );
  XOR U7624 ( .A(n3566), .B(n6104), .Z(n8484) );
  XOR U7625 ( .A(n8485), .B(n7359), .Z(n6104) );
  ANDN U7626 ( .B(n8420), .A(n8486), .Z(n8485) );
  XNOR U7627 ( .A(n8487), .B(n7365), .Z(n3566) );
  ANDN U7628 ( .B(n8415), .A(n8488), .Z(n8487) );
  XOR U7629 ( .A(n8489), .B(n7355), .Z(n2255) );
  ANDN U7630 ( .B(n8424), .A(n8490), .Z(n8489) );
  XNOR U7631 ( .A(n2500), .B(n8491), .Z(n1144) );
  IV U7632 ( .A(n4821), .Z(n2500) );
  XOR U7633 ( .A(n5923), .B(n6353), .Z(n4821) );
  XOR U7634 ( .A(n8492), .B(n8493), .Z(n6353) );
  XNOR U7635 ( .A(n3277), .B(n4725), .Z(n8493) );
  XOR U7636 ( .A(n8494), .B(n8495), .Z(n4725) );
  NOR U7637 ( .A(n8496), .B(n8497), .Z(n8494) );
  XOR U7638 ( .A(n8498), .B(n8499), .Z(n3277) );
  AND U7639 ( .A(n8500), .B(n8501), .Z(n8498) );
  XOR U7640 ( .A(n5613), .B(n8502), .Z(n8492) );
  XOR U7641 ( .A(n8503), .B(n2535), .Z(n8502) );
  XOR U7642 ( .A(n8504), .B(n8505), .Z(n2535) );
  ANDN U7643 ( .B(n8506), .A(n8507), .Z(n8504) );
  XOR U7644 ( .A(n8508), .B(n8509), .Z(n5613) );
  NOR U7645 ( .A(n8510), .B(n8511), .Z(n8508) );
  XOR U7646 ( .A(n8512), .B(n8513), .Z(n5923) );
  XNOR U7647 ( .A(n3805), .B(n5153), .Z(n8513) );
  XOR U7648 ( .A(n8514), .B(n8515), .Z(n5153) );
  ANDN U7649 ( .B(n8516), .A(n8517), .Z(n8514) );
  XOR U7650 ( .A(n8518), .B(n8519), .Z(n3805) );
  ANDN U7651 ( .B(n8520), .A(n8521), .Z(n8518) );
  XOR U7652 ( .A(n6412), .B(n8522), .Z(n8512) );
  XOR U7653 ( .A(n1756), .B(n8523), .Z(n8522) );
  XNOR U7654 ( .A(n8524), .B(n8525), .Z(n1756) );
  ANDN U7655 ( .B(n8526), .A(n8527), .Z(n8524) );
  XNOR U7656 ( .A(n8528), .B(n8529), .Z(n6412) );
  ANDN U7657 ( .B(n8530), .A(n8531), .Z(n8528) );
  XOR U7658 ( .A(n8532), .B(n6058), .Z(out[1040]) );
  XOR U7659 ( .A(n7525), .B(n2427), .Z(n6058) );
  XNOR U7660 ( .A(n8533), .B(n8534), .Z(n7525) );
  ANDN U7661 ( .B(n8535), .A(n8536), .Z(n8533) );
  ANDN U7662 ( .B(n1148), .A(n1149), .Z(n8532) );
  XNOR U7663 ( .A(n1901), .B(n8537), .Z(n1149) );
  IV U7664 ( .A(n5263), .Z(n1901) );
  XOR U7665 ( .A(n7350), .B(n6202), .Z(n5263) );
  XOR U7666 ( .A(n8538), .B(n8539), .Z(n6202) );
  XNOR U7667 ( .A(n4574), .B(n1987), .Z(n8539) );
  XOR U7668 ( .A(n8540), .B(n8541), .Z(n1987) );
  AND U7669 ( .A(n7505), .B(n8542), .Z(n8540) );
  XOR U7670 ( .A(n8543), .B(n8544), .Z(n4574) );
  NOR U7671 ( .A(n7513), .B(n7515), .Z(n8543) );
  XOR U7672 ( .A(n6109), .B(n8545), .Z(n8538) );
  XOR U7673 ( .A(n5608), .B(n3794), .Z(n8545) );
  XOR U7674 ( .A(n8546), .B(n8547), .Z(n3794) );
  ANDN U7675 ( .B(n7502), .A(n7500), .Z(n8546) );
  XNOR U7676 ( .A(n8548), .B(n8549), .Z(n5608) );
  ANDN U7677 ( .B(n7511), .A(n7509), .Z(n8548) );
  XOR U7678 ( .A(n8550), .B(n8551), .Z(n6109) );
  AND U7679 ( .A(n7498), .B(n7496), .Z(n8550) );
  XOR U7680 ( .A(n8552), .B(n8553), .Z(n7350) );
  XNOR U7681 ( .A(n4949), .B(n8554), .Z(n8553) );
  XOR U7682 ( .A(n8555), .B(n7443), .Z(n4949) );
  ANDN U7683 ( .B(n8471), .A(n8556), .Z(n8555) );
  XOR U7684 ( .A(n2262), .B(n8557), .Z(n8552) );
  XOR U7685 ( .A(n3568), .B(n6162), .Z(n8557) );
  XOR U7686 ( .A(n8558), .B(n7430), .Z(n6162) );
  ANDN U7687 ( .B(n8474), .A(n8559), .Z(n8558) );
  IV U7688 ( .A(n8560), .Z(n8474) );
  XNOR U7689 ( .A(n8561), .B(n7436), .Z(n3568) );
  NOR U7690 ( .A(n8562), .B(n8468), .Z(n8561) );
  XOR U7691 ( .A(n8563), .B(n7426), .Z(n2262) );
  XNOR U7692 ( .A(n2505), .B(n8565), .Z(n1148) );
  IV U7693 ( .A(n4826), .Z(n2505) );
  XOR U7694 ( .A(n5928), .B(n6357), .Z(n4826) );
  XOR U7695 ( .A(n8566), .B(n8567), .Z(n6357) );
  XOR U7696 ( .A(n3280), .B(n4752), .Z(n8567) );
  XOR U7697 ( .A(n8568), .B(n8569), .Z(n4752) );
  AND U7698 ( .A(n8570), .B(n8519), .Z(n8568) );
  IV U7699 ( .A(n8571), .Z(n8519) );
  XOR U7700 ( .A(n8572), .B(n8573), .Z(n3280) );
  ANDN U7701 ( .B(n8574), .A(n8525), .Z(n8572) );
  XOR U7702 ( .A(n5296), .B(n8575), .Z(n8566) );
  XOR U7703 ( .A(n8576), .B(n2542), .Z(n8575) );
  XOR U7704 ( .A(n8577), .B(n8578), .Z(n2542) );
  NOR U7705 ( .A(n8579), .B(n8580), .Z(n8577) );
  XNOR U7706 ( .A(n8581), .B(n8582), .Z(n5296) );
  NOR U7707 ( .A(n8583), .B(n8529), .Z(n8581) );
  XOR U7708 ( .A(n8584), .B(n8585), .Z(n5928) );
  XNOR U7709 ( .A(n3809), .B(n5155), .Z(n8585) );
  XNOR U7710 ( .A(n8586), .B(n8587), .Z(n5155) );
  ANDN U7711 ( .B(n8588), .A(n6476), .Z(n8586) );
  XNOR U7712 ( .A(n8589), .B(n8590), .Z(n3809) );
  ANDN U7713 ( .B(n8591), .A(n6463), .Z(n8589) );
  XNOR U7714 ( .A(n8592), .B(n8593), .Z(n8584) );
  XOR U7715 ( .A(n4196), .B(n1762), .Z(n8593) );
  XOR U7716 ( .A(n8594), .B(n8595), .Z(n1762) );
  ANDN U7717 ( .B(n8596), .A(n6467), .Z(n8594) );
  XNOR U7718 ( .A(n8597), .B(n8598), .Z(n4196) );
  ANDN U7719 ( .B(n8599), .A(n6480), .Z(n8597) );
  XOR U7720 ( .A(n8600), .B(n4125), .Z(out[103]) );
  IV U7721 ( .A(n4299), .Z(n4125) );
  XOR U7722 ( .A(n8601), .B(n3707), .Z(n4299) );
  XNOR U7723 ( .A(n7870), .B(n8602), .Z(n3707) );
  XOR U7724 ( .A(n8603), .B(n8604), .Z(n7870) );
  XOR U7725 ( .A(n4304), .B(n2193), .Z(n8604) );
  XOR U7726 ( .A(n8605), .B(n7953), .Z(n2193) );
  ANDN U7727 ( .B(n8606), .A(n8607), .Z(n8605) );
  XOR U7728 ( .A(n8608), .B(n7944), .Z(n4304) );
  IV U7729 ( .A(n8609), .Z(n7944) );
  XOR U7730 ( .A(n6038), .B(n8612), .Z(n8603) );
  XOR U7731 ( .A(n5556), .B(n3747), .Z(n8612) );
  XOR U7732 ( .A(n8613), .B(n7948), .Z(n3747) );
  NOR U7733 ( .A(n8614), .B(n8615), .Z(n8613) );
  XNOR U7734 ( .A(n8616), .B(n8617), .Z(n5556) );
  AND U7735 ( .A(n8618), .B(n8619), .Z(n8616) );
  XOR U7736 ( .A(n8620), .B(n7956), .Z(n6038) );
  ANDN U7737 ( .B(n8621), .A(n8622), .Z(n8620) );
  AND U7738 ( .A(n3528), .B(n3530), .Z(n8600) );
  XOR U7739 ( .A(n2345), .B(n8623), .Z(n3530) );
  IV U7740 ( .A(n4988), .Z(n2345) );
  XOR U7741 ( .A(n6252), .B(n8624), .Z(n4988) );
  XOR U7742 ( .A(n8625), .B(n8626), .Z(n6252) );
  XOR U7743 ( .A(n3204), .B(n6678), .Z(n8626) );
  XOR U7744 ( .A(n8627), .B(n8628), .Z(n6678) );
  ANDN U7745 ( .B(n8629), .A(n8630), .Z(n8627) );
  XNOR U7746 ( .A(n8631), .B(n8632), .Z(n3204) );
  ANDN U7747 ( .B(n8633), .A(n8634), .Z(n8631) );
  XOR U7748 ( .A(n5512), .B(n8635), .Z(n8625) );
  XOR U7749 ( .A(n8197), .B(n2378), .Z(n8635) );
  XNOR U7750 ( .A(n8636), .B(n8637), .Z(n2378) );
  ANDN U7751 ( .B(n8638), .A(n8639), .Z(n8636) );
  XNOR U7752 ( .A(n8640), .B(n8641), .Z(n8197) );
  ANDN U7753 ( .B(n8642), .A(n8643), .Z(n8640) );
  XNOR U7754 ( .A(n8644), .B(n8645), .Z(n5512) );
  ANDN U7755 ( .B(n8646), .A(n8647), .Z(n8644) );
  XOR U7756 ( .A(n7404), .B(n2413), .Z(n3528) );
  XNOR U7757 ( .A(n8648), .B(n8649), .Z(n2413) );
  XOR U7758 ( .A(n8650), .B(n8651), .Z(n7404) );
  NOR U7759 ( .A(n8652), .B(n8653), .Z(n8650) );
  XOR U7760 ( .A(n8654), .B(n6063), .Z(out[1039]) );
  XOR U7761 ( .A(n7624), .B(n2434), .Z(n6063) );
  XNOR U7762 ( .A(n8655), .B(n8656), .Z(n7624) );
  ANDN U7763 ( .B(n8657), .A(n8658), .Z(n8655) );
  ANDN U7764 ( .B(n1152), .A(n1153), .Z(n8654) );
  XNOR U7765 ( .A(n1906), .B(n8659), .Z(n1153) );
  IV U7766 ( .A(n5266), .Z(n1906) );
  XOR U7767 ( .A(n7421), .B(n6207), .Z(n5266) );
  XOR U7768 ( .A(n8660), .B(n8661), .Z(n6207) );
  XNOR U7769 ( .A(n4625), .B(n1991), .Z(n8661) );
  XOR U7770 ( .A(n8662), .B(n8663), .Z(n1991) );
  AND U7771 ( .A(n7579), .B(n7577), .Z(n8662) );
  XOR U7772 ( .A(n8664), .B(n8665), .Z(n4625) );
  NOR U7773 ( .A(n7587), .B(n7585), .Z(n8664) );
  IV U7774 ( .A(n8666), .Z(n7587) );
  XOR U7775 ( .A(n6114), .B(n8667), .Z(n8660) );
  XOR U7776 ( .A(n5612), .B(n3798), .Z(n8667) );
  XOR U7777 ( .A(n8668), .B(n8669), .Z(n3798) );
  ANDN U7778 ( .B(n7574), .A(n7572), .Z(n8668) );
  XOR U7779 ( .A(n8670), .B(n8671), .Z(n5612) );
  ANDN U7780 ( .B(n7583), .A(n7581), .Z(n8670) );
  XOR U7781 ( .A(n8672), .B(n8673), .Z(n6114) );
  AND U7782 ( .A(n7570), .B(n7568), .Z(n8672) );
  XOR U7783 ( .A(n8674), .B(n8675), .Z(n7421) );
  XNOR U7784 ( .A(n4952), .B(n8676), .Z(n8675) );
  XOR U7785 ( .A(n8677), .B(n7514), .Z(n4952) );
  ANDN U7786 ( .B(n8544), .A(n8678), .Z(n8677) );
  XOR U7787 ( .A(n2269), .B(n8679), .Z(n8674) );
  XOR U7788 ( .A(n3570), .B(n6217), .Z(n8679) );
  XOR U7789 ( .A(n8680), .B(n7501), .Z(n6217) );
  ANDN U7790 ( .B(n8547), .A(n8681), .Z(n8680) );
  XNOR U7791 ( .A(n8682), .B(n7507), .Z(n3570) );
  XOR U7792 ( .A(n8684), .B(n7497), .Z(n2269) );
  ANDN U7793 ( .B(n8551), .A(n8685), .Z(n8684) );
  XOR U7794 ( .A(n8686), .B(n2513), .Z(n1152) );
  XOR U7795 ( .A(n5939), .B(n6361), .Z(n2513) );
  XOR U7796 ( .A(n8687), .B(n8688), .Z(n6361) );
  XNOR U7797 ( .A(n3283), .B(n4776), .Z(n8688) );
  XOR U7798 ( .A(n8689), .B(n6464), .Z(n4776) );
  AND U7799 ( .A(n8590), .B(n6465), .Z(n8689) );
  XOR U7800 ( .A(n8690), .B(n6468), .Z(n3283) );
  ANDN U7801 ( .B(n6469), .A(n8595), .Z(n8690) );
  XOR U7802 ( .A(n5301), .B(n8691), .Z(n8687) );
  XOR U7803 ( .A(n6458), .B(n2553), .Z(n8691) );
  XOR U7804 ( .A(n8692), .B(n6473), .Z(n2553) );
  ANDN U7805 ( .B(n6474), .A(n8693), .Z(n8692) );
  XOR U7806 ( .A(n8694), .B(n6477), .Z(n6458) );
  AND U7807 ( .A(n8587), .B(n6478), .Z(n8694) );
  XNOR U7808 ( .A(n8695), .B(n6481), .Z(n5301) );
  AND U7809 ( .A(n8598), .B(n6482), .Z(n8695) );
  XOR U7810 ( .A(n8696), .B(n8697), .Z(n5939) );
  XOR U7811 ( .A(n3815), .B(n5158), .Z(n8697) );
  XOR U7812 ( .A(n8698), .B(n8699), .Z(n5158) );
  AND U7813 ( .A(n6502), .B(n8700), .Z(n8698) );
  XNOR U7814 ( .A(n8701), .B(n8702), .Z(n3815) );
  XOR U7815 ( .A(n4199), .B(n8704), .Z(n8696) );
  XOR U7816 ( .A(n1765), .B(n8705), .Z(n8704) );
  XNOR U7817 ( .A(n8706), .B(n8707), .Z(n1765) );
  ANDN U7818 ( .B(n8708), .A(n6493), .Z(n8706) );
  XNOR U7819 ( .A(n8709), .B(n8710), .Z(n4199) );
  XNOR U7820 ( .A(n8712), .B(n6068), .Z(out[1038]) );
  XNOR U7821 ( .A(n2438), .B(n7688), .Z(n6068) );
  XOR U7822 ( .A(n8713), .B(n8714), .Z(n7688) );
  ANDN U7823 ( .B(n8715), .A(n8716), .Z(n8713) );
  XNOR U7824 ( .A(n8717), .B(n8718), .Z(n2438) );
  ANDN U7825 ( .B(n1156), .A(n1157), .Z(n8712) );
  XNOR U7826 ( .A(n1914), .B(n8719), .Z(n1157) );
  IV U7827 ( .A(n5269), .Z(n1914) );
  XOR U7828 ( .A(n7492), .B(n6212), .Z(n5269) );
  XOR U7829 ( .A(n8720), .B(n8721), .Z(n6212) );
  XNOR U7830 ( .A(n4675), .B(n1994), .Z(n8721) );
  XOR U7831 ( .A(n8722), .B(n8723), .Z(n1994) );
  AND U7832 ( .A(n7648), .B(n7650), .Z(n8722) );
  XOR U7833 ( .A(n8724), .B(n8725), .Z(n4675) );
  AND U7834 ( .A(n7656), .B(n8726), .Z(n8724) );
  XOR U7835 ( .A(n6120), .B(n8727), .Z(n8720) );
  XOR U7836 ( .A(n5295), .B(n3803), .Z(n8727) );
  XNOR U7837 ( .A(n8728), .B(n8729), .Z(n3803) );
  ANDN U7838 ( .B(n7645), .A(n7643), .Z(n8728) );
  XNOR U7839 ( .A(n8730), .B(n8731), .Z(n5295) );
  AND U7840 ( .A(n7654), .B(n7652), .Z(n8730) );
  XOR U7841 ( .A(n8732), .B(n8733), .Z(n6120) );
  AND U7842 ( .A(n7639), .B(n8734), .Z(n8732) );
  XOR U7843 ( .A(n8735), .B(n8736), .Z(n7492) );
  XNOR U7844 ( .A(n4955), .B(n8737), .Z(n8736) );
  XOR U7845 ( .A(n8738), .B(n7586), .Z(n4955) );
  ANDN U7846 ( .B(n8665), .A(n8739), .Z(n8738) );
  XOR U7847 ( .A(n2276), .B(n8740), .Z(n8735) );
  XOR U7848 ( .A(n3572), .B(n6274), .Z(n8740) );
  XOR U7849 ( .A(n8741), .B(n7573), .Z(n6274) );
  ANDN U7850 ( .B(n8669), .A(n8742), .Z(n8741) );
  XOR U7851 ( .A(n8743), .B(n7578), .Z(n3572) );
  ANDN U7852 ( .B(n8663), .A(n8744), .Z(n8743) );
  XOR U7853 ( .A(n8745), .B(n7569), .Z(n2276) );
  ANDN U7854 ( .B(n8673), .A(n8746), .Z(n8745) );
  XNOR U7855 ( .A(n2519), .B(n8747), .Z(n1156) );
  IV U7856 ( .A(n4838), .Z(n2519) );
  XOR U7857 ( .A(n5944), .B(n6369), .Z(n4838) );
  XOR U7858 ( .A(n8748), .B(n8749), .Z(n6369) );
  XOR U7859 ( .A(n3287), .B(n4801), .Z(n8749) );
  XOR U7860 ( .A(n8750), .B(n6490), .Z(n4801) );
  ANDN U7861 ( .B(n6491), .A(n8702), .Z(n8750) );
  XNOR U7862 ( .A(n8751), .B(n6494), .Z(n3287) );
  ANDN U7863 ( .B(n6495), .A(n8707), .Z(n8751) );
  XOR U7864 ( .A(n5305), .B(n8752), .Z(n8748) );
  XOR U7865 ( .A(n6484), .B(n2560), .Z(n8752) );
  XNOR U7866 ( .A(n8753), .B(n6499), .Z(n2560) );
  ANDN U7867 ( .B(n6500), .A(n8754), .Z(n8753) );
  XNOR U7868 ( .A(n8755), .B(n6503), .Z(n6484) );
  ANDN U7869 ( .B(n6504), .A(n8699), .Z(n8755) );
  XNOR U7870 ( .A(n8756), .B(n6507), .Z(n5305) );
  ANDN U7871 ( .B(n6508), .A(n8710), .Z(n8756) );
  XOR U7872 ( .A(n8757), .B(n8758), .Z(n5944) );
  XOR U7873 ( .A(n3819), .B(n5161), .Z(n8758) );
  XOR U7874 ( .A(n8759), .B(n8760), .Z(n5161) );
  ANDN U7875 ( .B(n8761), .A(n6528), .Z(n8759) );
  XOR U7876 ( .A(n8762), .B(n8763), .Z(n3819) );
  ANDN U7877 ( .B(n8764), .A(n6515), .Z(n8762) );
  XOR U7878 ( .A(n4207), .B(n8765), .Z(n8757) );
  XOR U7879 ( .A(n1774), .B(n8766), .Z(n8765) );
  XNOR U7880 ( .A(n8767), .B(n8768), .Z(n1774) );
  ANDN U7881 ( .B(n8769), .A(n6519), .Z(n8767) );
  XNOR U7882 ( .A(n8770), .B(n8771), .Z(n4207) );
  ANDN U7883 ( .B(n8772), .A(n6532), .Z(n8770) );
  XOR U7884 ( .A(n8773), .B(n6073), .Z(out[1037]) );
  XOR U7885 ( .A(n2445), .B(n7763), .Z(n6073) );
  XOR U7886 ( .A(n8774), .B(n8775), .Z(n7763) );
  AND U7887 ( .A(n8776), .B(n8777), .Z(n8774) );
  ANDN U7888 ( .B(n6403), .A(n1161), .Z(n8773) );
  XNOR U7889 ( .A(n1919), .B(n8780), .Z(n1161) );
  IV U7890 ( .A(n5272), .Z(n1919) );
  XOR U7891 ( .A(n7564), .B(n6222), .Z(n5272) );
  XOR U7892 ( .A(n8781), .B(n8782), .Z(n6222) );
  XNOR U7893 ( .A(n4700), .B(n1997), .Z(n8782) );
  XOR U7894 ( .A(n8783), .B(n8784), .Z(n1997) );
  AND U7895 ( .A(n7721), .B(n8785), .Z(n8783) );
  XOR U7896 ( .A(n8786), .B(n8787), .Z(n4700) );
  ANDN U7897 ( .B(n7731), .A(n7729), .Z(n8786) );
  XOR U7898 ( .A(n6126), .B(n8788), .Z(n8781) );
  XOR U7899 ( .A(n5299), .B(n3807), .Z(n8788) );
  XOR U7900 ( .A(n8789), .B(n8790), .Z(n3807) );
  ANDN U7901 ( .B(n7718), .A(n7716), .Z(n8789) );
  XNOR U7902 ( .A(n8791), .B(n8792), .Z(n5299) );
  AND U7903 ( .A(n7727), .B(n7725), .Z(n8791) );
  XOR U7904 ( .A(n8793), .B(n8794), .Z(n6126) );
  ANDN U7905 ( .B(n8795), .A(n7712), .Z(n8793) );
  XOR U7906 ( .A(n8796), .B(n8797), .Z(n7564) );
  XNOR U7907 ( .A(n4958), .B(n8798), .Z(n8797) );
  XNOR U7908 ( .A(n8799), .B(n7658), .Z(n4958) );
  ANDN U7909 ( .B(n8725), .A(n8800), .Z(n8799) );
  XOR U7910 ( .A(n2283), .B(n8801), .Z(n8796) );
  XOR U7911 ( .A(n3574), .B(n6321), .Z(n8801) );
  XOR U7912 ( .A(n8802), .B(n7644), .Z(n6321) );
  NOR U7913 ( .A(n8729), .B(n8803), .Z(n8802) );
  XOR U7914 ( .A(n8804), .B(n7649), .Z(n3574) );
  ANDN U7915 ( .B(n8723), .A(n8805), .Z(n8804) );
  XNOR U7916 ( .A(n8806), .B(n7641), .Z(n2283) );
  ANDN U7917 ( .B(n8733), .A(n8807), .Z(n8806) );
  XNOR U7918 ( .A(n2526), .B(n8808), .Z(n6403) );
  XOR U7919 ( .A(n5949), .B(n6374), .Z(n2526) );
  XNOR U7920 ( .A(n8809), .B(n8810), .Z(n6374) );
  XNOR U7921 ( .A(n2567), .B(n5310), .Z(n8810) );
  XOR U7922 ( .A(n8811), .B(n6533), .Z(n5310) );
  ANDN U7923 ( .B(n6534), .A(n8771), .Z(n8811) );
  XOR U7924 ( .A(n8812), .B(n6525), .Z(n2567) );
  ANDN U7925 ( .B(n6526), .A(n8813), .Z(n8812) );
  XNOR U7926 ( .A(n3290), .B(n8814), .Z(n8809) );
  XOR U7927 ( .A(n4831), .B(n6510), .Z(n8814) );
  XOR U7928 ( .A(n8815), .B(n6529), .Z(n6510) );
  ANDN U7929 ( .B(n6530), .A(n8760), .Z(n8815) );
  XOR U7930 ( .A(n8816), .B(n6516), .Z(n4831) );
  AND U7931 ( .A(n8763), .B(n6517), .Z(n8816) );
  XOR U7932 ( .A(n8817), .B(n6520), .Z(n3290) );
  ANDN U7933 ( .B(n6521), .A(n8768), .Z(n8817) );
  XOR U7934 ( .A(n8818), .B(n8819), .Z(n5949) );
  XOR U7935 ( .A(n3823), .B(n5164), .Z(n8819) );
  XOR U7936 ( .A(n8820), .B(n8821), .Z(n5164) );
  ANDN U7937 ( .B(n8822), .A(n6562), .Z(n8820) );
  XNOR U7938 ( .A(n8823), .B(n8824), .Z(n3823) );
  ANDN U7939 ( .B(n8825), .A(n6541), .Z(n8823) );
  XOR U7940 ( .A(n4209), .B(n8826), .Z(n8818) );
  XOR U7941 ( .A(n1779), .B(n8827), .Z(n8826) );
  XNOR U7942 ( .A(n8828), .B(n8829), .Z(n1779) );
  ANDN U7943 ( .B(n8830), .A(n6545), .Z(n8828) );
  XNOR U7944 ( .A(n8831), .B(n8832), .Z(n4209) );
  ANDN U7945 ( .B(n8833), .A(n6566), .Z(n8831) );
  XOR U7946 ( .A(n8834), .B(n6078), .Z(out[1036]) );
  XOR U7947 ( .A(n7834), .B(n2455), .Z(n6078) );
  IV U7948 ( .A(n3239), .Z(n2455) );
  XNOR U7949 ( .A(n8835), .B(n8836), .Z(n3239) );
  XOR U7950 ( .A(n8837), .B(n8838), .Z(n7834) );
  NOR U7951 ( .A(n8839), .B(n8840), .Z(n8837) );
  ANDN U7952 ( .B(n1164), .A(n1165), .Z(n8834) );
  XNOR U7953 ( .A(n1923), .B(n8841), .Z(n1165) );
  IV U7954 ( .A(n5279), .Z(n1923) );
  XOR U7955 ( .A(n7635), .B(n6227), .Z(n5279) );
  XOR U7956 ( .A(n8842), .B(n8843), .Z(n6227) );
  XNOR U7957 ( .A(n4724), .B(n2004), .Z(n8843) );
  XNOR U7958 ( .A(n8844), .B(n8845), .Z(n2004) );
  ANDN U7959 ( .B(n7798), .A(n7796), .Z(n8844) );
  XOR U7960 ( .A(n8846), .B(n8847), .Z(n4724) );
  ANDN U7961 ( .B(n7805), .A(n7804), .Z(n8846) );
  XOR U7962 ( .A(n6132), .B(n8848), .Z(n8842) );
  XOR U7963 ( .A(n5303), .B(n3811), .Z(n8848) );
  XOR U7964 ( .A(n8849), .B(n8850), .Z(n3811) );
  XOR U7965 ( .A(n8851), .B(n8852), .Z(n5303) );
  AND U7966 ( .A(n7800), .B(n7802), .Z(n8851) );
  XOR U7967 ( .A(n8853), .B(n8854), .Z(n6132) );
  AND U7968 ( .A(n7787), .B(n7789), .Z(n8853) );
  IV U7969 ( .A(n8855), .Z(n7787) );
  XOR U7970 ( .A(n8856), .B(n8857), .Z(n7635) );
  XNOR U7971 ( .A(n4961), .B(n8858), .Z(n8857) );
  XOR U7972 ( .A(n8859), .B(n7730), .Z(n4961) );
  ANDN U7973 ( .B(n8787), .A(n8860), .Z(n8859) );
  XOR U7974 ( .A(n2290), .B(n8861), .Z(n8856) );
  XOR U7975 ( .A(n3402), .B(n6365), .Z(n8861) );
  XOR U7976 ( .A(n8862), .B(n7717), .Z(n6365) );
  ANDN U7977 ( .B(n8790), .A(n8863), .Z(n8862) );
  XOR U7978 ( .A(n8864), .B(n7722), .Z(n3402) );
  ANDN U7979 ( .B(n8784), .A(n8865), .Z(n8864) );
  XOR U7980 ( .A(n8866), .B(n7713), .Z(n2290) );
  XNOR U7981 ( .A(n2533), .B(n8868), .Z(n1164) );
  IV U7982 ( .A(n4845), .Z(n2533) );
  XOR U7983 ( .A(n5954), .B(n6377), .Z(n4845) );
  XOR U7984 ( .A(n8869), .B(n8870), .Z(n6377) );
  XNOR U7985 ( .A(n3293), .B(n4870), .Z(n8870) );
  XOR U7986 ( .A(n8871), .B(n6542), .Z(n4870) );
  ANDN U7987 ( .B(n6543), .A(n8824), .Z(n8871) );
  XOR U7988 ( .A(n8872), .B(n6546), .Z(n3293) );
  ANDN U7989 ( .B(n6547), .A(n8829), .Z(n8872) );
  XOR U7990 ( .A(n5319), .B(n8873), .Z(n8869) );
  XOR U7991 ( .A(n6536), .B(n2574), .Z(n8873) );
  XOR U7992 ( .A(n8874), .B(n6559), .Z(n2574) );
  ANDN U7993 ( .B(n6560), .A(n8875), .Z(n8874) );
  XOR U7994 ( .A(n8876), .B(n6563), .Z(n6536) );
  ANDN U7995 ( .B(n6564), .A(n8821), .Z(n8876) );
  XNOR U7996 ( .A(n8877), .B(n6567), .Z(n5319) );
  ANDN U7997 ( .B(n6568), .A(n8832), .Z(n8877) );
  XOR U7998 ( .A(n8878), .B(n8879), .Z(n5954) );
  XOR U7999 ( .A(n3827), .B(n5172), .Z(n8879) );
  XOR U8000 ( .A(n8880), .B(n8881), .Z(n5172) );
  ANDN U8001 ( .B(n8882), .A(n6588), .Z(n8880) );
  XOR U8002 ( .A(n8883), .B(n8884), .Z(n3827) );
  ANDN U8003 ( .B(n8885), .A(n6575), .Z(n8883) );
  XOR U8004 ( .A(n4211), .B(n8886), .Z(n8878) );
  XOR U8005 ( .A(n1783), .B(n8887), .Z(n8886) );
  XNOR U8006 ( .A(n8888), .B(n8889), .Z(n1783) );
  ANDN U8007 ( .B(n8890), .A(n6579), .Z(n8888) );
  XNOR U8008 ( .A(n8891), .B(n8892), .Z(n4211) );
  AND U8009 ( .A(n6592), .B(n8893), .Z(n8891) );
  XOR U8010 ( .A(n8894), .B(n6084), .Z(out[1035]) );
  XNOR U8011 ( .A(n7901), .B(n2462), .Z(n6084) );
  XOR U8012 ( .A(n8897), .B(n8898), .Z(n7901) );
  ANDN U8013 ( .B(n8899), .A(n8900), .Z(n8897) );
  ANDN U8014 ( .B(n1168), .A(n1169), .Z(n8894) );
  XNOR U8015 ( .A(n1927), .B(n8901), .Z(n1169) );
  IV U8016 ( .A(n5282), .Z(n1927) );
  XOR U8017 ( .A(n7708), .B(n6232), .Z(n5282) );
  XOR U8018 ( .A(n8902), .B(n8903), .Z(n6232) );
  XNOR U8019 ( .A(n4751), .B(n2008), .Z(n8903) );
  XOR U8020 ( .A(n8904), .B(n8905), .Z(n2008) );
  ANDN U8021 ( .B(n7860), .A(n7858), .Z(n8904) );
  XOR U8022 ( .A(n8906), .B(n8907), .Z(n4751) );
  ANDN U8023 ( .B(n7868), .A(n7866), .Z(n8906) );
  XOR U8024 ( .A(n6138), .B(n8908), .Z(n8902) );
  XOR U8025 ( .A(n5308), .B(n3817), .Z(n8908) );
  XOR U8026 ( .A(n8909), .B(n8910), .Z(n3817) );
  ANDN U8027 ( .B(n7855), .A(n7853), .Z(n8909) );
  XNOR U8028 ( .A(n8911), .B(n8912), .Z(n5308) );
  AND U8029 ( .A(n7864), .B(n7862), .Z(n8911) );
  XOR U8030 ( .A(n8913), .B(n8914), .Z(n6138) );
  ANDN U8031 ( .B(n7851), .A(n7849), .Z(n8913) );
  XOR U8032 ( .A(n8915), .B(n8916), .Z(n7708) );
  XNOR U8033 ( .A(n4964), .B(n8917), .Z(n8916) );
  XNOR U8034 ( .A(n8918), .B(n7806), .Z(n4964) );
  ANDN U8035 ( .B(n8847), .A(n8919), .Z(n8918) );
  XOR U8036 ( .A(n2297), .B(n8920), .Z(n8915) );
  XOR U8037 ( .A(n3404), .B(n6415), .Z(n8920) );
  XOR U8038 ( .A(n8921), .B(n7792), .Z(n6415) );
  ANDN U8039 ( .B(n8850), .A(n8922), .Z(n8921) );
  XOR U8040 ( .A(n8923), .B(n7797), .Z(n3404) );
  NOR U8041 ( .A(n8845), .B(n8924), .Z(n8923) );
  XOR U8042 ( .A(n8925), .B(n7788), .Z(n2297) );
  ANDN U8043 ( .B(n8854), .A(n8926), .Z(n8925) );
  XNOR U8044 ( .A(n2540), .B(n8927), .Z(n1168) );
  IV U8045 ( .A(n3485), .Z(n2540) );
  XOR U8046 ( .A(n5958), .B(n6381), .Z(n3485) );
  XOR U8047 ( .A(n8928), .B(n8929), .Z(n6381) );
  XNOR U8048 ( .A(n3297), .B(n4903), .Z(n8929) );
  XOR U8049 ( .A(n8930), .B(n6576), .Z(n4903) );
  AND U8050 ( .A(n8884), .B(n6577), .Z(n8930) );
  XOR U8051 ( .A(n8931), .B(n6580), .Z(n3297) );
  ANDN U8052 ( .B(n6581), .A(n8889), .Z(n8931) );
  XOR U8053 ( .A(n5324), .B(n8932), .Z(n8928) );
  XOR U8054 ( .A(n6570), .B(n2581), .Z(n8932) );
  XOR U8055 ( .A(n8933), .B(n6586), .Z(n2581) );
  NOR U8056 ( .A(n8934), .B(n6585), .Z(n8933) );
  XOR U8057 ( .A(n8935), .B(n6589), .Z(n6570) );
  ANDN U8058 ( .B(n6590), .A(n8881), .Z(n8935) );
  XNOR U8059 ( .A(n8936), .B(n6593), .Z(n5324) );
  ANDN U8060 ( .B(n6594), .A(n8892), .Z(n8936) );
  XOR U8061 ( .A(n8937), .B(n8938), .Z(n5958) );
  XOR U8062 ( .A(n3831), .B(n5175), .Z(n8938) );
  XOR U8063 ( .A(n8939), .B(n8940), .Z(n5175) );
  ANDN U8064 ( .B(n8941), .A(n6614), .Z(n8939) );
  XNOR U8065 ( .A(n8942), .B(n8943), .Z(n3831) );
  ANDN U8066 ( .B(n8944), .A(n6601), .Z(n8942) );
  XOR U8067 ( .A(n4214), .B(n8945), .Z(n8937) );
  XOR U8068 ( .A(n1787), .B(n8946), .Z(n8945) );
  XNOR U8069 ( .A(n8947), .B(n8948), .Z(n1787) );
  ANDN U8070 ( .B(n8949), .A(n6605), .Z(n8947) );
  XNOR U8071 ( .A(n8950), .B(n8951), .Z(n4214) );
  AND U8072 ( .A(n6618), .B(n8952), .Z(n8950) );
  XOR U8073 ( .A(n8953), .B(n6090), .Z(out[1034]) );
  XOR U8074 ( .A(n7971), .B(n2469), .Z(n6090) );
  XNOR U8075 ( .A(n8954), .B(n8955), .Z(n2469) );
  IV U8076 ( .A(n8956), .Z(n8954) );
  XNOR U8077 ( .A(n8957), .B(n8958), .Z(n7971) );
  ANDN U8078 ( .B(n8959), .A(n8960), .Z(n8957) );
  ANDN U8079 ( .B(n1172), .A(n1173), .Z(n8953) );
  XNOR U8080 ( .A(n1931), .B(n8961), .Z(n1173) );
  IV U8081 ( .A(n5285), .Z(n1931) );
  XOR U8082 ( .A(n7783), .B(n6237), .Z(n5285) );
  XOR U8083 ( .A(n8962), .B(n8963), .Z(n6237) );
  XNOR U8084 ( .A(n4775), .B(n2012), .Z(n8963) );
  XOR U8085 ( .A(n8964), .B(n8965), .Z(n2012) );
  ANDN U8086 ( .B(n7927), .A(n7925), .Z(n8964) );
  XOR U8087 ( .A(n8966), .B(n8967), .Z(n4775) );
  ANDN U8088 ( .B(n7935), .A(n7933), .Z(n8966) );
  XOR U8089 ( .A(n6144), .B(n8968), .Z(n8962) );
  XOR U8090 ( .A(n5317), .B(n3821), .Z(n8968) );
  XOR U8091 ( .A(n8969), .B(n8970), .Z(n3821) );
  XOR U8092 ( .A(n8971), .B(n8972), .Z(n5317) );
  AND U8093 ( .A(n7931), .B(n7929), .Z(n8971) );
  XOR U8094 ( .A(n8973), .B(n8974), .Z(n6144) );
  AND U8095 ( .A(n7916), .B(n7918), .Z(n8973) );
  XOR U8096 ( .A(n8975), .B(n8976), .Z(n7783) );
  XNOR U8097 ( .A(n4967), .B(n8977), .Z(n8976) );
  XOR U8098 ( .A(n8978), .B(n7867), .Z(n4967) );
  ANDN U8099 ( .B(n8907), .A(n8979), .Z(n8978) );
  XOR U8100 ( .A(n2304), .B(n8980), .Z(n8975) );
  XOR U8101 ( .A(n3406), .B(n6451), .Z(n8980) );
  XOR U8102 ( .A(n8981), .B(n7854), .Z(n6451) );
  ANDN U8103 ( .B(n8910), .A(n8982), .Z(n8981) );
  XOR U8104 ( .A(n8983), .B(n7859), .Z(n3406) );
  ANDN U8105 ( .B(n8905), .A(n8984), .Z(n8983) );
  XOR U8106 ( .A(n8985), .B(n7850), .Z(n2304) );
  XNOR U8107 ( .A(n2551), .B(n8987), .Z(n1172) );
  IV U8108 ( .A(n3488), .Z(n2551) );
  XOR U8109 ( .A(n5963), .B(n6385), .Z(n3488) );
  XOR U8110 ( .A(n8988), .B(n8989), .Z(n6385) );
  XNOR U8111 ( .A(n3300), .B(n4945), .Z(n8989) );
  XOR U8112 ( .A(n8990), .B(n6602), .Z(n4945) );
  ANDN U8113 ( .B(n6603), .A(n8943), .Z(n8990) );
  XOR U8114 ( .A(n8991), .B(n6606), .Z(n3300) );
  ANDN U8115 ( .B(n6607), .A(n8948), .Z(n8991) );
  XOR U8116 ( .A(n5331), .B(n8992), .Z(n8988) );
  XOR U8117 ( .A(n6596), .B(n2588), .Z(n8992) );
  XOR U8118 ( .A(n8993), .B(n6611), .Z(n2588) );
  ANDN U8119 ( .B(n6612), .A(n8994), .Z(n8993) );
  XOR U8120 ( .A(n8995), .B(n6615), .Z(n6596) );
  ANDN U8121 ( .B(n6616), .A(n8940), .Z(n8995) );
  XNOR U8122 ( .A(n8996), .B(n6619), .Z(n5331) );
  ANDN U8123 ( .B(n6620), .A(n8951), .Z(n8996) );
  XOR U8124 ( .A(n8997), .B(n8998), .Z(n5963) );
  XNOR U8125 ( .A(n3835), .B(n5178), .Z(n8998) );
  XOR U8126 ( .A(n8999), .B(n9000), .Z(n5178) );
  XOR U8127 ( .A(n9002), .B(n9003), .Z(n3835) );
  ANDN U8128 ( .B(n9004), .A(n6640), .Z(n9002) );
  XOR U8129 ( .A(n4216), .B(n9005), .Z(n8997) );
  XOR U8130 ( .A(n1791), .B(n9006), .Z(n9005) );
  XNOR U8131 ( .A(n9007), .B(n9008), .Z(n1791) );
  ANDN U8132 ( .B(n9009), .A(n6644), .Z(n9007) );
  XNOR U8133 ( .A(n9010), .B(n9011), .Z(n4216) );
  AND U8134 ( .A(n6627), .B(n9012), .Z(n9010) );
  XOR U8135 ( .A(n9013), .B(n6095), .Z(out[1033]) );
  XNOR U8136 ( .A(n8060), .B(n2480), .Z(n6095) );
  XNOR U8137 ( .A(n9016), .B(n9017), .Z(n8060) );
  AND U8138 ( .A(n9018), .B(n9019), .Z(n9016) );
  ANDN U8139 ( .B(n1180), .A(n1181), .Z(n9013) );
  XNOR U8140 ( .A(n1936), .B(n9020), .Z(n1181) );
  IV U8141 ( .A(n5288), .Z(n1936) );
  XOR U8142 ( .A(n7845), .B(n6242), .Z(n5288) );
  XOR U8143 ( .A(n9021), .B(n9022), .Z(n6242) );
  XNOR U8144 ( .A(n4800), .B(n2016), .Z(n9022) );
  XOR U8145 ( .A(n9023), .B(n9024), .Z(n2016) );
  ANDN U8146 ( .B(n8035), .A(n8033), .Z(n9023) );
  XOR U8147 ( .A(n9025), .B(n9026), .Z(n4800) );
  AND U8148 ( .A(n8041), .B(n9027), .Z(n9025) );
  XOR U8149 ( .A(n6149), .B(n9028), .Z(n9021) );
  XNOR U8150 ( .A(n5321), .B(n3825), .Z(n9028) );
  XNOR U8151 ( .A(n9029), .B(n9030), .Z(n3825) );
  XNOR U8152 ( .A(n9031), .B(n9032), .Z(n5321) );
  AND U8153 ( .A(n8039), .B(n8037), .Z(n9031) );
  XOR U8154 ( .A(n9033), .B(n9034), .Z(n6149) );
  AND U8155 ( .A(n8024), .B(n8026), .Z(n9033) );
  XOR U8156 ( .A(n9035), .B(n9036), .Z(n7845) );
  XNOR U8157 ( .A(n4970), .B(n9037), .Z(n9036) );
  XOR U8158 ( .A(n9038), .B(n7934), .Z(n4970) );
  ANDN U8159 ( .B(n8967), .A(n9039), .Z(n9038) );
  XOR U8160 ( .A(n2311), .B(n9040), .Z(n9035) );
  XOR U8161 ( .A(n3408), .B(n6677), .Z(n9040) );
  XOR U8162 ( .A(n9041), .B(n7921), .Z(n6677) );
  ANDN U8163 ( .B(n8970), .A(n9042), .Z(n9041) );
  XOR U8164 ( .A(n9043), .B(n7926), .Z(n3408) );
  ANDN U8165 ( .B(n8965), .A(n9044), .Z(n9043) );
  XOR U8166 ( .A(n9045), .B(n7917), .Z(n2311) );
  ANDN U8167 ( .B(n8974), .A(n9046), .Z(n9045) );
  XNOR U8168 ( .A(n2558), .B(n9047), .Z(n1180) );
  IV U8169 ( .A(n3491), .Z(n2558) );
  XOR U8170 ( .A(n5968), .B(n6389), .Z(n3491) );
  XOR U8171 ( .A(n9048), .B(n9049), .Z(n6389) );
  XNOR U8172 ( .A(n3303), .B(n4980), .Z(n9049) );
  XOR U8173 ( .A(n9050), .B(n6641), .Z(n4980) );
  AND U8174 ( .A(n9003), .B(n6642), .Z(n9050) );
  XOR U8175 ( .A(n9051), .B(n6646), .Z(n3303) );
  NOR U8176 ( .A(n9008), .B(n6645), .Z(n9051) );
  XOR U8177 ( .A(n5337), .B(n9052), .Z(n9048) );
  XOR U8178 ( .A(n6622), .B(n2595), .Z(n9052) );
  XNOR U8179 ( .A(n9053), .B(n6632), .Z(n2595) );
  ANDN U8180 ( .B(n6633), .A(n9054), .Z(n9053) );
  XOR U8181 ( .A(n9055), .B(n6637), .Z(n6622) );
  AND U8182 ( .A(n9000), .B(n6638), .Z(n9055) );
  XNOR U8183 ( .A(n9056), .B(n6628), .Z(n5337) );
  ANDN U8184 ( .B(n6629), .A(n9011), .Z(n9056) );
  XOR U8185 ( .A(n9057), .B(n9058), .Z(n5968) );
  XNOR U8186 ( .A(n3839), .B(n5182), .Z(n9058) );
  XNOR U8187 ( .A(n9059), .B(n7135), .Z(n5182) );
  ANDN U8188 ( .B(n7136), .A(n6662), .Z(n9059) );
  XNOR U8189 ( .A(n9060), .B(n9061), .Z(n3839) );
  ANDN U8190 ( .B(n9062), .A(n6666), .Z(n9060) );
  XOR U8191 ( .A(n4220), .B(n9063), .Z(n9057) );
  XNOR U8192 ( .A(n7115), .B(n1796), .Z(n9063) );
  XNOR U8193 ( .A(n9064), .B(n7132), .Z(n1796) );
  ANDN U8194 ( .B(n7133), .A(n6670), .Z(n9064) );
  XOR U8195 ( .A(n9065), .B(n7143), .Z(n7115) );
  ANDN U8196 ( .B(n7144), .A(n6657), .Z(n9065) );
  XNOR U8197 ( .A(n9066), .B(n7140), .Z(n4220) );
  AND U8198 ( .A(n6653), .B(n7141), .Z(n9066) );
  XOR U8199 ( .A(n9067), .B(n6101), .Z(out[1032]) );
  XOR U8200 ( .A(n8127), .B(n2487), .Z(n6101) );
  XNOR U8201 ( .A(n9068), .B(n9069), .Z(n2487) );
  XNOR U8202 ( .A(n9070), .B(n9071), .Z(n8127) );
  ANDN U8203 ( .B(n9072), .A(n9073), .Z(n9070) );
  ANDN U8204 ( .B(n1186), .A(n1184), .Z(n9067) );
  XOR U8205 ( .A(n2565), .B(n7137), .Z(n1184) );
  XNOR U8206 ( .A(n9074), .B(n6667), .Z(n7137) );
  ANDN U8207 ( .B(n9061), .A(n9062), .Z(n9074) );
  IV U8208 ( .A(n4858), .Z(n2565) );
  XOR U8209 ( .A(n6393), .B(n5973), .Z(n4858) );
  XOR U8210 ( .A(n9075), .B(n9076), .Z(n5973) );
  XNOR U8211 ( .A(n3843), .B(n5184), .Z(n9076) );
  XOR U8212 ( .A(n9077), .B(n9078), .Z(n5184) );
  NOR U8213 ( .A(n7119), .B(n6694), .Z(n9077) );
  XOR U8214 ( .A(round_reg[1327]), .B(n9079), .Z(n6694) );
  XNOR U8215 ( .A(round_reg[82]), .B(n9080), .Z(n7119) );
  XOR U8216 ( .A(n9081), .B(n9082), .Z(n3843) );
  NOR U8217 ( .A(n7128), .B(n6698), .Z(n9081) );
  XOR U8218 ( .A(round_reg[1420]), .B(n9083), .Z(n6698) );
  XOR U8219 ( .A(n4223), .B(n9084), .Z(n9075) );
  XOR U8220 ( .A(n1799), .B(n7172), .Z(n9084) );
  XOR U8221 ( .A(n9085), .B(n9086), .Z(n7172) );
  XOR U8222 ( .A(round_reg[1546]), .B(n9087), .Z(n6689) );
  XOR U8223 ( .A(round_reg[60]), .B(n9088), .Z(n7124) );
  XOR U8224 ( .A(n9089), .B(n9090), .Z(n1799) );
  NOR U8225 ( .A(n7126), .B(n6702), .Z(n9089) );
  XOR U8226 ( .A(round_reg[1481]), .B(n9091), .Z(n6702) );
  XNOR U8227 ( .A(round_reg[312]), .B(n9092), .Z(n7126) );
  XOR U8228 ( .A(n9093), .B(n7197), .Z(n4223) );
  NOR U8229 ( .A(n7121), .B(n6685), .Z(n9093) );
  XOR U8230 ( .A(round_reg[1390]), .B(n9094), .Z(n6685) );
  XOR U8231 ( .A(round_reg[141]), .B(n9095), .Z(n7121) );
  XOR U8232 ( .A(n9096), .B(n9097), .Z(n6393) );
  XNOR U8233 ( .A(n3310), .B(n5108), .Z(n9097) );
  XOR U8234 ( .A(n9098), .B(n6668), .Z(n5108) );
  NOR U8235 ( .A(n6667), .B(n9061), .Z(n9098) );
  XOR U8236 ( .A(round_reg[610]), .B(n9099), .Z(n9061) );
  XOR U8237 ( .A(round_reg[676]), .B(n9100), .Z(n6667) );
  XOR U8238 ( .A(n9101), .B(n9102), .Z(n3310) );
  NOR U8239 ( .A(n6671), .B(n7132), .Z(n9101) );
  XOR U8240 ( .A(round_reg[323]), .B(n9103), .Z(n7132) );
  XOR U8241 ( .A(round_reg[754]), .B(n9104), .Z(n6671) );
  XOR U8242 ( .A(n5342), .B(n9105), .Z(n9096) );
  XOR U8243 ( .A(n6648), .B(n2602), .Z(n9105) );
  XOR U8244 ( .A(n9106), .B(n9107), .Z(n2602) );
  NOR U8245 ( .A(n6658), .B(n7143), .Z(n9106) );
  XOR U8246 ( .A(round_reg[438]), .B(n9108), .Z(n7143) );
  XOR U8247 ( .A(round_reg[800]), .B(n9109), .Z(n6658) );
  XOR U8248 ( .A(n9110), .B(n9111), .Z(n6648) );
  NOR U8249 ( .A(n6663), .B(n7135), .Z(n9110) );
  XOR U8250 ( .A(round_reg[508]), .B(n9112), .Z(n7135) );
  XOR U8251 ( .A(round_reg[833]), .B(n9113), .Z(n6663) );
  XOR U8252 ( .A(n9114), .B(n6655), .Z(n5342) );
  XOR U8253 ( .A(round_reg[542]), .B(n9115), .Z(n7140) );
  XOR U8254 ( .A(round_reg[904]), .B(n9116), .Z(n6654) );
  XOR U8255 ( .A(n9117), .B(n1941), .Z(n1186) );
  XOR U8256 ( .A(n9118), .B(n9119), .Z(n7912) );
  XNOR U8257 ( .A(n4973), .B(n9120), .Z(n9119) );
  XOR U8258 ( .A(n9121), .B(n8042), .Z(n4973) );
  ANDN U8259 ( .B(n9026), .A(n9122), .Z(n9121) );
  XOR U8260 ( .A(n2318), .B(n9123), .Z(n9118) );
  XOR U8261 ( .A(n3410), .B(n6960), .Z(n9123) );
  XOR U8262 ( .A(n9124), .B(n8029), .Z(n6960) );
  ANDN U8263 ( .B(n9030), .A(n9125), .Z(n9124) );
  IV U8264 ( .A(n9126), .Z(n9030) );
  XOR U8265 ( .A(n9127), .B(n8034), .Z(n3410) );
  ANDN U8266 ( .B(n9024), .A(n9128), .Z(n9127) );
  XOR U8267 ( .A(n9129), .B(n8025), .Z(n2318) );
  ANDN U8268 ( .B(n9034), .A(n9130), .Z(n9129) );
  XNOR U8269 ( .A(n9131), .B(n9132), .Z(n6248) );
  XOR U8270 ( .A(n9133), .B(n3829), .Z(n9132) );
  XNOR U8271 ( .A(n9134), .B(n9135), .Z(n3829) );
  ANDN U8272 ( .B(n8081), .A(n8079), .Z(n9134) );
  XOR U8273 ( .A(n4830), .B(n9136), .Z(n9131) );
  XOR U8274 ( .A(n2020), .B(n5327), .Z(n9136) );
  XOR U8275 ( .A(n9137), .B(n9138), .Z(n5327) );
  ANDN U8276 ( .B(n8090), .A(n8088), .Z(n9137) );
  XOR U8277 ( .A(n9139), .B(n9140), .Z(n2020) );
  ANDN U8278 ( .B(n8086), .A(n8084), .Z(n9139) );
  XOR U8279 ( .A(n9141), .B(n9142), .Z(n4830) );
  ANDN U8280 ( .B(n8094), .A(n8092), .Z(n9141) );
  XOR U8281 ( .A(n9143), .B(n6112), .Z(out[1031]) );
  XOR U8282 ( .A(n8187), .B(n2492), .Z(n6112) );
  XNOR U8283 ( .A(n9144), .B(n9145), .Z(n2492) );
  XNOR U8284 ( .A(n9146), .B(n9147), .Z(n8187) );
  ANDN U8285 ( .B(n9148), .A(n9149), .Z(n9146) );
  AND U8286 ( .A(n1188), .B(n1190), .Z(n9143) );
  XOR U8287 ( .A(n9150), .B(n1946), .Z(n1190) );
  XOR U8288 ( .A(n9151), .B(n9152), .Z(n8020) );
  XNOR U8289 ( .A(n4976), .B(n9153), .Z(n9152) );
  XOR U8290 ( .A(n9154), .B(n8093), .Z(n4976) );
  ANDN U8291 ( .B(n9142), .A(n9155), .Z(n9154) );
  XOR U8292 ( .A(n2329), .B(n9156), .Z(n9151) );
  XOR U8293 ( .A(n3412), .B(n7293), .Z(n9156) );
  XOR U8294 ( .A(n9157), .B(n8080), .Z(n7293) );
  ANDN U8295 ( .B(n9135), .A(n9158), .Z(n9157) );
  XOR U8296 ( .A(n9159), .B(n8085), .Z(n3412) );
  ANDN U8297 ( .B(n9140), .A(n9160), .Z(n9159) );
  XOR U8298 ( .A(n9161), .B(n8076), .Z(n2329) );
  ANDN U8299 ( .B(n9162), .A(n9163), .Z(n9161) );
  XNOR U8300 ( .A(n9164), .B(n9165), .Z(n6253) );
  XOR U8301 ( .A(n9166), .B(n3833), .Z(n9165) );
  XNOR U8302 ( .A(n9167), .B(n9168), .Z(n3833) );
  ANDN U8303 ( .B(n9169), .A(n8010), .Z(n9167) );
  XOR U8304 ( .A(n4868), .B(n9170), .Z(n9164) );
  XOR U8305 ( .A(n2023), .B(n5334), .Z(n9170) );
  XNOR U8306 ( .A(n9171), .B(n9172), .Z(n5334) );
  XOR U8307 ( .A(n9174), .B(n9175), .Z(n2023) );
  NOR U8308 ( .A(n9176), .B(n8140), .Z(n9174) );
  XOR U8309 ( .A(n9177), .B(n9178), .Z(n4868) );
  XNOR U8310 ( .A(n7193), .B(n2573), .Z(n1188) );
  XOR U8311 ( .A(n5978), .B(n6397), .Z(n2573) );
  XOR U8312 ( .A(n9180), .B(n9181), .Z(n6397) );
  XOR U8313 ( .A(n3313), .B(n5519), .Z(n9181) );
  XOR U8314 ( .A(n9182), .B(n6699), .Z(n5519) );
  XOR U8315 ( .A(round_reg[1043]), .B(n9183), .Z(n6699) );
  AND U8316 ( .A(n6700), .B(n9082), .Z(n9182) );
  IV U8317 ( .A(n9184), .Z(n9082) );
  XNOR U8318 ( .A(n9185), .B(n6703), .Z(n3313) );
  XNOR U8319 ( .A(round_reg[1092]), .B(n9186), .Z(n6703) );
  AND U8320 ( .A(n6704), .B(n9090), .Z(n9185) );
  IV U8321 ( .A(n7191), .Z(n9090) );
  XNOR U8322 ( .A(round_reg[322]), .B(n9187), .Z(n7191) );
  XOR U8323 ( .A(round_reg[753]), .B(n9188), .Z(n6704) );
  XOR U8324 ( .A(n5347), .B(n9189), .Z(n9180) );
  XOR U8325 ( .A(n6680), .B(n2609), .Z(n9189) );
  XNOR U8326 ( .A(n9190), .B(n6690), .Z(n2609) );
  XOR U8327 ( .A(round_reg[1182]), .B(n9115), .Z(n6690) );
  AND U8328 ( .A(n6691), .B(n9086), .Z(n9190) );
  IV U8329 ( .A(n7189), .Z(n9086) );
  XOR U8330 ( .A(round_reg[437]), .B(n9191), .Z(n7189) );
  XOR U8331 ( .A(round_reg[799]), .B(n9192), .Z(n6691) );
  XNOR U8332 ( .A(n9193), .B(n6695), .Z(n6680) );
  XNOR U8333 ( .A(round_reg[1254]), .B(n9194), .Z(n6695) );
  AND U8334 ( .A(n6696), .B(n9078), .Z(n9193) );
  IV U8335 ( .A(n7195), .Z(n9078) );
  XNOR U8336 ( .A(round_reg[507]), .B(n9195), .Z(n7195) );
  XOR U8337 ( .A(round_reg[832]), .B(n9196), .Z(n6696) );
  XNOR U8338 ( .A(n9197), .B(n6686), .Z(n5347) );
  XOR U8339 ( .A(round_reg[1014]), .B(n9198), .Z(n6686) );
  AND U8340 ( .A(n6687), .B(n7197), .Z(n9197) );
  XOR U8341 ( .A(round_reg[541]), .B(n9199), .Z(n7197) );
  XOR U8342 ( .A(round_reg[903]), .B(n9200), .Z(n6687) );
  XOR U8343 ( .A(n9201), .B(n9202), .Z(n5978) );
  XNOR U8344 ( .A(n3847), .B(n5187), .Z(n9202) );
  XOR U8345 ( .A(n9203), .B(n9204), .Z(n5187) );
  ANDN U8346 ( .B(n7181), .A(n6720), .Z(n9203) );
  XNOR U8347 ( .A(round_reg[1326]), .B(n9205), .Z(n6720) );
  XOR U8348 ( .A(n9206), .B(n9207), .Z(n3847) );
  ANDN U8349 ( .B(n7178), .A(n6724), .Z(n9206) );
  XOR U8350 ( .A(round_reg[1419]), .B(n9208), .Z(n6724) );
  XNOR U8351 ( .A(n9209), .B(n9210), .Z(n9201) );
  XOR U8352 ( .A(n7225), .B(n1804), .Z(n9210) );
  XOR U8353 ( .A(n9211), .B(n9212), .Z(n1804) );
  ANDN U8354 ( .B(n7176), .A(n6728), .Z(n9211) );
  XNOR U8355 ( .A(round_reg[1480]), .B(n9213), .Z(n6728) );
  XOR U8356 ( .A(n9214), .B(n9215), .Z(n7225) );
  ANDN U8357 ( .B(n7185), .A(n6715), .Z(n9214) );
  XOR U8358 ( .A(round_reg[1545]), .B(n9216), .Z(n6715) );
  XNOR U8359 ( .A(n9217), .B(n6700), .Z(n7193) );
  XOR U8360 ( .A(round_reg[675]), .B(n9218), .Z(n6700) );
  AND U8361 ( .A(n7128), .B(n9184), .Z(n9217) );
  XOR U8362 ( .A(round_reg[609]), .B(n9219), .Z(n9184) );
  XOR U8363 ( .A(round_reg[200]), .B(n9213), .Z(n7128) );
  XOR U8364 ( .A(n9220), .B(n6117), .Z(out[1030]) );
  XOR U8365 ( .A(n8241), .B(n2499), .Z(n6117) );
  XNOR U8366 ( .A(n9221), .B(n9222), .Z(n2499) );
  XOR U8367 ( .A(n9223), .B(n9224), .Z(n8241) );
  ANDN U8368 ( .B(n9225), .A(n9226), .Z(n9223) );
  ANDN U8369 ( .B(n1192), .A(n1193), .Z(n9220) );
  XNOR U8370 ( .A(n9227), .B(n1951), .Z(n1193) );
  XOR U8371 ( .A(n9228), .B(n9229), .Z(n8071) );
  XNOR U8372 ( .A(n3414), .B(n4985), .Z(n9229) );
  XOR U8373 ( .A(n9230), .B(n8005), .Z(n4985) );
  AND U8374 ( .A(n9178), .B(n8006), .Z(n9230) );
  XOR U8375 ( .A(n9231), .B(n8141), .Z(n3414) );
  AND U8376 ( .A(n9175), .B(n8142), .Z(n9231) );
  XNOR U8377 ( .A(n7995), .B(n9232), .Z(n9228) );
  XOR U8378 ( .A(n7145), .B(n2339), .Z(n9232) );
  XNOR U8379 ( .A(n9233), .B(n8015), .Z(n2339) );
  AND U8380 ( .A(n9234), .B(n8016), .Z(n9233) );
  XOR U8381 ( .A(n9235), .B(n8001), .Z(n7145) );
  ANDN U8382 ( .B(n8002), .A(n9172), .Z(n9235) );
  XNOR U8383 ( .A(n9236), .B(n8011), .Z(n7995) );
  AND U8384 ( .A(n9168), .B(n8012), .Z(n9236) );
  XNOR U8385 ( .A(n9237), .B(n9238), .Z(n6258) );
  XNOR U8386 ( .A(n9239), .B(n3837), .Z(n9238) );
  XNOR U8387 ( .A(n9240), .B(n9241), .Z(n3837) );
  ANDN U8388 ( .B(n9242), .A(n8637), .Z(n9240) );
  XNOR U8389 ( .A(n4902), .B(n9243), .Z(n9237) );
  XNOR U8390 ( .A(n2027), .B(n5340), .Z(n9243) );
  XNOR U8391 ( .A(n9244), .B(n9245), .Z(n5340) );
  ANDN U8392 ( .B(n9246), .A(n8628), .Z(n9244) );
  XOR U8393 ( .A(n9247), .B(n9248), .Z(n2027) );
  ANDN U8394 ( .B(n9249), .A(n8641), .Z(n9247) );
  XOR U8395 ( .A(n9250), .B(n9251), .Z(n4902) );
  ANDN U8396 ( .B(n9252), .A(n8632), .Z(n9250) );
  XNOR U8397 ( .A(n9253), .B(n2580), .Z(n1192) );
  XNOR U8398 ( .A(n5984), .B(n6402), .Z(n2580) );
  XNOR U8399 ( .A(n9254), .B(n9255), .Z(n6402) );
  XOR U8400 ( .A(n2616), .B(n5351), .Z(n9255) );
  XOR U8401 ( .A(n9256), .B(n6712), .Z(n5351) );
  XOR U8402 ( .A(round_reg[1013]), .B(n9257), .Z(n6712) );
  ANDN U8403 ( .B(n6713), .A(n9258), .Z(n9256) );
  XNOR U8404 ( .A(n9259), .B(n6716), .Z(n2616) );
  XOR U8405 ( .A(round_reg[1181]), .B(n9260), .Z(n6716) );
  ANDN U8406 ( .B(n6717), .A(n9215), .Z(n9259) );
  XOR U8407 ( .A(n3316), .B(n9261), .Z(n9254) );
  XOR U8408 ( .A(n5893), .B(n6706), .Z(n9261) );
  XNOR U8409 ( .A(n9262), .B(n6721), .Z(n6706) );
  XOR U8410 ( .A(round_reg[1253]), .B(n9263), .Z(n6721) );
  ANDN U8411 ( .B(n6722), .A(n9204), .Z(n9262) );
  XNOR U8412 ( .A(n9264), .B(n6725), .Z(n5893) );
  XOR U8413 ( .A(round_reg[1042]), .B(n9080), .Z(n6725) );
  ANDN U8414 ( .B(n6726), .A(n9207), .Z(n9264) );
  XNOR U8415 ( .A(n9265), .B(n6729), .Z(n3316) );
  XOR U8416 ( .A(round_reg[1091]), .B(n9266), .Z(n6729) );
  ANDN U8417 ( .B(n6730), .A(n9212), .Z(n9265) );
  XOR U8418 ( .A(n9267), .B(n9268), .Z(n5984) );
  XNOR U8419 ( .A(n3851), .B(n5190), .Z(n9268) );
  XOR U8420 ( .A(n9269), .B(n7280), .Z(n5190) );
  ANDN U8421 ( .B(n7281), .A(n6746), .Z(n9269) );
  XOR U8422 ( .A(n9270), .B(n9271), .Z(n3851) );
  AND U8423 ( .A(n6750), .B(n9272), .Z(n9270) );
  XNOR U8424 ( .A(n4045), .B(n9273), .Z(n9267) );
  XOR U8425 ( .A(n7253), .B(n1808), .Z(n9273) );
  XOR U8426 ( .A(n9274), .B(n7275), .Z(n1808) );
  ANDN U8427 ( .B(n7276), .A(n6754), .Z(n9274) );
  XOR U8428 ( .A(n9275), .B(n7272), .Z(n7253) );
  ANDN U8429 ( .B(n7273), .A(n6741), .Z(n9275) );
  XOR U8430 ( .A(n9276), .B(n7283), .Z(n4045) );
  ANDN U8431 ( .B(n7284), .A(n6737), .Z(n9276) );
  XOR U8432 ( .A(n9277), .B(n4128), .Z(out[102]) );
  IV U8433 ( .A(n4302), .Z(n4128) );
  XOR U8434 ( .A(n7034), .B(n2578), .Z(n4302) );
  XNOR U8435 ( .A(n7937), .B(n9278), .Z(n2578) );
  XOR U8436 ( .A(n9279), .B(n9280), .Z(n7937) );
  XOR U8437 ( .A(n4307), .B(n2200), .Z(n9280) );
  XOR U8438 ( .A(n9281), .B(n9282), .Z(n2200) );
  ANDN U8439 ( .B(n9283), .A(n9284), .Z(n9281) );
  XNOR U8440 ( .A(n9285), .B(n9286), .Z(n4307) );
  XOR U8441 ( .A(n6050), .B(n9287), .Z(n9279) );
  XOR U8442 ( .A(n5561), .B(n3751), .Z(n9287) );
  XNOR U8443 ( .A(n9288), .B(n9289), .Z(n3751) );
  ANDN U8444 ( .B(n7032), .A(n7030), .Z(n9288) );
  XOR U8445 ( .A(n9290), .B(n9291), .Z(n5561) );
  XOR U8446 ( .A(n9292), .B(n9293), .Z(n6050) );
  ANDN U8447 ( .B(n7026), .A(n7028), .Z(n9292) );
  XOR U8448 ( .A(n9294), .B(n9283), .Z(n7034) );
  ANDN U8449 ( .B(n9284), .A(n9295), .Z(n9294) );
  AND U8450 ( .A(n3560), .B(n3562), .Z(n9277) );
  XOR U8451 ( .A(n2352), .B(n9296), .Z(n3562) );
  IV U8452 ( .A(n4993), .Z(n2352) );
  XOR U8453 ( .A(n6257), .B(n9297), .Z(n4993) );
  XOR U8454 ( .A(n9298), .B(n9299), .Z(n6257) );
  XNOR U8455 ( .A(n3207), .B(n6961), .Z(n9299) );
  XOR U8456 ( .A(n9300), .B(n9301), .Z(n6961) );
  ANDN U8457 ( .B(n9302), .A(n9303), .Z(n9300) );
  XNOR U8458 ( .A(n9304), .B(n9305), .Z(n3207) );
  NOR U8459 ( .A(n9306), .B(n9307), .Z(n9304) );
  XOR U8460 ( .A(n5516), .B(n9308), .Z(n9298) );
  XOR U8461 ( .A(n8251), .B(n2385), .Z(n9308) );
  XNOR U8462 ( .A(n9309), .B(n9310), .Z(n2385) );
  ANDN U8463 ( .B(n9311), .A(n9312), .Z(n9309) );
  XNOR U8464 ( .A(n9313), .B(n9314), .Z(n8251) );
  ANDN U8465 ( .B(n9315), .A(n9316), .Z(n9313) );
  XNOR U8466 ( .A(n9317), .B(n9318), .Z(n5516) );
  ANDN U8467 ( .B(n9319), .A(n9320), .Z(n9317) );
  XNOR U8468 ( .A(n7475), .B(n2420), .Z(n3560) );
  XNOR U8469 ( .A(n9321), .B(n9322), .Z(n2420) );
  XOR U8470 ( .A(n9323), .B(n9324), .Z(n7475) );
  ANDN U8471 ( .B(n9325), .A(n9326), .Z(n9323) );
  XOR U8472 ( .A(n9327), .B(n6123), .Z(out[1029]) );
  XOR U8473 ( .A(n8293), .B(n2508), .Z(n6123) );
  XNOR U8474 ( .A(n9328), .B(n9329), .Z(n2508) );
  XNOR U8475 ( .A(n9330), .B(n9331), .Z(n8293) );
  NOR U8476 ( .A(n9332), .B(n9333), .Z(n9330) );
  ANDN U8477 ( .B(n1196), .A(n1197), .Z(n9327) );
  XNOR U8478 ( .A(n9334), .B(n1957), .Z(n1197) );
  XOR U8479 ( .A(n9335), .B(n9336), .Z(n8137) );
  XNOR U8480 ( .A(n3416), .B(n4989), .Z(n9336) );
  XOR U8481 ( .A(n9337), .B(n8633), .Z(n4989) );
  ANDN U8482 ( .B(n8634), .A(n9251), .Z(n9337) );
  XOR U8483 ( .A(n9338), .B(n8642), .Z(n3416) );
  ANDN U8484 ( .B(n8643), .A(n9248), .Z(n9338) );
  XNOR U8485 ( .A(n8623), .B(n9339), .Z(n9335) );
  XOR U8486 ( .A(n7198), .B(n2346), .Z(n9339) );
  XOR U8487 ( .A(n9340), .B(n8646), .Z(n2346) );
  ANDN U8488 ( .B(n8647), .A(n9341), .Z(n9340) );
  XOR U8489 ( .A(n9342), .B(n8629), .Z(n7198) );
  ANDN U8490 ( .B(n8630), .A(n9245), .Z(n9342) );
  XOR U8491 ( .A(n9343), .B(n8638), .Z(n8623) );
  AND U8492 ( .A(n9241), .B(n8639), .Z(n9343) );
  XNOR U8493 ( .A(n9344), .B(n9345), .Z(n6263) );
  XNOR U8494 ( .A(n9346), .B(n3841), .Z(n9345) );
  XOR U8495 ( .A(n9347), .B(n9348), .Z(n3841) );
  ANDN U8496 ( .B(n9349), .A(n9310), .Z(n9347) );
  XNOR U8497 ( .A(n4944), .B(n9350), .Z(n9344) );
  XNOR U8498 ( .A(n2031), .B(n5345), .Z(n9350) );
  XNOR U8499 ( .A(n9351), .B(n9352), .Z(n5345) );
  AND U8500 ( .A(n9301), .B(n9353), .Z(n9351) );
  XNOR U8501 ( .A(n9354), .B(n9355), .Z(n2031) );
  ANDN U8502 ( .B(n9356), .A(n9314), .Z(n9354) );
  XOR U8503 ( .A(n9357), .B(n9358), .Z(n4944) );
  ANDN U8504 ( .B(n9359), .A(n9305), .Z(n9357) );
  XNOR U8505 ( .A(n7278), .B(n2587), .Z(n1196) );
  XNOR U8506 ( .A(n5993), .B(n6407), .Z(n2587) );
  XNOR U8507 ( .A(n9360), .B(n9361), .Z(n6407) );
  XOR U8508 ( .A(n2628), .B(n5355), .Z(n9361) );
  XOR U8509 ( .A(n9362), .B(n6738), .Z(n5355) );
  ANDN U8510 ( .B(n6739), .A(n7283), .Z(n9362) );
  XNOR U8511 ( .A(round_reg[539]), .B(n9363), .Z(n7283) );
  XOR U8512 ( .A(round_reg[901]), .B(n9364), .Z(n6739) );
  XNOR U8513 ( .A(n9365), .B(n6742), .Z(n2628) );
  ANDN U8514 ( .B(n6743), .A(n7272), .Z(n9365) );
  XNOR U8515 ( .A(round_reg[435]), .B(n9366), .Z(n7272) );
  XNOR U8516 ( .A(round_reg[797]), .B(n9367), .Z(n6743) );
  XOR U8517 ( .A(n3319), .B(n9368), .Z(n9360) );
  XOR U8518 ( .A(n6409), .B(n6732), .Z(n9368) );
  XNOR U8519 ( .A(n9369), .B(n6747), .Z(n6732) );
  ANDN U8520 ( .B(n6748), .A(n7280), .Z(n9369) );
  XNOR U8521 ( .A(round_reg[505]), .B(n9370), .Z(n7280) );
  XOR U8522 ( .A(round_reg[894]), .B(n9371), .Z(n6748) );
  XNOR U8523 ( .A(n9372), .B(n6751), .Z(n6409) );
  ANDN U8524 ( .B(n6752), .A(n9271), .Z(n9372) );
  XNOR U8525 ( .A(n9373), .B(n6755), .Z(n3319) );
  ANDN U8526 ( .B(n6756), .A(n7275), .Z(n9373) );
  XNOR U8527 ( .A(round_reg[320]), .B(n9374), .Z(n7275) );
  XOR U8528 ( .A(round_reg[751]), .B(n9375), .Z(n6756) );
  XOR U8529 ( .A(n9376), .B(n9377), .Z(n5993) );
  XOR U8530 ( .A(n3576), .B(n5193), .Z(n9377) );
  XOR U8531 ( .A(n9378), .B(n7344), .Z(n5193) );
  AND U8532 ( .A(n7263), .B(n6783), .Z(n9378) );
  IV U8533 ( .A(n7264), .Z(n6783) );
  XNOR U8534 ( .A(round_reg[1324]), .B(n9379), .Z(n7264) );
  XOR U8535 ( .A(round_reg[79]), .B(n9380), .Z(n7263) );
  XNOR U8536 ( .A(n9381), .B(n9382), .Z(n3576) );
  AND U8537 ( .A(n7266), .B(n6763), .Z(n9381) );
  XOR U8538 ( .A(round_reg[1417]), .B(n9383), .Z(n6763) );
  XNOR U8539 ( .A(n4048), .B(n9384), .Z(n9376) );
  XOR U8540 ( .A(n7321), .B(n1812), .Z(n9384) );
  XOR U8541 ( .A(n9385), .B(n7340), .Z(n1812) );
  AND U8542 ( .A(n7257), .B(n6767), .Z(n9385) );
  XOR U8543 ( .A(round_reg[1478]), .B(n9386), .Z(n6767) );
  XOR U8544 ( .A(round_reg[309]), .B(n9387), .Z(n7257) );
  XOR U8545 ( .A(n9388), .B(n7338), .Z(n7321) );
  AND U8546 ( .A(n6771), .B(n7268), .Z(n9388) );
  XOR U8547 ( .A(round_reg[57]), .B(n9389), .Z(n7268) );
  XOR U8548 ( .A(round_reg[1543]), .B(n9390), .Z(n6771) );
  XOR U8549 ( .A(n9391), .B(n7346), .Z(n4048) );
  AND U8550 ( .A(n7259), .B(n6787), .Z(n9391) );
  IV U8551 ( .A(n7260), .Z(n6787) );
  XNOR U8552 ( .A(round_reg[1387]), .B(n9392), .Z(n7260) );
  XNOR U8553 ( .A(round_reg[138]), .B(n9393), .Z(n7259) );
  XNOR U8554 ( .A(n9394), .B(n6752), .Z(n7278) );
  XOR U8555 ( .A(round_reg[673]), .B(n9395), .Z(n6752) );
  ANDN U8556 ( .B(n9271), .A(n9272), .Z(n9394) );
  XNOR U8557 ( .A(round_reg[607]), .B(n9396), .Z(n9271) );
  XOR U8558 ( .A(n9397), .B(n6129), .Z(out[1028]) );
  XOR U8559 ( .A(n8345), .B(n2515), .Z(n6129) );
  XNOR U8560 ( .A(n9398), .B(n9399), .Z(n2515) );
  XNOR U8561 ( .A(n9400), .B(n9401), .Z(n8345) );
  ANDN U8562 ( .B(n9402), .A(n9403), .Z(n9400) );
  ANDN U8563 ( .B(n1200), .A(n1201), .Z(n9397) );
  XNOR U8564 ( .A(n9404), .B(n1966), .Z(n1201) );
  XOR U8565 ( .A(n9405), .B(n9406), .Z(n8198) );
  XNOR U8566 ( .A(n3422), .B(n4994), .Z(n9406) );
  XNOR U8567 ( .A(n9407), .B(n9306), .Z(n4994) );
  ANDN U8568 ( .B(n9307), .A(n9358), .Z(n9407) );
  XOR U8569 ( .A(n9408), .B(n9315), .Z(n3422) );
  AND U8570 ( .A(n9355), .B(n9316), .Z(n9408) );
  XNOR U8571 ( .A(n9296), .B(n9409), .Z(n9405) );
  XOR U8572 ( .A(n7226), .B(n2353), .Z(n9409) );
  XOR U8573 ( .A(n9410), .B(n9319), .Z(n2353) );
  ANDN U8574 ( .B(n9320), .A(n9411), .Z(n9410) );
  XOR U8575 ( .A(n9412), .B(n9302), .Z(n7226) );
  ANDN U8576 ( .B(n9303), .A(n9352), .Z(n9412) );
  XOR U8577 ( .A(n9413), .B(n9311), .Z(n9296) );
  ANDN U8578 ( .B(n9312), .A(n9348), .Z(n9413) );
  XNOR U8579 ( .A(n9414), .B(n9415), .Z(n6269) );
  XNOR U8580 ( .A(n2035), .B(n3845), .Z(n9415) );
  XOR U8581 ( .A(n9416), .B(n9417), .Z(n3845) );
  ANDN U8582 ( .B(n9418), .A(n9419), .Z(n9416) );
  XOR U8583 ( .A(n9420), .B(n9421), .Z(n2035) );
  ANDN U8584 ( .B(n9422), .A(n9423), .Z(n9420) );
  XNOR U8585 ( .A(n9424), .B(n9425), .Z(n9414) );
  XNOR U8586 ( .A(n5349), .B(n4979), .Z(n9425) );
  XOR U8587 ( .A(n9426), .B(n9427), .Z(n4979) );
  NOR U8588 ( .A(n9428), .B(n9429), .Z(n9426) );
  XNOR U8589 ( .A(n9430), .B(n9431), .Z(n5349) );
  ANDN U8590 ( .B(n9432), .A(n9433), .Z(n9430) );
  XNOR U8591 ( .A(n7342), .B(n2594), .Z(n1200) );
  XNOR U8592 ( .A(n5998), .B(n6420), .Z(n2594) );
  XNOR U8593 ( .A(n9434), .B(n9435), .Z(n6420) );
  XNOR U8594 ( .A(n2636), .B(n5359), .Z(n9435) );
  XNOR U8595 ( .A(n9436), .B(n6788), .Z(n5359) );
  XNOR U8596 ( .A(round_reg[1011]), .B(n9437), .Z(n6788) );
  ANDN U8597 ( .B(n6789), .A(n7346), .Z(n9436) );
  XNOR U8598 ( .A(round_reg[538]), .B(n9438), .Z(n7346) );
  XOR U8599 ( .A(round_reg[900]), .B(n9439), .Z(n6789) );
  XNOR U8600 ( .A(n9440), .B(n6780), .Z(n2636) );
  XNOR U8601 ( .A(round_reg[1179]), .B(n9363), .Z(n6780) );
  ANDN U8602 ( .B(n6781), .A(n7338), .Z(n9440) );
  XNOR U8603 ( .A(round_reg[434]), .B(n9104), .Z(n7338) );
  XOR U8604 ( .A(round_reg[796]), .B(n9441), .Z(n6781) );
  XOR U8605 ( .A(n6758), .B(n9442), .Z(n9434) );
  XNOR U8606 ( .A(n5169), .B(n3322), .Z(n9442) );
  XNOR U8607 ( .A(n9443), .B(n6768), .Z(n3322) );
  XNOR U8608 ( .A(round_reg[1089]), .B(n9444), .Z(n6768) );
  ANDN U8609 ( .B(n6769), .A(n7340), .Z(n9443) );
  XNOR U8610 ( .A(round_reg[383]), .B(n9445), .Z(n7340) );
  XOR U8611 ( .A(round_reg[750]), .B(n9094), .Z(n6769) );
  XNOR U8612 ( .A(n9446), .B(n6764), .Z(n5169) );
  XNOR U8613 ( .A(round_reg[1040]), .B(n9447), .Z(n6764) );
  ANDN U8614 ( .B(n6765), .A(n9382), .Z(n9446) );
  XNOR U8615 ( .A(n9448), .B(n6784), .Z(n6758) );
  XOR U8616 ( .A(round_reg[1251]), .B(n9449), .Z(n6784) );
  ANDN U8617 ( .B(n6785), .A(n7344), .Z(n9448) );
  XNOR U8618 ( .A(round_reg[504]), .B(n9450), .Z(n7344) );
  XOR U8619 ( .A(round_reg[893]), .B(n9451), .Z(n6785) );
  XOR U8620 ( .A(n9452), .B(n9453), .Z(n5998) );
  XNOR U8621 ( .A(n1824), .B(n5197), .Z(n9453) );
  XNOR U8622 ( .A(n9454), .B(n7397), .Z(n5197) );
  ANDN U8623 ( .B(n7330), .A(n6805), .Z(n9454) );
  XNOR U8624 ( .A(round_reg[1323]), .B(n9455), .Z(n6805) );
  XOR U8625 ( .A(round_reg[78]), .B(n9456), .Z(n7330) );
  XNOR U8626 ( .A(n9457), .B(n7393), .Z(n1824) );
  ANDN U8627 ( .B(n7325), .A(n6813), .Z(n9457) );
  XNOR U8628 ( .A(round_reg[1477]), .B(n9458), .Z(n6813) );
  XOR U8629 ( .A(round_reg[308]), .B(n9459), .Z(n7325) );
  XNOR U8630 ( .A(n4051), .B(n9460), .Z(n9452) );
  XOR U8631 ( .A(n7374), .B(n3580), .Z(n9460) );
  XOR U8632 ( .A(n9461), .B(n9462), .Z(n3580) );
  ANDN U8633 ( .B(n7332), .A(n6809), .Z(n9461) );
  XNOR U8634 ( .A(round_reg[1416]), .B(n9463), .Z(n6809) );
  XNOR U8635 ( .A(n9464), .B(n7391), .Z(n7374) );
  ANDN U8636 ( .B(n7334), .A(n6800), .Z(n9464) );
  XOR U8637 ( .A(round_reg[1542]), .B(n9465), .Z(n6800) );
  XOR U8638 ( .A(round_reg[56]), .B(n9466), .Z(n7334) );
  XNOR U8639 ( .A(n9467), .B(n7399), .Z(n4051) );
  ANDN U8640 ( .B(n7327), .A(n6796), .Z(n9467) );
  XNOR U8641 ( .A(round_reg[1386]), .B(n9468), .Z(n6796) );
  XOR U8642 ( .A(round_reg[137]), .B(n9469), .Z(n7327) );
  XNOR U8643 ( .A(n9470), .B(n6765), .Z(n7342) );
  XOR U8644 ( .A(round_reg[672]), .B(n9471), .Z(n6765) );
  ANDN U8645 ( .B(n9382), .A(n7266), .Z(n9470) );
  XOR U8646 ( .A(round_reg[197]), .B(n9472), .Z(n7266) );
  XOR U8647 ( .A(round_reg[606]), .B(n9473), .Z(n9382) );
  XOR U8648 ( .A(n9474), .B(n6135), .Z(out[1027]) );
  XOR U8649 ( .A(n8397), .B(n2522), .Z(n6135) );
  XNOR U8650 ( .A(n9475), .B(n9476), .Z(n2522) );
  XNOR U8651 ( .A(n9477), .B(n9478), .Z(n8397) );
  ANDN U8652 ( .B(n9479), .A(n9480), .Z(n9477) );
  ANDN U8653 ( .B(n1204), .A(n1205), .Z(n9474) );
  XNOR U8654 ( .A(n9481), .B(n1971), .Z(n1205) );
  XOR U8655 ( .A(n9482), .B(n9483), .Z(n8252) );
  XNOR U8656 ( .A(n3424), .B(n4999), .Z(n9483) );
  XOR U8657 ( .A(n9484), .B(n9485), .Z(n4999) );
  ANDN U8658 ( .B(n9486), .A(n9427), .Z(n9484) );
  XOR U8659 ( .A(n9487), .B(n9488), .Z(n3424) );
  ANDN U8660 ( .B(n9489), .A(n9421), .Z(n9487) );
  XNOR U8661 ( .A(n9490), .B(n9491), .Z(n9482) );
  XOR U8662 ( .A(n7285), .B(n2360), .Z(n9491) );
  XOR U8663 ( .A(n9492), .B(n9493), .Z(n2360) );
  ANDN U8664 ( .B(n9494), .A(n9495), .Z(n9492) );
  XOR U8665 ( .A(n9496), .B(n9497), .Z(n7285) );
  ANDN U8666 ( .B(n9498), .A(n9431), .Z(n9496) );
  XNOR U8667 ( .A(n9499), .B(n9500), .Z(n6280) );
  XNOR U8668 ( .A(n2039), .B(n3849), .Z(n9500) );
  XOR U8669 ( .A(n9501), .B(n9502), .Z(n3849) );
  ANDN U8670 ( .B(n9503), .A(n9504), .Z(n9501) );
  XNOR U8671 ( .A(n9505), .B(n9506), .Z(n2039) );
  ANDN U8672 ( .B(n9507), .A(n9508), .Z(n9505) );
  XNOR U8673 ( .A(n9509), .B(n9510), .Z(n9499) );
  XNOR U8674 ( .A(n5353), .B(n5027), .Z(n9510) );
  XOR U8675 ( .A(n9511), .B(n9512), .Z(n5027) );
  ANDN U8676 ( .B(n9513), .A(n9514), .Z(n9511) );
  XNOR U8677 ( .A(n9515), .B(n9516), .Z(n5353) );
  ANDN U8678 ( .B(n9517), .A(n9518), .Z(n9515) );
  XNOR U8679 ( .A(n7395), .B(n2601), .Z(n1204) );
  XNOR U8680 ( .A(n6003), .B(n6424), .Z(n2601) );
  XNOR U8681 ( .A(n9519), .B(n9520), .Z(n6424) );
  XOR U8682 ( .A(n2642), .B(n5364), .Z(n9520) );
  XOR U8683 ( .A(n9521), .B(n6797), .Z(n5364) );
  XOR U8684 ( .A(round_reg[1010]), .B(n9522), .Z(n6797) );
  AND U8685 ( .A(n7399), .B(n6798), .Z(n9521) );
  XOR U8686 ( .A(round_reg[899]), .B(n9523), .Z(n6798) );
  XOR U8687 ( .A(round_reg[537]), .B(n9524), .Z(n7399) );
  XNOR U8688 ( .A(n9525), .B(n6801), .Z(n2642) );
  XOR U8689 ( .A(round_reg[1178]), .B(n9526), .Z(n6801) );
  AND U8690 ( .A(n7391), .B(n6802), .Z(n9525) );
  XOR U8691 ( .A(round_reg[795]), .B(n9527), .Z(n6802) );
  XNOR U8692 ( .A(round_reg[433]), .B(n9188), .Z(n7391) );
  XOR U8693 ( .A(n3326), .B(n9528), .Z(n9519) );
  XNOR U8694 ( .A(n5205), .B(n6791), .Z(n9528) );
  XNOR U8695 ( .A(n9529), .B(n6806), .Z(n6791) );
  XOR U8696 ( .A(round_reg[1250]), .B(n9099), .Z(n6806) );
  AND U8697 ( .A(n7397), .B(n6807), .Z(n9529) );
  XOR U8698 ( .A(round_reg[892]), .B(n9530), .Z(n6807) );
  XOR U8699 ( .A(round_reg[503]), .B(n9531), .Z(n7397) );
  XNOR U8700 ( .A(n9532), .B(n6811), .Z(n5205) );
  XNOR U8701 ( .A(round_reg[1039]), .B(n9380), .Z(n6811) );
  ANDN U8702 ( .B(n6810), .A(n9462), .Z(n9532) );
  XNOR U8703 ( .A(n9533), .B(n6814), .Z(n3326) );
  XOR U8704 ( .A(round_reg[1088]), .B(n9534), .Z(n6814) );
  AND U8705 ( .A(n7393), .B(n6815), .Z(n9533) );
  XOR U8706 ( .A(round_reg[749]), .B(n9535), .Z(n6815) );
  XOR U8707 ( .A(round_reg[382]), .B(n9536), .Z(n7393) );
  XOR U8708 ( .A(n9537), .B(n9538), .Z(n6003) );
  XNOR U8709 ( .A(n1828), .B(n5201), .Z(n9538) );
  XOR U8710 ( .A(n9539), .B(n7468), .Z(n5201) );
  ANDN U8711 ( .B(n7383), .A(n6831), .Z(n9539) );
  XNOR U8712 ( .A(round_reg[1322]), .B(n9540), .Z(n6831) );
  XOR U8713 ( .A(round_reg[77]), .B(n9541), .Z(n7383) );
  XOR U8714 ( .A(n9542), .B(n7464), .Z(n1828) );
  ANDN U8715 ( .B(n7385), .A(n6839), .Z(n9542) );
  XNOR U8716 ( .A(round_reg[1476]), .B(n9543), .Z(n6839) );
  XOR U8717 ( .A(round_reg[307]), .B(n9544), .Z(n7385) );
  XNOR U8718 ( .A(n4054), .B(n9545), .Z(n9537) );
  XOR U8719 ( .A(n7445), .B(n3584), .Z(n9545) );
  XOR U8720 ( .A(n9546), .B(n9547), .Z(n3584) );
  ANDN U8721 ( .B(n7378), .A(n6835), .Z(n9546) );
  XNOR U8722 ( .A(round_reg[1415]), .B(n9548), .Z(n6835) );
  XOR U8723 ( .A(n9549), .B(n7462), .Z(n7445) );
  ANDN U8724 ( .B(n7387), .A(n6826), .Z(n9549) );
  XOR U8725 ( .A(round_reg[1541]), .B(n9364), .Z(n6826) );
  XOR U8726 ( .A(round_reg[55]), .B(n9550), .Z(n7387) );
  XOR U8727 ( .A(n9551), .B(n7470), .Z(n4054) );
  ANDN U8728 ( .B(n7380), .A(n6822), .Z(n9551) );
  XNOR U8729 ( .A(round_reg[1385]), .B(n9552), .Z(n6822) );
  XNOR U8730 ( .A(round_reg[136]), .B(n9463), .Z(n7380) );
  XNOR U8731 ( .A(n9553), .B(n6810), .Z(n7395) );
  XOR U8732 ( .A(round_reg[671]), .B(n9554), .Z(n6810) );
  ANDN U8733 ( .B(n9462), .A(n7332), .Z(n9553) );
  XOR U8734 ( .A(round_reg[196]), .B(n9555), .Z(n7332) );
  XOR U8735 ( .A(round_reg[605]), .B(n9556), .Z(n9462) );
  XOR U8736 ( .A(n9557), .B(n6141), .Z(out[1026]) );
  XOR U8737 ( .A(n8450), .B(n2529), .Z(n6141) );
  XNOR U8738 ( .A(n9558), .B(n9559), .Z(n2529) );
  XNOR U8739 ( .A(n9560), .B(n9561), .Z(n8450) );
  ANDN U8740 ( .B(n9562), .A(n9563), .Z(n9560) );
  ANDN U8741 ( .B(n1208), .A(n1209), .Z(n9557) );
  XOR U8742 ( .A(n9564), .B(n1658), .Z(n1209) );
  XOR U8743 ( .A(n9565), .B(n9566), .Z(n8304) );
  XNOR U8744 ( .A(n3426), .B(n5003), .Z(n9566) );
  XOR U8745 ( .A(n9567), .B(n9568), .Z(n5003) );
  ANDN U8746 ( .B(n9569), .A(n9512), .Z(n9567) );
  XOR U8747 ( .A(n9570), .B(n9571), .Z(n3426) );
  AND U8748 ( .A(n9572), .B(n9506), .Z(n9570) );
  XNOR U8749 ( .A(n9573), .B(n9574), .Z(n9565) );
  XOR U8750 ( .A(n7347), .B(n2367), .Z(n9574) );
  XOR U8751 ( .A(n9575), .B(n9576), .Z(n2367) );
  AND U8752 ( .A(n9577), .B(n9578), .Z(n9575) );
  XOR U8753 ( .A(n9579), .B(n9580), .Z(n7347) );
  ANDN U8754 ( .B(n9581), .A(n9516), .Z(n9579) );
  XNOR U8755 ( .A(n9582), .B(n9583), .Z(n6285) );
  XNOR U8756 ( .A(n2047), .B(n3853), .Z(n9583) );
  XOR U8757 ( .A(n9584), .B(n9585), .Z(n3853) );
  ANDN U8758 ( .B(n9586), .A(n7412), .Z(n9584) );
  XOR U8759 ( .A(n9587), .B(n9588), .Z(n2047) );
  ANDN U8760 ( .B(n9589), .A(n8408), .Z(n9587) );
  XNOR U8761 ( .A(n9590), .B(n9591), .Z(n9582) );
  XOR U8762 ( .A(n5357), .B(n5078), .Z(n9591) );
  XOR U8763 ( .A(n9592), .B(n9593), .Z(n5078) );
  NOR U8764 ( .A(n7406), .B(n9594), .Z(n9592) );
  XNOR U8765 ( .A(n9595), .B(n9596), .Z(n5357) );
  ANDN U8766 ( .B(n9597), .A(n8651), .Z(n9595) );
  XNOR U8767 ( .A(n7466), .B(n2608), .Z(n1208) );
  XNOR U8768 ( .A(n6008), .B(n6428), .Z(n2608) );
  XNOR U8769 ( .A(n9598), .B(n9599), .Z(n6428) );
  XOR U8770 ( .A(n2649), .B(n5373), .Z(n9599) );
  XOR U8771 ( .A(n9600), .B(n6823), .Z(n5373) );
  XOR U8772 ( .A(round_reg[1009]), .B(n9601), .Z(n6823) );
  ANDN U8773 ( .B(n6824), .A(n7470), .Z(n9600) );
  XNOR U8774 ( .A(round_reg[536]), .B(n9602), .Z(n7470) );
  XOR U8775 ( .A(round_reg[898]), .B(n9603), .Z(n6824) );
  XNOR U8776 ( .A(n9604), .B(n6827), .Z(n2649) );
  XOR U8777 ( .A(round_reg[1177]), .B(n9605), .Z(n6827) );
  ANDN U8778 ( .B(n6828), .A(n7462), .Z(n9604) );
  XOR U8779 ( .A(round_reg[432]), .B(n9606), .Z(n7462) );
  XOR U8780 ( .A(round_reg[794]), .B(n9607), .Z(n6828) );
  XOR U8781 ( .A(n3330), .B(n9608), .Z(n9598) );
  XOR U8782 ( .A(n5243), .B(n6817), .Z(n9608) );
  XNOR U8783 ( .A(n9609), .B(n6832), .Z(n6817) );
  XOR U8784 ( .A(round_reg[1249]), .B(n9219), .Z(n6832) );
  ANDN U8785 ( .B(n6833), .A(n7468), .Z(n9609) );
  XNOR U8786 ( .A(round_reg[502]), .B(n9610), .Z(n7468) );
  XOR U8787 ( .A(round_reg[891]), .B(n9611), .Z(n6833) );
  XNOR U8788 ( .A(n9612), .B(n6836), .Z(n5243) );
  XOR U8789 ( .A(round_reg[1038]), .B(n9456), .Z(n6836) );
  ANDN U8790 ( .B(n6837), .A(n9547), .Z(n9612) );
  XNOR U8791 ( .A(n9613), .B(n6840), .Z(n3330) );
  XOR U8792 ( .A(round_reg[1151]), .B(n9614), .Z(n6840) );
  ANDN U8793 ( .B(n6841), .A(n7464), .Z(n9613) );
  XNOR U8794 ( .A(round_reg[381]), .B(n9615), .Z(n7464) );
  XOR U8795 ( .A(round_reg[748]), .B(n9616), .Z(n6841) );
  XOR U8796 ( .A(n9617), .B(n9618), .Z(n6008) );
  XNOR U8797 ( .A(n1832), .B(n5210), .Z(n9618) );
  XOR U8798 ( .A(n9619), .B(n7559), .Z(n5210) );
  ANDN U8799 ( .B(n7454), .A(n6857), .Z(n9619) );
  XNOR U8800 ( .A(round_reg[1321]), .B(n9620), .Z(n6857) );
  XOR U8801 ( .A(round_reg[76]), .B(n9621), .Z(n7454) );
  XOR U8802 ( .A(n9622), .B(n7555), .Z(n1832) );
  ANDN U8803 ( .B(n7456), .A(n6865), .Z(n9622) );
  XNOR U8804 ( .A(round_reg[1475]), .B(n9623), .Z(n6865) );
  XOR U8805 ( .A(round_reg[306]), .B(n9624), .Z(n7456) );
  XNOR U8806 ( .A(n4057), .B(n9625), .Z(n9617) );
  XOR U8807 ( .A(n7535), .B(n3589), .Z(n9625) );
  XOR U8808 ( .A(n9626), .B(n9627), .Z(n3589) );
  ANDN U8809 ( .B(n7449), .A(n6861), .Z(n9626) );
  XNOR U8810 ( .A(round_reg[1414]), .B(n9628), .Z(n6861) );
  ANDN U8811 ( .B(n7458), .A(n6852), .Z(n9629) );
  XOR U8812 ( .A(round_reg[1540]), .B(n9439), .Z(n6852) );
  XNOR U8813 ( .A(round_reg[54]), .B(n9630), .Z(n7458) );
  XNOR U8814 ( .A(n9631), .B(n7561), .Z(n4057) );
  ANDN U8815 ( .B(n7451), .A(n6848), .Z(n9631) );
  XNOR U8816 ( .A(round_reg[1384]), .B(n9632), .Z(n6848) );
  XOR U8817 ( .A(round_reg[135]), .B(n9633), .Z(n7451) );
  XNOR U8818 ( .A(n9634), .B(n6837), .Z(n7466) );
  XOR U8819 ( .A(round_reg[670]), .B(n9635), .Z(n6837) );
  ANDN U8820 ( .B(n9547), .A(n7378), .Z(n9634) );
  XOR U8821 ( .A(round_reg[195]), .B(n9636), .Z(n7378) );
  XNOR U8822 ( .A(round_reg[604]), .B(n9637), .Z(n9547) );
  XOR U8823 ( .A(n9638), .B(n6147), .Z(out[1025]) );
  XOR U8824 ( .A(n8503), .B(n2536), .Z(n6147) );
  XNOR U8825 ( .A(n9639), .B(n9640), .Z(n2536) );
  XNOR U8826 ( .A(n9641), .B(n9642), .Z(n8503) );
  ANDN U8827 ( .B(n1212), .A(n1213), .Z(n9638) );
  XNOR U8828 ( .A(n9645), .B(n1663), .Z(n1213) );
  XNOR U8829 ( .A(n9646), .B(n8356), .Z(n1663) );
  XOR U8830 ( .A(n9647), .B(n9648), .Z(n8356) );
  XNOR U8831 ( .A(n3428), .B(n5008), .Z(n9648) );
  XOR U8832 ( .A(n9649), .B(n7407), .Z(n5008) );
  ANDN U8833 ( .B(n7408), .A(n9593), .Z(n9649) );
  XOR U8834 ( .A(n9650), .B(n8409), .Z(n3428) );
  ANDN U8835 ( .B(n8410), .A(n9588), .Z(n9650) );
  XNOR U8836 ( .A(n2372), .B(n9651), .Z(n9647) );
  XOR U8837 ( .A(n3924), .B(n7400), .Z(n9651) );
  XNOR U8838 ( .A(n9652), .B(n8652), .Z(n7400) );
  AND U8839 ( .A(n9596), .B(n8653), .Z(n9652) );
  XNOR U8840 ( .A(n9653), .B(n7413), .Z(n3924) );
  ANDN U8841 ( .B(n7414), .A(n9585), .Z(n9653) );
  XNOR U8842 ( .A(n9654), .B(n7417), .Z(n2372) );
  ANDN U8843 ( .B(n7418), .A(n9655), .Z(n9654) );
  IV U8844 ( .A(n6290), .Z(n9646) );
  XNOR U8845 ( .A(n9656), .B(n9657), .Z(n6290) );
  XNOR U8846 ( .A(n2051), .B(n3578), .Z(n9657) );
  XOR U8847 ( .A(n9658), .B(n9659), .Z(n3578) );
  ANDN U8848 ( .B(n9660), .A(n7483), .Z(n9658) );
  XOR U8849 ( .A(n9661), .B(n9662), .Z(n2051) );
  ANDN U8850 ( .B(n9663), .A(n8461), .Z(n9661) );
  XNOR U8851 ( .A(n9664), .B(n9665), .Z(n9656) );
  XNOR U8852 ( .A(n5362), .B(n5112), .Z(n9665) );
  XNOR U8853 ( .A(n9666), .B(n9667), .Z(n5112) );
  ANDN U8854 ( .B(n9668), .A(n7477), .Z(n9666) );
  XNOR U8855 ( .A(n9669), .B(n9670), .Z(n5362) );
  AND U8856 ( .A(n9324), .B(n9671), .Z(n9669) );
  XNOR U8857 ( .A(n7557), .B(n2615), .Z(n1212) );
  XNOR U8858 ( .A(n6013), .B(n6432), .Z(n2615) );
  XNOR U8859 ( .A(n9672), .B(n9673), .Z(n6432) );
  XOR U8860 ( .A(n2656), .B(n5378), .Z(n9673) );
  XOR U8861 ( .A(n9674), .B(n6850), .Z(n5378) );
  XOR U8862 ( .A(round_reg[1008]), .B(n9675), .Z(n6850) );
  ANDN U8863 ( .B(n7561), .A(n6849), .Z(n9674) );
  XNOR U8864 ( .A(round_reg[897]), .B(n9676), .Z(n6849) );
  XOR U8865 ( .A(round_reg[535]), .B(n9677), .Z(n7561) );
  XNOR U8866 ( .A(n9678), .B(n6853), .Z(n2656) );
  XOR U8867 ( .A(round_reg[1176]), .B(n9679), .Z(n6853) );
  AND U8868 ( .A(n6854), .B(n7553), .Z(n9678) );
  XNOR U8869 ( .A(round_reg[431]), .B(n9375), .Z(n7553) );
  XOR U8870 ( .A(round_reg[793]), .B(n9680), .Z(n6854) );
  XOR U8871 ( .A(n3334), .B(n9681), .Z(n9672) );
  XNOR U8872 ( .A(n5276), .B(n6843), .Z(n9681) );
  XNOR U8873 ( .A(n9682), .B(n6858), .Z(n6843) );
  XOR U8874 ( .A(round_reg[1248]), .B(n9683), .Z(n6858) );
  ANDN U8875 ( .B(n6859), .A(n7559), .Z(n9682) );
  XNOR U8876 ( .A(round_reg[501]), .B(n9684), .Z(n7559) );
  XOR U8877 ( .A(round_reg[890]), .B(n9685), .Z(n6859) );
  XNOR U8878 ( .A(n9686), .B(n6863), .Z(n5276) );
  XNOR U8879 ( .A(round_reg[1037]), .B(n9541), .Z(n6863) );
  ANDN U8880 ( .B(n6862), .A(n9627), .Z(n9686) );
  XNOR U8881 ( .A(n9687), .B(n6866), .Z(n3334) );
  XOR U8882 ( .A(round_reg[1150]), .B(n9688), .Z(n6866) );
  ANDN U8883 ( .B(n6867), .A(n7555), .Z(n9687) );
  XNOR U8884 ( .A(round_reg[380]), .B(n9088), .Z(n7555) );
  XNOR U8885 ( .A(round_reg[747]), .B(n9392), .Z(n6867) );
  XOR U8886 ( .A(n9689), .B(n9690), .Z(n6013) );
  XNOR U8887 ( .A(n1836), .B(n5214), .Z(n9690) );
  XOR U8888 ( .A(n9691), .B(n7611), .Z(n5214) );
  ANDN U8889 ( .B(n6889), .A(n7544), .Z(n9691) );
  XNOR U8890 ( .A(round_reg[75]), .B(n9692), .Z(n7544) );
  XOR U8891 ( .A(round_reg[1320]), .B(n9693), .Z(n6889) );
  XNOR U8892 ( .A(n9694), .B(n7607), .Z(n1836) );
  ANDN U8893 ( .B(n7546), .A(n6897), .Z(n9694) );
  XNOR U8894 ( .A(round_reg[1474]), .B(n9695), .Z(n6897) );
  XOR U8895 ( .A(round_reg[305]), .B(n9696), .Z(n7546) );
  XNOR U8896 ( .A(n4060), .B(n9697), .Z(n9689) );
  XOR U8897 ( .A(n7588), .B(n3598), .Z(n9697) );
  XOR U8898 ( .A(n9698), .B(n9699), .Z(n3598) );
  ANDN U8899 ( .B(n7539), .A(n6893), .Z(n9698) );
  XNOR U8900 ( .A(round_reg[1413]), .B(n9700), .Z(n6893) );
  AND U8901 ( .A(n7548), .B(n7549), .Z(n9701) );
  XOR U8902 ( .A(round_reg[1539]), .B(n9702), .Z(n7549) );
  XNOR U8903 ( .A(round_reg[53]), .B(n9703), .Z(n7548) );
  XNOR U8904 ( .A(n9704), .B(n7613), .Z(n4060) );
  ANDN U8905 ( .B(n7541), .A(n6874), .Z(n9704) );
  XNOR U8906 ( .A(round_reg[1383]), .B(n9705), .Z(n6874) );
  XOR U8907 ( .A(round_reg[134]), .B(n9706), .Z(n7541) );
  XNOR U8908 ( .A(n9707), .B(n6862), .Z(n7557) );
  XOR U8909 ( .A(round_reg[669]), .B(n9708), .Z(n6862) );
  ANDN U8910 ( .B(n9627), .A(n7449), .Z(n9707) );
  XOR U8911 ( .A(round_reg[194]), .B(n9709), .Z(n7449) );
  XNOR U8912 ( .A(round_reg[603]), .B(n9710), .Z(n9627) );
  XOR U8913 ( .A(n9711), .B(n6152), .Z(out[1024]) );
  XOR U8914 ( .A(n8576), .B(n2543), .Z(n6152) );
  XNOR U8915 ( .A(n9712), .B(n9713), .Z(n2543) );
  XNOR U8916 ( .A(n9714), .B(n9715), .Z(n8576) );
  ANDN U8917 ( .B(n8515), .A(n9716), .Z(n9714) );
  ANDN U8918 ( .B(n1216), .A(n1217), .Z(n9711) );
  XNOR U8919 ( .A(n9717), .B(n1671), .Z(n1217) );
  XNOR U8920 ( .A(n9718), .B(n8648), .Z(n1671) );
  XOR U8921 ( .A(n9719), .B(n9720), .Z(n8648) );
  XNOR U8922 ( .A(n3430), .B(n5012), .Z(n9720) );
  XOR U8923 ( .A(n9721), .B(n7478), .Z(n5012) );
  AND U8924 ( .A(n9667), .B(n7479), .Z(n9721) );
  XOR U8925 ( .A(n9722), .B(n8462), .Z(n3430) );
  ANDN U8926 ( .B(n8463), .A(n9662), .Z(n9722) );
  XNOR U8927 ( .A(n2381), .B(n9723), .Z(n9719) );
  XOR U8928 ( .A(n7471), .B(n3927), .Z(n9723) );
  XOR U8929 ( .A(n9724), .B(n7484), .Z(n3927) );
  ANDN U8930 ( .B(n7485), .A(n9659), .Z(n9724) );
  XNOR U8931 ( .A(n9725), .B(n9326), .Z(n7471) );
  ANDN U8932 ( .B(n9726), .A(n9670), .Z(n9725) );
  XOR U8933 ( .A(n9727), .B(n7488), .Z(n2381) );
  AND U8934 ( .A(n9728), .B(n7489), .Z(n9727) );
  IV U8935 ( .A(n6294), .Z(n9718) );
  XNOR U8936 ( .A(n9729), .B(n9730), .Z(n6294) );
  XNOR U8937 ( .A(n2055), .B(n3582), .Z(n9730) );
  XOR U8938 ( .A(n9731), .B(n9732), .Z(n3582) );
  ANDN U8939 ( .B(n9733), .A(n7527), .Z(n9731) );
  XOR U8940 ( .A(n9734), .B(n9735), .Z(n2055) );
  ANDN U8941 ( .B(n9736), .A(n8534), .Z(n9734) );
  XNOR U8942 ( .A(n9737), .B(n9738), .Z(n9729) );
  XNOR U8943 ( .A(n5371), .B(n5137), .Z(n9738) );
  XOR U8944 ( .A(n9739), .B(n9740), .Z(n5137) );
  NOR U8945 ( .A(n7521), .B(n9741), .Z(n9739) );
  XNOR U8946 ( .A(n9742), .B(n9743), .Z(n5371) );
  AND U8947 ( .A(n9744), .B(n9745), .Z(n9742) );
  XNOR U8948 ( .A(n7609), .B(n2627), .Z(n1216) );
  XNOR U8949 ( .A(n6018), .B(n6436), .Z(n2627) );
  XNOR U8950 ( .A(n9746), .B(n9747), .Z(n6436) );
  XOR U8951 ( .A(n2663), .B(n5384), .Z(n9747) );
  XOR U8952 ( .A(n9748), .B(n6876), .Z(n5384) );
  XOR U8953 ( .A(round_reg[1007]), .B(n9079), .Z(n6876) );
  ANDN U8954 ( .B(n7613), .A(n6875), .Z(n9748) );
  XNOR U8955 ( .A(round_reg[896]), .B(n9749), .Z(n6875) );
  XOR U8956 ( .A(round_reg[534]), .B(n9750), .Z(n7613) );
  XNOR U8957 ( .A(n9751), .B(n6885), .Z(n2663) );
  XOR U8958 ( .A(round_reg[1175]), .B(n9752), .Z(n6885) );
  AND U8959 ( .A(n6886), .B(n7605), .Z(n9751) );
  XNOR U8960 ( .A(round_reg[430]), .B(n9094), .Z(n7605) );
  XOR U8961 ( .A(round_reg[792]), .B(n9753), .Z(n6886) );
  XOR U8962 ( .A(n3338), .B(n9754), .Z(n9746) );
  XNOR U8963 ( .A(n5315), .B(n6869), .Z(n9754) );
  XNOR U8964 ( .A(n9755), .B(n6891), .Z(n6869) );
  XOR U8965 ( .A(round_reg[1247]), .B(n9756), .Z(n6891) );
  NOR U8966 ( .A(n6890), .B(n7611), .Z(n9755) );
  XNOR U8967 ( .A(round_reg[500]), .B(n9757), .Z(n7611) );
  XNOR U8968 ( .A(round_reg[889]), .B(n9758), .Z(n6890) );
  XNOR U8969 ( .A(n9759), .B(n6895), .Z(n5315) );
  XNOR U8970 ( .A(round_reg[1036]), .B(n9621), .Z(n6895) );
  ANDN U8971 ( .B(n6894), .A(n9699), .Z(n9759) );
  XNOR U8972 ( .A(n9760), .B(n6899), .Z(n3338) );
  XOR U8973 ( .A(round_reg[1149]), .B(n9761), .Z(n6899) );
  ANDN U8974 ( .B(n7607), .A(n6898), .Z(n9760) );
  XOR U8975 ( .A(round_reg[746]), .B(n9468), .Z(n6898) );
  XOR U8976 ( .A(round_reg[379]), .B(n9762), .Z(n7607) );
  XOR U8977 ( .A(n9763), .B(n9764), .Z(n6018) );
  XNOR U8978 ( .A(n1840), .B(n5218), .Z(n9764) );
  XOR U8979 ( .A(n9765), .B(n7681), .Z(n5218) );
  ANDN U8980 ( .B(n7592), .A(n6915), .Z(n9765) );
  XNOR U8981 ( .A(round_reg[1319]), .B(n9766), .Z(n6915) );
  XOR U8982 ( .A(round_reg[74]), .B(n9767), .Z(n7592) );
  XOR U8983 ( .A(n9768), .B(n7677), .Z(n1840) );
  ANDN U8984 ( .B(n7599), .A(n6923), .Z(n9768) );
  XNOR U8985 ( .A(round_reg[1473]), .B(n9113), .Z(n6923) );
  XOR U8986 ( .A(round_reg[304]), .B(n9769), .Z(n7599) );
  XNOR U8987 ( .A(n4065), .B(n9770), .Z(n9763) );
  XOR U8988 ( .A(n7659), .B(n3602), .Z(n9770) );
  XOR U8989 ( .A(n9771), .B(n9772), .Z(n3602) );
  ANDN U8990 ( .B(n7597), .A(n6919), .Z(n9771) );
  XNOR U8991 ( .A(round_reg[1412]), .B(n9186), .Z(n6919) );
  XOR U8992 ( .A(n9773), .B(n9774), .Z(n7659) );
  ANDN U8993 ( .B(n7601), .A(n6910), .Z(n9773) );
  XOR U8994 ( .A(round_reg[1538]), .B(n9603), .Z(n6910) );
  XNOR U8995 ( .A(n9775), .B(n7683), .Z(n4065) );
  ANDN U8996 ( .B(n7594), .A(n6906), .Z(n9775) );
  XNOR U8997 ( .A(round_reg[1382]), .B(n9776), .Z(n6906) );
  XNOR U8998 ( .A(round_reg[133]), .B(n9700), .Z(n7594) );
  XNOR U8999 ( .A(n9777), .B(n6894), .Z(n7609) );
  XOR U9000 ( .A(round_reg[668]), .B(n9778), .Z(n6894) );
  ANDN U9001 ( .B(n9699), .A(n7539), .Z(n9777) );
  XOR U9002 ( .A(round_reg[193]), .B(n9779), .Z(n7539) );
  XNOR U9003 ( .A(round_reg[602]), .B(n9780), .Z(n9699) );
  XOR U9004 ( .A(n9781), .B(n6156), .Z(out[1023]) );
  XOR U9005 ( .A(n7679), .B(n2634), .Z(n6156) );
  XNOR U9006 ( .A(n9782), .B(n6920), .Z(n7679) );
  ANDN U9007 ( .B(n9772), .A(n7597), .Z(n9782) );
  XOR U9008 ( .A(round_reg[192]), .B(n9196), .Z(n7597) );
  ANDN U9009 ( .B(n5622), .A(n5620), .Z(n9781) );
  XNOR U9010 ( .A(n9783), .B(n1675), .Z(n5620) );
  XNOR U9011 ( .A(n9784), .B(n9321), .Z(n1675) );
  XOR U9012 ( .A(n9785), .B(n9786), .Z(n9321) );
  XNOR U9013 ( .A(n3432), .B(n5016), .Z(n9786) );
  XOR U9014 ( .A(n9787), .B(n7522), .Z(n5016) );
  ANDN U9015 ( .B(n7523), .A(n9740), .Z(n9787) );
  XOR U9016 ( .A(n9788), .B(n8535), .Z(n3432) );
  ANDN U9017 ( .B(n8536), .A(n9735), .Z(n9788) );
  XNOR U9018 ( .A(n2388), .B(n9789), .Z(n9785) );
  XOR U9019 ( .A(n7516), .B(n3932), .Z(n9789) );
  XOR U9020 ( .A(n9790), .B(n7528), .Z(n3932) );
  ANDN U9021 ( .B(n7529), .A(n9732), .Z(n9790) );
  XNOR U9022 ( .A(n9791), .B(n9792), .Z(n7516) );
  XOR U9023 ( .A(n9794), .B(n7532), .Z(n2388) );
  ANDN U9024 ( .B(n7533), .A(n9795), .Z(n9794) );
  IV U9025 ( .A(n6298), .Z(n9784) );
  XNOR U9026 ( .A(n9796), .B(n9797), .Z(n6298) );
  XNOR U9027 ( .A(n5376), .B(n3587), .Z(n9797) );
  XOR U9028 ( .A(n9798), .B(n9799), .Z(n3587) );
  NOR U9029 ( .A(n7626), .B(n9800), .Z(n9798) );
  XNOR U9030 ( .A(n9801), .B(n9802), .Z(n5376) );
  AND U9031 ( .A(n9803), .B(n9804), .Z(n9801) );
  XNOR U9032 ( .A(n9805), .B(n9806), .Z(n9796) );
  XOR U9033 ( .A(n2059), .B(n5167), .Z(n9806) );
  XOR U9034 ( .A(n9807), .B(n9808), .Z(n5167) );
  ANDN U9035 ( .B(n9809), .A(n7620), .Z(n9807) );
  XOR U9036 ( .A(n9810), .B(n9811), .Z(n2059) );
  ANDN U9037 ( .B(n9812), .A(n8656), .Z(n9810) );
  XNOR U9038 ( .A(n9133), .B(n5328), .Z(n5622) );
  XOR U9039 ( .A(n9813), .B(n8138), .Z(n5328) );
  XNOR U9040 ( .A(n9814), .B(n9815), .Z(n8138) );
  XOR U9041 ( .A(n5406), .B(n3793), .Z(n9815) );
  XOR U9042 ( .A(n9816), .B(n9817), .Z(n3793) );
  AND U9043 ( .A(n8015), .B(n8014), .Z(n9816) );
  XOR U9044 ( .A(round_reg[935]), .B(n9818), .Z(n8015) );
  XNOR U9045 ( .A(n9819), .B(n9820), .Z(n5406) );
  AND U9046 ( .A(n8011), .B(n8010), .Z(n9819) );
  XOR U9047 ( .A(round_reg[1214]), .B(n9371), .Z(n8010) );
  XOR U9048 ( .A(round_reg[831]), .B(n9821), .Z(n8011) );
  XOR U9049 ( .A(n6251), .B(n9822), .Z(n9814) );
  XNOR U9050 ( .A(n2239), .B(n4802), .Z(n9822) );
  XOR U9051 ( .A(n9823), .B(n9176), .Z(n4802) );
  ANDN U9052 ( .B(n8140), .A(n8141), .Z(n9823) );
  XNOR U9053 ( .A(round_reg[864]), .B(n9824), .Z(n8141) );
  XOR U9054 ( .A(round_reg[1222]), .B(n9465), .Z(n8140) );
  XNOR U9055 ( .A(n9825), .B(n9173), .Z(n2239) );
  ANDN U9056 ( .B(n8000), .A(n8001), .Z(n9825) );
  XNOR U9057 ( .A(round_reg[643]), .B(n9826), .Z(n8001) );
  XOR U9058 ( .A(round_reg[1075]), .B(n9827), .Z(n8000) );
  XOR U9059 ( .A(n9828), .B(n9179), .Z(n6251) );
  ANDN U9060 ( .B(n8004), .A(n8005), .Z(n9828) );
  XOR U9061 ( .A(round_reg[1124]), .B(n9830), .Z(n8004) );
  XOR U9062 ( .A(n9831), .B(n9162), .Z(n9133) );
  AND U9063 ( .A(n8075), .B(n9832), .Z(n9831) );
  XOR U9064 ( .A(n9833), .B(n6159), .Z(out[1022]) );
  XOR U9065 ( .A(n7754), .B(n2641), .Z(n6159) );
  XNOR U9066 ( .A(n6028), .B(n6676), .Z(n2641) );
  XNOR U9067 ( .A(n9834), .B(n9835), .Z(n6676) );
  XOR U9068 ( .A(n2677), .B(n5393), .Z(n9835) );
  XOR U9069 ( .A(n9836), .B(n6934), .Z(n5393) );
  XOR U9070 ( .A(round_reg[1005]), .B(n9837), .Z(n6934) );
  ANDN U9071 ( .B(n7758), .A(n6933), .Z(n9836) );
  XNOR U9072 ( .A(round_reg[958]), .B(n9838), .Z(n6933) );
  XNOR U9073 ( .A(n9839), .B(n6941), .Z(n2677) );
  XOR U9074 ( .A(round_reg[1173]), .B(n9840), .Z(n6941) );
  AND U9075 ( .A(n6942), .B(n7750), .Z(n9839) );
  XOR U9076 ( .A(round_reg[790]), .B(n9841), .Z(n6942) );
  XOR U9077 ( .A(n3352), .B(n9842), .Z(n9834) );
  XNOR U9078 ( .A(n5419), .B(n6927), .Z(n9842) );
  XNOR U9079 ( .A(n9843), .B(n6958), .Z(n6927) );
  XOR U9080 ( .A(round_reg[1245]), .B(n9556), .Z(n6958) );
  ANDN U9081 ( .B(n6959), .A(n7756), .Z(n9843) );
  XOR U9082 ( .A(round_reg[887]), .B(n9844), .Z(n6959) );
  XNOR U9083 ( .A(n9845), .B(n6948), .Z(n5419) );
  XNOR U9084 ( .A(round_reg[1034]), .B(n9767), .Z(n6948) );
  ANDN U9085 ( .B(n6947), .A(n9846), .Z(n9845) );
  XNOR U9086 ( .A(n9847), .B(n6951), .Z(n3352) );
  XNOR U9087 ( .A(round_reg[1147]), .B(n9195), .Z(n6951) );
  AND U9088 ( .A(n7752), .B(n6952), .Z(n9847) );
  XOR U9089 ( .A(n9848), .B(n9849), .Z(n6028) );
  XNOR U9090 ( .A(n1848), .B(n5225), .Z(n9849) );
  XOR U9091 ( .A(n9850), .B(n7818), .Z(n5225) );
  ANDN U9092 ( .B(n7736), .A(n7290), .Z(n9850) );
  XNOR U9093 ( .A(round_reg[1317]), .B(n9851), .Z(n7290) );
  XOR U9094 ( .A(round_reg[72]), .B(n9852), .Z(n7736) );
  XNOR U9095 ( .A(n9853), .B(n7814), .Z(n1848) );
  ANDN U9096 ( .B(n7744), .A(n6987), .Z(n9853) );
  XNOR U9097 ( .A(round_reg[1535]), .B(n9854), .Z(n6987) );
  XNOR U9098 ( .A(round_reg[302]), .B(n9855), .Z(n7744) );
  XNOR U9099 ( .A(n4071), .B(n9856), .Z(n9848) );
  XOR U9100 ( .A(n7807), .B(n3610), .Z(n9856) );
  XOR U9101 ( .A(n9857), .B(n9858), .Z(n3610) );
  ANDN U9102 ( .B(n7746), .A(n6983), .Z(n9857) );
  XNOR U9103 ( .A(n9860), .B(n7812), .Z(n7807) );
  AND U9104 ( .A(n7741), .B(n7742), .Z(n9860) );
  XNOR U9105 ( .A(round_reg[1536]), .B(n9749), .Z(n7742) );
  XNOR U9106 ( .A(round_reg[50]), .B(n9861), .Z(n7741) );
  XNOR U9107 ( .A(n9862), .B(n7820), .Z(n4071) );
  ANDN U9108 ( .B(n7738), .A(n6968), .Z(n9862) );
  XNOR U9109 ( .A(round_reg[1380]), .B(n9863), .Z(n6968) );
  XOR U9110 ( .A(round_reg[131]), .B(n9266), .Z(n7738) );
  XNOR U9111 ( .A(n9864), .B(n6947), .Z(n7754) );
  XOR U9112 ( .A(round_reg[666]), .B(n9865), .Z(n6947) );
  ANDN U9113 ( .B(n9846), .A(n7668), .Z(n9864) );
  ANDN U9114 ( .B(n5626), .A(n5624), .Z(n9833) );
  XOR U9115 ( .A(n9866), .B(n1680), .Z(n5624) );
  XNOR U9116 ( .A(n9867), .B(n6302), .Z(n1680) );
  XNOR U9117 ( .A(n9868), .B(n9869), .Z(n6302) );
  XNOR U9118 ( .A(n5381), .B(n3592), .Z(n9869) );
  XOR U9119 ( .A(n9870), .B(n9871), .Z(n3592) );
  ANDN U9120 ( .B(n9872), .A(n7703), .Z(n9870) );
  XNOR U9121 ( .A(n9873), .B(n9874), .Z(n5381) );
  ANDN U9122 ( .B(n9875), .A(n7699), .Z(n9873) );
  XNOR U9123 ( .A(n9876), .B(n9877), .Z(n9868) );
  XOR U9124 ( .A(n2062), .B(n5204), .Z(n9877) );
  XOR U9125 ( .A(n9878), .B(n9879), .Z(n5204) );
  ANDN U9126 ( .B(n9880), .A(n7690), .Z(n9878) );
  XOR U9127 ( .A(n9881), .B(n9882), .Z(n2062) );
  ANDN U9128 ( .B(n9883), .A(n8714), .Z(n9881) );
  XNOR U9129 ( .A(n9166), .B(n5335), .Z(n5626) );
  XOR U9130 ( .A(n9884), .B(n8199), .Z(n5335) );
  XNOR U9131 ( .A(n9885), .B(n9886), .Z(n8199) );
  XOR U9132 ( .A(n5410), .B(n3797), .Z(n9886) );
  XOR U9133 ( .A(n9887), .B(n9888), .Z(n3797) );
  ANDN U9134 ( .B(n8645), .A(n8646), .Z(n9887) );
  XNOR U9135 ( .A(round_reg[934]), .B(n9194), .Z(n8646) );
  IV U9136 ( .A(n9889), .Z(n9194) );
  XNOR U9137 ( .A(n9890), .B(n9242), .Z(n5410) );
  ANDN U9138 ( .B(n8637), .A(n8638), .Z(n9890) );
  XNOR U9139 ( .A(round_reg[830]), .B(n9891), .Z(n8638) );
  XOR U9140 ( .A(round_reg[1213]), .B(n9451), .Z(n8637) );
  XOR U9141 ( .A(n6256), .B(n9892), .Z(n9885) );
  XOR U9142 ( .A(n2253), .B(n4832), .Z(n9892) );
  XNOR U9143 ( .A(n9893), .B(n9249), .Z(n4832) );
  ANDN U9144 ( .B(n8641), .A(n8642), .Z(n9893) );
  XNOR U9145 ( .A(round_reg[863]), .B(n9894), .Z(n8642) );
  XOR U9146 ( .A(round_reg[1221]), .B(n9364), .Z(n8641) );
  XNOR U9147 ( .A(n9895), .B(n9246), .Z(n2253) );
  ANDN U9148 ( .B(n8628), .A(n8629), .Z(n9895) );
  XNOR U9149 ( .A(round_reg[642]), .B(n9187), .Z(n8629) );
  XOR U9150 ( .A(round_reg[1074]), .B(n9896), .Z(n8628) );
  XNOR U9151 ( .A(n9897), .B(n9252), .Z(n6256) );
  ANDN U9152 ( .B(n8632), .A(n8633), .Z(n9897) );
  XNOR U9153 ( .A(round_reg[720]), .B(n9898), .Z(n8633) );
  XNOR U9154 ( .A(round_reg[1123]), .B(n9899), .Z(n8632) );
  XOR U9155 ( .A(n9900), .B(n9234), .Z(n9166) );
  NOR U9156 ( .A(n9817), .B(n8014), .Z(n9900) );
  XOR U9157 ( .A(round_reg[982]), .B(n9901), .Z(n8014) );
  XOR U9158 ( .A(n9902), .B(n6169), .Z(out[1021]) );
  XOR U9159 ( .A(n7816), .B(n2648), .Z(n6169) );
  XNOR U9160 ( .A(n6034), .B(n6955), .Z(n2648) );
  XNOR U9161 ( .A(n9903), .B(n9904), .Z(n6955) );
  XOR U9162 ( .A(n2684), .B(n5398), .Z(n9904) );
  XOR U9163 ( .A(n9905), .B(n6970), .Z(n5398) );
  XNOR U9164 ( .A(round_reg[1004]), .B(n9379), .Z(n6970) );
  ANDN U9165 ( .B(n7820), .A(n6969), .Z(n9905) );
  XNOR U9166 ( .A(round_reg[957]), .B(n9906), .Z(n6969) );
  XOR U9167 ( .A(round_reg[531]), .B(n9907), .Z(n7820) );
  XNOR U9168 ( .A(n9908), .B(n6979), .Z(n2684) );
  XOR U9169 ( .A(round_reg[1172]), .B(n9909), .Z(n6979) );
  ANDN U9170 ( .B(n7812), .A(n6978), .Z(n9908) );
  XNOR U9171 ( .A(round_reg[789]), .B(n9910), .Z(n6978) );
  XOR U9172 ( .A(round_reg[427]), .B(n9392), .Z(n7812) );
  XOR U9173 ( .A(n3357), .B(n9911), .Z(n9903) );
  XNOR U9174 ( .A(n5469), .B(n6963), .Z(n9911) );
  XNOR U9175 ( .A(n9912), .B(n7291), .Z(n6963) );
  XNOR U9176 ( .A(round_reg[1244]), .B(n9637), .Z(n7291) );
  ANDN U9177 ( .B(n7292), .A(n7818), .Z(n9912) );
  XNOR U9178 ( .A(round_reg[497]), .B(n9913), .Z(n7818) );
  XOR U9179 ( .A(round_reg[886]), .B(n9914), .Z(n7292) );
  XNOR U9180 ( .A(n9915), .B(n6985), .Z(n5469) );
  XNOR U9181 ( .A(round_reg[1033]), .B(n9916), .Z(n6985) );
  ANDN U9182 ( .B(n6984), .A(n9858), .Z(n9915) );
  XNOR U9183 ( .A(n9917), .B(n6988), .Z(n3357) );
  XNOR U9184 ( .A(round_reg[1146]), .B(n9918), .Z(n6988) );
  AND U9185 ( .A(n7814), .B(n6989), .Z(n9917) );
  XOR U9186 ( .A(round_reg[743]), .B(n9919), .Z(n6989) );
  XNOR U9187 ( .A(round_reg[376]), .B(n9466), .Z(n7814) );
  XOR U9188 ( .A(n9920), .B(n9921), .Z(n6034) );
  XNOR U9189 ( .A(n5228), .B(n1853), .Z(n9921) );
  AND U9190 ( .A(n7876), .B(n7015), .Z(n9922) );
  XNOR U9191 ( .A(round_reg[1534]), .B(n9371), .Z(n7015) );
  XOR U9192 ( .A(round_reg[301]), .B(n9923), .Z(n7876) );
  XOR U9193 ( .A(n9924), .B(n7883), .Z(n5228) );
  ANDN U9194 ( .B(n7884), .A(n7985), .Z(n9924) );
  XNOR U9195 ( .A(round_reg[1316]), .B(n9100), .Z(n7985) );
  XOR U9196 ( .A(round_reg[71]), .B(n9925), .Z(n7884) );
  XNOR U9197 ( .A(n3614), .B(n9926), .Z(n9920) );
  XOR U9198 ( .A(n7869), .B(n4074), .Z(n9926) );
  XNOR U9199 ( .A(n9927), .B(n7887), .Z(n4074) );
  ANDN U9200 ( .B(n7886), .A(n6996), .Z(n9927) );
  XOR U9201 ( .A(round_reg[130]), .B(n9859), .Z(n7886) );
  XNOR U9202 ( .A(n9929), .B(n7880), .Z(n7869) );
  ANDN U9203 ( .B(n7990), .A(n7879), .Z(n9929) );
  XNOR U9204 ( .A(round_reg[49]), .B(n9601), .Z(n7879) );
  XNOR U9205 ( .A(round_reg[1599]), .B(n9930), .Z(n7990) );
  XOR U9206 ( .A(n9931), .B(n9932), .Z(n3614) );
  ANDN U9207 ( .B(n7011), .A(n7992), .Z(n9931) );
  XOR U9208 ( .A(round_reg[1409]), .B(n9444), .Z(n7011) );
  XNOR U9209 ( .A(n9933), .B(n6984), .Z(n7816) );
  XOR U9210 ( .A(round_reg[665]), .B(n9934), .Z(n6984) );
  ANDN U9211 ( .B(n9858), .A(n7746), .Z(n9933) );
  XOR U9212 ( .A(round_reg[254]), .B(n9371), .Z(n7746) );
  XNOR U9213 ( .A(round_reg[599]), .B(n9935), .Z(n9858) );
  NOR U9214 ( .A(n5629), .B(n5628), .Z(n9902) );
  XOR U9215 ( .A(n9936), .B(n1685), .Z(n5628) );
  XNOR U9216 ( .A(n9937), .B(n6306), .Z(n1685) );
  XNOR U9217 ( .A(n9938), .B(n9939), .Z(n6306) );
  XOR U9218 ( .A(n5386), .B(n3599), .Z(n9939) );
  XOR U9219 ( .A(n9940), .B(n9941), .Z(n3599) );
  ANDN U9220 ( .B(n7778), .A(n9942), .Z(n9940) );
  XNOR U9221 ( .A(n9943), .B(n9944), .Z(n5386) );
  AND U9222 ( .A(n9945), .B(n9946), .Z(n9943) );
  XOR U9223 ( .A(n9947), .B(n9948), .Z(n9938) );
  XOR U9224 ( .A(n2065), .B(n5242), .Z(n9948) );
  XNOR U9225 ( .A(n9949), .B(n9950), .Z(n5242) );
  NOR U9226 ( .A(n9951), .B(n7765), .Z(n9949) );
  XNOR U9227 ( .A(n9952), .B(n9953), .Z(n2065) );
  ANDN U9228 ( .B(n9954), .A(n8775), .Z(n9952) );
  XOR U9229 ( .A(n9239), .B(n2028), .Z(n5629) );
  XNOR U9230 ( .A(n7996), .B(n8253), .Z(n2028) );
  XNOR U9231 ( .A(n9955), .B(n9956), .Z(n8253) );
  XOR U9232 ( .A(n5414), .B(n3801), .Z(n9956) );
  XOR U9233 ( .A(n9957), .B(n9958), .Z(n3801) );
  ANDN U9234 ( .B(n9318), .A(n9319), .Z(n9957) );
  XNOR U9235 ( .A(round_reg[933]), .B(n9959), .Z(n9319) );
  XNOR U9236 ( .A(n9960), .B(n9349), .Z(n5414) );
  ANDN U9237 ( .B(n9310), .A(n9311), .Z(n9960) );
  XNOR U9238 ( .A(round_reg[829]), .B(n9961), .Z(n9311) );
  XOR U9239 ( .A(round_reg[1212]), .B(n9530), .Z(n9310) );
  XOR U9240 ( .A(n6261), .B(n9962), .Z(n9955) );
  XOR U9241 ( .A(n2260), .B(n4869), .Z(n9962) );
  XNOR U9242 ( .A(n9963), .B(n9356), .Z(n4869) );
  ANDN U9243 ( .B(n9314), .A(n9315), .Z(n9963) );
  XOR U9244 ( .A(round_reg[862]), .B(n9115), .Z(n9315) );
  XOR U9245 ( .A(round_reg[1220]), .B(n9439), .Z(n9314) );
  IV U9246 ( .A(n9964), .Z(n9439) );
  XNOR U9247 ( .A(n9965), .B(n9353), .Z(n2260) );
  NOR U9248 ( .A(n9301), .B(n9302), .Z(n9965) );
  XNOR U9249 ( .A(round_reg[641]), .B(n9966), .Z(n9302) );
  XNOR U9250 ( .A(round_reg[1073]), .B(n9188), .Z(n9301) );
  XNOR U9251 ( .A(n9967), .B(n9359), .Z(n6261) );
  AND U9252 ( .A(n9306), .B(n9305), .Z(n9967) );
  XOR U9253 ( .A(round_reg[1122]), .B(n9968), .Z(n9305) );
  XOR U9254 ( .A(round_reg[719]), .B(n9969), .Z(n9306) );
  XOR U9255 ( .A(n9970), .B(n9971), .Z(n7996) );
  XOR U9256 ( .A(n1956), .B(n9334), .Z(n9971) );
  XOR U9257 ( .A(n9972), .B(n8639), .Z(n9334) );
  XOR U9258 ( .A(round_reg[404]), .B(n9973), .Z(n8639) );
  NOR U9259 ( .A(n9241), .B(n9242), .Z(n9972) );
  XOR U9260 ( .A(round_reg[1577]), .B(n9974), .Z(n9242) );
  XNOR U9261 ( .A(round_reg[27]), .B(n9975), .Z(n9241) );
  XNOR U9262 ( .A(n9976), .B(n8634), .Z(n1956) );
  XOR U9263 ( .A(round_reg[353]), .B(n9395), .Z(n8634) );
  ANDN U9264 ( .B(n9251), .A(n9252), .Z(n9976) );
  XOR U9265 ( .A(round_reg[1512]), .B(n9977), .Z(n9252) );
  XNOR U9266 ( .A(round_reg[279]), .B(n9935), .Z(n9251) );
  XOR U9267 ( .A(n3710), .B(n9978), .Z(n9970) );
  XOR U9268 ( .A(n5094), .B(n4144), .Z(n9978) );
  XNOR U9269 ( .A(n9979), .B(n8647), .Z(n4144) );
  XOR U9270 ( .A(round_reg[572]), .B(n9530), .Z(n8647) );
  ANDN U9271 ( .B(n9341), .A(n9888), .Z(n9979) );
  XNOR U9272 ( .A(n9980), .B(n8643), .Z(n5094) );
  XOR U9273 ( .A(round_reg[474]), .B(n9607), .Z(n8643) );
  ANDN U9274 ( .B(n9248), .A(n9249), .Z(n9980) );
  XOR U9275 ( .A(round_reg[1294]), .B(n9981), .Z(n9249) );
  XOR U9276 ( .A(round_reg[113]), .B(n9188), .Z(n9248) );
  XNOR U9277 ( .A(n9982), .B(n8630), .Z(n3710) );
  XOR U9278 ( .A(round_reg[576]), .B(n9749), .Z(n8630) );
  ANDN U9279 ( .B(n9245), .A(n9246), .Z(n9982) );
  XOR U9280 ( .A(round_reg[1451]), .B(n9983), .Z(n9246) );
  XOR U9281 ( .A(round_reg[231]), .B(n9984), .Z(n9245) );
  XOR U9282 ( .A(n9985), .B(n9341), .Z(n9239) );
  XNOR U9283 ( .A(round_reg[172]), .B(n9986), .Z(n9341) );
  ANDN U9284 ( .B(n9888), .A(n8645), .Z(n9985) );
  XOR U9285 ( .A(round_reg[981]), .B(n9987), .Z(n8645) );
  XOR U9286 ( .A(round_reg[1357]), .B(n9541), .Z(n9888) );
  XOR U9287 ( .A(n9988), .B(n6174), .Z(out[1020]) );
  XNOR U9288 ( .A(n7873), .B(n2655), .Z(n6174) );
  XNOR U9289 ( .A(n6039), .B(n7288), .Z(n2655) );
  XNOR U9290 ( .A(n9989), .B(n9990), .Z(n7288) );
  XOR U9291 ( .A(n2691), .B(n5403), .Z(n9990) );
  XNOR U9292 ( .A(n9991), .B(n6998), .Z(n5403) );
  XNOR U9293 ( .A(round_reg[1003]), .B(n9992), .Z(n6998) );
  ANDN U9294 ( .B(n7887), .A(n6997), .Z(n9991) );
  XNOR U9295 ( .A(round_reg[956]), .B(n9993), .Z(n6997) );
  XOR U9296 ( .A(round_reg[530]), .B(n9994), .Z(n7887) );
  XNOR U9297 ( .A(n9995), .B(n7007), .Z(n2691) );
  XOR U9298 ( .A(round_reg[1171]), .B(n9996), .Z(n7007) );
  ANDN U9299 ( .B(n7880), .A(n7006), .Z(n9995) );
  XNOR U9300 ( .A(round_reg[788]), .B(n9997), .Z(n7006) );
  XOR U9301 ( .A(round_reg[426]), .B(n9468), .Z(n7880) );
  XOR U9302 ( .A(n3362), .B(n9998), .Z(n9989) );
  XNOR U9303 ( .A(n5526), .B(n6991), .Z(n9998) );
  XNOR U9304 ( .A(n9999), .B(n7986), .Z(n6991) );
  XOR U9305 ( .A(round_reg[1243]), .B(n10000), .Z(n7986) );
  ANDN U9306 ( .B(n7882), .A(n7883), .Z(n9999) );
  XNOR U9307 ( .A(round_reg[496]), .B(n10001), .Z(n7883) );
  XOR U9308 ( .A(round_reg[885]), .B(n10002), .Z(n7882) );
  XNOR U9309 ( .A(n10003), .B(n7013), .Z(n5526) );
  XNOR U9310 ( .A(round_reg[1032]), .B(n9852), .Z(n7013) );
  ANDN U9311 ( .B(n7012), .A(n9932), .Z(n10003) );
  XNOR U9312 ( .A(n10004), .B(n7016), .Z(n3362) );
  XOR U9313 ( .A(round_reg[1145]), .B(n10005), .Z(n7016) );
  AND U9314 ( .A(n7017), .B(n7875), .Z(n10004) );
  XNOR U9315 ( .A(round_reg[375]), .B(n9550), .Z(n7875) );
  XOR U9316 ( .A(round_reg[742]), .B(n10006), .Z(n7017) );
  XOR U9317 ( .A(n10007), .B(n10008), .Z(n6039) );
  XNOR U9318 ( .A(n5231), .B(n1857), .Z(n10008) );
  XOR U9319 ( .A(n10009), .B(n7943), .Z(n1857) );
  AND U9320 ( .A(n8611), .B(n8609), .Z(n10009) );
  XNOR U9321 ( .A(round_reg[300]), .B(n10010), .Z(n8609) );
  XOR U9322 ( .A(n10011), .B(n7952), .Z(n5231) );
  ANDN U9323 ( .B(n7953), .A(n8606), .Z(n10011) );
  XOR U9324 ( .A(round_reg[70]), .B(n10012), .Z(n7953) );
  XNOR U9325 ( .A(n3618), .B(n10013), .Z(n10007) );
  XOR U9326 ( .A(n7936), .B(n4077), .Z(n10013) );
  XNOR U9327 ( .A(n10014), .B(n7957), .Z(n4077) );
  NOR U9328 ( .A(n7956), .B(n8621), .Z(n10014) );
  XNOR U9329 ( .A(round_reg[129]), .B(n10015), .Z(n7956) );
  XNOR U9330 ( .A(n10016), .B(n7949), .Z(n7936) );
  ANDN U9331 ( .B(n8614), .A(n7948), .Z(n10016) );
  XNOR U9332 ( .A(round_reg[48]), .B(n9675), .Z(n7948) );
  XOR U9333 ( .A(n10017), .B(n10018), .Z(n3618) );
  ANDN U9334 ( .B(n8617), .A(n8619), .Z(n10017) );
  XOR U9335 ( .A(n10019), .B(n7012), .Z(n7873) );
  XNOR U9336 ( .A(round_reg[664]), .B(n10020), .Z(n7012) );
  AND U9337 ( .A(n7992), .B(n9932), .Z(n10019) );
  XNOR U9338 ( .A(round_reg[598]), .B(n10021), .Z(n9932) );
  XNOR U9339 ( .A(round_reg[253]), .B(n9451), .Z(n7992) );
  ANDN U9340 ( .B(n5632), .A(n5633), .Z(n9988) );
  XOR U9341 ( .A(n9346), .B(n2032), .Z(n5633) );
  XNOR U9342 ( .A(n8624), .B(n8305), .Z(n2032) );
  XNOR U9343 ( .A(n10022), .B(n10023), .Z(n8305) );
  XOR U9344 ( .A(n5422), .B(n3806), .Z(n10023) );
  XOR U9345 ( .A(n10024), .B(n10025), .Z(n3806) );
  ANDN U9346 ( .B(n10026), .A(n9493), .Z(n10024) );
  XNOR U9347 ( .A(n10027), .B(n9418), .Z(n5422) );
  ANDN U9348 ( .B(n9419), .A(n10028), .Z(n10027) );
  XNOR U9349 ( .A(n6267), .B(n10029), .Z(n10022) );
  XOR U9350 ( .A(n2267), .B(n4904), .Z(n10029) );
  XNOR U9351 ( .A(n10030), .B(n9422), .Z(n4904) );
  ANDN U9352 ( .B(n9423), .A(n9488), .Z(n10030) );
  XNOR U9353 ( .A(n10031), .B(n9432), .Z(n2267) );
  ANDN U9354 ( .B(n9433), .A(n9497), .Z(n10031) );
  XNOR U9355 ( .A(n10032), .B(n9429), .Z(n6267) );
  ANDN U9356 ( .B(n9428), .A(n9485), .Z(n10032) );
  XOR U9357 ( .A(n10033), .B(n10034), .Z(n8624) );
  XOR U9358 ( .A(n1965), .B(n9404), .Z(n10034) );
  XOR U9359 ( .A(n10035), .B(n9312), .Z(n9404) );
  XOR U9360 ( .A(round_reg[403]), .B(n9183), .Z(n9312) );
  ANDN U9361 ( .B(n9348), .A(n9349), .Z(n10035) );
  XOR U9362 ( .A(round_reg[1576]), .B(n10036), .Z(n9349) );
  XOR U9363 ( .A(round_reg[26]), .B(n9865), .Z(n9348) );
  XNOR U9364 ( .A(n10037), .B(n9307), .Z(n1965) );
  XOR U9365 ( .A(round_reg[352]), .B(n9471), .Z(n9307) );
  ANDN U9366 ( .B(n9358), .A(n9359), .Z(n10037) );
  XOR U9367 ( .A(round_reg[1511]), .B(n9984), .Z(n9359) );
  XNOR U9368 ( .A(round_reg[278]), .B(n10021), .Z(n9358) );
  XOR U9369 ( .A(n3714), .B(n10038), .Z(n10033) );
  XOR U9370 ( .A(n5096), .B(n4147), .Z(n10038) );
  XNOR U9371 ( .A(n10039), .B(n9320), .Z(n4147) );
  XOR U9372 ( .A(round_reg[571]), .B(n9611), .Z(n9320) );
  ANDN U9373 ( .B(n9411), .A(n9958), .Z(n10039) );
  XNOR U9374 ( .A(n10040), .B(n9316), .Z(n5096) );
  XNOR U9375 ( .A(round_reg[473]), .B(n10041), .Z(n9316) );
  NOR U9376 ( .A(n9355), .B(n9356), .Z(n10040) );
  XOR U9377 ( .A(round_reg[1293]), .B(n10042), .Z(n9356) );
  XNOR U9378 ( .A(round_reg[112]), .B(n9606), .Z(n9355) );
  XNOR U9379 ( .A(n10043), .B(n9303), .Z(n3714) );
  XOR U9380 ( .A(round_reg[639]), .B(n9930), .Z(n9303) );
  ANDN U9381 ( .B(n9352), .A(n9353), .Z(n10043) );
  XOR U9382 ( .A(round_reg[1450]), .B(n10044), .Z(n9353) );
  XOR U9383 ( .A(round_reg[230]), .B(n10045), .Z(n9352) );
  XOR U9384 ( .A(n10046), .B(n9411), .Z(n9346) );
  XNOR U9385 ( .A(round_reg[171]), .B(n10047), .Z(n9411) );
  ANDN U9386 ( .B(n9958), .A(n9318), .Z(n10046) );
  XOR U9387 ( .A(round_reg[980]), .B(n10048), .Z(n9318) );
  XOR U9388 ( .A(round_reg[1356]), .B(n9621), .Z(n9958) );
  XOR U9389 ( .A(n10049), .B(n1690), .Z(n5632) );
  XNOR U9390 ( .A(n8718), .B(n6310), .Z(n1690) );
  XNOR U9391 ( .A(n10050), .B(n10051), .Z(n6310) );
  XNOR U9392 ( .A(n5390), .B(n3604), .Z(n10051) );
  XOR U9393 ( .A(n10052), .B(n10053), .Z(n3604) );
  AND U9394 ( .A(n7836), .B(n10054), .Z(n10052) );
  IV U9395 ( .A(n10055), .Z(n7836) );
  XNOR U9396 ( .A(n10056), .B(n10057), .Z(n5390) );
  AND U9397 ( .A(n10058), .B(n7826), .Z(n10056) );
  XNOR U9398 ( .A(n10059), .B(n10060), .Z(n10050) );
  XOR U9399 ( .A(n2069), .B(n5275), .Z(n10060) );
  XNOR U9400 ( .A(n10061), .B(n10062), .Z(n5275) );
  ANDN U9401 ( .B(n7830), .A(n10063), .Z(n10061) );
  XNOR U9402 ( .A(n10064), .B(n10065), .Z(n2069) );
  AND U9403 ( .A(n10066), .B(n8838), .Z(n10064) );
  IV U9404 ( .A(n10067), .Z(n8838) );
  XOR U9405 ( .A(n10068), .B(n10069), .Z(n8718) );
  XNOR U9406 ( .A(n5030), .B(n7759), .Z(n10069) );
  XOR U9407 ( .A(n10070), .B(n7776), .Z(n7759) );
  ANDN U9408 ( .B(n7775), .A(n9944), .Z(n10070) );
  XNOR U9409 ( .A(n10071), .B(n7766), .Z(n5030) );
  ANDN U9410 ( .B(n7767), .A(n9950), .Z(n10071) );
  XOR U9411 ( .A(n2410), .B(n10072), .Z(n10068) );
  XOR U9412 ( .A(n3438), .B(n3941), .Z(n10072) );
  XNOR U9413 ( .A(n10073), .B(n7779), .Z(n3941) );
  ANDN U9414 ( .B(n7780), .A(n9941), .Z(n10073) );
  XNOR U9415 ( .A(n10074), .B(n8777), .Z(n3438) );
  NOR U9416 ( .A(n8776), .B(n9953), .Z(n10074) );
  XNOR U9417 ( .A(n10075), .B(n7771), .Z(n2410) );
  ANDN U9418 ( .B(n7772), .A(n10076), .Z(n10075) );
  XOR U9419 ( .A(n10077), .B(n4133), .Z(out[101]) );
  IV U9420 ( .A(n4305), .Z(n4133) );
  XOR U9421 ( .A(n7057), .B(n2585), .Z(n4305) );
  XNOR U9422 ( .A(n8046), .B(n10078), .Z(n2585) );
  XOR U9423 ( .A(n10079), .B(n10080), .Z(n8046) );
  XOR U9424 ( .A(n4310), .B(n2203), .Z(n10080) );
  XOR U9425 ( .A(n10081), .B(n8110), .Z(n2203) );
  ANDN U9426 ( .B(n10082), .A(n10083), .Z(n10081) );
  XOR U9427 ( .A(n10084), .B(n8102), .Z(n4310) );
  IV U9428 ( .A(n10085), .Z(n8102) );
  XOR U9429 ( .A(n6055), .B(n10086), .Z(n10079) );
  XOR U9430 ( .A(n5565), .B(n3755), .Z(n10086) );
  XNOR U9431 ( .A(n10087), .B(n8105), .Z(n3755) );
  ANDN U9432 ( .B(n7055), .A(n7053), .Z(n10087) );
  XOR U9433 ( .A(n10088), .B(n10089), .Z(n5565) );
  XOR U9434 ( .A(n10090), .B(n8112), .Z(n6055) );
  ANDN U9435 ( .B(n7049), .A(n7051), .Z(n10090) );
  XOR U9436 ( .A(n10091), .B(n10082), .Z(n7057) );
  ANDN U9437 ( .B(n10083), .A(n8108), .Z(n10091) );
  AND U9438 ( .A(n3594), .B(n3596), .Z(n10077) );
  XOR U9439 ( .A(n2359), .B(n9490), .Z(n3596) );
  XOR U9440 ( .A(n10092), .B(n10028), .Z(n9490) );
  ANDN U9441 ( .B(n10093), .A(n9417), .Z(n10092) );
  IV U9442 ( .A(n4998), .Z(n2359) );
  XOR U9443 ( .A(n6262), .B(n10094), .Z(n4998) );
  XOR U9444 ( .A(n10095), .B(n10096), .Z(n6262) );
  XOR U9445 ( .A(n3210), .B(n7294), .Z(n10096) );
  XOR U9446 ( .A(n10097), .B(n9433), .Z(n7294) );
  XOR U9447 ( .A(round_reg[1072]), .B(n9606), .Z(n9433) );
  ANDN U9448 ( .B(n9497), .A(n9498), .Z(n10097) );
  XNOR U9449 ( .A(round_reg[640]), .B(n9374), .Z(n9497) );
  XNOR U9450 ( .A(n10098), .B(n9428), .Z(n3210) );
  XOR U9451 ( .A(round_reg[1121]), .B(n10099), .Z(n9428) );
  ANDN U9452 ( .B(n9485), .A(n9486), .Z(n10098) );
  XOR U9453 ( .A(n5529), .B(n10100), .Z(n10095) );
  XOR U9454 ( .A(n8303), .B(n2394), .Z(n10100) );
  XNOR U9455 ( .A(n10101), .B(n9419), .Z(n2394) );
  XOR U9456 ( .A(round_reg[1211]), .B(n9611), .Z(n9419) );
  ANDN U9457 ( .B(n10028), .A(n10093), .Z(n10101) );
  XNOR U9458 ( .A(round_reg[828]), .B(n10102), .Z(n10028) );
  XNOR U9459 ( .A(n10103), .B(n9423), .Z(n8303) );
  XOR U9460 ( .A(round_reg[1219]), .B(n9523), .Z(n9423) );
  ANDN U9461 ( .B(n9488), .A(n9489), .Z(n10103) );
  XNOR U9462 ( .A(round_reg[861]), .B(n9199), .Z(n9488) );
  XNOR U9463 ( .A(n10104), .B(n10026), .Z(n5529) );
  ANDN U9464 ( .B(n9493), .A(n9494), .Z(n10104) );
  XNOR U9465 ( .A(round_reg[932]), .B(n10105), .Z(n9493) );
  XNOR U9466 ( .A(n7519), .B(n2427), .Z(n3594) );
  XNOR U9467 ( .A(n9867), .B(n10106), .Z(n2427) );
  XOR U9468 ( .A(n10107), .B(n10108), .Z(n9867) );
  XNOR U9469 ( .A(n3434), .B(n5020), .Z(n10108) );
  XOR U9470 ( .A(n10109), .B(n7621), .Z(n5020) );
  ANDN U9471 ( .B(n7622), .A(n9808), .Z(n10109) );
  XOR U9472 ( .A(n10110), .B(n8657), .Z(n3434) );
  ANDN U9473 ( .B(n8658), .A(n9811), .Z(n10110) );
  XNOR U9474 ( .A(n2393), .B(n10111), .Z(n10107) );
  XOR U9475 ( .A(n7614), .B(n3935), .Z(n10111) );
  XOR U9476 ( .A(n10112), .B(n7628), .Z(n3935) );
  NOR U9477 ( .A(n7627), .B(n9799), .Z(n10112) );
  XNOR U9478 ( .A(n10113), .B(n10114), .Z(n7614) );
  AND U9479 ( .A(n9802), .B(n10115), .Z(n10113) );
  XOR U9480 ( .A(n10116), .B(n7631), .Z(n2393) );
  ANDN U9481 ( .B(n7632), .A(n10117), .Z(n10116) );
  XOR U9482 ( .A(n10118), .B(n9744), .Z(n7519) );
  ANDN U9483 ( .B(n9793), .A(n9792), .Z(n10118) );
  XOR U9484 ( .A(n10119), .B(n6179), .Z(out[1019]) );
  XNOR U9485 ( .A(n7940), .B(n2662), .Z(n6179) );
  XNOR U9486 ( .A(n6051), .B(n7981), .Z(n2662) );
  XNOR U9487 ( .A(n10120), .B(n10121), .Z(n7981) );
  XNOR U9488 ( .A(n10122), .B(n5407), .Z(n10121) );
  XNOR U9489 ( .A(n10123), .B(n8622), .Z(n5407) );
  ANDN U9490 ( .B(n7957), .A(n7955), .Z(n10123) );
  XOR U9491 ( .A(round_reg[529]), .B(n10124), .Z(n7957) );
  XOR U9492 ( .A(n7019), .B(n10125), .Z(n10120) );
  XNOR U9493 ( .A(n2223), .B(n3367), .Z(n10125) );
  XNOR U9494 ( .A(n10126), .B(n8610), .Z(n3367) );
  ANDN U9495 ( .B(n7942), .A(n7943), .Z(n10126) );
  XOR U9496 ( .A(round_reg[374]), .B(n9198), .Z(n7943) );
  XOR U9497 ( .A(n10127), .B(n8615), .Z(n2223) );
  ANDN U9498 ( .B(n7949), .A(n7947), .Z(n10127) );
  XOR U9499 ( .A(round_reg[425]), .B(n9552), .Z(n7949) );
  XNOR U9500 ( .A(n10128), .B(n8607), .Z(n7019) );
  ANDN U9501 ( .B(n7951), .A(n7952), .Z(n10128) );
  XNOR U9502 ( .A(round_reg[495]), .B(n10129), .Z(n7952) );
  XOR U9503 ( .A(n10130), .B(n10131), .Z(n6051) );
  XNOR U9504 ( .A(n5233), .B(n1861), .Z(n10131) );
  XOR U9505 ( .A(n10132), .B(n10133), .Z(n1861) );
  AND U9506 ( .A(n9286), .B(n7040), .Z(n10132) );
  XNOR U9507 ( .A(round_reg[1532]), .B(n9530), .Z(n7040) );
  XOR U9508 ( .A(n10134), .B(n10135), .Z(n5233) );
  ANDN U9509 ( .B(n9282), .A(n9283), .Z(n10134) );
  XNOR U9510 ( .A(round_reg[1314]), .B(n10136), .Z(n9283) );
  XNOR U9511 ( .A(n3622), .B(n10137), .Z(n10130) );
  XOR U9512 ( .A(n8044), .B(n4080), .Z(n10137) );
  XNOR U9513 ( .A(n10138), .B(n10139), .Z(n4080) );
  NOR U9514 ( .A(n9293), .B(n7026), .Z(n10138) );
  XNOR U9515 ( .A(round_reg[1377]), .B(n10140), .Z(n7026) );
  XNOR U9516 ( .A(n10141), .B(n10142), .Z(n8044) );
  AND U9517 ( .A(n7030), .B(n9289), .Z(n10141) );
  XNOR U9518 ( .A(round_reg[1597]), .B(n9906), .Z(n7030) );
  XNOR U9519 ( .A(n10143), .B(n10144), .Z(n3622) );
  ANDN U9520 ( .B(n7036), .A(n9291), .Z(n10143) );
  XOR U9521 ( .A(round_reg[1471]), .B(n9821), .Z(n7036) );
  IV U9522 ( .A(n9614), .Z(n9821) );
  XOR U9523 ( .A(n10145), .B(n10146), .Z(n7940) );
  ANDN U9524 ( .B(n10018), .A(n8617), .Z(n10145) );
  XOR U9525 ( .A(round_reg[252]), .B(n9530), .Z(n8617) );
  XNOR U9526 ( .A(n10147), .B(n10148), .Z(n9530) );
  ANDN U9527 ( .B(n5636), .A(n5637), .Z(n10119) );
  XOR U9528 ( .A(n9424), .B(n2036), .Z(n5637) );
  XNOR U9529 ( .A(n9297), .B(n8357), .Z(n2036) );
  XNOR U9530 ( .A(n10149), .B(n10150), .Z(n8357) );
  XOR U9531 ( .A(n5426), .B(n3810), .Z(n10150) );
  XOR U9532 ( .A(n10151), .B(n10152), .Z(n3810) );
  ANDN U9533 ( .B(n10153), .A(n9576), .Z(n10151) );
  XNOR U9534 ( .A(n10154), .B(n9503), .Z(n5426) );
  ANDN U9535 ( .B(n9504), .A(n10155), .Z(n10154) );
  XOR U9536 ( .A(n6278), .B(n10156), .Z(n10149) );
  XOR U9537 ( .A(n2274), .B(n4946), .Z(n10156) );
  XNOR U9538 ( .A(n10157), .B(n9507), .Z(n4946) );
  ANDN U9539 ( .B(n9508), .A(n9571), .Z(n10157) );
  XNOR U9540 ( .A(n10158), .B(n9517), .Z(n2274) );
  ANDN U9541 ( .B(n9518), .A(n9580), .Z(n10158) );
  XNOR U9542 ( .A(n10159), .B(n9513), .Z(n6278) );
  ANDN U9543 ( .B(n9514), .A(n9568), .Z(n10159) );
  XOR U9544 ( .A(n10160), .B(n10161), .Z(n9297) );
  XOR U9545 ( .A(n1970), .B(n9481), .Z(n10161) );
  XOR U9546 ( .A(n10162), .B(n10093), .Z(n9481) );
  XOR U9547 ( .A(round_reg[402]), .B(n9080), .Z(n10093) );
  ANDN U9548 ( .B(n9417), .A(n9418), .Z(n10162) );
  XNOR U9549 ( .A(round_reg[1575]), .B(n9818), .Z(n9418) );
  XOR U9550 ( .A(round_reg[25]), .B(n9934), .Z(n9417) );
  XNOR U9551 ( .A(n10163), .B(n9486), .Z(n1970) );
  XOR U9552 ( .A(round_reg[351]), .B(n9554), .Z(n9486) );
  AND U9553 ( .A(n9429), .B(n9427), .Z(n10163) );
  XNOR U9554 ( .A(round_reg[277]), .B(n10164), .Z(n9427) );
  XNOR U9555 ( .A(round_reg[1510]), .B(n10045), .Z(n9429) );
  XOR U9556 ( .A(n3718), .B(n10165), .Z(n10160) );
  XOR U9557 ( .A(n5098), .B(n4150), .Z(n10165) );
  XNOR U9558 ( .A(n10166), .B(n9494), .Z(n4150) );
  XOR U9559 ( .A(round_reg[570]), .B(n9685), .Z(n9494) );
  ANDN U9560 ( .B(n9495), .A(n10025), .Z(n10166) );
  XNOR U9561 ( .A(n10167), .B(n9489), .Z(n5098) );
  XOR U9562 ( .A(round_reg[472]), .B(n9753), .Z(n9489) );
  ANDN U9563 ( .B(n9421), .A(n9422), .Z(n10167) );
  XOR U9564 ( .A(round_reg[1292]), .B(n10168), .Z(n9422) );
  XOR U9565 ( .A(round_reg[111]), .B(n9375), .Z(n9421) );
  XNOR U9566 ( .A(n10169), .B(n9498), .Z(n3718) );
  XOR U9567 ( .A(round_reg[638]), .B(n9838), .Z(n9498) );
  ANDN U9568 ( .B(n9431), .A(n9432), .Z(n10169) );
  XOR U9569 ( .A(round_reg[1449]), .B(n10170), .Z(n9432) );
  XOR U9570 ( .A(round_reg[229]), .B(n10171), .Z(n9431) );
  XOR U9571 ( .A(n10172), .B(n9495), .Z(n9424) );
  XNOR U9572 ( .A(round_reg[170]), .B(n10173), .Z(n9495) );
  ANDN U9573 ( .B(n10025), .A(n10026), .Z(n10172) );
  XOR U9574 ( .A(round_reg[979]), .B(n10174), .Z(n10026) );
  XOR U9575 ( .A(round_reg[1355]), .B(n9692), .Z(n10025) );
  XOR U9576 ( .A(n10175), .B(n1695), .Z(n5636) );
  XNOR U9577 ( .A(n8778), .B(n6314), .Z(n1695) );
  XNOR U9578 ( .A(n10176), .B(n10177), .Z(n6314) );
  XNOR U9579 ( .A(n5395), .B(n3608), .Z(n10177) );
  XOR U9580 ( .A(n10178), .B(n10179), .Z(n3608) );
  ANDN U9581 ( .B(n7903), .A(n10180), .Z(n10178) );
  XNOR U9582 ( .A(n10181), .B(n10182), .Z(n5395) );
  AND U9583 ( .A(n7893), .B(n10183), .Z(n10181) );
  XNOR U9584 ( .A(n10184), .B(n10185), .Z(n10176) );
  XOR U9585 ( .A(n2072), .B(n5313), .Z(n10185) );
  XNOR U9586 ( .A(n10186), .B(n10187), .Z(n5313) );
  ANDN U9587 ( .B(n7897), .A(n10188), .Z(n10186) );
  XNOR U9588 ( .A(n10189), .B(n10190), .Z(n2072) );
  ANDN U9589 ( .B(n8898), .A(n10191), .Z(n10189) );
  XOR U9590 ( .A(n10192), .B(n10193), .Z(n8778) );
  XOR U9591 ( .A(n5034), .B(n7821), .Z(n10193) );
  XNOR U9592 ( .A(n10194), .B(n7827), .Z(n7821) );
  AND U9593 ( .A(n10057), .B(n7828), .Z(n10194) );
  XOR U9594 ( .A(n10195), .B(n7831), .Z(n5034) );
  ANDN U9595 ( .B(n7832), .A(n10062), .Z(n10195) );
  XOR U9596 ( .A(n2417), .B(n10196), .Z(n10192) );
  XOR U9597 ( .A(n3440), .B(n3944), .Z(n10196) );
  XOR U9598 ( .A(n10197), .B(n7838), .Z(n3944) );
  NOR U9599 ( .A(n7837), .B(n10053), .Z(n10197) );
  XOR U9600 ( .A(n10198), .B(n8839), .Z(n3440) );
  ANDN U9601 ( .B(n8840), .A(n10065), .Z(n10198) );
  XOR U9602 ( .A(n10199), .B(n10200), .Z(n2417) );
  AND U9603 ( .A(n10201), .B(n7842), .Z(n10199) );
  XOR U9604 ( .A(n10202), .B(n6184), .Z(out[1018]) );
  XOR U9605 ( .A(n10203), .B(n2669), .Z(n6184) );
  XNOR U9606 ( .A(n6056), .B(n8602), .Z(n2669) );
  XNOR U9607 ( .A(n10204), .B(n10205), .Z(n8602) );
  XNOR U9608 ( .A(n5617), .B(n5411), .Z(n10205) );
  XNOR U9609 ( .A(n10206), .B(n7028), .Z(n5411) );
  XOR U9610 ( .A(round_reg[1001]), .B(n10207), .Z(n7028) );
  ANDN U9611 ( .B(n10139), .A(n7027), .Z(n10206) );
  XOR U9612 ( .A(n10208), .B(n7038), .Z(n5617) );
  XNOR U9613 ( .A(round_reg[1030]), .B(n10012), .Z(n7038) );
  ANDN U9614 ( .B(n10144), .A(n7037), .Z(n10208) );
  XOR U9615 ( .A(n7021), .B(n10209), .Z(n10204) );
  XNOR U9616 ( .A(n2230), .B(n3370), .Z(n10209) );
  XNOR U9617 ( .A(n10210), .B(n7041), .Z(n3370) );
  XOR U9618 ( .A(round_reg[1143]), .B(n10211), .Z(n7041) );
  AND U9619 ( .A(n7042), .B(n10212), .Z(n10210) );
  XNOR U9620 ( .A(n10213), .B(n7032), .Z(n2230) );
  XNOR U9621 ( .A(round_reg[1169]), .B(n10214), .Z(n7032) );
  ANDN U9622 ( .B(n10142), .A(n7031), .Z(n10213) );
  XNOR U9623 ( .A(n10215), .B(n9284), .Z(n7021) );
  XOR U9624 ( .A(round_reg[1241]), .B(n10216), .Z(n9284) );
  ANDN U9625 ( .B(n9295), .A(n10135), .Z(n10215) );
  XOR U9626 ( .A(n10217), .B(n10218), .Z(n6056) );
  XNOR U9627 ( .A(n5237), .B(n1869), .Z(n10218) );
  XOR U9628 ( .A(n10219), .B(n8101), .Z(n1869) );
  AND U9629 ( .A(n7063), .B(n10085), .Z(n10219) );
  XNOR U9630 ( .A(round_reg[298]), .B(n10220), .Z(n10085) );
  XNOR U9631 ( .A(round_reg[1531]), .B(n9611), .Z(n7063) );
  XOR U9632 ( .A(n10221), .B(n8109), .Z(n5237) );
  ANDN U9633 ( .B(n8110), .A(n10082), .Z(n10221) );
  XNOR U9634 ( .A(round_reg[1313]), .B(n10222), .Z(n10082) );
  XOR U9635 ( .A(round_reg[68]), .B(n10223), .Z(n8110) );
  XNOR U9636 ( .A(n3626), .B(n10224), .Z(n10217) );
  XOR U9637 ( .A(n8095), .B(n4084), .Z(n10224) );
  XNOR U9638 ( .A(n10225), .B(n8113), .Z(n4084) );
  NOR U9639 ( .A(n8112), .B(n7049), .Z(n10225) );
  XNOR U9640 ( .A(round_reg[1376]), .B(n10226), .Z(n7049) );
  XNOR U9641 ( .A(round_reg[191]), .B(n9614), .Z(n8112) );
  XNOR U9642 ( .A(n10227), .B(n8106), .Z(n8095) );
  AND U9643 ( .A(n7053), .B(n8105), .Z(n10227) );
  XNOR U9644 ( .A(round_reg[46]), .B(n9205), .Z(n8105) );
  XNOR U9645 ( .A(round_reg[1596]), .B(n9993), .Z(n7053) );
  XNOR U9646 ( .A(n10228), .B(n10229), .Z(n3626) );
  ANDN U9647 ( .B(n7059), .A(n10089), .Z(n10228) );
  XOR U9648 ( .A(round_reg[1470]), .B(n9891), .Z(n7059) );
  IV U9649 ( .A(n9688), .Z(n9891) );
  NOR U9650 ( .A(n5641), .B(n5640), .Z(n10202) );
  XOR U9651 ( .A(n10230), .B(n1700), .Z(n5640) );
  XNOR U9652 ( .A(n8836), .B(n6318), .Z(n1700) );
  XNOR U9653 ( .A(n10231), .B(n10232), .Z(n6318) );
  XOR U9654 ( .A(n5400), .B(n3612), .Z(n10232) );
  XOR U9655 ( .A(n10233), .B(n10234), .Z(n3612) );
  AND U9656 ( .A(n10235), .B(n7973), .Z(n10233) );
  XNOR U9657 ( .A(n10236), .B(n10237), .Z(n5400) );
  AND U9658 ( .A(n10238), .B(n7963), .Z(n10236) );
  XNOR U9659 ( .A(n10239), .B(n10240), .Z(n10231) );
  XOR U9660 ( .A(n2075), .B(n5367), .Z(n10240) );
  XNOR U9661 ( .A(n10241), .B(n10242), .Z(n5367) );
  ANDN U9662 ( .B(n7967), .A(n10243), .Z(n10241) );
  XNOR U9663 ( .A(n10244), .B(n10245), .Z(n2075) );
  ANDN U9664 ( .B(n8958), .A(n10246), .Z(n10244) );
  XOR U9665 ( .A(n10247), .B(n10248), .Z(n8836) );
  XNOR U9666 ( .A(n3446), .B(n5039), .Z(n10248) );
  XOR U9667 ( .A(n10249), .B(n7898), .Z(n5039) );
  ANDN U9668 ( .B(n7899), .A(n10187), .Z(n10249) );
  XOR U9669 ( .A(n10250), .B(n8899), .Z(n3446) );
  ANDN U9670 ( .B(n8900), .A(n10190), .Z(n10250) );
  XNOR U9671 ( .A(n3947), .B(n10251), .Z(n10247) );
  XOR U9672 ( .A(n7888), .B(n2425), .Z(n10251) );
  XOR U9673 ( .A(n10252), .B(n7908), .Z(n2425) );
  AND U9674 ( .A(n10253), .B(n7909), .Z(n10252) );
  XNOR U9675 ( .A(n10254), .B(n7894), .Z(n7888) );
  AND U9676 ( .A(n10182), .B(n7895), .Z(n10254) );
  XOR U9677 ( .A(n10255), .B(n7905), .Z(n3947) );
  NOR U9678 ( .A(n7904), .B(n10179), .Z(n10255) );
  XOR U9679 ( .A(n9509), .B(n2040), .Z(n5641) );
  XNOR U9680 ( .A(n10094), .B(n8649), .Z(n2040) );
  XNOR U9681 ( .A(n10256), .B(n10257), .Z(n8649) );
  XOR U9682 ( .A(n5430), .B(n3816), .Z(n10257) );
  XOR U9683 ( .A(n10258), .B(n10259), .Z(n3816) );
  AND U9684 ( .A(n7417), .B(n7416), .Z(n10258) );
  XOR U9685 ( .A(round_reg[930]), .B(n10260), .Z(n7417) );
  XNOR U9686 ( .A(n10261), .B(n9586), .Z(n5430) );
  AND U9687 ( .A(n7413), .B(n7412), .Z(n10261) );
  XNOR U9688 ( .A(round_reg[1209]), .B(n10262), .Z(n7412) );
  XOR U9689 ( .A(round_reg[826]), .B(n9918), .Z(n7413) );
  XNOR U9690 ( .A(n6283), .B(n10263), .Z(n10256) );
  XOR U9691 ( .A(n2281), .B(n4981), .Z(n10263) );
  XNOR U9692 ( .A(n10264), .B(n9589), .Z(n4981) );
  ANDN U9693 ( .B(n8408), .A(n8409), .Z(n10264) );
  XNOR U9694 ( .A(round_reg[859]), .B(n9363), .Z(n8409) );
  IV U9695 ( .A(n10265), .Z(n9363) );
  XOR U9696 ( .A(round_reg[1217]), .B(n9676), .Z(n8408) );
  XNOR U9697 ( .A(n10266), .B(n9597), .Z(n2281) );
  AND U9698 ( .A(n8652), .B(n8651), .Z(n10266) );
  XOR U9699 ( .A(round_reg[1070]), .B(n9094), .Z(n8651) );
  XOR U9700 ( .A(round_reg[702]), .B(n9536), .Z(n8652) );
  XNOR U9701 ( .A(n10267), .B(n9594), .Z(n6283) );
  ANDN U9702 ( .B(n7406), .A(n7407), .Z(n10267) );
  XOR U9703 ( .A(round_reg[716]), .B(n9621), .Z(n7407) );
  XOR U9704 ( .A(round_reg[1119]), .B(n9192), .Z(n7406) );
  XOR U9705 ( .A(n10268), .B(n10269), .Z(n10094) );
  XNOR U9706 ( .A(n1657), .B(n9564), .Z(n10269) );
  XOR U9707 ( .A(n10270), .B(n10271), .Z(n9564) );
  ANDN U9708 ( .B(n9502), .A(n9503), .Z(n10270) );
  XOR U9709 ( .A(round_reg[1574]), .B(n9889), .Z(n9503) );
  XNOR U9710 ( .A(n10272), .B(n9569), .Z(n1657) );
  ANDN U9711 ( .B(n9512), .A(n9513), .Z(n10272) );
  XOR U9712 ( .A(round_reg[1509]), .B(n10171), .Z(n9513) );
  XNOR U9713 ( .A(round_reg[276]), .B(n10273), .Z(n9512) );
  XOR U9714 ( .A(n3722), .B(n10274), .Z(n10268) );
  XOR U9715 ( .A(n5100), .B(n4153), .Z(n10274) );
  XNOR U9716 ( .A(n10275), .B(n9578), .Z(n4153) );
  NOR U9717 ( .A(n9577), .B(n10152), .Z(n10275) );
  XNOR U9718 ( .A(n10276), .B(n9572), .Z(n5100) );
  XOR U9719 ( .A(round_reg[1291]), .B(n10277), .Z(n9507) );
  XNOR U9720 ( .A(round_reg[110]), .B(n9094), .Z(n9506) );
  XNOR U9721 ( .A(n10278), .B(n10279), .Z(n9094) );
  XNOR U9722 ( .A(n10280), .B(n9581), .Z(n3722) );
  ANDN U9723 ( .B(n9516), .A(n9517), .Z(n10280) );
  XOR U9724 ( .A(round_reg[1448]), .B(n10281), .Z(n9517) );
  XOR U9725 ( .A(round_reg[228]), .B(n10282), .Z(n9516) );
  XNOR U9726 ( .A(n10283), .B(n9577), .Z(n9509) );
  XOR U9727 ( .A(round_reg[169]), .B(n10284), .Z(n9577) );
  ANDN U9728 ( .B(n10152), .A(n10153), .Z(n10283) );
  XOR U9729 ( .A(round_reg[1354]), .B(n9767), .Z(n10152) );
  XOR U9730 ( .A(n10285), .B(n6189), .Z(out[1017]) );
  XOR U9731 ( .A(n8099), .B(n2676), .Z(n6189) );
  XNOR U9732 ( .A(n6061), .B(n9278), .Z(n2676) );
  XNOR U9733 ( .A(n10286), .B(n10287), .Z(n9278) );
  XNOR U9734 ( .A(n5662), .B(n5415), .Z(n10287) );
  XNOR U9735 ( .A(n10288), .B(n7051), .Z(n5415) );
  XOR U9736 ( .A(round_reg[1000]), .B(n10289), .Z(n7051) );
  ANDN U9737 ( .B(n8113), .A(n7050), .Z(n10288) );
  XNOR U9738 ( .A(round_reg[953]), .B(n10290), .Z(n7050) );
  XOR U9739 ( .A(round_reg[527]), .B(n10291), .Z(n8113) );
  XNOR U9740 ( .A(n10292), .B(n7061), .Z(n5662) );
  XOR U9741 ( .A(round_reg[1029]), .B(n10293), .Z(n7061) );
  ANDN U9742 ( .B(n10229), .A(n7060), .Z(n10292) );
  XOR U9743 ( .A(n7044), .B(n10294), .Z(n10286) );
  XNOR U9744 ( .A(n2237), .B(n3373), .Z(n10294) );
  XNOR U9745 ( .A(n10295), .B(n7064), .Z(n3373) );
  XOR U9746 ( .A(round_reg[1142]), .B(n10296), .Z(n7064) );
  ANDN U9747 ( .B(n7065), .A(n8101), .Z(n10295) );
  XOR U9748 ( .A(round_reg[372]), .B(n10297), .Z(n8101) );
  XOR U9749 ( .A(round_reg[739]), .B(n9928), .Z(n7065) );
  XNOR U9750 ( .A(n10298), .B(n7055), .Z(n2237) );
  XNOR U9751 ( .A(round_reg[1168]), .B(n10299), .Z(n7055) );
  ANDN U9752 ( .B(n8106), .A(n7054), .Z(n10298) );
  XNOR U9753 ( .A(round_reg[785]), .B(n10300), .Z(n7054) );
  XOR U9754 ( .A(round_reg[423]), .B(n9705), .Z(n8106) );
  IV U9755 ( .A(n9919), .Z(n9705) );
  XNOR U9756 ( .A(n10301), .B(n10083), .Z(n7044) );
  XOR U9757 ( .A(round_reg[1240]), .B(n10302), .Z(n10083) );
  ANDN U9758 ( .B(n8108), .A(n8109), .Z(n10301) );
  XNOR U9759 ( .A(round_reg[493]), .B(n10303), .Z(n8109) );
  XOR U9760 ( .A(round_reg[882]), .B(n10304), .Z(n8108) );
  XOR U9761 ( .A(n10305), .B(n10306), .Z(n6061) );
  XNOR U9762 ( .A(n5239), .B(n1873), .Z(n10306) );
  XNOR U9763 ( .A(n10307), .B(n8149), .Z(n1873) );
  ANDN U9764 ( .B(n7086), .A(n8148), .Z(n10307) );
  XOR U9765 ( .A(n10308), .B(n8157), .Z(n5239) );
  ANDN U9766 ( .B(n10309), .A(n8156), .Z(n10308) );
  XNOR U9767 ( .A(n3630), .B(n10310), .Z(n10305) );
  XOR U9768 ( .A(n8143), .B(n4088), .Z(n10310) );
  XNOR U9769 ( .A(n10311), .B(n8160), .Z(n4088) );
  NOR U9770 ( .A(n7072), .B(n8159), .Z(n10311) );
  XNOR U9771 ( .A(n10312), .B(n8153), .Z(n8143) );
  AND U9772 ( .A(n8152), .B(n7076), .Z(n10312) );
  XNOR U9773 ( .A(n10313), .B(n10314), .Z(n3630) );
  ANDN U9774 ( .B(n7082), .A(n10315), .Z(n10313) );
  XOR U9775 ( .A(n10316), .B(n7060), .Z(n8099) );
  XNOR U9776 ( .A(round_reg[661]), .B(n9987), .Z(n7060) );
  XOR U9777 ( .A(round_reg[595]), .B(n10317), .Z(n10229) );
  XNOR U9778 ( .A(round_reg[250]), .B(n9685), .Z(n10089) );
  NOR U9779 ( .A(n5646), .B(n5644), .Z(n10285) );
  XOR U9780 ( .A(n10318), .B(n1705), .Z(n5644) );
  XNOR U9781 ( .A(n8895), .B(n6326), .Z(n1705) );
  XNOR U9782 ( .A(n10319), .B(n10320), .Z(n6326) );
  XNOR U9783 ( .A(n5405), .B(n3616), .Z(n10320) );
  XOR U9784 ( .A(n10321), .B(n10322), .Z(n3616) );
  NOR U9785 ( .A(n8062), .B(n10323), .Z(n10321) );
  XNOR U9786 ( .A(n10324), .B(n10325), .Z(n5405) );
  ANDN U9787 ( .B(n10326), .A(n8052), .Z(n10324) );
  XNOR U9788 ( .A(n10327), .B(n10328), .Z(n10319) );
  XOR U9789 ( .A(n2079), .B(n5417), .Z(n10328) );
  XNOR U9790 ( .A(n10329), .B(n10330), .Z(n5417) );
  ANDN U9791 ( .B(n8056), .A(n10331), .Z(n10329) );
  XNOR U9792 ( .A(n10332), .B(n10333), .Z(n2079) );
  NOR U9793 ( .A(n9017), .B(n10334), .Z(n10332) );
  XOR U9794 ( .A(n10335), .B(n10336), .Z(n8895) );
  XNOR U9795 ( .A(n3448), .B(n5044), .Z(n10336) );
  XOR U9796 ( .A(n10337), .B(n7968), .Z(n5044) );
  ANDN U9797 ( .B(n7969), .A(n10242), .Z(n10337) );
  XOR U9798 ( .A(n10338), .B(n8959), .Z(n3448) );
  ANDN U9799 ( .B(n8960), .A(n10245), .Z(n10338) );
  XNOR U9800 ( .A(n3962), .B(n10339), .Z(n10335) );
  XOR U9801 ( .A(n7958), .B(n2432), .Z(n10339) );
  XOR U9802 ( .A(n10340), .B(n7978), .Z(n2432) );
  AND U9803 ( .A(n10341), .B(n7979), .Z(n10340) );
  XOR U9804 ( .A(n10342), .B(n10343), .Z(n7958) );
  ANDN U9805 ( .B(n7965), .A(n10237), .Z(n10342) );
  XOR U9806 ( .A(n10344), .B(n7975), .Z(n3962) );
  NOR U9807 ( .A(n7974), .B(n10234), .Z(n10344) );
  XOR U9808 ( .A(n9590), .B(n2048), .Z(n5646) );
  XNOR U9809 ( .A(n10345), .B(n9322), .Z(n2048) );
  XNOR U9810 ( .A(n10346), .B(n10347), .Z(n9322) );
  XOR U9811 ( .A(n5435), .B(n3820), .Z(n10347) );
  XOR U9812 ( .A(n10348), .B(n10349), .Z(n3820) );
  ANDN U9813 ( .B(n7487), .A(n7488), .Z(n10348) );
  XOR U9814 ( .A(round_reg[929]), .B(n9219), .Z(n7488) );
  XNOR U9815 ( .A(n10350), .B(n9660), .Z(n5435) );
  ANDN U9816 ( .B(n7483), .A(n7484), .Z(n10350) );
  XNOR U9817 ( .A(round_reg[825]), .B(n9370), .Z(n7484) );
  XOR U9818 ( .A(round_reg[1208]), .B(n10351), .Z(n7483) );
  XOR U9819 ( .A(n6288), .B(n10352), .Z(n10346) );
  XOR U9820 ( .A(n2288), .B(n5028), .Z(n10352) );
  XNOR U9821 ( .A(n10353), .B(n9663), .Z(n5028) );
  ANDN U9822 ( .B(n8461), .A(n8462), .Z(n10353) );
  XNOR U9823 ( .A(round_reg[858]), .B(n9438), .Z(n8462) );
  XOR U9824 ( .A(round_reg[1216]), .B(n9749), .Z(n8461) );
  XNOR U9825 ( .A(n10354), .B(n9671), .Z(n2288) );
  ANDN U9826 ( .B(n9326), .A(n9324), .Z(n10354) );
  XNOR U9827 ( .A(round_reg[1069]), .B(n9535), .Z(n9324) );
  XOR U9828 ( .A(round_reg[701]), .B(n9615), .Z(n9326) );
  XNOR U9829 ( .A(n10355), .B(n9668), .Z(n6288) );
  ANDN U9830 ( .B(n7477), .A(n7478), .Z(n10355) );
  XNOR U9831 ( .A(round_reg[715]), .B(n10356), .Z(n7478) );
  XOR U9832 ( .A(round_reg[1118]), .B(n10357), .Z(n7477) );
  XOR U9833 ( .A(n10358), .B(n9655), .Z(n9590) );
  ANDN U9834 ( .B(n10259), .A(n7416), .Z(n10358) );
  XOR U9835 ( .A(round_reg[977]), .B(n10359), .Z(n7416) );
  XOR U9836 ( .A(n10360), .B(n6194), .Z(out[1016]) );
  XOR U9837 ( .A(n8146), .B(n2683), .Z(n6194) );
  XNOR U9838 ( .A(n6066), .B(n10078), .Z(n2683) );
  XNOR U9839 ( .A(n10361), .B(n10362), .Z(n10078) );
  XNOR U9840 ( .A(n5708), .B(n5423), .Z(n10362) );
  XNOR U9841 ( .A(n10363), .B(n7074), .Z(n5423) );
  ANDN U9842 ( .B(n8160), .A(n7073), .Z(n10363) );
  XNOR U9843 ( .A(round_reg[952]), .B(n9092), .Z(n7073) );
  XOR U9844 ( .A(round_reg[526]), .B(n10364), .Z(n8160) );
  XOR U9845 ( .A(n10365), .B(n10366), .Z(n5708) );
  ANDN U9846 ( .B(n10314), .A(n7083), .Z(n10365) );
  XOR U9847 ( .A(n7067), .B(n10367), .Z(n10361) );
  XNOR U9848 ( .A(n2244), .B(n3376), .Z(n10367) );
  XNOR U9849 ( .A(n10368), .B(n7087), .Z(n3376) );
  AND U9850 ( .A(n8149), .B(n7088), .Z(n10368) );
  XNOR U9851 ( .A(round_reg[738]), .B(n10369), .Z(n7088) );
  XNOR U9852 ( .A(round_reg[371]), .B(n10370), .Z(n8149) );
  XNOR U9853 ( .A(n10371), .B(n7078), .Z(n2244) );
  ANDN U9854 ( .B(n8153), .A(n7077), .Z(n10371) );
  XNOR U9855 ( .A(round_reg[784]), .B(n10372), .Z(n7077) );
  XOR U9856 ( .A(round_reg[422]), .B(n9776), .Z(n8153) );
  XNOR U9857 ( .A(n10373), .B(n10374), .Z(n7067) );
  ANDN U9858 ( .B(n8155), .A(n8157), .Z(n10373) );
  XNOR U9859 ( .A(round_reg[492]), .B(n9986), .Z(n8157) );
  XOR U9860 ( .A(n10375), .B(n10376), .Z(n6066) );
  XNOR U9861 ( .A(n5247), .B(n1877), .Z(n10376) );
  XNOR U9862 ( .A(n10377), .B(n8205), .Z(n1877) );
  NOR U9863 ( .A(n7112), .B(n8166), .Z(n10377) );
  XNOR U9864 ( .A(round_reg[296]), .B(n10036), .Z(n8166) );
  XNOR U9865 ( .A(round_reg[1529]), .B(n10262), .Z(n7112) );
  IV U9866 ( .A(n9758), .Z(n10262) );
  XOR U9867 ( .A(n10378), .B(n8211), .Z(n5247) );
  ANDN U9868 ( .B(n8164), .A(n7108), .Z(n10378) );
  XOR U9869 ( .A(round_reg[66]), .B(n10379), .Z(n8164) );
  XNOR U9870 ( .A(n3634), .B(n10380), .Z(n10375) );
  XOR U9871 ( .A(n8200), .B(n4092), .Z(n10380) );
  XNOR U9872 ( .A(n10381), .B(n8213), .Z(n4092) );
  ANDN U9873 ( .B(n8173), .A(n7095), .Z(n10381) );
  XNOR U9874 ( .A(round_reg[1374]), .B(n10382), .Z(n7095) );
  XOR U9875 ( .A(round_reg[189]), .B(n9761), .Z(n8173) );
  XNOR U9876 ( .A(n10383), .B(n8208), .Z(n8200) );
  ANDN U9877 ( .B(n8209), .A(n7099), .Z(n10383) );
  XOR U9878 ( .A(round_reg[1594]), .B(n10384), .Z(n7099) );
  XNOR U9879 ( .A(round_reg[44]), .B(n9379), .Z(n8209) );
  XNOR U9880 ( .A(n10385), .B(n10386), .Z(n3634) );
  ANDN U9881 ( .B(n8171), .A(n7104), .Z(n10385) );
  XNOR U9882 ( .A(round_reg[1468]), .B(n10102), .Z(n7104) );
  XOR U9883 ( .A(n10387), .B(n7083), .Z(n8146) );
  XNOR U9884 ( .A(round_reg[660]), .B(n10048), .Z(n7083) );
  XOR U9885 ( .A(round_reg[594]), .B(n10388), .Z(n10314) );
  NOR U9886 ( .A(n5649), .B(n5648), .Z(n10360) );
  XOR U9887 ( .A(n10389), .B(n1710), .Z(n5648) );
  XNOR U9888 ( .A(n8955), .B(n6330), .Z(n1710) );
  XNOR U9889 ( .A(n10390), .B(n10391), .Z(n6330) );
  XNOR U9890 ( .A(n5409), .B(n3620), .Z(n10391) );
  XOR U9891 ( .A(n10392), .B(n10393), .Z(n3620) );
  NOR U9892 ( .A(n8129), .B(n10394), .Z(n10392) );
  XNOR U9893 ( .A(n10395), .B(n10396), .Z(n5409) );
  AND U9894 ( .A(n8119), .B(n10397), .Z(n10395) );
  XNOR U9895 ( .A(n10398), .B(n10399), .Z(n10390) );
  XOR U9896 ( .A(n2086), .B(n5467), .Z(n10399) );
  XNOR U9897 ( .A(n10400), .B(n10401), .Z(n5467) );
  ANDN U9898 ( .B(n8123), .A(n10402), .Z(n10400) );
  XNOR U9899 ( .A(n10403), .B(n10404), .Z(n2086) );
  ANDN U9900 ( .B(n10405), .A(n9071), .Z(n10403) );
  XOR U9901 ( .A(n10406), .B(n10407), .Z(n8955) );
  XNOR U9902 ( .A(n3450), .B(n5049), .Z(n10407) );
  XOR U9903 ( .A(n10408), .B(n8057), .Z(n5049) );
  ANDN U9904 ( .B(n8058), .A(n10330), .Z(n10408) );
  XOR U9905 ( .A(n10409), .B(n9019), .Z(n3450) );
  NOR U9906 ( .A(n9018), .B(n10333), .Z(n10409) );
  XNOR U9907 ( .A(n3995), .B(n10410), .Z(n10406) );
  XOR U9908 ( .A(n8047), .B(n2441), .Z(n10410) );
  XOR U9909 ( .A(n10411), .B(n8067), .Z(n2441) );
  AND U9910 ( .A(n10412), .B(n8068), .Z(n10411) );
  XOR U9911 ( .A(n10413), .B(n10414), .Z(n8047) );
  AND U9912 ( .A(n10325), .B(n8054), .Z(n10413) );
  XOR U9913 ( .A(n10415), .B(n8064), .Z(n3995) );
  NOR U9914 ( .A(n8063), .B(n10322), .Z(n10415) );
  XOR U9915 ( .A(n9664), .B(n2052), .Z(n5649) );
  XNOR U9916 ( .A(n7401), .B(n10106), .Z(n2052) );
  XNOR U9917 ( .A(n10416), .B(n10417), .Z(n10106) );
  XOR U9918 ( .A(n5439), .B(n3824), .Z(n10417) );
  XOR U9919 ( .A(n10418), .B(n10419), .Z(n3824) );
  ANDN U9920 ( .B(n7531), .A(n7532), .Z(n10418) );
  XNOR U9921 ( .A(round_reg[928]), .B(n10420), .Z(n7532) );
  XNOR U9922 ( .A(n10421), .B(n9733), .Z(n5439) );
  ANDN U9923 ( .B(n7527), .A(n7528), .Z(n10421) );
  XNOR U9924 ( .A(round_reg[824]), .B(n9450), .Z(n7528) );
  IV U9925 ( .A(n10422), .Z(n9450) );
  XOR U9926 ( .A(round_reg[1207]), .B(n9844), .Z(n7527) );
  XNOR U9927 ( .A(n6292), .B(n10423), .Z(n10416) );
  XOR U9928 ( .A(n2295), .B(n5079), .Z(n10423) );
  XNOR U9929 ( .A(n10424), .B(n9736), .Z(n5079) );
  ANDN U9930 ( .B(n8534), .A(n8535), .Z(n10424) );
  XNOR U9931 ( .A(round_reg[857]), .B(n9524), .Z(n8535) );
  XOR U9932 ( .A(round_reg[1279]), .B(n9930), .Z(n8534) );
  XNOR U9933 ( .A(n10425), .B(n9745), .Z(n2295) );
  ANDN U9934 ( .B(n9792), .A(n9744), .Z(n10425) );
  XNOR U9935 ( .A(round_reg[1068]), .B(n9616), .Z(n9744) );
  XOR U9936 ( .A(round_reg[700]), .B(n9088), .Z(n9792) );
  XNOR U9937 ( .A(n10426), .B(n9741), .Z(n6292) );
  ANDN U9938 ( .B(n7521), .A(n7522), .Z(n10426) );
  XNOR U9939 ( .A(round_reg[714]), .B(n10427), .Z(n7522) );
  XNOR U9940 ( .A(round_reg[1117]), .B(n9367), .Z(n7521) );
  XOR U9941 ( .A(n10428), .B(n10429), .Z(n7401) );
  XOR U9942 ( .A(n1670), .B(n9717), .Z(n10429) );
  XOR U9943 ( .A(n10430), .B(n7485), .Z(n9717) );
  XOR U9944 ( .A(round_reg[399]), .B(n9380), .Z(n7485) );
  ANDN U9945 ( .B(n9659), .A(n9660), .Z(n10430) );
  XOR U9946 ( .A(round_reg[1572]), .B(n10431), .Z(n9660) );
  XOR U9947 ( .A(round_reg[22]), .B(n9901), .Z(n9659) );
  XNOR U9948 ( .A(n10432), .B(n7479), .Z(n1670) );
  XOR U9949 ( .A(round_reg[348]), .B(n9778), .Z(n7479) );
  NOR U9950 ( .A(n9667), .B(n9668), .Z(n10432) );
  XOR U9951 ( .A(round_reg[1507]), .B(n10433), .Z(n9668) );
  XOR U9952 ( .A(round_reg[274]), .B(n10388), .Z(n9667) );
  XOR U9953 ( .A(n3732), .B(n10434), .Z(n10428) );
  XOR U9954 ( .A(n5104), .B(n4160), .Z(n10434) );
  XNOR U9955 ( .A(n10435), .B(n7489), .Z(n4160) );
  XNOR U9956 ( .A(round_reg[567]), .B(n10436), .Z(n7489) );
  NOR U9957 ( .A(n9728), .B(n10349), .Z(n10435) );
  XNOR U9958 ( .A(n10437), .B(n8463), .Z(n5104) );
  XOR U9959 ( .A(round_reg[469]), .B(n9910), .Z(n8463) );
  ANDN U9960 ( .B(n9662), .A(n9663), .Z(n10437) );
  XNOR U9961 ( .A(round_reg[1289]), .B(n10438), .Z(n9663) );
  XOR U9962 ( .A(round_reg[108]), .B(n9616), .Z(n9662) );
  XOR U9963 ( .A(n10439), .B(n9325), .Z(n3732) );
  IV U9964 ( .A(n9726), .Z(n9325) );
  XNOR U9965 ( .A(round_reg[635]), .B(n10440), .Z(n9726) );
  ANDN U9966 ( .B(n9670), .A(n9671), .Z(n10439) );
  XOR U9967 ( .A(round_reg[1446]), .B(n10441), .Z(n9671) );
  XOR U9968 ( .A(round_reg[226]), .B(n10442), .Z(n9670) );
  XNOR U9969 ( .A(n10443), .B(n9728), .Z(n9664) );
  XOR U9970 ( .A(round_reg[167]), .B(n10444), .Z(n9728) );
  ANDN U9971 ( .B(n10349), .A(n7487), .Z(n10443) );
  XOR U9972 ( .A(round_reg[976]), .B(n10445), .Z(n7487) );
  XOR U9973 ( .A(round_reg[1352]), .B(n9852), .Z(n10349) );
  XOR U9974 ( .A(n10446), .B(n6199), .Z(out[1015]) );
  XOR U9975 ( .A(n8203), .B(n2690), .Z(n6199) );
  XNOR U9976 ( .A(n6071), .B(n10447), .Z(n2690) );
  XOR U9977 ( .A(n10448), .B(n10449), .Z(n6071) );
  XNOR U9978 ( .A(n5249), .B(n1881), .Z(n10449) );
  XNOR U9979 ( .A(n10450), .B(n8272), .Z(n1881) );
  ANDN U9980 ( .B(n7169), .A(n8219), .Z(n10450) );
  XOR U9981 ( .A(round_reg[295]), .B(n9818), .Z(n8219) );
  XOR U9982 ( .A(round_reg[1528]), .B(n10451), .Z(n7169) );
  XNOR U9983 ( .A(n10452), .B(n8277), .Z(n5249) );
  ANDN U9984 ( .B(n8217), .A(n7165), .Z(n10452) );
  XNOR U9985 ( .A(round_reg[1310]), .B(n10453), .Z(n7165) );
  XOR U9986 ( .A(round_reg[65]), .B(n10454), .Z(n8217) );
  XOR U9987 ( .A(n3643), .B(n10455), .Z(n10448) );
  XNOR U9988 ( .A(n8254), .B(n4095), .Z(n10455) );
  XNOR U9989 ( .A(n10456), .B(n8279), .Z(n4095) );
  NOR U9990 ( .A(n8227), .B(n7152), .Z(n10456) );
  XNOR U9991 ( .A(round_reg[1373]), .B(n10457), .Z(n7152) );
  XNOR U9992 ( .A(round_reg[188]), .B(n9112), .Z(n8227) );
  XOR U9993 ( .A(n10458), .B(n8275), .Z(n8254) );
  ANDN U9994 ( .B(n8223), .A(n7156), .Z(n10458) );
  XOR U9995 ( .A(round_reg[1593]), .B(n10290), .Z(n7156) );
  XOR U9996 ( .A(round_reg[43]), .B(n9992), .Z(n8223) );
  XNOR U9997 ( .A(n10459), .B(n10460), .Z(n3643) );
  ANDN U9998 ( .B(n8225), .A(n7161), .Z(n10459) );
  XNOR U9999 ( .A(round_reg[1467]), .B(n9195), .Z(n7161) );
  XOR U10000 ( .A(n10461), .B(n7105), .Z(n8203) );
  NOR U10001 ( .A(n10386), .B(n8171), .Z(n10461) );
  XOR U10002 ( .A(round_reg[248]), .B(n10351), .Z(n8171) );
  NOR U10003 ( .A(n5653), .B(n5652), .Z(n10446) );
  XOR U10004 ( .A(n10462), .B(n1715), .Z(n5652) );
  XNOR U10005 ( .A(n9014), .B(n6334), .Z(n1715) );
  XNOR U10006 ( .A(n10463), .B(n10464), .Z(n6334) );
  XNOR U10007 ( .A(n5413), .B(n3624), .Z(n10464) );
  XOR U10008 ( .A(n10465), .B(n10466), .Z(n3624) );
  NOR U10009 ( .A(n8189), .B(n10467), .Z(n10465) );
  XNOR U10010 ( .A(n10468), .B(n10469), .Z(n5413) );
  AND U10011 ( .A(n8179), .B(n10470), .Z(n10468) );
  XNOR U10012 ( .A(n10471), .B(n10472), .Z(n10463) );
  XOR U10013 ( .A(n2089), .B(n5524), .Z(n10472) );
  XOR U10014 ( .A(n10473), .B(n10474), .Z(n5524) );
  ANDN U10015 ( .B(n8183), .A(n10475), .Z(n10473) );
  XOR U10016 ( .A(n10476), .B(n10477), .Z(n2089) );
  NOR U10017 ( .A(n9147), .B(n10478), .Z(n10476) );
  XOR U10018 ( .A(n10479), .B(n10480), .Z(n9014) );
  XNOR U10019 ( .A(n3452), .B(n5054), .Z(n10480) );
  XOR U10020 ( .A(n10481), .B(n8124), .Z(n5054) );
  ANDN U10021 ( .B(n8125), .A(n10401), .Z(n10481) );
  XNOR U10022 ( .A(n10482), .B(n9073), .Z(n3452) );
  NOR U10023 ( .A(n10404), .B(n9072), .Z(n10482) );
  XNOR U10024 ( .A(n4029), .B(n10483), .Z(n10479) );
  XOR U10025 ( .A(n8114), .B(n2448), .Z(n10483) );
  XOR U10026 ( .A(n10484), .B(n8134), .Z(n2448) );
  AND U10027 ( .A(n10485), .B(n8135), .Z(n10484) );
  XNOR U10028 ( .A(n10486), .B(n8121), .Z(n8114) );
  AND U10029 ( .A(n10396), .B(n8120), .Z(n10486) );
  XOR U10030 ( .A(n10487), .B(n8131), .Z(n4029) );
  NOR U10031 ( .A(n8130), .B(n10393), .Z(n10487) );
  XOR U10032 ( .A(n9737), .B(n2056), .Z(n5653) );
  XNOR U10033 ( .A(n7472), .B(n10488), .Z(n2056) );
  XOR U10034 ( .A(n10489), .B(n10490), .Z(n7472) );
  XOR U10035 ( .A(n3736), .B(n5106), .Z(n10490) );
  XOR U10036 ( .A(n10491), .B(n8536), .Z(n5106) );
  XOR U10037 ( .A(round_reg[468]), .B(n9997), .Z(n8536) );
  ANDN U10038 ( .B(n9735), .A(n9736), .Z(n10491) );
  XOR U10039 ( .A(round_reg[1288]), .B(n10492), .Z(n9736) );
  XNOR U10040 ( .A(round_reg[107]), .B(n9392), .Z(n9735) );
  XOR U10041 ( .A(n10493), .B(n9793), .Z(n3736) );
  XOR U10042 ( .A(round_reg[634]), .B(n10494), .Z(n9793) );
  ANDN U10043 ( .B(n9743), .A(n9745), .Z(n10493) );
  XOR U10044 ( .A(round_reg[1445]), .B(n10495), .Z(n9745) );
  XOR U10045 ( .A(round_reg[225]), .B(n10496), .Z(n9743) );
  XOR U10046 ( .A(n4163), .B(n10497), .Z(n10489) );
  XOR U10047 ( .A(n1674), .B(n9783), .Z(n10497) );
  XNOR U10048 ( .A(n10498), .B(n7529), .Z(n9783) );
  XOR U10049 ( .A(round_reg[398]), .B(n9456), .Z(n7529) );
  ANDN U10050 ( .B(n9732), .A(n9733), .Z(n10498) );
  XOR U10051 ( .A(round_reg[1571]), .B(n9449), .Z(n9733) );
  XOR U10052 ( .A(round_reg[21]), .B(n9987), .Z(n9732) );
  XNOR U10053 ( .A(n10499), .B(n7523), .Z(n1674) );
  XOR U10054 ( .A(round_reg[347]), .B(n9975), .Z(n7523) );
  AND U10055 ( .A(n9741), .B(n9740), .Z(n10499) );
  XNOR U10056 ( .A(round_reg[273]), .B(n10500), .Z(n9740) );
  XNOR U10057 ( .A(round_reg[1506]), .B(n10442), .Z(n9741) );
  XNOR U10058 ( .A(n10501), .B(n7533), .Z(n4163) );
  XOR U10059 ( .A(round_reg[566]), .B(n9914), .Z(n7533) );
  ANDN U10060 ( .B(n9795), .A(n10419), .Z(n10501) );
  XOR U10061 ( .A(n10502), .B(n9795), .Z(n9737) );
  XNOR U10062 ( .A(round_reg[166]), .B(n10503), .Z(n9795) );
  ANDN U10063 ( .B(n10419), .A(n7531), .Z(n10502) );
  XOR U10064 ( .A(round_reg[975]), .B(n10504), .Z(n7531) );
  XOR U10065 ( .A(round_reg[1351]), .B(n9925), .Z(n10419) );
  XOR U10066 ( .A(n10505), .B(n6204), .Z(out[1014]) );
  XOR U10067 ( .A(n8270), .B(n4925), .Z(n6204) );
  XOR U10068 ( .A(n6167), .B(n6077), .Z(n4925) );
  XNOR U10069 ( .A(n10506), .B(n10507), .Z(n6077) );
  XNOR U10070 ( .A(n3647), .B(n4100), .Z(n10507) );
  XNOR U10071 ( .A(n10508), .B(n8331), .Z(n4100) );
  NOR U10072 ( .A(n8267), .B(n7205), .Z(n10508) );
  XNOR U10073 ( .A(round_reg[1372]), .B(n10509), .Z(n7205) );
  XOR U10074 ( .A(round_reg[187]), .B(n9195), .Z(n8267) );
  XOR U10075 ( .A(n10510), .B(n10511), .Z(n3647) );
  ANDN U10076 ( .B(n7214), .A(n8265), .Z(n10510) );
  XOR U10077 ( .A(round_reg[1466]), .B(n9918), .Z(n7214) );
  XOR U10078 ( .A(n5252), .B(n10512), .Z(n10506) );
  XNOR U10079 ( .A(n8306), .B(n1886), .Z(n10512) );
  XNOR U10080 ( .A(n10513), .B(n8324), .Z(n1886) );
  ANDN U10081 ( .B(n7222), .A(n8260), .Z(n10513) );
  XNOR U10082 ( .A(round_reg[294]), .B(n9889), .Z(n8260) );
  XOR U10083 ( .A(round_reg[1527]), .B(n10436), .Z(n7222) );
  IV U10084 ( .A(n9844), .Z(n10436) );
  XOR U10085 ( .A(n10514), .B(n8327), .Z(n8306) );
  ANDN U10086 ( .B(n7209), .A(n8263), .Z(n10514) );
  XNOR U10087 ( .A(round_reg[42]), .B(n10515), .Z(n8263) );
  XNOR U10088 ( .A(round_reg[1592]), .B(n9092), .Z(n7209) );
  XNOR U10089 ( .A(n10516), .B(n8329), .Z(n5252) );
  ANDN U10090 ( .B(n8258), .A(n7218), .Z(n10516) );
  XNOR U10091 ( .A(round_reg[1309]), .B(n10517), .Z(n7218) );
  XOR U10092 ( .A(round_reg[64]), .B(n10518), .Z(n8258) );
  XOR U10093 ( .A(n10519), .B(n10520), .Z(n6167) );
  XNOR U10094 ( .A(n3382), .B(n5777), .Z(n10520) );
  XNOR U10095 ( .A(n10521), .B(n7162), .Z(n5777) );
  XNOR U10096 ( .A(round_reg[1026]), .B(n10522), .Z(n7162) );
  ANDN U10097 ( .B(n7163), .A(n10460), .Z(n10521) );
  XOR U10098 ( .A(n10523), .B(n8220), .Z(n3382) );
  IV U10099 ( .A(n7170), .Z(n8220) );
  XNOR U10100 ( .A(round_reg[1139]), .B(n10524), .Z(n7170) );
  ANDN U10101 ( .B(n7171), .A(n8272), .Z(n10523) );
  XOR U10102 ( .A(round_reg[369]), .B(n9601), .Z(n8272) );
  XNOR U10103 ( .A(round_reg[736]), .B(n10226), .Z(n7171) );
  XOR U10104 ( .A(n5431), .B(n10525), .Z(n10519) );
  XOR U10105 ( .A(n7147), .B(n2264), .Z(n10525) );
  XNOR U10106 ( .A(n10526), .B(n7157), .Z(n2264) );
  XOR U10107 ( .A(round_reg[1165]), .B(n10527), .Z(n7157) );
  ANDN U10108 ( .B(n7158), .A(n8275), .Z(n10526) );
  XOR U10109 ( .A(round_reg[420]), .B(n10528), .Z(n8275) );
  XNOR U10110 ( .A(n10530), .B(n7166), .Z(n7147) );
  XOR U10111 ( .A(round_reg[1237]), .B(n10531), .Z(n7166) );
  ANDN U10112 ( .B(n7167), .A(n8277), .Z(n10530) );
  XOR U10113 ( .A(round_reg[490]), .B(n10044), .Z(n8277) );
  XOR U10114 ( .A(round_reg[879]), .B(n10532), .Z(n7167) );
  XNOR U10115 ( .A(n10533), .B(n7153), .Z(n5431) );
  XOR U10116 ( .A(round_reg[997]), .B(n10534), .Z(n7153) );
  ANDN U10117 ( .B(n7154), .A(n8279), .Z(n10533) );
  XOR U10118 ( .A(round_reg[524]), .B(n10535), .Z(n8279) );
  XNOR U10119 ( .A(round_reg[950]), .B(n10536), .Z(n7154) );
  XOR U10120 ( .A(n10537), .B(n7163), .Z(n8270) );
  XNOR U10121 ( .A(round_reg[658]), .B(n10538), .Z(n7163) );
  ANDN U10122 ( .B(n10460), .A(n8225), .Z(n10537) );
  XOR U10123 ( .A(round_reg[247]), .B(n9844), .Z(n8225) );
  XOR U10124 ( .A(n10539), .B(n10540), .Z(n9844) );
  XOR U10125 ( .A(round_reg[592]), .B(n10541), .Z(n10460) );
  ANDN U10126 ( .B(n5658), .A(n5656), .Z(n10505) );
  XNOR U10127 ( .A(n10542), .B(n1724), .Z(n5656) );
  XOR U10128 ( .A(n10543), .B(n10544), .Z(n9068) );
  XNOR U10129 ( .A(n3454), .B(n5059), .Z(n10544) );
  XNOR U10130 ( .A(n10545), .B(n8185), .Z(n5059) );
  NOR U10131 ( .A(n10474), .B(n8184), .Z(n10545) );
  XNOR U10132 ( .A(n10546), .B(n9149), .Z(n3454) );
  NOR U10133 ( .A(n10477), .B(n9148), .Z(n10546) );
  XNOR U10134 ( .A(n4063), .B(n10547), .Z(n10543) );
  XOR U10135 ( .A(n8174), .B(n2453), .Z(n10547) );
  XOR U10136 ( .A(n10548), .B(n8194), .Z(n2453) );
  ANDN U10137 ( .B(n8195), .A(n10549), .Z(n10548) );
  XNOR U10138 ( .A(n10550), .B(n8181), .Z(n8174) );
  AND U10139 ( .A(n10469), .B(n8180), .Z(n10550) );
  XOR U10140 ( .A(n10551), .B(n8191), .Z(n4063) );
  NOR U10141 ( .A(n8190), .B(n10466), .Z(n10551) );
  XNOR U10142 ( .A(n10552), .B(n10553), .Z(n6338) );
  XNOR U10143 ( .A(n5421), .B(n3628), .Z(n10553) );
  XNOR U10144 ( .A(n10554), .B(n10555), .Z(n3628) );
  ANDN U10145 ( .B(n10556), .A(n8243), .Z(n10554) );
  XNOR U10146 ( .A(n10557), .B(n10558), .Z(n5421) );
  ANDN U10147 ( .B(n8233), .A(n10559), .Z(n10557) );
  XNOR U10148 ( .A(n10560), .B(n10561), .Z(n10552) );
  XOR U10149 ( .A(n2093), .B(n5569), .Z(n10561) );
  XOR U10150 ( .A(n10562), .B(n10563), .Z(n5569) );
  ANDN U10151 ( .B(n8237), .A(n10564), .Z(n10562) );
  XOR U10152 ( .A(n10565), .B(n10566), .Z(n2093) );
  ANDN U10153 ( .B(n9224), .A(n10567), .Z(n10565) );
  XOR U10154 ( .A(n9805), .B(n5168), .Z(n5658) );
  XOR U10155 ( .A(n8717), .B(n7534), .Z(n5168) );
  XNOR U10156 ( .A(n10568), .B(n10569), .Z(n7534) );
  XOR U10157 ( .A(n9866), .B(n4166), .Z(n10569) );
  XOR U10158 ( .A(n10570), .B(n7632), .Z(n4166) );
  XOR U10159 ( .A(round_reg[565]), .B(n10002), .Z(n7632) );
  ANDN U10160 ( .B(n10117), .A(n10571), .Z(n10570) );
  XOR U10161 ( .A(n10572), .B(n7627), .Z(n9866) );
  XNOR U10162 ( .A(round_reg[397]), .B(n9541), .Z(n7627) );
  IV U10163 ( .A(n10573), .Z(n9541) );
  AND U10164 ( .A(n9800), .B(n9799), .Z(n10572) );
  XNOR U10165 ( .A(round_reg[20]), .B(n10574), .Z(n9799) );
  XOR U10166 ( .A(n3740), .B(n10575), .Z(n10568) );
  XOR U10167 ( .A(n5116), .B(n1679), .Z(n10575) );
  XNOR U10168 ( .A(n10576), .B(n7622), .Z(n1679) );
  XOR U10169 ( .A(round_reg[346]), .B(n9865), .Z(n7622) );
  ANDN U10170 ( .B(n9808), .A(n9809), .Z(n10576) );
  XNOR U10171 ( .A(round_reg[272]), .B(n10577), .Z(n9808) );
  XNOR U10172 ( .A(n10578), .B(n8658), .Z(n5116) );
  XNOR U10173 ( .A(round_reg[467]), .B(n10579), .Z(n8658) );
  ANDN U10174 ( .B(n9811), .A(n9812), .Z(n10578) );
  XNOR U10175 ( .A(round_reg[106]), .B(n9468), .Z(n9811) );
  XNOR U10176 ( .A(n10580), .B(n10115), .Z(n3740) );
  NOR U10177 ( .A(n9802), .B(n9804), .Z(n10580) );
  XNOR U10178 ( .A(round_reg[224]), .B(n10581), .Z(n9802) );
  XOR U10179 ( .A(n10582), .B(n10583), .Z(n8717) );
  XOR U10180 ( .A(n6300), .B(n2309), .Z(n10583) );
  XOR U10181 ( .A(n10584), .B(n9875), .Z(n2309) );
  ANDN U10182 ( .B(n7699), .A(n7700), .Z(n10584) );
  XNOR U10183 ( .A(round_reg[1066]), .B(n9468), .Z(n7699) );
  XNOR U10184 ( .A(n10585), .B(n10586), .Z(n9468) );
  XNOR U10185 ( .A(n10587), .B(n9880), .Z(n6300) );
  ANDN U10186 ( .B(n7690), .A(n7691), .Z(n10587) );
  XNOR U10187 ( .A(round_reg[1115]), .B(n10588), .Z(n7690) );
  XOR U10188 ( .A(n3832), .B(n10589), .Z(n10582) );
  XOR U10189 ( .A(n5138), .B(n5449), .Z(n10589) );
  XNOR U10190 ( .A(n10590), .B(n9872), .Z(n5449) );
  ANDN U10191 ( .B(n7703), .A(n7705), .Z(n10590) );
  XOR U10192 ( .A(round_reg[1205]), .B(n10002), .Z(n7703) );
  XNOR U10193 ( .A(n10591), .B(n9883), .Z(n5138) );
  ANDN U10194 ( .B(n8714), .A(n8715), .Z(n10591) );
  XNOR U10195 ( .A(round_reg[1277]), .B(n10592), .Z(n8714) );
  XOR U10196 ( .A(n10593), .B(n10594), .Z(n3832) );
  ANDN U10197 ( .B(n7695), .A(n7696), .Z(n10593) );
  XOR U10198 ( .A(n10595), .B(n10117), .Z(n9805) );
  XNOR U10199 ( .A(round_reg[165]), .B(n10596), .Z(n10117) );
  ANDN U10200 ( .B(n10571), .A(n7630), .Z(n10595) );
  XOR U10201 ( .A(n10597), .B(n6209), .Z(out[1013]) );
  XOR U10202 ( .A(n8322), .B(n3555), .Z(n6209) );
  XOR U10203 ( .A(n6172), .B(n6083), .Z(n3555) );
  XNOR U10204 ( .A(n10598), .B(n10599), .Z(n6083) );
  XNOR U10205 ( .A(n3651), .B(n4103), .Z(n10599) );
  XNOR U10206 ( .A(n10600), .B(n8383), .Z(n4103) );
  NOR U10207 ( .A(n8319), .B(n7233), .Z(n10600) );
  XNOR U10208 ( .A(round_reg[1371]), .B(n10601), .Z(n7233) );
  XOR U10209 ( .A(round_reg[186]), .B(n9918), .Z(n8319) );
  XOR U10210 ( .A(n10602), .B(n10603), .Z(n3651) );
  ANDN U10211 ( .B(n7246), .A(n8317), .Z(n10602) );
  XOR U10212 ( .A(round_reg[1465]), .B(n9370), .Z(n7246) );
  IV U10213 ( .A(n10005), .Z(n9370) );
  XOR U10214 ( .A(n5255), .B(n10604), .Z(n10598) );
  XNOR U10215 ( .A(n8358), .B(n1890), .Z(n10604) );
  XOR U10216 ( .A(n10605), .B(n8376), .Z(n1890) );
  ANDN U10217 ( .B(n7250), .A(n8312), .Z(n10605) );
  XNOR U10218 ( .A(round_reg[293]), .B(n9263), .Z(n8312) );
  XOR U10219 ( .A(round_reg[1526]), .B(n10606), .Z(n7250) );
  XNOR U10220 ( .A(n10607), .B(n8379), .Z(n8358) );
  ANDN U10221 ( .B(n7237), .A(n8315), .Z(n10607) );
  XNOR U10222 ( .A(round_reg[41]), .B(n10207), .Z(n8315) );
  XNOR U10223 ( .A(round_reg[1591]), .B(n10608), .Z(n7237) );
  XNOR U10224 ( .A(n10609), .B(n8381), .Z(n5255) );
  ANDN U10225 ( .B(n8310), .A(n7242), .Z(n10609) );
  XNOR U10226 ( .A(round_reg[1308]), .B(n10610), .Z(n7242) );
  XOR U10227 ( .A(round_reg[127]), .B(n10611), .Z(n8310) );
  XOR U10228 ( .A(n10612), .B(n10613), .Z(n6172) );
  XNOR U10229 ( .A(n3386), .B(n5808), .Z(n10613) );
  XNOR U10230 ( .A(n10614), .B(n7215), .Z(n5808) );
  XNOR U10231 ( .A(round_reg[1025]), .B(n10615), .Z(n7215) );
  AND U10232 ( .A(n10511), .B(n7216), .Z(n10614) );
  XNOR U10233 ( .A(n10616), .B(n7223), .Z(n3386) );
  XNOR U10234 ( .A(round_reg[1138]), .B(n10617), .Z(n7223) );
  ANDN U10235 ( .B(n7224), .A(n8324), .Z(n10616) );
  XOR U10236 ( .A(round_reg[368]), .B(n9675), .Z(n8324) );
  XNOR U10237 ( .A(round_reg[735]), .B(n10618), .Z(n7224) );
  XOR U10238 ( .A(n5434), .B(n10619), .Z(n10612) );
  XOR U10239 ( .A(n7200), .B(n2271), .Z(n10619) );
  XOR U10240 ( .A(n10620), .B(n7211), .Z(n2271) );
  XNOR U10241 ( .A(round_reg[1164]), .B(n10535), .Z(n7211) );
  XOR U10242 ( .A(round_reg[419]), .B(n9928), .Z(n8327) );
  XOR U10243 ( .A(round_reg[781]), .B(n9095), .Z(n7210) );
  XNOR U10244 ( .A(n10621), .B(n7219), .Z(n7200) );
  XOR U10245 ( .A(round_reg[1236]), .B(n10622), .Z(n7219) );
  ANDN U10246 ( .B(n7220), .A(n8329), .Z(n10621) );
  XOR U10247 ( .A(round_reg[489]), .B(n10170), .Z(n8329) );
  XNOR U10248 ( .A(round_reg[878]), .B(n10623), .Z(n7220) );
  XNOR U10249 ( .A(n10624), .B(n7206), .Z(n5434) );
  XOR U10250 ( .A(round_reg[996]), .B(n10625), .Z(n7206) );
  ANDN U10251 ( .B(n7207), .A(n8331), .Z(n10624) );
  XOR U10252 ( .A(round_reg[523]), .B(n10626), .Z(n8331) );
  XNOR U10253 ( .A(round_reg[949]), .B(n10627), .Z(n7207) );
  XOR U10254 ( .A(n10628), .B(n7216), .Z(n8322) );
  XNOR U10255 ( .A(round_reg[657]), .B(n10629), .Z(n7216) );
  ANDN U10256 ( .B(n8265), .A(n10511), .Z(n10628) );
  XNOR U10257 ( .A(round_reg[591]), .B(n10630), .Z(n10511) );
  XNOR U10258 ( .A(round_reg[246]), .B(n9914), .Z(n8265) );
  ANDN U10259 ( .B(n5668), .A(n5666), .Z(n10597) );
  XNOR U10260 ( .A(n10631), .B(n1728), .Z(n5666) );
  XOR U10261 ( .A(n10632), .B(n10633), .Z(n9144) );
  XNOR U10262 ( .A(n3456), .B(n5064), .Z(n10633) );
  XOR U10263 ( .A(n10634), .B(n8238), .Z(n5064) );
  ANDN U10264 ( .B(n8239), .A(n10563), .Z(n10634) );
  XNOR U10265 ( .A(n10635), .B(n9226), .Z(n3456) );
  NOR U10266 ( .A(n10566), .B(n9225), .Z(n10635) );
  XNOR U10267 ( .A(n4098), .B(n10636), .Z(n10632) );
  XOR U10268 ( .A(n8228), .B(n2460), .Z(n10636) );
  XNOR U10269 ( .A(n10637), .B(n8249), .Z(n2460) );
  AND U10270 ( .A(n10638), .B(n8248), .Z(n10637) );
  XNOR U10271 ( .A(n10639), .B(n8235), .Z(n8228) );
  AND U10272 ( .A(n10558), .B(n8234), .Z(n10639) );
  XOR U10273 ( .A(n10640), .B(n8245), .Z(n4098) );
  ANDN U10274 ( .B(n10555), .A(n8244), .Z(n10640) );
  XNOR U10275 ( .A(n10641), .B(n10642), .Z(n6342) );
  XNOR U10276 ( .A(n5425), .B(n3632), .Z(n10642) );
  XOR U10277 ( .A(n10643), .B(n10644), .Z(n3632) );
  ANDN U10278 ( .B(n10645), .A(n8295), .Z(n10643) );
  XNOR U10279 ( .A(n10646), .B(n10647), .Z(n5425) );
  ANDN U10280 ( .B(n8285), .A(n10648), .Z(n10646) );
  XNOR U10281 ( .A(n10649), .B(n10650), .Z(n10641) );
  XOR U10282 ( .A(n2097), .B(n4226), .Z(n10650) );
  XNOR U10283 ( .A(n10651), .B(n10652), .Z(n4226) );
  ANDN U10284 ( .B(n8289), .A(n10653), .Z(n10651) );
  XOR U10285 ( .A(n10654), .B(n10655), .Z(n2097) );
  NOR U10286 ( .A(n9331), .B(n10656), .Z(n10654) );
  XOR U10287 ( .A(n9876), .B(n5382), .Z(n5668) );
  XOR U10288 ( .A(n7615), .B(n8779), .Z(n5382) );
  XNOR U10289 ( .A(n10657), .B(n10658), .Z(n8779) );
  XOR U10290 ( .A(n5455), .B(n3836), .Z(n10658) );
  XOR U10291 ( .A(n10659), .B(n10660), .Z(n3836) );
  ANDN U10292 ( .B(n7770), .A(n7771), .Z(n10659) );
  XOR U10293 ( .A(round_reg[925]), .B(n9556), .Z(n7771) );
  XOR U10294 ( .A(n10661), .B(n9942), .Z(n5455) );
  XOR U10295 ( .A(round_reg[821]), .B(n10662), .Z(n7779) );
  XOR U10296 ( .A(round_reg[1204]), .B(n10663), .Z(n7778) );
  XOR U10297 ( .A(n6304), .B(n10664), .Z(n10657) );
  XOR U10298 ( .A(n2316), .B(n5170), .Z(n10664) );
  XNOR U10299 ( .A(n10665), .B(n9954), .Z(n5170) );
  ANDN U10300 ( .B(n8775), .A(n8777), .Z(n10665) );
  XOR U10301 ( .A(round_reg[854]), .B(n10666), .Z(n8777) );
  XNOR U10302 ( .A(round_reg[1276]), .B(n10667), .Z(n8775) );
  XNOR U10303 ( .A(n10668), .B(n9945), .Z(n2316) );
  AND U10304 ( .A(n7776), .B(n7774), .Z(n10668) );
  IV U10305 ( .A(n9946), .Z(n7774) );
  XOR U10306 ( .A(round_reg[1065]), .B(n9552), .Z(n9946) );
  XNOR U10307 ( .A(round_reg[697]), .B(n9389), .Z(n7776) );
  XOR U10308 ( .A(n10669), .B(n9951), .Z(n6304) );
  ANDN U10309 ( .B(n7765), .A(n7766), .Z(n10669) );
  XOR U10310 ( .A(round_reg[711]), .B(n9925), .Z(n7766) );
  XNOR U10311 ( .A(round_reg[1114]), .B(n10670), .Z(n7765) );
  XOR U10312 ( .A(n10671), .B(n10672), .Z(n7615) );
  XOR U10313 ( .A(n3745), .B(n5118), .Z(n10672) );
  XOR U10314 ( .A(n10673), .B(n8716), .Z(n5118) );
  ANDN U10315 ( .B(n9882), .A(n9883), .Z(n10673) );
  XOR U10316 ( .A(round_reg[1286]), .B(n10674), .Z(n9883) );
  XNOR U10317 ( .A(n10675), .B(n7701), .Z(n3745) );
  XOR U10318 ( .A(round_reg[1443]), .B(n10676), .Z(n9875) );
  XOR U10319 ( .A(n4169), .B(n10677), .Z(n10671) );
  XOR U10320 ( .A(n1684), .B(n9936), .Z(n10677) );
  XOR U10321 ( .A(n10678), .B(n7704), .Z(n9936) );
  ANDN U10322 ( .B(n9871), .A(n9872), .Z(n10678) );
  XOR U10323 ( .A(round_reg[1569]), .B(n9219), .Z(n9872) );
  XNOR U10324 ( .A(n10679), .B(n7692), .Z(n1684) );
  ANDN U10325 ( .B(n9879), .A(n9880), .Z(n10679) );
  XOR U10326 ( .A(round_reg[1504]), .B(n10581), .Z(n9880) );
  XNOR U10327 ( .A(n10680), .B(n7697), .Z(n4169) );
  XNOR U10328 ( .A(n10682), .B(n10681), .Z(n9876) );
  NOR U10329 ( .A(n7695), .B(n10594), .Z(n10682) );
  XNOR U10330 ( .A(round_reg[1349]), .B(n10293), .Z(n10594) );
  XNOR U10331 ( .A(round_reg[973]), .B(n10683), .Z(n7695) );
  XOR U10332 ( .A(n10684), .B(n6214), .Z(out[1012]) );
  XOR U10333 ( .A(n8374), .B(n3558), .Z(n6214) );
  XOR U10334 ( .A(n6178), .B(n6089), .Z(n3558) );
  XNOR U10335 ( .A(n10685), .B(n10686), .Z(n6089) );
  XNOR U10336 ( .A(n3655), .B(n4106), .Z(n10686) );
  XOR U10337 ( .A(n10687), .B(n8436), .Z(n4106) );
  NOR U10338 ( .A(n8371), .B(n7301), .Z(n10687) );
  XNOR U10339 ( .A(round_reg[1370]), .B(n10688), .Z(n7301) );
  XNOR U10340 ( .A(round_reg[185]), .B(n10005), .Z(n8371) );
  XOR U10341 ( .A(n10689), .B(n10690), .Z(n10005) );
  XOR U10342 ( .A(n10691), .B(n10692), .Z(n3655) );
  AND U10343 ( .A(n7314), .B(n8369), .Z(n10691) );
  XNOR U10344 ( .A(round_reg[1464]), .B(n10422), .Z(n7314) );
  XNOR U10345 ( .A(n5258), .B(n10693), .Z(n10685) );
  XOR U10346 ( .A(n8411), .B(n1894), .Z(n10693) );
  XNOR U10347 ( .A(n10694), .B(n8429), .Z(n1894) );
  ANDN U10348 ( .B(n7318), .A(n8364), .Z(n10694) );
  XNOR U10349 ( .A(round_reg[292]), .B(n10431), .Z(n8364) );
  XNOR U10350 ( .A(round_reg[1525]), .B(n10002), .Z(n7318) );
  XNOR U10351 ( .A(n10695), .B(n8432), .Z(n8411) );
  ANDN U10352 ( .B(n7305), .A(n8367), .Z(n10695) );
  XNOR U10353 ( .A(round_reg[40]), .B(n10289), .Z(n8367) );
  XNOR U10354 ( .A(round_reg[1590]), .B(n10696), .Z(n7305) );
  XNOR U10355 ( .A(n10697), .B(n8434), .Z(n5258) );
  ANDN U10356 ( .B(n7310), .A(n8362), .Z(n10697) );
  XNOR U10357 ( .A(round_reg[126]), .B(n10698), .Z(n8362) );
  XNOR U10358 ( .A(round_reg[1307]), .B(n9975), .Z(n7310) );
  XOR U10359 ( .A(n10699), .B(n10700), .Z(n6178) );
  XOR U10360 ( .A(n3394), .B(n5835), .Z(n10700) );
  XOR U10361 ( .A(n10701), .B(n7247), .Z(n5835) );
  XOR U10362 ( .A(round_reg[1024]), .B(n10518), .Z(n7247) );
  AND U10363 ( .A(n7248), .B(n10603), .Z(n10701) );
  XNOR U10364 ( .A(n10702), .B(n7251), .Z(n3394) );
  XNOR U10365 ( .A(round_reg[1137]), .B(n9913), .Z(n7251) );
  AND U10366 ( .A(n8376), .B(n7252), .Z(n10702) );
  XNOR U10367 ( .A(round_reg[734]), .B(n10382), .Z(n7252) );
  XNOR U10368 ( .A(round_reg[367]), .B(n9079), .Z(n8376) );
  XOR U10369 ( .A(n5440), .B(n10703), .Z(n10699) );
  XOR U10370 ( .A(n7228), .B(n2278), .Z(n10703) );
  XOR U10371 ( .A(n10704), .B(n7239), .Z(n2278) );
  XNOR U10372 ( .A(round_reg[1163]), .B(n10626), .Z(n7239) );
  ANDN U10373 ( .B(n8379), .A(n7238), .Z(n10704) );
  XOR U10374 ( .A(round_reg[780]), .B(n10705), .Z(n7238) );
  XOR U10375 ( .A(round_reg[418]), .B(n10369), .Z(n8379) );
  XOR U10376 ( .A(n10706), .B(n7244), .Z(n7228) );
  XNOR U10377 ( .A(round_reg[1235]), .B(n10707), .Z(n7244) );
  XOR U10378 ( .A(round_reg[488]), .B(n10281), .Z(n8381) );
  XOR U10379 ( .A(round_reg[877]), .B(n10708), .Z(n7243) );
  XNOR U10380 ( .A(n10709), .B(n7234), .Z(n5440) );
  XOR U10381 ( .A(round_reg[995]), .B(n9218), .Z(n7234) );
  ANDN U10382 ( .B(n7235), .A(n8383), .Z(n10709) );
  XOR U10383 ( .A(round_reg[522]), .B(n10710), .Z(n8383) );
  XNOR U10384 ( .A(round_reg[948]), .B(n10711), .Z(n7235) );
  XOR U10385 ( .A(n10712), .B(n7248), .Z(n8374) );
  XOR U10386 ( .A(round_reg[656]), .B(n10445), .Z(n7248) );
  XNOR U10387 ( .A(round_reg[590]), .B(n10713), .Z(n10603) );
  XNOR U10388 ( .A(round_reg[245]), .B(n10002), .Z(n8317) );
  XNOR U10389 ( .A(n10714), .B(n10715), .Z(n10002) );
  ANDN U10390 ( .B(n5672), .A(n5670), .Z(n10684) );
  XNOR U10391 ( .A(n10716), .B(n1732), .Z(n5670) );
  XOR U10392 ( .A(n10717), .B(n10718), .Z(n9221) );
  XNOR U10393 ( .A(n3458), .B(n5069), .Z(n10718) );
  XOR U10394 ( .A(n10719), .B(n8290), .Z(n5069) );
  AND U10395 ( .A(n10652), .B(n8291), .Z(n10719) );
  XNOR U10396 ( .A(n10720), .B(n9332), .Z(n3458) );
  ANDN U10397 ( .B(n9333), .A(n10655), .Z(n10720) );
  XNOR U10398 ( .A(n4130), .B(n10721), .Z(n10717) );
  XOR U10399 ( .A(n8280), .B(n2467), .Z(n10721) );
  XOR U10400 ( .A(n10722), .B(n8300), .Z(n2467) );
  AND U10401 ( .A(n10723), .B(n8301), .Z(n10722) );
  XNOR U10402 ( .A(n10724), .B(n8287), .Z(n8280) );
  AND U10403 ( .A(n10647), .B(n10725), .Z(n10724) );
  XOR U10404 ( .A(n10726), .B(n8297), .Z(n4130) );
  NOR U10405 ( .A(n8296), .B(n10644), .Z(n10726) );
  XNOR U10406 ( .A(n10727), .B(n10728), .Z(n6346) );
  XNOR U10407 ( .A(n5429), .B(n3636), .Z(n10728) );
  XNOR U10408 ( .A(n10729), .B(n10730), .Z(n3636) );
  XNOR U10409 ( .A(n10732), .B(n10733), .Z(n5429) );
  ANDN U10410 ( .B(n8337), .A(n10734), .Z(n10732) );
  XNOR U10411 ( .A(n10735), .B(n10736), .Z(n10727) );
  XOR U10412 ( .A(n2100), .B(n4229), .Z(n10736) );
  XNOR U10413 ( .A(n10737), .B(n10738), .Z(n4229) );
  ANDN U10414 ( .B(n8341), .A(n10739), .Z(n10737) );
  XOR U10415 ( .A(n10740), .B(n10741), .Z(n2100) );
  NOR U10416 ( .A(n9401), .B(n10742), .Z(n10740) );
  XNOR U10417 ( .A(n9947), .B(n2066), .Z(n5672) );
  XNOR U10418 ( .A(n7685), .B(n8835), .Z(n2066) );
  XNOR U10419 ( .A(n10743), .B(n10744), .Z(n8835) );
  XOR U10420 ( .A(n5460), .B(n3840), .Z(n10744) );
  XOR U10421 ( .A(n10745), .B(n10746), .Z(n3840) );
  IV U10422 ( .A(n7841), .Z(n10200) );
  XNOR U10423 ( .A(round_reg[924]), .B(n9637), .Z(n7841) );
  XOR U10424 ( .A(n10054), .B(n10747), .Z(n5460) );
  XOR U10425 ( .A(n10748), .B(n10749), .Z(n10747) );
  NAND U10426 ( .A(n10750), .B(n10751), .Z(n10749) );
  AND U10427 ( .A(n6883), .B(n4340), .Z(n10751) );
  IV U10428 ( .A(rc_i[3]), .Z(n4340) );
  AND U10429 ( .A(n4635), .B(n4608), .Z(n6883) );
  IV U10430 ( .A(rc_i[6]), .Z(n4608) );
  IV U10431 ( .A(rc_i[5]), .Z(n4635) );
  AND U10432 ( .A(n4566), .B(n4491), .Z(n10750) );
  IV U10433 ( .A(rc_i[11]), .Z(n4491) );
  IV U10434 ( .A(rc_i[10]), .Z(n4566) );
  AND U10435 ( .A(n7838), .B(n10055), .Z(n10748) );
  XNOR U10436 ( .A(round_reg[1203]), .B(n10752), .Z(n10055) );
  XOR U10437 ( .A(round_reg[820]), .B(n9757), .Z(n7838) );
  XOR U10438 ( .A(n6308), .B(n10753), .Z(n10743) );
  XOR U10439 ( .A(n2327), .B(n5206), .Z(n10753) );
  XNOR U10440 ( .A(n10754), .B(n10066), .Z(n5206) );
  AND U10441 ( .A(n8839), .B(n10067), .Z(n10754) );
  XNOR U10442 ( .A(round_reg[1275]), .B(n10440), .Z(n10067) );
  XOR U10443 ( .A(round_reg[853]), .B(n10755), .Z(n8839) );
  XNOR U10444 ( .A(n10756), .B(n10058), .Z(n2327) );
  XOR U10445 ( .A(round_reg[1064]), .B(n9632), .Z(n7826) );
  XNOR U10446 ( .A(round_reg[696]), .B(n9466), .Z(n7827) );
  XOR U10447 ( .A(n10757), .B(n10063), .Z(n6308) );
  XOR U10448 ( .A(round_reg[1113]), .B(n10041), .Z(n7830) );
  XOR U10449 ( .A(round_reg[710]), .B(n10758), .Z(n7831) );
  XOR U10450 ( .A(n10759), .B(n10760), .Z(n7685) );
  XNOR U10451 ( .A(n3749), .B(n5120), .Z(n10760) );
  XNOR U10452 ( .A(n10761), .B(n8776), .Z(n5120) );
  XOR U10453 ( .A(round_reg[465]), .B(n10762), .Z(n8776) );
  ANDN U10454 ( .B(n9953), .A(n9954), .Z(n10761) );
  XOR U10455 ( .A(round_reg[1285]), .B(n10763), .Z(n9954) );
  XNOR U10456 ( .A(round_reg[104]), .B(n9632), .Z(n9953) );
  XOR U10457 ( .A(n10764), .B(n7775), .Z(n3749) );
  XOR U10458 ( .A(round_reg[631]), .B(n10608), .Z(n7775) );
  ANDN U10459 ( .B(n9944), .A(n9945), .Z(n10764) );
  XOR U10460 ( .A(round_reg[1442]), .B(n9968), .Z(n9945) );
  XOR U10461 ( .A(round_reg[222]), .B(n9115), .Z(n9944) );
  XNOR U10462 ( .A(n4172), .B(n10765), .Z(n10759) );
  XOR U10463 ( .A(n1689), .B(n10049), .Z(n10765) );
  XOR U10464 ( .A(n10766), .B(n7780), .Z(n10049) );
  XNOR U10465 ( .A(round_reg[395]), .B(n10356), .Z(n7780) );
  AND U10466 ( .A(n9942), .B(n9941), .Z(n10766) );
  XOR U10467 ( .A(round_reg[18]), .B(n10767), .Z(n9941) );
  XNOR U10468 ( .A(round_reg[1568]), .B(n9683), .Z(n9942) );
  XOR U10469 ( .A(n10768), .B(n7767), .Z(n1689) );
  XNOR U10470 ( .A(round_reg[344]), .B(n10020), .Z(n7767) );
  AND U10471 ( .A(n9951), .B(n9950), .Z(n10768) );
  XOR U10472 ( .A(round_reg[270]), .B(n10713), .Z(n9950) );
  XOR U10473 ( .A(round_reg[1503]), .B(n9894), .Z(n9951) );
  XOR U10474 ( .A(n10769), .B(n7772), .Z(n4172) );
  XNOR U10475 ( .A(round_reg[563]), .B(n10752), .Z(n7772) );
  ANDN U10476 ( .B(n10076), .A(n10660), .Z(n10769) );
  XNOR U10477 ( .A(n10770), .B(n10076), .Z(n9947) );
  XOR U10478 ( .A(round_reg[163]), .B(n10676), .Z(n10076) );
  ANDN U10479 ( .B(n10660), .A(n7770), .Z(n10770) );
  XNOR U10480 ( .A(round_reg[972]), .B(n10771), .Z(n7770) );
  XOR U10481 ( .A(round_reg[1348]), .B(n10223), .Z(n10660) );
  XOR U10482 ( .A(n10772), .B(n6224), .Z(out[1011]) );
  XOR U10483 ( .A(n8427), .B(n6046), .Z(n6224) );
  XOR U10484 ( .A(n6183), .B(n6094), .Z(n6046) );
  XNOR U10485 ( .A(n10773), .B(n10774), .Z(n6094) );
  XNOR U10486 ( .A(n3659), .B(n4109), .Z(n10774) );
  XNOR U10487 ( .A(n10775), .B(n8490), .Z(n4109) );
  NOR U10488 ( .A(n7354), .B(n8424), .Z(n10775) );
  XNOR U10489 ( .A(round_reg[184]), .B(n10422), .Z(n8424) );
  XNOR U10490 ( .A(round_reg[1369]), .B(n10776), .Z(n7354) );
  XNOR U10491 ( .A(n10777), .B(n10778), .Z(n3659) );
  ANDN U10492 ( .B(n7367), .A(n8422), .Z(n10777) );
  XNOR U10493 ( .A(round_reg[1463]), .B(n10211), .Z(n7367) );
  XNOR U10494 ( .A(n5261), .B(n10779), .Z(n10773) );
  XOR U10495 ( .A(n8464), .B(n1898), .Z(n10779) );
  XNOR U10496 ( .A(n10780), .B(n8483), .Z(n1898) );
  ANDN U10497 ( .B(n7371), .A(n8417), .Z(n10780) );
  XNOR U10498 ( .A(round_reg[291]), .B(n9449), .Z(n8417) );
  XNOR U10499 ( .A(round_reg[1524]), .B(n10781), .Z(n7371) );
  XNOR U10500 ( .A(n10782), .B(n8486), .Z(n8464) );
  ANDN U10501 ( .B(n7358), .A(n8420), .Z(n10782) );
  XNOR U10502 ( .A(round_reg[39]), .B(n10783), .Z(n8420) );
  XNOR U10503 ( .A(round_reg[1589]), .B(n9387), .Z(n7358) );
  XNOR U10504 ( .A(n10784), .B(n8488), .Z(n5261) );
  ANDN U10505 ( .B(n7363), .A(n8415), .Z(n10784) );
  XNOR U10506 ( .A(round_reg[125]), .B(n10785), .Z(n8415) );
  XNOR U10507 ( .A(round_reg[1306]), .B(n9865), .Z(n7363) );
  XOR U10508 ( .A(n10786), .B(n10787), .Z(n6183) );
  XNOR U10509 ( .A(n3398), .B(n5866), .Z(n10787) );
  XOR U10510 ( .A(n10788), .B(n7315), .Z(n5866) );
  XNOR U10511 ( .A(round_reg[1087]), .B(n10611), .Z(n7315) );
  ANDN U10512 ( .B(n7316), .A(n10692), .Z(n10788) );
  XNOR U10513 ( .A(n10789), .B(n7319), .Z(n3398) );
  XOR U10514 ( .A(round_reg[1136]), .B(n10790), .Z(n7319) );
  AND U10515 ( .A(n8429), .B(n7320), .Z(n10789) );
  XNOR U10516 ( .A(round_reg[733]), .B(n10457), .Z(n7320) );
  XNOR U10517 ( .A(round_reg[366]), .B(n10791), .Z(n8429) );
  XNOR U10518 ( .A(n5444), .B(n10792), .Z(n10786) );
  XNOR U10519 ( .A(n7296), .B(n2285), .Z(n10792) );
  XNOR U10520 ( .A(n10793), .B(n7307), .Z(n2285) );
  XNOR U10521 ( .A(round_reg[1162]), .B(n10710), .Z(n7307) );
  ANDN U10522 ( .B(n8432), .A(n7306), .Z(n10793) );
  XNOR U10523 ( .A(round_reg[779]), .B(n9208), .Z(n7306) );
  XOR U10524 ( .A(round_reg[417]), .B(n10140), .Z(n8432) );
  XNOR U10525 ( .A(n10794), .B(n7311), .Z(n7296) );
  XOR U10526 ( .A(round_reg[1234]), .B(n10795), .Z(n7311) );
  AND U10527 ( .A(n8434), .B(n7312), .Z(n10794) );
  XOR U10528 ( .A(round_reg[876]), .B(n10796), .Z(n7312) );
  XNOR U10529 ( .A(round_reg[487]), .B(n10797), .Z(n8434) );
  XNOR U10530 ( .A(n10798), .B(n7303), .Z(n5444) );
  XNOR U10531 ( .A(round_reg[994]), .B(n10799), .Z(n7303) );
  NOR U10532 ( .A(n7302), .B(n8436), .Z(n10798) );
  XNOR U10533 ( .A(round_reg[521]), .B(n10800), .Z(n8436) );
  XNOR U10534 ( .A(round_reg[947]), .B(n9544), .Z(n7302) );
  XOR U10535 ( .A(n10801), .B(n7316), .Z(n8427) );
  XOR U10536 ( .A(round_reg[655]), .B(n10504), .Z(n7316) );
  ANDN U10537 ( .B(n10692), .A(n8369), .Z(n10801) );
  XNOR U10538 ( .A(round_reg[244]), .B(n10663), .Z(n8369) );
  IV U10539 ( .A(n10781), .Z(n10663) );
  XOR U10540 ( .A(round_reg[589]), .B(n10802), .Z(n10692) );
  ANDN U10541 ( .B(n5676), .A(n5674), .Z(n10772) );
  XNOR U10542 ( .A(n10803), .B(n1737), .Z(n5674) );
  XOR U10543 ( .A(n10804), .B(n10805), .Z(n9328) );
  XNOR U10544 ( .A(n3460), .B(n5074), .Z(n10805) );
  XOR U10545 ( .A(n10806), .B(n8342), .Z(n5074) );
  AND U10546 ( .A(n10738), .B(n8343), .Z(n10806) );
  XNOR U10547 ( .A(n10807), .B(n9403), .Z(n3460) );
  NOR U10548 ( .A(n10741), .B(n9402), .Z(n10807) );
  XNOR U10549 ( .A(n4158), .B(n10808), .Z(n10804) );
  XOR U10550 ( .A(n8332), .B(n2478), .Z(n10808) );
  XNOR U10551 ( .A(n10809), .B(n8353), .Z(n2478) );
  AND U10552 ( .A(n10810), .B(n8352), .Z(n10809) );
  XNOR U10553 ( .A(n10811), .B(n8339), .Z(n8332) );
  AND U10554 ( .A(n10733), .B(n8338), .Z(n10811) );
  XOR U10555 ( .A(n10812), .B(n8349), .Z(n4158) );
  ANDN U10556 ( .B(n10730), .A(n8348), .Z(n10812) );
  XNOR U10557 ( .A(n10813), .B(n10814), .Z(n6350) );
  XNOR U10558 ( .A(n5433), .B(n3645), .Z(n10814) );
  XOR U10559 ( .A(n10815), .B(n10816), .Z(n3645) );
  NOR U10560 ( .A(n8399), .B(n10817), .Z(n10815) );
  XNOR U10561 ( .A(n10818), .B(n10819), .Z(n5433) );
  NOR U10562 ( .A(n8389), .B(n10820), .Z(n10818) );
  XNOR U10563 ( .A(n10821), .B(n10822), .Z(n10813) );
  XOR U10564 ( .A(n2104), .B(n4235), .Z(n10822) );
  XNOR U10565 ( .A(n10823), .B(n10824), .Z(n4235) );
  ANDN U10566 ( .B(n8393), .A(n10825), .Z(n10823) );
  XOR U10567 ( .A(n10826), .B(n10827), .Z(n2104) );
  NOR U10568 ( .A(n9478), .B(n10828), .Z(n10826) );
  XOR U10569 ( .A(n10059), .B(n5391), .Z(n5676) );
  XOR U10570 ( .A(n7760), .B(n8896), .Z(n5391) );
  XNOR U10571 ( .A(n10829), .B(n10830), .Z(n8896) );
  XOR U10572 ( .A(n5464), .B(n3844), .Z(n10830) );
  XOR U10573 ( .A(n10831), .B(n10832), .Z(n3844) );
  XNOR U10574 ( .A(round_reg[923]), .B(n9710), .Z(n7908) );
  XOR U10575 ( .A(n10833), .B(n10180), .Z(n5464) );
  XNOR U10576 ( .A(round_reg[819]), .B(n10524), .Z(n7905) );
  XOR U10577 ( .A(round_reg[1202]), .B(n10834), .Z(n7903) );
  XOR U10578 ( .A(n6312), .B(n10835), .Z(n10829) );
  XOR U10579 ( .A(n2334), .B(n5244), .Z(n10835) );
  XOR U10580 ( .A(n10836), .B(n10191), .Z(n5244) );
  XNOR U10581 ( .A(round_reg[852]), .B(n10837), .Z(n8899) );
  XOR U10582 ( .A(round_reg[1274]), .B(n10494), .Z(n8898) );
  XNOR U10583 ( .A(n10838), .B(n10183), .Z(n2334) );
  ANDN U10584 ( .B(n7894), .A(n7893), .Z(n10838) );
  XNOR U10585 ( .A(round_reg[1063]), .B(n9919), .Z(n7893) );
  XNOR U10586 ( .A(round_reg[695]), .B(n9550), .Z(n7894) );
  XOR U10587 ( .A(n10839), .B(n10188), .Z(n6312) );
  XOR U10588 ( .A(round_reg[1112]), .B(n10840), .Z(n7897) );
  XOR U10589 ( .A(n10841), .B(n10842), .Z(n7760) );
  XNOR U10590 ( .A(n3753), .B(n5122), .Z(n10842) );
  XOR U10591 ( .A(n10843), .B(n8840), .Z(n5122) );
  XNOR U10592 ( .A(round_reg[464]), .B(n10844), .Z(n8840) );
  ANDN U10593 ( .B(n10065), .A(n10066), .Z(n10843) );
  XOR U10594 ( .A(round_reg[1284]), .B(n10845), .Z(n10066) );
  XOR U10595 ( .A(round_reg[103]), .B(n9919), .Z(n10065) );
  XOR U10596 ( .A(n10846), .B(n10847), .Z(n9919) );
  XOR U10597 ( .A(n10848), .B(n7828), .Z(n3753) );
  XNOR U10598 ( .A(round_reg[630]), .B(n10536), .Z(n7828) );
  IV U10599 ( .A(n10696), .Z(n10536) );
  NOR U10600 ( .A(n10058), .B(n10057), .Z(n10848) );
  XNOR U10601 ( .A(round_reg[221]), .B(n9260), .Z(n10057) );
  XOR U10602 ( .A(round_reg[1441]), .B(n10099), .Z(n10058) );
  XNOR U10603 ( .A(n4175), .B(n10849), .Z(n10841) );
  XOR U10604 ( .A(n1694), .B(n10175), .Z(n10849) );
  XNOR U10605 ( .A(n10850), .B(n7837), .Z(n10175) );
  XNOR U10606 ( .A(round_reg[394]), .B(n9767), .Z(n7837) );
  IV U10607 ( .A(n10427), .Z(n9767) );
  XNOR U10608 ( .A(n10851), .B(n10852), .Z(n10427) );
  XOR U10609 ( .A(round_reg[1567]), .B(n9756), .Z(n10054) );
  XOR U10610 ( .A(round_reg[17]), .B(n10359), .Z(n10053) );
  XOR U10611 ( .A(n10853), .B(n7832), .Z(n1694) );
  XNOR U10612 ( .A(round_reg[343]), .B(n10854), .Z(n7832) );
  AND U10613 ( .A(n10063), .B(n10062), .Z(n10853) );
  XOR U10614 ( .A(round_reg[269]), .B(n10802), .Z(n10062) );
  XNOR U10615 ( .A(round_reg[1502]), .B(n9115), .Z(n10063) );
  XNOR U10616 ( .A(n10855), .B(n10856), .Z(n9115) );
  XOR U10617 ( .A(n10857), .B(n7842), .Z(n4175) );
  XNOR U10618 ( .A(round_reg[562]), .B(n10834), .Z(n7842) );
  NOR U10619 ( .A(n10746), .B(n10201), .Z(n10857) );
  XNOR U10620 ( .A(n10858), .B(n10201), .Z(n10059) );
  XNOR U10621 ( .A(round_reg[162]), .B(n9968), .Z(n10201) );
  AND U10622 ( .A(n10746), .B(n7840), .Z(n10858) );
  XOR U10623 ( .A(round_reg[971]), .B(n10859), .Z(n7840) );
  XOR U10624 ( .A(round_reg[1347]), .B(n10860), .Z(n10746) );
  XOR U10625 ( .A(n10861), .B(n6229), .Z(out[1010]) );
  XNOR U10626 ( .A(n8481), .B(n6105), .Z(n6229) );
  XOR U10627 ( .A(n6099), .B(n6188), .Z(n6105) );
  XNOR U10628 ( .A(n10862), .B(n10863), .Z(n6188) );
  XNOR U10629 ( .A(n2292), .B(n5448), .Z(n10863) );
  XNOR U10630 ( .A(n10864), .B(n7356), .Z(n5448) );
  XNOR U10631 ( .A(round_reg[993]), .B(n9395), .Z(n7356) );
  ANDN U10632 ( .B(n8490), .A(n7355), .Z(n10864) );
  XNOR U10633 ( .A(round_reg[946]), .B(n9624), .Z(n7355) );
  XOR U10634 ( .A(round_reg[520]), .B(n9213), .Z(n8490) );
  XNOR U10635 ( .A(n10865), .B(n7360), .Z(n2292) );
  XNOR U10636 ( .A(round_reg[1161]), .B(n9091), .Z(n7360) );
  ANDN U10637 ( .B(n8486), .A(n7359), .Z(n10865) );
  XOR U10638 ( .A(round_reg[778]), .B(n9393), .Z(n7359) );
  XOR U10639 ( .A(round_reg[416]), .B(n10226), .Z(n8486) );
  XOR U10640 ( .A(n3151), .B(n10866), .Z(n10862) );
  XOR U10641 ( .A(n5901), .B(n7349), .Z(n10866) );
  XNOR U10642 ( .A(n10867), .B(n7364), .Z(n7349) );
  XNOR U10643 ( .A(round_reg[1233]), .B(n10500), .Z(n7364) );
  AND U10644 ( .A(n8488), .B(n7365), .Z(n10867) );
  XOR U10645 ( .A(round_reg[875]), .B(n10868), .Z(n7365) );
  XNOR U10646 ( .A(round_reg[486]), .B(n10441), .Z(n8488) );
  XOR U10647 ( .A(n10869), .B(n7369), .Z(n5901) );
  XNOR U10648 ( .A(round_reg[1086]), .B(n10698), .Z(n7369) );
  ANDN U10649 ( .B(n10778), .A(n7368), .Z(n10869) );
  XNOR U10650 ( .A(n10870), .B(n7372), .Z(n3151) );
  XOR U10651 ( .A(round_reg[1135]), .B(n10871), .Z(n7372) );
  AND U10652 ( .A(n8483), .B(n7373), .Z(n10870) );
  XOR U10653 ( .A(round_reg[732]), .B(n10872), .Z(n7373) );
  XNOR U10654 ( .A(round_reg[365]), .B(n9837), .Z(n8483) );
  IV U10655 ( .A(n10873), .Z(n9837) );
  XOR U10656 ( .A(n10874), .B(n10875), .Z(n6099) );
  XNOR U10657 ( .A(n5264), .B(n1902), .Z(n10875) );
  XNOR U10658 ( .A(n10876), .B(n8556), .Z(n1902) );
  ANDN U10659 ( .B(n7442), .A(n8471), .Z(n10876) );
  XNOR U10660 ( .A(round_reg[290]), .B(n9099), .Z(n8471) );
  XOR U10661 ( .A(round_reg[1523]), .B(n10752), .Z(n7442) );
  XNOR U10662 ( .A(n10877), .B(n8562), .Z(n5264) );
  ANDN U10663 ( .B(n8468), .A(n7434), .Z(n10877) );
  XOR U10664 ( .A(round_reg[1305]), .B(n9934), .Z(n7434) );
  XNOR U10665 ( .A(round_reg[124]), .B(n10878), .Z(n8468) );
  XNOR U10666 ( .A(n3663), .B(n10879), .Z(n10874) );
  XOR U10667 ( .A(n8537), .B(n4112), .Z(n10879) );
  XNOR U10668 ( .A(n10880), .B(n8564), .Z(n4112) );
  NOR U10669 ( .A(n8478), .B(n7425), .Z(n10880) );
  XNOR U10670 ( .A(round_reg[1368]), .B(n10881), .Z(n7425) );
  XNOR U10671 ( .A(round_reg[183]), .B(n10211), .Z(n8478) );
  XNOR U10672 ( .A(n10882), .B(n8559), .Z(n8537) );
  AND U10673 ( .A(n7429), .B(n8560), .Z(n10882) );
  XNOR U10674 ( .A(round_reg[38]), .B(n10883), .Z(n8560) );
  XNOR U10675 ( .A(round_reg[1588]), .B(n9459), .Z(n7429) );
  XNOR U10676 ( .A(n10884), .B(n10885), .Z(n3663) );
  AND U10677 ( .A(n7438), .B(n8476), .Z(n10884) );
  XNOR U10678 ( .A(round_reg[1462]), .B(n10296), .Z(n7438) );
  XOR U10679 ( .A(n10886), .B(n7368), .Z(n8481) );
  XNOR U10680 ( .A(round_reg[654]), .B(n9981), .Z(n7368) );
  ANDN U10681 ( .B(n8422), .A(n10778), .Z(n10886) );
  XOR U10682 ( .A(round_reg[588]), .B(n10887), .Z(n10778) );
  XOR U10683 ( .A(round_reg[243]), .B(n10752), .Z(n8422) );
  ANDN U10684 ( .B(n5680), .A(n5678), .Z(n10861) );
  XNOR U10685 ( .A(n10888), .B(n1742), .Z(n5678) );
  XOR U10686 ( .A(n10889), .B(n10890), .Z(n9398) );
  XNOR U10687 ( .A(n3462), .B(n5083), .Z(n10890) );
  XOR U10688 ( .A(n10891), .B(n8395), .Z(n5083) );
  ANDN U10689 ( .B(n10824), .A(n8394), .Z(n10891) );
  XNOR U10690 ( .A(n10892), .B(n9480), .Z(n3462) );
  NOR U10691 ( .A(n10827), .B(n9479), .Z(n10892) );
  XNOR U10692 ( .A(n4185), .B(n10893), .Z(n10889) );
  XOR U10693 ( .A(n8384), .B(n2485), .Z(n10893) );
  XNOR U10694 ( .A(n10894), .B(n8405), .Z(n2485) );
  AND U10695 ( .A(n10895), .B(n8404), .Z(n10894) );
  XOR U10696 ( .A(n10896), .B(n10897), .Z(n8384) );
  AND U10697 ( .A(n10819), .B(n8391), .Z(n10896) );
  XNOR U10698 ( .A(n10898), .B(n8401), .Z(n4185) );
  NOR U10699 ( .A(n10816), .B(n8400), .Z(n10898) );
  XNOR U10700 ( .A(n10899), .B(n10900), .Z(n6354) );
  XNOR U10701 ( .A(n5438), .B(n3649), .Z(n10900) );
  XOR U10702 ( .A(n10901), .B(n10902), .Z(n3649) );
  ANDN U10703 ( .B(n10903), .A(n8452), .Z(n10901) );
  XNOR U10704 ( .A(n10904), .B(n10905), .Z(n5438) );
  ANDN U10705 ( .B(n8442), .A(n10906), .Z(n10904) );
  XNOR U10706 ( .A(n10907), .B(n10908), .Z(n10899) );
  XOR U10707 ( .A(n2107), .B(n4238), .Z(n10908) );
  XNOR U10708 ( .A(n10909), .B(n10910), .Z(n4238) );
  ANDN U10709 ( .B(n8446), .A(n10911), .Z(n10909) );
  XOR U10710 ( .A(n10912), .B(n10913), .Z(n2107) );
  NOR U10711 ( .A(n9561), .B(n10914), .Z(n10912) );
  XOR U10712 ( .A(n10184), .B(n5396), .Z(n5680) );
  XOR U10713 ( .A(n7822), .B(n8956), .Z(n5396) );
  XNOR U10714 ( .A(n10915), .B(n10916), .Z(n8956) );
  XOR U10715 ( .A(n5474), .B(n3848), .Z(n10916) );
  XOR U10716 ( .A(n10917), .B(n10918), .Z(n3848) );
  XNOR U10717 ( .A(round_reg[922]), .B(n9780), .Z(n7978) );
  XNOR U10718 ( .A(n10919), .B(n10235), .Z(n5474) );
  XNOR U10719 ( .A(round_reg[818]), .B(n10617), .Z(n7975) );
  XOR U10720 ( .A(round_reg[1201]), .B(n10920), .Z(n7973) );
  XOR U10721 ( .A(n6316), .B(n10921), .Z(n10915) );
  XOR U10722 ( .A(n2341), .B(n5277), .Z(n10921) );
  XOR U10723 ( .A(n10922), .B(n10246), .Z(n5277) );
  NOR U10724 ( .A(n8959), .B(n8958), .Z(n10922) );
  XOR U10725 ( .A(round_reg[1273]), .B(n10923), .Z(n8958) );
  XNOR U10726 ( .A(round_reg[851]), .B(n9907), .Z(n8959) );
  XNOR U10727 ( .A(n10924), .B(n10238), .Z(n2341) );
  XOR U10728 ( .A(round_reg[1062]), .B(n9776), .Z(n7963) );
  IV U10729 ( .A(n10006), .Z(n9776) );
  IV U10730 ( .A(n10343), .Z(n7964) );
  XOR U10731 ( .A(round_reg[694]), .B(n9198), .Z(n10343) );
  IV U10732 ( .A(n9630), .Z(n9198) );
  XOR U10733 ( .A(n10925), .B(n10243), .Z(n6316) );
  XNOR U10734 ( .A(round_reg[708]), .B(n10926), .Z(n7968) );
  XOR U10735 ( .A(round_reg[1111]), .B(n10927), .Z(n7967) );
  XOR U10736 ( .A(n10928), .B(n10929), .Z(n7822) );
  XOR U10737 ( .A(n3757), .B(n5124), .Z(n10929) );
  XOR U10738 ( .A(n10930), .B(n8900), .Z(n5124) );
  XOR U10739 ( .A(round_reg[463]), .B(n10931), .Z(n8900) );
  AND U10740 ( .A(n10191), .B(n10190), .Z(n10930) );
  XOR U10741 ( .A(round_reg[102]), .B(n10006), .Z(n10190) );
  XOR U10742 ( .A(n10932), .B(n10933), .Z(n10006) );
  XNOR U10743 ( .A(round_reg[1283]), .B(n9103), .Z(n10191) );
  XNOR U10744 ( .A(n10934), .B(n7895), .Z(n3757) );
  XNOR U10745 ( .A(round_reg[629]), .B(n10627), .Z(n7895) );
  NOR U10746 ( .A(n10182), .B(n10183), .Z(n10934) );
  XOR U10747 ( .A(round_reg[1440]), .B(n10935), .Z(n10183) );
  XNOR U10748 ( .A(round_reg[220]), .B(n10936), .Z(n10182) );
  XOR U10749 ( .A(n4178), .B(n10937), .Z(n10928) );
  XOR U10750 ( .A(n1699), .B(n10230), .Z(n10937) );
  XOR U10751 ( .A(n10938), .B(n7904), .Z(n10230) );
  XNOR U10752 ( .A(round_reg[393]), .B(n9916), .Z(n7904) );
  AND U10753 ( .A(n10180), .B(n10179), .Z(n10938) );
  XNOR U10754 ( .A(round_reg[16]), .B(n10939), .Z(n10179) );
  XNOR U10755 ( .A(round_reg[1566]), .B(n9473), .Z(n10180) );
  XNOR U10756 ( .A(n10940), .B(n7899), .Z(n1699) );
  XOR U10757 ( .A(round_reg[342]), .B(n9901), .Z(n7899) );
  AND U10758 ( .A(n10188), .B(n10187), .Z(n10940) );
  XOR U10759 ( .A(round_reg[268]), .B(n10941), .Z(n10187) );
  XNOR U10760 ( .A(round_reg[1501]), .B(n9260), .Z(n10188) );
  IV U10761 ( .A(n9199), .Z(n9260) );
  XOR U10762 ( .A(n10942), .B(n10943), .Z(n9199) );
  XNOR U10763 ( .A(n10944), .B(n7909), .Z(n4178) );
  XOR U10764 ( .A(round_reg[561]), .B(n10945), .Z(n7909) );
  NOR U10765 ( .A(n10253), .B(n10832), .Z(n10944) );
  XNOR U10766 ( .A(n10946), .B(n10253), .Z(n10184) );
  XNOR U10767 ( .A(round_reg[161]), .B(n10099), .Z(n10253) );
  AND U10768 ( .A(n10832), .B(n7907), .Z(n10946) );
  XOR U10769 ( .A(round_reg[970]), .B(n10947), .Z(n7907) );
  XOR U10770 ( .A(round_reg[1346]), .B(n10379), .Z(n10832) );
  XOR U10771 ( .A(n10948), .B(n4136), .Z(out[100]) );
  IV U10772 ( .A(n4308), .Z(n4136) );
  XOR U10773 ( .A(n7080), .B(n2592), .Z(n4308) );
  XNOR U10774 ( .A(n8096), .B(n10447), .Z(n2592) );
  XNOR U10775 ( .A(n10949), .B(n10950), .Z(n10447) );
  XNOR U10776 ( .A(n5743), .B(n5427), .Z(n10950) );
  XNOR U10777 ( .A(n10951), .B(n7097), .Z(n5427) );
  XNOR U10778 ( .A(round_reg[998]), .B(n10883), .Z(n7097) );
  ANDN U10779 ( .B(n8213), .A(n7096), .Z(n10951) );
  XNOR U10780 ( .A(round_reg[951]), .B(n10608), .Z(n7096) );
  XNOR U10781 ( .A(n10952), .B(n7106), .Z(n5743) );
  XOR U10782 ( .A(round_reg[1027]), .B(n10860), .Z(n7106) );
  ANDN U10783 ( .B(n10386), .A(n7105), .Z(n10952) );
  XNOR U10784 ( .A(round_reg[659]), .B(n10174), .Z(n7105) );
  XOR U10785 ( .A(round_reg[593]), .B(n10500), .Z(n10386) );
  XOR U10786 ( .A(n7090), .B(n10953), .Z(n10949) );
  XNOR U10787 ( .A(n2258), .B(n3379), .Z(n10953) );
  XNOR U10788 ( .A(n10954), .B(n7113), .Z(n3379) );
  XOR U10789 ( .A(round_reg[1140]), .B(n10955), .Z(n7113) );
  AND U10790 ( .A(n8205), .B(n7114), .Z(n10954) );
  XNOR U10791 ( .A(round_reg[737]), .B(n10140), .Z(n7114) );
  XNOR U10792 ( .A(round_reg[370]), .B(n9522), .Z(n8205) );
  XOR U10793 ( .A(n10956), .B(n7101), .Z(n2258) );
  XOR U10794 ( .A(round_reg[1166]), .B(n10957), .Z(n7101) );
  ANDN U10795 ( .B(n8208), .A(n7100), .Z(n10956) );
  XNOR U10796 ( .A(round_reg[783]), .B(n10931), .Z(n7100) );
  XOR U10797 ( .A(round_reg[421]), .B(n10958), .Z(n8208) );
  XNOR U10798 ( .A(n10959), .B(n7109), .Z(n7090) );
  XOR U10799 ( .A(round_reg[1238]), .B(n10960), .Z(n7109) );
  ANDN U10800 ( .B(n7110), .A(n8211), .Z(n10959) );
  XNOR U10801 ( .A(round_reg[491]), .B(n10047), .Z(n8211) );
  XOR U10802 ( .A(round_reg[880]), .B(n10961), .Z(n7110) );
  XOR U10803 ( .A(n10962), .B(n10963), .Z(n8096) );
  XNOR U10804 ( .A(n4314), .B(n2206), .Z(n10963) );
  XOR U10805 ( .A(n10964), .B(n8156), .Z(n2206) );
  XNOR U10806 ( .A(round_reg[67]), .B(n10860), .Z(n8156) );
  XOR U10807 ( .A(n10965), .B(n8148), .Z(n4314) );
  XNOR U10808 ( .A(round_reg[297]), .B(n9974), .Z(n8148) );
  XOR U10809 ( .A(round_reg[1141]), .B(n10662), .Z(n7087) );
  XNOR U10810 ( .A(round_reg[1530]), .B(n9685), .Z(n7086) );
  XOR U10811 ( .A(n6060), .B(n10966), .Z(n10962) );
  XOR U10812 ( .A(n5572), .B(n3759), .Z(n10966) );
  XNOR U10813 ( .A(n10967), .B(n8152), .Z(n3759) );
  XNOR U10814 ( .A(round_reg[45]), .B(n10873), .Z(n8152) );
  XOR U10815 ( .A(round_reg[1595]), .B(n10440), .Z(n7076) );
  XNOR U10816 ( .A(round_reg[1167]), .B(n10968), .Z(n7078) );
  XOR U10817 ( .A(n10969), .B(n10315), .Z(n5572) );
  XNOR U10818 ( .A(round_reg[249]), .B(n9758), .Z(n10315) );
  ANDN U10819 ( .B(n10366), .A(n7082), .Z(n10969) );
  XOR U10820 ( .A(round_reg[1469]), .B(n9961), .Z(n7082) );
  IV U10821 ( .A(n7084), .Z(n10366) );
  XOR U10822 ( .A(round_reg[1028]), .B(n10223), .Z(n7084) );
  XOR U10823 ( .A(n10970), .B(n8159), .Z(n6060) );
  XNOR U10824 ( .A(round_reg[190]), .B(n9688), .Z(n8159) );
  ANDN U10825 ( .B(n7072), .A(n7074), .Z(n10970) );
  XOR U10826 ( .A(round_reg[999]), .B(n10783), .Z(n7074) );
  XNOR U10827 ( .A(round_reg[1375]), .B(n10618), .Z(n7072) );
  XNOR U10828 ( .A(n10971), .B(n10309), .Z(n7080) );
  XOR U10829 ( .A(round_reg[1312]), .B(n10972), .Z(n10309) );
  ANDN U10830 ( .B(n10374), .A(n8155), .Z(n10971) );
  XOR U10831 ( .A(round_reg[881]), .B(n10945), .Z(n8155) );
  XNOR U10832 ( .A(round_reg[1239]), .B(n9935), .Z(n10374) );
  AND U10833 ( .A(n3638), .B(n3640), .Z(n10948) );
  XOR U10834 ( .A(n2366), .B(n9573), .Z(n3640) );
  XOR U10835 ( .A(n10973), .B(n10155), .Z(n9573) );
  NOR U10836 ( .A(n10271), .B(n9502), .Z(n10973) );
  XNOR U10837 ( .A(round_reg[24]), .B(n10020), .Z(n9502) );
  IV U10838 ( .A(n5002), .Z(n2366) );
  XOR U10839 ( .A(n6268), .B(n10345), .Z(n5002) );
  XOR U10840 ( .A(n10974), .B(n10975), .Z(n10345) );
  XOR U10841 ( .A(n1662), .B(n9645), .Z(n10975) );
  XOR U10842 ( .A(n10976), .B(n7414), .Z(n9645) );
  XOR U10843 ( .A(round_reg[400]), .B(n9447), .Z(n7414) );
  ANDN U10844 ( .B(n9585), .A(n9586), .Z(n10976) );
  XOR U10845 ( .A(round_reg[1573]), .B(n9263), .Z(n9586) );
  XOR U10846 ( .A(round_reg[23]), .B(n10977), .Z(n9585) );
  XNOR U10847 ( .A(n10978), .B(n7408), .Z(n1662) );
  XOR U10848 ( .A(round_reg[349]), .B(n9708), .Z(n7408) );
  AND U10849 ( .A(n9594), .B(n9593), .Z(n10978) );
  XNOR U10850 ( .A(round_reg[275]), .B(n10317), .Z(n9593) );
  XNOR U10851 ( .A(round_reg[1508]), .B(n10282), .Z(n9594) );
  XOR U10852 ( .A(n3728), .B(n10979), .Z(n10974) );
  XOR U10853 ( .A(n5102), .B(n4156), .Z(n10979) );
  XNOR U10854 ( .A(n10980), .B(n7418), .Z(n4156) );
  XOR U10855 ( .A(round_reg[568]), .B(n10351), .Z(n7418) );
  ANDN U10856 ( .B(n9655), .A(n10259), .Z(n10980) );
  XOR U10857 ( .A(round_reg[1353]), .B(n9916), .Z(n10259) );
  XNOR U10858 ( .A(round_reg[168]), .B(n10981), .Z(n9655) );
  XNOR U10859 ( .A(n10982), .B(n8410), .Z(n5102) );
  XOR U10860 ( .A(round_reg[470]), .B(n9841), .Z(n8410) );
  ANDN U10861 ( .B(n9588), .A(n9589), .Z(n10982) );
  XOR U10862 ( .A(round_reg[1290]), .B(n10983), .Z(n9589) );
  XNOR U10863 ( .A(round_reg[109]), .B(n10984), .Z(n9588) );
  XNOR U10864 ( .A(n10985), .B(n8653), .Z(n3728) );
  XOR U10865 ( .A(round_reg[636]), .B(n9993), .Z(n8653) );
  IV U10866 ( .A(n10667), .Z(n9993) );
  NOR U10867 ( .A(n9596), .B(n9597), .Z(n10985) );
  XOR U10868 ( .A(round_reg[1447]), .B(n10797), .Z(n9597) );
  XNOR U10869 ( .A(round_reg[227]), .B(n10433), .Z(n9596) );
  XOR U10870 ( .A(n10986), .B(n10987), .Z(n6268) );
  XOR U10871 ( .A(n3213), .B(n8017), .Z(n10987) );
  XOR U10872 ( .A(n10988), .B(n9518), .Z(n8017) );
  XOR U10873 ( .A(round_reg[1071]), .B(n9375), .Z(n9518) );
  ANDN U10874 ( .B(n9580), .A(n9581), .Z(n10988) );
  XOR U10875 ( .A(round_reg[637]), .B(n9906), .Z(n9581) );
  IV U10876 ( .A(n10592), .Z(n9906) );
  XNOR U10877 ( .A(round_reg[703]), .B(n9445), .Z(n9580) );
  XNOR U10878 ( .A(n10989), .B(n9514), .Z(n3213) );
  XOR U10879 ( .A(round_reg[1120]), .B(n10935), .Z(n9514) );
  ANDN U10880 ( .B(n9568), .A(n9569), .Z(n10989) );
  XOR U10881 ( .A(round_reg[350]), .B(n9635), .Z(n9569) );
  XNOR U10882 ( .A(round_reg[717]), .B(n10573), .Z(n9568) );
  XNOR U10883 ( .A(n10990), .B(n10991), .Z(n10573) );
  XOR U10884 ( .A(n5533), .B(n10992), .Z(n10986) );
  XOR U10885 ( .A(n8355), .B(n2403), .Z(n10992) );
  XNOR U10886 ( .A(n10993), .B(n9504), .Z(n2403) );
  XOR U10887 ( .A(round_reg[1210]), .B(n9685), .Z(n9504) );
  XOR U10888 ( .A(n10994), .B(n10995), .Z(n9685) );
  AND U10889 ( .A(n10271), .B(n10155), .Z(n10993) );
  XNOR U10890 ( .A(round_reg[827]), .B(n9195), .Z(n10155) );
  XNOR U10891 ( .A(n10996), .B(n10997), .Z(n9195) );
  XNOR U10892 ( .A(round_reg[401]), .B(n9829), .Z(n10271) );
  XNOR U10893 ( .A(n10998), .B(n9508), .Z(n8355) );
  XOR U10894 ( .A(round_reg[1218]), .B(n9603), .Z(n9508) );
  IV U10895 ( .A(n10999), .Z(n9603) );
  ANDN U10896 ( .B(n9571), .A(n9572), .Z(n10998) );
  XOR U10897 ( .A(round_reg[471]), .B(n11000), .Z(n9572) );
  XNOR U10898 ( .A(round_reg[860]), .B(n11001), .Z(n9571) );
  XNOR U10899 ( .A(n11002), .B(n10153), .Z(n5533) );
  XOR U10900 ( .A(round_reg[978]), .B(n10767), .Z(n10153) );
  ANDN U10901 ( .B(n9576), .A(n9578), .Z(n11002) );
  XOR U10902 ( .A(round_reg[569]), .B(n9758), .Z(n9578) );
  XNOR U10903 ( .A(round_reg[931]), .B(n11005), .Z(n9576) );
  XNOR U10904 ( .A(n7618), .B(n2434), .Z(n3638) );
  XNOR U10905 ( .A(n9937), .B(n10488), .Z(n2434) );
  XNOR U10906 ( .A(n11006), .B(n11007), .Z(n10488) );
  XNOR U10907 ( .A(n5443), .B(n3828), .Z(n11007) );
  XOR U10908 ( .A(n11008), .B(n10571), .Z(n3828) );
  XOR U10909 ( .A(round_reg[1350]), .B(n10012), .Z(n10571) );
  ANDN U10910 ( .B(n7630), .A(n7631), .Z(n11008) );
  XNOR U10911 ( .A(round_reg[927]), .B(n9396), .Z(n7631) );
  XOR U10912 ( .A(round_reg[974]), .B(n9981), .Z(n7630) );
  XNOR U10913 ( .A(n11009), .B(n9800), .Z(n5443) );
  XNOR U10914 ( .A(round_reg[1570]), .B(n9099), .Z(n9800) );
  IV U10915 ( .A(n10260), .Z(n9099) );
  XNOR U10916 ( .A(n11010), .B(n11011), .Z(n10260) );
  ANDN U10917 ( .B(n7626), .A(n7628), .Z(n11009) );
  XNOR U10918 ( .A(round_reg[823]), .B(n9531), .Z(n7628) );
  IV U10919 ( .A(n10211), .Z(n9531) );
  XOR U10920 ( .A(n11012), .B(n11013), .Z(n10211) );
  XOR U10921 ( .A(round_reg[1206]), .B(n9914), .Z(n7626) );
  IV U10922 ( .A(n10606), .Z(n9914) );
  XNOR U10923 ( .A(n11014), .B(n11015), .Z(n10606) );
  XOR U10924 ( .A(n6296), .B(n11016), .Z(n11006) );
  XOR U10925 ( .A(n2302), .B(n5113), .Z(n11016) );
  XNOR U10926 ( .A(n11017), .B(n9812), .Z(n5113) );
  XOR U10927 ( .A(round_reg[1287]), .B(n11018), .Z(n9812) );
  ANDN U10928 ( .B(n8656), .A(n8657), .Z(n11017) );
  XNOR U10929 ( .A(round_reg[856]), .B(n9602), .Z(n8657) );
  XOR U10930 ( .A(round_reg[1278]), .B(n9838), .Z(n8656) );
  XNOR U10931 ( .A(n11019), .B(n9804), .Z(n2302) );
  XOR U10932 ( .A(round_reg[1444]), .B(n9830), .Z(n9804) );
  ANDN U10933 ( .B(n10114), .A(n9803), .Z(n11019) );
  XNOR U10934 ( .A(n11020), .B(n9809), .Z(n6296) );
  XOR U10935 ( .A(round_reg[1505]), .B(n10496), .Z(n9809) );
  ANDN U10936 ( .B(n7620), .A(n7621), .Z(n11020) );
  XNOR U10937 ( .A(round_reg[713]), .B(n11021), .Z(n7621) );
  XOR U10938 ( .A(round_reg[1116]), .B(n9441), .Z(n7620) );
  XOR U10939 ( .A(n11022), .B(n11023), .Z(n9937) );
  XNOR U10940 ( .A(n3436), .B(n5024), .Z(n11023) );
  XNOR U10941 ( .A(n11024), .B(n7691), .Z(n5024) );
  XOR U10942 ( .A(round_reg[712]), .B(n9852), .Z(n7691) );
  ANDN U10943 ( .B(n7692), .A(n9879), .Z(n11024) );
  XNOR U10944 ( .A(round_reg[271]), .B(n11025), .Z(n9879) );
  XOR U10945 ( .A(round_reg[345]), .B(n9934), .Z(n7692) );
  XNOR U10946 ( .A(n11026), .B(n8715), .Z(n3436) );
  XOR U10947 ( .A(round_reg[855]), .B(n9752), .Z(n8715) );
  ANDN U10948 ( .B(n8716), .A(n9882), .Z(n11026) );
  XNOR U10949 ( .A(round_reg[105]), .B(n9552), .Z(n9882) );
  XOR U10950 ( .A(round_reg[466]), .B(n11027), .Z(n8716) );
  XOR U10951 ( .A(n2406), .B(n11028), .Z(n11022) );
  XOR U10952 ( .A(n7684), .B(n3938), .Z(n11028) );
  XOR U10953 ( .A(n11029), .B(n7705), .Z(n3938) );
  XOR U10954 ( .A(round_reg[822]), .B(n10296), .Z(n7705) );
  NOR U10955 ( .A(n7704), .B(n9871), .Z(n11029) );
  XNOR U10956 ( .A(round_reg[19]), .B(n11030), .Z(n9871) );
  XNOR U10957 ( .A(round_reg[396]), .B(n9621), .Z(n7704) );
  XOR U10958 ( .A(n11033), .B(n7700), .Z(n7684) );
  XOR U10959 ( .A(round_reg[698]), .B(n11034), .Z(n7700) );
  AND U10960 ( .A(n7701), .B(n9874), .Z(n11033) );
  XOR U10961 ( .A(round_reg[223]), .B(n9894), .Z(n9874) );
  XOR U10962 ( .A(round_reg[632]), .B(n9092), .Z(n7701) );
  XNOR U10963 ( .A(n11035), .B(n7696), .Z(n2406) );
  XOR U10964 ( .A(round_reg[926]), .B(n9473), .Z(n7696) );
  AND U10965 ( .A(n7697), .B(n10681), .Z(n11035) );
  XNOR U10966 ( .A(round_reg[164]), .B(n9830), .Z(n10681) );
  XOR U10967 ( .A(round_reg[564]), .B(n10781), .Z(n7697) );
  XOR U10968 ( .A(n11036), .B(n9803), .Z(n7618) );
  XOR U10969 ( .A(round_reg[1067]), .B(n9392), .Z(n9803) );
  XOR U10970 ( .A(n11037), .B(n11038), .Z(n9392) );
  NOR U10971 ( .A(n10115), .B(n10114), .Z(n11036) );
  XOR U10972 ( .A(round_reg[699]), .B(n9762), .Z(n10114) );
  XNOR U10973 ( .A(round_reg[633]), .B(n10923), .Z(n10115) );
  XOR U10974 ( .A(n11039), .B(n6234), .Z(out[1009]) );
  XOR U10975 ( .A(n8554), .B(n2263), .Z(n6234) );
  XNOR U10976 ( .A(n6110), .B(n6193), .Z(n2263) );
  XNOR U10977 ( .A(n11040), .B(n11041), .Z(n6193) );
  XNOR U10978 ( .A(n2299), .B(n5454), .Z(n11041) );
  XOR U10979 ( .A(n11042), .B(n7427), .Z(n5454) );
  XOR U10980 ( .A(round_reg[992]), .B(n9471), .Z(n7427) );
  ANDN U10981 ( .B(n8564), .A(n7426), .Z(n11042) );
  XNOR U10982 ( .A(round_reg[945]), .B(n9696), .Z(n7426) );
  XOR U10983 ( .A(round_reg[519]), .B(n11043), .Z(n8564) );
  XNOR U10984 ( .A(n11044), .B(n7431), .Z(n2299) );
  XNOR U10985 ( .A(round_reg[1160]), .B(n11045), .Z(n7431) );
  ANDN U10986 ( .B(n8559), .A(n7430), .Z(n11044) );
  XNOR U10987 ( .A(round_reg[777]), .B(n9469), .Z(n7430) );
  IV U10988 ( .A(n9383), .Z(n9469) );
  XOR U10989 ( .A(round_reg[415]), .B(n10618), .Z(n8559) );
  XOR U10990 ( .A(n3155), .B(n11046), .Z(n11040) );
  XOR U10991 ( .A(n5934), .B(n7420), .Z(n11046) );
  XOR U10992 ( .A(n11047), .B(n8469), .Z(n7420) );
  IV U10993 ( .A(n7435), .Z(n8469) );
  XOR U10994 ( .A(round_reg[1232]), .B(n10541), .Z(n7435) );
  AND U10995 ( .A(n8562), .B(n7436), .Z(n11047) );
  XOR U10996 ( .A(round_reg[874]), .B(n11048), .Z(n7436) );
  XNOR U10997 ( .A(round_reg[485]), .B(n10495), .Z(n8562) );
  XOR U10998 ( .A(n11049), .B(n7440), .Z(n5934) );
  XNOR U10999 ( .A(round_reg[1085]), .B(n10785), .Z(n7440) );
  ANDN U11000 ( .B(n10885), .A(n7439), .Z(n11049) );
  XNOR U11001 ( .A(n11050), .B(n7444), .Z(n3155) );
  XOR U11002 ( .A(round_reg[1134]), .B(n11051), .Z(n7444) );
  ANDN U11003 ( .B(n8556), .A(n7443), .Z(n11050) );
  XOR U11004 ( .A(round_reg[364]), .B(n9379), .Z(n8556) );
  XOR U11005 ( .A(n11052), .B(n11053), .Z(n6110) );
  XNOR U11006 ( .A(n5267), .B(n1907), .Z(n11053) );
  XNOR U11007 ( .A(n11054), .B(n8678), .Z(n1907) );
  ANDN U11008 ( .B(n7513), .A(n8544), .Z(n11054) );
  XNOR U11009 ( .A(round_reg[289]), .B(n9219), .Z(n8544) );
  XNOR U11010 ( .A(n11055), .B(n11056), .Z(n9219) );
  XNOR U11011 ( .A(round_reg[1522]), .B(n10304), .Z(n7513) );
  XNOR U11012 ( .A(n11057), .B(n8683), .Z(n5267) );
  NOR U11013 ( .A(n7505), .B(n8541), .Z(n11057) );
  XNOR U11014 ( .A(round_reg[123]), .B(n11058), .Z(n8541) );
  XNOR U11015 ( .A(round_reg[1304]), .B(n10020), .Z(n7505) );
  XNOR U11016 ( .A(n3667), .B(n11059), .Z(n11052) );
  XOR U11017 ( .A(n8659), .B(n4115), .Z(n11059) );
  XNOR U11018 ( .A(n11060), .B(n8685), .Z(n4115) );
  NOR U11019 ( .A(n7496), .B(n8551), .Z(n11060) );
  XNOR U11020 ( .A(round_reg[182]), .B(n10296), .Z(n8551) );
  IV U11021 ( .A(n9610), .Z(n10296) );
  XOR U11022 ( .A(n11061), .B(n11062), .Z(n9610) );
  XNOR U11023 ( .A(round_reg[1367]), .B(n11063), .Z(n7496) );
  XNOR U11024 ( .A(n11064), .B(n8681), .Z(n8659) );
  ANDN U11025 ( .B(n7500), .A(n8547), .Z(n11064) );
  XNOR U11026 ( .A(round_reg[37]), .B(n10534), .Z(n8547) );
  XNOR U11027 ( .A(round_reg[1587]), .B(n9544), .Z(n7500) );
  XNOR U11028 ( .A(n11065), .B(n11066), .Z(n3667) );
  AND U11029 ( .A(n7509), .B(n8549), .Z(n11065) );
  XNOR U11030 ( .A(round_reg[1461]), .B(n10662), .Z(n7509) );
  XOR U11031 ( .A(n11067), .B(n7439), .Z(n8554) );
  XNOR U11032 ( .A(round_reg[653]), .B(n10042), .Z(n7439) );
  NOR U11033 ( .A(n8476), .B(n10885), .Z(n11067) );
  XOR U11034 ( .A(round_reg[587]), .B(n11068), .Z(n10885) );
  XNOR U11035 ( .A(round_reg[242]), .B(n10834), .Z(n8476) );
  IV U11036 ( .A(n10304), .Z(n10834) );
  XOR U11037 ( .A(n11069), .B(n11070), .Z(n10304) );
  ANDN U11038 ( .B(n5684), .A(n5682), .Z(n11039) );
  XNOR U11039 ( .A(n11071), .B(n1747), .Z(n5682) );
  XOR U11040 ( .A(n11072), .B(n11073), .Z(n9475) );
  XNOR U11041 ( .A(n3464), .B(n5088), .Z(n11073) );
  XOR U11042 ( .A(n11074), .B(n8447), .Z(n5088) );
  AND U11043 ( .A(n10910), .B(n8448), .Z(n11074) );
  XOR U11044 ( .A(n11075), .B(n9562), .Z(n3464) );
  ANDN U11045 ( .B(n9563), .A(n10913), .Z(n11075) );
  XNOR U11046 ( .A(n4204), .B(n11076), .Z(n11072) );
  XOR U11047 ( .A(n8437), .B(n2494), .Z(n11076) );
  XNOR U11048 ( .A(n11077), .B(n8458), .Z(n2494) );
  AND U11049 ( .A(n11078), .B(n8457), .Z(n11077) );
  XNOR U11050 ( .A(n11079), .B(n8444), .Z(n8437) );
  AND U11051 ( .A(n10905), .B(n11080), .Z(n11079) );
  XNOR U11052 ( .A(n11081), .B(n8454), .Z(n4204) );
  ANDN U11053 ( .B(n11082), .A(n8453), .Z(n11081) );
  XNOR U11054 ( .A(n11083), .B(n11084), .Z(n6358) );
  XNOR U11055 ( .A(n5442), .B(n3653), .Z(n11084) );
  XOR U11056 ( .A(n11085), .B(n11086), .Z(n3653) );
  AND U11057 ( .A(n8505), .B(n11087), .Z(n11085) );
  XNOR U11058 ( .A(n11088), .B(n11089), .Z(n5442) );
  ANDN U11059 ( .B(n8495), .A(n11090), .Z(n11088) );
  XNOR U11060 ( .A(n11091), .B(n11092), .Z(n11083) );
  XOR U11061 ( .A(n2110), .B(n4240), .Z(n11092) );
  XNOR U11062 ( .A(n11093), .B(n11094), .Z(n4240) );
  AND U11063 ( .A(n8499), .B(n11095), .Z(n11093) );
  XOR U11064 ( .A(n11096), .B(n11097), .Z(n2110) );
  NOR U11065 ( .A(n9642), .B(n11098), .Z(n11096) );
  XOR U11066 ( .A(n10239), .B(n5401), .Z(n5684) );
  XOR U11067 ( .A(n7889), .B(n9015), .Z(n5401) );
  XNOR U11068 ( .A(n11099), .B(n11100), .Z(n9015) );
  XNOR U11069 ( .A(n5480), .B(n3852), .Z(n11100) );
  XOR U11070 ( .A(n11101), .B(n11102), .Z(n3852) );
  ANDN U11071 ( .B(n8066), .A(n8067), .Z(n11101) );
  XNOR U11072 ( .A(round_reg[921]), .B(n11103), .Z(n8067) );
  XNOR U11073 ( .A(n11104), .B(n10323), .Z(n5480) );
  ANDN U11074 ( .B(n8062), .A(n8064), .Z(n11104) );
  XNOR U11075 ( .A(round_reg[817]), .B(n9913), .Z(n8064) );
  XOR U11076 ( .A(round_reg[1200]), .B(n10961), .Z(n8062) );
  XNOR U11077 ( .A(n6324), .B(n11105), .Z(n11099) );
  XNOR U11078 ( .A(n2348), .B(n5314), .Z(n11105) );
  XNOR U11079 ( .A(n11106), .B(n10334), .Z(n5314) );
  ANDN U11080 ( .B(n9017), .A(n9019), .Z(n11106) );
  XNOR U11081 ( .A(round_reg[850]), .B(n9994), .Z(n9019) );
  IV U11082 ( .A(n11107), .Z(n9994) );
  XOR U11083 ( .A(round_reg[1272]), .B(n9092), .Z(n9017) );
  XNOR U11084 ( .A(n11109), .B(n11110), .Z(n11013) );
  XNOR U11085 ( .A(round_reg[1527]), .B(round_reg[1207]), .Z(n11110) );
  XOR U11086 ( .A(round_reg[247]), .B(n11111), .Z(n11109) );
  XOR U11087 ( .A(round_reg[887]), .B(round_reg[567]), .Z(n11111) );
  XNOR U11088 ( .A(n11112), .B(n10326), .Z(n2348) );
  AND U11089 ( .A(n8052), .B(n8053), .Z(n11112) );
  IV U11090 ( .A(n10414), .Z(n8053) );
  XOR U11091 ( .A(round_reg[693]), .B(n9257), .Z(n10414) );
  XOR U11092 ( .A(round_reg[1061]), .B(n11113), .Z(n8052) );
  XNOR U11093 ( .A(n11114), .B(n10331), .Z(n6324) );
  NOR U11094 ( .A(n8056), .B(n8057), .Z(n11114) );
  XNOR U11095 ( .A(round_reg[707]), .B(n11115), .Z(n8057) );
  XNOR U11096 ( .A(round_reg[1110]), .B(n9841), .Z(n8056) );
  XOR U11097 ( .A(n11116), .B(n11117), .Z(n7889) );
  XOR U11098 ( .A(n3761), .B(n5126), .Z(n11117) );
  XOR U11099 ( .A(n11118), .B(n8960), .Z(n5126) );
  XOR U11100 ( .A(round_reg[462]), .B(n10529), .Z(n8960) );
  AND U11101 ( .A(n10246), .B(n10245), .Z(n11118) );
  XOR U11102 ( .A(round_reg[101]), .B(n11113), .Z(n10245) );
  XOR U11103 ( .A(round_reg[1282]), .B(n9187), .Z(n10246) );
  XNOR U11104 ( .A(n11119), .B(n7965), .Z(n3761) );
  XNOR U11105 ( .A(round_reg[628]), .B(n10711), .Z(n7965) );
  IV U11106 ( .A(n9459), .Z(n10711) );
  ANDN U11107 ( .B(n10237), .A(n10238), .Z(n11119) );
  XOR U11108 ( .A(round_reg[1439]), .B(n9192), .Z(n10238) );
  XOR U11109 ( .A(round_reg[219]), .B(n10265), .Z(n10237) );
  XOR U11110 ( .A(n4186), .B(n11120), .Z(n11116) );
  XOR U11111 ( .A(n1704), .B(n10318), .Z(n11120) );
  XOR U11112 ( .A(n11121), .B(n7974), .Z(n10318) );
  XNOR U11113 ( .A(round_reg[392]), .B(n9852), .Z(n7974) );
  XOR U11114 ( .A(n11122), .B(n11123), .Z(n9852) );
  ANDN U11115 ( .B(n10234), .A(n10235), .Z(n11121) );
  XOR U11116 ( .A(round_reg[1565]), .B(n9556), .Z(n10235) );
  XNOR U11117 ( .A(n11124), .B(n7969), .Z(n1704) );
  XOR U11118 ( .A(round_reg[341]), .B(n9987), .Z(n7969) );
  AND U11119 ( .A(n10243), .B(n10242), .Z(n11124) );
  XOR U11120 ( .A(round_reg[267]), .B(n11125), .Z(n10242) );
  XNOR U11121 ( .A(round_reg[1500]), .B(n10936), .Z(n10243) );
  XNOR U11122 ( .A(n11126), .B(n7979), .Z(n4186) );
  XOR U11123 ( .A(round_reg[560]), .B(n10961), .Z(n7979) );
  NOR U11124 ( .A(n10341), .B(n10918), .Z(n11126) );
  XNOR U11125 ( .A(n11127), .B(n10341), .Z(n10239) );
  XNOR U11126 ( .A(round_reg[160]), .B(n10935), .Z(n10341) );
  IV U11127 ( .A(n9109), .Z(n10935) );
  AND U11128 ( .A(n10918), .B(n7977), .Z(n11127) );
  XOR U11129 ( .A(round_reg[969]), .B(n10438), .Z(n7977) );
  XOR U11130 ( .A(round_reg[1345]), .B(n10454), .Z(n10918) );
  XOR U11131 ( .A(n11128), .B(n6239), .Z(out[1008]) );
  XOR U11132 ( .A(n8676), .B(n2270), .Z(n6239) );
  XNOR U11133 ( .A(n6115), .B(n6198), .Z(n2270) );
  XNOR U11134 ( .A(n11129), .B(n11130), .Z(n6198) );
  XNOR U11135 ( .A(n2306), .B(n5459), .Z(n11130) );
  XNOR U11136 ( .A(n11131), .B(n7498), .Z(n5459) );
  XNOR U11137 ( .A(round_reg[991]), .B(n9554), .Z(n7498) );
  ANDN U11138 ( .B(n8685), .A(n7497), .Z(n11131) );
  XNOR U11139 ( .A(round_reg[944]), .B(n9769), .Z(n7497) );
  XOR U11140 ( .A(round_reg[518]), .B(n9386), .Z(n8685) );
  XNOR U11141 ( .A(n11132), .B(n7502), .Z(n2306) );
  XNOR U11142 ( .A(round_reg[1159]), .B(n11133), .Z(n7502) );
  ANDN U11143 ( .B(n8681), .A(n7501), .Z(n11132) );
  XOR U11144 ( .A(round_reg[776]), .B(n9463), .Z(n7501) );
  XOR U11145 ( .A(round_reg[414]), .B(n10382), .Z(n8681) );
  XOR U11146 ( .A(n3163), .B(n11134), .Z(n11129) );
  XOR U11147 ( .A(n5989), .B(n7491), .Z(n11134) );
  XOR U11148 ( .A(n11135), .B(n8542), .Z(n7491) );
  IV U11149 ( .A(n7506), .Z(n8542) );
  XOR U11150 ( .A(round_reg[1231]), .B(n10630), .Z(n7506) );
  AND U11151 ( .A(n7507), .B(n8683), .Z(n11135) );
  XNOR U11152 ( .A(round_reg[484]), .B(n9830), .Z(n8683) );
  XOR U11153 ( .A(round_reg[873]), .B(n11136), .Z(n7507) );
  XOR U11154 ( .A(n11137), .B(n7511), .Z(n5989) );
  XNOR U11155 ( .A(round_reg[1084]), .B(n11138), .Z(n7511) );
  ANDN U11156 ( .B(n11066), .A(n7510), .Z(n11137) );
  XNOR U11157 ( .A(n11139), .B(n7515), .Z(n3163) );
  XOR U11158 ( .A(round_reg[1133]), .B(n11140), .Z(n7515) );
  ANDN U11159 ( .B(n8678), .A(n7514), .Z(n11139) );
  XNOR U11160 ( .A(round_reg[730]), .B(n11141), .Z(n7514) );
  XOR U11161 ( .A(round_reg[363]), .B(n9455), .Z(n8678) );
  XOR U11162 ( .A(n11142), .B(n11143), .Z(n6115) );
  XNOR U11163 ( .A(n5270), .B(n1915), .Z(n11143) );
  XNOR U11164 ( .A(n11144), .B(n8739), .Z(n1915) );
  ANDN U11165 ( .B(n7585), .A(n8665), .Z(n11144) );
  XNOR U11166 ( .A(round_reg[288]), .B(n9683), .Z(n8665) );
  IV U11167 ( .A(n10420), .Z(n9683) );
  XNOR U11168 ( .A(round_reg[1521]), .B(n10945), .Z(n7585) );
  XNOR U11169 ( .A(n11145), .B(n8744), .Z(n5270) );
  NOR U11170 ( .A(n7577), .B(n8663), .Z(n11145) );
  XNOR U11171 ( .A(round_reg[122]), .B(n11146), .Z(n8663) );
  XNOR U11172 ( .A(round_reg[1303]), .B(n10854), .Z(n7577) );
  XNOR U11173 ( .A(n3671), .B(n11147), .Z(n11142) );
  XOR U11174 ( .A(n8719), .B(n4118), .Z(n11147) );
  XNOR U11175 ( .A(n11148), .B(n8746), .Z(n4118) );
  NOR U11176 ( .A(n7568), .B(n8673), .Z(n11148) );
  XNOR U11177 ( .A(round_reg[181]), .B(n10662), .Z(n8673) );
  IV U11178 ( .A(n9684), .Z(n10662) );
  XNOR U11179 ( .A(round_reg[1366]), .B(n11151), .Z(n7568) );
  XNOR U11180 ( .A(n11152), .B(n8742), .Z(n8719) );
  ANDN U11181 ( .B(n7572), .A(n8669), .Z(n11152) );
  XNOR U11182 ( .A(round_reg[36]), .B(n10625), .Z(n8669) );
  IV U11183 ( .A(n9100), .Z(n10625) );
  XNOR U11184 ( .A(round_reg[1586]), .B(n9624), .Z(n7572) );
  XNOR U11185 ( .A(n11153), .B(n11154), .Z(n3671) );
  ANDN U11186 ( .B(n7581), .A(n8671), .Z(n11153) );
  XNOR U11187 ( .A(round_reg[1460]), .B(n10955), .Z(n7581) );
  XOR U11188 ( .A(n11155), .B(n7510), .Z(n8676) );
  XNOR U11189 ( .A(round_reg[652]), .B(n10168), .Z(n7510) );
  NOR U11190 ( .A(n8549), .B(n11066), .Z(n11155) );
  XOR U11191 ( .A(round_reg[586]), .B(n11156), .Z(n11066) );
  XNOR U11192 ( .A(round_reg[241]), .B(n10920), .Z(n8549) );
  IV U11193 ( .A(n10945), .Z(n10920) );
  XOR U11194 ( .A(n11157), .B(n11158), .Z(n10945) );
  NOR U11195 ( .A(n5687), .B(n5686), .Z(n11128) );
  XNOR U11196 ( .A(n11159), .B(n1752), .Z(n5686) );
  XOR U11197 ( .A(n11160), .B(n11161), .Z(n9558) );
  XNOR U11198 ( .A(n3470), .B(n4822), .Z(n11161) );
  XOR U11199 ( .A(n11162), .B(n8501), .Z(n4822) );
  ANDN U11200 ( .B(n11094), .A(n8500), .Z(n11162) );
  XNOR U11201 ( .A(n11163), .B(n9644), .Z(n3470) );
  NOR U11202 ( .A(n11097), .B(n9643), .Z(n11163) );
  XNOR U11203 ( .A(n4232), .B(n11164), .Z(n11160) );
  XOR U11204 ( .A(n8491), .B(n2501), .Z(n11164) );
  XNOR U11205 ( .A(n11165), .B(n8511), .Z(n2501) );
  AND U11206 ( .A(n11166), .B(n8510), .Z(n11165) );
  XNOR U11207 ( .A(n11167), .B(n8497), .Z(n8491) );
  AND U11208 ( .A(n11089), .B(n8496), .Z(n11167) );
  XNOR U11209 ( .A(n11168), .B(n8507), .Z(n4232) );
  ANDN U11210 ( .B(n11169), .A(n8506), .Z(n11168) );
  XNOR U11211 ( .A(n11170), .B(n11171), .Z(n6362) );
  XOR U11212 ( .A(n5447), .B(n3657), .Z(n11171) );
  XNOR U11213 ( .A(n11172), .B(n11173), .Z(n3657) );
  AND U11214 ( .A(n8578), .B(n11174), .Z(n11172) );
  XNOR U11215 ( .A(n11175), .B(n8520), .Z(n5447) );
  ANDN U11216 ( .B(n8521), .A(n8569), .Z(n11175) );
  XNOR U11217 ( .A(n4242), .B(n11176), .Z(n11170) );
  XOR U11218 ( .A(n5921), .B(n2115), .Z(n11176) );
  XOR U11219 ( .A(n11177), .B(n8516), .Z(n2115) );
  ANDN U11220 ( .B(n8517), .A(n9715), .Z(n11177) );
  XOR U11221 ( .A(n11178), .B(n8530), .Z(n5921) );
  ANDN U11222 ( .B(n8531), .A(n8582), .Z(n11178) );
  XOR U11223 ( .A(n11179), .B(n8526), .Z(n4242) );
  AND U11224 ( .A(n8573), .B(n8527), .Z(n11179) );
  XOR U11225 ( .A(n10327), .B(n2080), .Z(n5687) );
  XNOR U11226 ( .A(n7959), .B(n9069), .Z(n2080) );
  XNOR U11227 ( .A(n11180), .B(n11181), .Z(n9069) );
  XNOR U11228 ( .A(n5485), .B(n3577), .Z(n11181) );
  XOR U11229 ( .A(n11182), .B(n11183), .Z(n3577) );
  ANDN U11230 ( .B(n8133), .A(n8134), .Z(n11182) );
  XNOR U11231 ( .A(round_reg[920]), .B(n11184), .Z(n8134) );
  XNOR U11232 ( .A(n11185), .B(n10394), .Z(n5485) );
  ANDN U11233 ( .B(n8129), .A(n8131), .Z(n11185) );
  XNOR U11234 ( .A(round_reg[816]), .B(n10001), .Z(n8131) );
  XOR U11235 ( .A(round_reg[1199]), .B(n10532), .Z(n8129) );
  XNOR U11236 ( .A(n6328), .B(n11186), .Z(n11180) );
  XOR U11237 ( .A(n2355), .B(n5369), .Z(n11186) );
  XNOR U11238 ( .A(n11187), .B(n10405), .Z(n5369) );
  AND U11239 ( .A(n9073), .B(n9071), .Z(n11187) );
  XOR U11240 ( .A(round_reg[1271]), .B(n10608), .Z(n9071) );
  XNOR U11241 ( .A(round_reg[849]), .B(n10214), .Z(n9073) );
  XNOR U11242 ( .A(n11188), .B(n10397), .Z(n2355) );
  ANDN U11243 ( .B(n8121), .A(n8119), .Z(n11188) );
  XNOR U11244 ( .A(round_reg[1060]), .B(n10528), .Z(n8119) );
  XOR U11245 ( .A(round_reg[692]), .B(n11189), .Z(n8121) );
  XNOR U11246 ( .A(n11190), .B(n10402), .Z(n6328) );
  NOR U11247 ( .A(n8123), .B(n8124), .Z(n11190) );
  XNOR U11248 ( .A(round_reg[706]), .B(n10522), .Z(n8124) );
  XNOR U11249 ( .A(round_reg[1109]), .B(n9910), .Z(n8123) );
  XOR U11250 ( .A(n11191), .B(n11192), .Z(n7959) );
  XNOR U11251 ( .A(n3765), .B(n5128), .Z(n11192) );
  XOR U11252 ( .A(n11193), .B(n9018), .Z(n5128) );
  XNOR U11253 ( .A(round_reg[461]), .B(n11194), .Z(n9018) );
  AND U11254 ( .A(n10334), .B(n10333), .Z(n11193) );
  XNOR U11255 ( .A(round_reg[100]), .B(n9863), .Z(n10333) );
  IV U11256 ( .A(n10528), .Z(n9863) );
  XOR U11257 ( .A(round_reg[1281]), .B(n9966), .Z(n10334) );
  XNOR U11258 ( .A(n11195), .B(n8054), .Z(n3765) );
  XNOR U11259 ( .A(round_reg[627]), .B(n11196), .Z(n8054) );
  NOR U11260 ( .A(n10325), .B(n10326), .Z(n11195) );
  XOR U11261 ( .A(round_reg[1438]), .B(n10357), .Z(n10326) );
  XNOR U11262 ( .A(round_reg[218]), .B(n9526), .Z(n10325) );
  XOR U11263 ( .A(n4205), .B(n11197), .Z(n11191) );
  XOR U11264 ( .A(n1709), .B(n10389), .Z(n11197) );
  XOR U11265 ( .A(n11198), .B(n8063), .Z(n10389) );
  XNOR U11266 ( .A(round_reg[391]), .B(n9925), .Z(n8063) );
  AND U11267 ( .A(n10323), .B(n10322), .Z(n11198) );
  XNOR U11268 ( .A(round_reg[14]), .B(n11199), .Z(n10322) );
  XOR U11269 ( .A(round_reg[1564]), .B(n9637), .Z(n10323) );
  XNOR U11270 ( .A(n11200), .B(n8058), .Z(n1709) );
  XOR U11271 ( .A(round_reg[340]), .B(n10048), .Z(n8058) );
  AND U11272 ( .A(n10331), .B(n10330), .Z(n11200) );
  XOR U11273 ( .A(round_reg[266]), .B(n9087), .Z(n10330) );
  XNOR U11274 ( .A(round_reg[1499]), .B(n10265), .Z(n10331) );
  XOR U11275 ( .A(n11201), .B(n11202), .Z(n10265) );
  XNOR U11276 ( .A(n11203), .B(n8068), .Z(n4205) );
  XOR U11277 ( .A(round_reg[559]), .B(n10532), .Z(n8068) );
  NOR U11278 ( .A(n10412), .B(n11102), .Z(n11203) );
  XNOR U11279 ( .A(n11204), .B(n10412), .Z(n10327) );
  XNOR U11280 ( .A(round_reg[159]), .B(n9192), .Z(n10412) );
  IV U11281 ( .A(n11205), .Z(n9192) );
  ANDN U11282 ( .B(n11102), .A(n8066), .Z(n11204) );
  XOR U11283 ( .A(round_reg[968]), .B(n10492), .Z(n8066) );
  XOR U11284 ( .A(round_reg[1344]), .B(n10518), .Z(n11102) );
  XOR U11285 ( .A(n11206), .B(n6244), .Z(out[1007]) );
  XOR U11286 ( .A(n8737), .B(n2277), .Z(n6244) );
  XNOR U11287 ( .A(n6121), .B(n6203), .Z(n2277) );
  XNOR U11288 ( .A(n11207), .B(n11208), .Z(n6203) );
  XNOR U11289 ( .A(n2313), .B(n5463), .Z(n11208) );
  XNOR U11290 ( .A(n11209), .B(n7570), .Z(n5463) );
  XNOR U11291 ( .A(round_reg[990]), .B(n9635), .Z(n7570) );
  ANDN U11292 ( .B(n8746), .A(n7569), .Z(n11209) );
  XOR U11293 ( .A(round_reg[943]), .B(n11210), .Z(n7569) );
  XOR U11294 ( .A(round_reg[517]), .B(n9458), .Z(n8746) );
  XNOR U11295 ( .A(n11211), .B(n7574), .Z(n2313) );
  XNOR U11296 ( .A(round_reg[1158]), .B(n11212), .Z(n7574) );
  ANDN U11297 ( .B(n8742), .A(n7573), .Z(n11211) );
  XNOR U11298 ( .A(round_reg[775]), .B(n9633), .Z(n7573) );
  XOR U11299 ( .A(round_reg[413]), .B(n10457), .Z(n8742) );
  XOR U11300 ( .A(n3167), .B(n11213), .Z(n11207) );
  XNOR U11301 ( .A(n6047), .B(n7563), .Z(n11213) );
  XNOR U11302 ( .A(n11214), .B(n7579), .Z(n7563) );
  XNOR U11303 ( .A(round_reg[1230]), .B(n10713), .Z(n7579) );
  ANDN U11304 ( .B(n8744), .A(n7578), .Z(n11214) );
  XNOR U11305 ( .A(round_reg[872]), .B(n9977), .Z(n7578) );
  XOR U11306 ( .A(round_reg[483]), .B(n9899), .Z(n8744) );
  XOR U11307 ( .A(n11215), .B(n7583), .Z(n6047) );
  XNOR U11308 ( .A(round_reg[1083]), .B(n11058), .Z(n7583) );
  ANDN U11309 ( .B(n11154), .A(n7582), .Z(n11215) );
  XOR U11310 ( .A(n11216), .B(n8666), .Z(n3167) );
  XOR U11311 ( .A(round_reg[1132]), .B(n9986), .Z(n8666) );
  ANDN U11312 ( .B(n8739), .A(n7586), .Z(n11216) );
  XOR U11313 ( .A(round_reg[729]), .B(n10776), .Z(n7586) );
  XOR U11314 ( .A(round_reg[362]), .B(n9540), .Z(n8739) );
  XOR U11315 ( .A(n11217), .B(n11218), .Z(n6121) );
  XNOR U11316 ( .A(n5273), .B(n1920), .Z(n11218) );
  XNOR U11317 ( .A(n11219), .B(n8800), .Z(n1920) );
  NOR U11318 ( .A(n7656), .B(n8725), .Z(n11219) );
  XNOR U11319 ( .A(round_reg[287]), .B(n9756), .Z(n8725) );
  IV U11320 ( .A(n9396), .Z(n9756) );
  XNOR U11321 ( .A(n11220), .B(n11221), .Z(n9396) );
  XOR U11322 ( .A(round_reg[1520]), .B(n10961), .Z(n7656) );
  XNOR U11323 ( .A(n11222), .B(n8805), .Z(n5273) );
  NOR U11324 ( .A(n7648), .B(n8723), .Z(n11222) );
  XNOR U11325 ( .A(round_reg[121]), .B(n11223), .Z(n8723) );
  XOR U11326 ( .A(round_reg[1302]), .B(n9901), .Z(n7648) );
  XNOR U11327 ( .A(n3675), .B(n11224), .Z(n11217) );
  XOR U11328 ( .A(n8780), .B(n4121), .Z(n11224) );
  XNOR U11329 ( .A(n11225), .B(n8807), .Z(n4121) );
  NOR U11330 ( .A(n7639), .B(n8733), .Z(n11225) );
  XNOR U11331 ( .A(round_reg[180]), .B(n10955), .Z(n8733) );
  IV U11332 ( .A(n9757), .Z(n10955) );
  XNOR U11333 ( .A(n11226), .B(n11227), .Z(n9757) );
  XOR U11334 ( .A(round_reg[1365]), .B(n11228), .Z(n7639) );
  XNOR U11335 ( .A(n11229), .B(n8803), .Z(n8780) );
  AND U11336 ( .A(n7643), .B(n8729), .Z(n11229) );
  XNOR U11337 ( .A(round_reg[35]), .B(n11230), .Z(n8729) );
  XNOR U11338 ( .A(round_reg[1585]), .B(n9696), .Z(n7643) );
  XNOR U11339 ( .A(n11231), .B(n11232), .Z(n3675) );
  ANDN U11340 ( .B(n8731), .A(n7652), .Z(n11231) );
  XNOR U11341 ( .A(round_reg[1459]), .B(n10524), .Z(n7652) );
  XOR U11342 ( .A(n11233), .B(n7582), .Z(n8737) );
  XNOR U11343 ( .A(round_reg[651]), .B(n10277), .Z(n7582) );
  ANDN U11344 ( .B(n8671), .A(n11154), .Z(n11233) );
  XOR U11345 ( .A(round_reg[585]), .B(n11234), .Z(n11154) );
  XNOR U11346 ( .A(round_reg[240]), .B(n10961), .Z(n8671) );
  XNOR U11347 ( .A(n11235), .B(n11236), .Z(n10961) );
  NOR U11348 ( .A(n5691), .B(n5690), .Z(n11206) );
  XNOR U11349 ( .A(n8523), .B(n1757), .Z(n5690) );
  XOR U11350 ( .A(n11237), .B(n11238), .Z(n9639) );
  XNOR U11351 ( .A(n3472), .B(n4827), .Z(n11238) );
  XOR U11352 ( .A(n11239), .B(n8574), .Z(n4827) );
  ANDN U11353 ( .B(n8525), .A(n8526), .Z(n11239) );
  XNOR U11354 ( .A(round_reg[257]), .B(n11240), .Z(n8526) );
  XOR U11355 ( .A(round_reg[331]), .B(n10277), .Z(n8525) );
  IV U11356 ( .A(n10859), .Z(n10277) );
  XNOR U11357 ( .A(n11241), .B(n9716), .Z(n3472) );
  NOR U11358 ( .A(n8516), .B(n8515), .Z(n11241) );
  XNOR U11359 ( .A(round_reg[452]), .B(n11242), .Z(n8515) );
  XNOR U11360 ( .A(round_reg[91]), .B(n10601), .Z(n8516) );
  XNOR U11361 ( .A(n4258), .B(n11243), .Z(n11237) );
  XOR U11362 ( .A(n8565), .B(n2506), .Z(n11243) );
  XNOR U11363 ( .A(n11244), .B(n8583), .Z(n2506) );
  ANDN U11364 ( .B(n8529), .A(n8530), .Z(n11244) );
  XNOR U11365 ( .A(round_reg[150]), .B(n11245), .Z(n8530) );
  XOR U11366 ( .A(round_reg[550]), .B(n10045), .Z(n8529) );
  XOR U11367 ( .A(n11246), .B(n8570), .Z(n8565) );
  IV U11368 ( .A(n11247), .Z(n8570) );
  ANDN U11369 ( .B(n8571), .A(n8520), .Z(n11246) );
  XOR U11370 ( .A(round_reg[209]), .B(n10214), .Z(n8520) );
  XNOR U11371 ( .A(round_reg[618]), .B(n10220), .Z(n8571) );
  XNOR U11372 ( .A(n11248), .B(n8580), .Z(n4258) );
  AND U11373 ( .A(n11173), .B(n8579), .Z(n11248) );
  XNOR U11374 ( .A(n11249), .B(n11250), .Z(n6370) );
  XNOR U11375 ( .A(n5453), .B(n3661), .Z(n11250) );
  XNOR U11376 ( .A(n11251), .B(n11252), .Z(n3661) );
  ANDN U11377 ( .B(n6472), .A(n6473), .Z(n11251) );
  XOR U11378 ( .A(round_reg[1190]), .B(n10045), .Z(n6473) );
  XNOR U11379 ( .A(n11253), .B(n8591), .Z(n5453) );
  ANDN U11380 ( .B(n6463), .A(n6464), .Z(n11253) );
  XNOR U11381 ( .A(round_reg[1051]), .B(n10601), .Z(n6464) );
  XOR U11382 ( .A(round_reg[1428]), .B(n9997), .Z(n6463) );
  XOR U11383 ( .A(n4245), .B(n11254), .Z(n11249) );
  XNOR U11384 ( .A(n5926), .B(n2119), .Z(n11254) );
  XNOR U11385 ( .A(n11255), .B(n8588), .Z(n2119) );
  ANDN U11386 ( .B(n6476), .A(n6477), .Z(n11255) );
  XNOR U11387 ( .A(round_reg[1262]), .B(n9855), .Z(n6477) );
  XOR U11388 ( .A(round_reg[1335]), .B(n9550), .Z(n6476) );
  XOR U11389 ( .A(n11256), .B(n8599), .Z(n5926) );
  ANDN U11390 ( .B(n6480), .A(n6481), .Z(n11256) );
  XNOR U11391 ( .A(round_reg[1022]), .B(n9536), .Z(n6481) );
  XOR U11392 ( .A(round_reg[1398]), .B(n9108), .Z(n6480) );
  XNOR U11393 ( .A(n11257), .B(n8596), .Z(n4245) );
  ANDN U11394 ( .B(n6467), .A(n6468), .Z(n11257) );
  XNOR U11395 ( .A(round_reg[1100]), .B(n10705), .Z(n6468) );
  XOR U11396 ( .A(round_reg[1489]), .B(n10214), .Z(n6467) );
  IV U11397 ( .A(n10124), .Z(n10214) );
  XNOR U11398 ( .A(n11258), .B(n11259), .Z(n10124) );
  XNOR U11399 ( .A(n11260), .B(n8579), .Z(n8523) );
  XNOR U11400 ( .A(round_reg[446]), .B(n11261), .Z(n8579) );
  NOR U11401 ( .A(n11173), .B(n11174), .Z(n11260) );
  XNOR U11402 ( .A(round_reg[5]), .B(n10763), .Z(n11173) );
  XOR U11403 ( .A(n10398), .B(n2087), .Z(n5691) );
  XNOR U11404 ( .A(n8048), .B(n9145), .Z(n2087) );
  XNOR U11405 ( .A(n11262), .B(n11263), .Z(n9145) );
  XNOR U11406 ( .A(n5490), .B(n3581), .Z(n11263) );
  XOR U11407 ( .A(n11264), .B(n11265), .Z(n3581) );
  ANDN U11408 ( .B(n8193), .A(n8194), .Z(n11264) );
  XNOR U11409 ( .A(round_reg[919]), .B(n9935), .Z(n8194) );
  XNOR U11410 ( .A(n11266), .B(n10467), .Z(n5490) );
  ANDN U11411 ( .B(n8189), .A(n8191), .Z(n11266) );
  XNOR U11412 ( .A(round_reg[815]), .B(n10129), .Z(n8191) );
  XOR U11413 ( .A(round_reg[1198]), .B(n11267), .Z(n8189) );
  XNOR U11414 ( .A(n6332), .B(n11268), .Z(n11262) );
  XNOR U11415 ( .A(n2362), .B(n5418), .Z(n11268) );
  XNOR U11416 ( .A(n11269), .B(n10478), .Z(n5418) );
  AND U11417 ( .A(n9149), .B(n9147), .Z(n11269) );
  XOR U11418 ( .A(round_reg[1270]), .B(n10696), .Z(n9147) );
  XNOR U11419 ( .A(round_reg[848]), .B(n10299), .Z(n9149) );
  XNOR U11420 ( .A(n11270), .B(n10470), .Z(n2362) );
  ANDN U11421 ( .B(n8181), .A(n8179), .Z(n11270) );
  XNOR U11422 ( .A(round_reg[1059]), .B(n9928), .Z(n8179) );
  XOR U11423 ( .A(round_reg[691]), .B(n9437), .Z(n8181) );
  XNOR U11424 ( .A(n11271), .B(n10475), .Z(n6332) );
  ANDN U11425 ( .B(n8185), .A(n8183), .Z(n11271) );
  XNOR U11426 ( .A(round_reg[1108]), .B(n9997), .Z(n8183) );
  XOR U11427 ( .A(round_reg[705]), .B(n10615), .Z(n8185) );
  XOR U11428 ( .A(n11272), .B(n11273), .Z(n8048) );
  XNOR U11429 ( .A(n3772), .B(n5130), .Z(n11273) );
  XOR U11430 ( .A(n11274), .B(n9072), .Z(n5130) );
  XNOR U11431 ( .A(round_reg[460]), .B(n9083), .Z(n9072) );
  ANDN U11432 ( .B(n10404), .A(n10405), .Z(n11274) );
  XOR U11433 ( .A(round_reg[1280]), .B(n11275), .Z(n10405) );
  XOR U11434 ( .A(round_reg[99]), .B(n9928), .Z(n10404) );
  XOR U11435 ( .A(n11010), .B(n11276), .Z(n9928) );
  XOR U11436 ( .A(n11277), .B(n11278), .Z(n11010) );
  XNOR U11437 ( .A(round_reg[34]), .B(round_reg[1314]), .Z(n11278) );
  XOR U11438 ( .A(round_reg[354]), .B(n11279), .Z(n11277) );
  XOR U11439 ( .A(round_reg[994]), .B(round_reg[674]), .Z(n11279) );
  XNOR U11440 ( .A(n11280), .B(n8120), .Z(n3772) );
  XNOR U11441 ( .A(round_reg[626]), .B(n11281), .Z(n8120) );
  NOR U11442 ( .A(n10396), .B(n10397), .Z(n11280) );
  XNOR U11443 ( .A(round_reg[1437]), .B(n9367), .Z(n10397) );
  XNOR U11444 ( .A(round_reg[217]), .B(n9605), .Z(n10396) );
  XOR U11445 ( .A(n4233), .B(n11282), .Z(n11272) );
  XOR U11446 ( .A(n1714), .B(n10462), .Z(n11282) );
  XOR U11447 ( .A(n11283), .B(n8130), .Z(n10462) );
  XNOR U11448 ( .A(round_reg[390]), .B(n10012), .Z(n8130) );
  IV U11449 ( .A(n10758), .Z(n10012) );
  XNOR U11450 ( .A(n11284), .B(n11285), .Z(n10758) );
  AND U11451 ( .A(n10394), .B(n10393), .Z(n11283) );
  XNOR U11452 ( .A(round_reg[13]), .B(n10683), .Z(n10393) );
  IV U11453 ( .A(n10042), .Z(n10683) );
  XNOR U11454 ( .A(round_reg[1563]), .B(n10000), .Z(n10394) );
  XNOR U11455 ( .A(n11286), .B(n8125), .Z(n1714) );
  XOR U11456 ( .A(round_reg[339]), .B(n10174), .Z(n8125) );
  AND U11457 ( .A(n10402), .B(n10401), .Z(n11286) );
  XOR U11458 ( .A(round_reg[265]), .B(n9216), .Z(n10401) );
  XNOR U11459 ( .A(round_reg[1498]), .B(n9526), .Z(n10402) );
  IV U11460 ( .A(n9438), .Z(n9526) );
  XNOR U11461 ( .A(n11287), .B(n11288), .Z(n9438) );
  XNOR U11462 ( .A(n11289), .B(n8135), .Z(n4233) );
  XOR U11463 ( .A(round_reg[558]), .B(n11267), .Z(n8135) );
  NOR U11464 ( .A(n10485), .B(n11183), .Z(n11289) );
  XNOR U11465 ( .A(n11290), .B(n10485), .Z(n10398) );
  XNOR U11466 ( .A(round_reg[158]), .B(n10357), .Z(n10485) );
  ANDN U11467 ( .B(n11183), .A(n8133), .Z(n11290) );
  XOR U11468 ( .A(round_reg[967]), .B(n11018), .Z(n8133) );
  XOR U11469 ( .A(round_reg[1407]), .B(n10611), .Z(n11183) );
  XOR U11470 ( .A(n11291), .B(n6249), .Z(out[1006]) );
  XOR U11471 ( .A(n8798), .B(n2284), .Z(n6249) );
  XNOR U11472 ( .A(n6127), .B(n6208), .Z(n2284) );
  XNOR U11473 ( .A(n11292), .B(n11293), .Z(n6208) );
  XOR U11474 ( .A(n2320), .B(n5473), .Z(n11293) );
  XOR U11475 ( .A(n11294), .B(n8734), .Z(n5473) );
  IV U11476 ( .A(n7640), .Z(n8734) );
  XOR U11477 ( .A(round_reg[989]), .B(n9708), .Z(n7640) );
  AND U11478 ( .A(n8807), .B(n7641), .Z(n11294) );
  XOR U11479 ( .A(round_reg[942]), .B(n11295), .Z(n7641) );
  XNOR U11480 ( .A(round_reg[516]), .B(n9555), .Z(n8807) );
  XNOR U11481 ( .A(n11296), .B(n7645), .Z(n2320) );
  XNOR U11482 ( .A(round_reg[1157]), .B(n9472), .Z(n7645) );
  ANDN U11483 ( .B(n8803), .A(n7644), .Z(n11296) );
  XNOR U11484 ( .A(round_reg[774]), .B(n9706), .Z(n7644) );
  XOR U11485 ( .A(round_reg[412]), .B(n10509), .Z(n8803) );
  XOR U11486 ( .A(n3171), .B(n11297), .Z(n11292) );
  XNOR U11487 ( .A(n6106), .B(n7634), .Z(n11297) );
  XOR U11488 ( .A(n11298), .B(n7650), .Z(n7634) );
  XNOR U11489 ( .A(round_reg[1229]), .B(n10802), .Z(n7650) );
  ANDN U11490 ( .B(n8805), .A(n7649), .Z(n11298) );
  XNOR U11491 ( .A(round_reg[871]), .B(n9984), .Z(n7649) );
  XOR U11492 ( .A(round_reg[482]), .B(n11299), .Z(n8805) );
  XNOR U11493 ( .A(n11300), .B(n7654), .Z(n6106) );
  XNOR U11494 ( .A(round_reg[1082]), .B(n11146), .Z(n7654) );
  ANDN U11495 ( .B(n11232), .A(n7653), .Z(n11300) );
  XOR U11496 ( .A(n11301), .B(n8726), .Z(n3171) );
  IV U11497 ( .A(n7657), .Z(n8726) );
  XOR U11498 ( .A(round_reg[1131]), .B(n9983), .Z(n7657) );
  AND U11499 ( .A(n8800), .B(n7658), .Z(n11301) );
  XOR U11500 ( .A(round_reg[728]), .B(n11302), .Z(n7658) );
  XNOR U11501 ( .A(round_reg[361]), .B(n10207), .Z(n8800) );
  XOR U11502 ( .A(n11303), .B(n11304), .Z(n6127) );
  XNOR U11503 ( .A(n5280), .B(n1924), .Z(n11304) );
  XNOR U11504 ( .A(n11305), .B(n8860), .Z(n1924) );
  ANDN U11505 ( .B(n7729), .A(n8787), .Z(n11305) );
  XNOR U11506 ( .A(round_reg[286]), .B(n9473), .Z(n8787) );
  XNOR U11507 ( .A(round_reg[1519]), .B(n10532), .Z(n7729) );
  IV U11508 ( .A(n11306), .Z(n10532) );
  XNOR U11509 ( .A(n11307), .B(n8865), .Z(n5280) );
  NOR U11510 ( .A(n7721), .B(n8784), .Z(n11307) );
  XNOR U11511 ( .A(round_reg[120]), .B(n11308), .Z(n8784) );
  XOR U11512 ( .A(round_reg[1301]), .B(n9987), .Z(n7721) );
  XOR U11513 ( .A(n11309), .B(n11310), .Z(n9987) );
  XNOR U11514 ( .A(n3679), .B(n11311), .Z(n11303) );
  XOR U11515 ( .A(n8841), .B(n4124), .Z(n11311) );
  XNOR U11516 ( .A(n11312), .B(n8867), .Z(n4124) );
  ANDN U11517 ( .B(n7712), .A(n8794), .Z(n11312) );
  XOR U11518 ( .A(round_reg[179]), .B(n10524), .Z(n8794) );
  XOR U11519 ( .A(round_reg[1364]), .B(n11313), .Z(n7712) );
  XNOR U11520 ( .A(n11314), .B(n8863), .Z(n8841) );
  ANDN U11521 ( .B(n7716), .A(n8790), .Z(n11314) );
  XNOR U11522 ( .A(round_reg[34]), .B(n10799), .Z(n8790) );
  XNOR U11523 ( .A(round_reg[1584]), .B(n9769), .Z(n7716) );
  XNOR U11524 ( .A(n11315), .B(n11316), .Z(n3679) );
  ANDN U11525 ( .B(n8792), .A(n7725), .Z(n11315) );
  XNOR U11526 ( .A(round_reg[1458]), .B(n10617), .Z(n7725) );
  XOR U11527 ( .A(n11317), .B(n7653), .Z(n8798) );
  XNOR U11528 ( .A(round_reg[650]), .B(n10983), .Z(n7653) );
  IV U11529 ( .A(n10947), .Z(n10983) );
  NOR U11530 ( .A(n8731), .B(n11232), .Z(n11317) );
  XOR U11531 ( .A(round_reg[584]), .B(n9116), .Z(n11232) );
  XNOR U11532 ( .A(round_reg[239]), .B(n11306), .Z(n8731) );
  XOR U11533 ( .A(n10278), .B(n11318), .Z(n11306) );
  XOR U11534 ( .A(n11319), .B(n11320), .Z(n10278) );
  XNOR U11535 ( .A(round_reg[1454]), .B(round_reg[1134]), .Z(n11320) );
  XOR U11536 ( .A(round_reg[174]), .B(n11321), .Z(n11319) );
  XOR U11537 ( .A(round_reg[814]), .B(round_reg[494]), .Z(n11321) );
  ANDN U11538 ( .B(n5694), .A(n5696), .Z(n11291) );
  XOR U11539 ( .A(n10471), .B(n2090), .Z(n5696) );
  XNOR U11540 ( .A(n8115), .B(n9222), .Z(n2090) );
  XNOR U11541 ( .A(n11322), .B(n11323), .Z(n9222) );
  XOR U11542 ( .A(n5494), .B(n3585), .Z(n11323) );
  XOR U11543 ( .A(n11324), .B(n11325), .Z(n3585) );
  ANDN U11544 ( .B(n8249), .A(n8247), .Z(n11324) );
  XOR U11545 ( .A(round_reg[918]), .B(n10021), .Z(n8249) );
  XOR U11546 ( .A(n11326), .B(n11327), .Z(n5494) );
  ANDN U11547 ( .B(n8243), .A(n8245), .Z(n11326) );
  XNOR U11548 ( .A(round_reg[814]), .B(n11328), .Z(n8245) );
  XOR U11549 ( .A(round_reg[1197]), .B(n11329), .Z(n8243) );
  XNOR U11550 ( .A(n6336), .B(n11330), .Z(n11322) );
  XOR U11551 ( .A(n2369), .B(n5468), .Z(n11330) );
  XNOR U11552 ( .A(n11331), .B(n10567), .Z(n5468) );
  ANDN U11553 ( .B(n9226), .A(n9224), .Z(n11331) );
  XNOR U11554 ( .A(round_reg[1269]), .B(n9387), .Z(n9224) );
  IV U11555 ( .A(n10627), .Z(n9387) );
  XNOR U11556 ( .A(n11332), .B(n11227), .Z(n10627) );
  XNOR U11557 ( .A(n11333), .B(n11334), .Z(n11227) );
  XNOR U11558 ( .A(round_reg[1524]), .B(round_reg[1204]), .Z(n11334) );
  XOR U11559 ( .A(round_reg[244]), .B(n11335), .Z(n11333) );
  XOR U11560 ( .A(round_reg[884]), .B(round_reg[564]), .Z(n11335) );
  XOR U11561 ( .A(round_reg[847]), .B(n10291), .Z(n9226) );
  XNOR U11562 ( .A(n11336), .B(n10559), .Z(n2369) );
  ANDN U11563 ( .B(n8235), .A(n8233), .Z(n11336) );
  XOR U11564 ( .A(round_reg[1058]), .B(n10369), .Z(n8233) );
  XOR U11565 ( .A(round_reg[690]), .B(n9861), .Z(n8235) );
  XNOR U11566 ( .A(n11337), .B(n10564), .Z(n6336) );
  NOR U11567 ( .A(n8237), .B(n8238), .Z(n11337) );
  XOR U11568 ( .A(round_reg[1107]), .B(n10579), .Z(n8237) );
  XOR U11569 ( .A(n11338), .B(n11339), .Z(n8115) );
  XNOR U11570 ( .A(n3776), .B(n5132), .Z(n11339) );
  XOR U11571 ( .A(n11340), .B(n9148), .Z(n5132) );
  XNOR U11572 ( .A(round_reg[459]), .B(n9208), .Z(n9148) );
  AND U11573 ( .A(n10478), .B(n10477), .Z(n11340) );
  XNOR U11574 ( .A(round_reg[98]), .B(n10369), .Z(n10477) );
  XNOR U11575 ( .A(round_reg[1343]), .B(n11341), .Z(n10478) );
  XNOR U11576 ( .A(n11342), .B(n8180), .Z(n3776) );
  XNOR U11577 ( .A(round_reg[625]), .B(n11343), .Z(n8180) );
  NOR U11578 ( .A(n10469), .B(n10470), .Z(n11342) );
  XOR U11579 ( .A(round_reg[1436]), .B(n9441), .Z(n10470) );
  XNOR U11580 ( .A(round_reg[216]), .B(n9679), .Z(n10469) );
  XOR U11581 ( .A(n4257), .B(n11344), .Z(n11338) );
  XOR U11582 ( .A(n1723), .B(n10542), .Z(n11344) );
  XOR U11583 ( .A(n11345), .B(n8190), .Z(n10542) );
  XNOR U11584 ( .A(round_reg[389]), .B(n10293), .Z(n8190) );
  AND U11585 ( .A(n10467), .B(n10466), .Z(n11345) );
  XNOR U11586 ( .A(round_reg[12]), .B(n10771), .Z(n10466) );
  XNOR U11587 ( .A(round_reg[1562]), .B(n11346), .Z(n10467) );
  XOR U11588 ( .A(n11347), .B(n8184), .Z(n1723) );
  XNOR U11589 ( .A(round_reg[338]), .B(n10767), .Z(n8184) );
  AND U11590 ( .A(n10475), .B(n10474), .Z(n11347) );
  XNOR U11591 ( .A(round_reg[264]), .B(n9116), .Z(n10474) );
  XNOR U11592 ( .A(round_reg[1497]), .B(n9605), .Z(n10475) );
  IV U11593 ( .A(n9524), .Z(n9605) );
  XOR U11594 ( .A(n11348), .B(n11349), .Z(n9524) );
  XNOR U11595 ( .A(n11350), .B(n8195), .Z(n4257) );
  XNOR U11596 ( .A(round_reg[557]), .B(n10708), .Z(n8195) );
  ANDN U11597 ( .B(n10549), .A(n11265), .Z(n11350) );
  XOR U11598 ( .A(n11351), .B(n10549), .Z(n10471) );
  XNOR U11599 ( .A(round_reg[157]), .B(n9367), .Z(n10549) );
  ANDN U11600 ( .B(n11265), .A(n8193), .Z(n11351) );
  XOR U11601 ( .A(round_reg[966]), .B(n10674), .Z(n8193) );
  XOR U11602 ( .A(round_reg[1406]), .B(n10698), .Z(n11265) );
  IV U11603 ( .A(n11261), .Z(n10698) );
  XOR U11604 ( .A(n5156), .B(n8592), .Z(n5694) );
  XOR U11605 ( .A(n11352), .B(n8693), .Z(n8592) );
  ANDN U11606 ( .B(n11252), .A(n6472), .Z(n11352) );
  XOR U11607 ( .A(round_reg[1554]), .B(n10795), .Z(n6472) );
  IV U11608 ( .A(n10388), .Z(n10795) );
  XOR U11609 ( .A(n9712), .B(n6373), .Z(n5156) );
  XOR U11610 ( .A(n11353), .B(n11354), .Z(n6373) );
  XNOR U11611 ( .A(n5937), .B(n2124), .Z(n11354) );
  XOR U11612 ( .A(n11355), .B(n11356), .Z(n2124) );
  NOR U11613 ( .A(n6502), .B(n6503), .Z(n11355) );
  XOR U11614 ( .A(round_reg[1261]), .B(n9923), .Z(n6503) );
  XOR U11615 ( .A(round_reg[1334]), .B(n9630), .Z(n6502) );
  XOR U11616 ( .A(n11012), .B(n10714), .Z(n9630) );
  XOR U11617 ( .A(n11357), .B(n11358), .Z(n10714) );
  XNOR U11618 ( .A(round_reg[1589]), .B(round_reg[1269]), .Z(n11358) );
  XOR U11619 ( .A(round_reg[309]), .B(n11359), .Z(n11357) );
  XOR U11620 ( .A(round_reg[949]), .B(round_reg[629]), .Z(n11359) );
  XOR U11621 ( .A(n11360), .B(n11361), .Z(n11012) );
  XNOR U11622 ( .A(round_reg[118]), .B(round_reg[1078]), .Z(n11361) );
  XOR U11623 ( .A(round_reg[1398]), .B(n11362), .Z(n11360) );
  XOR U11624 ( .A(round_reg[758]), .B(round_reg[438]), .Z(n11362) );
  XOR U11625 ( .A(n11363), .B(n8711), .Z(n5937) );
  NOR U11626 ( .A(n6506), .B(n6507), .Z(n11363) );
  XNOR U11627 ( .A(round_reg[1021]), .B(n9615), .Z(n6507) );
  XNOR U11628 ( .A(round_reg[1397]), .B(n9191), .Z(n6506) );
  XOR U11629 ( .A(n3665), .B(n11364), .Z(n11353) );
  XOR U11630 ( .A(n4247), .B(n5458), .Z(n11364) );
  XOR U11631 ( .A(n11365), .B(n8703), .Z(n5458) );
  NOR U11632 ( .A(n6489), .B(n6490), .Z(n11365) );
  XNOR U11633 ( .A(round_reg[1050]), .B(n10688), .Z(n6490) );
  XOR U11634 ( .A(round_reg[1427]), .B(n10579), .Z(n6489) );
  XOR U11635 ( .A(n11366), .B(n11367), .Z(n4247) );
  ANDN U11636 ( .B(n6493), .A(n6494), .Z(n11366) );
  XOR U11637 ( .A(round_reg[1099]), .B(n9208), .Z(n6494) );
  XNOR U11638 ( .A(round_reg[1488]), .B(n11368), .Z(n6493) );
  XOR U11639 ( .A(n11369), .B(n11370), .Z(n3665) );
  NOR U11640 ( .A(n6498), .B(n6499), .Z(n11369) );
  XNOR U11641 ( .A(round_reg[1189]), .B(n11371), .Z(n6499) );
  XOR U11642 ( .A(n11372), .B(n11373), .Z(n9712) );
  XOR U11643 ( .A(n4835), .B(n8686), .Z(n11373) );
  XOR U11644 ( .A(n11374), .B(n6465), .Z(n8686) );
  XOR U11645 ( .A(round_reg[683]), .B(n9992), .Z(n6465) );
  IV U11646 ( .A(n9455), .Z(n9992) );
  XOR U11647 ( .A(n11375), .B(n11376), .Z(n9455) );
  NOR U11648 ( .A(n8590), .B(n8591), .Z(n11374) );
  XOR U11649 ( .A(round_reg[208]), .B(n10299), .Z(n8591) );
  IV U11650 ( .A(n11368), .Z(n10299) );
  XOR U11651 ( .A(round_reg[617]), .B(n11377), .Z(n8590) );
  XNOR U11652 ( .A(n11378), .B(n6469), .Z(n4835) );
  XOR U11653 ( .A(round_reg[761]), .B(n11223), .Z(n6469) );
  ANDN U11654 ( .B(n8595), .A(n8596), .Z(n11378) );
  XOR U11655 ( .A(round_reg[256]), .B(n9749), .Z(n8596) );
  XNOR U11656 ( .A(round_reg[330]), .B(n10947), .Z(n8595) );
  XOR U11657 ( .A(n2512), .B(n11381), .Z(n11372) );
  XOR U11658 ( .A(n3474), .B(n4289), .Z(n11381) );
  XNOR U11659 ( .A(n11382), .B(n6474), .Z(n4289) );
  XOR U11660 ( .A(round_reg[807]), .B(n10797), .Z(n6474) );
  ANDN U11661 ( .B(n8693), .A(n11252), .Z(n11382) );
  XOR U11662 ( .A(round_reg[4]), .B(n10845), .Z(n11252) );
  XNOR U11663 ( .A(round_reg[445]), .B(n11383), .Z(n8693) );
  XNOR U11664 ( .A(n11384), .B(n6478), .Z(n3474) );
  XOR U11665 ( .A(round_reg[840]), .B(n11045), .Z(n6478) );
  IV U11666 ( .A(n9213), .Z(n11045) );
  XOR U11667 ( .A(n11385), .B(n11386), .Z(n9213) );
  NOR U11668 ( .A(n8587), .B(n8588), .Z(n11384) );
  XOR U11669 ( .A(round_reg[90]), .B(n11141), .Z(n8588) );
  IV U11670 ( .A(n10688), .Z(n11141) );
  XOR U11671 ( .A(round_reg[451]), .B(n11387), .Z(n8587) );
  XNOR U11672 ( .A(n11388), .B(n6482), .Z(n2512) );
  XOR U11673 ( .A(round_reg[911]), .B(n10630), .Z(n6482) );
  IV U11674 ( .A(n11025), .Z(n10630) );
  NOR U11675 ( .A(n8598), .B(n8599), .Z(n11388) );
  XOR U11676 ( .A(round_reg[149]), .B(n9910), .Z(n8599) );
  XOR U11677 ( .A(round_reg[549]), .B(n11371), .Z(n8598) );
  IV U11678 ( .A(n10171), .Z(n11371) );
  XOR U11679 ( .A(n11389), .B(n6254), .Z(out[1005]) );
  XOR U11680 ( .A(n8858), .B(n2291), .Z(n6254) );
  XNOR U11681 ( .A(n6133), .B(n6213), .Z(n2291) );
  XNOR U11682 ( .A(n11390), .B(n11391), .Z(n6213) );
  XOR U11683 ( .A(n2331), .B(n5479), .Z(n11391) );
  XOR U11684 ( .A(n11392), .B(n8795), .Z(n5479) );
  IV U11685 ( .A(n7714), .Z(n8795) );
  XOR U11686 ( .A(round_reg[988]), .B(n9778), .Z(n7714) );
  ANDN U11687 ( .B(n8867), .A(n7713), .Z(n11392) );
  XNOR U11688 ( .A(round_reg[941]), .B(n9923), .Z(n7713) );
  XOR U11689 ( .A(round_reg[515]), .B(n9623), .Z(n8867) );
  IV U11690 ( .A(n9636), .Z(n9623) );
  XNOR U11691 ( .A(n11393), .B(n7718), .Z(n2331) );
  XNOR U11692 ( .A(round_reg[1156]), .B(n9555), .Z(n7718) );
  ANDN U11693 ( .B(n8863), .A(n7717), .Z(n11393) );
  XOR U11694 ( .A(round_reg[773]), .B(n9700), .Z(n7717) );
  XOR U11695 ( .A(round_reg[411]), .B(n10601), .Z(n8863) );
  XOR U11696 ( .A(n3175), .B(n11396), .Z(n11390) );
  XNOR U11697 ( .A(n6163), .B(n7707), .Z(n11396) );
  XOR U11698 ( .A(n11397), .B(n8785), .Z(n7707) );
  IV U11699 ( .A(n7723), .Z(n8785) );
  XOR U11700 ( .A(round_reg[1228]), .B(n10941), .Z(n7723) );
  ANDN U11701 ( .B(n8865), .A(n7722), .Z(n11397) );
  XNOR U11702 ( .A(round_reg[870]), .B(n10045), .Z(n7722) );
  XOR U11703 ( .A(round_reg[481]), .B(n11400), .Z(n8865) );
  XNOR U11704 ( .A(n11401), .B(n7727), .Z(n6163) );
  XNOR U11705 ( .A(round_reg[1081]), .B(n11223), .Z(n7727) );
  ANDN U11706 ( .B(n11316), .A(n7726), .Z(n11401) );
  XOR U11707 ( .A(n11402), .B(n7731), .Z(n3175) );
  XNOR U11708 ( .A(round_reg[1130]), .B(n10044), .Z(n7731) );
  ANDN U11709 ( .B(n8860), .A(n7730), .Z(n11402) );
  XOR U11710 ( .A(round_reg[727]), .B(n11063), .Z(n7730) );
  XOR U11711 ( .A(round_reg[360]), .B(n9693), .Z(n8860) );
  XOR U11712 ( .A(n11403), .B(n11404), .Z(n6133) );
  XNOR U11713 ( .A(n5283), .B(n1928), .Z(n11404) );
  XNOR U11714 ( .A(n11405), .B(n8919), .Z(n1928) );
  ANDN U11715 ( .B(n7804), .A(n8847), .Z(n11405) );
  XNOR U11716 ( .A(round_reg[285]), .B(n9556), .Z(n8847) );
  XNOR U11717 ( .A(n11406), .B(n11407), .Z(n9556) );
  XNOR U11718 ( .A(round_reg[1518]), .B(n11267), .Z(n7804) );
  XNOR U11719 ( .A(n11408), .B(n8924), .Z(n5283) );
  AND U11720 ( .A(n7796), .B(n8845), .Z(n11408) );
  XNOR U11721 ( .A(round_reg[1300]), .B(n10048), .Z(n7796) );
  IV U11722 ( .A(n10574), .Z(n10048) );
  XNOR U11723 ( .A(n11410), .B(n11411), .Z(n10574) );
  XNOR U11724 ( .A(n3685), .B(n11412), .Z(n11403) );
  XOR U11725 ( .A(n8901), .B(n4127), .Z(n11412) );
  XNOR U11726 ( .A(n11413), .B(n8926), .Z(n4127) );
  ANDN U11727 ( .B(n8855), .A(n8854), .Z(n11413) );
  XNOR U11728 ( .A(round_reg[178]), .B(n11414), .Z(n8854) );
  XNOR U11729 ( .A(round_reg[1363]), .B(n9183), .Z(n8855) );
  XNOR U11730 ( .A(n11415), .B(n8922), .Z(n8901) );
  ANDN U11731 ( .B(n7791), .A(n8850), .Z(n11415) );
  XNOR U11732 ( .A(round_reg[33]), .B(n9395), .Z(n8850) );
  IV U11733 ( .A(n10222), .Z(n9395) );
  XNOR U11734 ( .A(n11416), .B(n11417), .Z(n10222) );
  XOR U11735 ( .A(round_reg[1583]), .B(n11210), .Z(n7791) );
  XNOR U11736 ( .A(n11418), .B(n11419), .Z(n3685) );
  NOR U11737 ( .A(n7800), .B(n8852), .Z(n11418) );
  XNOR U11738 ( .A(round_reg[1457]), .B(n9913), .Z(n7800) );
  XOR U11739 ( .A(n11420), .B(n7726), .Z(n8858) );
  XNOR U11740 ( .A(round_reg[649]), .B(n11421), .Z(n7726) );
  NOR U11741 ( .A(n8792), .B(n11316), .Z(n11420) );
  XOR U11742 ( .A(round_reg[583]), .B(n9390), .Z(n11316) );
  XNOR U11743 ( .A(round_reg[238]), .B(n10623), .Z(n8792) );
  IV U11744 ( .A(n11267), .Z(n10623) );
  XOR U11745 ( .A(n11422), .B(n11423), .Z(n11267) );
  NOR U11746 ( .A(n5700), .B(n5698), .Z(n11389) );
  XNOR U11747 ( .A(n8705), .B(n5159), .Z(n5698) );
  XNOR U11748 ( .A(n11424), .B(n11425), .Z(n6459) );
  XNOR U11749 ( .A(n4327), .B(n2520), .Z(n11425) );
  XNOR U11750 ( .A(n11426), .B(n6508), .Z(n2520) );
  XOR U11751 ( .A(round_reg[910]), .B(n10713), .Z(n6508) );
  AND U11752 ( .A(n8710), .B(n8711), .Z(n11426) );
  XNOR U11753 ( .A(round_reg[148]), .B(n9997), .Z(n8711) );
  XNOR U11754 ( .A(n11427), .B(n11428), .Z(n9997) );
  XOR U11755 ( .A(round_reg[548]), .B(n10282), .Z(n8710) );
  XNOR U11756 ( .A(n11429), .B(n6500), .Z(n4327) );
  XOR U11757 ( .A(round_reg[806]), .B(n10441), .Z(n6500) );
  AND U11758 ( .A(n8754), .B(n11370), .Z(n11429) );
  XOR U11759 ( .A(n3477), .B(n11430), .Z(n11424) );
  XNOR U11760 ( .A(n8747), .B(n4839), .Z(n11430) );
  XNOR U11761 ( .A(n11431), .B(n6495), .Z(n4839) );
  XOR U11762 ( .A(round_reg[760]), .B(n11308), .Z(n6495) );
  AND U11763 ( .A(n8707), .B(n11367), .Z(n11431) );
  IV U11764 ( .A(n8708), .Z(n11367) );
  XOR U11765 ( .A(round_reg[319]), .B(n9930), .Z(n8708) );
  XOR U11766 ( .A(round_reg[329]), .B(n11421), .Z(n8707) );
  IV U11767 ( .A(n10438), .Z(n11421) );
  XOR U11768 ( .A(n11432), .B(n6491), .Z(n8747) );
  XOR U11769 ( .A(round_reg[682]), .B(n10515), .Z(n6491) );
  AND U11770 ( .A(n8702), .B(n8703), .Z(n11432) );
  XOR U11771 ( .A(round_reg[207]), .B(n10291), .Z(n8703) );
  XOR U11772 ( .A(round_reg[616]), .B(n10036), .Z(n8702) );
  XNOR U11773 ( .A(n11433), .B(n6504), .Z(n3477) );
  XOR U11774 ( .A(round_reg[839]), .B(n11133), .Z(n6504) );
  AND U11775 ( .A(n8699), .B(n11356), .Z(n11433) );
  IV U11776 ( .A(n8700), .Z(n11356) );
  XNOR U11777 ( .A(round_reg[89]), .B(n10776), .Z(n8700) );
  XOR U11778 ( .A(round_reg[450]), .B(n9859), .Z(n8699) );
  XNOR U11779 ( .A(n11434), .B(n11435), .Z(n6378) );
  XOR U11780 ( .A(n5462), .B(n3669), .Z(n11435) );
  XOR U11781 ( .A(n11436), .B(n11437), .Z(n3669) );
  ANDN U11782 ( .B(n6524), .A(n6525), .Z(n11436) );
  XOR U11783 ( .A(round_reg[1188]), .B(n10282), .Z(n6525) );
  XNOR U11784 ( .A(n11438), .B(n8764), .Z(n5462) );
  ANDN U11785 ( .B(n6515), .A(n6516), .Z(n11438) );
  XNOR U11786 ( .A(round_reg[1049]), .B(n10776), .Z(n6516) );
  XOR U11787 ( .A(round_reg[1426]), .B(n11027), .Z(n6515) );
  XNOR U11788 ( .A(n4249), .B(n11439), .Z(n11434) );
  XOR U11789 ( .A(n5942), .B(n2128), .Z(n11439) );
  XOR U11790 ( .A(n11440), .B(n8761), .Z(n2128) );
  ANDN U11791 ( .B(n6528), .A(n6529), .Z(n11440) );
  XNOR U11792 ( .A(round_reg[1260]), .B(n10010), .Z(n6529) );
  XOR U11793 ( .A(round_reg[1333]), .B(n9257), .Z(n6528) );
  XOR U11794 ( .A(n11441), .B(n8772), .Z(n5942) );
  ANDN U11795 ( .B(n6532), .A(n6533), .Z(n11441) );
  XOR U11796 ( .A(round_reg[1020]), .B(n11442), .Z(n6533) );
  XOR U11797 ( .A(round_reg[1396]), .B(n11443), .Z(n6532) );
  XOR U11798 ( .A(n11444), .B(n8769), .Z(n4249) );
  ANDN U11799 ( .B(n6519), .A(n6520), .Z(n11444) );
  XNOR U11800 ( .A(round_reg[1098]), .B(n9393), .Z(n6520) );
  XOR U11801 ( .A(round_reg[1487]), .B(n10968), .Z(n6519) );
  IV U11802 ( .A(n10291), .Z(n10968) );
  XNOR U11803 ( .A(n11447), .B(n8754), .Z(n8705) );
  XOR U11804 ( .A(round_reg[444]), .B(n11138), .Z(n8754) );
  XOR U11805 ( .A(round_reg[3]), .B(n9826), .Z(n11370) );
  XOR U11806 ( .A(round_reg[1553]), .B(n10500), .Z(n6498) );
  XOR U11807 ( .A(n10560), .B(n2094), .Z(n5700) );
  XNOR U11808 ( .A(n8175), .B(n9329), .Z(n2094) );
  XNOR U11809 ( .A(n11448), .B(n11449), .Z(n9329) );
  XOR U11810 ( .A(n5498), .B(n3590), .Z(n11449) );
  XOR U11811 ( .A(n11450), .B(n11451), .Z(n3590) );
  ANDN U11812 ( .B(n8299), .A(n8300), .Z(n11450) );
  XNOR U11813 ( .A(round_reg[917]), .B(n10164), .Z(n8300) );
  XNOR U11814 ( .A(n11452), .B(n10645), .Z(n5498) );
  ANDN U11815 ( .B(n8295), .A(n8297), .Z(n11452) );
  XNOR U11816 ( .A(round_reg[813]), .B(n10303), .Z(n8297) );
  IV U11817 ( .A(n11140), .Z(n10303) );
  XOR U11818 ( .A(round_reg[1196]), .B(n10796), .Z(n8295) );
  XOR U11819 ( .A(n6340), .B(n11453), .Z(n11448) );
  XOR U11820 ( .A(n2376), .B(n5525), .Z(n11453) );
  XNOR U11821 ( .A(n11454), .B(n10656), .Z(n5525) );
  AND U11822 ( .A(n9332), .B(n9331), .Z(n11454) );
  XOR U11823 ( .A(round_reg[1268]), .B(n9459), .Z(n9331) );
  XOR U11824 ( .A(n11455), .B(n11456), .Z(n9459) );
  XNOR U11825 ( .A(round_reg[846]), .B(n10957), .Z(n9332) );
  XNOR U11826 ( .A(n11457), .B(n10648), .Z(n2376) );
  ANDN U11827 ( .B(n8287), .A(n8285), .Z(n11457) );
  XOR U11828 ( .A(round_reg[1057]), .B(n10140), .Z(n8285) );
  XOR U11829 ( .A(round_reg[689]), .B(n11458), .Z(n8287) );
  XOR U11830 ( .A(n11459), .B(n10653), .Z(n6340) );
  NOR U11831 ( .A(n8289), .B(n8290), .Z(n11459) );
  XNOR U11832 ( .A(round_reg[767]), .B(n11460), .Z(n8290) );
  XNOR U11833 ( .A(round_reg[1106]), .B(n11027), .Z(n8289) );
  XOR U11834 ( .A(n11461), .B(n11462), .Z(n8175) );
  XNOR U11835 ( .A(n3780), .B(n5135), .Z(n11462) );
  XOR U11836 ( .A(n11463), .B(n9225), .Z(n5135) );
  XOR U11837 ( .A(round_reg[458]), .B(n9393), .Z(n9225) );
  AND U11838 ( .A(n10567), .B(n10566), .Z(n11463) );
  XNOR U11839 ( .A(round_reg[97]), .B(n10140), .Z(n10566) );
  XNOR U11840 ( .A(n11464), .B(n11465), .Z(n10140) );
  XOR U11841 ( .A(round_reg[1342]), .B(n9536), .Z(n10567) );
  XNOR U11842 ( .A(n11466), .B(n8234), .Z(n3780) );
  XNOR U11843 ( .A(round_reg[624]), .B(n11467), .Z(n8234) );
  ANDN U11844 ( .B(n10559), .A(n10558), .Z(n11466) );
  XNOR U11845 ( .A(round_reg[215]), .B(n9752), .Z(n10558) );
  XNOR U11846 ( .A(round_reg[1435]), .B(n9527), .Z(n10559) );
  XOR U11847 ( .A(n4288), .B(n11468), .Z(n11461) );
  XOR U11848 ( .A(n1727), .B(n10631), .Z(n11468) );
  XOR U11849 ( .A(n11469), .B(n8244), .Z(n10631) );
  XNOR U11850 ( .A(round_reg[388]), .B(n10223), .Z(n8244) );
  IV U11851 ( .A(n10926), .Z(n10223) );
  XNOR U11852 ( .A(n11470), .B(n11471), .Z(n10926) );
  ANDN U11853 ( .B(n11327), .A(n10555), .Z(n11469) );
  XOR U11854 ( .A(round_reg[11]), .B(n10859), .Z(n10555) );
  XOR U11855 ( .A(n11472), .B(n11473), .Z(n10859) );
  IV U11856 ( .A(n10556), .Z(n11327) );
  XOR U11857 ( .A(round_reg[1561]), .B(n10216), .Z(n10556) );
  XNOR U11858 ( .A(n11474), .B(n8239), .Z(n1727) );
  XOR U11859 ( .A(round_reg[337]), .B(n10359), .Z(n8239) );
  AND U11860 ( .A(n10564), .B(n10563), .Z(n11474) );
  XNOR U11861 ( .A(round_reg[263]), .B(n9390), .Z(n10563) );
  XNOR U11862 ( .A(round_reg[1496]), .B(n9679), .Z(n10564) );
  IV U11863 ( .A(n9602), .Z(n9679) );
  XNOR U11864 ( .A(n11475), .B(n11476), .Z(n9602) );
  XNOR U11865 ( .A(n11477), .B(n8248), .Z(n4288) );
  XOR U11866 ( .A(round_reg[556]), .B(n10796), .Z(n8248) );
  NOR U11867 ( .A(n10638), .B(n11325), .Z(n11477) );
  XNOR U11868 ( .A(n11478), .B(n10638), .Z(n10560) );
  XNOR U11869 ( .A(round_reg[156]), .B(n9441), .Z(n10638) );
  IV U11870 ( .A(n11479), .Z(n9441) );
  AND U11871 ( .A(n8247), .B(n11325), .Z(n11478) );
  XOR U11872 ( .A(round_reg[1405]), .B(n10785), .Z(n11325) );
  IV U11873 ( .A(n11383), .Z(n10785) );
  XNOR U11874 ( .A(round_reg[965]), .B(n10763), .Z(n8247) );
  XOR U11875 ( .A(n11480), .B(n6259), .Z(out[1004]) );
  XOR U11876 ( .A(n8917), .B(n2298), .Z(n6259) );
  XNOR U11877 ( .A(n6139), .B(n6223), .Z(n2298) );
  XNOR U11878 ( .A(n11481), .B(n11482), .Z(n6223) );
  XOR U11879 ( .A(n2336), .B(n5484), .Z(n11482) );
  XOR U11880 ( .A(n11483), .B(n7789), .Z(n5484) );
  XNOR U11881 ( .A(round_reg[987]), .B(n9975), .Z(n7789) );
  ANDN U11882 ( .B(n8926), .A(n7788), .Z(n11483) );
  XOR U11883 ( .A(round_reg[940]), .B(n10010), .Z(n7788) );
  XOR U11884 ( .A(round_reg[514]), .B(n9695), .Z(n8926) );
  XNOR U11885 ( .A(n11484), .B(n7793), .Z(n2336) );
  XNOR U11886 ( .A(round_reg[1155]), .B(n9636), .Z(n7793) );
  ANDN U11887 ( .B(n8922), .A(n7792), .Z(n11484) );
  XNOR U11888 ( .A(round_reg[772]), .B(n11242), .Z(n7792) );
  XOR U11889 ( .A(round_reg[410]), .B(n10688), .Z(n8922) );
  XNOR U11890 ( .A(n11486), .B(n11487), .Z(n11202) );
  XNOR U11891 ( .A(round_reg[1434]), .B(round_reg[1114]), .Z(n11487) );
  XOR U11892 ( .A(round_reg[154]), .B(n11488), .Z(n11486) );
  XOR U11893 ( .A(round_reg[794]), .B(round_reg[474]), .Z(n11488) );
  XOR U11894 ( .A(n3179), .B(n11489), .Z(n11481) );
  XOR U11895 ( .A(n6218), .B(n7782), .Z(n11489) );
  XOR U11896 ( .A(n11490), .B(n7798), .Z(n7782) );
  XNOR U11897 ( .A(round_reg[1227]), .B(n11125), .Z(n7798) );
  ANDN U11898 ( .B(n8924), .A(n7797), .Z(n11490) );
  XNOR U11899 ( .A(round_reg[869]), .B(n10171), .Z(n7797) );
  XOR U11900 ( .A(round_reg[480]), .B(n9109), .Z(n8924) );
  XOR U11901 ( .A(n11493), .B(n11494), .Z(n11055) );
  XNOR U11902 ( .A(round_reg[1504]), .B(round_reg[1184]), .Z(n11494) );
  XOR U11903 ( .A(round_reg[224]), .B(n11495), .Z(n11493) );
  XOR U11904 ( .A(round_reg[864]), .B(round_reg[544]), .Z(n11495) );
  XOR U11905 ( .A(n11497), .B(n7802), .Z(n6218) );
  XNOR U11906 ( .A(round_reg[1080]), .B(n11308), .Z(n7802) );
  ANDN U11907 ( .B(n11419), .A(n7801), .Z(n11497) );
  XOR U11908 ( .A(n11498), .B(n7805), .Z(n3179) );
  XNOR U11909 ( .A(round_reg[1129]), .B(n10170), .Z(n7805) );
  IV U11910 ( .A(n10284), .Z(n10170) );
  AND U11911 ( .A(n8919), .B(n7806), .Z(n11498) );
  XOR U11912 ( .A(round_reg[726]), .B(n11499), .Z(n7806) );
  XNOR U11913 ( .A(round_reg[359]), .B(n10783), .Z(n8919) );
  XOR U11914 ( .A(n11500), .B(n11501), .Z(n6139) );
  XNOR U11915 ( .A(n5286), .B(n1932), .Z(n11501) );
  XNOR U11916 ( .A(n11502), .B(n8979), .Z(n1932) );
  ANDN U11917 ( .B(n7866), .A(n8907), .Z(n11502) );
  XOR U11918 ( .A(round_reg[284]), .B(n9637), .Z(n8907) );
  XNOR U11919 ( .A(n11503), .B(n11504), .Z(n9637) );
  XNOR U11920 ( .A(round_reg[1517]), .B(n11329), .Z(n7866) );
  XNOR U11921 ( .A(n11505), .B(n8984), .Z(n5286) );
  ANDN U11922 ( .B(n7858), .A(n8905), .Z(n11505) );
  XNOR U11923 ( .A(round_reg[118]), .B(n9108), .Z(n8905) );
  XNOR U11924 ( .A(round_reg[1299]), .B(n10174), .Z(n7858) );
  IV U11925 ( .A(n11030), .Z(n10174) );
  XNOR U11926 ( .A(n11428), .B(n11506), .Z(n11030) );
  XOR U11927 ( .A(n11507), .B(n11508), .Z(n11428) );
  XNOR U11928 ( .A(round_reg[1363]), .B(round_reg[1043]), .Z(n11508) );
  XOR U11929 ( .A(round_reg[403]), .B(n11509), .Z(n11507) );
  XOR U11930 ( .A(round_reg[83]), .B(round_reg[723]), .Z(n11509) );
  XNOR U11931 ( .A(n3689), .B(n11510), .Z(n11500) );
  XOR U11932 ( .A(n8961), .B(n4132), .Z(n11510) );
  XNOR U11933 ( .A(n11511), .B(n8986), .Z(n4132) );
  ANDN U11934 ( .B(n7849), .A(n8914), .Z(n11511) );
  XOR U11935 ( .A(round_reg[177]), .B(n9913), .Z(n8914) );
  XNOR U11936 ( .A(n11512), .B(n11513), .Z(n9913) );
  XOR U11937 ( .A(round_reg[1362]), .B(n11514), .Z(n7849) );
  XNOR U11938 ( .A(n11515), .B(n8982), .Z(n8961) );
  ANDN U11939 ( .B(n7853), .A(n8910), .Z(n11515) );
  XNOR U11940 ( .A(round_reg[32]), .B(n9471), .Z(n8910) );
  IV U11941 ( .A(n10972), .Z(n9471) );
  XOR U11942 ( .A(n11516), .B(n11517), .Z(n10972) );
  XNOR U11943 ( .A(round_reg[1582]), .B(n11295), .Z(n7853) );
  XNOR U11944 ( .A(n11518), .B(n11519), .Z(n3689) );
  ANDN U11945 ( .B(n8912), .A(n7862), .Z(n11518) );
  XNOR U11946 ( .A(round_reg[1456]), .B(n10001), .Z(n7862) );
  IV U11947 ( .A(n10790), .Z(n10001) );
  XOR U11948 ( .A(n11520), .B(n7801), .Z(n8917) );
  XNOR U11949 ( .A(round_reg[648]), .B(n10492), .Z(n7801) );
  ANDN U11950 ( .B(n8852), .A(n11419), .Z(n11520) );
  XOR U11951 ( .A(round_reg[582]), .B(n11521), .Z(n11419) );
  XNOR U11952 ( .A(round_reg[237]), .B(n11329), .Z(n8852) );
  IV U11953 ( .A(n10708), .Z(n11329) );
  XNOR U11954 ( .A(n11522), .B(n11523), .Z(n10708) );
  NOR U11955 ( .A(n5704), .B(n5702), .Z(n11480) );
  XNOR U11956 ( .A(n8766), .B(n5162), .Z(n5702) );
  XNOR U11957 ( .A(n11524), .B(n11525), .Z(n6485) );
  XNOR U11958 ( .A(n4748), .B(n2527), .Z(n11525) );
  XNOR U11959 ( .A(n11526), .B(n6534), .Z(n2527) );
  XOR U11960 ( .A(round_reg[909]), .B(n10802), .Z(n6534) );
  ANDN U11961 ( .B(n8771), .A(n8772), .Z(n11526) );
  XNOR U11962 ( .A(round_reg[147]), .B(n10579), .Z(n8772) );
  XOR U11963 ( .A(round_reg[547]), .B(n10433), .Z(n8771) );
  XNOR U11964 ( .A(n11527), .B(n6526), .Z(n4748) );
  XOR U11965 ( .A(round_reg[805]), .B(n10495), .Z(n6526) );
  ANDN U11966 ( .B(n8813), .A(n11437), .Z(n11527) );
  XOR U11967 ( .A(n3480), .B(n11528), .Z(n11524) );
  XNOR U11968 ( .A(n8808), .B(n4842), .Z(n11528) );
  XNOR U11969 ( .A(n11529), .B(n6521), .Z(n4842) );
  XOR U11970 ( .A(round_reg[759]), .B(n11409), .Z(n6521) );
  ANDN U11971 ( .B(n8768), .A(n8769), .Z(n11529) );
  XNOR U11972 ( .A(round_reg[318]), .B(n11530), .Z(n8769) );
  XOR U11973 ( .A(round_reg[328]), .B(n10492), .Z(n8768) );
  XOR U11974 ( .A(n11531), .B(n6517), .Z(n8808) );
  XOR U11975 ( .A(round_reg[681]), .B(n10207), .Z(n6517) );
  IV U11976 ( .A(n9620), .Z(n10207) );
  XNOR U11977 ( .A(n11532), .B(n11533), .Z(n9620) );
  NOR U11978 ( .A(n8763), .B(n8764), .Z(n11531) );
  XNOR U11979 ( .A(round_reg[206]), .B(n10364), .Z(n8764) );
  XOR U11980 ( .A(round_reg[615]), .B(n9818), .Z(n8763) );
  XNOR U11981 ( .A(n11534), .B(n6530), .Z(n3480) );
  XOR U11982 ( .A(round_reg[838]), .B(n11212), .Z(n6530) );
  ANDN U11983 ( .B(n8760), .A(n8761), .Z(n11534) );
  XNOR U11984 ( .A(round_reg[88]), .B(n10881), .Z(n8761) );
  XOR U11985 ( .A(round_reg[449]), .B(n10015), .Z(n8760) );
  XNOR U11986 ( .A(n11535), .B(n11536), .Z(n6382) );
  XOR U11987 ( .A(n5472), .B(n3673), .Z(n11536) );
  XOR U11988 ( .A(n11537), .B(n11538), .Z(n3673) );
  ANDN U11989 ( .B(n6549), .A(n6559), .Z(n11537) );
  XNOR U11990 ( .A(round_reg[1187]), .B(n11539), .Z(n6559) );
  XNOR U11991 ( .A(n11540), .B(n8825), .Z(n5472) );
  ANDN U11992 ( .B(n6541), .A(n6542), .Z(n11540) );
  XNOR U11993 ( .A(round_reg[1048]), .B(n10881), .Z(n6542) );
  XOR U11994 ( .A(round_reg[1425]), .B(n10300), .Z(n6541) );
  XNOR U11995 ( .A(n4251), .B(n11541), .Z(n11535) );
  XOR U11996 ( .A(n5947), .B(n2132), .Z(n11541) );
  XOR U11997 ( .A(n11542), .B(n8822), .Z(n2132) );
  ANDN U11998 ( .B(n6562), .A(n6563), .Z(n11542) );
  XNOR U11999 ( .A(round_reg[1259]), .B(n11543), .Z(n6563) );
  XOR U12000 ( .A(round_reg[1332]), .B(n10297), .Z(n6562) );
  XOR U12001 ( .A(n11544), .B(n8833), .Z(n5947) );
  ANDN U12002 ( .B(n6566), .A(n6567), .Z(n11544) );
  XOR U12003 ( .A(round_reg[1019]), .B(n11545), .Z(n6567) );
  XOR U12004 ( .A(round_reg[1395]), .B(n9827), .Z(n6566) );
  XOR U12005 ( .A(n11546), .B(n8830), .Z(n4251) );
  ANDN U12006 ( .B(n6545), .A(n6546), .Z(n11546) );
  XNOR U12007 ( .A(round_reg[1097]), .B(n9383), .Z(n6546) );
  XOR U12008 ( .A(round_reg[1486]), .B(n10957), .Z(n6545) );
  IV U12009 ( .A(n10364), .Z(n10957) );
  XOR U12010 ( .A(n11547), .B(n10990), .Z(n10364) );
  XOR U12011 ( .A(n11548), .B(n11549), .Z(n10990) );
  XNOR U12012 ( .A(round_reg[141]), .B(round_reg[1101]), .Z(n11549) );
  XOR U12013 ( .A(round_reg[1421]), .B(n11550), .Z(n11548) );
  XOR U12014 ( .A(round_reg[781]), .B(round_reg[461]), .Z(n11550) );
  XNOR U12015 ( .A(n11551), .B(n8813), .Z(n8766) );
  XOR U12016 ( .A(round_reg[443]), .B(n11058), .Z(n8813) );
  ANDN U12017 ( .B(n11437), .A(n6524), .Z(n11551) );
  XOR U12018 ( .A(round_reg[1552]), .B(n10541), .Z(n6524) );
  XNOR U12019 ( .A(round_reg[2]), .B(n9187), .Z(n11437) );
  XOR U12020 ( .A(n10649), .B(n2098), .Z(n5704) );
  XNOR U12021 ( .A(n8229), .B(n9399), .Z(n2098) );
  XNOR U12022 ( .A(n11552), .B(n11553), .Z(n9399) );
  XOR U12023 ( .A(n5502), .B(n3600), .Z(n11553) );
  XOR U12024 ( .A(n11554), .B(n11555), .Z(n3600) );
  ANDN U12025 ( .B(n8353), .A(n8351), .Z(n11554) );
  XOR U12026 ( .A(round_reg[916]), .B(n10273), .Z(n8353) );
  XOR U12027 ( .A(n11556), .B(n10731), .Z(n5502) );
  ANDN U12028 ( .B(n8347), .A(n8349), .Z(n11556) );
  XNOR U12029 ( .A(round_reg[812]), .B(n9986), .Z(n8349) );
  XOR U12030 ( .A(round_reg[1195]), .B(n10868), .Z(n8347) );
  XOR U12031 ( .A(n6344), .B(n11557), .Z(n11552) );
  XOR U12032 ( .A(n2383), .B(n5570), .Z(n11557) );
  XNOR U12033 ( .A(n11558), .B(n10742), .Z(n5570) );
  AND U12034 ( .A(n9403), .B(n9401), .Z(n11558) );
  XOR U12035 ( .A(round_reg[1267]), .B(n9544), .Z(n9401) );
  IV U12036 ( .A(n11196), .Z(n9544) );
  XNOR U12037 ( .A(n11559), .B(n11560), .Z(n11196) );
  XNOR U12038 ( .A(round_reg[845]), .B(n10527), .Z(n9403) );
  XNOR U12039 ( .A(n11561), .B(n10734), .Z(n2383) );
  ANDN U12040 ( .B(n8339), .A(n8337), .Z(n11561) );
  XOR U12041 ( .A(round_reg[1056]), .B(n10226), .Z(n8337) );
  XOR U12042 ( .A(round_reg[688]), .B(n11562), .Z(n8339) );
  XOR U12043 ( .A(n11563), .B(n10739), .Z(n6344) );
  NOR U12044 ( .A(n8341), .B(n8342), .Z(n11563) );
  XNOR U12045 ( .A(round_reg[766]), .B(n11261), .Z(n8342) );
  XOR U12046 ( .A(n11564), .B(n11565), .Z(n11261) );
  XNOR U12047 ( .A(round_reg[1105]), .B(n10300), .Z(n8341) );
  IV U12048 ( .A(n10762), .Z(n10300) );
  XOR U12049 ( .A(n11566), .B(n11567), .Z(n8229) );
  XNOR U12050 ( .A(n3784), .B(n5140), .Z(n11567) );
  XNOR U12051 ( .A(n11568), .B(n9333), .Z(n5140) );
  XNOR U12052 ( .A(round_reg[457]), .B(n9383), .Z(n9333) );
  XOR U12053 ( .A(n11569), .B(n11570), .Z(n9383) );
  AND U12054 ( .A(n10656), .B(n10655), .Z(n11568) );
  XNOR U12055 ( .A(round_reg[96]), .B(n10226), .Z(n10655) );
  XOR U12056 ( .A(n11571), .B(n11220), .Z(n10226) );
  XOR U12057 ( .A(n11572), .B(n11573), .Z(n11220) );
  XNOR U12058 ( .A(round_reg[31]), .B(round_reg[1311]), .Z(n11573) );
  XOR U12059 ( .A(round_reg[351]), .B(n11574), .Z(n11572) );
  XOR U12060 ( .A(round_reg[991]), .B(round_reg[671]), .Z(n11574) );
  XNOR U12061 ( .A(round_reg[1341]), .B(n11575), .Z(n10656) );
  XOR U12062 ( .A(n11576), .B(n8286), .Z(n3784) );
  IV U12063 ( .A(n10725), .Z(n8286) );
  XNOR U12064 ( .A(round_reg[623]), .B(n11210), .Z(n10725) );
  ANDN U12065 ( .B(n10648), .A(n10647), .Z(n11576) );
  XNOR U12066 ( .A(round_reg[214]), .B(n10666), .Z(n10647) );
  XNOR U12067 ( .A(round_reg[1434]), .B(n9607), .Z(n10648) );
  XOR U12068 ( .A(n4328), .B(n11577), .Z(n11566) );
  XOR U12069 ( .A(n1731), .B(n10716), .Z(n11577) );
  XOR U12070 ( .A(n11578), .B(n8296), .Z(n10716) );
  XNOR U12071 ( .A(round_reg[387]), .B(n10860), .Z(n8296) );
  IV U12072 ( .A(n11115), .Z(n10860) );
  XNOR U12073 ( .A(n11579), .B(n11580), .Z(n11115) );
  ANDN U12074 ( .B(n10644), .A(n10645), .Z(n11578) );
  XOR U12075 ( .A(round_reg[1560]), .B(n10302), .Z(n10645) );
  XNOR U12076 ( .A(round_reg[10]), .B(n10947), .Z(n10644) );
  XOR U12077 ( .A(n11581), .B(n11582), .Z(n10947) );
  XNOR U12078 ( .A(n11583), .B(n8291), .Z(n1731) );
  XOR U12079 ( .A(round_reg[336]), .B(n10445), .Z(n8291) );
  ANDN U12080 ( .B(n10653), .A(n10652), .Z(n11583) );
  XNOR U12081 ( .A(round_reg[262]), .B(n9465), .Z(n10652) );
  XNOR U12082 ( .A(round_reg[1495]), .B(n9752), .Z(n10653) );
  IV U12083 ( .A(n9677), .Z(n9752) );
  XNOR U12084 ( .A(n11586), .B(n8301), .Z(n4328) );
  XOR U12085 ( .A(round_reg[555]), .B(n10868), .Z(n8301) );
  NOR U12086 ( .A(n10723), .B(n11451), .Z(n11586) );
  XNOR U12087 ( .A(n11587), .B(n10723), .Z(n10649) );
  XNOR U12088 ( .A(round_reg[155]), .B(n9527), .Z(n10723) );
  ANDN U12089 ( .B(n11451), .A(n8299), .Z(n11587) );
  XOR U12090 ( .A(round_reg[964]), .B(n10845), .Z(n8299) );
  XOR U12091 ( .A(round_reg[1404]), .B(n11138), .Z(n11451) );
  XOR U12092 ( .A(n11588), .B(n6264), .Z(out[1003]) );
  XOR U12093 ( .A(n8977), .B(n2305), .Z(n6264) );
  XNOR U12094 ( .A(n6145), .B(n6228), .Z(n2305) );
  XNOR U12095 ( .A(n11589), .B(n11590), .Z(n6228) );
  XOR U12096 ( .A(n2343), .B(n5489), .Z(n11590) );
  XOR U12097 ( .A(n11591), .B(n7851), .Z(n5489) );
  XNOR U12098 ( .A(round_reg[986]), .B(n9865), .Z(n7851) );
  XOR U12099 ( .A(n11349), .B(n11592), .Z(n9865) );
  XOR U12100 ( .A(n11593), .B(n11594), .Z(n11349) );
  XNOR U12101 ( .A(round_reg[1561]), .B(round_reg[1241]), .Z(n11594) );
  XOR U12102 ( .A(round_reg[281]), .B(n11595), .Z(n11593) );
  XOR U12103 ( .A(round_reg[921]), .B(round_reg[601]), .Z(n11595) );
  ANDN U12104 ( .B(n8986), .A(n7850), .Z(n11591) );
  XNOR U12105 ( .A(round_reg[939]), .B(n11596), .Z(n7850) );
  XOR U12106 ( .A(round_reg[513]), .B(n9113), .Z(n8986) );
  IV U12107 ( .A(n9779), .Z(n9113) );
  XNOR U12108 ( .A(n11597), .B(n7855), .Z(n2343) );
  XNOR U12109 ( .A(round_reg[1154]), .B(n9709), .Z(n7855) );
  ANDN U12110 ( .B(n8982), .A(n7854), .Z(n11597) );
  XNOR U12111 ( .A(round_reg[771]), .B(n9266), .Z(n7854) );
  XOR U12112 ( .A(round_reg[409]), .B(n10776), .Z(n8982) );
  XOR U12113 ( .A(n11598), .B(n11287), .Z(n10776) );
  XOR U12114 ( .A(n11599), .B(n11600), .Z(n11287) );
  XNOR U12115 ( .A(round_reg[1433]), .B(round_reg[1113]), .Z(n11600) );
  XOR U12116 ( .A(round_reg[153]), .B(n11601), .Z(n11599) );
  XOR U12117 ( .A(round_reg[793]), .B(round_reg[473]), .Z(n11601) );
  XOR U12118 ( .A(n3182), .B(n11602), .Z(n11589) );
  XNOR U12119 ( .A(n6275), .B(n7844), .Z(n11602) );
  XOR U12120 ( .A(n11603), .B(n7860), .Z(n7844) );
  XNOR U12121 ( .A(round_reg[1226]), .B(n9087), .Z(n7860) );
  ANDN U12122 ( .B(n8984), .A(n7859), .Z(n11603) );
  XNOR U12123 ( .A(round_reg[868]), .B(n10282), .Z(n7859) );
  XOR U12124 ( .A(n11604), .B(n11276), .Z(n10282) );
  XNOR U12125 ( .A(n11605), .B(n11606), .Z(n11276) );
  XNOR U12126 ( .A(round_reg[1443]), .B(round_reg[1123]), .Z(n11606) );
  XOR U12127 ( .A(round_reg[163]), .B(n11607), .Z(n11605) );
  XOR U12128 ( .A(round_reg[803]), .B(round_reg[483]), .Z(n11607) );
  XOR U12129 ( .A(round_reg[479]), .B(n11205), .Z(n8984) );
  XNOR U12130 ( .A(n11608), .B(n11609), .Z(n11205) );
  XNOR U12131 ( .A(n11610), .B(n7864), .Z(n6275) );
  XNOR U12132 ( .A(round_reg[1079]), .B(n11409), .Z(n7864) );
  ANDN U12133 ( .B(n11519), .A(n7863), .Z(n11610) );
  XOR U12134 ( .A(n11611), .B(n7868), .Z(n3182) );
  XNOR U12135 ( .A(round_reg[1128]), .B(n10281), .Z(n7868) );
  IV U12136 ( .A(n10981), .Z(n10281) );
  ANDN U12137 ( .B(n8979), .A(n7867), .Z(n11611) );
  XNOR U12138 ( .A(round_reg[725]), .B(n11228), .Z(n7867) );
  XOR U12139 ( .A(round_reg[358]), .B(n10883), .Z(n8979) );
  XOR U12140 ( .A(n11612), .B(n11613), .Z(n6145) );
  XNOR U12141 ( .A(n5289), .B(n1937), .Z(n11613) );
  XNOR U12142 ( .A(n11614), .B(n9039), .Z(n1937) );
  ANDN U12143 ( .B(n7933), .A(n8967), .Z(n11614) );
  XNOR U12144 ( .A(round_reg[283]), .B(n10000), .Z(n8967) );
  IV U12145 ( .A(n9710), .Z(n10000) );
  XNOR U12146 ( .A(n11615), .B(n11616), .Z(n9710) );
  XNOR U12147 ( .A(round_reg[1516]), .B(n10796), .Z(n7933) );
  XNOR U12148 ( .A(n11617), .B(n9044), .Z(n5289) );
  ANDN U12149 ( .B(n7925), .A(n8965), .Z(n11617) );
  XNOR U12150 ( .A(round_reg[117]), .B(n9191), .Z(n8965) );
  XNOR U12151 ( .A(round_reg[1298]), .B(n10767), .Z(n7925) );
  IV U12152 ( .A(n10538), .Z(n10767) );
  XNOR U12153 ( .A(n11618), .B(n11259), .Z(n10538) );
  XNOR U12154 ( .A(n11619), .B(n11620), .Z(n11259) );
  XNOR U12155 ( .A(round_reg[1553]), .B(round_reg[1233]), .Z(n11620) );
  XOR U12156 ( .A(round_reg[273]), .B(n11621), .Z(n11619) );
  XOR U12157 ( .A(round_reg[913]), .B(round_reg[593]), .Z(n11621) );
  XNOR U12158 ( .A(n3693), .B(n11622), .Z(n11612) );
  XOR U12159 ( .A(n9020), .B(n4135), .Z(n11622) );
  XNOR U12160 ( .A(n11623), .B(n9046), .Z(n4135) );
  NOR U12161 ( .A(n7916), .B(n8974), .Z(n11623) );
  XNOR U12162 ( .A(round_reg[176]), .B(n10790), .Z(n8974) );
  XOR U12163 ( .A(n11624), .B(n11625), .Z(n10790) );
  XOR U12164 ( .A(round_reg[1361]), .B(n9829), .Z(n7916) );
  XNOR U12165 ( .A(n11626), .B(n9042), .Z(n9020) );
  ANDN U12166 ( .B(n7920), .A(n8970), .Z(n11626) );
  XNOR U12167 ( .A(round_reg[31]), .B(n9554), .Z(n8970) );
  XOR U12168 ( .A(n10855), .B(n11496), .Z(n9554) );
  XNOR U12169 ( .A(n11627), .B(n11628), .Z(n11496) );
  XNOR U12170 ( .A(round_reg[1375]), .B(round_reg[1055]), .Z(n11628) );
  XOR U12171 ( .A(round_reg[415]), .B(n11629), .Z(n11627) );
  XOR U12172 ( .A(round_reg[95]), .B(round_reg[735]), .Z(n11629) );
  XOR U12173 ( .A(n11630), .B(n11631), .Z(n10855) );
  XNOR U12174 ( .A(round_reg[1566]), .B(round_reg[1246]), .Z(n11631) );
  XOR U12175 ( .A(round_reg[286]), .B(n11632), .Z(n11630) );
  XOR U12176 ( .A(round_reg[926]), .B(round_reg[606]), .Z(n11632) );
  XNOR U12177 ( .A(round_reg[1581]), .B(n9923), .Z(n7920) );
  XNOR U12178 ( .A(n11633), .B(n11634), .Z(n3693) );
  NOR U12179 ( .A(n7929), .B(n8972), .Z(n11633) );
  XNOR U12180 ( .A(round_reg[1455]), .B(n10129), .Z(n7929) );
  IV U12181 ( .A(n10871), .Z(n10129) );
  XOR U12182 ( .A(n11635), .B(n7863), .Z(n8977) );
  XNOR U12183 ( .A(round_reg[647]), .B(n11018), .Z(n7863) );
  NOR U12184 ( .A(n8912), .B(n11519), .Z(n11635) );
  XOR U12185 ( .A(round_reg[581]), .B(n11636), .Z(n11519) );
  XOR U12186 ( .A(n11037), .B(n11637), .Z(n10796) );
  XOR U12187 ( .A(n11638), .B(n11639), .Z(n11037) );
  XNOR U12188 ( .A(round_reg[1451]), .B(round_reg[1131]), .Z(n11639) );
  XOR U12189 ( .A(round_reg[171]), .B(n11640), .Z(n11638) );
  XOR U12190 ( .A(round_reg[811]), .B(round_reg[491]), .Z(n11640) );
  NOR U12191 ( .A(n5714), .B(n5712), .Z(n11588) );
  XNOR U12192 ( .A(n8827), .B(n5165), .Z(n5712) );
  XNOR U12193 ( .A(n11641), .B(n11642), .Z(n6511) );
  XNOR U12194 ( .A(n5109), .B(n2534), .Z(n11642) );
  XNOR U12195 ( .A(n11643), .B(n6568), .Z(n2534) );
  XOR U12196 ( .A(round_reg[908]), .B(n10941), .Z(n6568) );
  IV U12197 ( .A(n10887), .Z(n10941) );
  ANDN U12198 ( .B(n8832), .A(n8833), .Z(n11643) );
  XNOR U12199 ( .A(round_reg[146]), .B(n11644), .Z(n8833) );
  XOR U12200 ( .A(round_reg[546]), .B(n10442), .Z(n8832) );
  XNOR U12201 ( .A(n11645), .B(n6560), .Z(n5109) );
  XOR U12202 ( .A(round_reg[804]), .B(n9830), .Z(n6560) );
  XOR U12203 ( .A(n11646), .B(n11647), .Z(n9830) );
  ANDN U12204 ( .B(n8875), .A(n11538), .Z(n11645) );
  XOR U12205 ( .A(n3482), .B(n11648), .Z(n11641) );
  XNOR U12206 ( .A(n8868), .B(n4846), .Z(n11648) );
  XNOR U12207 ( .A(n11649), .B(n6547), .Z(n4846) );
  XOR U12208 ( .A(round_reg[758]), .B(n9108), .Z(n6547) );
  ANDN U12209 ( .B(n8829), .A(n8830), .Z(n11649) );
  XNOR U12210 ( .A(round_reg[317]), .B(n10592), .Z(n8830) );
  XOR U12211 ( .A(n11650), .B(n11564), .Z(n10592) );
  XOR U12212 ( .A(n11651), .B(n11652), .Z(n11564) );
  XNOR U12213 ( .A(round_reg[1341]), .B(round_reg[1021]), .Z(n11652) );
  XOR U12214 ( .A(round_reg[381]), .B(n11653), .Z(n11651) );
  XOR U12215 ( .A(round_reg[701]), .B(round_reg[61]), .Z(n11653) );
  XOR U12216 ( .A(round_reg[327]), .B(n11018), .Z(n8829) );
  XOR U12217 ( .A(n11654), .B(n6543), .Z(n8868) );
  XOR U12218 ( .A(round_reg[680]), .B(n10289), .Z(n6543) );
  IV U12219 ( .A(n9693), .Z(n10289) );
  XNOR U12220 ( .A(n11655), .B(n11656), .Z(n9693) );
  ANDN U12221 ( .B(n8824), .A(n8825), .Z(n11654) );
  XOR U12222 ( .A(round_reg[205]), .B(n10527), .Z(n8825) );
  XOR U12223 ( .A(round_reg[614]), .B(n9889), .Z(n8824) );
  XNOR U12224 ( .A(n11658), .B(n11659), .Z(n10847) );
  XNOR U12225 ( .A(round_reg[358]), .B(round_reg[1318]), .Z(n11659) );
  XOR U12226 ( .A(round_reg[38]), .B(n11660), .Z(n11658) );
  XOR U12227 ( .A(round_reg[998]), .B(round_reg[678]), .Z(n11660) );
  XNOR U12228 ( .A(n11661), .B(n6564), .Z(n3482) );
  XOR U12229 ( .A(round_reg[837]), .B(n9472), .Z(n6564) );
  IV U12230 ( .A(n9458), .Z(n9472) );
  XNOR U12231 ( .A(n11662), .B(n11471), .Z(n9458) );
  XNOR U12232 ( .A(n11663), .B(n11664), .Z(n11471) );
  XNOR U12233 ( .A(round_reg[132]), .B(round_reg[1092]), .Z(n11664) );
  XOR U12234 ( .A(round_reg[1412]), .B(n11665), .Z(n11663) );
  XOR U12235 ( .A(round_reg[772]), .B(round_reg[452]), .Z(n11665) );
  ANDN U12236 ( .B(n8821), .A(n8822), .Z(n11661) );
  XNOR U12237 ( .A(round_reg[87]), .B(n11063), .Z(n8822) );
  XOR U12238 ( .A(round_reg[448]), .B(n9534), .Z(n8821) );
  XNOR U12239 ( .A(n11666), .B(n11667), .Z(n6386) );
  XOR U12240 ( .A(n5478), .B(n3677), .Z(n11667) );
  XOR U12241 ( .A(n11668), .B(n11669), .Z(n3677) );
  ANDN U12242 ( .B(n6584), .A(n6586), .Z(n11668) );
  XNOR U12243 ( .A(round_reg[1186]), .B(n11670), .Z(n6586) );
  XNOR U12244 ( .A(n11671), .B(n8885), .Z(n5478) );
  ANDN U12245 ( .B(n6575), .A(n6576), .Z(n11671) );
  XNOR U12246 ( .A(round_reg[1047]), .B(n11063), .Z(n6576) );
  XOR U12247 ( .A(round_reg[1424]), .B(n10372), .Z(n6575) );
  XNOR U12248 ( .A(n4253), .B(n11672), .Z(n11666) );
  XOR U12249 ( .A(n5952), .B(n2136), .Z(n11672) );
  XOR U12250 ( .A(n11673), .B(n8882), .Z(n2136) );
  ANDN U12251 ( .B(n6588), .A(n6589), .Z(n11673) );
  XNOR U12252 ( .A(round_reg[1258]), .B(n10220), .Z(n6589) );
  XOR U12253 ( .A(round_reg[1331]), .B(n10370), .Z(n6588) );
  IV U12254 ( .A(n9437), .Z(n10370) );
  XOR U12255 ( .A(n11674), .B(n8893), .Z(n5952) );
  NOR U12256 ( .A(n6592), .B(n6593), .Z(n11674) );
  XNOR U12257 ( .A(round_reg[1018]), .B(n11675), .Z(n6593) );
  XNOR U12258 ( .A(round_reg[1394]), .B(n9896), .Z(n6592) );
  XOR U12259 ( .A(n11676), .B(n8890), .Z(n4253) );
  ANDN U12260 ( .B(n6579), .A(n6580), .Z(n11676) );
  XNOR U12261 ( .A(round_reg[1096]), .B(n9463), .Z(n6580) );
  XOR U12262 ( .A(round_reg[1485]), .B(n10527), .Z(n6579) );
  XOR U12263 ( .A(n11677), .B(n11032), .Z(n10527) );
  XNOR U12264 ( .A(n11678), .B(n11679), .Z(n11032) );
  XNOR U12265 ( .A(round_reg[140]), .B(round_reg[1100]), .Z(n11679) );
  XOR U12266 ( .A(round_reg[1420]), .B(n11680), .Z(n11678) );
  XOR U12267 ( .A(round_reg[780]), .B(round_reg[460]), .Z(n11680) );
  XNOR U12268 ( .A(n11681), .B(n8875), .Z(n8827) );
  XOR U12269 ( .A(round_reg[442]), .B(n11146), .Z(n8875) );
  ANDN U12270 ( .B(n11538), .A(n6549), .Z(n11681) );
  XNOR U12271 ( .A(round_reg[1551]), .B(n11025), .Z(n6549) );
  XOR U12272 ( .A(n11682), .B(n11683), .Z(n11025) );
  XNOR U12273 ( .A(round_reg[1]), .B(n9966), .Z(n11538) );
  XOR U12274 ( .A(n10735), .B(n2101), .Z(n5714) );
  XNOR U12275 ( .A(n8281), .B(n9476), .Z(n2101) );
  XNOR U12276 ( .A(n11684), .B(n11685), .Z(n9476) );
  XNOR U12277 ( .A(n5507), .B(n3603), .Z(n11685) );
  XOR U12278 ( .A(n11686), .B(n11687), .Z(n3603) );
  ANDN U12279 ( .B(n8405), .A(n8403), .Z(n11686) );
  XOR U12280 ( .A(round_reg[915]), .B(n10317), .Z(n8405) );
  XNOR U12281 ( .A(n11688), .B(n10817), .Z(n5507) );
  AND U12282 ( .A(n8401), .B(n8399), .Z(n11688) );
  XOR U12283 ( .A(round_reg[1194]), .B(n11048), .Z(n8399) );
  XNOR U12284 ( .A(round_reg[811]), .B(n9983), .Z(n8401) );
  IV U12285 ( .A(n10047), .Z(n9983) );
  XNOR U12286 ( .A(n11689), .B(n11690), .Z(n10047) );
  XNOR U12287 ( .A(n6348), .B(n11691), .Z(n11684) );
  XOR U12288 ( .A(n2390), .B(n5616), .Z(n11691) );
  XNOR U12289 ( .A(n11692), .B(n10828), .Z(n5616) );
  AND U12290 ( .A(n9480), .B(n9478), .Z(n11692) );
  XOR U12291 ( .A(round_reg[1266]), .B(n9624), .Z(n9478) );
  IV U12292 ( .A(n11281), .Z(n9624) );
  XOR U12293 ( .A(n11693), .B(n11512), .Z(n11281) );
  XOR U12294 ( .A(n11694), .B(n11695), .Z(n11512) );
  XNOR U12295 ( .A(round_reg[1521]), .B(round_reg[1201]), .Z(n11695) );
  XOR U12296 ( .A(round_reg[241]), .B(n11696), .Z(n11694) );
  XOR U12297 ( .A(round_reg[881]), .B(round_reg[561]), .Z(n11696) );
  XNOR U12298 ( .A(round_reg[844]), .B(n10535), .Z(n9480) );
  XNOR U12299 ( .A(n11697), .B(n10820), .Z(n2390) );
  AND U12300 ( .A(n8389), .B(n8390), .Z(n11697) );
  IV U12301 ( .A(n10897), .Z(n8390) );
  XOR U12302 ( .A(round_reg[687]), .B(n9079), .Z(n10897) );
  IV U12303 ( .A(n11698), .Z(n9079) );
  XOR U12304 ( .A(round_reg[1055]), .B(n11699), .Z(n8389) );
  XNOR U12305 ( .A(n11700), .B(n10825), .Z(n6348) );
  NOR U12306 ( .A(n8393), .B(n8395), .Z(n11700) );
  XNOR U12307 ( .A(round_reg[765]), .B(n11383), .Z(n8395) );
  XOR U12308 ( .A(n11701), .B(n11702), .Z(n11383) );
  XNOR U12309 ( .A(round_reg[1104]), .B(n10372), .Z(n8393) );
  IV U12310 ( .A(n10844), .Z(n10372) );
  XOR U12311 ( .A(n11703), .B(n11704), .Z(n8281) );
  XNOR U12312 ( .A(n3788), .B(n5143), .Z(n11704) );
  XOR U12313 ( .A(n11705), .B(n9402), .Z(n5143) );
  XOR U12314 ( .A(round_reg[456]), .B(n9463), .Z(n9402) );
  XNOR U12315 ( .A(n11706), .B(n11707), .Z(n9463) );
  AND U12316 ( .A(n10742), .B(n10741), .Z(n11705) );
  XNOR U12317 ( .A(round_reg[95]), .B(n10618), .Z(n10741) );
  IV U12318 ( .A(n11699), .Z(n10618) );
  XOR U12319 ( .A(n11708), .B(n11709), .Z(n11699) );
  XNOR U12320 ( .A(round_reg[1340]), .B(n11442), .Z(n10742) );
  IV U12321 ( .A(n9088), .Z(n11442) );
  XOR U12322 ( .A(n11710), .B(n11711), .Z(n9088) );
  XNOR U12323 ( .A(n11712), .B(n8338), .Z(n3788) );
  XNOR U12324 ( .A(round_reg[622]), .B(n9855), .Z(n8338) );
  IV U12325 ( .A(n11295), .Z(n9855) );
  ANDN U12326 ( .B(n10734), .A(n10733), .Z(n11712) );
  XNOR U12327 ( .A(round_reg[213]), .B(n9840), .Z(n10733) );
  XNOR U12328 ( .A(round_reg[1433]), .B(n9680), .Z(n10734) );
  XOR U12329 ( .A(n4749), .B(n11715), .Z(n11703) );
  XOR U12330 ( .A(n1736), .B(n10803), .Z(n11715) );
  XOR U12331 ( .A(n11716), .B(n8348), .Z(n10803) );
  XNOR U12332 ( .A(round_reg[386]), .B(n10379), .Z(n8348) );
  IV U12333 ( .A(n10522), .Z(n10379) );
  ANDN U12334 ( .B(n10731), .A(n10730), .Z(n11716) );
  XOR U12335 ( .A(round_reg[9]), .B(n10438), .Z(n10730) );
  XOR U12336 ( .A(n11386), .B(n11719), .Z(n10438) );
  XOR U12337 ( .A(n11720), .B(n11721), .Z(n11386) );
  XNOR U12338 ( .A(round_reg[1544]), .B(round_reg[1224]), .Z(n11721) );
  XOR U12339 ( .A(round_reg[264]), .B(n11722), .Z(n11720) );
  XOR U12340 ( .A(round_reg[904]), .B(round_reg[584]), .Z(n11722) );
  XOR U12341 ( .A(round_reg[1559]), .B(n9935), .Z(n10731) );
  XNOR U12342 ( .A(n11723), .B(n11724), .Z(n9935) );
  XNOR U12343 ( .A(n11725), .B(n8343), .Z(n1736) );
  XOR U12344 ( .A(round_reg[335]), .B(n10504), .Z(n8343) );
  ANDN U12345 ( .B(n10739), .A(n10738), .Z(n11725) );
  XNOR U12346 ( .A(round_reg[261]), .B(n9364), .Z(n10738) );
  IV U12347 ( .A(n11636), .Z(n9364) );
  XOR U12348 ( .A(n11726), .B(n11284), .Z(n11636) );
  XOR U12349 ( .A(n11727), .B(n11728), .Z(n11284) );
  XNOR U12350 ( .A(round_reg[325]), .B(round_reg[1285]), .Z(n11728) );
  XOR U12351 ( .A(round_reg[5]), .B(n11729), .Z(n11727) );
  XOR U12352 ( .A(round_reg[965]), .B(round_reg[645]), .Z(n11729) );
  XNOR U12353 ( .A(round_reg[1494]), .B(n10666), .Z(n10739) );
  XNOR U12354 ( .A(n11730), .B(n8352), .Z(n4749) );
  XOR U12355 ( .A(round_reg[554]), .B(n11048), .Z(n8352) );
  NOR U12356 ( .A(n10810), .B(n11555), .Z(n11730) );
  XNOR U12357 ( .A(n11731), .B(n10810), .Z(n10735) );
  XNOR U12358 ( .A(round_reg[154]), .B(n9607), .Z(n10810) );
  IV U12359 ( .A(n10670), .Z(n9607) );
  XOR U12360 ( .A(n11615), .B(n11732), .Z(n10670) );
  XOR U12361 ( .A(n11733), .B(n11734), .Z(n11615) );
  XNOR U12362 ( .A(round_reg[1498]), .B(round_reg[1178]), .Z(n11734) );
  XOR U12363 ( .A(round_reg[218]), .B(n11735), .Z(n11733) );
  XOR U12364 ( .A(round_reg[858]), .B(round_reg[538]), .Z(n11735) );
  AND U12365 ( .A(n8351), .B(n11555), .Z(n11731) );
  XOR U12366 ( .A(round_reg[1403]), .B(n11058), .Z(n11555) );
  IV U12367 ( .A(n11736), .Z(n11058) );
  XNOR U12368 ( .A(round_reg[963]), .B(n9103), .Z(n8351) );
  IV U12369 ( .A(n9826), .Z(n9103) );
  XOR U12370 ( .A(n11737), .B(n11738), .Z(n9826) );
  XOR U12371 ( .A(n11739), .B(n6270), .Z(out[1002]) );
  XOR U12372 ( .A(n9037), .B(n2312), .Z(n6270) );
  XNOR U12373 ( .A(n6150), .B(n6233), .Z(n2312) );
  XNOR U12374 ( .A(n11740), .B(n11741), .Z(n6233) );
  XOR U12375 ( .A(n2350), .B(n5495), .Z(n11741) );
  XOR U12376 ( .A(n11742), .B(n7918), .Z(n5495) );
  XNOR U12377 ( .A(round_reg[985]), .B(n9934), .Z(n7918) );
  XNOR U12378 ( .A(n11732), .B(n11475), .Z(n9934) );
  XOR U12379 ( .A(n11743), .B(n11744), .Z(n11475) );
  XNOR U12380 ( .A(round_reg[1560]), .B(round_reg[1240]), .Z(n11744) );
  XOR U12381 ( .A(round_reg[280]), .B(n11745), .Z(n11743) );
  XOR U12382 ( .A(round_reg[920]), .B(round_reg[600]), .Z(n11745) );
  XOR U12383 ( .A(n11746), .B(n11747), .Z(n11732) );
  XNOR U12384 ( .A(round_reg[1369]), .B(round_reg[1049]), .Z(n11747) );
  XOR U12385 ( .A(round_reg[409]), .B(n11748), .Z(n11746) );
  XOR U12386 ( .A(round_reg[89]), .B(round_reg[729]), .Z(n11748) );
  ANDN U12387 ( .B(n9046), .A(n7917), .Z(n11742) );
  XOR U12388 ( .A(round_reg[938]), .B(n10220), .Z(n7917) );
  XOR U12389 ( .A(round_reg[512]), .B(n11749), .Z(n9046) );
  XNOR U12390 ( .A(n11750), .B(n7922), .Z(n2350) );
  XNOR U12391 ( .A(round_reg[1153]), .B(n9779), .Z(n7922) );
  ANDN U12392 ( .B(n9042), .A(n7921), .Z(n11750) );
  XNOR U12393 ( .A(round_reg[770]), .B(n9859), .Z(n7921) );
  XOR U12394 ( .A(round_reg[408]), .B(n10881), .Z(n9042) );
  IV U12395 ( .A(n11302), .Z(n10881) );
  XOR U12396 ( .A(n11348), .B(n11724), .Z(n11302) );
  XNOR U12397 ( .A(n11753), .B(n11754), .Z(n11724) );
  XNOR U12398 ( .A(round_reg[23]), .B(round_reg[1303]), .Z(n11754) );
  XOR U12399 ( .A(round_reg[343]), .B(n11755), .Z(n11753) );
  XOR U12400 ( .A(round_reg[983]), .B(round_reg[663]), .Z(n11755) );
  XOR U12401 ( .A(n11756), .B(n11757), .Z(n11348) );
  XNOR U12402 ( .A(round_reg[1432]), .B(round_reg[1112]), .Z(n11757) );
  XOR U12403 ( .A(round_reg[152]), .B(n11758), .Z(n11756) );
  XOR U12404 ( .A(round_reg[792]), .B(round_reg[472]), .Z(n11758) );
  XOR U12405 ( .A(n3185), .B(n11759), .Z(n11740) );
  XNOR U12406 ( .A(n6322), .B(n7911), .Z(n11759) );
  XOR U12407 ( .A(n11760), .B(n7927), .Z(n7911) );
  XNOR U12408 ( .A(round_reg[1225]), .B(n9216), .Z(n7927) );
  ANDN U12409 ( .B(n9044), .A(n7926), .Z(n11760) );
  XNOR U12410 ( .A(round_reg[867]), .B(n10433), .Z(n7926) );
  IV U12411 ( .A(n11539), .Z(n10433) );
  XNOR U12412 ( .A(n11761), .B(n11762), .Z(n11539) );
  XOR U12413 ( .A(round_reg[478]), .B(n11763), .Z(n9044) );
  XNOR U12414 ( .A(n11764), .B(n7931), .Z(n6322) );
  XNOR U12415 ( .A(round_reg[1078]), .B(n9108), .Z(n7931) );
  XOR U12416 ( .A(n11765), .B(n11766), .Z(n11332) );
  XNOR U12417 ( .A(round_reg[1333]), .B(round_reg[1013]), .Z(n11766) );
  XOR U12418 ( .A(round_reg[373]), .B(n11767), .Z(n11765) );
  XOR U12419 ( .A(round_reg[693]), .B(round_reg[53]), .Z(n11767) );
  XNOR U12420 ( .A(n11768), .B(n11769), .Z(n10540) );
  XNOR U12421 ( .A(round_reg[1462]), .B(round_reg[1142]), .Z(n11769) );
  XOR U12422 ( .A(round_reg[182]), .B(n11770), .Z(n11768) );
  XOR U12423 ( .A(round_reg[822]), .B(round_reg[502]), .Z(n11770) );
  ANDN U12424 ( .B(n11634), .A(n7930), .Z(n11764) );
  XOR U12425 ( .A(n11771), .B(n7935), .Z(n3185) );
  XNOR U12426 ( .A(round_reg[1127]), .B(n10797), .Z(n7935) );
  IV U12427 ( .A(n10444), .Z(n10797) );
  XOR U12428 ( .A(n11772), .B(n11773), .Z(n10444) );
  ANDN U12429 ( .B(n9039), .A(n7934), .Z(n11771) );
  XNOR U12430 ( .A(round_reg[724]), .B(n9973), .Z(n7934) );
  IV U12431 ( .A(n11313), .Z(n9973) );
  XOR U12432 ( .A(round_reg[357]), .B(n9851), .Z(n9039) );
  XOR U12433 ( .A(n11774), .B(n11775), .Z(n6150) );
  XNOR U12434 ( .A(n5291), .B(n1942), .Z(n11775) );
  XNOR U12435 ( .A(n11776), .B(n9122), .Z(n1942) );
  NOR U12436 ( .A(n8041), .B(n9026), .Z(n11776) );
  XNOR U12437 ( .A(round_reg[282]), .B(n11346), .Z(n9026) );
  XOR U12438 ( .A(round_reg[1515]), .B(n10868), .Z(n8041) );
  XNOR U12439 ( .A(n11777), .B(n9128), .Z(n5291) );
  ANDN U12440 ( .B(n8033), .A(n9024), .Z(n11777) );
  XNOR U12441 ( .A(round_reg[116]), .B(n11443), .Z(n9024) );
  XNOR U12442 ( .A(round_reg[1297]), .B(n10359), .Z(n8033) );
  IV U12443 ( .A(n10629), .Z(n10359) );
  XOR U12444 ( .A(n11778), .B(n11779), .Z(n10629) );
  XNOR U12445 ( .A(n3697), .B(n11780), .Z(n11774) );
  XOR U12446 ( .A(n9117), .B(n4138), .Z(n11780) );
  XNOR U12447 ( .A(n11781), .B(n9130), .Z(n4138) );
  NOR U12448 ( .A(n8024), .B(n9034), .Z(n11781) );
  XNOR U12449 ( .A(round_reg[175]), .B(n10871), .Z(n9034) );
  XOR U12450 ( .A(n11782), .B(n11783), .Z(n10871) );
  XOR U12451 ( .A(round_reg[1360]), .B(n9447), .Z(n8024) );
  XNOR U12452 ( .A(n11784), .B(n9125), .Z(n9117) );
  AND U12453 ( .A(n8028), .B(n9126), .Z(n11784) );
  XOR U12454 ( .A(round_reg[30]), .B(n9635), .Z(n9126) );
  IV U12455 ( .A(n10453), .Z(n9635) );
  XNOR U12456 ( .A(n10943), .B(n11609), .Z(n10453) );
  XNOR U12457 ( .A(n11785), .B(n11786), .Z(n11609) );
  XNOR U12458 ( .A(round_reg[1374]), .B(round_reg[1054]), .Z(n11786) );
  XOR U12459 ( .A(round_reg[414]), .B(n11787), .Z(n11785) );
  XOR U12460 ( .A(round_reg[94]), .B(round_reg[734]), .Z(n11787) );
  XOR U12461 ( .A(n11788), .B(n11789), .Z(n10943) );
  XNOR U12462 ( .A(round_reg[1565]), .B(round_reg[1245]), .Z(n11789) );
  XOR U12463 ( .A(round_reg[285]), .B(n11790), .Z(n11788) );
  XOR U12464 ( .A(round_reg[925]), .B(round_reg[605]), .Z(n11790) );
  XOR U12465 ( .A(round_reg[1580]), .B(n10010), .Z(n8028) );
  XNOR U12466 ( .A(n11791), .B(n11792), .Z(n3697) );
  ANDN U12467 ( .B(n9032), .A(n8037), .Z(n11791) );
  XNOR U12468 ( .A(round_reg[1454]), .B(n11328), .Z(n8037) );
  XOR U12469 ( .A(n11793), .B(n7930), .Z(n9037) );
  XNOR U12470 ( .A(round_reg[646]), .B(n10674), .Z(n7930) );
  ANDN U12471 ( .B(n8972), .A(n11634), .Z(n11793) );
  XOR U12472 ( .A(round_reg[580]), .B(n9964), .Z(n11634) );
  XNOR U12473 ( .A(round_reg[235]), .B(n10868), .Z(n8972) );
  XOR U12474 ( .A(n11794), .B(n10586), .Z(n10868) );
  XNOR U12475 ( .A(n11795), .B(n11796), .Z(n10586) );
  XNOR U12476 ( .A(round_reg[1450]), .B(round_reg[1130]), .Z(n11796) );
  XOR U12477 ( .A(round_reg[170]), .B(n11797), .Z(n11795) );
  XOR U12478 ( .A(round_reg[810]), .B(round_reg[490]), .Z(n11797) );
  NOR U12479 ( .A(n5718), .B(n5716), .Z(n11739) );
  XNOR U12480 ( .A(n8887), .B(n5173), .Z(n5716) );
  XNOR U12481 ( .A(n11798), .B(n11799), .Z(n6537) );
  XNOR U12482 ( .A(n5521), .B(n2541), .Z(n11799) );
  XNOR U12483 ( .A(n11800), .B(n6594), .Z(n2541) );
  XOR U12484 ( .A(round_reg[907]), .B(n11125), .Z(n6594) );
  ANDN U12485 ( .B(n8892), .A(n8893), .Z(n11800) );
  XNOR U12486 ( .A(round_reg[145]), .B(n10762), .Z(n8893) );
  XNOR U12487 ( .A(n11801), .B(n11802), .Z(n10762) );
  XOR U12488 ( .A(round_reg[545]), .B(n10496), .Z(n8892) );
  XOR U12489 ( .A(n11803), .B(n6585), .Z(n5521) );
  XNOR U12490 ( .A(round_reg[803]), .B(n10676), .Z(n6585) );
  IV U12491 ( .A(n9899), .Z(n10676) );
  XOR U12492 ( .A(n11804), .B(n11805), .Z(n9899) );
  ANDN U12493 ( .B(n8934), .A(n11669), .Z(n11803) );
  XOR U12494 ( .A(n3486), .B(n11806), .Z(n11798) );
  XNOR U12495 ( .A(n8927), .B(n4849), .Z(n11806) );
  XNOR U12496 ( .A(n11807), .B(n6581), .Z(n4849) );
  XOR U12497 ( .A(round_reg[757]), .B(n9191), .Z(n6581) );
  ANDN U12498 ( .B(n8889), .A(n8890), .Z(n11807) );
  XNOR U12499 ( .A(round_reg[316]), .B(n10667), .Z(n8890) );
  XNOR U12500 ( .A(n11702), .B(n10997), .Z(n10667) );
  XNOR U12501 ( .A(n11808), .B(n11809), .Z(n10997) );
  XNOR U12502 ( .A(round_reg[1531]), .B(round_reg[1211]), .Z(n11809) );
  XOR U12503 ( .A(round_reg[251]), .B(n11810), .Z(n11808) );
  XOR U12504 ( .A(round_reg[891]), .B(round_reg[571]), .Z(n11810) );
  XOR U12505 ( .A(n11811), .B(n11812), .Z(n11702) );
  XNOR U12506 ( .A(round_reg[1340]), .B(round_reg[1020]), .Z(n11812) );
  XOR U12507 ( .A(round_reg[380]), .B(n11813), .Z(n11811) );
  XOR U12508 ( .A(round_reg[700]), .B(round_reg[60]), .Z(n11813) );
  XOR U12509 ( .A(round_reg[326]), .B(n10674), .Z(n8889) );
  XOR U12510 ( .A(n11814), .B(n6577), .Z(n8927) );
  XOR U12511 ( .A(round_reg[679]), .B(n10783), .Z(n6577) );
  IV U12512 ( .A(n9766), .Z(n10783) );
  XNOR U12513 ( .A(n11398), .B(n11815), .Z(n9766) );
  XOR U12514 ( .A(n11816), .B(n11817), .Z(n11398) );
  XNOR U12515 ( .A(round_reg[1574]), .B(round_reg[1254]), .Z(n11817) );
  XOR U12516 ( .A(round_reg[294]), .B(n11818), .Z(n11816) );
  XOR U12517 ( .A(round_reg[934]), .B(round_reg[614]), .Z(n11818) );
  NOR U12518 ( .A(n8884), .B(n8885), .Z(n11814) );
  XNOR U12519 ( .A(round_reg[204]), .B(n11819), .Z(n8885) );
  XNOR U12520 ( .A(round_reg[613]), .B(n9263), .Z(n8884) );
  IV U12521 ( .A(n9959), .Z(n9263) );
  XNOR U12522 ( .A(n11646), .B(n10933), .Z(n9959) );
  XNOR U12523 ( .A(n11820), .B(n11821), .Z(n10933) );
  XNOR U12524 ( .A(round_reg[357]), .B(round_reg[1317]), .Z(n11821) );
  XOR U12525 ( .A(round_reg[37]), .B(n11822), .Z(n11820) );
  XOR U12526 ( .A(round_reg[997]), .B(round_reg[677]), .Z(n11822) );
  XOR U12527 ( .A(n11823), .B(n11824), .Z(n11646) );
  XNOR U12528 ( .A(round_reg[1508]), .B(round_reg[1188]), .Z(n11824) );
  XOR U12529 ( .A(round_reg[228]), .B(n11825), .Z(n11823) );
  XOR U12530 ( .A(round_reg[868]), .B(round_reg[548]), .Z(n11825) );
  XNOR U12531 ( .A(n11826), .B(n6590), .Z(n3486) );
  XOR U12532 ( .A(round_reg[836]), .B(n9555), .Z(n6590) );
  IV U12533 ( .A(n9543), .Z(n9555) );
  XOR U12534 ( .A(n11827), .B(n11579), .Z(n9543) );
  XOR U12535 ( .A(n11828), .B(n11829), .Z(n11579) );
  XNOR U12536 ( .A(round_reg[131]), .B(round_reg[1091]), .Z(n11829) );
  XOR U12537 ( .A(round_reg[1411]), .B(n11830), .Z(n11828) );
  XOR U12538 ( .A(round_reg[771]), .B(round_reg[451]), .Z(n11830) );
  ANDN U12539 ( .B(n8881), .A(n8882), .Z(n11826) );
  XNOR U12540 ( .A(round_reg[86]), .B(n11151), .Z(n8882) );
  XOR U12541 ( .A(round_reg[511]), .B(n9614), .Z(n8881) );
  XOR U12542 ( .A(n11831), .B(n11380), .Z(n9614) );
  XNOR U12543 ( .A(n11832), .B(n11833), .Z(n11380) );
  XNOR U12544 ( .A(round_reg[1535]), .B(round_reg[1215]), .Z(n11833) );
  XOR U12545 ( .A(round_reg[255]), .B(n11834), .Z(n11832) );
  XOR U12546 ( .A(round_reg[895]), .B(round_reg[575]), .Z(n11834) );
  XNOR U12547 ( .A(n11835), .B(n11836), .Z(n6390) );
  XOR U12548 ( .A(n5483), .B(n3681), .Z(n11836) );
  XOR U12549 ( .A(n11837), .B(n11838), .Z(n3681) );
  ANDN U12550 ( .B(n6610), .A(n6611), .Z(n11837) );
  XNOR U12551 ( .A(n11839), .B(n8944), .Z(n5483) );
  ANDN U12552 ( .B(n6601), .A(n6602), .Z(n11839) );
  XNOR U12553 ( .A(round_reg[1046]), .B(n11151), .Z(n6602) );
  XOR U12554 ( .A(round_reg[1423]), .B(n10931), .Z(n6601) );
  XNOR U12555 ( .A(n4255), .B(n11840), .Z(n11835) );
  XOR U12556 ( .A(n5957), .B(n2140), .Z(n11840) );
  XOR U12557 ( .A(n11841), .B(n8941), .Z(n2140) );
  ANDN U12558 ( .B(n6614), .A(n6615), .Z(n11841) );
  XNOR U12559 ( .A(round_reg[1257]), .B(n11377), .Z(n6615) );
  XOR U12560 ( .A(round_reg[1330]), .B(n9522), .Z(n6614) );
  IV U12561 ( .A(n9861), .Z(n9522) );
  XNOR U12562 ( .A(n11842), .B(n11158), .Z(n9861) );
  XNOR U12563 ( .A(n11843), .B(n11844), .Z(n11158) );
  XNOR U12564 ( .A(round_reg[1585]), .B(round_reg[1265]), .Z(n11844) );
  XOR U12565 ( .A(round_reg[305]), .B(n11845), .Z(n11843) );
  XOR U12566 ( .A(round_reg[945]), .B(round_reg[625]), .Z(n11845) );
  XOR U12567 ( .A(n11846), .B(n8952), .Z(n5957) );
  NOR U12568 ( .A(n6618), .B(n6619), .Z(n11846) );
  XNOR U12569 ( .A(round_reg[1017]), .B(n11847), .Z(n6619) );
  XNOR U12570 ( .A(round_reg[1393]), .B(n9188), .Z(n6618) );
  XNOR U12571 ( .A(n11849), .B(n11850), .Z(n11070) );
  XNOR U12572 ( .A(round_reg[1457]), .B(round_reg[1137]), .Z(n11850) );
  XOR U12573 ( .A(round_reg[177]), .B(n11851), .Z(n11849) );
  XOR U12574 ( .A(round_reg[817]), .B(round_reg[497]), .Z(n11851) );
  XOR U12575 ( .A(n11852), .B(n8949), .Z(n4255) );
  ANDN U12576 ( .B(n6605), .A(n6606), .Z(n11852) );
  XNOR U12577 ( .A(round_reg[1095]), .B(n9548), .Z(n6606) );
  IV U12578 ( .A(n9633), .Z(n9548) );
  XOR U12579 ( .A(round_reg[1484]), .B(n10535), .Z(n6605) );
  IV U12580 ( .A(n11819), .Z(n10535) );
  XNOR U12581 ( .A(n11853), .B(n11854), .Z(n11819) );
  XNOR U12582 ( .A(n11855), .B(n8934), .Z(n8887) );
  XOR U12583 ( .A(round_reg[441]), .B(n11223), .Z(n8934) );
  ANDN U12584 ( .B(n11669), .A(n6584), .Z(n11855) );
  XOR U12585 ( .A(round_reg[1550]), .B(n10713), .Z(n6584) );
  XOR U12586 ( .A(n11856), .B(n11857), .Z(n10713) );
  XNOR U12587 ( .A(round_reg[0]), .B(n9374), .Z(n11669) );
  IV U12588 ( .A(n11275), .Z(n9374) );
  XOR U12589 ( .A(n10821), .B(n2105), .Z(n5718) );
  XNOR U12590 ( .A(n8333), .B(n9559), .Z(n2105) );
  XNOR U12591 ( .A(n11858), .B(n11859), .Z(n9559) );
  XOR U12592 ( .A(n5513), .B(n3607), .Z(n11859) );
  XOR U12593 ( .A(n11860), .B(n11861), .Z(n3607) );
  ANDN U12594 ( .B(n8458), .A(n8456), .Z(n11860) );
  XOR U12595 ( .A(round_reg[914]), .B(n10388), .Z(n8458) );
  XOR U12596 ( .A(n11801), .B(n11862), .Z(n10388) );
  XOR U12597 ( .A(n11863), .B(n11864), .Z(n11801) );
  XNOR U12598 ( .A(round_reg[1489]), .B(round_reg[1169]), .Z(n11864) );
  XOR U12599 ( .A(round_reg[209]), .B(n11865), .Z(n11863) );
  XOR U12600 ( .A(round_reg[849]), .B(round_reg[529]), .Z(n11865) );
  XOR U12601 ( .A(n11866), .B(n11867), .Z(n5513) );
  AND U12602 ( .A(n8454), .B(n8452), .Z(n11866) );
  XOR U12603 ( .A(round_reg[1193]), .B(n11136), .Z(n8452) );
  XNOR U12604 ( .A(round_reg[810]), .B(n10044), .Z(n8454) );
  IV U12605 ( .A(n10173), .Z(n10044) );
  XOR U12606 ( .A(n11868), .B(n11532), .Z(n10173) );
  XOR U12607 ( .A(n11869), .B(n11870), .Z(n11532) );
  XNOR U12608 ( .A(round_reg[1065]), .B(round_reg[105]), .Z(n11870) );
  XOR U12609 ( .A(round_reg[1385]), .B(n11871), .Z(n11869) );
  XOR U12610 ( .A(round_reg[745]), .B(round_reg[425]), .Z(n11871) );
  XOR U12611 ( .A(n6352), .B(n11872), .Z(n11858) );
  XOR U12612 ( .A(n2401), .B(n5660), .Z(n11872) );
  XNOR U12613 ( .A(n11873), .B(n10914), .Z(n5660) );
  ANDN U12614 ( .B(n9561), .A(n9562), .Z(n11873) );
  XOR U12615 ( .A(round_reg[843]), .B(n10626), .Z(n9562) );
  XOR U12616 ( .A(round_reg[1265]), .B(n9696), .Z(n9561) );
  IV U12617 ( .A(n11343), .Z(n9696) );
  XNOR U12618 ( .A(n11874), .B(n11625), .Z(n11343) );
  XNOR U12619 ( .A(n11875), .B(n11876), .Z(n11625) );
  XNOR U12620 ( .A(round_reg[1520]), .B(round_reg[1200]), .Z(n11876) );
  XOR U12621 ( .A(round_reg[240]), .B(n11877), .Z(n11875) );
  XOR U12622 ( .A(round_reg[880]), .B(round_reg[560]), .Z(n11877) );
  XNOR U12623 ( .A(n11878), .B(n10906), .Z(n2401) );
  ANDN U12624 ( .B(n8444), .A(n8442), .Z(n11878) );
  XOR U12625 ( .A(round_reg[1054]), .B(n10382), .Z(n8442) );
  XOR U12626 ( .A(round_reg[686]), .B(n9205), .Z(n8444) );
  XOR U12627 ( .A(n11879), .B(n10911), .Z(n6352) );
  NOR U12628 ( .A(n8446), .B(n8447), .Z(n11879) );
  XNOR U12629 ( .A(round_reg[764]), .B(n10878), .Z(n8447) );
  IV U12630 ( .A(n11138), .Z(n10878) );
  XOR U12631 ( .A(n11880), .B(n11881), .Z(n11138) );
  XNOR U12632 ( .A(round_reg[1103]), .B(n10931), .Z(n8446) );
  IV U12633 ( .A(n11882), .Z(n10931) );
  XOR U12634 ( .A(n11883), .B(n11884), .Z(n8333) );
  XNOR U12635 ( .A(n3792), .B(n5146), .Z(n11884) );
  XOR U12636 ( .A(n11885), .B(n9479), .Z(n5146) );
  XNOR U12637 ( .A(round_reg[455]), .B(n9633), .Z(n9479) );
  XOR U12638 ( .A(n11886), .B(n11887), .Z(n9633) );
  AND U12639 ( .A(n10828), .B(n10827), .Z(n11885) );
  XNOR U12640 ( .A(round_reg[94]), .B(n10382), .Z(n10827) );
  XNOR U12641 ( .A(n11407), .B(n11888), .Z(n10382) );
  XOR U12642 ( .A(n11889), .B(n11890), .Z(n11407) );
  XNOR U12643 ( .A(round_reg[29]), .B(round_reg[1309]), .Z(n11890) );
  XOR U12644 ( .A(round_reg[349]), .B(n11891), .Z(n11889) );
  XOR U12645 ( .A(round_reg[989]), .B(round_reg[669]), .Z(n11891) );
  XNOR U12646 ( .A(round_reg[1339]), .B(n11545), .Z(n10828) );
  XNOR U12647 ( .A(n11892), .B(n8391), .Z(n3792) );
  XOR U12648 ( .A(round_reg[621]), .B(n9923), .Z(n8391) );
  XOR U12649 ( .A(n10279), .B(n11893), .Z(n9923) );
  XOR U12650 ( .A(n11894), .B(n11895), .Z(n10279) );
  XNOR U12651 ( .A(round_reg[1325]), .B(round_reg[1005]), .Z(n11895) );
  XOR U12652 ( .A(round_reg[365]), .B(n11896), .Z(n11894) );
  XOR U12653 ( .A(round_reg[685]), .B(round_reg[45]), .Z(n11896) );
  ANDN U12654 ( .B(n10820), .A(n10819), .Z(n11892) );
  XNOR U12655 ( .A(round_reg[212]), .B(n9909), .Z(n10819) );
  XNOR U12656 ( .A(round_reg[1432]), .B(n9753), .Z(n10820) );
  XOR U12657 ( .A(n5110), .B(n11897), .Z(n11883) );
  XOR U12658 ( .A(n1741), .B(n10888), .Z(n11897) );
  XOR U12659 ( .A(n11898), .B(n8400), .Z(n10888) );
  XNOR U12660 ( .A(round_reg[385]), .B(n10454), .Z(n8400) );
  IV U12661 ( .A(n10615), .Z(n10454) );
  XNOR U12662 ( .A(n11379), .B(n11899), .Z(n10615) );
  XOR U12663 ( .A(n11900), .B(n11901), .Z(n11379) );
  XNOR U12664 ( .A(round_reg[1280]), .B(round_reg[0]), .Z(n11901) );
  XOR U12665 ( .A(round_reg[320]), .B(n11902), .Z(n11900) );
  XOR U12666 ( .A(round_reg[960]), .B(round_reg[640]), .Z(n11902) );
  AND U12667 ( .A(n10817), .B(n10816), .Z(n11898) );
  XOR U12668 ( .A(n11570), .B(n11903), .Z(n10492) );
  XOR U12669 ( .A(n11904), .B(n11905), .Z(n11570) );
  XNOR U12670 ( .A(round_reg[1352]), .B(round_reg[1032]), .Z(n11905) );
  XOR U12671 ( .A(round_reg[392]), .B(n11906), .Z(n11904) );
  XOR U12672 ( .A(round_reg[72]), .B(round_reg[712]), .Z(n11906) );
  XNOR U12673 ( .A(round_reg[1558]), .B(n10960), .Z(n10817) );
  IV U12674 ( .A(n10021), .Z(n10960) );
  XOR U12675 ( .A(n11907), .B(n11908), .Z(n10021) );
  XOR U12676 ( .A(n11909), .B(n8394), .Z(n1741) );
  XNOR U12677 ( .A(round_reg[334]), .B(n9981), .Z(n8394) );
  IV U12678 ( .A(n11199), .Z(n9981) );
  XNOR U12679 ( .A(n11677), .B(n11910), .Z(n11199) );
  XOR U12680 ( .A(n11911), .B(n11912), .Z(n11677) );
  XNOR U12681 ( .A(round_reg[1549]), .B(round_reg[1229]), .Z(n11912) );
  XOR U12682 ( .A(round_reg[269]), .B(n11913), .Z(n11911) );
  XOR U12683 ( .A(round_reg[909]), .B(round_reg[589]), .Z(n11913) );
  XOR U12684 ( .A(round_reg[260]), .B(n9964), .Z(n10824) );
  XOR U12685 ( .A(n11914), .B(n11915), .Z(n9964) );
  XNOR U12686 ( .A(round_reg[1493]), .B(n9840), .Z(n10825) );
  XNOR U12687 ( .A(n11916), .B(n8404), .Z(n5110) );
  XOR U12688 ( .A(round_reg[553]), .B(n11136), .Z(n8404) );
  NOR U12689 ( .A(n10895), .B(n11687), .Z(n11916) );
  XNOR U12690 ( .A(n11917), .B(n10895), .Z(n10821) );
  XNOR U12691 ( .A(round_reg[153]), .B(n9680), .Z(n10895) );
  IV U12692 ( .A(n10041), .Z(n9680) );
  XNOR U12693 ( .A(n11918), .B(n11919), .Z(n10041) );
  AND U12694 ( .A(n8403), .B(n11687), .Z(n11917) );
  XOR U12695 ( .A(round_reg[1402]), .B(n11146), .Z(n11687) );
  IV U12696 ( .A(n11920), .Z(n11146) );
  XOR U12697 ( .A(round_reg[962]), .B(n9187), .Z(n8403) );
  XOR U12698 ( .A(n11921), .B(n11751), .Z(n9187) );
  XNOR U12699 ( .A(n11922), .B(n11923), .Z(n11751) );
  XNOR U12700 ( .A(round_reg[1537]), .B(round_reg[1217]), .Z(n11923) );
  XOR U12701 ( .A(round_reg[257]), .B(n11924), .Z(n11922) );
  XOR U12702 ( .A(round_reg[897]), .B(round_reg[577]), .Z(n11924) );
  XOR U12703 ( .A(n11925), .B(n6281), .Z(out[1001]) );
  XOR U12704 ( .A(n9120), .B(n2319), .Z(n6281) );
  XNOR U12705 ( .A(n9813), .B(n6238), .Z(n2319) );
  XNOR U12706 ( .A(n11926), .B(n11927), .Z(n6238) );
  XOR U12707 ( .A(n2357), .B(n5499), .Z(n11927) );
  XOR U12708 ( .A(n11928), .B(n8026), .Z(n5499) );
  XOR U12709 ( .A(round_reg[984]), .B(n10020), .Z(n8026) );
  XOR U12710 ( .A(n11584), .B(n11918), .Z(n10020) );
  XOR U12711 ( .A(n11929), .B(n11930), .Z(n11918) );
  XNOR U12712 ( .A(round_reg[1368]), .B(round_reg[1048]), .Z(n11930) );
  XOR U12713 ( .A(round_reg[408]), .B(n11931), .Z(n11929) );
  XOR U12714 ( .A(round_reg[88]), .B(round_reg[728]), .Z(n11931) );
  XOR U12715 ( .A(n11932), .B(n11933), .Z(n11584) );
  XNOR U12716 ( .A(round_reg[1559]), .B(round_reg[1239]), .Z(n11933) );
  XOR U12717 ( .A(round_reg[279]), .B(n11934), .Z(n11932) );
  XOR U12718 ( .A(round_reg[919]), .B(round_reg[599]), .Z(n11934) );
  ANDN U12719 ( .B(n9130), .A(n8025), .Z(n11928) );
  XNOR U12720 ( .A(round_reg[937]), .B(n9974), .Z(n8025) );
  IV U12721 ( .A(n11377), .Z(n9974) );
  XOR U12722 ( .A(n10585), .B(n11935), .Z(n11377) );
  XOR U12723 ( .A(n11936), .B(n11937), .Z(n10585) );
  XNOR U12724 ( .A(round_reg[1321]), .B(round_reg[1001]), .Z(n11937) );
  XOR U12725 ( .A(round_reg[361]), .B(n11938), .Z(n11936) );
  XOR U12726 ( .A(round_reg[681]), .B(round_reg[41]), .Z(n11938) );
  XOR U12727 ( .A(round_reg[575]), .B(n9854), .Z(n9130) );
  XNOR U12728 ( .A(n11939), .B(n8030), .Z(n2357) );
  XNOR U12729 ( .A(round_reg[1152]), .B(n9196), .Z(n8030) );
  IV U12730 ( .A(n11749), .Z(n9196) );
  ANDN U12731 ( .B(n9125), .A(n8029), .Z(n11939) );
  XNOR U12732 ( .A(round_reg[769]), .B(n10015), .Z(n8029) );
  IV U12733 ( .A(n9444), .Z(n10015) );
  XOR U12734 ( .A(n11940), .B(n11941), .Z(n9444) );
  XOR U12735 ( .A(round_reg[407]), .B(n11063), .Z(n9125) );
  XNOR U12736 ( .A(n11908), .B(n11476), .Z(n11063) );
  XNOR U12737 ( .A(n11942), .B(n11943), .Z(n11476) );
  XNOR U12738 ( .A(round_reg[1431]), .B(round_reg[1111]), .Z(n11943) );
  XOR U12739 ( .A(round_reg[151]), .B(n11944), .Z(n11942) );
  XOR U12740 ( .A(round_reg[791]), .B(round_reg[471]), .Z(n11944) );
  XOR U12741 ( .A(n11945), .B(n11946), .Z(n11908) );
  XNOR U12742 ( .A(round_reg[22]), .B(round_reg[1302]), .Z(n11946) );
  XOR U12743 ( .A(round_reg[342]), .B(n11947), .Z(n11945) );
  XOR U12744 ( .A(round_reg[982]), .B(round_reg[662]), .Z(n11947) );
  XOR U12745 ( .A(n3188), .B(n11948), .Z(n11926) );
  XNOR U12746 ( .A(n6366), .B(n8019), .Z(n11948) );
  XOR U12747 ( .A(n11949), .B(n8035), .Z(n8019) );
  XNOR U12748 ( .A(round_reg[1224]), .B(n11950), .Z(n8035) );
  ANDN U12749 ( .B(n9128), .A(n8034), .Z(n11949) );
  XNOR U12750 ( .A(round_reg[866]), .B(n10442), .Z(n8034) );
  IV U12751 ( .A(n11670), .Z(n10442) );
  XOR U12752 ( .A(n11951), .B(n11464), .Z(n11670) );
  XOR U12753 ( .A(n11952), .B(n11953), .Z(n11464) );
  XNOR U12754 ( .A(round_reg[1441]), .B(round_reg[1121]), .Z(n11953) );
  XOR U12755 ( .A(round_reg[161]), .B(n11954), .Z(n11952) );
  XOR U12756 ( .A(round_reg[801]), .B(round_reg[481]), .Z(n11954) );
  XOR U12757 ( .A(round_reg[477]), .B(n9367), .Z(n9128) );
  XNOR U12758 ( .A(n11955), .B(n11956), .Z(n9367) );
  XNOR U12759 ( .A(n11957), .B(n8039), .Z(n6366) );
  XNOR U12760 ( .A(round_reg[1077]), .B(n9191), .Z(n8039) );
  XOR U12761 ( .A(n11958), .B(n11959), .Z(n11014) );
  XNOR U12762 ( .A(round_reg[1461]), .B(round_reg[1141]), .Z(n11959) );
  XOR U12763 ( .A(round_reg[181]), .B(n11960), .Z(n11958) );
  XOR U12764 ( .A(round_reg[821]), .B(round_reg[501]), .Z(n11960) );
  XNOR U12765 ( .A(n11961), .B(n11962), .Z(n11456) );
  XNOR U12766 ( .A(round_reg[1332]), .B(round_reg[1012]), .Z(n11962) );
  XOR U12767 ( .A(round_reg[372]), .B(n11963), .Z(n11961) );
  XOR U12768 ( .A(round_reg[692]), .B(round_reg[52]), .Z(n11963) );
  ANDN U12769 ( .B(n11792), .A(n8038), .Z(n11957) );
  XOR U12770 ( .A(n11964), .B(n9027), .Z(n3188) );
  IV U12771 ( .A(n8043), .Z(n9027) );
  XOR U12772 ( .A(round_reg[1126]), .B(n10441), .Z(n8043) );
  IV U12773 ( .A(n10503), .Z(n10441) );
  XNOR U12774 ( .A(n11965), .B(n11966), .Z(n10503) );
  ANDN U12775 ( .B(n9122), .A(n8042), .Z(n11964) );
  XNOR U12776 ( .A(round_reg[723]), .B(n9183), .Z(n8042) );
  XOR U12777 ( .A(round_reg[356]), .B(n9100), .Z(n9122) );
  XOR U12778 ( .A(n11761), .B(n11967), .Z(n9100) );
  XOR U12779 ( .A(n11968), .B(n11969), .Z(n11761) );
  XNOR U12780 ( .A(round_reg[1571]), .B(round_reg[1251]), .Z(n11969) );
  XOR U12781 ( .A(round_reg[291]), .B(n11970), .Z(n11968) );
  XOR U12782 ( .A(round_reg[931]), .B(round_reg[611]), .Z(n11970) );
  XOR U12783 ( .A(n11971), .B(n11972), .Z(n9813) );
  XNOR U12784 ( .A(n5293), .B(n1947), .Z(n11972) );
  XNOR U12785 ( .A(n11973), .B(n9155), .Z(n1947) );
  ANDN U12786 ( .B(n8092), .A(n9142), .Z(n11973) );
  XNOR U12787 ( .A(round_reg[281]), .B(n10216), .Z(n9142) );
  IV U12788 ( .A(n11103), .Z(n10216) );
  XNOR U12789 ( .A(round_reg[1514]), .B(n11048), .Z(n8092) );
  XNOR U12790 ( .A(n11974), .B(n9160), .Z(n5293) );
  ANDN U12791 ( .B(n8084), .A(n9140), .Z(n11974) );
  XNOR U12792 ( .A(round_reg[115]), .B(n9827), .Z(n9140) );
  XNOR U12793 ( .A(round_reg[1296]), .B(n10445), .Z(n8084) );
  IV U12794 ( .A(n10939), .Z(n10445) );
  XNOR U12795 ( .A(n11445), .B(n11802), .Z(n10939) );
  XNOR U12796 ( .A(n11975), .B(n11976), .Z(n11802) );
  XNOR U12797 ( .A(round_reg[1360]), .B(round_reg[1040]), .Z(n11976) );
  XOR U12798 ( .A(round_reg[400]), .B(n11977), .Z(n11975) );
  XOR U12799 ( .A(round_reg[80]), .B(round_reg[720]), .Z(n11977) );
  XOR U12800 ( .A(n11978), .B(n11979), .Z(n11445) );
  XNOR U12801 ( .A(round_reg[1551]), .B(round_reg[1231]), .Z(n11979) );
  XOR U12802 ( .A(round_reg[271]), .B(n11980), .Z(n11978) );
  XOR U12803 ( .A(round_reg[911]), .B(round_reg[591]), .Z(n11980) );
  XNOR U12804 ( .A(n3701), .B(n11981), .Z(n11971) );
  XOR U12805 ( .A(n9150), .B(n4140), .Z(n11981) );
  XNOR U12806 ( .A(n11982), .B(n9163), .Z(n4140) );
  NOR U12807 ( .A(n8075), .B(n9162), .Z(n11982) );
  XNOR U12808 ( .A(round_reg[174]), .B(n11051), .Z(n9162) );
  XOR U12809 ( .A(round_reg[1359]), .B(n9380), .Z(n8075) );
  IV U12810 ( .A(n9969), .Z(n9380) );
  XNOR U12811 ( .A(n11983), .B(n11857), .Z(n9969) );
  XNOR U12812 ( .A(n11984), .B(n11985), .Z(n11857) );
  XNOR U12813 ( .A(round_reg[14]), .B(round_reg[1294]), .Z(n11985) );
  XOR U12814 ( .A(round_reg[334]), .B(n11986), .Z(n11984) );
  XOR U12815 ( .A(round_reg[974]), .B(round_reg[654]), .Z(n11986) );
  XNOR U12816 ( .A(n11987), .B(n9158), .Z(n9150) );
  ANDN U12817 ( .B(n8079), .A(n9135), .Z(n11987) );
  XNOR U12818 ( .A(round_reg[29]), .B(n9708), .Z(n9135) );
  IV U12819 ( .A(n10517), .Z(n9708) );
  XOR U12820 ( .A(n11988), .B(n11989), .Z(n10517) );
  XNOR U12821 ( .A(round_reg[1579]), .B(n11596), .Z(n8079) );
  XNOR U12822 ( .A(n11990), .B(n11991), .Z(n3701) );
  ANDN U12823 ( .B(n8088), .A(n9138), .Z(n11990) );
  XNOR U12824 ( .A(round_reg[1453]), .B(n11140), .Z(n8088) );
  XOR U12825 ( .A(n11992), .B(n8038), .Z(n9120) );
  XNOR U12826 ( .A(round_reg[645]), .B(n10763), .Z(n8038) );
  NOR U12827 ( .A(n9032), .B(n11792), .Z(n11992) );
  XOR U12828 ( .A(round_reg[579]), .B(n9702), .Z(n11792) );
  XOR U12829 ( .A(n11375), .B(n11993), .Z(n11048) );
  XOR U12830 ( .A(n11994), .B(n11995), .Z(n11375) );
  XNOR U12831 ( .A(round_reg[1578]), .B(round_reg[1258]), .Z(n11995) );
  XOR U12832 ( .A(round_reg[298]), .B(n11996), .Z(n11994) );
  XOR U12833 ( .A(round_reg[938]), .B(round_reg[618]), .Z(n11996) );
  NOR U12834 ( .A(n5722), .B(n5720), .Z(n11925) );
  XNOR U12835 ( .A(n8946), .B(n5176), .Z(n5720) );
  XOR U12836 ( .A(n11997), .B(n6571), .Z(n5176) );
  XNOR U12837 ( .A(n11998), .B(n11999), .Z(n6571) );
  XNOR U12838 ( .A(n5895), .B(n2552), .Z(n11999) );
  XNOR U12839 ( .A(n12000), .B(n6620), .Z(n2552) );
  XOR U12840 ( .A(round_reg[906]), .B(n9087), .Z(n6620) );
  IV U12841 ( .A(n11156), .Z(n9087) );
  XOR U12842 ( .A(n11569), .B(n12001), .Z(n11156) );
  XOR U12843 ( .A(n12002), .B(n12003), .Z(n11569) );
  XNOR U12844 ( .A(round_reg[1481]), .B(round_reg[1161]), .Z(n12003) );
  XOR U12845 ( .A(round_reg[201]), .B(n12004), .Z(n12002) );
  XOR U12846 ( .A(round_reg[841]), .B(round_reg[521]), .Z(n12004) );
  ANDN U12847 ( .B(n8951), .A(n8952), .Z(n12000) );
  XNOR U12848 ( .A(round_reg[144]), .B(n10844), .Z(n8952) );
  XNOR U12849 ( .A(n12005), .B(n12006), .Z(n10844) );
  XOR U12850 ( .A(round_reg[544]), .B(n10581), .Z(n8951) );
  XNOR U12851 ( .A(n12007), .B(n6612), .Z(n5895) );
  XOR U12852 ( .A(round_reg[802]), .B(n9968), .Z(n6612) );
  IV U12853 ( .A(n11299), .Z(n9968) );
  XNOR U12854 ( .A(n12008), .B(n11417), .Z(n11299) );
  XNOR U12855 ( .A(n12009), .B(n12010), .Z(n11417) );
  XNOR U12856 ( .A(round_reg[1377]), .B(round_reg[1057]), .Z(n12010) );
  XOR U12857 ( .A(round_reg[417]), .B(n12011), .Z(n12009) );
  XOR U12858 ( .A(round_reg[97]), .B(round_reg[737]), .Z(n12011) );
  ANDN U12859 ( .B(n8994), .A(n11838), .Z(n12007) );
  XOR U12860 ( .A(n3489), .B(n12012), .Z(n11998) );
  XNOR U12861 ( .A(n8987), .B(n4852), .Z(n12012) );
  XNOR U12862 ( .A(n12013), .B(n6607), .Z(n4852) );
  XOR U12863 ( .A(round_reg[756]), .B(n11443), .Z(n6607) );
  ANDN U12864 ( .B(n8948), .A(n8949), .Z(n12013) );
  XNOR U12865 ( .A(round_reg[315]), .B(n10440), .Z(n8949) );
  XOR U12866 ( .A(round_reg[325]), .B(n10763), .Z(n8948) );
  XOR U12867 ( .A(n11827), .B(n12014), .Z(n10763) );
  XOR U12868 ( .A(n12015), .B(n12016), .Z(n11827) );
  XNOR U12869 ( .A(round_reg[1540]), .B(round_reg[1220]), .Z(n12016) );
  XOR U12870 ( .A(round_reg[260]), .B(n12017), .Z(n12015) );
  XOR U12871 ( .A(round_reg[900]), .B(round_reg[580]), .Z(n12017) );
  XOR U12872 ( .A(n12018), .B(n6603), .Z(n8987) );
  XNOR U12873 ( .A(round_reg[678]), .B(n10883), .Z(n6603) );
  ANDN U12874 ( .B(n8943), .A(n8944), .Z(n12018) );
  XOR U12875 ( .A(round_reg[203]), .B(n10626), .Z(n8944) );
  XOR U12876 ( .A(round_reg[612]), .B(n10431), .Z(n8943) );
  XNOR U12877 ( .A(n12019), .B(n6616), .Z(n3489) );
  XOR U12878 ( .A(round_reg[835]), .B(n9636), .Z(n6616) );
  XOR U12879 ( .A(n12020), .B(n11718), .Z(n9636) );
  XNOR U12880 ( .A(n12021), .B(n12022), .Z(n11718) );
  XNOR U12881 ( .A(round_reg[130]), .B(round_reg[1090]), .Z(n12022) );
  XOR U12882 ( .A(round_reg[1410]), .B(n12023), .Z(n12021) );
  XOR U12883 ( .A(round_reg[770]), .B(round_reg[450]), .Z(n12023) );
  ANDN U12884 ( .B(n8940), .A(n8941), .Z(n12019) );
  XNOR U12885 ( .A(round_reg[85]), .B(n12024), .Z(n8941) );
  XOR U12886 ( .A(round_reg[510]), .B(n9688), .Z(n8940) );
  XOR U12887 ( .A(n12025), .B(n12026), .Z(n9688) );
  IV U12888 ( .A(n6394), .Z(n11997) );
  XNOR U12889 ( .A(n12027), .B(n12028), .Z(n6394) );
  XOR U12890 ( .A(n5488), .B(n3687), .Z(n12028) );
  AND U12891 ( .A(n6632), .B(n6631), .Z(n12029) );
  XNOR U12892 ( .A(round_reg[1184]), .B(n10581), .Z(n6632) );
  IV U12893 ( .A(n9824), .Z(n10581) );
  XOR U12894 ( .A(n12031), .B(n12032), .Z(n11416) );
  XNOR U12895 ( .A(round_reg[1568]), .B(round_reg[1248]), .Z(n12032) );
  XOR U12896 ( .A(round_reg[288]), .B(n12033), .Z(n12031) );
  XOR U12897 ( .A(round_reg[928]), .B(round_reg[608]), .Z(n12033) );
  XNOR U12898 ( .A(n12034), .B(n12035), .Z(n11709) );
  XNOR U12899 ( .A(round_reg[1439]), .B(round_reg[1119]), .Z(n12035) );
  XOR U12900 ( .A(round_reg[159]), .B(n12036), .Z(n12034) );
  XOR U12901 ( .A(round_reg[799]), .B(round_reg[479]), .Z(n12036) );
  XNOR U12902 ( .A(n12037), .B(n9004), .Z(n5488) );
  ANDN U12903 ( .B(n6640), .A(n6641), .Z(n12037) );
  XNOR U12904 ( .A(round_reg[1045]), .B(n12024), .Z(n6641) );
  XOR U12905 ( .A(round_reg[1422]), .B(n10529), .Z(n6640) );
  XNOR U12906 ( .A(n4260), .B(n12038), .Z(n12027) );
  XOR U12907 ( .A(n5962), .B(n2144), .Z(n12038) );
  XNOR U12908 ( .A(n12039), .B(n9001), .Z(n2144) );
  ANDN U12909 ( .B(n6636), .A(n6637), .Z(n12039) );
  XNOR U12910 ( .A(round_reg[1256]), .B(n12040), .Z(n6637) );
  XOR U12911 ( .A(round_reg[1329]), .B(n9601), .Z(n6636) );
  IV U12912 ( .A(n11458), .Z(n9601) );
  XOR U12913 ( .A(n12041), .B(n11235), .Z(n11458) );
  XOR U12914 ( .A(n12042), .B(n12043), .Z(n11235) );
  XNOR U12915 ( .A(round_reg[1584]), .B(round_reg[1264]), .Z(n12043) );
  XOR U12916 ( .A(round_reg[304]), .B(n12044), .Z(n12042) );
  XOR U12917 ( .A(round_reg[944]), .B(round_reg[624]), .Z(n12044) );
  XOR U12918 ( .A(n12045), .B(n9012), .Z(n5962) );
  NOR U12919 ( .A(n6627), .B(n6628), .Z(n12045) );
  XNOR U12920 ( .A(round_reg[1016]), .B(n12046), .Z(n6628) );
  XNOR U12921 ( .A(round_reg[1392]), .B(n9606), .Z(n6627) );
  XOR U12922 ( .A(n12047), .B(n9009), .Z(n4260) );
  ANDN U12923 ( .B(n6644), .A(n6646), .Z(n12047) );
  XNOR U12924 ( .A(round_reg[1094]), .B(n9628), .Z(n6646) );
  XOR U12925 ( .A(round_reg[1483]), .B(n10626), .Z(n6644) );
  XOR U12926 ( .A(n12048), .B(n10852), .Z(n10626) );
  XNOR U12927 ( .A(n12049), .B(n12050), .Z(n10852) );
  XNOR U12928 ( .A(round_reg[138]), .B(round_reg[1098]), .Z(n12050) );
  XOR U12929 ( .A(round_reg[1418]), .B(n12051), .Z(n12049) );
  XOR U12930 ( .A(round_reg[778]), .B(round_reg[458]), .Z(n12051) );
  XNOR U12931 ( .A(n12052), .B(n8994), .Z(n8946) );
  XOR U12932 ( .A(round_reg[440]), .B(n11308), .Z(n8994) );
  ANDN U12933 ( .B(n11838), .A(n6610), .Z(n12052) );
  XOR U12934 ( .A(round_reg[1549]), .B(n10802), .Z(n6610) );
  XOR U12935 ( .A(n12053), .B(n12054), .Z(n10802) );
  XNOR U12936 ( .A(round_reg[63]), .B(n9445), .Z(n11838) );
  IV U12937 ( .A(n11341), .Z(n9445) );
  XOR U12938 ( .A(n10907), .B(n2108), .Z(n5722) );
  XNOR U12939 ( .A(n8385), .B(n9640), .Z(n2108) );
  XNOR U12940 ( .A(n12055), .B(n12056), .Z(n9640) );
  XOR U12941 ( .A(n5517), .B(n3611), .Z(n12056) );
  XOR U12942 ( .A(n12057), .B(n12058), .Z(n3611) );
  ANDN U12943 ( .B(n8511), .A(n8509), .Z(n12057) );
  XOR U12944 ( .A(round_reg[913]), .B(n10500), .Z(n8511) );
  XOR U12945 ( .A(n12059), .B(n12005), .Z(n10500) );
  XOR U12946 ( .A(n12060), .B(n12061), .Z(n12005) );
  XNOR U12947 ( .A(round_reg[1488]), .B(round_reg[1168]), .Z(n12061) );
  XOR U12948 ( .A(round_reg[208]), .B(n12062), .Z(n12060) );
  XOR U12949 ( .A(round_reg[848]), .B(round_reg[528]), .Z(n12062) );
  XOR U12950 ( .A(n12063), .B(n12064), .Z(n5517) );
  ANDN U12951 ( .B(n8507), .A(n8505), .Z(n12063) );
  XNOR U12952 ( .A(round_reg[1192]), .B(n9977), .Z(n8505) );
  XOR U12953 ( .A(round_reg[809]), .B(n10284), .Z(n8507) );
  XNOR U12954 ( .A(n12065), .B(n11656), .Z(n10284) );
  XNOR U12955 ( .A(n12066), .B(n12067), .Z(n11656) );
  XNOR U12956 ( .A(round_reg[1064]), .B(round_reg[104]), .Z(n12067) );
  XOR U12957 ( .A(round_reg[1384]), .B(n12068), .Z(n12066) );
  XOR U12958 ( .A(round_reg[744]), .B(round_reg[424]), .Z(n12068) );
  XOR U12959 ( .A(n6356), .B(n12069), .Z(n12055) );
  XOR U12960 ( .A(n2408), .B(n5706), .Z(n12069) );
  XNOR U12961 ( .A(n12070), .B(n11098), .Z(n5706) );
  AND U12962 ( .A(n9642), .B(n9644), .Z(n12070) );
  XNOR U12963 ( .A(round_reg[842]), .B(n10710), .Z(n9644) );
  XOR U12964 ( .A(round_reg[1264]), .B(n9769), .Z(n9642) );
  IV U12965 ( .A(n11467), .Z(n9769) );
  XNOR U12966 ( .A(n11848), .B(n11783), .Z(n11467) );
  XNOR U12967 ( .A(n12071), .B(n12072), .Z(n11783) );
  XNOR U12968 ( .A(round_reg[1519]), .B(round_reg[1199]), .Z(n12072) );
  XOR U12969 ( .A(round_reg[239]), .B(n12073), .Z(n12071) );
  XOR U12970 ( .A(round_reg[879]), .B(round_reg[559]), .Z(n12073) );
  XOR U12971 ( .A(n12074), .B(n12075), .Z(n11848) );
  XNOR U12972 ( .A(round_reg[1328]), .B(round_reg[1008]), .Z(n12075) );
  XOR U12973 ( .A(round_reg[368]), .B(n12076), .Z(n12074) );
  XOR U12974 ( .A(round_reg[688]), .B(round_reg[48]), .Z(n12076) );
  XNOR U12975 ( .A(n12077), .B(n11090), .Z(n2408) );
  ANDN U12976 ( .B(n8497), .A(n8495), .Z(n12077) );
  XOR U12977 ( .A(round_reg[1053]), .B(n10457), .Z(n8495) );
  XOR U12978 ( .A(round_reg[685]), .B(n10873), .Z(n8497) );
  XOR U12979 ( .A(n12078), .B(n12079), .Z(n6356) );
  NOR U12980 ( .A(n8499), .B(n8501), .Z(n12078) );
  XNOR U12981 ( .A(round_reg[763]), .B(n11736), .Z(n8501) );
  XNOR U12982 ( .A(n10148), .B(n12080), .Z(n11736) );
  XOR U12983 ( .A(n12081), .B(n12082), .Z(n10148) );
  XNOR U12984 ( .A(round_reg[1467]), .B(round_reg[1147]), .Z(n12082) );
  XOR U12985 ( .A(round_reg[187]), .B(n12083), .Z(n12081) );
  XOR U12986 ( .A(round_reg[827]), .B(round_reg[507]), .Z(n12083) );
  XNOR U12987 ( .A(round_reg[1102]), .B(n10529), .Z(n8499) );
  XOR U12988 ( .A(n12084), .B(n12085), .Z(n8385) );
  XNOR U12989 ( .A(n3796), .B(n5149), .Z(n12085) );
  XNOR U12990 ( .A(n12086), .B(n9563), .Z(n5149) );
  XNOR U12991 ( .A(round_reg[454]), .B(n9628), .Z(n9563) );
  IV U12992 ( .A(n9706), .Z(n9628) );
  XOR U12993 ( .A(n12087), .B(n12014), .Z(n9706) );
  XNOR U12994 ( .A(n12088), .B(n12089), .Z(n12014) );
  XNOR U12995 ( .A(round_reg[1349]), .B(round_reg[1029]), .Z(n12089) );
  XOR U12996 ( .A(round_reg[389]), .B(n12090), .Z(n12088) );
  XOR U12997 ( .A(round_reg[709]), .B(round_reg[69]), .Z(n12090) );
  AND U12998 ( .A(n10914), .B(n10913), .Z(n12086) );
  XNOR U12999 ( .A(round_reg[93]), .B(n10457), .Z(n10913) );
  XNOR U13000 ( .A(n10856), .B(n11504), .Z(n10457) );
  XNOR U13001 ( .A(n12091), .B(n12092), .Z(n11504) );
  XNOR U13002 ( .A(round_reg[28]), .B(round_reg[1308]), .Z(n12092) );
  XOR U13003 ( .A(round_reg[348]), .B(n12093), .Z(n12091) );
  XOR U13004 ( .A(round_reg[988]), .B(round_reg[668]), .Z(n12093) );
  XOR U13005 ( .A(n12094), .B(n12095), .Z(n10856) );
  XNOR U13006 ( .A(round_reg[1437]), .B(round_reg[1117]), .Z(n12095) );
  XOR U13007 ( .A(round_reg[157]), .B(n12096), .Z(n12094) );
  XOR U13008 ( .A(round_reg[797]), .B(round_reg[477]), .Z(n12096) );
  XNOR U13009 ( .A(round_reg[1338]), .B(n11034), .Z(n10914) );
  XOR U13010 ( .A(n12097), .B(n8443), .Z(n3796) );
  IV U13011 ( .A(n11080), .Z(n8443) );
  XNOR U13012 ( .A(round_reg[620]), .B(n10010), .Z(n11080) );
  XNOR U13013 ( .A(n12098), .B(n11690), .Z(n10010) );
  XNOR U13014 ( .A(n12099), .B(n12100), .Z(n11690) );
  XNOR U13015 ( .A(round_reg[1515]), .B(round_reg[1195]), .Z(n12100) );
  XOR U13016 ( .A(round_reg[235]), .B(n12101), .Z(n12099) );
  XOR U13017 ( .A(round_reg[875]), .B(round_reg[555]), .Z(n12101) );
  ANDN U13018 ( .B(n10906), .A(n10905), .Z(n12097) );
  XNOR U13019 ( .A(round_reg[211]), .B(n9996), .Z(n10905) );
  XNOR U13020 ( .A(round_reg[1431]), .B(n11000), .Z(n10906) );
  XOR U13021 ( .A(n5522), .B(n12102), .Z(n12084) );
  XOR U13022 ( .A(n1746), .B(n11071), .Z(n12102) );
  XOR U13023 ( .A(n12103), .B(n8453), .Z(n11071) );
  XNOR U13024 ( .A(round_reg[384]), .B(n10518), .Z(n8453) );
  XOR U13025 ( .A(n12104), .B(n11752), .Z(n10518) );
  XNOR U13026 ( .A(n12105), .B(n12106), .Z(n11752) );
  XNOR U13027 ( .A(round_reg[128]), .B(round_reg[1088]), .Z(n12106) );
  XOR U13028 ( .A(round_reg[1408]), .B(n12107), .Z(n12105) );
  XOR U13029 ( .A(round_reg[768]), .B(round_reg[448]), .Z(n12107) );
  AND U13030 ( .A(n10902), .B(n11867), .Z(n12103) );
  IV U13031 ( .A(n10903), .Z(n11867) );
  XOR U13032 ( .A(round_reg[1557]), .B(n10531), .Z(n10903) );
  IV U13033 ( .A(n10164), .Z(n10531) );
  IV U13034 ( .A(n11082), .Z(n10902) );
  XNOR U13035 ( .A(round_reg[7]), .B(n11018), .Z(n11082) );
  XOR U13036 ( .A(n12108), .B(n11707), .Z(n11018) );
  XNOR U13037 ( .A(n12109), .B(n12110), .Z(n11707) );
  XNOR U13038 ( .A(round_reg[1351]), .B(round_reg[1031]), .Z(n12110) );
  XOR U13039 ( .A(round_reg[391]), .B(n12111), .Z(n12109) );
  XOR U13040 ( .A(round_reg[71]), .B(round_reg[711]), .Z(n12111) );
  XNOR U13041 ( .A(n12112), .B(n8448), .Z(n1746) );
  XOR U13042 ( .A(round_reg[333]), .B(n10042), .Z(n8448) );
  XNOR U13043 ( .A(n12113), .B(n12114), .Z(n11854) );
  XNOR U13044 ( .A(round_reg[1548]), .B(round_reg[1228]), .Z(n12114) );
  XOR U13045 ( .A(round_reg[268]), .B(n12115), .Z(n12113) );
  XOR U13046 ( .A(round_reg[908]), .B(round_reg[588]), .Z(n12115) );
  ANDN U13047 ( .B(n10911), .A(n10910), .Z(n12112) );
  XNOR U13048 ( .A(round_reg[259]), .B(n9523), .Z(n10910) );
  IV U13049 ( .A(n9702), .Z(n9523) );
  XOR U13050 ( .A(n12117), .B(n11470), .Z(n9702) );
  XOR U13051 ( .A(n12118), .B(n12119), .Z(n11470) );
  XNOR U13052 ( .A(round_reg[323]), .B(round_reg[1283]), .Z(n12119) );
  XOR U13053 ( .A(round_reg[3]), .B(n12120), .Z(n12118) );
  XOR U13054 ( .A(round_reg[963]), .B(round_reg[643]), .Z(n12120) );
  XNOR U13055 ( .A(round_reg[1492]), .B(n9909), .Z(n10911) );
  IV U13056 ( .A(n10837), .Z(n9909) );
  XNOR U13057 ( .A(n12121), .B(n8457), .Z(n5522) );
  XNOR U13058 ( .A(round_reg[552]), .B(n12122), .Z(n8457) );
  NOR U13059 ( .A(n11078), .B(n11861), .Z(n12121) );
  XNOR U13060 ( .A(n12123), .B(n11078), .Z(n10907) );
  XNOR U13061 ( .A(round_reg[152]), .B(n9753), .Z(n11078) );
  IV U13062 ( .A(n10840), .Z(n9753) );
  XNOR U13063 ( .A(n12124), .B(n12125), .Z(n10840) );
  AND U13064 ( .A(n8456), .B(n11861), .Z(n12123) );
  XOR U13065 ( .A(round_reg[1401]), .B(n11223), .Z(n11861) );
  XOR U13066 ( .A(n11108), .B(n10994), .Z(n11223) );
  XOR U13067 ( .A(n12126), .B(n12127), .Z(n10994) );
  XNOR U13068 ( .A(round_reg[1465]), .B(round_reg[1145]), .Z(n12127) );
  XOR U13069 ( .A(round_reg[185]), .B(n12128), .Z(n12126) );
  XOR U13070 ( .A(round_reg[825]), .B(round_reg[505]), .Z(n12128) );
  XNOR U13071 ( .A(n12129), .B(n12130), .Z(n11108) );
  XNOR U13072 ( .A(round_reg[1336]), .B(round_reg[1016]), .Z(n12130) );
  XOR U13073 ( .A(round_reg[376]), .B(n12131), .Z(n12129) );
  XOR U13074 ( .A(round_reg[696]), .B(round_reg[56]), .Z(n12131) );
  XOR U13075 ( .A(round_reg[961]), .B(n9966), .Z(n8456) );
  XOR U13076 ( .A(n12132), .B(n6286), .Z(out[1000]) );
  XOR U13077 ( .A(n9153), .B(n2330), .Z(n6286) );
  XNOR U13078 ( .A(n9884), .B(n6243), .Z(n2330) );
  XNOR U13079 ( .A(n12133), .B(n12134), .Z(n6243) );
  XOR U13080 ( .A(n2364), .B(n5504), .Z(n12134) );
  XOR U13081 ( .A(n12135), .B(n9832), .Z(n5504) );
  IV U13082 ( .A(n8077), .Z(n9832) );
  XOR U13083 ( .A(round_reg[983]), .B(n10977), .Z(n8077) );
  ANDN U13084 ( .B(n9163), .A(n8076), .Z(n12135) );
  XNOR U13085 ( .A(round_reg[936]), .B(n10036), .Z(n8076) );
  IV U13086 ( .A(n12040), .Z(n10036) );
  XOR U13087 ( .A(n11772), .B(n12136), .Z(n12040) );
  XOR U13088 ( .A(n12137), .B(n12138), .Z(n11772) );
  XNOR U13089 ( .A(round_reg[1511]), .B(round_reg[1191]), .Z(n12138) );
  XOR U13090 ( .A(round_reg[231]), .B(n12139), .Z(n12137) );
  XOR U13091 ( .A(round_reg[871]), .B(round_reg[551]), .Z(n12139) );
  XNOR U13092 ( .A(round_reg[574]), .B(n9371), .Z(n9163) );
  XOR U13093 ( .A(n11701), .B(n12140), .Z(n9371) );
  XOR U13094 ( .A(n12141), .B(n12142), .Z(n11701) );
  XNOR U13095 ( .A(round_reg[1469]), .B(round_reg[1149]), .Z(n12142) );
  XOR U13096 ( .A(round_reg[189]), .B(n12143), .Z(n12141) );
  XOR U13097 ( .A(round_reg[829]), .B(round_reg[509]), .Z(n12143) );
  XNOR U13098 ( .A(n12144), .B(n8081), .Z(n2364) );
  XNOR U13099 ( .A(round_reg[1215]), .B(n12145), .Z(n8081) );
  ANDN U13100 ( .B(n9158), .A(n8080), .Z(n12144) );
  XNOR U13101 ( .A(round_reg[768]), .B(n9534), .Z(n8080) );
  XOR U13102 ( .A(round_reg[406]), .B(n11151), .Z(n9158) );
  IV U13103 ( .A(n11499), .Z(n11151) );
  XOR U13104 ( .A(n12146), .B(n11585), .Z(n11499) );
  XNOR U13105 ( .A(n12147), .B(n12148), .Z(n11585) );
  XNOR U13106 ( .A(round_reg[1430]), .B(round_reg[1110]), .Z(n12148) );
  XOR U13107 ( .A(round_reg[150]), .B(n12149), .Z(n12147) );
  XOR U13108 ( .A(round_reg[790]), .B(round_reg[470]), .Z(n12149) );
  XOR U13109 ( .A(n3191), .B(n12150), .Z(n12133) );
  XOR U13110 ( .A(n6416), .B(n8070), .Z(n12150) );
  XOR U13111 ( .A(n12151), .B(n8086), .Z(n8070) );
  XNOR U13112 ( .A(round_reg[1223]), .B(n9200), .Z(n8086) );
  IV U13113 ( .A(n9390), .Z(n9200) );
  XOR U13114 ( .A(n12087), .B(n11122), .Z(n9390) );
  XOR U13115 ( .A(n12152), .B(n12153), .Z(n11122) );
  XNOR U13116 ( .A(round_reg[327]), .B(round_reg[1287]), .Z(n12153) );
  XOR U13117 ( .A(round_reg[647]), .B(n12154), .Z(n12152) );
  XOR U13118 ( .A(round_reg[967]), .B(round_reg[7]), .Z(n12154) );
  XOR U13119 ( .A(n12155), .B(n12156), .Z(n12087) );
  XNOR U13120 ( .A(round_reg[1478]), .B(round_reg[1158]), .Z(n12156) );
  XOR U13121 ( .A(round_reg[198]), .B(n12157), .Z(n12155) );
  XOR U13122 ( .A(round_reg[838]), .B(round_reg[518]), .Z(n12157) );
  ANDN U13123 ( .B(n9160), .A(n8085), .Z(n12151) );
  XNOR U13124 ( .A(round_reg[865]), .B(n10496), .Z(n8085) );
  XOR U13125 ( .A(n11571), .B(n12158), .Z(n10496) );
  XOR U13126 ( .A(n12159), .B(n12160), .Z(n11571) );
  XNOR U13127 ( .A(round_reg[1440]), .B(round_reg[1120]), .Z(n12160) );
  XOR U13128 ( .A(round_reg[160]), .B(n12161), .Z(n12159) );
  XOR U13129 ( .A(round_reg[800]), .B(round_reg[480]), .Z(n12161) );
  XOR U13130 ( .A(round_reg[476]), .B(n11479), .Z(n9160) );
  XOR U13131 ( .A(n11406), .B(n12162), .Z(n11479) );
  XOR U13132 ( .A(n12163), .B(n12164), .Z(n11406) );
  XNOR U13133 ( .A(round_reg[1500]), .B(round_reg[1180]), .Z(n12164) );
  XOR U13134 ( .A(round_reg[220]), .B(n12165), .Z(n12163) );
  XOR U13135 ( .A(round_reg[860]), .B(round_reg[540]), .Z(n12165) );
  XOR U13136 ( .A(n12166), .B(n8090), .Z(n6416) );
  XNOR U13137 ( .A(round_reg[1076]), .B(n11443), .Z(n8090) );
  IV U13138 ( .A(n12167), .Z(n11443) );
  ANDN U13139 ( .B(n11991), .A(n8089), .Z(n12166) );
  XOR U13140 ( .A(n12168), .B(n8094), .Z(n3191) );
  XNOR U13141 ( .A(round_reg[1125]), .B(n10495), .Z(n8094) );
  IV U13142 ( .A(n10596), .Z(n10495) );
  XNOR U13143 ( .A(n11967), .B(n11657), .Z(n10596) );
  XNOR U13144 ( .A(n12169), .B(n12170), .Z(n11657) );
  XNOR U13145 ( .A(round_reg[1509]), .B(round_reg[1189]), .Z(n12170) );
  XOR U13146 ( .A(round_reg[229]), .B(n12171), .Z(n12169) );
  XOR U13147 ( .A(round_reg[869]), .B(round_reg[549]), .Z(n12171) );
  XOR U13148 ( .A(n12172), .B(n12173), .Z(n11967) );
  XNOR U13149 ( .A(round_reg[1060]), .B(round_reg[100]), .Z(n12173) );
  XOR U13150 ( .A(round_reg[1380]), .B(n12174), .Z(n12172) );
  XOR U13151 ( .A(round_reg[740]), .B(round_reg[420]), .Z(n12174) );
  ANDN U13152 ( .B(n9155), .A(n8093), .Z(n12168) );
  XNOR U13153 ( .A(round_reg[722]), .B(n9080), .Z(n8093) );
  IV U13154 ( .A(n11514), .Z(n9080) );
  XOR U13155 ( .A(n12059), .B(n12175), .Z(n11514) );
  XOR U13156 ( .A(n12176), .B(n12177), .Z(n12059) );
  XNOR U13157 ( .A(round_reg[17]), .B(round_reg[1297]), .Z(n12177) );
  XOR U13158 ( .A(round_reg[337]), .B(n12178), .Z(n12176) );
  XOR U13159 ( .A(round_reg[977]), .B(round_reg[657]), .Z(n12178) );
  XOR U13160 ( .A(round_reg[355]), .B(n11230), .Z(n9155) );
  XOR U13161 ( .A(n12179), .B(n12180), .Z(n9884) );
  XNOR U13162 ( .A(n5092), .B(n1952), .Z(n12180) );
  XNOR U13163 ( .A(n12181), .B(n8006), .Z(n1952) );
  XOR U13164 ( .A(round_reg[354]), .B(n10799), .Z(n8006) );
  ANDN U13165 ( .B(n9179), .A(n9178), .Z(n12181) );
  XNOR U13166 ( .A(round_reg[280]), .B(n10302), .Z(n9178) );
  XNOR U13167 ( .A(round_reg[1513]), .B(n11136), .Z(n9179) );
  XNOR U13168 ( .A(n12182), .B(n8142), .Z(n5092) );
  XOR U13169 ( .A(round_reg[475]), .B(n9527), .Z(n8142) );
  IV U13170 ( .A(n10588), .Z(n9527) );
  XNOR U13171 ( .A(n11503), .B(n11592), .Z(n10588) );
  XNOR U13172 ( .A(n12183), .B(n12184), .Z(n11592) );
  XNOR U13173 ( .A(round_reg[1370]), .B(round_reg[1050]), .Z(n12184) );
  XOR U13174 ( .A(round_reg[410]), .B(n12185), .Z(n12183) );
  XOR U13175 ( .A(round_reg[90]), .B(round_reg[730]), .Z(n12185) );
  XOR U13176 ( .A(n12186), .B(n12187), .Z(n11503) );
  XNOR U13177 ( .A(round_reg[1499]), .B(round_reg[1179]), .Z(n12187) );
  XOR U13178 ( .A(round_reg[219]), .B(n12188), .Z(n12186) );
  XOR U13179 ( .A(round_reg[859]), .B(round_reg[539]), .Z(n12188) );
  ANDN U13180 ( .B(n9176), .A(n9175), .Z(n12182) );
  XNOR U13181 ( .A(round_reg[114]), .B(n9896), .Z(n9175) );
  IV U13182 ( .A(n9104), .Z(n9896) );
  XOR U13183 ( .A(n12189), .B(n11874), .Z(n9104) );
  XOR U13184 ( .A(n12190), .B(n12191), .Z(n11874) );
  XNOR U13185 ( .A(round_reg[1329]), .B(round_reg[1009]), .Z(n12191) );
  XOR U13186 ( .A(round_reg[369]), .B(n12192), .Z(n12190) );
  XOR U13187 ( .A(round_reg[689]), .B(round_reg[49]), .Z(n12192) );
  XNOR U13188 ( .A(round_reg[1295]), .B(n10504), .Z(n9176) );
  XOR U13189 ( .A(n11547), .B(n12006), .Z(n10504) );
  XNOR U13190 ( .A(n12193), .B(n12194), .Z(n12006) );
  XNOR U13191 ( .A(round_reg[1359]), .B(round_reg[1039]), .Z(n12194) );
  XOR U13192 ( .A(round_reg[399]), .B(n12195), .Z(n12193) );
  XOR U13193 ( .A(round_reg[79]), .B(round_reg[719]), .Z(n12195) );
  XOR U13194 ( .A(n12196), .B(n12197), .Z(n11547) );
  XNOR U13195 ( .A(round_reg[1550]), .B(round_reg[1230]), .Z(n12197) );
  XOR U13196 ( .A(round_reg[270]), .B(n12198), .Z(n12196) );
  XOR U13197 ( .A(round_reg[910]), .B(round_reg[590]), .Z(n12198) );
  XOR U13198 ( .A(n3705), .B(n12199), .Z(n12179) );
  XNOR U13199 ( .A(n9227), .B(n4142), .Z(n12199) );
  XNOR U13200 ( .A(n12200), .B(n8016), .Z(n4142) );
  XOR U13201 ( .A(round_reg[573]), .B(n9451), .Z(n8016) );
  ANDN U13202 ( .B(n9817), .A(n9234), .Z(n12200) );
  XNOR U13203 ( .A(round_reg[173]), .B(n11140), .Z(n9234) );
  XOR U13204 ( .A(n12201), .B(n11714), .Z(n11140) );
  XNOR U13205 ( .A(n12202), .B(n12203), .Z(n11714) );
  XNOR U13206 ( .A(round_reg[1517]), .B(round_reg[1197]), .Z(n12203) );
  XOR U13207 ( .A(round_reg[237]), .B(n12204), .Z(n12202) );
  XOR U13208 ( .A(round_reg[877]), .B(round_reg[557]), .Z(n12204) );
  XNOR U13209 ( .A(round_reg[1358]), .B(n9456), .Z(n9817) );
  XOR U13210 ( .A(n12053), .B(n11446), .Z(n9456) );
  XNOR U13211 ( .A(n12205), .B(n12206), .Z(n11446) );
  XNOR U13212 ( .A(round_reg[1422]), .B(round_reg[1102]), .Z(n12206) );
  XOR U13213 ( .A(round_reg[142]), .B(n12207), .Z(n12205) );
  XOR U13214 ( .A(round_reg[782]), .B(round_reg[462]), .Z(n12207) );
  XOR U13215 ( .A(n12208), .B(n12209), .Z(n12053) );
  XNOR U13216 ( .A(round_reg[13]), .B(round_reg[1293]), .Z(n12209) );
  XOR U13217 ( .A(round_reg[333]), .B(n12210), .Z(n12208) );
  XOR U13218 ( .A(round_reg[973]), .B(round_reg[653]), .Z(n12210) );
  XOR U13219 ( .A(n12211), .B(n8012), .Z(n9227) );
  XOR U13220 ( .A(round_reg[405]), .B(n11228), .Z(n8012) );
  IV U13221 ( .A(n12024), .Z(n11228) );
  XNOR U13222 ( .A(n12212), .B(n12213), .Z(n12024) );
  NOR U13223 ( .A(n9169), .B(n9168), .Z(n12211) );
  XNOR U13224 ( .A(round_reg[28]), .B(n9778), .Z(n9168) );
  IV U13225 ( .A(n10610), .Z(n9778) );
  XNOR U13226 ( .A(n11201), .B(n11956), .Z(n10610) );
  XNOR U13227 ( .A(n12214), .B(n12215), .Z(n11956) );
  XNOR U13228 ( .A(round_reg[1372]), .B(round_reg[1052]), .Z(n12215) );
  XOR U13229 ( .A(round_reg[412]), .B(n12216), .Z(n12214) );
  XOR U13230 ( .A(round_reg[92]), .B(round_reg[732]), .Z(n12216) );
  XOR U13231 ( .A(n12217), .B(n12218), .Z(n11201) );
  XNOR U13232 ( .A(round_reg[1563]), .B(round_reg[1243]), .Z(n12218) );
  XOR U13233 ( .A(round_reg[283]), .B(n12219), .Z(n12217) );
  XOR U13234 ( .A(round_reg[923]), .B(round_reg[603]), .Z(n12219) );
  IV U13235 ( .A(n9820), .Z(n9169) );
  XOR U13236 ( .A(round_reg[1578]), .B(n10220), .Z(n9820) );
  XOR U13237 ( .A(n11038), .B(n12065), .Z(n10220) );
  XOR U13238 ( .A(n12220), .B(n12221), .Z(n12065) );
  XNOR U13239 ( .A(round_reg[1513]), .B(round_reg[1193]), .Z(n12221) );
  XOR U13240 ( .A(round_reg[233]), .B(n12222), .Z(n12220) );
  XOR U13241 ( .A(round_reg[873]), .B(round_reg[553]), .Z(n12222) );
  XOR U13242 ( .A(n12223), .B(n12224), .Z(n11038) );
  XNOR U13243 ( .A(round_reg[1322]), .B(round_reg[1002]), .Z(n12224) );
  XOR U13244 ( .A(round_reg[362]), .B(n12225), .Z(n12223) );
  XOR U13245 ( .A(round_reg[682]), .B(round_reg[42]), .Z(n12225) );
  XNOR U13246 ( .A(n12226), .B(n8002), .Z(n3705) );
  XOR U13247 ( .A(round_reg[577]), .B(n9676), .Z(n8002) );
  AND U13248 ( .A(n9172), .B(n9173), .Z(n12226) );
  XOR U13249 ( .A(round_reg[1452]), .B(n9986), .Z(n9173) );
  XNOR U13250 ( .A(n11376), .B(n11893), .Z(n9986) );
  XNOR U13251 ( .A(n12227), .B(n12228), .Z(n11893) );
  XNOR U13252 ( .A(round_reg[1516]), .B(round_reg[1196]), .Z(n12228) );
  XOR U13253 ( .A(round_reg[236]), .B(n12229), .Z(n12227) );
  XOR U13254 ( .A(round_reg[876]), .B(round_reg[556]), .Z(n12229) );
  XOR U13255 ( .A(n12230), .B(n12231), .Z(n11376) );
  XNOR U13256 ( .A(round_reg[107]), .B(round_reg[1067]), .Z(n12231) );
  XOR U13257 ( .A(round_reg[1387]), .B(n12232), .Z(n12230) );
  XOR U13258 ( .A(round_reg[747]), .B(round_reg[427]), .Z(n12232) );
  XOR U13259 ( .A(round_reg[232]), .B(n9977), .Z(n9172) );
  IV U13260 ( .A(n12122), .Z(n9977) );
  XNOR U13261 ( .A(n10846), .B(n11533), .Z(n12122) );
  XNOR U13262 ( .A(n12233), .B(n12234), .Z(n11533) );
  XNOR U13263 ( .A(round_reg[1576]), .B(round_reg[1256]), .Z(n12234) );
  XOR U13264 ( .A(round_reg[296]), .B(n12235), .Z(n12233) );
  XOR U13265 ( .A(round_reg[936]), .B(round_reg[616]), .Z(n12235) );
  XOR U13266 ( .A(n12236), .B(n12237), .Z(n10846) );
  XNOR U13267 ( .A(round_reg[1447]), .B(round_reg[1127]), .Z(n12237) );
  XOR U13268 ( .A(round_reg[167]), .B(n12238), .Z(n12236) );
  XOR U13269 ( .A(round_reg[807]), .B(round_reg[487]), .Z(n12238) );
  XOR U13270 ( .A(n12239), .B(n8089), .Z(n9153) );
  XNOR U13271 ( .A(round_reg[644]), .B(n10845), .Z(n8089) );
  ANDN U13272 ( .B(n9138), .A(n11991), .Z(n12239) );
  XOR U13273 ( .A(round_reg[578]), .B(n10999), .Z(n11991) );
  XNOR U13274 ( .A(round_reg[233]), .B(n11136), .Z(n9138) );
  XOR U13275 ( .A(n12240), .B(n12241), .Z(n11136) );
  NOR U13276 ( .A(n5726), .B(n5724), .Z(n12132) );
  XNOR U13277 ( .A(n9006), .B(n5179), .Z(n5724) );
  XNOR U13278 ( .A(n12242), .B(n12243), .Z(n6597) );
  XNOR U13279 ( .A(n6411), .B(n2559), .Z(n12243) );
  XNOR U13280 ( .A(n12244), .B(n6629), .Z(n2559) );
  XOR U13281 ( .A(round_reg[905]), .B(n9216), .Z(n6629) );
  IV U13282 ( .A(n11234), .Z(n9216) );
  XOR U13283 ( .A(n11706), .B(n10851), .Z(n11234) );
  XOR U13284 ( .A(n12245), .B(n12246), .Z(n10851) );
  XNOR U13285 ( .A(round_reg[329]), .B(round_reg[1289]), .Z(n12246) );
  XOR U13286 ( .A(round_reg[649]), .B(n12247), .Z(n12245) );
  XOR U13287 ( .A(round_reg[9]), .B(round_reg[969]), .Z(n12247) );
  XOR U13288 ( .A(n12248), .B(n12249), .Z(n11706) );
  XNOR U13289 ( .A(round_reg[1480]), .B(round_reg[1160]), .Z(n12249) );
  XOR U13290 ( .A(round_reg[200]), .B(n12250), .Z(n12248) );
  XOR U13291 ( .A(round_reg[840]), .B(round_reg[520]), .Z(n12250) );
  ANDN U13292 ( .B(n9011), .A(n9012), .Z(n12244) );
  XNOR U13293 ( .A(round_reg[143]), .B(n11882), .Z(n9012) );
  XNOR U13294 ( .A(n12251), .B(n11910), .Z(n11882) );
  XNOR U13295 ( .A(n12252), .B(n12253), .Z(n11910) );
  XNOR U13296 ( .A(round_reg[1358]), .B(round_reg[1038]), .Z(n12253) );
  XOR U13297 ( .A(round_reg[398]), .B(n12254), .Z(n12252) );
  XOR U13298 ( .A(round_reg[78]), .B(round_reg[718]), .Z(n12254) );
  XNOR U13299 ( .A(round_reg[543]), .B(n9894), .Z(n9011) );
  XNOR U13300 ( .A(n12255), .B(n6633), .Z(n6411) );
  XOR U13301 ( .A(round_reg[801]), .B(n10099), .Z(n6633) );
  IV U13302 ( .A(n11400), .Z(n10099) );
  XNOR U13303 ( .A(n11517), .B(n11011), .Z(n11400) );
  XNOR U13304 ( .A(n12256), .B(n12257), .Z(n11011) );
  XNOR U13305 ( .A(round_reg[1505]), .B(round_reg[1185]), .Z(n12257) );
  XOR U13306 ( .A(round_reg[225]), .B(n12258), .Z(n12256) );
  XOR U13307 ( .A(round_reg[865]), .B(round_reg[545]), .Z(n12258) );
  XOR U13308 ( .A(n12259), .B(n12260), .Z(n11517) );
  XNOR U13309 ( .A(round_reg[1376]), .B(round_reg[1056]), .Z(n12260) );
  XOR U13310 ( .A(round_reg[416]), .B(n12261), .Z(n12259) );
  XOR U13311 ( .A(round_reg[96]), .B(round_reg[736]), .Z(n12261) );
  AND U13312 ( .A(n9054), .B(n12030), .Z(n12255) );
  XOR U13313 ( .A(n3492), .B(n12262), .Z(n12242) );
  XNOR U13314 ( .A(n9047), .B(n4855), .Z(n12262) );
  XOR U13315 ( .A(n12263), .B(n6645), .Z(n4855) );
  XNOR U13316 ( .A(round_reg[755]), .B(n9827), .Z(n6645) );
  IV U13317 ( .A(n9366), .Z(n9827) );
  XOR U13318 ( .A(n12264), .B(n11693), .Z(n9366) );
  XOR U13319 ( .A(n12265), .B(n12266), .Z(n11693) );
  XNOR U13320 ( .A(round_reg[1330]), .B(round_reg[1010]), .Z(n12266) );
  XOR U13321 ( .A(round_reg[370]), .B(n12267), .Z(n12265) );
  XOR U13322 ( .A(round_reg[690]), .B(round_reg[50]), .Z(n12267) );
  ANDN U13323 ( .B(n9008), .A(n9009), .Z(n12263) );
  XNOR U13324 ( .A(round_reg[314]), .B(n10494), .Z(n9009) );
  IV U13325 ( .A(n10384), .Z(n10494) );
  XOR U13326 ( .A(round_reg[324]), .B(n10845), .Z(n9008) );
  XNOR U13327 ( .A(n12268), .B(n12020), .Z(n10845) );
  XOR U13328 ( .A(n12269), .B(n12270), .Z(n12020) );
  XNOR U13329 ( .A(round_reg[1539]), .B(round_reg[1219]), .Z(n12270) );
  XOR U13330 ( .A(round_reg[259]), .B(n12271), .Z(n12269) );
  XOR U13331 ( .A(round_reg[899]), .B(round_reg[579]), .Z(n12271) );
  XOR U13332 ( .A(n12272), .B(n6642), .Z(n9047) );
  XOR U13333 ( .A(round_reg[677]), .B(n10534), .Z(n6642) );
  IV U13334 ( .A(n9851), .Z(n10534) );
  XNOR U13335 ( .A(n11604), .B(n11966), .Z(n9851) );
  XNOR U13336 ( .A(n12273), .B(n12274), .Z(n11966) );
  XNOR U13337 ( .A(round_reg[1061]), .B(round_reg[101]), .Z(n12274) );
  XOR U13338 ( .A(round_reg[1381]), .B(n12275), .Z(n12273) );
  XOR U13339 ( .A(round_reg[741]), .B(round_reg[421]), .Z(n12275) );
  XOR U13340 ( .A(n12276), .B(n12277), .Z(n11604) );
  XNOR U13341 ( .A(round_reg[1572]), .B(round_reg[1252]), .Z(n12277) );
  XOR U13342 ( .A(round_reg[292]), .B(n12278), .Z(n12276) );
  XOR U13343 ( .A(round_reg[932]), .B(round_reg[612]), .Z(n12278) );
  NOR U13344 ( .A(n9003), .B(n9004), .Z(n12272) );
  XOR U13345 ( .A(round_reg[202]), .B(n10710), .Z(n9004) );
  XNOR U13346 ( .A(round_reg[611]), .B(n9449), .Z(n9003) );
  IV U13347 ( .A(n11005), .Z(n9449) );
  XOR U13348 ( .A(n12279), .B(n12008), .Z(n11005) );
  XOR U13349 ( .A(n12280), .B(n12281), .Z(n12008) );
  XNOR U13350 ( .A(round_reg[1506]), .B(round_reg[1186]), .Z(n12281) );
  XOR U13351 ( .A(round_reg[226]), .B(n12282), .Z(n12280) );
  XOR U13352 ( .A(round_reg[866]), .B(round_reg[546]), .Z(n12282) );
  XNOR U13353 ( .A(n12283), .B(n6638), .Z(n3492) );
  XOR U13354 ( .A(round_reg[834]), .B(n9709), .Z(n6638) );
  IV U13355 ( .A(n9695), .Z(n9709) );
  XNOR U13356 ( .A(n11738), .B(n11899), .Z(n9695) );
  XNOR U13357 ( .A(n12284), .B(n12285), .Z(n11899) );
  XNOR U13358 ( .A(round_reg[129]), .B(round_reg[1089]), .Z(n12285) );
  XOR U13359 ( .A(round_reg[1409]), .B(n12286), .Z(n12284) );
  XOR U13360 ( .A(round_reg[769]), .B(round_reg[449]), .Z(n12286) );
  XOR U13361 ( .A(n12287), .B(n12288), .Z(n11738) );
  XNOR U13362 ( .A(round_reg[1538]), .B(round_reg[1218]), .Z(n12288) );
  XOR U13363 ( .A(round_reg[258]), .B(n12289), .Z(n12287) );
  XOR U13364 ( .A(round_reg[898]), .B(round_reg[578]), .Z(n12289) );
  ANDN U13365 ( .B(n9001), .A(n9000), .Z(n12283) );
  XNOR U13366 ( .A(round_reg[509]), .B(n9761), .Z(n9000) );
  IV U13367 ( .A(n9961), .Z(n9761) );
  XOR U13368 ( .A(n11711), .B(n12290), .Z(n9961) );
  XOR U13369 ( .A(n12291), .B(n12292), .Z(n11711) );
  XNOR U13370 ( .A(round_reg[124]), .B(round_reg[1084]), .Z(n12292) );
  XOR U13371 ( .A(round_reg[1404]), .B(n12293), .Z(n12291) );
  XOR U13372 ( .A(round_reg[764]), .B(round_reg[444]), .Z(n12293) );
  XOR U13373 ( .A(round_reg[84]), .B(n11313), .Z(n9001) );
  XNOR U13374 ( .A(n12294), .B(n12295), .Z(n6398) );
  XNOR U13375 ( .A(n3690), .B(n5493), .Z(n12295) );
  XNOR U13376 ( .A(n12296), .B(n9062), .Z(n5493) );
  XOR U13377 ( .A(round_reg[201]), .B(n9091), .Z(n9062) );
  AND U13378 ( .A(n6666), .B(n6668), .Z(n12296) );
  XOR U13379 ( .A(round_reg[1044]), .B(n11313), .Z(n6668) );
  XOR U13380 ( .A(n12297), .B(n12298), .Z(n11313) );
  XOR U13381 ( .A(round_reg[1421]), .B(n11194), .Z(n6666) );
  XNOR U13382 ( .A(n12299), .B(n7144), .Z(n3690) );
  XOR U13383 ( .A(round_reg[61]), .B(n11575), .Z(n7144) );
  IV U13384 ( .A(n9615), .Z(n11575) );
  XNOR U13385 ( .A(n10147), .B(n12026), .Z(n9615) );
  XNOR U13386 ( .A(n12300), .B(n12301), .Z(n12026) );
  XNOR U13387 ( .A(round_reg[125]), .B(round_reg[1085]), .Z(n12301) );
  XOR U13388 ( .A(round_reg[1405]), .B(n12302), .Z(n12300) );
  XOR U13389 ( .A(round_reg[765]), .B(round_reg[445]), .Z(n12302) );
  XOR U13390 ( .A(n12303), .B(n12304), .Z(n10147) );
  XNOR U13391 ( .A(round_reg[1596]), .B(round_reg[1276]), .Z(n12304) );
  XOR U13392 ( .A(round_reg[316]), .B(n12305), .Z(n12303) );
  XOR U13393 ( .A(round_reg[956]), .B(round_reg[636]), .Z(n12305) );
  AND U13394 ( .A(n6657), .B(n9107), .Z(n12299) );
  IV U13395 ( .A(n6659), .Z(n9107) );
  XNOR U13396 ( .A(round_reg[1183]), .B(n9894), .Z(n6659) );
  XNOR U13397 ( .A(n11516), .B(n11888), .Z(n9894) );
  XNOR U13398 ( .A(n12306), .B(n12307), .Z(n11888) );
  XNOR U13399 ( .A(round_reg[1438]), .B(round_reg[1118]), .Z(n12307) );
  XOR U13400 ( .A(round_reg[158]), .B(n12308), .Z(n12306) );
  XOR U13401 ( .A(round_reg[798]), .B(round_reg[478]), .Z(n12308) );
  XOR U13402 ( .A(n12309), .B(n12310), .Z(n11516) );
  XNOR U13403 ( .A(round_reg[1567]), .B(round_reg[1247]), .Z(n12310) );
  XOR U13404 ( .A(round_reg[287]), .B(n12311), .Z(n12309) );
  XOR U13405 ( .A(round_reg[927]), .B(round_reg[607]), .Z(n12311) );
  XOR U13406 ( .A(round_reg[1547]), .B(n11125), .Z(n6657) );
  IV U13407 ( .A(n11068), .Z(n11125) );
  XNOR U13408 ( .A(n11031), .B(n12312), .Z(n11068) );
  XOR U13409 ( .A(n12313), .B(n12314), .Z(n11031) );
  XNOR U13410 ( .A(round_reg[1291]), .B(round_reg[11]), .Z(n12314) );
  XOR U13411 ( .A(round_reg[331]), .B(n12315), .Z(n12313) );
  XOR U13412 ( .A(round_reg[971]), .B(round_reg[651]), .Z(n12315) );
  XOR U13413 ( .A(n4262), .B(n12316), .Z(n12294) );
  XNOR U13414 ( .A(n5967), .B(n2148), .Z(n12316) );
  XNOR U13415 ( .A(n12317), .B(n7136), .Z(n2148) );
  XOR U13416 ( .A(round_reg[83]), .B(n9183), .Z(n7136) );
  XNOR U13417 ( .A(n11862), .B(n12318), .Z(n9183) );
  XOR U13418 ( .A(n12319), .B(n12320), .Z(n11862) );
  XNOR U13419 ( .A(round_reg[18]), .B(round_reg[1298]), .Z(n12320) );
  XOR U13420 ( .A(round_reg[338]), .B(n12321), .Z(n12319) );
  XOR U13421 ( .A(round_reg[978]), .B(round_reg[658]), .Z(n12321) );
  AND U13422 ( .A(n6662), .B(n9111), .Z(n12317) );
  IV U13423 ( .A(n6664), .Z(n9111) );
  XNOR U13424 ( .A(round_reg[1255]), .B(n9818), .Z(n6664) );
  XOR U13425 ( .A(n12322), .B(n11965), .Z(n9818) );
  XOR U13426 ( .A(n12323), .B(n12324), .Z(n11965) );
  XNOR U13427 ( .A(round_reg[1510]), .B(round_reg[1190]), .Z(n12324) );
  XOR U13428 ( .A(round_reg[230]), .B(n12325), .Z(n12323) );
  XOR U13429 ( .A(round_reg[870]), .B(round_reg[550]), .Z(n12325) );
  XOR U13430 ( .A(round_reg[1328]), .B(n9675), .Z(n6662) );
  IV U13431 ( .A(n11562), .Z(n9675) );
  XNOR U13432 ( .A(n11318), .B(n11513), .Z(n11562) );
  XNOR U13433 ( .A(n12326), .B(n12327), .Z(n11513) );
  XNOR U13434 ( .A(round_reg[112]), .B(round_reg[1072]), .Z(n12327) );
  XOR U13435 ( .A(round_reg[1392]), .B(n12328), .Z(n12326) );
  XOR U13436 ( .A(round_reg[752]), .B(round_reg[432]), .Z(n12328) );
  XOR U13437 ( .A(n12329), .B(n12330), .Z(n11318) );
  XNOR U13438 ( .A(round_reg[1583]), .B(round_reg[1263]), .Z(n12330) );
  XOR U13439 ( .A(round_reg[303]), .B(n12331), .Z(n12329) );
  XOR U13440 ( .A(round_reg[943]), .B(round_reg[623]), .Z(n12331) );
  XOR U13441 ( .A(n12332), .B(n7141), .Z(n5967) );
  XOR U13442 ( .A(round_reg[142]), .B(n10529), .Z(n7141) );
  XOR U13443 ( .A(n11683), .B(n12116), .Z(n10529) );
  XNOR U13444 ( .A(n12333), .B(n12334), .Z(n12116) );
  XNOR U13445 ( .A(round_reg[1357]), .B(round_reg[1037]), .Z(n12334) );
  XOR U13446 ( .A(round_reg[397]), .B(n12335), .Z(n12333) );
  XOR U13447 ( .A(round_reg[77]), .B(round_reg[717]), .Z(n12335) );
  XOR U13448 ( .A(n12336), .B(n12337), .Z(n11683) );
  XNOR U13449 ( .A(round_reg[1486]), .B(round_reg[1166]), .Z(n12337) );
  XOR U13450 ( .A(round_reg[206]), .B(n12338), .Z(n12336) );
  XOR U13451 ( .A(round_reg[846]), .B(round_reg[526]), .Z(n12338) );
  ANDN U13452 ( .B(n6655), .A(n6653), .Z(n12332) );
  XNOR U13453 ( .A(round_reg[1391]), .B(n9375), .Z(n6653) );
  XOR U13454 ( .A(n11236), .B(n11713), .Z(n9375) );
  XNOR U13455 ( .A(n12339), .B(n12340), .Z(n11713) );
  XNOR U13456 ( .A(round_reg[1326]), .B(round_reg[1006]), .Z(n12340) );
  XOR U13457 ( .A(round_reg[366]), .B(n12341), .Z(n12339) );
  XOR U13458 ( .A(round_reg[686]), .B(round_reg[46]), .Z(n12341) );
  XOR U13459 ( .A(n12342), .B(n12343), .Z(n11236) );
  XNOR U13460 ( .A(round_reg[1455]), .B(round_reg[1135]), .Z(n12343) );
  XOR U13461 ( .A(round_reg[175]), .B(n12344), .Z(n12342) );
  XOR U13462 ( .A(round_reg[815]), .B(round_reg[495]), .Z(n12344) );
  XNOR U13463 ( .A(round_reg[1015]), .B(n9550), .Z(n6655) );
  XOR U13464 ( .A(n12345), .B(n11015), .Z(n9550) );
  XNOR U13465 ( .A(n12346), .B(n12347), .Z(n11015) );
  XNOR U13466 ( .A(round_reg[1590]), .B(round_reg[1270]), .Z(n12347) );
  XOR U13467 ( .A(round_reg[310]), .B(n12348), .Z(n12346) );
  XOR U13468 ( .A(round_reg[950]), .B(round_reg[630]), .Z(n12348) );
  XNOR U13469 ( .A(n12349), .B(n7133), .Z(n4262) );
  XOR U13470 ( .A(round_reg[313]), .B(n10290), .Z(n7133) );
  IV U13471 ( .A(n10923), .Z(n10290) );
  AND U13472 ( .A(n6670), .B(n9102), .Z(n12349) );
  IV U13473 ( .A(n6672), .Z(n9102) );
  XNOR U13474 ( .A(round_reg[1093]), .B(n9700), .Z(n6672) );
  XOR U13475 ( .A(round_reg[1482]), .B(n10710), .Z(n6670) );
  XOR U13476 ( .A(n11473), .B(n12352), .Z(n10710) );
  XOR U13477 ( .A(n12353), .B(n12354), .Z(n11473) );
  XNOR U13478 ( .A(round_reg[1546]), .B(round_reg[1226]), .Z(n12354) );
  XOR U13479 ( .A(round_reg[266]), .B(n12355), .Z(n12353) );
  XOR U13480 ( .A(round_reg[906]), .B(round_reg[586]), .Z(n12355) );
  XNOR U13481 ( .A(n12356), .B(n9054), .Z(n9006) );
  XOR U13482 ( .A(round_reg[439]), .B(n11409), .Z(n9054) );
  NOR U13483 ( .A(n12030), .B(n6631), .Z(n12356) );
  XNOR U13484 ( .A(round_reg[1548]), .B(n10887), .Z(n6631) );
  XNOR U13485 ( .A(n12357), .B(n10991), .Z(n10887) );
  XNOR U13486 ( .A(n12358), .B(n12359), .Z(n10991) );
  XNOR U13487 ( .A(round_reg[12]), .B(round_reg[1292]), .Z(n12359) );
  XOR U13488 ( .A(round_reg[332]), .B(n12360), .Z(n12358) );
  XOR U13489 ( .A(round_reg[972]), .B(round_reg[652]), .Z(n12360) );
  XOR U13490 ( .A(round_reg[62]), .B(n9536), .Z(n12030) );
  XOR U13491 ( .A(n12361), .B(n11831), .Z(n9536) );
  XOR U13492 ( .A(n12362), .B(n12363), .Z(n11831) );
  XNOR U13493 ( .A(round_reg[126]), .B(round_reg[1086]), .Z(n12363) );
  XOR U13494 ( .A(round_reg[1406]), .B(n12364), .Z(n12362) );
  XOR U13495 ( .A(round_reg[766]), .B(round_reg[446]), .Z(n12364) );
  XOR U13496 ( .A(n11091), .B(n2111), .Z(n5726) );
  XNOR U13497 ( .A(n8438), .B(n9713), .Z(n2111) );
  XNOR U13498 ( .A(n12365), .B(n12366), .Z(n9713) );
  XOR U13499 ( .A(n5530), .B(n3615), .Z(n12366) );
  XOR U13500 ( .A(n12367), .B(n8531), .Z(n3615) );
  XOR U13501 ( .A(round_reg[1399]), .B(n11409), .Z(n8531) );
  XOR U13502 ( .A(n12368), .B(n12369), .Z(n11409) );
  AND U13503 ( .A(n8583), .B(n8582), .Z(n12367) );
  XOR U13504 ( .A(round_reg[1023]), .B(n11341), .Z(n8582) );
  XNOR U13505 ( .A(n12371), .B(n12372), .Z(n12140) );
  XNOR U13506 ( .A(round_reg[1598]), .B(round_reg[1278]), .Z(n12372) );
  XOR U13507 ( .A(round_reg[318]), .B(n12373), .Z(n12371) );
  XOR U13508 ( .A(round_reg[958]), .B(round_reg[638]), .Z(n12373) );
  XNOR U13509 ( .A(round_reg[912]), .B(n10541), .Z(n8583) );
  IV U13510 ( .A(n10577), .Z(n10541) );
  XOR U13511 ( .A(n12374), .B(n12251), .Z(n10577) );
  XOR U13512 ( .A(n12375), .B(n12376), .Z(n12251) );
  XNOR U13513 ( .A(round_reg[1487]), .B(round_reg[1167]), .Z(n12376) );
  XOR U13514 ( .A(round_reg[207]), .B(n12377), .Z(n12375) );
  XOR U13515 ( .A(round_reg[847]), .B(round_reg[527]), .Z(n12377) );
  XNOR U13516 ( .A(n12378), .B(n11174), .Z(n5530) );
  XOR U13517 ( .A(round_reg[1555]), .B(n10707), .Z(n11174) );
  IV U13518 ( .A(n10317), .Z(n10707) );
  XNOR U13519 ( .A(n12298), .B(n12379), .Z(n10317) );
  XOR U13520 ( .A(n12380), .B(n12381), .Z(n12298) );
  XNOR U13521 ( .A(round_reg[19]), .B(round_reg[1299]), .Z(n12381) );
  XOR U13522 ( .A(round_reg[339]), .B(n12382), .Z(n12380) );
  XOR U13523 ( .A(round_reg[979]), .B(round_reg[659]), .Z(n12382) );
  ANDN U13524 ( .B(n8580), .A(n8578), .Z(n12378) );
  XNOR U13525 ( .A(round_reg[1191]), .B(n9984), .Z(n8578) );
  IV U13526 ( .A(n12383), .Z(n9984) );
  XOR U13527 ( .A(round_reg[808]), .B(n10981), .Z(n8580) );
  XNOR U13528 ( .A(n11935), .B(n11815), .Z(n10981) );
  XNOR U13529 ( .A(n12384), .B(n12385), .Z(n11815) );
  XNOR U13530 ( .A(round_reg[1063]), .B(round_reg[103]), .Z(n12385) );
  XOR U13531 ( .A(round_reg[1383]), .B(n12386), .Z(n12384) );
  XOR U13532 ( .A(round_reg[743]), .B(round_reg[423]), .Z(n12386) );
  XOR U13533 ( .A(n12387), .B(n12388), .Z(n11935) );
  XNOR U13534 ( .A(round_reg[1512]), .B(round_reg[1192]), .Z(n12388) );
  XOR U13535 ( .A(round_reg[232]), .B(n12389), .Z(n12387) );
  XOR U13536 ( .A(round_reg[872]), .B(round_reg[552]), .Z(n12389) );
  XOR U13537 ( .A(n6360), .B(n12390), .Z(n12365) );
  XOR U13538 ( .A(n2415), .B(n5741), .Z(n12390) );
  XNOR U13539 ( .A(n12391), .B(n8517), .Z(n5741) );
  XOR U13540 ( .A(round_reg[1336]), .B(n9466), .Z(n8517) );
  IV U13541 ( .A(n12046), .Z(n9466) );
  XOR U13542 ( .A(n10689), .B(n10539), .Z(n12046) );
  XOR U13543 ( .A(n12392), .B(n12393), .Z(n10539) );
  XNOR U13544 ( .A(round_reg[1591]), .B(round_reg[1271]), .Z(n12393) );
  XOR U13545 ( .A(round_reg[311]), .B(n12394), .Z(n12392) );
  XOR U13546 ( .A(round_reg[951]), .B(round_reg[631]), .Z(n12394) );
  XOR U13547 ( .A(n12395), .B(n12396), .Z(n10689) );
  XNOR U13548 ( .A(round_reg[120]), .B(round_reg[1080]), .Z(n12396) );
  XOR U13549 ( .A(round_reg[1400]), .B(n12397), .Z(n12395) );
  XOR U13550 ( .A(round_reg[760]), .B(round_reg[440]), .Z(n12397) );
  AND U13551 ( .A(n9716), .B(n9715), .Z(n12391) );
  XNOR U13552 ( .A(round_reg[1263]), .B(n11210), .Z(n9715) );
  XNOR U13553 ( .A(round_reg[841]), .B(n9091), .Z(n9716) );
  IV U13554 ( .A(n10800), .Z(n9091) );
  XNOR U13555 ( .A(n11581), .B(n11123), .Z(n10800) );
  XNOR U13556 ( .A(n12398), .B(n12399), .Z(n11123) );
  XNOR U13557 ( .A(round_reg[136]), .B(round_reg[1096]), .Z(n12399) );
  XOR U13558 ( .A(round_reg[1416]), .B(n12400), .Z(n12398) );
  XOR U13559 ( .A(round_reg[776]), .B(round_reg[456]), .Z(n12400) );
  XOR U13560 ( .A(n12401), .B(n12402), .Z(n11581) );
  XNOR U13561 ( .A(round_reg[1545]), .B(round_reg[1225]), .Z(n12402) );
  XOR U13562 ( .A(round_reg[265]), .B(n12403), .Z(n12401) );
  XOR U13563 ( .A(round_reg[905]), .B(round_reg[585]), .Z(n12403) );
  XNOR U13564 ( .A(n12404), .B(n8521), .Z(n2415) );
  XOR U13565 ( .A(round_reg[1429]), .B(n9910), .Z(n8521) );
  XNOR U13566 ( .A(n11907), .B(n11410), .Z(n9910) );
  XOR U13567 ( .A(n12405), .B(n12406), .Z(n11410) );
  XNOR U13568 ( .A(round_reg[1364]), .B(round_reg[1044]), .Z(n12406) );
  XOR U13569 ( .A(round_reg[404]), .B(n12407), .Z(n12405) );
  XOR U13570 ( .A(round_reg[84]), .B(round_reg[724]), .Z(n12407) );
  XOR U13571 ( .A(n12408), .B(n12409), .Z(n11907) );
  XNOR U13572 ( .A(round_reg[1493]), .B(round_reg[1173]), .Z(n12409) );
  XOR U13573 ( .A(round_reg[213]), .B(n12410), .Z(n12408) );
  XOR U13574 ( .A(round_reg[853]), .B(round_reg[533]), .Z(n12410) );
  AND U13575 ( .A(n8569), .B(n11247), .Z(n12404) );
  XOR U13576 ( .A(round_reg[684]), .B(n9379), .Z(n11247) );
  XOR U13577 ( .A(n12201), .B(n11794), .Z(n9379) );
  XOR U13578 ( .A(n12411), .B(n12412), .Z(n11794) );
  XNOR U13579 ( .A(round_reg[1579]), .B(round_reg[1259]), .Z(n12412) );
  XOR U13580 ( .A(round_reg[299]), .B(n12413), .Z(n12411) );
  XOR U13581 ( .A(round_reg[939]), .B(round_reg[619]), .Z(n12413) );
  XOR U13582 ( .A(n12414), .B(n12415), .Z(n12201) );
  XNOR U13583 ( .A(round_reg[108]), .B(round_reg[1068]), .Z(n12415) );
  XOR U13584 ( .A(round_reg[1388]), .B(n12416), .Z(n12414) );
  XOR U13585 ( .A(round_reg[748]), .B(round_reg[428]), .Z(n12416) );
  XOR U13586 ( .A(round_reg[1052]), .B(n10872), .Z(n8569) );
  XNOR U13587 ( .A(n12417), .B(n8527), .Z(n6360) );
  XOR U13588 ( .A(round_reg[1490]), .B(n11107), .Z(n8527) );
  NOR U13589 ( .A(n8573), .B(n8574), .Z(n12417) );
  XNOR U13590 ( .A(round_reg[762]), .B(n11920), .Z(n8574) );
  XNOR U13591 ( .A(n12350), .B(n12418), .Z(n11920) );
  XOR U13592 ( .A(n12419), .B(n12420), .Z(n12350) );
  XNOR U13593 ( .A(round_reg[1337]), .B(round_reg[1017]), .Z(n12420) );
  XOR U13594 ( .A(round_reg[377]), .B(n12421), .Z(n12419) );
  XOR U13595 ( .A(round_reg[697]), .B(round_reg[57]), .Z(n12421) );
  XNOR U13596 ( .A(round_reg[1101]), .B(n11194), .Z(n8573) );
  IV U13597 ( .A(n9095), .Z(n11194) );
  XOR U13598 ( .A(n11856), .B(n12422), .Z(n9095) );
  XOR U13599 ( .A(n12423), .B(n12424), .Z(n11856) );
  XNOR U13600 ( .A(round_reg[1485]), .B(round_reg[1165]), .Z(n12424) );
  XOR U13601 ( .A(round_reg[205]), .B(n12425), .Z(n12423) );
  XOR U13602 ( .A(round_reg[845]), .B(round_reg[525]), .Z(n12425) );
  XOR U13603 ( .A(n12426), .B(n12427), .Z(n8438) );
  XNOR U13604 ( .A(n3800), .B(n5151), .Z(n12427) );
  XOR U13605 ( .A(n12428), .B(n9643), .Z(n5151) );
  XOR U13606 ( .A(round_reg[453]), .B(n9700), .Z(n9643) );
  XOR U13607 ( .A(n12268), .B(n12429), .Z(n9700) );
  XOR U13608 ( .A(n12430), .B(n12431), .Z(n12268) );
  XNOR U13609 ( .A(round_reg[1348]), .B(round_reg[1028]), .Z(n12431) );
  XOR U13610 ( .A(round_reg[388]), .B(n12432), .Z(n12430) );
  XOR U13611 ( .A(round_reg[708]), .B(round_reg[68]), .Z(n12432) );
  AND U13612 ( .A(n11098), .B(n11097), .Z(n12428) );
  XNOR U13613 ( .A(round_reg[92]), .B(n10509), .Z(n11097) );
  IV U13614 ( .A(n10872), .Z(n10509) );
  XOR U13615 ( .A(n10942), .B(n11616), .Z(n10872) );
  XNOR U13616 ( .A(n12433), .B(n12434), .Z(n11616) );
  XNOR U13617 ( .A(round_reg[27]), .B(round_reg[1307]), .Z(n12434) );
  XOR U13618 ( .A(round_reg[347]), .B(n12435), .Z(n12433) );
  XOR U13619 ( .A(round_reg[987]), .B(round_reg[667]), .Z(n12435) );
  XOR U13620 ( .A(n12436), .B(n12437), .Z(n10942) );
  XNOR U13621 ( .A(round_reg[1436]), .B(round_reg[1116]), .Z(n12437) );
  XOR U13622 ( .A(round_reg[156]), .B(n12438), .Z(n12436) );
  XOR U13623 ( .A(round_reg[796]), .B(round_reg[476]), .Z(n12438) );
  XNOR U13624 ( .A(round_reg[1337]), .B(n9389), .Z(n11098) );
  XNOR U13625 ( .A(n12439), .B(n8496), .Z(n3800) );
  XNOR U13626 ( .A(round_reg[619]), .B(n11543), .Z(n8496) );
  ANDN U13627 ( .B(n11090), .A(n11089), .Z(n12439) );
  XNOR U13628 ( .A(round_reg[210]), .B(n11107), .Z(n11089) );
  XNOR U13629 ( .A(round_reg[1430]), .B(n9841), .Z(n11090) );
  IV U13630 ( .A(n11245), .Z(n9841) );
  XOR U13631 ( .A(n11723), .B(n11309), .Z(n11245) );
  XOR U13632 ( .A(n12440), .B(n12441), .Z(n11309) );
  XNOR U13633 ( .A(round_reg[1365]), .B(round_reg[1045]), .Z(n12441) );
  XOR U13634 ( .A(round_reg[405]), .B(n12442), .Z(n12440) );
  XOR U13635 ( .A(round_reg[85]), .B(round_reg[725]), .Z(n12442) );
  XOR U13636 ( .A(n12443), .B(n12444), .Z(n11723) );
  XNOR U13637 ( .A(round_reg[1494]), .B(round_reg[1174]), .Z(n12444) );
  XOR U13638 ( .A(round_reg[214]), .B(n12445), .Z(n12443) );
  XOR U13639 ( .A(round_reg[854]), .B(round_reg[534]), .Z(n12445) );
  XOR U13640 ( .A(n5896), .B(n12446), .Z(n12426) );
  XOR U13641 ( .A(n1751), .B(n11159), .Z(n12446) );
  XOR U13642 ( .A(n12447), .B(n8506), .Z(n11159) );
  XNOR U13643 ( .A(round_reg[447]), .B(n10611), .Z(n8506) );
  IV U13644 ( .A(n11460), .Z(n10611) );
  XNOR U13645 ( .A(n12448), .B(n12449), .Z(n11460) );
  AND U13646 ( .A(n11086), .B(n12064), .Z(n12447) );
  IV U13647 ( .A(n11087), .Z(n12064) );
  XOR U13648 ( .A(round_reg[1556]), .B(n10622), .Z(n11087) );
  IV U13649 ( .A(n11169), .Z(n11086) );
  XNOR U13650 ( .A(round_reg[6]), .B(n10674), .Z(n11169) );
  XOR U13651 ( .A(n12450), .B(n12451), .Z(n11662) );
  XNOR U13652 ( .A(round_reg[1541]), .B(round_reg[1221]), .Z(n12451) );
  XOR U13653 ( .A(round_reg[261]), .B(n12452), .Z(n12450) );
  XOR U13654 ( .A(round_reg[901]), .B(round_reg[581]), .Z(n12452) );
  XNOR U13655 ( .A(n12453), .B(n12454), .Z(n11887) );
  XNOR U13656 ( .A(round_reg[1350]), .B(round_reg[1030]), .Z(n12454) );
  XOR U13657 ( .A(round_reg[390]), .B(n12455), .Z(n12453) );
  XOR U13658 ( .A(round_reg[710]), .B(round_reg[70]), .Z(n12455) );
  XOR U13659 ( .A(n12456), .B(n8500), .Z(n1751) );
  XNOR U13660 ( .A(round_reg[332]), .B(n10168), .Z(n8500) );
  IV U13661 ( .A(n10771), .Z(n10168) );
  XOR U13662 ( .A(n12422), .B(n12048), .Z(n10771) );
  XOR U13663 ( .A(n12457), .B(n12458), .Z(n12048) );
  XNOR U13664 ( .A(round_reg[1547]), .B(round_reg[1227]), .Z(n12458) );
  XOR U13665 ( .A(round_reg[267]), .B(n12459), .Z(n12457) );
  XOR U13666 ( .A(round_reg[907]), .B(round_reg[587]), .Z(n12459) );
  XOR U13667 ( .A(n12460), .B(n12461), .Z(n12422) );
  XNOR U13668 ( .A(round_reg[1356]), .B(round_reg[1036]), .Z(n12461) );
  XOR U13669 ( .A(round_reg[396]), .B(n12462), .Z(n12460) );
  XOR U13670 ( .A(round_reg[76]), .B(round_reg[716]), .Z(n12462) );
  ANDN U13671 ( .B(n12079), .A(n11094), .Z(n12456) );
  XOR U13672 ( .A(round_reg[258]), .B(n10999), .Z(n11094) );
  XNOR U13673 ( .A(n11941), .B(n11580), .Z(n10999) );
  XNOR U13674 ( .A(n12463), .B(n12464), .Z(n11580) );
  XNOR U13675 ( .A(round_reg[2]), .B(round_reg[1282]), .Z(n12464) );
  XOR U13676 ( .A(round_reg[322]), .B(n12465), .Z(n12463) );
  XOR U13677 ( .A(round_reg[962]), .B(round_reg[642]), .Z(n12465) );
  XOR U13678 ( .A(n12466), .B(n12467), .Z(n11941) );
  XNOR U13679 ( .A(round_reg[1473]), .B(round_reg[1153]), .Z(n12467) );
  XOR U13680 ( .A(round_reg[193]), .B(n12468), .Z(n12466) );
  XOR U13681 ( .A(round_reg[833]), .B(round_reg[513]), .Z(n12468) );
  IV U13682 ( .A(n11095), .Z(n12079) );
  XOR U13683 ( .A(round_reg[1491]), .B(n9996), .Z(n11095) );
  IV U13684 ( .A(n9907), .Z(n9996) );
  XNOR U13685 ( .A(n12175), .B(n11411), .Z(n9907) );
  XNOR U13686 ( .A(n12469), .B(n12470), .Z(n11411) );
  XNOR U13687 ( .A(round_reg[1555]), .B(round_reg[1235]), .Z(n12470) );
  XOR U13688 ( .A(round_reg[275]), .B(n12471), .Z(n12469) );
  XOR U13689 ( .A(round_reg[915]), .B(round_reg[595]), .Z(n12471) );
  XOR U13690 ( .A(n12472), .B(n12473), .Z(n12175) );
  XNOR U13691 ( .A(round_reg[1426]), .B(round_reg[1106]), .Z(n12473) );
  XOR U13692 ( .A(round_reg[146]), .B(n12474), .Z(n12472) );
  XOR U13693 ( .A(round_reg[786]), .B(round_reg[466]), .Z(n12474) );
  XNOR U13694 ( .A(n12475), .B(n8510), .Z(n5896) );
  XNOR U13695 ( .A(round_reg[551]), .B(n12383), .Z(n8510) );
  XOR U13696 ( .A(n10932), .B(n11655), .Z(n12383) );
  XOR U13697 ( .A(n12476), .B(n12477), .Z(n11655) );
  XNOR U13698 ( .A(round_reg[1575]), .B(round_reg[1255]), .Z(n12477) );
  XOR U13699 ( .A(round_reg[295]), .B(n12478), .Z(n12476) );
  XOR U13700 ( .A(round_reg[935]), .B(round_reg[615]), .Z(n12478) );
  XOR U13701 ( .A(n12479), .B(n12480), .Z(n10932) );
  XNOR U13702 ( .A(round_reg[1446]), .B(round_reg[1126]), .Z(n12480) );
  XOR U13703 ( .A(round_reg[166]), .B(n12481), .Z(n12479) );
  XOR U13704 ( .A(round_reg[806]), .B(round_reg[486]), .Z(n12481) );
  NOR U13705 ( .A(n11166), .B(n12058), .Z(n12475) );
  XNOR U13706 ( .A(n12482), .B(n11166), .Z(n11091) );
  XNOR U13707 ( .A(round_reg[151]), .B(n11000), .Z(n11166) );
  AND U13708 ( .A(n8509), .B(n12058), .Z(n12482) );
  XOR U13709 ( .A(round_reg[1400]), .B(n11308), .Z(n12058) );
  XOR U13710 ( .A(n11003), .B(n12483), .Z(n11308) );
  XOR U13711 ( .A(n12484), .B(n12485), .Z(n11003) );
  XNOR U13712 ( .A(round_reg[1464]), .B(round_reg[1144]), .Z(n12485) );
  XOR U13713 ( .A(round_reg[184]), .B(n12486), .Z(n12484) );
  XOR U13714 ( .A(round_reg[824]), .B(round_reg[504]), .Z(n12486) );
  XNOR U13715 ( .A(round_reg[960]), .B(n11275), .Z(n8509) );
  XOR U13716 ( .A(n11940), .B(n12487), .Z(n11275) );
  XOR U13717 ( .A(n12488), .B(n12489), .Z(n11940) );
  XNOR U13718 ( .A(round_reg[1344]), .B(round_reg[1024]), .Z(n12489) );
  XOR U13719 ( .A(round_reg[384]), .B(n12490), .Z(n12488) );
  XOR U13720 ( .A(round_reg[704]), .B(round_reg[64]), .Z(n12490) );
  XOR U13721 ( .A(n12491), .B(n2622), .Z(out[0]) );
  XNOR U13722 ( .A(n2222), .B(n10122), .Z(n2622) );
  XOR U13723 ( .A(n12492), .B(n8618), .Z(n10122) );
  ANDN U13724 ( .B(n10146), .A(n10018), .Z(n12492) );
  XNOR U13725 ( .A(round_reg[597]), .B(n10164), .Z(n10018) );
  XOR U13726 ( .A(n11427), .B(n12146), .Z(n10164) );
  XOR U13727 ( .A(n12493), .B(n12494), .Z(n12146) );
  XNOR U13728 ( .A(round_reg[21]), .B(round_reg[1301]), .Z(n12494) );
  XOR U13729 ( .A(round_reg[341]), .B(n12495), .Z(n12493) );
  XOR U13730 ( .A(round_reg[981]), .B(round_reg[661]), .Z(n12495) );
  XOR U13731 ( .A(n12496), .B(n12497), .Z(n11427) );
  XNOR U13732 ( .A(round_reg[1492]), .B(round_reg[1172]), .Z(n12497) );
  XOR U13733 ( .A(round_reg[212]), .B(n12498), .Z(n12496) );
  XOR U13734 ( .A(round_reg[852]), .B(round_reg[532]), .Z(n12498) );
  XOR U13735 ( .A(n8045), .B(n6035), .Z(n2222) );
  XNOR U13736 ( .A(n12499), .B(n12500), .Z(n6035) );
  XNOR U13737 ( .A(n5300), .B(n3706), .Z(n12500) );
  XOR U13738 ( .A(n12501), .B(n8621), .Z(n3706) );
  XNOR U13739 ( .A(round_reg[1378]), .B(n10369), .Z(n8621) );
  XNOR U13740 ( .A(n11056), .B(n11762), .Z(n10369) );
  XNOR U13741 ( .A(n12502), .B(n12503), .Z(n11762) );
  XNOR U13742 ( .A(round_reg[1442]), .B(round_reg[1122]), .Z(n12503) );
  XOR U13743 ( .A(round_reg[162]), .B(n12504), .Z(n12502) );
  XOR U13744 ( .A(round_reg[802]), .B(round_reg[482]), .Z(n12504) );
  XOR U13745 ( .A(n12505), .B(n12506), .Z(n11056) );
  XNOR U13746 ( .A(round_reg[33]), .B(round_reg[1313]), .Z(n12506) );
  XOR U13747 ( .A(round_reg[353]), .B(n12507), .Z(n12505) );
  XOR U13748 ( .A(round_reg[993]), .B(round_reg[673]), .Z(n12507) );
  AND U13749 ( .A(n7955), .B(n8622), .Z(n12501) );
  XOR U13750 ( .A(round_reg[1002]), .B(n10515), .Z(n8622) );
  IV U13751 ( .A(n9540), .Z(n10515) );
  XNOR U13752 ( .A(n11689), .B(n12241), .Z(n9540) );
  XNOR U13753 ( .A(n12508), .B(n12509), .Z(n12241) );
  XNOR U13754 ( .A(round_reg[1577]), .B(round_reg[1257]), .Z(n12509) );
  XOR U13755 ( .A(round_reg[297]), .B(n12510), .Z(n12508) );
  XOR U13756 ( .A(round_reg[937]), .B(round_reg[617]), .Z(n12510) );
  XOR U13757 ( .A(n12511), .B(n12512), .Z(n11689) );
  XNOR U13758 ( .A(round_reg[106]), .B(round_reg[1066]), .Z(n12512) );
  XOR U13759 ( .A(round_reg[1386]), .B(n12513), .Z(n12511) );
  XOR U13760 ( .A(round_reg[746]), .B(round_reg[426]), .Z(n12513) );
  XOR U13761 ( .A(round_reg[955]), .B(n10440), .Z(n7955) );
  XNOR U13762 ( .A(n12514), .B(n11881), .Z(n10440) );
  XNOR U13763 ( .A(n12515), .B(n12516), .Z(n11881) );
  XNOR U13764 ( .A(round_reg[1339]), .B(round_reg[1019]), .Z(n12516) );
  XOR U13765 ( .A(round_reg[379]), .B(n12517), .Z(n12515) );
  XOR U13766 ( .A(round_reg[699]), .B(round_reg[59]), .Z(n12517) );
  XNOR U13767 ( .A(n12518), .B(n8614), .Z(n5300) );
  XNOR U13768 ( .A(round_reg[1598]), .B(n9838), .Z(n8614) );
  IV U13769 ( .A(n11530), .Z(n9838) );
  XNOR U13770 ( .A(n12290), .B(n12449), .Z(n11530) );
  XNOR U13771 ( .A(n12519), .B(n12520), .Z(n12449) );
  XNOR U13772 ( .A(round_reg[1342]), .B(round_reg[1022]), .Z(n12520) );
  XOR U13773 ( .A(round_reg[382]), .B(n12521), .Z(n12519) );
  XOR U13774 ( .A(round_reg[702]), .B(round_reg[62]), .Z(n12521) );
  XOR U13775 ( .A(n12522), .B(n12523), .Z(n12290) );
  XNOR U13776 ( .A(round_reg[1533]), .B(round_reg[1213]), .Z(n12523) );
  XOR U13777 ( .A(round_reg[253]), .B(n12524), .Z(n12522) );
  XOR U13778 ( .A(round_reg[893]), .B(round_reg[573]), .Z(n12524) );
  AND U13779 ( .A(n7947), .B(n8615), .Z(n12518) );
  XOR U13780 ( .A(round_reg[1170]), .B(n11107), .Z(n8615) );
  XNOR U13781 ( .A(n12525), .B(n12526), .Z(n11506) );
  XNOR U13782 ( .A(round_reg[1554]), .B(round_reg[1234]), .Z(n12526) );
  XOR U13783 ( .A(round_reg[274]), .B(n12527), .Z(n12525) );
  XOR U13784 ( .A(round_reg[914]), .B(round_reg[594]), .Z(n12527) );
  XOR U13785 ( .A(round_reg[787]), .B(n10579), .Z(n7947) );
  XOR U13786 ( .A(n12529), .B(n11618), .Z(n10579) );
  XOR U13787 ( .A(n12530), .B(n12531), .Z(n11618) );
  XNOR U13788 ( .A(round_reg[1362]), .B(round_reg[1042]), .Z(n12531) );
  XOR U13789 ( .A(round_reg[402]), .B(n12532), .Z(n12530) );
  XOR U13790 ( .A(round_reg[82]), .B(round_reg[722]), .Z(n12532) );
  XNOR U13791 ( .A(n6454), .B(n12533), .Z(n12499) );
  XOR U13792 ( .A(n2570), .B(n8601), .Z(n12533) );
  XOR U13793 ( .A(n12534), .B(n8606), .Z(n8601) );
  XNOR U13794 ( .A(round_reg[1315]), .B(n11230), .Z(n8606) );
  IV U13795 ( .A(n9218), .Z(n11230) );
  XOR U13796 ( .A(n11951), .B(n11647), .Z(n9218) );
  XNOR U13797 ( .A(n12535), .B(n12536), .Z(n11647) );
  XNOR U13798 ( .A(round_reg[1379]), .B(round_reg[1059]), .Z(n12536) );
  XOR U13799 ( .A(round_reg[419]), .B(n12537), .Z(n12535) );
  XOR U13800 ( .A(round_reg[99]), .B(round_reg[739]), .Z(n12537) );
  XOR U13801 ( .A(n12538), .B(n12539), .Z(n11951) );
  XNOR U13802 ( .A(round_reg[1570]), .B(round_reg[1250]), .Z(n12539) );
  XOR U13803 ( .A(round_reg[290]), .B(n12540), .Z(n12538) );
  XOR U13804 ( .A(round_reg[930]), .B(round_reg[610]), .Z(n12540) );
  ANDN U13805 ( .B(n8607), .A(n7951), .Z(n12534) );
  XOR U13806 ( .A(round_reg[884]), .B(n10781), .Z(n7951) );
  XOR U13807 ( .A(n12264), .B(n12541), .Z(n10781) );
  XOR U13808 ( .A(n12542), .B(n12543), .Z(n12264) );
  XNOR U13809 ( .A(round_reg[1459]), .B(round_reg[1139]), .Z(n12543) );
  XOR U13810 ( .A(round_reg[179]), .B(n12544), .Z(n12542) );
  XOR U13811 ( .A(round_reg[819]), .B(round_reg[499]), .Z(n12544) );
  XOR U13812 ( .A(round_reg[1242]), .B(n11346), .Z(n8607) );
  IV U13813 ( .A(n9780), .Z(n11346) );
  XNOR U13814 ( .A(n11394), .B(n11919), .Z(n9780) );
  XNOR U13815 ( .A(n12545), .B(n12546), .Z(n11919) );
  XNOR U13816 ( .A(round_reg[1497]), .B(round_reg[1177]), .Z(n12546) );
  XOR U13817 ( .A(round_reg[217]), .B(n12547), .Z(n12545) );
  XOR U13818 ( .A(round_reg[857]), .B(round_reg[537]), .Z(n12547) );
  XOR U13819 ( .A(n12548), .B(n12549), .Z(n11394) );
  XNOR U13820 ( .A(round_reg[26]), .B(round_reg[1306]), .Z(n12549) );
  XOR U13821 ( .A(round_reg[346]), .B(n12550), .Z(n12548) );
  XOR U13822 ( .A(round_reg[986]), .B(round_reg[666]), .Z(n12550) );
  XOR U13823 ( .A(n12551), .B(n8619), .Z(n2570) );
  XNOR U13824 ( .A(round_reg[1408]), .B(n12552), .Z(n8619) );
  NOR U13825 ( .A(n10146), .B(n8618), .Z(n12551) );
  XNOR U13826 ( .A(round_reg[1031]), .B(n9925), .Z(n8618) );
  XOR U13827 ( .A(n11385), .B(n12553), .Z(n9925) );
  XOR U13828 ( .A(n12554), .B(n12555), .Z(n11385) );
  XNOR U13829 ( .A(round_reg[135]), .B(round_reg[1095]), .Z(n12555) );
  XOR U13830 ( .A(round_reg[1415]), .B(n12556), .Z(n12554) );
  XOR U13831 ( .A(round_reg[775]), .B(round_reg[455]), .Z(n12556) );
  XOR U13832 ( .A(round_reg[663]), .B(n10977), .Z(n10146) );
  IV U13833 ( .A(n10854), .Z(n10977) );
  XOR U13834 ( .A(n12557), .B(n12124), .Z(n10854) );
  XOR U13835 ( .A(n12558), .B(n12559), .Z(n12124) );
  XNOR U13836 ( .A(round_reg[1367]), .B(round_reg[1047]), .Z(n12559) );
  XOR U13837 ( .A(round_reg[407]), .B(n12560), .Z(n12558) );
  XOR U13838 ( .A(round_reg[87]), .B(round_reg[727]), .Z(n12560) );
  XNOR U13839 ( .A(n12561), .B(n8611), .Z(n6454) );
  XNOR U13840 ( .A(round_reg[1533]), .B(n9451), .Z(n8611) );
  XNOR U13841 ( .A(n11880), .B(n12361), .Z(n9451) );
  XOR U13842 ( .A(n12562), .B(n12563), .Z(n12361) );
  XNOR U13843 ( .A(round_reg[1597]), .B(round_reg[1277]), .Z(n12563) );
  XOR U13844 ( .A(round_reg[317]), .B(n12564), .Z(n12562) );
  XOR U13845 ( .A(round_reg[957]), .B(round_reg[637]), .Z(n12564) );
  XOR U13846 ( .A(n12565), .B(n12566), .Z(n11880) );
  XNOR U13847 ( .A(round_reg[1468]), .B(round_reg[1148]), .Z(n12566) );
  XOR U13848 ( .A(round_reg[188]), .B(n12567), .Z(n12565) );
  XOR U13849 ( .A(round_reg[828]), .B(round_reg[508]), .Z(n12567) );
  ANDN U13850 ( .B(n8610), .A(n7942), .Z(n12561) );
  XOR U13851 ( .A(round_reg[741]), .B(n11113), .Z(n7942) );
  XOR U13852 ( .A(round_reg[1144]), .B(n10422), .Z(n8610) );
  XOR U13853 ( .A(n12345), .B(n12351), .Z(n10422) );
  XNOR U13854 ( .A(n12568), .B(n12569), .Z(n12351) );
  XNOR U13855 ( .A(round_reg[1528]), .B(round_reg[1208]), .Z(n12569) );
  XOR U13856 ( .A(round_reg[248]), .B(n12570), .Z(n12568) );
  XOR U13857 ( .A(round_reg[888]), .B(round_reg[568]), .Z(n12570) );
  XOR U13858 ( .A(n12571), .B(n12572), .Z(n12345) );
  XNOR U13859 ( .A(round_reg[119]), .B(round_reg[1079]), .Z(n12572) );
  XOR U13860 ( .A(round_reg[1399]), .B(n12573), .Z(n12571) );
  XOR U13861 ( .A(round_reg[759]), .B(round_reg[439]), .Z(n12573) );
  XOR U13862 ( .A(n12574), .B(n12575), .Z(n8045) );
  XNOR U13863 ( .A(n4910), .B(n10203), .Z(n12575) );
  XOR U13864 ( .A(n12576), .B(n7037), .Z(n10203) );
  XNOR U13865 ( .A(round_reg[662]), .B(n9901), .Z(n7037) );
  XOR U13866 ( .A(round_reg[596]), .B(n10273), .Z(n10144) );
  IV U13867 ( .A(n10622), .Z(n10273) );
  XOR U13868 ( .A(n12529), .B(n12213), .Z(n10622) );
  XNOR U13869 ( .A(n12579), .B(n12580), .Z(n12213) );
  XNOR U13870 ( .A(round_reg[20]), .B(round_reg[1300]), .Z(n12580) );
  XOR U13871 ( .A(round_reg[340]), .B(n12581), .Z(n12579) );
  XOR U13872 ( .A(round_reg[980]), .B(round_reg[660]), .Z(n12581) );
  XOR U13873 ( .A(n12582), .B(n12583), .Z(n12529) );
  XNOR U13874 ( .A(round_reg[1491]), .B(round_reg[1171]), .Z(n12583) );
  XOR U13875 ( .A(round_reg[211]), .B(n12584), .Z(n12582) );
  XOR U13876 ( .A(round_reg[851]), .B(round_reg[531]), .Z(n12584) );
  XNOR U13877 ( .A(round_reg[251]), .B(n9611), .Z(n9291) );
  XOR U13878 ( .A(n11710), .B(n12418), .Z(n9611) );
  XNOR U13879 ( .A(n12585), .B(n12586), .Z(n12418) );
  XNOR U13880 ( .A(round_reg[1466]), .B(round_reg[1146]), .Z(n12586) );
  XOR U13881 ( .A(round_reg[186]), .B(n12587), .Z(n12585) );
  XOR U13882 ( .A(round_reg[826]), .B(round_reg[506]), .Z(n12587) );
  XOR U13883 ( .A(n12588), .B(n12589), .Z(n11710) );
  XNOR U13884 ( .A(round_reg[1595]), .B(round_reg[1275]), .Z(n12589) );
  XOR U13885 ( .A(round_reg[315]), .B(n12590), .Z(n12588) );
  XOR U13886 ( .A(round_reg[955]), .B(round_reg[635]), .Z(n12590) );
  XNOR U13887 ( .A(n12591), .B(n7042), .Z(n4910) );
  XOR U13888 ( .A(round_reg[740]), .B(n10528), .Z(n7042) );
  XOR U13889 ( .A(n12279), .B(n11491), .Z(n10528) );
  XNOR U13890 ( .A(n12592), .B(n12593), .Z(n11491) );
  XNOR U13891 ( .A(round_reg[1444]), .B(round_reg[1124]), .Z(n12593) );
  XOR U13892 ( .A(round_reg[164]), .B(n12594), .Z(n12592) );
  XOR U13893 ( .A(round_reg[804]), .B(round_reg[484]), .Z(n12594) );
  XOR U13894 ( .A(n12595), .B(n12596), .Z(n12279) );
  XNOR U13895 ( .A(round_reg[355]), .B(round_reg[1315]), .Z(n12596) );
  XOR U13896 ( .A(round_reg[35]), .B(n12597), .Z(n12595) );
  XOR U13897 ( .A(round_reg[995]), .B(round_reg[675]), .Z(n12597) );
  NOR U13898 ( .A(n10212), .B(n9286), .Z(n12591) );
  XNOR U13899 ( .A(round_reg[299]), .B(n11543), .Z(n9286) );
  IV U13900 ( .A(n11596), .Z(n11543) );
  XOR U13901 ( .A(n11868), .B(n12598), .Z(n11596) );
  XOR U13902 ( .A(n12599), .B(n12600), .Z(n11868) );
  XNOR U13903 ( .A(round_reg[1514]), .B(round_reg[1194]), .Z(n12600) );
  XOR U13904 ( .A(round_reg[234]), .B(n12601), .Z(n12599) );
  XOR U13905 ( .A(round_reg[874]), .B(round_reg[554]), .Z(n12601) );
  IV U13906 ( .A(n10133), .Z(n10212) );
  XOR U13907 ( .A(round_reg[373]), .B(n9257), .Z(n10133) );
  IV U13908 ( .A(n9703), .Z(n9257) );
  XNOR U13909 ( .A(n11061), .B(n12541), .Z(n9703) );
  XNOR U13910 ( .A(n12602), .B(n12603), .Z(n12541) );
  XNOR U13911 ( .A(round_reg[1588]), .B(round_reg[1268]), .Z(n12603) );
  XOR U13912 ( .A(round_reg[308]), .B(n12604), .Z(n12602) );
  XOR U13913 ( .A(round_reg[948]), .B(round_reg[628]), .Z(n12604) );
  XOR U13914 ( .A(n12605), .B(n12606), .Z(n11061) );
  XNOR U13915 ( .A(round_reg[117]), .B(round_reg[1077]), .Z(n12606) );
  XOR U13916 ( .A(round_reg[1397]), .B(n12607), .Z(n12605) );
  XOR U13917 ( .A(round_reg[757]), .B(round_reg[437]), .Z(n12607) );
  XOR U13918 ( .A(n2668), .B(n12608), .Z(n12574) );
  XOR U13919 ( .A(n3541), .B(n5776), .Z(n12608) );
  XOR U13920 ( .A(n12609), .B(n7031), .Z(n5776) );
  XNOR U13921 ( .A(round_reg[786]), .B(n11027), .Z(n7031) );
  IV U13922 ( .A(n11644), .Z(n11027) );
  XNOR U13923 ( .A(n11779), .B(n12379), .Z(n11644) );
  XNOR U13924 ( .A(n12610), .B(n12611), .Z(n12379) );
  XNOR U13925 ( .A(round_reg[1490]), .B(round_reg[1170]), .Z(n12611) );
  XOR U13926 ( .A(round_reg[210]), .B(n12612), .Z(n12610) );
  XOR U13927 ( .A(round_reg[850]), .B(round_reg[530]), .Z(n12612) );
  XOR U13928 ( .A(n12613), .B(n12614), .Z(n11779) );
  XNOR U13929 ( .A(round_reg[1361]), .B(round_reg[1041]), .Z(n12614) );
  XOR U13930 ( .A(round_reg[401]), .B(n12615), .Z(n12613) );
  XOR U13931 ( .A(round_reg[81]), .B(round_reg[721]), .Z(n12615) );
  NOR U13932 ( .A(n9289), .B(n10142), .Z(n12609) );
  XOR U13933 ( .A(round_reg[424]), .B(n9632), .Z(n10142) );
  XOR U13934 ( .A(n12322), .B(n12240), .Z(n9632) );
  XOR U13935 ( .A(n12616), .B(n12617), .Z(n12240) );
  XNOR U13936 ( .A(round_reg[1448]), .B(round_reg[1128]), .Z(n12617) );
  XOR U13937 ( .A(round_reg[168]), .B(n12618), .Z(n12616) );
  XOR U13938 ( .A(round_reg[808]), .B(round_reg[488]), .Z(n12618) );
  XOR U13939 ( .A(n12619), .B(n12620), .Z(n12322) );
  XNOR U13940 ( .A(round_reg[359]), .B(round_reg[1319]), .Z(n12620) );
  XOR U13941 ( .A(round_reg[39]), .B(n12621), .Z(n12619) );
  XOR U13942 ( .A(round_reg[999]), .B(round_reg[679]), .Z(n12621) );
  XNOR U13943 ( .A(round_reg[47]), .B(n11698), .Z(n9289) );
  XNOR U13944 ( .A(n11624), .B(n11423), .Z(n11698) );
  XNOR U13945 ( .A(n12622), .B(n12623), .Z(n11423) );
  XNOR U13946 ( .A(round_reg[1582]), .B(round_reg[1262]), .Z(n12623) );
  XOR U13947 ( .A(round_reg[302]), .B(n12624), .Z(n12622) );
  XOR U13948 ( .A(round_reg[942]), .B(round_reg[622]), .Z(n12624) );
  XOR U13949 ( .A(n12625), .B(n12626), .Z(n11624) );
  XNOR U13950 ( .A(round_reg[111]), .B(round_reg[1071]), .Z(n12626) );
  XOR U13951 ( .A(round_reg[1391]), .B(n12627), .Z(n12625) );
  XOR U13952 ( .A(round_reg[751]), .B(round_reg[431]), .Z(n12627) );
  XNOR U13953 ( .A(n12628), .B(n9295), .Z(n3541) );
  XNOR U13954 ( .A(round_reg[883]), .B(n10752), .Z(n9295) );
  XNOR U13955 ( .A(n12189), .B(n12629), .Z(n10752) );
  XOR U13956 ( .A(n12630), .B(n12631), .Z(n12189) );
  XNOR U13957 ( .A(round_reg[1458]), .B(round_reg[1138]), .Z(n12631) );
  XOR U13958 ( .A(round_reg[178]), .B(n12632), .Z(n12630) );
  XOR U13959 ( .A(round_reg[818]), .B(round_reg[498]), .Z(n12632) );
  ANDN U13960 ( .B(n10135), .A(n9282), .Z(n12628) );
  XOR U13961 ( .A(round_reg[69]), .B(n10293), .Z(n9282) );
  XOR U13962 ( .A(n11915), .B(n12633), .Z(n10293) );
  XOR U13963 ( .A(n12634), .B(n12635), .Z(n11915) );
  XNOR U13964 ( .A(round_reg[324]), .B(round_reg[1284]), .Z(n12635) );
  XOR U13965 ( .A(round_reg[4]), .B(n12636), .Z(n12634) );
  XOR U13966 ( .A(round_reg[964]), .B(round_reg[644]), .Z(n12636) );
  XNOR U13967 ( .A(round_reg[494]), .B(n11328), .Z(n10135) );
  IV U13968 ( .A(n11051), .Z(n11328) );
  XOR U13969 ( .A(n12637), .B(n12638), .Z(n11051) );
  XOR U13970 ( .A(n12639), .B(n7027), .Z(n2668) );
  XNOR U13971 ( .A(round_reg[954]), .B(n10384), .Z(n7027) );
  XNOR U13972 ( .A(n12640), .B(n12641), .Z(n12080) );
  XNOR U13973 ( .A(round_reg[1338]), .B(round_reg[1018]), .Z(n12641) );
  XOR U13974 ( .A(round_reg[378]), .B(n12642), .Z(n12640) );
  XOR U13975 ( .A(round_reg[698]), .B(round_reg[58]), .Z(n12642) );
  XNOR U13976 ( .A(n12643), .B(n12644), .Z(n10690) );
  XNOR U13977 ( .A(round_reg[1529]), .B(round_reg[1209]), .Z(n12644) );
  XOR U13978 ( .A(round_reg[249]), .B(n12645), .Z(n12643) );
  XOR U13979 ( .A(round_reg[889]), .B(round_reg[569]), .Z(n12645) );
  XOR U13980 ( .A(round_reg[528]), .B(n11368), .Z(n10139) );
  XOR U13981 ( .A(n11778), .B(n11983), .Z(n11368) );
  XOR U13982 ( .A(n12646), .B(n12647), .Z(n11983) );
  XNOR U13983 ( .A(round_reg[1423]), .B(round_reg[1103]), .Z(n12647) );
  XOR U13984 ( .A(round_reg[143]), .B(n12648), .Z(n12646) );
  XOR U13985 ( .A(round_reg[783]), .B(round_reg[463]), .Z(n12648) );
  XOR U13986 ( .A(n12649), .B(n12650), .Z(n11778) );
  XNOR U13987 ( .A(round_reg[1552]), .B(round_reg[1232]), .Z(n12650) );
  XOR U13988 ( .A(round_reg[272]), .B(n12651), .Z(n12649) );
  XOR U13989 ( .A(round_reg[912]), .B(round_reg[592]), .Z(n12651) );
  XNOR U13990 ( .A(round_reg[128]), .B(n9534), .Z(n9293) );
  IV U13991 ( .A(n12552), .Z(n9534) );
  XNOR U13992 ( .A(n12652), .B(n12370), .Z(n12552) );
  XNOR U13993 ( .A(n12653), .B(n12654), .Z(n12370) );
  XNOR U13994 ( .A(round_reg[127]), .B(round_reg[1087]), .Z(n12654) );
  XOR U13995 ( .A(round_reg[1407]), .B(n12655), .Z(n12653) );
  XOR U13996 ( .A(round_reg[767]), .B(round_reg[447]), .Z(n12655) );
  AND U13997 ( .A(n4043), .B(n4041), .Z(n12491) );
  XOR U13998 ( .A(n7675), .B(n2634), .Z(n4041) );
  XNOR U13999 ( .A(n6023), .B(n6450), .Z(n2634) );
  XNOR U14000 ( .A(n12656), .B(n12657), .Z(n6450) );
  XOR U14001 ( .A(n2670), .B(n5388), .Z(n12657) );
  XOR U14002 ( .A(n12658), .B(n6908), .Z(n5388) );
  XOR U14003 ( .A(round_reg[1006]), .B(n10791), .Z(n6908) );
  IV U14004 ( .A(n9205), .Z(n10791) );
  XNOR U14005 ( .A(n11782), .B(n11523), .Z(n9205) );
  XNOR U14006 ( .A(n12659), .B(n12660), .Z(n11523) );
  XNOR U14007 ( .A(round_reg[1581]), .B(round_reg[1261]), .Z(n12660) );
  XOR U14008 ( .A(round_reg[301]), .B(n12661), .Z(n12659) );
  XOR U14009 ( .A(round_reg[941]), .B(round_reg[621]), .Z(n12661) );
  XOR U14010 ( .A(n12662), .B(n12663), .Z(n11782) );
  XNOR U14011 ( .A(round_reg[110]), .B(round_reg[1070]), .Z(n12663) );
  XOR U14012 ( .A(round_reg[1390]), .B(n12664), .Z(n12662) );
  XOR U14013 ( .A(round_reg[750]), .B(round_reg[430]), .Z(n12664) );
  ANDN U14014 ( .B(n7683), .A(n6907), .Z(n12658) );
  XNOR U14015 ( .A(round_reg[959]), .B(n9930), .Z(n6907) );
  XNOR U14016 ( .A(n12025), .B(n12104), .Z(n9930) );
  XOR U14017 ( .A(n12665), .B(n12666), .Z(n12104) );
  XNOR U14018 ( .A(round_reg[1343]), .B(round_reg[1023]), .Z(n12666) );
  XOR U14019 ( .A(round_reg[383]), .B(n12667), .Z(n12665) );
  XOR U14020 ( .A(round_reg[703]), .B(round_reg[63]), .Z(n12667) );
  XOR U14021 ( .A(n12668), .B(n12669), .Z(n12025) );
  XNOR U14022 ( .A(round_reg[1534]), .B(round_reg[1214]), .Z(n12669) );
  XOR U14023 ( .A(round_reg[254]), .B(n12670), .Z(n12668) );
  XOR U14024 ( .A(round_reg[894]), .B(round_reg[574]), .Z(n12670) );
  XOR U14025 ( .A(round_reg[533]), .B(n10755), .Z(n7683) );
  IV U14026 ( .A(n9840), .Z(n10755) );
  XOR U14027 ( .A(n12297), .B(n12578), .Z(n9840) );
  XNOR U14028 ( .A(n12671), .B(n12672), .Z(n12578) );
  XNOR U14029 ( .A(round_reg[1557]), .B(round_reg[1237]), .Z(n12672) );
  XOR U14030 ( .A(round_reg[277]), .B(n12673), .Z(n12671) );
  XOR U14031 ( .A(round_reg[917]), .B(round_reg[597]), .Z(n12673) );
  XOR U14032 ( .A(n12674), .B(n12675), .Z(n12297) );
  XNOR U14033 ( .A(round_reg[1428]), .B(round_reg[1108]), .Z(n12675) );
  XOR U14034 ( .A(round_reg[148]), .B(n12676), .Z(n12674) );
  XOR U14035 ( .A(round_reg[788]), .B(round_reg[468]), .Z(n12676) );
  XNOR U14036 ( .A(n12677), .B(n6911), .Z(n2670) );
  XOR U14037 ( .A(round_reg[1174]), .B(n10666), .Z(n6911) );
  IV U14038 ( .A(n9750), .Z(n10666) );
  XOR U14039 ( .A(n12557), .B(n12212), .Z(n9750) );
  XOR U14040 ( .A(n12678), .B(n12679), .Z(n12212) );
  XNOR U14041 ( .A(round_reg[1429]), .B(round_reg[1109]), .Z(n12679) );
  XOR U14042 ( .A(round_reg[149]), .B(n12680), .Z(n12678) );
  XOR U14043 ( .A(round_reg[789]), .B(round_reg[469]), .Z(n12680) );
  XOR U14044 ( .A(n12681), .B(n12682), .Z(n12557) );
  XNOR U14045 ( .A(round_reg[1558]), .B(round_reg[1238]), .Z(n12682) );
  XOR U14046 ( .A(round_reg[278]), .B(n12683), .Z(n12681) );
  XOR U14047 ( .A(round_reg[918]), .B(round_reg[598]), .Z(n12683) );
  AND U14048 ( .A(n6912), .B(n12684), .Z(n12677) );
  XNOR U14049 ( .A(n3343), .B(n12685), .Z(n12656) );
  XNOR U14050 ( .A(n5368), .B(n6901), .Z(n12685) );
  XNOR U14051 ( .A(n12686), .B(n6917), .Z(n6901) );
  XOR U14052 ( .A(round_reg[1246]), .B(n9473), .Z(n6917) );
  XNOR U14053 ( .A(n11955), .B(n11708), .Z(n9473) );
  XOR U14054 ( .A(n12687), .B(n12688), .Z(n11708) );
  XNOR U14055 ( .A(round_reg[30]), .B(round_reg[1310]), .Z(n12688) );
  XOR U14056 ( .A(round_reg[350]), .B(n12689), .Z(n12687) );
  XOR U14057 ( .A(round_reg[990]), .B(round_reg[670]), .Z(n12689) );
  XOR U14058 ( .A(n12690), .B(n12691), .Z(n11955) );
  XNOR U14059 ( .A(round_reg[1501]), .B(round_reg[1181]), .Z(n12691) );
  XOR U14060 ( .A(round_reg[221]), .B(n12692), .Z(n12690) );
  XOR U14061 ( .A(round_reg[861]), .B(round_reg[541]), .Z(n12692) );
  NOR U14062 ( .A(n6916), .B(n7681), .Z(n12686) );
  XNOR U14063 ( .A(round_reg[499]), .B(n10524), .Z(n7681) );
  XOR U14064 ( .A(n11455), .B(n11842), .Z(n10524) );
  XOR U14065 ( .A(n12693), .B(n12694), .Z(n11842) );
  XNOR U14066 ( .A(round_reg[114]), .B(round_reg[1074]), .Z(n12694) );
  XOR U14067 ( .A(round_reg[1394]), .B(n12695), .Z(n12693) );
  XOR U14068 ( .A(round_reg[754]), .B(round_reg[434]), .Z(n12695) );
  XOR U14069 ( .A(n12696), .B(n12697), .Z(n11455) );
  XNOR U14070 ( .A(round_reg[1523]), .B(round_reg[1203]), .Z(n12697) );
  XOR U14071 ( .A(round_reg[243]), .B(n12698), .Z(n12696) );
  XOR U14072 ( .A(round_reg[883]), .B(round_reg[563]), .Z(n12698) );
  XNOR U14073 ( .A(round_reg[888]), .B(n10351), .Z(n6916) );
  IV U14074 ( .A(n10451), .Z(n10351) );
  XNOR U14075 ( .A(n12699), .B(n12369), .Z(n10451) );
  XNOR U14076 ( .A(n12700), .B(n12701), .Z(n12369) );
  XNOR U14077 ( .A(round_reg[1463]), .B(round_reg[1143]), .Z(n12701) );
  XOR U14078 ( .A(round_reg[183]), .B(n12702), .Z(n12700) );
  XOR U14079 ( .A(round_reg[823]), .B(round_reg[503]), .Z(n12702) );
  XNOR U14080 ( .A(n12703), .B(n6921), .Z(n5368) );
  XNOR U14081 ( .A(round_reg[1035]), .B(n9692), .Z(n6921) );
  IV U14082 ( .A(n10356), .Z(n9692) );
  XOR U14083 ( .A(n12001), .B(n11853), .Z(n10356) );
  XOR U14084 ( .A(n12704), .B(n12705), .Z(n11853) );
  XNOR U14085 ( .A(round_reg[139]), .B(round_reg[1099]), .Z(n12705) );
  XOR U14086 ( .A(round_reg[1419]), .B(n12706), .Z(n12704) );
  XOR U14087 ( .A(round_reg[779]), .B(round_reg[459]), .Z(n12706) );
  XOR U14088 ( .A(n12707), .B(n12708), .Z(n12001) );
  XNOR U14089 ( .A(round_reg[1290]), .B(round_reg[10]), .Z(n12708) );
  XOR U14090 ( .A(round_reg[330]), .B(n12709), .Z(n12707) );
  XOR U14091 ( .A(round_reg[970]), .B(round_reg[650]), .Z(n12709) );
  ANDN U14092 ( .B(n6920), .A(n9772), .Z(n12703) );
  XNOR U14093 ( .A(round_reg[601]), .B(n11103), .Z(n9772) );
  XNOR U14094 ( .A(n11485), .B(n12125), .Z(n11103) );
  XNOR U14095 ( .A(n12710), .B(n12711), .Z(n12125) );
  XNOR U14096 ( .A(round_reg[1496]), .B(round_reg[1176]), .Z(n12711) );
  XOR U14097 ( .A(round_reg[216]), .B(n12712), .Z(n12710) );
  XOR U14098 ( .A(round_reg[856]), .B(round_reg[536]), .Z(n12712) );
  XOR U14099 ( .A(n12713), .B(n12714), .Z(n11485) );
  XNOR U14100 ( .A(round_reg[25]), .B(round_reg[1305]), .Z(n12714) );
  XOR U14101 ( .A(round_reg[345]), .B(n12715), .Z(n12713) );
  XOR U14102 ( .A(round_reg[985]), .B(round_reg[665]), .Z(n12715) );
  XOR U14103 ( .A(round_reg[667]), .B(n9975), .Z(n6920) );
  XOR U14104 ( .A(n12162), .B(n11288), .Z(n9975) );
  XNOR U14105 ( .A(n12716), .B(n12717), .Z(n11288) );
  XNOR U14106 ( .A(round_reg[1562]), .B(round_reg[1242]), .Z(n12717) );
  XOR U14107 ( .A(round_reg[282]), .B(n12718), .Z(n12716) );
  XOR U14108 ( .A(round_reg[922]), .B(round_reg[602]), .Z(n12718) );
  XOR U14109 ( .A(n12719), .B(n12720), .Z(n12162) );
  XNOR U14110 ( .A(round_reg[1371]), .B(round_reg[1051]), .Z(n12720) );
  XOR U14111 ( .A(round_reg[411]), .B(n12721), .Z(n12719) );
  XOR U14112 ( .A(round_reg[91]), .B(round_reg[731]), .Z(n12721) );
  XNOR U14113 ( .A(n12722), .B(n6925), .Z(n3343) );
  XNOR U14114 ( .A(round_reg[1148]), .B(n9112), .Z(n6925) );
  IV U14115 ( .A(n10102), .Z(n9112) );
  XOR U14116 ( .A(n12723), .B(n11650), .Z(n10102) );
  XOR U14117 ( .A(n12724), .B(n12725), .Z(n11650) );
  XNOR U14118 ( .A(round_reg[1532]), .B(round_reg[1212]), .Z(n12725) );
  XOR U14119 ( .A(round_reg[252]), .B(n12726), .Z(n12724) );
  XOR U14120 ( .A(round_reg[892]), .B(round_reg[572]), .Z(n12726) );
  ANDN U14121 ( .B(n6924), .A(n7677), .Z(n12722) );
  XNOR U14122 ( .A(round_reg[378]), .B(n11675), .Z(n7677) );
  XNOR U14123 ( .A(round_reg[745]), .B(n9552), .Z(n6924) );
  XNOR U14124 ( .A(n12136), .B(n11993), .Z(n9552) );
  XNOR U14125 ( .A(n12727), .B(n12728), .Z(n11993) );
  XNOR U14126 ( .A(round_reg[1449]), .B(round_reg[1129]), .Z(n12728) );
  XOR U14127 ( .A(round_reg[169]), .B(n12729), .Z(n12727) );
  XOR U14128 ( .A(round_reg[809]), .B(round_reg[489]), .Z(n12729) );
  XOR U14129 ( .A(n12730), .B(n12731), .Z(n12136) );
  XNOR U14130 ( .A(round_reg[1320]), .B(round_reg[1000]), .Z(n12731) );
  XOR U14131 ( .A(round_reg[360]), .B(n12732), .Z(n12730) );
  XOR U14132 ( .A(round_reg[680]), .B(round_reg[40]), .Z(n12732) );
  XOR U14133 ( .A(n12733), .B(n12734), .Z(n6023) );
  XNOR U14134 ( .A(n1844), .B(n5221), .Z(n12734) );
  XOR U14135 ( .A(n12735), .B(n7756), .Z(n5221) );
  XNOR U14136 ( .A(round_reg[498]), .B(n10617), .Z(n7756) );
  IV U14137 ( .A(n11414), .Z(n10617) );
  XOR U14138 ( .A(n12041), .B(n11560), .Z(n11414) );
  XNOR U14139 ( .A(n12736), .B(n12737), .Z(n11560) );
  XNOR U14140 ( .A(round_reg[1522]), .B(round_reg[1202]), .Z(n12737) );
  XOR U14141 ( .A(round_reg[242]), .B(n12738), .Z(n12736) );
  XOR U14142 ( .A(round_reg[882]), .B(round_reg[562]), .Z(n12738) );
  XOR U14143 ( .A(n12739), .B(n12740), .Z(n12041) );
  XNOR U14144 ( .A(round_reg[113]), .B(round_reg[1073]), .Z(n12740) );
  XOR U14145 ( .A(round_reg[1393]), .B(n12741), .Z(n12739) );
  XOR U14146 ( .A(round_reg[753]), .B(round_reg[433]), .Z(n12741) );
  ANDN U14147 ( .B(n7663), .A(n6957), .Z(n12735) );
  XNOR U14148 ( .A(round_reg[1318]), .B(n10883), .Z(n6957) );
  XNOR U14149 ( .A(n11773), .B(n11492), .Z(n10883) );
  XNOR U14150 ( .A(n12742), .B(n12743), .Z(n11492) );
  XNOR U14151 ( .A(round_reg[1573]), .B(round_reg[1253]), .Z(n12743) );
  XOR U14152 ( .A(round_reg[293]), .B(n12744), .Z(n12742) );
  XOR U14153 ( .A(round_reg[933]), .B(round_reg[613]), .Z(n12744) );
  XOR U14154 ( .A(n12745), .B(n12746), .Z(n11773) );
  XNOR U14155 ( .A(round_reg[1062]), .B(round_reg[102]), .Z(n12746) );
  XOR U14156 ( .A(round_reg[1382]), .B(n12747), .Z(n12745) );
  XOR U14157 ( .A(round_reg[742]), .B(round_reg[422]), .Z(n12747) );
  XOR U14158 ( .A(round_reg[73]), .B(n9916), .Z(n7663) );
  IV U14159 ( .A(n11021), .Z(n9916) );
  XNOR U14160 ( .A(n12748), .B(n12352), .Z(n11021) );
  XNOR U14161 ( .A(n12749), .B(n12750), .Z(n12352) );
  XNOR U14162 ( .A(round_reg[137]), .B(round_reg[1097]), .Z(n12750) );
  XOR U14163 ( .A(round_reg[1417]), .B(n12751), .Z(n12749) );
  XOR U14164 ( .A(round_reg[777]), .B(round_reg[457]), .Z(n12751) );
  XNOR U14165 ( .A(n12752), .B(n7752), .Z(n1844) );
  XNOR U14166 ( .A(round_reg[377]), .B(n9389), .Z(n7752) );
  IV U14167 ( .A(n11847), .Z(n9389) );
  XOR U14168 ( .A(n12699), .B(n12753), .Z(n11847) );
  XOR U14169 ( .A(n12754), .B(n12755), .Z(n12699) );
  XNOR U14170 ( .A(round_reg[1592]), .B(round_reg[1272]), .Z(n12755) );
  XOR U14171 ( .A(round_reg[312]), .B(n12756), .Z(n12754) );
  XOR U14172 ( .A(round_reg[952]), .B(round_reg[632]), .Z(n12756) );
  ANDN U14173 ( .B(n7670), .A(n6950), .Z(n12752) );
  XNOR U14174 ( .A(round_reg[1472]), .B(n11749), .Z(n6950) );
  XOR U14175 ( .A(n12757), .B(n12448), .Z(n11749) );
  XOR U14176 ( .A(n12758), .B(n12759), .Z(n12448) );
  XNOR U14177 ( .A(round_reg[1471]), .B(round_reg[1151]), .Z(n12759) );
  XOR U14178 ( .A(round_reg[191]), .B(n12760), .Z(n12758) );
  XOR U14179 ( .A(round_reg[831]), .B(round_reg[511]), .Z(n12760) );
  XNOR U14180 ( .A(round_reg[303]), .B(n11210), .Z(n7670) );
  XNOR U14181 ( .A(n12761), .B(n12638), .Z(n11210) );
  XNOR U14182 ( .A(n12762), .B(n12763), .Z(n12638) );
  XNOR U14183 ( .A(round_reg[1518]), .B(round_reg[1198]), .Z(n12763) );
  XOR U14184 ( .A(round_reg[238]), .B(n12764), .Z(n12762) );
  XOR U14185 ( .A(round_reg[878]), .B(round_reg[558]), .Z(n12764) );
  XNOR U14186 ( .A(n4068), .B(n12765), .Z(n12733) );
  XOR U14187 ( .A(n7732), .B(n3606), .Z(n12765) );
  XOR U14188 ( .A(n12766), .B(n9846), .Z(n3606) );
  XNOR U14189 ( .A(round_reg[600]), .B(n11184), .Z(n9846) );
  IV U14190 ( .A(n10302), .Z(n11184) );
  XOR U14191 ( .A(n11598), .B(n12767), .Z(n10302) );
  XOR U14192 ( .A(n12768), .B(n12769), .Z(n11598) );
  XNOR U14193 ( .A(round_reg[24]), .B(round_reg[1304]), .Z(n12769) );
  XOR U14194 ( .A(round_reg[344]), .B(n12770), .Z(n12768) );
  XOR U14195 ( .A(round_reg[984]), .B(round_reg[664]), .Z(n12770) );
  ANDN U14196 ( .B(n7668), .A(n6946), .Z(n12766) );
  XNOR U14197 ( .A(round_reg[1411]), .B(n11387), .Z(n6946) );
  IV U14198 ( .A(n9266), .Z(n11387) );
  XOR U14199 ( .A(n11914), .B(n11921), .Z(n9266) );
  XNOR U14200 ( .A(n12771), .B(n12772), .Z(n11921) );
  XNOR U14201 ( .A(round_reg[1346]), .B(round_reg[1026]), .Z(n12772) );
  XOR U14202 ( .A(round_reg[386]), .B(n12773), .Z(n12771) );
  XOR U14203 ( .A(round_reg[706]), .B(round_reg[66]), .Z(n12773) );
  XOR U14204 ( .A(n12774), .B(n12775), .Z(n11914) );
  XNOR U14205 ( .A(round_reg[1475]), .B(round_reg[1155]), .Z(n12775) );
  XOR U14206 ( .A(round_reg[195]), .B(n12776), .Z(n12774) );
  XOR U14207 ( .A(round_reg[835]), .B(round_reg[515]), .Z(n12776) );
  XOR U14208 ( .A(round_reg[255]), .B(n12145), .Z(n7668) );
  XNOR U14209 ( .A(round_reg[428]), .B(n9616), .Z(n7750) );
  AND U14210 ( .A(n7672), .B(n12778), .Z(n12777) );
  IV U14211 ( .A(n6935), .Z(n12778) );
  XOR U14212 ( .A(round_reg[1537]), .B(n9676), .Z(n6935) );
  IV U14213 ( .A(n11240), .Z(n9676) );
  XOR U14214 ( .A(n12779), .B(n12780), .Z(n12652) );
  XNOR U14215 ( .A(round_reg[1472]), .B(round_reg[1152]), .Z(n12780) );
  XOR U14216 ( .A(round_reg[192]), .B(n12781), .Z(n12779) );
  XOR U14217 ( .A(round_reg[832]), .B(round_reg[512]), .Z(n12781) );
  XNOR U14218 ( .A(n12782), .B(n12783), .Z(n11717) );
  XNOR U14219 ( .A(round_reg[1]), .B(round_reg[1281]), .Z(n12783) );
  XOR U14220 ( .A(round_reg[321]), .B(n12784), .Z(n12782) );
  XOR U14221 ( .A(round_reg[961]), .B(round_reg[641]), .Z(n12784) );
  XNOR U14222 ( .A(round_reg[51]), .B(n9437), .Z(n7672) );
  XOR U14223 ( .A(n11226), .B(n11069), .Z(n9437) );
  XOR U14224 ( .A(n12785), .B(n12786), .Z(n11069) );
  XNOR U14225 ( .A(round_reg[1586]), .B(round_reg[1266]), .Z(n12786) );
  XOR U14226 ( .A(round_reg[306]), .B(n12787), .Z(n12785) );
  XOR U14227 ( .A(round_reg[946]), .B(round_reg[626]), .Z(n12787) );
  XOR U14228 ( .A(n12788), .B(n12789), .Z(n11226) );
  XNOR U14229 ( .A(round_reg[115]), .B(round_reg[1075]), .Z(n12789) );
  XOR U14230 ( .A(round_reg[1395]), .B(n12790), .Z(n12788) );
  XOR U14231 ( .A(round_reg[755]), .B(round_reg[435]), .Z(n12790) );
  XNOR U14232 ( .A(n12791), .B(n7758), .Z(n4068) );
  XOR U14233 ( .A(round_reg[532]), .B(n10837), .Z(n7758) );
  XNOR U14234 ( .A(n12318), .B(n11310), .Z(n10837) );
  XNOR U14235 ( .A(n12792), .B(n12793), .Z(n11310) );
  XNOR U14236 ( .A(round_reg[1556]), .B(round_reg[1236]), .Z(n12793) );
  XOR U14237 ( .A(round_reg[276]), .B(n12794), .Z(n12792) );
  XOR U14238 ( .A(round_reg[916]), .B(round_reg[596]), .Z(n12794) );
  XOR U14239 ( .A(n12795), .B(n12796), .Z(n12318) );
  XNOR U14240 ( .A(round_reg[1427]), .B(round_reg[1107]), .Z(n12796) );
  XOR U14241 ( .A(round_reg[147]), .B(n12797), .Z(n12795) );
  XOR U14242 ( .A(round_reg[787]), .B(round_reg[467]), .Z(n12797) );
  ANDN U14243 ( .B(n7665), .A(n6932), .Z(n12791) );
  XNOR U14244 ( .A(round_reg[1381]), .B(n10958), .Z(n6932) );
  IV U14245 ( .A(n11113), .Z(n10958) );
  XOR U14246 ( .A(n12798), .B(n11399), .Z(n11113) );
  XNOR U14247 ( .A(n12799), .B(n12800), .Z(n11399) );
  XNOR U14248 ( .A(round_reg[1445]), .B(round_reg[1125]), .Z(n12800) );
  XOR U14249 ( .A(round_reg[165]), .B(n12801), .Z(n12799) );
  XOR U14250 ( .A(round_reg[805]), .B(round_reg[485]), .Z(n12801) );
  XOR U14251 ( .A(round_reg[132]), .B(n11242), .Z(n7665) );
  IV U14252 ( .A(n9186), .Z(n11242) );
  XOR U14253 ( .A(n11737), .B(n11726), .Z(n9186) );
  XOR U14254 ( .A(n12802), .B(n12803), .Z(n11726) );
  XNOR U14255 ( .A(round_reg[1476]), .B(round_reg[1156]), .Z(n12803) );
  XOR U14256 ( .A(round_reg[196]), .B(n12804), .Z(n12802) );
  XOR U14257 ( .A(round_reg[836]), .B(round_reg[516]), .Z(n12804) );
  XOR U14258 ( .A(n12805), .B(n12806), .Z(n11737) );
  XNOR U14259 ( .A(round_reg[1347]), .B(round_reg[1027]), .Z(n12806) );
  XOR U14260 ( .A(round_reg[387]), .B(n12807), .Z(n12805) );
  XOR U14261 ( .A(round_reg[707]), .B(round_reg[67]), .Z(n12807) );
  XOR U14262 ( .A(n12808), .B(n6912), .Z(n7675) );
  XOR U14263 ( .A(round_reg[791]), .B(n11000), .Z(n6912) );
  IV U14264 ( .A(n10927), .Z(n11000) );
  XNOR U14265 ( .A(n12577), .B(n12767), .Z(n10927) );
  XNOR U14266 ( .A(n12809), .B(n12810), .Z(n12767) );
  XNOR U14267 ( .A(round_reg[1495]), .B(round_reg[1175]), .Z(n12810) );
  XOR U14268 ( .A(round_reg[215]), .B(n12811), .Z(n12809) );
  XOR U14269 ( .A(round_reg[855]), .B(round_reg[535]), .Z(n12811) );
  XOR U14270 ( .A(n12812), .B(n12813), .Z(n12577) );
  XNOR U14271 ( .A(round_reg[1366]), .B(round_reg[1046]), .Z(n12813) );
  XOR U14272 ( .A(round_reg[406]), .B(n12814), .Z(n12812) );
  XOR U14273 ( .A(round_reg[86]), .B(round_reg[726]), .Z(n12814) );
  NOR U14274 ( .A(n12684), .B(n7601), .Z(n12808) );
  XNOR U14275 ( .A(round_reg[52]), .B(n11189), .Z(n7601) );
  IV U14276 ( .A(n9774), .Z(n12684) );
  XOR U14277 ( .A(round_reg[429]), .B(n9535), .Z(n9774) );
  IV U14278 ( .A(n10984), .Z(n9535) );
  XOR U14279 ( .A(n1803), .B(n9209), .Z(n4043) );
  XOR U14280 ( .A(n12815), .B(n9258), .Z(n9209) );
  AND U14281 ( .A(n6711), .B(n7183), .Z(n12815) );
  XOR U14282 ( .A(round_reg[1389]), .B(n10984), .Z(n6711) );
  XOR U14283 ( .A(n11422), .B(n12098), .Z(n10984) );
  XOR U14284 ( .A(n12816), .B(n12817), .Z(n12098) );
  XNOR U14285 ( .A(round_reg[1324]), .B(round_reg[1004]), .Z(n12817) );
  XOR U14286 ( .A(round_reg[364]), .B(n12818), .Z(n12816) );
  XOR U14287 ( .A(round_reg[684]), .B(round_reg[44]), .Z(n12818) );
  XOR U14288 ( .A(n12819), .B(n12820), .Z(n11422) );
  XNOR U14289 ( .A(round_reg[1453]), .B(round_reg[1133]), .Z(n12820) );
  XOR U14290 ( .A(round_reg[173]), .B(n12821), .Z(n12819) );
  XOR U14291 ( .A(round_reg[813]), .B(round_reg[493]), .Z(n12821) );
  IV U14292 ( .A(n5186), .Z(n1803) );
  XOR U14293 ( .A(n6681), .B(n6419), .Z(n5186) );
  XOR U14294 ( .A(n12822), .B(n12823), .Z(n6419) );
  XOR U14295 ( .A(n5982), .B(n4270), .Z(n12823) );
  XOR U14296 ( .A(n12824), .B(n7276), .Z(n4270) );
  XOR U14297 ( .A(round_reg[310]), .B(n10696), .Z(n7276) );
  XOR U14298 ( .A(n12368), .B(n11150), .Z(n10696) );
  XNOR U14299 ( .A(n12825), .B(n12826), .Z(n11150) );
  XNOR U14300 ( .A(round_reg[1525]), .B(round_reg[1205]), .Z(n12826) );
  XOR U14301 ( .A(round_reg[245]), .B(n12827), .Z(n12825) );
  XOR U14302 ( .A(round_reg[885]), .B(round_reg[565]), .Z(n12827) );
  XOR U14303 ( .A(n12828), .B(n12829), .Z(n12368) );
  XNOR U14304 ( .A(round_reg[1334]), .B(round_reg[1014]), .Z(n12829) );
  XOR U14305 ( .A(round_reg[374]), .B(n12830), .Z(n12828) );
  XOR U14306 ( .A(round_reg[694]), .B(round_reg[54]), .Z(n12830) );
  ANDN U14307 ( .B(n6754), .A(n6755), .Z(n12824) );
  XOR U14308 ( .A(round_reg[1090]), .B(n9859), .Z(n6755) );
  XOR U14309 ( .A(n12117), .B(n12831), .Z(n9859) );
  XOR U14310 ( .A(n12832), .B(n12833), .Z(n12117) );
  XNOR U14311 ( .A(round_reg[1474]), .B(round_reg[1154]), .Z(n12833) );
  XOR U14312 ( .A(round_reg[194]), .B(n12834), .Z(n12832) );
  XOR U14313 ( .A(round_reg[834]), .B(round_reg[514]), .Z(n12834) );
  XNOR U14314 ( .A(round_reg[1479]), .B(n11043), .Z(n6754) );
  IV U14315 ( .A(n11133), .Z(n11043) );
  XNOR U14316 ( .A(n12835), .B(n7284), .Z(n5982) );
  XOR U14317 ( .A(round_reg[139]), .B(n9208), .Z(n7284) );
  XNOR U14318 ( .A(n11582), .B(n12357), .Z(n9208) );
  XOR U14319 ( .A(n12836), .B(n12837), .Z(n12357) );
  XNOR U14320 ( .A(round_reg[1483]), .B(round_reg[1163]), .Z(n12837) );
  XOR U14321 ( .A(round_reg[203]), .B(n12838), .Z(n12836) );
  XOR U14322 ( .A(round_reg[843]), .B(round_reg[523]), .Z(n12838) );
  XOR U14323 ( .A(n12839), .B(n12840), .Z(n11582) );
  XNOR U14324 ( .A(round_reg[1354]), .B(round_reg[1034]), .Z(n12840) );
  XOR U14325 ( .A(round_reg[394]), .B(n12841), .Z(n12839) );
  XOR U14326 ( .A(round_reg[74]), .B(round_reg[714]), .Z(n12841) );
  ANDN U14327 ( .B(n6737), .A(n6738), .Z(n12835) );
  XOR U14328 ( .A(round_reg[1012]), .B(n10297), .Z(n6738) );
  IV U14329 ( .A(n11189), .Z(n10297) );
  XNOR U14330 ( .A(n11149), .B(n12629), .Z(n11189) );
  XNOR U14331 ( .A(n12842), .B(n12843), .Z(n12629) );
  XNOR U14332 ( .A(round_reg[1587]), .B(round_reg[1267]), .Z(n12843) );
  XOR U14333 ( .A(round_reg[307]), .B(n12844), .Z(n12842) );
  XOR U14334 ( .A(round_reg[947]), .B(round_reg[627]), .Z(n12844) );
  XOR U14335 ( .A(n12845), .B(n12846), .Z(n11149) );
  XNOR U14336 ( .A(round_reg[116]), .B(round_reg[1076]), .Z(n12846) );
  XOR U14337 ( .A(round_reg[1396]), .B(n12847), .Z(n12845) );
  XOR U14338 ( .A(round_reg[756]), .B(round_reg[436]), .Z(n12847) );
  XOR U14339 ( .A(round_reg[1388]), .B(n9616), .Z(n6737) );
  XOR U14340 ( .A(n12848), .B(n12849), .Z(n11522) );
  XNOR U14341 ( .A(round_reg[1452]), .B(round_reg[1132]), .Z(n12849) );
  XOR U14342 ( .A(round_reg[172]), .B(n12850), .Z(n12848) );
  XOR U14343 ( .A(round_reg[812]), .B(round_reg[492]), .Z(n12850) );
  XNOR U14344 ( .A(n12851), .B(n12852), .Z(n12598) );
  XNOR U14345 ( .A(round_reg[1323]), .B(round_reg[1003]), .Z(n12852) );
  XOR U14346 ( .A(round_reg[363]), .B(n12853), .Z(n12851) );
  XOR U14347 ( .A(round_reg[683]), .B(round_reg[43]), .Z(n12853) );
  XOR U14348 ( .A(n3703), .B(n12854), .Z(n12822) );
  XOR U14349 ( .A(n5506), .B(n2158), .Z(n12854) );
  XNOR U14350 ( .A(n12855), .B(n7281), .Z(n2158) );
  XOR U14351 ( .A(round_reg[80]), .B(n9447), .Z(n7281) );
  IV U14352 ( .A(n9898), .Z(n9447) );
  XOR U14353 ( .A(n11682), .B(n11258), .Z(n9898) );
  XOR U14354 ( .A(n12856), .B(n12857), .Z(n11258) );
  XNOR U14355 ( .A(round_reg[1424]), .B(round_reg[1104]), .Z(n12857) );
  XOR U14356 ( .A(round_reg[144]), .B(n12858), .Z(n12856) );
  XOR U14357 ( .A(round_reg[784]), .B(round_reg[464]), .Z(n12858) );
  XOR U14358 ( .A(n12859), .B(n12860), .Z(n11682) );
  XNOR U14359 ( .A(round_reg[15]), .B(round_reg[1295]), .Z(n12860) );
  XOR U14360 ( .A(round_reg[335]), .B(n12861), .Z(n12859) );
  XOR U14361 ( .A(round_reg[975]), .B(round_reg[655]), .Z(n12861) );
  ANDN U14362 ( .B(n6746), .A(n6747), .Z(n12855) );
  XOR U14363 ( .A(round_reg[1252]), .B(n10431), .Z(n6747) );
  IV U14364 ( .A(n10105), .Z(n10431) );
  XOR U14365 ( .A(n11804), .B(n12798), .Z(n10105) );
  XOR U14366 ( .A(n12862), .B(n12863), .Z(n12798) );
  XNOR U14367 ( .A(round_reg[356]), .B(round_reg[1316]), .Z(n12863) );
  XOR U14368 ( .A(round_reg[36]), .B(n12864), .Z(n12862) );
  XOR U14369 ( .A(round_reg[996]), .B(round_reg[676]), .Z(n12864) );
  XOR U14370 ( .A(n12865), .B(n12866), .Z(n11804) );
  XNOR U14371 ( .A(round_reg[1507]), .B(round_reg[1187]), .Z(n12866) );
  XOR U14372 ( .A(round_reg[227]), .B(n12867), .Z(n12865) );
  XOR U14373 ( .A(round_reg[867]), .B(round_reg[547]), .Z(n12867) );
  XNOR U14374 ( .A(round_reg[1325]), .B(n10873), .Z(n6746) );
  XNOR U14375 ( .A(n12637), .B(n11637), .Z(n10873) );
  XNOR U14376 ( .A(n12868), .B(n12869), .Z(n11637) );
  XNOR U14377 ( .A(round_reg[1580]), .B(round_reg[1260]), .Z(n12869) );
  XOR U14378 ( .A(round_reg[300]), .B(n12870), .Z(n12868) );
  XOR U14379 ( .A(round_reg[940]), .B(round_reg[620]), .Z(n12870) );
  XOR U14380 ( .A(n12871), .B(n12872), .Z(n12637) );
  XNOR U14381 ( .A(round_reg[109]), .B(round_reg[1069]), .Z(n12872) );
  XOR U14382 ( .A(round_reg[1389]), .B(n12873), .Z(n12871) );
  XOR U14383 ( .A(round_reg[749]), .B(round_reg[429]), .Z(n12873) );
  XNOR U14384 ( .A(n12874), .B(n9272), .Z(n5506) );
  XOR U14385 ( .A(round_reg[198]), .B(n11212), .Z(n9272) );
  IV U14386 ( .A(n9386), .Z(n11212) );
  XOR U14387 ( .A(n12875), .B(n12876), .Z(n12108) );
  XNOR U14388 ( .A(round_reg[1542]), .B(round_reg[1222]), .Z(n12876) );
  XOR U14389 ( .A(round_reg[262]), .B(n12877), .Z(n12875) );
  XOR U14390 ( .A(round_reg[902]), .B(round_reg[582]), .Z(n12877) );
  XNOR U14391 ( .A(n12878), .B(n12879), .Z(n12633) );
  XNOR U14392 ( .A(round_reg[133]), .B(round_reg[1093]), .Z(n12879) );
  XOR U14393 ( .A(round_reg[1413]), .B(n12880), .Z(n12878) );
  XOR U14394 ( .A(round_reg[773]), .B(round_reg[453]), .Z(n12880) );
  NOR U14395 ( .A(n6750), .B(n6751), .Z(n12874) );
  XOR U14396 ( .A(round_reg[1041]), .B(n9829), .Z(n6751) );
  XOR U14397 ( .A(round_reg[1418]), .B(n9393), .Z(n6750) );
  XNOR U14398 ( .A(n11719), .B(n12312), .Z(n9393) );
  XNOR U14399 ( .A(n12881), .B(n12882), .Z(n12312) );
  XNOR U14400 ( .A(round_reg[1482]), .B(round_reg[1162]), .Z(n12882) );
  XOR U14401 ( .A(round_reg[202]), .B(n12883), .Z(n12881) );
  XOR U14402 ( .A(round_reg[842]), .B(round_reg[522]), .Z(n12883) );
  XOR U14403 ( .A(n12884), .B(n12885), .Z(n11719) );
  XNOR U14404 ( .A(round_reg[1353]), .B(round_reg[1033]), .Z(n12885) );
  XOR U14405 ( .A(round_reg[393]), .B(n12886), .Z(n12884) );
  XOR U14406 ( .A(round_reg[73]), .B(round_reg[713]), .Z(n12886) );
  XNOR U14407 ( .A(n12887), .B(n7273), .Z(n3703) );
  XOR U14408 ( .A(round_reg[58]), .B(n11034), .Z(n7273) );
  IV U14409 ( .A(n11675), .Z(n11034) );
  XOR U14410 ( .A(n10996), .B(n11004), .Z(n11675) );
  XOR U14411 ( .A(n12888), .B(n12889), .Z(n11004) );
  XNOR U14412 ( .A(round_reg[1593]), .B(round_reg[1273]), .Z(n12889) );
  XOR U14413 ( .A(round_reg[313]), .B(n12890), .Z(n12888) );
  XOR U14414 ( .A(round_reg[953]), .B(round_reg[633]), .Z(n12890) );
  XOR U14415 ( .A(n12891), .B(n12892), .Z(n10996) );
  XNOR U14416 ( .A(round_reg[122]), .B(round_reg[1082]), .Z(n12892) );
  XOR U14417 ( .A(round_reg[1402]), .B(n12893), .Z(n12891) );
  XOR U14418 ( .A(round_reg[762]), .B(round_reg[442]), .Z(n12893) );
  ANDN U14419 ( .B(n6741), .A(n6742), .Z(n12887) );
  XOR U14420 ( .A(round_reg[1180]), .B(n10936), .Z(n6742) );
  XOR U14421 ( .A(round_reg[1544]), .B(n11950), .Z(n6741) );
  IV U14422 ( .A(n9116), .Z(n11950) );
  XOR U14423 ( .A(n11886), .B(n12748), .Z(n9116) );
  XOR U14424 ( .A(n12894), .B(n12895), .Z(n12748) );
  XNOR U14425 ( .A(round_reg[328]), .B(round_reg[1288]), .Z(n12895) );
  XOR U14426 ( .A(round_reg[648]), .B(n12896), .Z(n12894) );
  XOR U14427 ( .A(round_reg[968]), .B(round_reg[8]), .Z(n12896) );
  XOR U14428 ( .A(n12897), .B(n12898), .Z(n11886) );
  XNOR U14429 ( .A(round_reg[1479]), .B(round_reg[1159]), .Z(n12898) );
  XOR U14430 ( .A(round_reg[199]), .B(n12899), .Z(n12897) );
  XOR U14431 ( .A(round_reg[839]), .B(round_reg[519]), .Z(n12899) );
  XOR U14432 ( .A(n12900), .B(n12901), .Z(n6681) );
  XOR U14433 ( .A(n4865), .B(n4016), .Z(n12901) );
  XOR U14434 ( .A(n12902), .B(n6717), .Z(n4016) );
  XOR U14435 ( .A(round_reg[798]), .B(n10357), .Z(n6717) );
  IV U14436 ( .A(n11763), .Z(n10357) );
  XNOR U14437 ( .A(n11989), .B(n11221), .Z(n11763) );
  XNOR U14438 ( .A(n12903), .B(n12904), .Z(n11221) );
  XNOR U14439 ( .A(round_reg[1502]), .B(round_reg[1182]), .Z(n12904) );
  XOR U14440 ( .A(round_reg[222]), .B(n12905), .Z(n12903) );
  XOR U14441 ( .A(round_reg[862]), .B(round_reg[542]), .Z(n12905) );
  XOR U14442 ( .A(n12906), .B(n12907), .Z(n11989) );
  XNOR U14443 ( .A(round_reg[1373]), .B(round_reg[1053]), .Z(n12907) );
  XOR U14444 ( .A(round_reg[413]), .B(n12908), .Z(n12906) );
  XOR U14445 ( .A(round_reg[93]), .B(round_reg[733]), .Z(n12908) );
  ANDN U14446 ( .B(n9215), .A(n7185), .Z(n12902) );
  XOR U14447 ( .A(round_reg[59]), .B(n11545), .Z(n7185) );
  IV U14448 ( .A(n9762), .Z(n11545) );
  XNOR U14449 ( .A(n12723), .B(n10995), .Z(n9762) );
  XNOR U14450 ( .A(n12909), .B(n12910), .Z(n10995) );
  XNOR U14451 ( .A(round_reg[1594]), .B(round_reg[1274]), .Z(n12910) );
  XOR U14452 ( .A(round_reg[314]), .B(n12911), .Z(n12909) );
  XOR U14453 ( .A(round_reg[954]), .B(round_reg[634]), .Z(n12911) );
  XOR U14454 ( .A(n12912), .B(n12913), .Z(n12723) );
  XNOR U14455 ( .A(round_reg[123]), .B(round_reg[1083]), .Z(n12913) );
  XOR U14456 ( .A(round_reg[1403]), .B(n12914), .Z(n12912) );
  XOR U14457 ( .A(round_reg[763]), .B(round_reg[443]), .Z(n12914) );
  XNOR U14458 ( .A(round_reg[436]), .B(n12167), .Z(n9215) );
  XOR U14459 ( .A(n10715), .B(n11559), .Z(n12167) );
  XOR U14460 ( .A(n12915), .B(n12916), .Z(n11559) );
  XNOR U14461 ( .A(round_reg[1331]), .B(round_reg[1011]), .Z(n12916) );
  XOR U14462 ( .A(round_reg[371]), .B(n12917), .Z(n12915) );
  XOR U14463 ( .A(round_reg[691]), .B(round_reg[51]), .Z(n12917) );
  XOR U14464 ( .A(n12918), .B(n12919), .Z(n10715) );
  XNOR U14465 ( .A(round_reg[1460]), .B(round_reg[1140]), .Z(n12919) );
  XOR U14466 ( .A(round_reg[180]), .B(n12920), .Z(n12918) );
  XOR U14467 ( .A(round_reg[820]), .B(round_reg[500]), .Z(n12920) );
  XNOR U14468 ( .A(n12921), .B(n6730), .Z(n4865) );
  XOR U14469 ( .A(round_reg[752]), .B(n9606), .Z(n6730) );
  XNOR U14470 ( .A(n11157), .B(n12761), .Z(n9606) );
  XOR U14471 ( .A(n12922), .B(n12923), .Z(n12761) );
  XNOR U14472 ( .A(round_reg[1327]), .B(round_reg[1007]), .Z(n12923) );
  XOR U14473 ( .A(round_reg[367]), .B(n12924), .Z(n12922) );
  XOR U14474 ( .A(round_reg[687]), .B(round_reg[47]), .Z(n12924) );
  XOR U14475 ( .A(n12925), .B(n12926), .Z(n11157) );
  XNOR U14476 ( .A(round_reg[1456]), .B(round_reg[1136]), .Z(n12926) );
  XOR U14477 ( .A(round_reg[176]), .B(n12927), .Z(n12925) );
  XOR U14478 ( .A(round_reg[816]), .B(round_reg[496]), .Z(n12927) );
  ANDN U14479 ( .B(n9212), .A(n7176), .Z(n12921) );
  XOR U14480 ( .A(round_reg[311]), .B(n10608), .Z(n7176) );
  XOR U14481 ( .A(n11062), .B(n12483), .Z(n10608) );
  XNOR U14482 ( .A(n12928), .B(n12929), .Z(n12483) );
  XNOR U14483 ( .A(round_reg[1335]), .B(round_reg[1015]), .Z(n12929) );
  XOR U14484 ( .A(round_reg[375]), .B(n12930), .Z(n12928) );
  XOR U14485 ( .A(round_reg[695]), .B(round_reg[55]), .Z(n12930) );
  XOR U14486 ( .A(n12931), .B(n12932), .Z(n11062) );
  XNOR U14487 ( .A(round_reg[1526]), .B(round_reg[1206]), .Z(n12932) );
  XOR U14488 ( .A(round_reg[246]), .B(n12933), .Z(n12931) );
  XOR U14489 ( .A(round_reg[886]), .B(round_reg[566]), .Z(n12933) );
  XNOR U14490 ( .A(round_reg[321]), .B(n9966), .Z(n9212) );
  XNOR U14491 ( .A(n12757), .B(n12831), .Z(n9966) );
  XNOR U14492 ( .A(n12934), .B(n12935), .Z(n12831) );
  XNOR U14493 ( .A(round_reg[1345]), .B(round_reg[1025]), .Z(n12935) );
  XOR U14494 ( .A(round_reg[385]), .B(n12936), .Z(n12934) );
  XOR U14495 ( .A(round_reg[705]), .B(round_reg[65]), .Z(n12936) );
  XOR U14496 ( .A(n12937), .B(n12938), .Z(n12757) );
  XNOR U14497 ( .A(round_reg[1536]), .B(round_reg[1216]), .Z(n12938) );
  XOR U14498 ( .A(round_reg[256]), .B(n12939), .Z(n12937) );
  XOR U14499 ( .A(round_reg[896]), .B(round_reg[576]), .Z(n12939) );
  XOR U14500 ( .A(n2579), .B(n12940), .Z(n12900) );
  XOR U14501 ( .A(n3502), .B(n9253), .Z(n12940) );
  XNOR U14502 ( .A(n12941), .B(n6726), .Z(n9253) );
  XOR U14503 ( .A(round_reg[674]), .B(n10799), .Z(n6726) );
  IV U14504 ( .A(n10136), .Z(n10799) );
  XNOR U14505 ( .A(n11805), .B(n12158), .Z(n10136) );
  XNOR U14506 ( .A(n12942), .B(n12943), .Z(n12158) );
  XNOR U14507 ( .A(round_reg[1569]), .B(round_reg[1249]), .Z(n12943) );
  XOR U14508 ( .A(round_reg[289]), .B(n12944), .Z(n12942) );
  XOR U14509 ( .A(round_reg[929]), .B(round_reg[609]), .Z(n12944) );
  XOR U14510 ( .A(n12945), .B(n12946), .Z(n11805) );
  XNOR U14511 ( .A(round_reg[1378]), .B(round_reg[1058]), .Z(n12946) );
  XOR U14512 ( .A(round_reg[418]), .B(n12947), .Z(n12945) );
  XOR U14513 ( .A(round_reg[98]), .B(round_reg[738]), .Z(n12947) );
  ANDN U14514 ( .B(n9207), .A(n7178), .Z(n12941) );
  XOR U14515 ( .A(round_reg[199]), .B(n11133), .Z(n7178) );
  XNOR U14516 ( .A(n12948), .B(n12949), .Z(n11285) );
  XNOR U14517 ( .A(round_reg[134]), .B(round_reg[1094]), .Z(n12949) );
  XOR U14518 ( .A(round_reg[1414]), .B(n12950), .Z(n12948) );
  XOR U14519 ( .A(round_reg[774]), .B(round_reg[454]), .Z(n12950) );
  XNOR U14520 ( .A(n12951), .B(n12952), .Z(n11903) );
  XNOR U14521 ( .A(round_reg[1543]), .B(round_reg[1223]), .Z(n12952) );
  XOR U14522 ( .A(round_reg[263]), .B(n12953), .Z(n12951) );
  XOR U14523 ( .A(round_reg[903]), .B(round_reg[583]), .Z(n12953) );
  XNOR U14524 ( .A(round_reg[608]), .B(n10420), .Z(n9207) );
  XNOR U14525 ( .A(n11608), .B(n11465), .Z(n10420) );
  XNOR U14526 ( .A(n12954), .B(n12955), .Z(n11465) );
  XNOR U14527 ( .A(round_reg[32]), .B(round_reg[1312]), .Z(n12955) );
  XOR U14528 ( .A(round_reg[352]), .B(n12956), .Z(n12954) );
  XOR U14529 ( .A(round_reg[992]), .B(round_reg[672]), .Z(n12956) );
  XOR U14530 ( .A(n12957), .B(n12958), .Z(n11608) );
  XNOR U14531 ( .A(round_reg[1503]), .B(round_reg[1183]), .Z(n12958) );
  XOR U14532 ( .A(round_reg[223]), .B(n12959), .Z(n12957) );
  XOR U14533 ( .A(round_reg[863]), .B(round_reg[543]), .Z(n12959) );
  XNOR U14534 ( .A(n12960), .B(n6722), .Z(n3502) );
  XOR U14535 ( .A(round_reg[895]), .B(n12145), .Z(n6722) );
  IV U14536 ( .A(n9854), .Z(n12145) );
  XNOR U14537 ( .A(n11565), .B(n12487), .Z(n9854) );
  XNOR U14538 ( .A(n12961), .B(n12962), .Z(n12487) );
  XNOR U14539 ( .A(round_reg[1599]), .B(round_reg[1279]), .Z(n12962) );
  XOR U14540 ( .A(round_reg[319]), .B(n12963), .Z(n12961) );
  XOR U14541 ( .A(round_reg[959]), .B(round_reg[639]), .Z(n12963) );
  XOR U14542 ( .A(n12964), .B(n12965), .Z(n11565) );
  XNOR U14543 ( .A(round_reg[1470]), .B(round_reg[1150]), .Z(n12965) );
  XOR U14544 ( .A(round_reg[190]), .B(n12966), .Z(n12964) );
  XOR U14545 ( .A(round_reg[830]), .B(round_reg[510]), .Z(n12966) );
  ANDN U14546 ( .B(n9204), .A(n7181), .Z(n12960) );
  XOR U14547 ( .A(round_reg[81]), .B(n9829), .Z(n7181) );
  XOR U14548 ( .A(n12374), .B(n12528), .Z(n9829) );
  XNOR U14549 ( .A(n12967), .B(n12968), .Z(n12528) );
  XNOR U14550 ( .A(round_reg[1425]), .B(round_reg[1105]), .Z(n12968) );
  XOR U14551 ( .A(round_reg[145]), .B(n12969), .Z(n12967) );
  XOR U14552 ( .A(round_reg[785]), .B(round_reg[465]), .Z(n12969) );
  XOR U14553 ( .A(n12970), .B(n12971), .Z(n12374) );
  XNOR U14554 ( .A(round_reg[16]), .B(round_reg[1296]), .Z(n12971) );
  XOR U14555 ( .A(round_reg[336]), .B(n12972), .Z(n12970) );
  XOR U14556 ( .A(round_reg[976]), .B(round_reg[656]), .Z(n12972) );
  XNOR U14557 ( .A(round_reg[506]), .B(n9918), .Z(n9204) );
  XOR U14558 ( .A(n12973), .B(n12974), .Z(n12514) );
  XNOR U14559 ( .A(round_reg[1530]), .B(round_reg[1210]), .Z(n12974) );
  XOR U14560 ( .A(round_reg[250]), .B(n12975), .Z(n12973) );
  XOR U14561 ( .A(round_reg[890]), .B(round_reg[570]), .Z(n12975) );
  XOR U14562 ( .A(n12976), .B(n12977), .Z(n12753) );
  XNOR U14563 ( .A(round_reg[121]), .B(round_reg[1081]), .Z(n12977) );
  XOR U14564 ( .A(round_reg[1401]), .B(n12978), .Z(n12976) );
  XOR U14565 ( .A(round_reg[761]), .B(round_reg[441]), .Z(n12978) );
  XNOR U14566 ( .A(n12979), .B(n6713), .Z(n2579) );
  XOR U14567 ( .A(round_reg[902]), .B(n9465), .Z(n6713) );
  IV U14568 ( .A(n11521), .Z(n9465) );
  XNOR U14569 ( .A(n12429), .B(n12553), .Z(n11521) );
  XNOR U14570 ( .A(n12980), .B(n12981), .Z(n12553) );
  XNOR U14571 ( .A(round_reg[326]), .B(round_reg[1286]), .Z(n12981) );
  XOR U14572 ( .A(round_reg[646]), .B(n12982), .Z(n12980) );
  XOR U14573 ( .A(round_reg[966]), .B(round_reg[6]), .Z(n12982) );
  XOR U14574 ( .A(n12983), .B(n12984), .Z(n12429) );
  XNOR U14575 ( .A(round_reg[1477]), .B(round_reg[1157]), .Z(n12984) );
  XOR U14576 ( .A(round_reg[197]), .B(n12985), .Z(n12983) );
  XOR U14577 ( .A(round_reg[837]), .B(round_reg[517]), .Z(n12985) );
  ANDN U14578 ( .B(n9258), .A(n7183), .Z(n12979) );
  XOR U14579 ( .A(round_reg[140]), .B(n9083), .Z(n7183) );
  IV U14580 ( .A(n10705), .Z(n9083) );
  XOR U14581 ( .A(n12986), .B(n12987), .Z(n11472) );
  XNOR U14582 ( .A(round_reg[1355]), .B(round_reg[1035]), .Z(n12987) );
  XOR U14583 ( .A(round_reg[395]), .B(n12988), .Z(n12986) );
  XOR U14584 ( .A(round_reg[75]), .B(round_reg[715]), .Z(n12988) );
  XNOR U14585 ( .A(n12989), .B(n12990), .Z(n12054) );
  XNOR U14586 ( .A(round_reg[1484]), .B(round_reg[1164]), .Z(n12990) );
  XOR U14587 ( .A(round_reg[204]), .B(n12991), .Z(n12989) );
  XOR U14588 ( .A(round_reg[844]), .B(round_reg[524]), .Z(n12991) );
  XNOR U14589 ( .A(round_reg[540]), .B(n11001), .Z(n9258) );
  IV U14590 ( .A(n10936), .Z(n11001) );
  XOR U14591 ( .A(n11988), .B(n11395), .Z(n10936) );
  XNOR U14592 ( .A(n12992), .B(n12993), .Z(n11395) );
  XNOR U14593 ( .A(round_reg[1435]), .B(round_reg[1115]), .Z(n12993) );
  XOR U14594 ( .A(round_reg[155]), .B(n12994), .Z(n12992) );
  XOR U14595 ( .A(round_reg[795]), .B(round_reg[475]), .Z(n12994) );
  XOR U14596 ( .A(n12995), .B(n12996), .Z(n11988) );
  XNOR U14597 ( .A(round_reg[1564]), .B(round_reg[1244]), .Z(n12996) );
  XOR U14598 ( .A(round_reg[284]), .B(n12997), .Z(n12995) );
  XOR U14599 ( .A(round_reg[924]), .B(round_reg[604]), .Z(n12997) );
  IV U14600 ( .A(init), .Z(n1038) );
endmodule

