
module mult_N128_CC64 ( clk, rst, a, b, c );
  input [127:0] a;
  input [1:0] b;
  output [255:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654;
  wire   [255:0] sreg;

  DFF \sreg_reg[253]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(sreg[253]) );
  DFF \sreg_reg[252]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(sreg[252]) );
  DFF \sreg_reg[251]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(sreg[251]) );
  DFF \sreg_reg[250]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(sreg[250]) );
  DFF \sreg_reg[249]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(sreg[249]) );
  DFF \sreg_reg[248]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(sreg[248]) );
  DFF \sreg_reg[247]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(sreg[247]) );
  DFF \sreg_reg[246]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(sreg[246]) );
  DFF \sreg_reg[245]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(sreg[245]) );
  DFF \sreg_reg[244]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(sreg[244]) );
  DFF \sreg_reg[243]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(sreg[243]) );
  DFF \sreg_reg[242]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(sreg[242]) );
  DFF \sreg_reg[241]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(sreg[241]) );
  DFF \sreg_reg[240]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(sreg[240]) );
  DFF \sreg_reg[239]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(sreg[239]) );
  DFF \sreg_reg[238]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(sreg[238]) );
  DFF \sreg_reg[237]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(sreg[237]) );
  DFF \sreg_reg[236]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(sreg[236]) );
  DFF \sreg_reg[235]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(sreg[235]) );
  DFF \sreg_reg[234]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(sreg[234]) );
  DFF \sreg_reg[233]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(sreg[233]) );
  DFF \sreg_reg[232]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(sreg[232]) );
  DFF \sreg_reg[231]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(sreg[231]) );
  DFF \sreg_reg[230]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(sreg[230]) );
  DFF \sreg_reg[229]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(sreg[229]) );
  DFF \sreg_reg[228]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(sreg[228]) );
  DFF \sreg_reg[227]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(sreg[227]) );
  DFF \sreg_reg[226]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(sreg[226]) );
  DFF \sreg_reg[225]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(sreg[225]) );
  DFF \sreg_reg[224]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(sreg[224]) );
  DFF \sreg_reg[223]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(sreg[223]) );
  DFF \sreg_reg[222]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(sreg[222]) );
  DFF \sreg_reg[221]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(sreg[221]) );
  DFF \sreg_reg[220]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(sreg[220]) );
  DFF \sreg_reg[219]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(sreg[219]) );
  DFF \sreg_reg[218]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(sreg[218]) );
  DFF \sreg_reg[217]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(sreg[217]) );
  DFF \sreg_reg[216]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(sreg[216]) );
  DFF \sreg_reg[215]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(sreg[215]) );
  DFF \sreg_reg[214]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(sreg[214]) );
  DFF \sreg_reg[213]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(sreg[213]) );
  DFF \sreg_reg[212]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(sreg[212]) );
  DFF \sreg_reg[211]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(sreg[211]) );
  DFF \sreg_reg[210]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(sreg[210]) );
  DFF \sreg_reg[209]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(sreg[209]) );
  DFF \sreg_reg[208]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(sreg[208]) );
  DFF \sreg_reg[207]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(sreg[207]) );
  DFF \sreg_reg[206]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(sreg[206]) );
  DFF \sreg_reg[205]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(sreg[205]) );
  DFF \sreg_reg[204]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(sreg[204]) );
  DFF \sreg_reg[203]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(sreg[203]) );
  DFF \sreg_reg[202]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(sreg[202]) );
  DFF \sreg_reg[201]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(sreg[201]) );
  DFF \sreg_reg[200]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(sreg[200]) );
  DFF \sreg_reg[199]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(sreg[199]) );
  DFF \sreg_reg[198]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(sreg[198]) );
  DFF \sreg_reg[197]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(sreg[197]) );
  DFF \sreg_reg[196]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(sreg[196]) );
  DFF \sreg_reg[195]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(sreg[195]) );
  DFF \sreg_reg[194]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(sreg[194]) );
  DFF \sreg_reg[193]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(sreg[193]) );
  DFF \sreg_reg[192]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(sreg[192]) );
  DFF \sreg_reg[191]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(sreg[191]) );
  DFF \sreg_reg[190]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(sreg[190]) );
  DFF \sreg_reg[189]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(sreg[189]) );
  DFF \sreg_reg[188]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(sreg[188]) );
  DFF \sreg_reg[187]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(sreg[187]) );
  DFF \sreg_reg[186]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(sreg[186]) );
  DFF \sreg_reg[185]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(sreg[185]) );
  DFF \sreg_reg[184]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(sreg[184]) );
  DFF \sreg_reg[183]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(sreg[183]) );
  DFF \sreg_reg[182]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(sreg[182]) );
  DFF \sreg_reg[181]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(sreg[181]) );
  DFF \sreg_reg[180]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(sreg[180]) );
  DFF \sreg_reg[179]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(sreg[179]) );
  DFF \sreg_reg[178]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(sreg[178]) );
  DFF \sreg_reg[177]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(sreg[177]) );
  DFF \sreg_reg[176]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(sreg[176]) );
  DFF \sreg_reg[175]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(sreg[175]) );
  DFF \sreg_reg[174]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(sreg[174]) );
  DFF \sreg_reg[173]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(sreg[173]) );
  DFF \sreg_reg[172]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(sreg[172]) );
  DFF \sreg_reg[171]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(sreg[171]) );
  DFF \sreg_reg[170]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(sreg[170]) );
  DFF \sreg_reg[169]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(sreg[169]) );
  DFF \sreg_reg[168]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(sreg[168]) );
  DFF \sreg_reg[167]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(sreg[167]) );
  DFF \sreg_reg[166]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(sreg[166]) );
  DFF \sreg_reg[165]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(sreg[165]) );
  DFF \sreg_reg[164]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(sreg[164]) );
  DFF \sreg_reg[163]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(sreg[163]) );
  DFF \sreg_reg[162]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(sreg[162]) );
  DFF \sreg_reg[161]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(sreg[161]) );
  DFF \sreg_reg[160]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(sreg[160]) );
  DFF \sreg_reg[159]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(sreg[159]) );
  DFF \sreg_reg[158]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(sreg[158]) );
  DFF \sreg_reg[157]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(sreg[157]) );
  DFF \sreg_reg[156]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(sreg[156]) );
  DFF \sreg_reg[155]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(sreg[155]) );
  DFF \sreg_reg[154]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(sreg[154]) );
  DFF \sreg_reg[153]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(sreg[153]) );
  DFF \sreg_reg[152]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(sreg[152]) );
  DFF \sreg_reg[151]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(sreg[151]) );
  DFF \sreg_reg[150]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(sreg[150]) );
  DFF \sreg_reg[149]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(sreg[149]) );
  DFF \sreg_reg[148]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(sreg[148]) );
  DFF \sreg_reg[147]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(sreg[147]) );
  DFF \sreg_reg[146]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(sreg[146]) );
  DFF \sreg_reg[145]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(sreg[145]) );
  DFF \sreg_reg[144]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(sreg[144]) );
  DFF \sreg_reg[143]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(sreg[143]) );
  DFF \sreg_reg[142]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(sreg[142]) );
  DFF \sreg_reg[141]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(sreg[141]) );
  DFF \sreg_reg[140]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(sreg[140]) );
  DFF \sreg_reg[139]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(sreg[139]) );
  DFF \sreg_reg[138]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(sreg[138]) );
  DFF \sreg_reg[137]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(sreg[137]) );
  DFF \sreg_reg[136]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(sreg[136]) );
  DFF \sreg_reg[135]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(sreg[135]) );
  DFF \sreg_reg[134]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(sreg[134]) );
  DFF \sreg_reg[133]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(sreg[133]) );
  DFF \sreg_reg[132]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(sreg[132]) );
  DFF \sreg_reg[131]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(sreg[131]) );
  DFF \sreg_reg[130]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(sreg[130]) );
  DFF \sreg_reg[129]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(sreg[129]) );
  DFF \sreg_reg[128]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(sreg[128]) );
  DFF \sreg_reg[127]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(sreg[127]) );
  DFF \sreg_reg[126]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(sreg[126]) );
  DFF \sreg_reg[125]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[125]) );
  DFF \sreg_reg[124]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[124]) );
  DFF \sreg_reg[123]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[123]) );
  DFF \sreg_reg[122]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[122]) );
  DFF \sreg_reg[121]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[121]) );
  DFF \sreg_reg[120]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[120]) );
  DFF \sreg_reg[119]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[118]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[117]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[116]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[115]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[114]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[113]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[112]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[111]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[110]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[109]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[108]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[107]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[106]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[105]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[104]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[103]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[102]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[101]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[100]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[99]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[98]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[97]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[96]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[95]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[94]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[93]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[92]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[91]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[90]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[89]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[88]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[87]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[86]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[85]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[84]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[83]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[82]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[81]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[80]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[79]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[78]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[77]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[76]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[75]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[74]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[73]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[72]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[71]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[70]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[69]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[68]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[67]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[66]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[65]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[64]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[63]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[62]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[3]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[2]), .CLK(clk), .RST(rst), .Q(c[0]) );
  NAND U5 ( .A(n1632), .B(n1630), .Z(n1) );
  XOR U6 ( .A(n1632), .B(n1630), .Z(n2) );
  NANDN U7 ( .A(n1631), .B(n2), .Z(n3) );
  NAND U8 ( .A(n1), .B(n3), .Z(n1639) );
  NAND U9 ( .A(n1639), .B(n1637), .Z(n4) );
  XOR U10 ( .A(n1639), .B(n1637), .Z(n5) );
  NANDN U11 ( .A(n1638), .B(n5), .Z(n6) );
  NAND U12 ( .A(n4), .B(n6), .Z(n1647) );
  NAND U13 ( .A(n785), .B(n783), .Z(n7) );
  XOR U14 ( .A(n785), .B(n783), .Z(n8) );
  NANDN U15 ( .A(n784), .B(n8), .Z(n9) );
  NAND U16 ( .A(n7), .B(n9), .Z(n792) );
  NAND U17 ( .A(n806), .B(n804), .Z(n10) );
  XOR U18 ( .A(n806), .B(n804), .Z(n11) );
  NANDN U19 ( .A(n805), .B(n11), .Z(n12) );
  NAND U20 ( .A(n10), .B(n12), .Z(n813) );
  NAND U21 ( .A(n827), .B(n825), .Z(n13) );
  XOR U22 ( .A(n827), .B(n825), .Z(n14) );
  NANDN U23 ( .A(n826), .B(n14), .Z(n15) );
  NAND U24 ( .A(n13), .B(n15), .Z(n834) );
  NAND U25 ( .A(n848), .B(n846), .Z(n16) );
  XOR U26 ( .A(n848), .B(n846), .Z(n17) );
  NANDN U27 ( .A(n847), .B(n17), .Z(n18) );
  NAND U28 ( .A(n16), .B(n18), .Z(n855) );
  NAND U29 ( .A(n869), .B(n867), .Z(n19) );
  XOR U30 ( .A(n869), .B(n867), .Z(n20) );
  NANDN U31 ( .A(n868), .B(n20), .Z(n21) );
  NAND U32 ( .A(n19), .B(n21), .Z(n876) );
  NAND U33 ( .A(n890), .B(n888), .Z(n22) );
  XOR U34 ( .A(n890), .B(n888), .Z(n23) );
  NANDN U35 ( .A(n889), .B(n23), .Z(n24) );
  NAND U36 ( .A(n22), .B(n24), .Z(n897) );
  NAND U37 ( .A(n911), .B(n909), .Z(n25) );
  XOR U38 ( .A(n911), .B(n909), .Z(n26) );
  NANDN U39 ( .A(n910), .B(n26), .Z(n27) );
  NAND U40 ( .A(n25), .B(n27), .Z(n918) );
  NAND U41 ( .A(n932), .B(n930), .Z(n28) );
  XOR U42 ( .A(n932), .B(n930), .Z(n29) );
  NANDN U43 ( .A(n931), .B(n29), .Z(n30) );
  NAND U44 ( .A(n28), .B(n30), .Z(n939) );
  NAND U45 ( .A(n955), .B(n953), .Z(n31) );
  XOR U46 ( .A(n955), .B(n953), .Z(n32) );
  NANDN U47 ( .A(n954), .B(n32), .Z(n33) );
  NAND U48 ( .A(n31), .B(n33), .Z(n960) );
  NAND U49 ( .A(n974), .B(n972), .Z(n34) );
  XOR U50 ( .A(n974), .B(n972), .Z(n35) );
  NANDN U51 ( .A(n973), .B(n35), .Z(n36) );
  NAND U52 ( .A(n34), .B(n36), .Z(n981) );
  NAND U53 ( .A(n995), .B(n993), .Z(n37) );
  XOR U54 ( .A(n995), .B(n993), .Z(n38) );
  NANDN U55 ( .A(n994), .B(n38), .Z(n39) );
  NAND U56 ( .A(n37), .B(n39), .Z(n1002) );
  NAND U57 ( .A(n1016), .B(n1014), .Z(n40) );
  XOR U58 ( .A(n1016), .B(n1014), .Z(n41) );
  NANDN U59 ( .A(n1015), .B(n41), .Z(n42) );
  NAND U60 ( .A(n40), .B(n42), .Z(n1023) );
  NAND U61 ( .A(n1037), .B(n1035), .Z(n43) );
  XOR U62 ( .A(n1037), .B(n1035), .Z(n44) );
  NANDN U63 ( .A(n1036), .B(n44), .Z(n45) );
  NAND U64 ( .A(n43), .B(n45), .Z(n1044) );
  NAND U65 ( .A(n1058), .B(n1056), .Z(n46) );
  XOR U66 ( .A(n1058), .B(n1056), .Z(n47) );
  NANDN U67 ( .A(n1057), .B(n47), .Z(n48) );
  NAND U68 ( .A(n46), .B(n48), .Z(n1065) );
  NAND U69 ( .A(n1079), .B(n1077), .Z(n49) );
  XOR U70 ( .A(n1079), .B(n1077), .Z(n50) );
  NANDN U71 ( .A(n1078), .B(n50), .Z(n51) );
  NAND U72 ( .A(n49), .B(n51), .Z(n1086) );
  NAND U73 ( .A(n1100), .B(n1098), .Z(n52) );
  XOR U74 ( .A(n1100), .B(n1098), .Z(n53) );
  NANDN U75 ( .A(n1099), .B(n53), .Z(n54) );
  NAND U76 ( .A(n52), .B(n54), .Z(n1107) );
  NAND U77 ( .A(n1121), .B(n1119), .Z(n55) );
  XOR U78 ( .A(n1121), .B(n1119), .Z(n56) );
  NANDN U79 ( .A(n1120), .B(n56), .Z(n57) );
  NAND U80 ( .A(n55), .B(n57), .Z(n1128) );
  NAND U81 ( .A(n1142), .B(n1140), .Z(n58) );
  XOR U82 ( .A(n1142), .B(n1140), .Z(n59) );
  NANDN U83 ( .A(n1141), .B(n59), .Z(n60) );
  NAND U84 ( .A(n58), .B(n60), .Z(n1149) );
  NAND U85 ( .A(n1163), .B(n1161), .Z(n61) );
  XOR U86 ( .A(n1163), .B(n1161), .Z(n62) );
  NANDN U87 ( .A(n1162), .B(n62), .Z(n63) );
  NAND U88 ( .A(n61), .B(n63), .Z(n1170) );
  NAND U89 ( .A(n1184), .B(n1182), .Z(n64) );
  XOR U90 ( .A(n1184), .B(n1182), .Z(n65) );
  NANDN U91 ( .A(n1183), .B(n65), .Z(n66) );
  NAND U92 ( .A(n64), .B(n66), .Z(n1191) );
  NAND U93 ( .A(n1205), .B(n1203), .Z(n67) );
  XOR U94 ( .A(n1205), .B(n1203), .Z(n68) );
  NANDN U95 ( .A(n1204), .B(n68), .Z(n69) );
  NAND U96 ( .A(n67), .B(n69), .Z(n1212) );
  NAND U97 ( .A(n1226), .B(n1224), .Z(n70) );
  XOR U98 ( .A(n1226), .B(n1224), .Z(n71) );
  NANDN U99 ( .A(n1225), .B(n71), .Z(n72) );
  NAND U100 ( .A(n70), .B(n72), .Z(n1233) );
  NAND U101 ( .A(n1247), .B(n1245), .Z(n73) );
  XOR U102 ( .A(n1247), .B(n1245), .Z(n74) );
  NANDN U103 ( .A(n1246), .B(n74), .Z(n75) );
  NAND U104 ( .A(n73), .B(n75), .Z(n1254) );
  NAND U105 ( .A(n1268), .B(n1266), .Z(n76) );
  XOR U106 ( .A(n1268), .B(n1266), .Z(n77) );
  NANDN U107 ( .A(n1267), .B(n77), .Z(n78) );
  NAND U108 ( .A(n76), .B(n78), .Z(n1275) );
  NAND U109 ( .A(n1289), .B(n1287), .Z(n79) );
  XOR U110 ( .A(n1289), .B(n1287), .Z(n80) );
  NANDN U111 ( .A(n1288), .B(n80), .Z(n81) );
  NAND U112 ( .A(n79), .B(n81), .Z(n1296) );
  NAND U113 ( .A(n1310), .B(n1308), .Z(n82) );
  XOR U114 ( .A(n1310), .B(n1308), .Z(n83) );
  NANDN U115 ( .A(n1309), .B(n83), .Z(n84) );
  NAND U116 ( .A(n82), .B(n84), .Z(n1317) );
  NAND U117 ( .A(n1331), .B(n1329), .Z(n85) );
  XOR U118 ( .A(n1331), .B(n1329), .Z(n86) );
  NANDN U119 ( .A(n1330), .B(n86), .Z(n87) );
  NAND U120 ( .A(n85), .B(n87), .Z(n1338) );
  NAND U121 ( .A(n1352), .B(n1350), .Z(n88) );
  XOR U122 ( .A(n1352), .B(n1350), .Z(n89) );
  NANDN U123 ( .A(n1351), .B(n89), .Z(n90) );
  NAND U124 ( .A(n88), .B(n90), .Z(n1359) );
  NAND U125 ( .A(n1373), .B(n1371), .Z(n91) );
  XOR U126 ( .A(n1373), .B(n1371), .Z(n92) );
  NANDN U127 ( .A(n1372), .B(n92), .Z(n93) );
  NAND U128 ( .A(n91), .B(n93), .Z(n1380) );
  NAND U129 ( .A(n1394), .B(n1392), .Z(n94) );
  XOR U130 ( .A(n1394), .B(n1392), .Z(n95) );
  NANDN U131 ( .A(n1393), .B(n95), .Z(n96) );
  NAND U132 ( .A(n94), .B(n96), .Z(n1401) );
  NAND U133 ( .A(n1415), .B(n1413), .Z(n97) );
  XOR U134 ( .A(n1415), .B(n1413), .Z(n98) );
  NANDN U135 ( .A(n1414), .B(n98), .Z(n99) );
  NAND U136 ( .A(n97), .B(n99), .Z(n1422) );
  NAND U137 ( .A(n1436), .B(n1434), .Z(n100) );
  XOR U138 ( .A(n1436), .B(n1434), .Z(n101) );
  NANDN U139 ( .A(n1435), .B(n101), .Z(n102) );
  NAND U140 ( .A(n100), .B(n102), .Z(n1443) );
  NAND U141 ( .A(n1457), .B(n1455), .Z(n103) );
  XOR U142 ( .A(n1457), .B(n1455), .Z(n104) );
  NANDN U143 ( .A(n1456), .B(n104), .Z(n105) );
  NAND U144 ( .A(n103), .B(n105), .Z(n1464) );
  NAND U145 ( .A(n1478), .B(n1476), .Z(n106) );
  XOR U146 ( .A(n1478), .B(n1476), .Z(n107) );
  NANDN U147 ( .A(n1477), .B(n107), .Z(n108) );
  NAND U148 ( .A(n106), .B(n108), .Z(n1485) );
  NAND U149 ( .A(n1499), .B(n1497), .Z(n109) );
  XOR U150 ( .A(n1499), .B(n1497), .Z(n110) );
  NANDN U151 ( .A(n1498), .B(n110), .Z(n111) );
  NAND U152 ( .A(n109), .B(n111), .Z(n1506) );
  NAND U153 ( .A(n1520), .B(n1518), .Z(n112) );
  XOR U154 ( .A(n1520), .B(n1518), .Z(n113) );
  NANDN U155 ( .A(n1519), .B(n113), .Z(n114) );
  NAND U156 ( .A(n112), .B(n114), .Z(n1527) );
  NAND U157 ( .A(n1541), .B(n1539), .Z(n115) );
  XOR U158 ( .A(n1541), .B(n1539), .Z(n116) );
  NANDN U159 ( .A(n1540), .B(n116), .Z(n117) );
  NAND U160 ( .A(n115), .B(n117), .Z(n1548) );
  NAND U161 ( .A(n1562), .B(n1560), .Z(n118) );
  XOR U162 ( .A(n1562), .B(n1560), .Z(n119) );
  NANDN U163 ( .A(n1561), .B(n119), .Z(n120) );
  NAND U164 ( .A(n118), .B(n120), .Z(n1569) );
  NAND U165 ( .A(n1583), .B(n1581), .Z(n121) );
  XOR U166 ( .A(n1583), .B(n1581), .Z(n122) );
  NANDN U167 ( .A(n1582), .B(n122), .Z(n123) );
  NAND U168 ( .A(n121), .B(n123), .Z(n1590) );
  NAND U169 ( .A(n1604), .B(n1602), .Z(n124) );
  XOR U170 ( .A(n1604), .B(n1602), .Z(n125) );
  NANDN U171 ( .A(n1603), .B(n125), .Z(n126) );
  NAND U172 ( .A(n124), .B(n126), .Z(n1611) );
  NAND U173 ( .A(n1625), .B(n1623), .Z(n127) );
  XOR U174 ( .A(n1625), .B(n1623), .Z(n128) );
  NANDN U175 ( .A(n1624), .B(n128), .Z(n129) );
  NAND U176 ( .A(n127), .B(n129), .Z(n1632) );
  NAND U177 ( .A(n781), .B(n780), .Z(n130) );
  XOR U178 ( .A(n781), .B(n780), .Z(n131) );
  NANDN U179 ( .A(sreg[129]), .B(n131), .Z(n132) );
  NAND U180 ( .A(n130), .B(n132), .Z(n788) );
  NAND U181 ( .A(n802), .B(n801), .Z(n133) );
  XOR U182 ( .A(n802), .B(n801), .Z(n134) );
  NANDN U183 ( .A(sreg[132]), .B(n134), .Z(n135) );
  NAND U184 ( .A(n133), .B(n135), .Z(n809) );
  NAND U185 ( .A(n823), .B(n822), .Z(n136) );
  XOR U186 ( .A(n823), .B(n822), .Z(n137) );
  NANDN U187 ( .A(sreg[135]), .B(n137), .Z(n138) );
  NAND U188 ( .A(n136), .B(n138), .Z(n830) );
  NAND U189 ( .A(n844), .B(n843), .Z(n139) );
  XOR U190 ( .A(n844), .B(n843), .Z(n140) );
  NANDN U191 ( .A(sreg[138]), .B(n140), .Z(n141) );
  NAND U192 ( .A(n139), .B(n141), .Z(n851) );
  NAND U193 ( .A(n865), .B(n864), .Z(n142) );
  XOR U194 ( .A(n865), .B(n864), .Z(n143) );
  NANDN U195 ( .A(sreg[141]), .B(n143), .Z(n144) );
  NAND U196 ( .A(n142), .B(n144), .Z(n872) );
  NAND U197 ( .A(n886), .B(n885), .Z(n145) );
  XOR U198 ( .A(n886), .B(n885), .Z(n146) );
  NANDN U199 ( .A(sreg[144]), .B(n146), .Z(n147) );
  NAND U200 ( .A(n145), .B(n147), .Z(n893) );
  NAND U201 ( .A(n907), .B(n906), .Z(n148) );
  XOR U202 ( .A(n907), .B(n906), .Z(n149) );
  NANDN U203 ( .A(sreg[147]), .B(n149), .Z(n150) );
  NAND U204 ( .A(n148), .B(n150), .Z(n914) );
  NAND U205 ( .A(n928), .B(n927), .Z(n151) );
  XOR U206 ( .A(n928), .B(n927), .Z(n152) );
  NANDN U207 ( .A(sreg[150]), .B(n152), .Z(n153) );
  NAND U208 ( .A(n151), .B(n153), .Z(n935) );
  NAND U209 ( .A(n949), .B(n948), .Z(n154) );
  XOR U210 ( .A(n949), .B(n948), .Z(n155) );
  NANDN U211 ( .A(sreg[153]), .B(n155), .Z(n156) );
  NAND U212 ( .A(n154), .B(n156), .Z(n952) );
  NAND U213 ( .A(n970), .B(n969), .Z(n157) );
  XOR U214 ( .A(n970), .B(n969), .Z(n158) );
  NANDN U215 ( .A(sreg[156]), .B(n158), .Z(n159) );
  NAND U216 ( .A(n157), .B(n159), .Z(n977) );
  NAND U217 ( .A(n991), .B(n990), .Z(n160) );
  XOR U218 ( .A(n991), .B(n990), .Z(n161) );
  NANDN U219 ( .A(sreg[159]), .B(n161), .Z(n162) );
  NAND U220 ( .A(n160), .B(n162), .Z(n998) );
  NAND U221 ( .A(n1012), .B(n1011), .Z(n163) );
  XOR U222 ( .A(n1012), .B(n1011), .Z(n164) );
  NANDN U223 ( .A(sreg[162]), .B(n164), .Z(n165) );
  NAND U224 ( .A(n163), .B(n165), .Z(n1019) );
  NAND U225 ( .A(n1033), .B(n1032), .Z(n166) );
  XOR U226 ( .A(n1033), .B(n1032), .Z(n167) );
  NANDN U227 ( .A(sreg[165]), .B(n167), .Z(n168) );
  NAND U228 ( .A(n166), .B(n168), .Z(n1040) );
  NAND U229 ( .A(n1054), .B(n1053), .Z(n169) );
  XOR U230 ( .A(n1054), .B(n1053), .Z(n170) );
  NANDN U231 ( .A(sreg[168]), .B(n170), .Z(n171) );
  NAND U232 ( .A(n169), .B(n171), .Z(n1061) );
  NAND U233 ( .A(n1075), .B(n1074), .Z(n172) );
  XOR U234 ( .A(n1075), .B(n1074), .Z(n173) );
  NANDN U235 ( .A(sreg[171]), .B(n173), .Z(n174) );
  NAND U236 ( .A(n172), .B(n174), .Z(n1082) );
  NAND U237 ( .A(n1096), .B(n1095), .Z(n175) );
  XOR U238 ( .A(n1096), .B(n1095), .Z(n176) );
  NANDN U239 ( .A(sreg[174]), .B(n176), .Z(n177) );
  NAND U240 ( .A(n175), .B(n177), .Z(n1103) );
  NAND U241 ( .A(n1117), .B(n1116), .Z(n178) );
  XOR U242 ( .A(n1117), .B(n1116), .Z(n179) );
  NANDN U243 ( .A(sreg[177]), .B(n179), .Z(n180) );
  NAND U244 ( .A(n178), .B(n180), .Z(n1124) );
  NAND U245 ( .A(n1138), .B(n1137), .Z(n181) );
  XOR U246 ( .A(n1138), .B(n1137), .Z(n182) );
  NANDN U247 ( .A(sreg[180]), .B(n182), .Z(n183) );
  NAND U248 ( .A(n181), .B(n183), .Z(n1145) );
  NAND U249 ( .A(n1159), .B(n1158), .Z(n184) );
  XOR U250 ( .A(n1159), .B(n1158), .Z(n185) );
  NANDN U251 ( .A(sreg[183]), .B(n185), .Z(n186) );
  NAND U252 ( .A(n184), .B(n186), .Z(n1166) );
  NAND U253 ( .A(n1180), .B(n1179), .Z(n187) );
  XOR U254 ( .A(n1180), .B(n1179), .Z(n188) );
  NANDN U255 ( .A(sreg[186]), .B(n188), .Z(n189) );
  NAND U256 ( .A(n187), .B(n189), .Z(n1187) );
  NAND U257 ( .A(n1201), .B(n1200), .Z(n190) );
  XOR U258 ( .A(n1201), .B(n1200), .Z(n191) );
  NANDN U259 ( .A(sreg[189]), .B(n191), .Z(n192) );
  NAND U260 ( .A(n190), .B(n192), .Z(n1208) );
  NAND U261 ( .A(n1222), .B(n1221), .Z(n193) );
  XOR U262 ( .A(n1222), .B(n1221), .Z(n194) );
  NANDN U263 ( .A(sreg[192]), .B(n194), .Z(n195) );
  NAND U264 ( .A(n193), .B(n195), .Z(n1229) );
  NAND U265 ( .A(n1243), .B(n1242), .Z(n196) );
  XOR U266 ( .A(n1243), .B(n1242), .Z(n197) );
  NANDN U267 ( .A(sreg[195]), .B(n197), .Z(n198) );
  NAND U268 ( .A(n196), .B(n198), .Z(n1250) );
  NAND U269 ( .A(n1264), .B(n1263), .Z(n199) );
  XOR U270 ( .A(n1264), .B(n1263), .Z(n200) );
  NANDN U271 ( .A(sreg[198]), .B(n200), .Z(n201) );
  NAND U272 ( .A(n199), .B(n201), .Z(n1271) );
  NAND U273 ( .A(n1285), .B(n1284), .Z(n202) );
  XOR U274 ( .A(n1285), .B(n1284), .Z(n203) );
  NANDN U275 ( .A(sreg[201]), .B(n203), .Z(n204) );
  NAND U276 ( .A(n202), .B(n204), .Z(n1292) );
  NAND U277 ( .A(n1306), .B(n1305), .Z(n205) );
  XOR U278 ( .A(n1306), .B(n1305), .Z(n206) );
  NANDN U279 ( .A(sreg[204]), .B(n206), .Z(n207) );
  NAND U280 ( .A(n205), .B(n207), .Z(n1313) );
  NAND U281 ( .A(n1327), .B(n1326), .Z(n208) );
  XOR U282 ( .A(n1327), .B(n1326), .Z(n209) );
  NANDN U283 ( .A(sreg[207]), .B(n209), .Z(n210) );
  NAND U284 ( .A(n208), .B(n210), .Z(n1334) );
  NAND U285 ( .A(n1348), .B(n1347), .Z(n211) );
  XOR U286 ( .A(n1348), .B(n1347), .Z(n212) );
  NANDN U287 ( .A(sreg[210]), .B(n212), .Z(n213) );
  NAND U288 ( .A(n211), .B(n213), .Z(n1355) );
  NAND U289 ( .A(n1369), .B(n1368), .Z(n214) );
  XOR U290 ( .A(n1369), .B(n1368), .Z(n215) );
  NANDN U291 ( .A(sreg[213]), .B(n215), .Z(n216) );
  NAND U292 ( .A(n214), .B(n216), .Z(n1376) );
  NAND U293 ( .A(n1390), .B(n1389), .Z(n217) );
  XOR U294 ( .A(n1390), .B(n1389), .Z(n218) );
  NANDN U295 ( .A(sreg[216]), .B(n218), .Z(n219) );
  NAND U296 ( .A(n217), .B(n219), .Z(n1397) );
  NAND U297 ( .A(n1411), .B(n1410), .Z(n220) );
  XOR U298 ( .A(n1411), .B(n1410), .Z(n221) );
  NANDN U299 ( .A(sreg[219]), .B(n221), .Z(n222) );
  NAND U300 ( .A(n220), .B(n222), .Z(n1418) );
  NAND U301 ( .A(n1432), .B(n1431), .Z(n223) );
  XOR U302 ( .A(n1432), .B(n1431), .Z(n224) );
  NANDN U303 ( .A(sreg[222]), .B(n224), .Z(n225) );
  NAND U304 ( .A(n223), .B(n225), .Z(n1439) );
  NAND U305 ( .A(n1453), .B(n1452), .Z(n226) );
  XOR U306 ( .A(n1453), .B(n1452), .Z(n227) );
  NANDN U307 ( .A(sreg[225]), .B(n227), .Z(n228) );
  NAND U308 ( .A(n226), .B(n228), .Z(n1460) );
  NAND U309 ( .A(n1474), .B(n1473), .Z(n229) );
  XOR U310 ( .A(n1474), .B(n1473), .Z(n230) );
  NANDN U311 ( .A(sreg[228]), .B(n230), .Z(n231) );
  NAND U312 ( .A(n229), .B(n231), .Z(n1481) );
  NAND U313 ( .A(n1495), .B(n1494), .Z(n232) );
  XOR U314 ( .A(n1495), .B(n1494), .Z(n233) );
  NANDN U315 ( .A(sreg[231]), .B(n233), .Z(n234) );
  NAND U316 ( .A(n232), .B(n234), .Z(n1502) );
  NAND U317 ( .A(n1516), .B(n1515), .Z(n235) );
  XOR U318 ( .A(n1516), .B(n1515), .Z(n236) );
  NANDN U319 ( .A(sreg[234]), .B(n236), .Z(n237) );
  NAND U320 ( .A(n235), .B(n237), .Z(n1523) );
  NAND U321 ( .A(n1537), .B(n1536), .Z(n238) );
  XOR U322 ( .A(n1537), .B(n1536), .Z(n239) );
  NANDN U323 ( .A(sreg[237]), .B(n239), .Z(n240) );
  NAND U324 ( .A(n238), .B(n240), .Z(n1544) );
  NAND U325 ( .A(n1558), .B(n1557), .Z(n241) );
  XOR U326 ( .A(n1558), .B(n1557), .Z(n242) );
  NANDN U327 ( .A(sreg[240]), .B(n242), .Z(n243) );
  NAND U328 ( .A(n241), .B(n243), .Z(n1565) );
  NAND U329 ( .A(n1579), .B(n1578), .Z(n244) );
  XOR U330 ( .A(n1579), .B(n1578), .Z(n245) );
  NANDN U331 ( .A(sreg[243]), .B(n245), .Z(n246) );
  NAND U332 ( .A(n244), .B(n246), .Z(n1586) );
  NAND U333 ( .A(n1600), .B(n1599), .Z(n247) );
  XOR U334 ( .A(n1600), .B(n1599), .Z(n248) );
  NANDN U335 ( .A(sreg[246]), .B(n248), .Z(n249) );
  NAND U336 ( .A(n247), .B(n249), .Z(n1607) );
  NAND U337 ( .A(n1621), .B(n1620), .Z(n250) );
  XOR U338 ( .A(n1621), .B(n1620), .Z(n251) );
  NANDN U339 ( .A(sreg[249]), .B(n251), .Z(n252) );
  NAND U340 ( .A(n250), .B(n252), .Z(n1628) );
  NAND U341 ( .A(n1641), .B(n1640), .Z(n253) );
  XOR U342 ( .A(n1641), .B(n1640), .Z(n254) );
  NANDN U343 ( .A(sreg[252]), .B(n254), .Z(n255) );
  NAND U344 ( .A(n253), .B(n255), .Z(n1644) );
  NAND U345 ( .A(n792), .B(n790), .Z(n256) );
  XOR U346 ( .A(n792), .B(n790), .Z(n257) );
  NANDN U347 ( .A(n791), .B(n257), .Z(n258) );
  NAND U348 ( .A(n256), .B(n258), .Z(n799) );
  NAND U349 ( .A(n813), .B(n811), .Z(n259) );
  XOR U350 ( .A(n813), .B(n811), .Z(n260) );
  NANDN U351 ( .A(n812), .B(n260), .Z(n261) );
  NAND U352 ( .A(n259), .B(n261), .Z(n820) );
  NAND U353 ( .A(n834), .B(n832), .Z(n262) );
  XOR U354 ( .A(n834), .B(n832), .Z(n263) );
  NANDN U355 ( .A(n833), .B(n263), .Z(n264) );
  NAND U356 ( .A(n262), .B(n264), .Z(n841) );
  NAND U357 ( .A(n855), .B(n853), .Z(n265) );
  XOR U358 ( .A(n855), .B(n853), .Z(n266) );
  NANDN U359 ( .A(n854), .B(n266), .Z(n267) );
  NAND U360 ( .A(n265), .B(n267), .Z(n862) );
  NAND U361 ( .A(n876), .B(n874), .Z(n268) );
  XOR U362 ( .A(n876), .B(n874), .Z(n269) );
  NANDN U363 ( .A(n875), .B(n269), .Z(n270) );
  NAND U364 ( .A(n268), .B(n270), .Z(n883) );
  NAND U365 ( .A(n897), .B(n895), .Z(n271) );
  XOR U366 ( .A(n897), .B(n895), .Z(n272) );
  NANDN U367 ( .A(n896), .B(n272), .Z(n273) );
  NAND U368 ( .A(n271), .B(n273), .Z(n904) );
  NAND U369 ( .A(n918), .B(n916), .Z(n274) );
  XOR U370 ( .A(n918), .B(n916), .Z(n275) );
  NANDN U371 ( .A(n917), .B(n275), .Z(n276) );
  NAND U372 ( .A(n274), .B(n276), .Z(n925) );
  NAND U373 ( .A(n939), .B(n937), .Z(n277) );
  XOR U374 ( .A(n939), .B(n937), .Z(n278) );
  NANDN U375 ( .A(n938), .B(n278), .Z(n279) );
  NAND U376 ( .A(n277), .B(n279), .Z(n946) );
  NAND U377 ( .A(n960), .B(n958), .Z(n280) );
  XOR U378 ( .A(n960), .B(n958), .Z(n281) );
  NANDN U379 ( .A(n959), .B(n281), .Z(n282) );
  NAND U380 ( .A(n280), .B(n282), .Z(n967) );
  NAND U381 ( .A(n981), .B(n979), .Z(n283) );
  XOR U382 ( .A(n981), .B(n979), .Z(n284) );
  NANDN U383 ( .A(n980), .B(n284), .Z(n285) );
  NAND U384 ( .A(n283), .B(n285), .Z(n988) );
  NAND U385 ( .A(n1002), .B(n1000), .Z(n286) );
  XOR U386 ( .A(n1002), .B(n1000), .Z(n287) );
  NANDN U387 ( .A(n1001), .B(n287), .Z(n288) );
  NAND U388 ( .A(n286), .B(n288), .Z(n1009) );
  NAND U389 ( .A(n1023), .B(n1021), .Z(n289) );
  XOR U390 ( .A(n1023), .B(n1021), .Z(n290) );
  NANDN U391 ( .A(n1022), .B(n290), .Z(n291) );
  NAND U392 ( .A(n289), .B(n291), .Z(n1030) );
  NAND U393 ( .A(n1044), .B(n1042), .Z(n292) );
  XOR U394 ( .A(n1044), .B(n1042), .Z(n293) );
  NANDN U395 ( .A(n1043), .B(n293), .Z(n294) );
  NAND U396 ( .A(n292), .B(n294), .Z(n1051) );
  NAND U397 ( .A(n1065), .B(n1063), .Z(n295) );
  XOR U398 ( .A(n1065), .B(n1063), .Z(n296) );
  NANDN U399 ( .A(n1064), .B(n296), .Z(n297) );
  NAND U400 ( .A(n295), .B(n297), .Z(n1072) );
  NAND U401 ( .A(n1086), .B(n1084), .Z(n298) );
  XOR U402 ( .A(n1086), .B(n1084), .Z(n299) );
  NANDN U403 ( .A(n1085), .B(n299), .Z(n300) );
  NAND U404 ( .A(n298), .B(n300), .Z(n1093) );
  NAND U405 ( .A(n1107), .B(n1105), .Z(n301) );
  XOR U406 ( .A(n1107), .B(n1105), .Z(n302) );
  NANDN U407 ( .A(n1106), .B(n302), .Z(n303) );
  NAND U408 ( .A(n301), .B(n303), .Z(n1114) );
  NAND U409 ( .A(n1128), .B(n1126), .Z(n304) );
  XOR U410 ( .A(n1128), .B(n1126), .Z(n305) );
  NANDN U411 ( .A(n1127), .B(n305), .Z(n306) );
  NAND U412 ( .A(n304), .B(n306), .Z(n1135) );
  NAND U413 ( .A(n1149), .B(n1147), .Z(n307) );
  XOR U414 ( .A(n1149), .B(n1147), .Z(n308) );
  NANDN U415 ( .A(n1148), .B(n308), .Z(n309) );
  NAND U416 ( .A(n307), .B(n309), .Z(n1156) );
  NAND U417 ( .A(n1170), .B(n1168), .Z(n310) );
  XOR U418 ( .A(n1170), .B(n1168), .Z(n311) );
  NANDN U419 ( .A(n1169), .B(n311), .Z(n312) );
  NAND U420 ( .A(n310), .B(n312), .Z(n1177) );
  NAND U421 ( .A(n1191), .B(n1189), .Z(n313) );
  XOR U422 ( .A(n1191), .B(n1189), .Z(n314) );
  NANDN U423 ( .A(n1190), .B(n314), .Z(n315) );
  NAND U424 ( .A(n313), .B(n315), .Z(n1198) );
  NAND U425 ( .A(n1212), .B(n1210), .Z(n316) );
  XOR U426 ( .A(n1212), .B(n1210), .Z(n317) );
  NANDN U427 ( .A(n1211), .B(n317), .Z(n318) );
  NAND U428 ( .A(n316), .B(n318), .Z(n1219) );
  NAND U429 ( .A(n1233), .B(n1231), .Z(n319) );
  XOR U430 ( .A(n1233), .B(n1231), .Z(n320) );
  NANDN U431 ( .A(n1232), .B(n320), .Z(n321) );
  NAND U432 ( .A(n319), .B(n321), .Z(n1240) );
  NAND U433 ( .A(n1254), .B(n1252), .Z(n322) );
  XOR U434 ( .A(n1254), .B(n1252), .Z(n323) );
  NANDN U435 ( .A(n1253), .B(n323), .Z(n324) );
  NAND U436 ( .A(n322), .B(n324), .Z(n1261) );
  NAND U437 ( .A(n1275), .B(n1273), .Z(n325) );
  XOR U438 ( .A(n1275), .B(n1273), .Z(n326) );
  NANDN U439 ( .A(n1274), .B(n326), .Z(n327) );
  NAND U440 ( .A(n325), .B(n327), .Z(n1282) );
  NAND U441 ( .A(n1296), .B(n1294), .Z(n328) );
  XOR U442 ( .A(n1296), .B(n1294), .Z(n329) );
  NANDN U443 ( .A(n1295), .B(n329), .Z(n330) );
  NAND U444 ( .A(n328), .B(n330), .Z(n1303) );
  NAND U445 ( .A(n1317), .B(n1315), .Z(n331) );
  XOR U446 ( .A(n1317), .B(n1315), .Z(n332) );
  NANDN U447 ( .A(n1316), .B(n332), .Z(n333) );
  NAND U448 ( .A(n331), .B(n333), .Z(n1324) );
  NAND U449 ( .A(n1338), .B(n1336), .Z(n334) );
  XOR U450 ( .A(n1338), .B(n1336), .Z(n335) );
  NANDN U451 ( .A(n1337), .B(n335), .Z(n336) );
  NAND U452 ( .A(n334), .B(n336), .Z(n1345) );
  NAND U453 ( .A(n1359), .B(n1357), .Z(n337) );
  XOR U454 ( .A(n1359), .B(n1357), .Z(n338) );
  NANDN U455 ( .A(n1358), .B(n338), .Z(n339) );
  NAND U456 ( .A(n337), .B(n339), .Z(n1366) );
  NAND U457 ( .A(n1380), .B(n1378), .Z(n340) );
  XOR U458 ( .A(n1380), .B(n1378), .Z(n341) );
  NANDN U459 ( .A(n1379), .B(n341), .Z(n342) );
  NAND U460 ( .A(n340), .B(n342), .Z(n1387) );
  NAND U461 ( .A(n1401), .B(n1399), .Z(n343) );
  XOR U462 ( .A(n1401), .B(n1399), .Z(n344) );
  NANDN U463 ( .A(n1400), .B(n344), .Z(n345) );
  NAND U464 ( .A(n343), .B(n345), .Z(n1408) );
  NAND U465 ( .A(n1422), .B(n1420), .Z(n346) );
  XOR U466 ( .A(n1422), .B(n1420), .Z(n347) );
  NANDN U467 ( .A(n1421), .B(n347), .Z(n348) );
  NAND U468 ( .A(n346), .B(n348), .Z(n1429) );
  NAND U469 ( .A(n1443), .B(n1441), .Z(n349) );
  XOR U470 ( .A(n1443), .B(n1441), .Z(n350) );
  NANDN U471 ( .A(n1442), .B(n350), .Z(n351) );
  NAND U472 ( .A(n349), .B(n351), .Z(n1450) );
  NAND U473 ( .A(n1464), .B(n1462), .Z(n352) );
  XOR U474 ( .A(n1464), .B(n1462), .Z(n353) );
  NANDN U475 ( .A(n1463), .B(n353), .Z(n354) );
  NAND U476 ( .A(n352), .B(n354), .Z(n1471) );
  NAND U477 ( .A(n1485), .B(n1483), .Z(n355) );
  XOR U478 ( .A(n1485), .B(n1483), .Z(n356) );
  NANDN U479 ( .A(n1484), .B(n356), .Z(n357) );
  NAND U480 ( .A(n355), .B(n357), .Z(n1492) );
  NAND U481 ( .A(n1506), .B(n1504), .Z(n358) );
  XOR U482 ( .A(n1506), .B(n1504), .Z(n359) );
  NANDN U483 ( .A(n1505), .B(n359), .Z(n360) );
  NAND U484 ( .A(n358), .B(n360), .Z(n1513) );
  NAND U485 ( .A(n1527), .B(n1525), .Z(n361) );
  XOR U486 ( .A(n1527), .B(n1525), .Z(n362) );
  NANDN U487 ( .A(n1526), .B(n362), .Z(n363) );
  NAND U488 ( .A(n361), .B(n363), .Z(n1534) );
  NAND U489 ( .A(n1548), .B(n1546), .Z(n364) );
  XOR U490 ( .A(n1548), .B(n1546), .Z(n365) );
  NANDN U491 ( .A(n1547), .B(n365), .Z(n366) );
  NAND U492 ( .A(n364), .B(n366), .Z(n1555) );
  NAND U493 ( .A(n1569), .B(n1567), .Z(n367) );
  XOR U494 ( .A(n1569), .B(n1567), .Z(n368) );
  NANDN U495 ( .A(n1568), .B(n368), .Z(n369) );
  NAND U496 ( .A(n367), .B(n369), .Z(n1576) );
  NAND U497 ( .A(n1590), .B(n1588), .Z(n370) );
  XOR U498 ( .A(n1590), .B(n1588), .Z(n371) );
  NANDN U499 ( .A(n1589), .B(n371), .Z(n372) );
  NAND U500 ( .A(n370), .B(n372), .Z(n1597) );
  NAND U501 ( .A(n1611), .B(n1609), .Z(n373) );
  XOR U502 ( .A(n1611), .B(n1609), .Z(n374) );
  NANDN U503 ( .A(n1610), .B(n374), .Z(n375) );
  NAND U504 ( .A(n373), .B(n375), .Z(n1618) );
  NAND U505 ( .A(n788), .B(n787), .Z(n376) );
  XOR U506 ( .A(n788), .B(n787), .Z(n377) );
  NANDN U507 ( .A(sreg[130]), .B(n377), .Z(n378) );
  NAND U508 ( .A(n376), .B(n378), .Z(n795) );
  NAND U509 ( .A(n809), .B(n808), .Z(n379) );
  XOR U510 ( .A(n809), .B(n808), .Z(n380) );
  NANDN U511 ( .A(sreg[133]), .B(n380), .Z(n381) );
  NAND U512 ( .A(n379), .B(n381), .Z(n816) );
  NAND U513 ( .A(n830), .B(n829), .Z(n382) );
  XOR U514 ( .A(n830), .B(n829), .Z(n383) );
  NANDN U515 ( .A(sreg[136]), .B(n383), .Z(n384) );
  NAND U516 ( .A(n382), .B(n384), .Z(n837) );
  NAND U517 ( .A(n851), .B(n850), .Z(n385) );
  XOR U518 ( .A(n851), .B(n850), .Z(n386) );
  NANDN U519 ( .A(sreg[139]), .B(n386), .Z(n387) );
  NAND U520 ( .A(n385), .B(n387), .Z(n858) );
  NAND U521 ( .A(n872), .B(n871), .Z(n388) );
  XOR U522 ( .A(n872), .B(n871), .Z(n389) );
  NANDN U523 ( .A(sreg[142]), .B(n389), .Z(n390) );
  NAND U524 ( .A(n388), .B(n390), .Z(n879) );
  NAND U525 ( .A(n893), .B(n892), .Z(n391) );
  XOR U526 ( .A(n893), .B(n892), .Z(n392) );
  NANDN U527 ( .A(sreg[145]), .B(n392), .Z(n393) );
  NAND U528 ( .A(n391), .B(n393), .Z(n900) );
  NAND U529 ( .A(n914), .B(n913), .Z(n394) );
  XOR U530 ( .A(n914), .B(n913), .Z(n395) );
  NANDN U531 ( .A(sreg[148]), .B(n395), .Z(n396) );
  NAND U532 ( .A(n394), .B(n396), .Z(n921) );
  NAND U533 ( .A(n935), .B(n934), .Z(n397) );
  XOR U534 ( .A(n935), .B(n934), .Z(n398) );
  NANDN U535 ( .A(sreg[151]), .B(n398), .Z(n399) );
  NAND U536 ( .A(n397), .B(n399), .Z(n942) );
  NAND U537 ( .A(n952), .B(n951), .Z(n400) );
  XOR U538 ( .A(n952), .B(n951), .Z(n401) );
  NANDN U539 ( .A(sreg[154]), .B(n401), .Z(n402) );
  NAND U540 ( .A(n400), .B(n402), .Z(n962) );
  NAND U541 ( .A(n977), .B(n976), .Z(n403) );
  XOR U542 ( .A(n977), .B(n976), .Z(n404) );
  NANDN U543 ( .A(sreg[157]), .B(n404), .Z(n405) );
  NAND U544 ( .A(n403), .B(n405), .Z(n984) );
  NAND U545 ( .A(n998), .B(n997), .Z(n406) );
  XOR U546 ( .A(n998), .B(n997), .Z(n407) );
  NANDN U547 ( .A(sreg[160]), .B(n407), .Z(n408) );
  NAND U548 ( .A(n406), .B(n408), .Z(n1005) );
  NAND U549 ( .A(n1019), .B(n1018), .Z(n409) );
  XOR U550 ( .A(n1019), .B(n1018), .Z(n410) );
  NANDN U551 ( .A(sreg[163]), .B(n410), .Z(n411) );
  NAND U552 ( .A(n409), .B(n411), .Z(n1026) );
  NAND U553 ( .A(n1040), .B(n1039), .Z(n412) );
  XOR U554 ( .A(n1040), .B(n1039), .Z(n413) );
  NANDN U555 ( .A(sreg[166]), .B(n413), .Z(n414) );
  NAND U556 ( .A(n412), .B(n414), .Z(n1047) );
  NAND U557 ( .A(n1061), .B(n1060), .Z(n415) );
  XOR U558 ( .A(n1061), .B(n1060), .Z(n416) );
  NANDN U559 ( .A(sreg[169]), .B(n416), .Z(n417) );
  NAND U560 ( .A(n415), .B(n417), .Z(n1068) );
  NAND U561 ( .A(n1082), .B(n1081), .Z(n418) );
  XOR U562 ( .A(n1082), .B(n1081), .Z(n419) );
  NANDN U563 ( .A(sreg[172]), .B(n419), .Z(n420) );
  NAND U564 ( .A(n418), .B(n420), .Z(n1089) );
  NAND U565 ( .A(n1103), .B(n1102), .Z(n421) );
  XOR U566 ( .A(n1103), .B(n1102), .Z(n422) );
  NANDN U567 ( .A(sreg[175]), .B(n422), .Z(n423) );
  NAND U568 ( .A(n421), .B(n423), .Z(n1110) );
  NAND U569 ( .A(n1124), .B(n1123), .Z(n424) );
  XOR U570 ( .A(n1124), .B(n1123), .Z(n425) );
  NANDN U571 ( .A(sreg[178]), .B(n425), .Z(n426) );
  NAND U572 ( .A(n424), .B(n426), .Z(n1131) );
  NAND U573 ( .A(n1145), .B(n1144), .Z(n427) );
  XOR U574 ( .A(n1145), .B(n1144), .Z(n428) );
  NANDN U575 ( .A(sreg[181]), .B(n428), .Z(n429) );
  NAND U576 ( .A(n427), .B(n429), .Z(n1152) );
  NAND U577 ( .A(n1166), .B(n1165), .Z(n430) );
  XOR U578 ( .A(n1166), .B(n1165), .Z(n431) );
  NANDN U579 ( .A(sreg[184]), .B(n431), .Z(n432) );
  NAND U580 ( .A(n430), .B(n432), .Z(n1173) );
  NAND U581 ( .A(n1187), .B(n1186), .Z(n433) );
  XOR U582 ( .A(n1187), .B(n1186), .Z(n434) );
  NANDN U583 ( .A(sreg[187]), .B(n434), .Z(n435) );
  NAND U584 ( .A(n433), .B(n435), .Z(n1194) );
  NAND U585 ( .A(n1208), .B(n1207), .Z(n436) );
  XOR U586 ( .A(n1208), .B(n1207), .Z(n437) );
  NANDN U587 ( .A(sreg[190]), .B(n437), .Z(n438) );
  NAND U588 ( .A(n436), .B(n438), .Z(n1215) );
  NAND U589 ( .A(n1229), .B(n1228), .Z(n439) );
  XOR U590 ( .A(n1229), .B(n1228), .Z(n440) );
  NANDN U591 ( .A(sreg[193]), .B(n440), .Z(n441) );
  NAND U592 ( .A(n439), .B(n441), .Z(n1236) );
  NAND U593 ( .A(n1250), .B(n1249), .Z(n442) );
  XOR U594 ( .A(n1250), .B(n1249), .Z(n443) );
  NANDN U595 ( .A(sreg[196]), .B(n443), .Z(n444) );
  NAND U596 ( .A(n442), .B(n444), .Z(n1257) );
  NAND U597 ( .A(n1271), .B(n1270), .Z(n445) );
  XOR U598 ( .A(n1271), .B(n1270), .Z(n446) );
  NANDN U599 ( .A(sreg[199]), .B(n446), .Z(n447) );
  NAND U600 ( .A(n445), .B(n447), .Z(n1278) );
  NAND U601 ( .A(n1292), .B(n1291), .Z(n448) );
  XOR U602 ( .A(n1292), .B(n1291), .Z(n449) );
  NANDN U603 ( .A(sreg[202]), .B(n449), .Z(n450) );
  NAND U604 ( .A(n448), .B(n450), .Z(n1299) );
  NAND U605 ( .A(n1313), .B(n1312), .Z(n451) );
  XOR U606 ( .A(n1313), .B(n1312), .Z(n452) );
  NANDN U607 ( .A(sreg[205]), .B(n452), .Z(n453) );
  NAND U608 ( .A(n451), .B(n453), .Z(n1320) );
  NAND U609 ( .A(n1334), .B(n1333), .Z(n454) );
  XOR U610 ( .A(n1334), .B(n1333), .Z(n455) );
  NANDN U611 ( .A(sreg[208]), .B(n455), .Z(n456) );
  NAND U612 ( .A(n454), .B(n456), .Z(n1341) );
  NAND U613 ( .A(n1355), .B(n1354), .Z(n457) );
  XOR U614 ( .A(n1355), .B(n1354), .Z(n458) );
  NANDN U615 ( .A(sreg[211]), .B(n458), .Z(n459) );
  NAND U616 ( .A(n457), .B(n459), .Z(n1362) );
  NAND U617 ( .A(n1376), .B(n1375), .Z(n460) );
  XOR U618 ( .A(n1376), .B(n1375), .Z(n461) );
  NANDN U619 ( .A(sreg[214]), .B(n461), .Z(n462) );
  NAND U620 ( .A(n460), .B(n462), .Z(n1383) );
  NAND U621 ( .A(n1397), .B(n1396), .Z(n463) );
  XOR U622 ( .A(n1397), .B(n1396), .Z(n464) );
  NANDN U623 ( .A(sreg[217]), .B(n464), .Z(n465) );
  NAND U624 ( .A(n463), .B(n465), .Z(n1404) );
  NAND U625 ( .A(n1418), .B(n1417), .Z(n466) );
  XOR U626 ( .A(n1418), .B(n1417), .Z(n467) );
  NANDN U627 ( .A(sreg[220]), .B(n467), .Z(n468) );
  NAND U628 ( .A(n466), .B(n468), .Z(n1425) );
  NAND U629 ( .A(n1439), .B(n1438), .Z(n469) );
  XOR U630 ( .A(n1439), .B(n1438), .Z(n470) );
  NANDN U631 ( .A(sreg[223]), .B(n470), .Z(n471) );
  NAND U632 ( .A(n469), .B(n471), .Z(n1446) );
  NAND U633 ( .A(n1460), .B(n1459), .Z(n472) );
  XOR U634 ( .A(n1460), .B(n1459), .Z(n473) );
  NANDN U635 ( .A(sreg[226]), .B(n473), .Z(n474) );
  NAND U636 ( .A(n472), .B(n474), .Z(n1467) );
  NAND U637 ( .A(n1481), .B(n1480), .Z(n475) );
  XOR U638 ( .A(n1481), .B(n1480), .Z(n476) );
  NANDN U639 ( .A(sreg[229]), .B(n476), .Z(n477) );
  NAND U640 ( .A(n475), .B(n477), .Z(n1488) );
  NAND U641 ( .A(n1502), .B(n1501), .Z(n478) );
  XOR U642 ( .A(n1502), .B(n1501), .Z(n479) );
  NANDN U643 ( .A(sreg[232]), .B(n479), .Z(n480) );
  NAND U644 ( .A(n478), .B(n480), .Z(n1509) );
  NAND U645 ( .A(n1523), .B(n1522), .Z(n481) );
  XOR U646 ( .A(n1523), .B(n1522), .Z(n482) );
  NANDN U647 ( .A(sreg[235]), .B(n482), .Z(n483) );
  NAND U648 ( .A(n481), .B(n483), .Z(n1530) );
  NAND U649 ( .A(n1544), .B(n1543), .Z(n484) );
  XOR U650 ( .A(n1544), .B(n1543), .Z(n485) );
  NANDN U651 ( .A(sreg[238]), .B(n485), .Z(n486) );
  NAND U652 ( .A(n484), .B(n486), .Z(n1551) );
  NAND U653 ( .A(n1565), .B(n1564), .Z(n487) );
  XOR U654 ( .A(n1565), .B(n1564), .Z(n488) );
  NANDN U655 ( .A(sreg[241]), .B(n488), .Z(n489) );
  NAND U656 ( .A(n487), .B(n489), .Z(n1572) );
  NAND U657 ( .A(n1586), .B(n1585), .Z(n490) );
  XOR U658 ( .A(n1586), .B(n1585), .Z(n491) );
  NANDN U659 ( .A(sreg[244]), .B(n491), .Z(n492) );
  NAND U660 ( .A(n490), .B(n492), .Z(n1593) );
  NAND U661 ( .A(n1607), .B(n1606), .Z(n493) );
  XOR U662 ( .A(n1607), .B(n1606), .Z(n494) );
  NANDN U663 ( .A(sreg[247]), .B(n494), .Z(n495) );
  NAND U664 ( .A(n493), .B(n495), .Z(n1614) );
  NAND U665 ( .A(n1628), .B(n1627), .Z(n496) );
  XOR U666 ( .A(n1628), .B(n1627), .Z(n497) );
  NANDN U667 ( .A(sreg[250]), .B(n497), .Z(n498) );
  NAND U668 ( .A(n496), .B(n498), .Z(n1635) );
  NAND U669 ( .A(n1644), .B(n1643), .Z(n499) );
  XOR U670 ( .A(n1644), .B(n1643), .Z(n500) );
  NANDN U671 ( .A(sreg[253]), .B(n500), .Z(n501) );
  NAND U672 ( .A(n499), .B(n501), .Z(n1653) );
  OR U673 ( .A(n776), .B(n778), .Z(n502) );
  NANDN U674 ( .A(n777), .B(n502), .Z(n503) );
  NANDN U675 ( .A(n778), .B(n777), .Z(n504) );
  NAND U676 ( .A(n775), .B(n504), .Z(n505) );
  NAND U677 ( .A(n503), .B(n505), .Z(n785) );
  NAND U678 ( .A(n799), .B(n797), .Z(n506) );
  XOR U679 ( .A(n799), .B(n797), .Z(n507) );
  NANDN U680 ( .A(n798), .B(n507), .Z(n508) );
  NAND U681 ( .A(n506), .B(n508), .Z(n806) );
  NAND U682 ( .A(n820), .B(n818), .Z(n509) );
  XOR U683 ( .A(n820), .B(n818), .Z(n510) );
  NANDN U684 ( .A(n819), .B(n510), .Z(n511) );
  NAND U685 ( .A(n509), .B(n511), .Z(n827) );
  NAND U686 ( .A(n841), .B(n839), .Z(n512) );
  XOR U687 ( .A(n841), .B(n839), .Z(n513) );
  NANDN U688 ( .A(n840), .B(n513), .Z(n514) );
  NAND U689 ( .A(n512), .B(n514), .Z(n848) );
  NAND U690 ( .A(n862), .B(n860), .Z(n515) );
  XOR U691 ( .A(n862), .B(n860), .Z(n516) );
  NANDN U692 ( .A(n861), .B(n516), .Z(n517) );
  NAND U693 ( .A(n515), .B(n517), .Z(n869) );
  NAND U694 ( .A(n883), .B(n881), .Z(n518) );
  XOR U695 ( .A(n883), .B(n881), .Z(n519) );
  NANDN U696 ( .A(n882), .B(n519), .Z(n520) );
  NAND U697 ( .A(n518), .B(n520), .Z(n890) );
  NAND U698 ( .A(n904), .B(n902), .Z(n521) );
  XOR U699 ( .A(n904), .B(n902), .Z(n522) );
  NANDN U700 ( .A(n903), .B(n522), .Z(n523) );
  NAND U701 ( .A(n521), .B(n523), .Z(n911) );
  NAND U702 ( .A(n925), .B(n923), .Z(n524) );
  XOR U703 ( .A(n925), .B(n923), .Z(n525) );
  NANDN U704 ( .A(n924), .B(n525), .Z(n526) );
  NAND U705 ( .A(n524), .B(n526), .Z(n932) );
  NAND U706 ( .A(n946), .B(n944), .Z(n527) );
  XOR U707 ( .A(n946), .B(n944), .Z(n528) );
  NANDN U708 ( .A(n945), .B(n528), .Z(n529) );
  NAND U709 ( .A(n527), .B(n529), .Z(n955) );
  NAND U710 ( .A(n967), .B(n965), .Z(n530) );
  XOR U711 ( .A(n967), .B(n965), .Z(n531) );
  NANDN U712 ( .A(n966), .B(n531), .Z(n532) );
  NAND U713 ( .A(n530), .B(n532), .Z(n974) );
  NAND U714 ( .A(n988), .B(n986), .Z(n533) );
  XOR U715 ( .A(n988), .B(n986), .Z(n534) );
  NANDN U716 ( .A(n987), .B(n534), .Z(n535) );
  NAND U717 ( .A(n533), .B(n535), .Z(n995) );
  NAND U718 ( .A(n1009), .B(n1007), .Z(n536) );
  XOR U719 ( .A(n1009), .B(n1007), .Z(n537) );
  NANDN U720 ( .A(n1008), .B(n537), .Z(n538) );
  NAND U721 ( .A(n536), .B(n538), .Z(n1016) );
  NAND U722 ( .A(n1030), .B(n1028), .Z(n539) );
  XOR U723 ( .A(n1030), .B(n1028), .Z(n540) );
  NANDN U724 ( .A(n1029), .B(n540), .Z(n541) );
  NAND U725 ( .A(n539), .B(n541), .Z(n1037) );
  NAND U726 ( .A(n1051), .B(n1049), .Z(n542) );
  XOR U727 ( .A(n1051), .B(n1049), .Z(n543) );
  NANDN U728 ( .A(n1050), .B(n543), .Z(n544) );
  NAND U729 ( .A(n542), .B(n544), .Z(n1058) );
  NAND U730 ( .A(n1072), .B(n1070), .Z(n545) );
  XOR U731 ( .A(n1072), .B(n1070), .Z(n546) );
  NANDN U732 ( .A(n1071), .B(n546), .Z(n547) );
  NAND U733 ( .A(n545), .B(n547), .Z(n1079) );
  NAND U734 ( .A(n1093), .B(n1091), .Z(n548) );
  XOR U735 ( .A(n1093), .B(n1091), .Z(n549) );
  NANDN U736 ( .A(n1092), .B(n549), .Z(n550) );
  NAND U737 ( .A(n548), .B(n550), .Z(n1100) );
  NAND U738 ( .A(n1114), .B(n1112), .Z(n551) );
  XOR U739 ( .A(n1114), .B(n1112), .Z(n552) );
  NANDN U740 ( .A(n1113), .B(n552), .Z(n553) );
  NAND U741 ( .A(n551), .B(n553), .Z(n1121) );
  NAND U742 ( .A(n1135), .B(n1133), .Z(n554) );
  XOR U743 ( .A(n1135), .B(n1133), .Z(n555) );
  NANDN U744 ( .A(n1134), .B(n555), .Z(n556) );
  NAND U745 ( .A(n554), .B(n556), .Z(n1142) );
  NAND U746 ( .A(n1156), .B(n1154), .Z(n557) );
  XOR U747 ( .A(n1156), .B(n1154), .Z(n558) );
  NANDN U748 ( .A(n1155), .B(n558), .Z(n559) );
  NAND U749 ( .A(n557), .B(n559), .Z(n1163) );
  NAND U750 ( .A(n1177), .B(n1175), .Z(n560) );
  XOR U751 ( .A(n1177), .B(n1175), .Z(n561) );
  NANDN U752 ( .A(n1176), .B(n561), .Z(n562) );
  NAND U753 ( .A(n560), .B(n562), .Z(n1184) );
  NAND U754 ( .A(n1198), .B(n1196), .Z(n563) );
  XOR U755 ( .A(n1198), .B(n1196), .Z(n564) );
  NANDN U756 ( .A(n1197), .B(n564), .Z(n565) );
  NAND U757 ( .A(n563), .B(n565), .Z(n1205) );
  NAND U758 ( .A(n1219), .B(n1217), .Z(n566) );
  XOR U759 ( .A(n1219), .B(n1217), .Z(n567) );
  NANDN U760 ( .A(n1218), .B(n567), .Z(n568) );
  NAND U761 ( .A(n566), .B(n568), .Z(n1226) );
  NAND U762 ( .A(n1240), .B(n1238), .Z(n569) );
  XOR U763 ( .A(n1240), .B(n1238), .Z(n570) );
  NANDN U764 ( .A(n1239), .B(n570), .Z(n571) );
  NAND U765 ( .A(n569), .B(n571), .Z(n1247) );
  NAND U766 ( .A(n1261), .B(n1259), .Z(n572) );
  XOR U767 ( .A(n1261), .B(n1259), .Z(n573) );
  NANDN U768 ( .A(n1260), .B(n573), .Z(n574) );
  NAND U769 ( .A(n572), .B(n574), .Z(n1268) );
  NAND U770 ( .A(n1282), .B(n1280), .Z(n575) );
  XOR U771 ( .A(n1282), .B(n1280), .Z(n576) );
  NANDN U772 ( .A(n1281), .B(n576), .Z(n577) );
  NAND U773 ( .A(n575), .B(n577), .Z(n1289) );
  NAND U774 ( .A(n1303), .B(n1301), .Z(n578) );
  XOR U775 ( .A(n1303), .B(n1301), .Z(n579) );
  NANDN U776 ( .A(n1302), .B(n579), .Z(n580) );
  NAND U777 ( .A(n578), .B(n580), .Z(n1310) );
  NAND U778 ( .A(n1324), .B(n1322), .Z(n581) );
  XOR U779 ( .A(n1324), .B(n1322), .Z(n582) );
  NANDN U780 ( .A(n1323), .B(n582), .Z(n583) );
  NAND U781 ( .A(n581), .B(n583), .Z(n1331) );
  NAND U782 ( .A(n1345), .B(n1343), .Z(n584) );
  XOR U783 ( .A(n1345), .B(n1343), .Z(n585) );
  NANDN U784 ( .A(n1344), .B(n585), .Z(n586) );
  NAND U785 ( .A(n584), .B(n586), .Z(n1352) );
  NAND U786 ( .A(n1366), .B(n1364), .Z(n587) );
  XOR U787 ( .A(n1366), .B(n1364), .Z(n588) );
  NANDN U788 ( .A(n1365), .B(n588), .Z(n589) );
  NAND U789 ( .A(n587), .B(n589), .Z(n1373) );
  NAND U790 ( .A(n1387), .B(n1385), .Z(n590) );
  XOR U791 ( .A(n1387), .B(n1385), .Z(n591) );
  NANDN U792 ( .A(n1386), .B(n591), .Z(n592) );
  NAND U793 ( .A(n590), .B(n592), .Z(n1394) );
  NAND U794 ( .A(n1408), .B(n1406), .Z(n593) );
  XOR U795 ( .A(n1408), .B(n1406), .Z(n594) );
  NANDN U796 ( .A(n1407), .B(n594), .Z(n595) );
  NAND U797 ( .A(n593), .B(n595), .Z(n1415) );
  NAND U798 ( .A(n1429), .B(n1427), .Z(n596) );
  XOR U799 ( .A(n1429), .B(n1427), .Z(n597) );
  NANDN U800 ( .A(n1428), .B(n597), .Z(n598) );
  NAND U801 ( .A(n596), .B(n598), .Z(n1436) );
  NAND U802 ( .A(n1450), .B(n1448), .Z(n599) );
  XOR U803 ( .A(n1450), .B(n1448), .Z(n600) );
  NANDN U804 ( .A(n1449), .B(n600), .Z(n601) );
  NAND U805 ( .A(n599), .B(n601), .Z(n1457) );
  NAND U806 ( .A(n1471), .B(n1469), .Z(n602) );
  XOR U807 ( .A(n1471), .B(n1469), .Z(n603) );
  NANDN U808 ( .A(n1470), .B(n603), .Z(n604) );
  NAND U809 ( .A(n602), .B(n604), .Z(n1478) );
  NAND U810 ( .A(n1492), .B(n1490), .Z(n605) );
  XOR U811 ( .A(n1492), .B(n1490), .Z(n606) );
  NANDN U812 ( .A(n1491), .B(n606), .Z(n607) );
  NAND U813 ( .A(n605), .B(n607), .Z(n1499) );
  NAND U814 ( .A(n1513), .B(n1511), .Z(n608) );
  XOR U815 ( .A(n1513), .B(n1511), .Z(n609) );
  NANDN U816 ( .A(n1512), .B(n609), .Z(n610) );
  NAND U817 ( .A(n608), .B(n610), .Z(n1520) );
  NAND U818 ( .A(n1534), .B(n1532), .Z(n611) );
  XOR U819 ( .A(n1534), .B(n1532), .Z(n612) );
  NANDN U820 ( .A(n1533), .B(n612), .Z(n613) );
  NAND U821 ( .A(n611), .B(n613), .Z(n1541) );
  NAND U822 ( .A(n1555), .B(n1553), .Z(n614) );
  XOR U823 ( .A(n1555), .B(n1553), .Z(n615) );
  NANDN U824 ( .A(n1554), .B(n615), .Z(n616) );
  NAND U825 ( .A(n614), .B(n616), .Z(n1562) );
  NAND U826 ( .A(n1576), .B(n1574), .Z(n617) );
  XOR U827 ( .A(n1576), .B(n1574), .Z(n618) );
  NANDN U828 ( .A(n1575), .B(n618), .Z(n619) );
  NAND U829 ( .A(n617), .B(n619), .Z(n1583) );
  NAND U830 ( .A(n1597), .B(n1595), .Z(n620) );
  XOR U831 ( .A(n1597), .B(n1595), .Z(n621) );
  NANDN U832 ( .A(n1596), .B(n621), .Z(n622) );
  NAND U833 ( .A(n620), .B(n622), .Z(n1604) );
  NAND U834 ( .A(n1618), .B(n1616), .Z(n623) );
  XOR U835 ( .A(n1618), .B(n1616), .Z(n624) );
  NANDN U836 ( .A(n1617), .B(n624), .Z(n625) );
  NAND U837 ( .A(n623), .B(n625), .Z(n1625) );
  NAND U838 ( .A(n795), .B(n794), .Z(n626) );
  XOR U839 ( .A(n795), .B(n794), .Z(n627) );
  NANDN U840 ( .A(sreg[131]), .B(n627), .Z(n628) );
  NAND U841 ( .A(n626), .B(n628), .Z(n802) );
  NAND U842 ( .A(n816), .B(n815), .Z(n629) );
  XOR U843 ( .A(n816), .B(n815), .Z(n630) );
  NANDN U844 ( .A(sreg[134]), .B(n630), .Z(n631) );
  NAND U845 ( .A(n629), .B(n631), .Z(n823) );
  NAND U846 ( .A(n837), .B(n836), .Z(n632) );
  XOR U847 ( .A(n837), .B(n836), .Z(n633) );
  NANDN U848 ( .A(sreg[137]), .B(n633), .Z(n634) );
  NAND U849 ( .A(n632), .B(n634), .Z(n844) );
  NAND U850 ( .A(n858), .B(n857), .Z(n635) );
  XOR U851 ( .A(n858), .B(n857), .Z(n636) );
  NANDN U852 ( .A(sreg[140]), .B(n636), .Z(n637) );
  NAND U853 ( .A(n635), .B(n637), .Z(n865) );
  NAND U854 ( .A(n879), .B(n878), .Z(n638) );
  XOR U855 ( .A(n879), .B(n878), .Z(n639) );
  NANDN U856 ( .A(sreg[143]), .B(n639), .Z(n640) );
  NAND U857 ( .A(n638), .B(n640), .Z(n886) );
  NAND U858 ( .A(n900), .B(n899), .Z(n641) );
  XOR U859 ( .A(n900), .B(n899), .Z(n642) );
  NANDN U860 ( .A(sreg[146]), .B(n642), .Z(n643) );
  NAND U861 ( .A(n641), .B(n643), .Z(n907) );
  NAND U862 ( .A(n921), .B(n920), .Z(n644) );
  XOR U863 ( .A(n921), .B(n920), .Z(n645) );
  NANDN U864 ( .A(sreg[149]), .B(n645), .Z(n646) );
  NAND U865 ( .A(n644), .B(n646), .Z(n928) );
  NAND U866 ( .A(n942), .B(n941), .Z(n647) );
  XOR U867 ( .A(n942), .B(n941), .Z(n648) );
  NANDN U868 ( .A(sreg[152]), .B(n648), .Z(n649) );
  NAND U869 ( .A(n647), .B(n649), .Z(n949) );
  XOR U870 ( .A(n963), .B(sreg[155]), .Z(n650) );
  NANDN U871 ( .A(n962), .B(n650), .Z(n651) );
  NAND U872 ( .A(n963), .B(sreg[155]), .Z(n652) );
  AND U873 ( .A(n651), .B(n652), .Z(n970) );
  NAND U874 ( .A(n984), .B(n983), .Z(n653) );
  XOR U875 ( .A(n984), .B(n983), .Z(n654) );
  NANDN U876 ( .A(sreg[158]), .B(n654), .Z(n655) );
  NAND U877 ( .A(n653), .B(n655), .Z(n991) );
  NAND U878 ( .A(n1005), .B(n1004), .Z(n656) );
  XOR U879 ( .A(n1005), .B(n1004), .Z(n657) );
  NANDN U880 ( .A(sreg[161]), .B(n657), .Z(n658) );
  NAND U881 ( .A(n656), .B(n658), .Z(n1012) );
  NAND U882 ( .A(n1026), .B(n1025), .Z(n659) );
  XOR U883 ( .A(n1026), .B(n1025), .Z(n660) );
  NANDN U884 ( .A(sreg[164]), .B(n660), .Z(n661) );
  NAND U885 ( .A(n659), .B(n661), .Z(n1033) );
  NAND U886 ( .A(n1047), .B(n1046), .Z(n662) );
  XOR U887 ( .A(n1047), .B(n1046), .Z(n663) );
  NANDN U888 ( .A(sreg[167]), .B(n663), .Z(n664) );
  NAND U889 ( .A(n662), .B(n664), .Z(n1054) );
  NAND U890 ( .A(n1068), .B(n1067), .Z(n665) );
  XOR U891 ( .A(n1068), .B(n1067), .Z(n666) );
  NANDN U892 ( .A(sreg[170]), .B(n666), .Z(n667) );
  NAND U893 ( .A(n665), .B(n667), .Z(n1075) );
  NAND U894 ( .A(n1089), .B(n1088), .Z(n668) );
  XOR U895 ( .A(n1089), .B(n1088), .Z(n669) );
  NANDN U896 ( .A(sreg[173]), .B(n669), .Z(n670) );
  NAND U897 ( .A(n668), .B(n670), .Z(n1096) );
  NAND U898 ( .A(n1110), .B(n1109), .Z(n671) );
  XOR U899 ( .A(n1110), .B(n1109), .Z(n672) );
  NANDN U900 ( .A(sreg[176]), .B(n672), .Z(n673) );
  NAND U901 ( .A(n671), .B(n673), .Z(n1117) );
  NAND U902 ( .A(n1131), .B(n1130), .Z(n674) );
  XOR U903 ( .A(n1131), .B(n1130), .Z(n675) );
  NANDN U904 ( .A(sreg[179]), .B(n675), .Z(n676) );
  NAND U905 ( .A(n674), .B(n676), .Z(n1138) );
  NAND U906 ( .A(n1152), .B(n1151), .Z(n677) );
  XOR U907 ( .A(n1152), .B(n1151), .Z(n678) );
  NANDN U908 ( .A(sreg[182]), .B(n678), .Z(n679) );
  NAND U909 ( .A(n677), .B(n679), .Z(n1159) );
  NAND U910 ( .A(n1173), .B(n1172), .Z(n680) );
  XOR U911 ( .A(n1173), .B(n1172), .Z(n681) );
  NANDN U912 ( .A(sreg[185]), .B(n681), .Z(n682) );
  NAND U913 ( .A(n680), .B(n682), .Z(n1180) );
  NAND U914 ( .A(n1194), .B(n1193), .Z(n683) );
  XOR U915 ( .A(n1194), .B(n1193), .Z(n684) );
  NANDN U916 ( .A(sreg[188]), .B(n684), .Z(n685) );
  NAND U917 ( .A(n683), .B(n685), .Z(n1201) );
  NAND U918 ( .A(n1215), .B(n1214), .Z(n686) );
  XOR U919 ( .A(n1215), .B(n1214), .Z(n687) );
  NANDN U920 ( .A(sreg[191]), .B(n687), .Z(n688) );
  NAND U921 ( .A(n686), .B(n688), .Z(n1222) );
  NAND U922 ( .A(n1236), .B(n1235), .Z(n689) );
  XOR U923 ( .A(n1236), .B(n1235), .Z(n690) );
  NANDN U924 ( .A(sreg[194]), .B(n690), .Z(n691) );
  NAND U925 ( .A(n689), .B(n691), .Z(n1243) );
  NAND U926 ( .A(n1257), .B(n1256), .Z(n692) );
  XOR U927 ( .A(n1257), .B(n1256), .Z(n693) );
  NANDN U928 ( .A(sreg[197]), .B(n693), .Z(n694) );
  NAND U929 ( .A(n692), .B(n694), .Z(n1264) );
  NAND U930 ( .A(n1278), .B(n1277), .Z(n695) );
  XOR U931 ( .A(n1278), .B(n1277), .Z(n696) );
  NANDN U932 ( .A(sreg[200]), .B(n696), .Z(n697) );
  NAND U933 ( .A(n695), .B(n697), .Z(n1285) );
  NAND U934 ( .A(n1299), .B(n1298), .Z(n698) );
  XOR U935 ( .A(n1299), .B(n1298), .Z(n699) );
  NANDN U936 ( .A(sreg[203]), .B(n699), .Z(n700) );
  NAND U937 ( .A(n698), .B(n700), .Z(n1306) );
  NAND U938 ( .A(n1320), .B(n1319), .Z(n701) );
  XOR U939 ( .A(n1320), .B(n1319), .Z(n702) );
  NANDN U940 ( .A(sreg[206]), .B(n702), .Z(n703) );
  NAND U941 ( .A(n701), .B(n703), .Z(n1327) );
  NAND U942 ( .A(n1341), .B(n1340), .Z(n704) );
  XOR U943 ( .A(n1341), .B(n1340), .Z(n705) );
  NANDN U944 ( .A(sreg[209]), .B(n705), .Z(n706) );
  NAND U945 ( .A(n704), .B(n706), .Z(n1348) );
  NAND U946 ( .A(n1362), .B(n1361), .Z(n707) );
  XOR U947 ( .A(n1362), .B(n1361), .Z(n708) );
  NANDN U948 ( .A(sreg[212]), .B(n708), .Z(n709) );
  NAND U949 ( .A(n707), .B(n709), .Z(n1369) );
  NAND U950 ( .A(n1383), .B(n1382), .Z(n710) );
  XOR U951 ( .A(n1383), .B(n1382), .Z(n711) );
  NANDN U952 ( .A(sreg[215]), .B(n711), .Z(n712) );
  NAND U953 ( .A(n710), .B(n712), .Z(n1390) );
  NAND U954 ( .A(n1404), .B(n1403), .Z(n713) );
  XOR U955 ( .A(n1404), .B(n1403), .Z(n714) );
  NANDN U956 ( .A(sreg[218]), .B(n714), .Z(n715) );
  NAND U957 ( .A(n713), .B(n715), .Z(n1411) );
  NAND U958 ( .A(n1425), .B(n1424), .Z(n716) );
  XOR U959 ( .A(n1425), .B(n1424), .Z(n717) );
  NANDN U960 ( .A(sreg[221]), .B(n717), .Z(n718) );
  NAND U961 ( .A(n716), .B(n718), .Z(n1432) );
  NAND U962 ( .A(n1446), .B(n1445), .Z(n719) );
  XOR U963 ( .A(n1446), .B(n1445), .Z(n720) );
  NANDN U964 ( .A(sreg[224]), .B(n720), .Z(n721) );
  NAND U965 ( .A(n719), .B(n721), .Z(n1453) );
  NAND U966 ( .A(n1467), .B(n1466), .Z(n722) );
  XOR U967 ( .A(n1467), .B(n1466), .Z(n723) );
  NANDN U968 ( .A(sreg[227]), .B(n723), .Z(n724) );
  NAND U969 ( .A(n722), .B(n724), .Z(n1474) );
  NAND U970 ( .A(n1488), .B(n1487), .Z(n725) );
  XOR U971 ( .A(n1488), .B(n1487), .Z(n726) );
  NANDN U972 ( .A(sreg[230]), .B(n726), .Z(n727) );
  NAND U973 ( .A(n725), .B(n727), .Z(n1495) );
  NAND U974 ( .A(n1509), .B(n1508), .Z(n728) );
  XOR U975 ( .A(n1509), .B(n1508), .Z(n729) );
  NANDN U976 ( .A(sreg[233]), .B(n729), .Z(n730) );
  NAND U977 ( .A(n728), .B(n730), .Z(n1516) );
  NAND U978 ( .A(n1530), .B(n1529), .Z(n731) );
  XOR U979 ( .A(n1530), .B(n1529), .Z(n732) );
  NANDN U980 ( .A(sreg[236]), .B(n732), .Z(n733) );
  NAND U981 ( .A(n731), .B(n733), .Z(n1537) );
  NAND U982 ( .A(n1551), .B(n1550), .Z(n734) );
  XOR U983 ( .A(n1551), .B(n1550), .Z(n735) );
  NANDN U984 ( .A(sreg[239]), .B(n735), .Z(n736) );
  NAND U985 ( .A(n734), .B(n736), .Z(n1558) );
  NAND U986 ( .A(n1572), .B(n1571), .Z(n737) );
  XOR U987 ( .A(n1572), .B(n1571), .Z(n738) );
  NANDN U988 ( .A(sreg[242]), .B(n738), .Z(n739) );
  NAND U989 ( .A(n737), .B(n739), .Z(n1579) );
  NAND U990 ( .A(n1593), .B(n1592), .Z(n740) );
  XOR U991 ( .A(n1593), .B(n1592), .Z(n741) );
  NANDN U992 ( .A(sreg[245]), .B(n741), .Z(n742) );
  NAND U993 ( .A(n740), .B(n742), .Z(n1600) );
  NAND U994 ( .A(n1614), .B(n1613), .Z(n743) );
  XOR U995 ( .A(n1614), .B(n1613), .Z(n744) );
  NANDN U996 ( .A(sreg[248]), .B(n744), .Z(n745) );
  NAND U997 ( .A(n743), .B(n745), .Z(n1621) );
  NAND U998 ( .A(n1635), .B(n1634), .Z(n746) );
  XOR U999 ( .A(n1635), .B(n1634), .Z(n747) );
  NANDN U1000 ( .A(sreg[251]), .B(n747), .Z(n748) );
  NAND U1001 ( .A(n746), .B(n748), .Z(n1641) );
  XOR U1002 ( .A(n1654), .B(n1653), .Z(n749) );
  NANDN U1003 ( .A(n1652), .B(n749), .Z(n750) );
  NAND U1004 ( .A(n1653), .B(n1654), .Z(n751) );
  AND U1005 ( .A(n750), .B(n751), .Z(c[255]) );
  AND U1006 ( .A(b[0]), .B(a[0]), .Z(n752) );
  XOR U1007 ( .A(n752), .B(sreg[126]), .Z(c[126]) );
  AND U1008 ( .A(b[0]), .B(a[1]), .Z(n776) );
  NAND U1009 ( .A(b[1]), .B(a[0]), .Z(n764) );
  XOR U1010 ( .A(n776), .B(n764), .Z(n759) );
  AND U1011 ( .A(n752), .B(sreg[126]), .Z(n758) );
  IV U1012 ( .A(n758), .Z(n757) );
  XNOR U1013 ( .A(sreg[127]), .B(n757), .Z(n753) );
  XNOR U1014 ( .A(n759), .B(n753), .Z(c[127]) );
  ANDN U1015 ( .B(n776), .A(n764), .Z(n778) );
  AND U1016 ( .A(a[2]), .B(b[0]), .Z(n755) );
  NAND U1017 ( .A(a[1]), .B(b[1]), .Z(n754) );
  XNOR U1018 ( .A(n755), .B(n754), .Z(n756) );
  XNOR U1019 ( .A(n778), .B(n756), .Z(n770) );
  IV U1020 ( .A(n770), .Z(n768) );
  NANDN U1021 ( .A(sreg[127]), .B(n757), .Z(n762) );
  AND U1022 ( .A(sreg[127]), .B(n758), .Z(n760) );
  NANDN U1023 ( .A(n760), .B(n759), .Z(n761) );
  AND U1024 ( .A(n762), .B(n761), .Z(n769) );
  XNOR U1025 ( .A(n768), .B(n769), .Z(n763) );
  XNOR U1026 ( .A(sreg[128]), .B(n763), .Z(c[128]) );
  AND U1027 ( .A(b[0]), .B(a[3]), .Z(n775) );
  NAND U1028 ( .A(b[1]), .B(a[2]), .Z(n777) );
  XNOR U1029 ( .A(n776), .B(n777), .Z(n766) );
  NAND U1030 ( .A(n776), .B(n764), .Z(n765) );
  NAND U1031 ( .A(n766), .B(n765), .Z(n767) );
  XOR U1032 ( .A(n775), .B(n767), .Z(n780) );
  NAND U1033 ( .A(n768), .B(n769), .Z(n773) );
  ANDN U1034 ( .B(n770), .A(n769), .Z(n771) );
  NANDN U1035 ( .A(n771), .B(sreg[128]), .Z(n772) );
  AND U1036 ( .A(n773), .B(n772), .Z(n781) );
  XNOR U1037 ( .A(n781), .B(sreg[129]), .Z(n774) );
  XNOR U1038 ( .A(n780), .B(n774), .Z(c[129]) );
  NAND U1039 ( .A(b[0]), .B(a[4]), .Z(n784) );
  AND U1040 ( .A(b[1]), .B(a[3]), .Z(n783) );
  XNOR U1041 ( .A(n785), .B(n783), .Z(n779) );
  XNOR U1042 ( .A(n784), .B(n779), .Z(n787) );
  XNOR U1043 ( .A(n788), .B(sreg[130]), .Z(n782) );
  XNOR U1044 ( .A(n787), .B(n782), .Z(c[130]) );
  NAND U1045 ( .A(b[0]), .B(a[5]), .Z(n791) );
  AND U1046 ( .A(b[1]), .B(a[4]), .Z(n790) );
  XNOR U1047 ( .A(n792), .B(n790), .Z(n786) );
  XNOR U1048 ( .A(n791), .B(n786), .Z(n794) );
  XNOR U1049 ( .A(n795), .B(sreg[131]), .Z(n789) );
  XNOR U1050 ( .A(n794), .B(n789), .Z(c[131]) );
  NAND U1051 ( .A(b[0]), .B(a[6]), .Z(n798) );
  AND U1052 ( .A(b[1]), .B(a[5]), .Z(n797) );
  XNOR U1053 ( .A(n799), .B(n797), .Z(n793) );
  XNOR U1054 ( .A(n798), .B(n793), .Z(n801) );
  XNOR U1055 ( .A(n802), .B(sreg[132]), .Z(n796) );
  XNOR U1056 ( .A(n801), .B(n796), .Z(c[132]) );
  NAND U1057 ( .A(b[0]), .B(a[7]), .Z(n805) );
  AND U1058 ( .A(b[1]), .B(a[6]), .Z(n804) );
  XNOR U1059 ( .A(n806), .B(n804), .Z(n800) );
  XNOR U1060 ( .A(n805), .B(n800), .Z(n808) );
  XNOR U1061 ( .A(n809), .B(sreg[133]), .Z(n803) );
  XNOR U1062 ( .A(n808), .B(n803), .Z(c[133]) );
  NAND U1063 ( .A(b[0]), .B(a[8]), .Z(n812) );
  AND U1064 ( .A(b[1]), .B(a[7]), .Z(n811) );
  XNOR U1065 ( .A(n813), .B(n811), .Z(n807) );
  XNOR U1066 ( .A(n812), .B(n807), .Z(n815) );
  XNOR U1067 ( .A(n816), .B(sreg[134]), .Z(n810) );
  XNOR U1068 ( .A(n815), .B(n810), .Z(c[134]) );
  NAND U1069 ( .A(b[0]), .B(a[9]), .Z(n819) );
  AND U1070 ( .A(b[1]), .B(a[8]), .Z(n818) );
  XNOR U1071 ( .A(n820), .B(n818), .Z(n814) );
  XNOR U1072 ( .A(n819), .B(n814), .Z(n822) );
  XNOR U1073 ( .A(n823), .B(sreg[135]), .Z(n817) );
  XNOR U1074 ( .A(n822), .B(n817), .Z(c[135]) );
  NAND U1075 ( .A(b[0]), .B(a[10]), .Z(n826) );
  AND U1076 ( .A(b[1]), .B(a[9]), .Z(n825) );
  XNOR U1077 ( .A(n827), .B(n825), .Z(n821) );
  XNOR U1078 ( .A(n826), .B(n821), .Z(n829) );
  XNOR U1079 ( .A(n830), .B(sreg[136]), .Z(n824) );
  XNOR U1080 ( .A(n829), .B(n824), .Z(c[136]) );
  NAND U1081 ( .A(b[0]), .B(a[11]), .Z(n833) );
  AND U1082 ( .A(b[1]), .B(a[10]), .Z(n832) );
  XNOR U1083 ( .A(n834), .B(n832), .Z(n828) );
  XNOR U1084 ( .A(n833), .B(n828), .Z(n836) );
  XNOR U1085 ( .A(n837), .B(sreg[137]), .Z(n831) );
  XNOR U1086 ( .A(n836), .B(n831), .Z(c[137]) );
  NAND U1087 ( .A(b[0]), .B(a[12]), .Z(n840) );
  AND U1088 ( .A(b[1]), .B(a[11]), .Z(n839) );
  XNOR U1089 ( .A(n841), .B(n839), .Z(n835) );
  XNOR U1090 ( .A(n840), .B(n835), .Z(n843) );
  XNOR U1091 ( .A(n844), .B(sreg[138]), .Z(n838) );
  XNOR U1092 ( .A(n843), .B(n838), .Z(c[138]) );
  NAND U1093 ( .A(b[0]), .B(a[13]), .Z(n847) );
  AND U1094 ( .A(b[1]), .B(a[12]), .Z(n846) );
  XNOR U1095 ( .A(n848), .B(n846), .Z(n842) );
  XNOR U1096 ( .A(n847), .B(n842), .Z(n850) );
  XNOR U1097 ( .A(n851), .B(sreg[139]), .Z(n845) );
  XNOR U1098 ( .A(n850), .B(n845), .Z(c[139]) );
  NAND U1099 ( .A(b[0]), .B(a[14]), .Z(n854) );
  AND U1100 ( .A(b[1]), .B(a[13]), .Z(n853) );
  XNOR U1101 ( .A(n855), .B(n853), .Z(n849) );
  XNOR U1102 ( .A(n854), .B(n849), .Z(n857) );
  XNOR U1103 ( .A(n858), .B(sreg[140]), .Z(n852) );
  XNOR U1104 ( .A(n857), .B(n852), .Z(c[140]) );
  NAND U1105 ( .A(b[0]), .B(a[15]), .Z(n861) );
  AND U1106 ( .A(b[1]), .B(a[14]), .Z(n860) );
  XNOR U1107 ( .A(n862), .B(n860), .Z(n856) );
  XNOR U1108 ( .A(n861), .B(n856), .Z(n864) );
  XNOR U1109 ( .A(n865), .B(sreg[141]), .Z(n859) );
  XNOR U1110 ( .A(n864), .B(n859), .Z(c[141]) );
  NAND U1111 ( .A(b[0]), .B(a[16]), .Z(n868) );
  AND U1112 ( .A(b[1]), .B(a[15]), .Z(n867) );
  XNOR U1113 ( .A(n869), .B(n867), .Z(n863) );
  XNOR U1114 ( .A(n868), .B(n863), .Z(n871) );
  XNOR U1115 ( .A(n872), .B(sreg[142]), .Z(n866) );
  XNOR U1116 ( .A(n871), .B(n866), .Z(c[142]) );
  NAND U1117 ( .A(b[0]), .B(a[17]), .Z(n875) );
  AND U1118 ( .A(b[1]), .B(a[16]), .Z(n874) );
  XNOR U1119 ( .A(n876), .B(n874), .Z(n870) );
  XNOR U1120 ( .A(n875), .B(n870), .Z(n878) );
  XNOR U1121 ( .A(n879), .B(sreg[143]), .Z(n873) );
  XNOR U1122 ( .A(n878), .B(n873), .Z(c[143]) );
  NAND U1123 ( .A(b[0]), .B(a[18]), .Z(n882) );
  AND U1124 ( .A(b[1]), .B(a[17]), .Z(n881) );
  XNOR U1125 ( .A(n883), .B(n881), .Z(n877) );
  XNOR U1126 ( .A(n882), .B(n877), .Z(n885) );
  XNOR U1127 ( .A(n886), .B(sreg[144]), .Z(n880) );
  XNOR U1128 ( .A(n885), .B(n880), .Z(c[144]) );
  NAND U1129 ( .A(b[0]), .B(a[19]), .Z(n889) );
  AND U1130 ( .A(b[1]), .B(a[18]), .Z(n888) );
  XNOR U1131 ( .A(n890), .B(n888), .Z(n884) );
  XNOR U1132 ( .A(n889), .B(n884), .Z(n892) );
  XNOR U1133 ( .A(n893), .B(sreg[145]), .Z(n887) );
  XNOR U1134 ( .A(n892), .B(n887), .Z(c[145]) );
  NAND U1135 ( .A(b[0]), .B(a[20]), .Z(n896) );
  AND U1136 ( .A(b[1]), .B(a[19]), .Z(n895) );
  XNOR U1137 ( .A(n897), .B(n895), .Z(n891) );
  XNOR U1138 ( .A(n896), .B(n891), .Z(n899) );
  XNOR U1139 ( .A(n900), .B(sreg[146]), .Z(n894) );
  XNOR U1140 ( .A(n899), .B(n894), .Z(c[146]) );
  NAND U1141 ( .A(b[0]), .B(a[21]), .Z(n903) );
  AND U1142 ( .A(b[1]), .B(a[20]), .Z(n902) );
  XNOR U1143 ( .A(n904), .B(n902), .Z(n898) );
  XNOR U1144 ( .A(n903), .B(n898), .Z(n906) );
  XNOR U1145 ( .A(n907), .B(sreg[147]), .Z(n901) );
  XNOR U1146 ( .A(n906), .B(n901), .Z(c[147]) );
  NAND U1147 ( .A(b[0]), .B(a[22]), .Z(n910) );
  AND U1148 ( .A(b[1]), .B(a[21]), .Z(n909) );
  XNOR U1149 ( .A(n911), .B(n909), .Z(n905) );
  XNOR U1150 ( .A(n910), .B(n905), .Z(n913) );
  XNOR U1151 ( .A(n914), .B(sreg[148]), .Z(n908) );
  XNOR U1152 ( .A(n913), .B(n908), .Z(c[148]) );
  NAND U1153 ( .A(b[0]), .B(a[23]), .Z(n917) );
  AND U1154 ( .A(b[1]), .B(a[22]), .Z(n916) );
  XNOR U1155 ( .A(n918), .B(n916), .Z(n912) );
  XNOR U1156 ( .A(n917), .B(n912), .Z(n920) );
  XNOR U1157 ( .A(n921), .B(sreg[149]), .Z(n915) );
  XNOR U1158 ( .A(n920), .B(n915), .Z(c[149]) );
  NAND U1159 ( .A(b[0]), .B(a[24]), .Z(n924) );
  AND U1160 ( .A(b[1]), .B(a[23]), .Z(n923) );
  XNOR U1161 ( .A(n925), .B(n923), .Z(n919) );
  XNOR U1162 ( .A(n924), .B(n919), .Z(n927) );
  XNOR U1163 ( .A(n928), .B(sreg[150]), .Z(n922) );
  XNOR U1164 ( .A(n927), .B(n922), .Z(c[150]) );
  NAND U1165 ( .A(b[0]), .B(a[25]), .Z(n931) );
  AND U1166 ( .A(b[1]), .B(a[24]), .Z(n930) );
  XNOR U1167 ( .A(n932), .B(n930), .Z(n926) );
  XNOR U1168 ( .A(n931), .B(n926), .Z(n934) );
  XNOR U1169 ( .A(n935), .B(sreg[151]), .Z(n929) );
  XNOR U1170 ( .A(n934), .B(n929), .Z(c[151]) );
  NAND U1171 ( .A(b[0]), .B(a[26]), .Z(n938) );
  AND U1172 ( .A(b[1]), .B(a[25]), .Z(n937) );
  XNOR U1173 ( .A(n939), .B(n937), .Z(n933) );
  XNOR U1174 ( .A(n938), .B(n933), .Z(n941) );
  XNOR U1175 ( .A(n942), .B(sreg[152]), .Z(n936) );
  XNOR U1176 ( .A(n941), .B(n936), .Z(c[152]) );
  NAND U1177 ( .A(b[0]), .B(a[27]), .Z(n945) );
  AND U1178 ( .A(b[1]), .B(a[26]), .Z(n944) );
  XNOR U1179 ( .A(n946), .B(n944), .Z(n940) );
  XNOR U1180 ( .A(n945), .B(n940), .Z(n948) );
  XNOR U1181 ( .A(n949), .B(sreg[153]), .Z(n943) );
  XNOR U1182 ( .A(n948), .B(n943), .Z(c[153]) );
  NAND U1183 ( .A(b[0]), .B(a[28]), .Z(n954) );
  AND U1184 ( .A(b[1]), .B(a[27]), .Z(n953) );
  XNOR U1185 ( .A(n955), .B(n953), .Z(n947) );
  XNOR U1186 ( .A(n954), .B(n947), .Z(n951) );
  XNOR U1187 ( .A(n952), .B(sreg[154]), .Z(n950) );
  XNOR U1188 ( .A(n951), .B(n950), .Z(c[154]) );
  NAND U1189 ( .A(b[0]), .B(a[29]), .Z(n959) );
  AND U1190 ( .A(b[1]), .B(a[28]), .Z(n958) );
  XNOR U1191 ( .A(n960), .B(n958), .Z(n956) );
  XOR U1192 ( .A(n959), .B(n956), .Z(n963) );
  XNOR U1193 ( .A(n963), .B(sreg[155]), .Z(n957) );
  XOR U1194 ( .A(n962), .B(n957), .Z(c[155]) );
  NAND U1195 ( .A(b[0]), .B(a[30]), .Z(n966) );
  AND U1196 ( .A(b[1]), .B(a[29]), .Z(n965) );
  XNOR U1197 ( .A(n967), .B(n965), .Z(n961) );
  XNOR U1198 ( .A(n966), .B(n961), .Z(n969) );
  XNOR U1199 ( .A(n970), .B(sreg[156]), .Z(n964) );
  XNOR U1200 ( .A(n969), .B(n964), .Z(c[156]) );
  NAND U1201 ( .A(b[0]), .B(a[31]), .Z(n973) );
  AND U1202 ( .A(b[1]), .B(a[30]), .Z(n972) );
  XNOR U1203 ( .A(n974), .B(n972), .Z(n968) );
  XNOR U1204 ( .A(n973), .B(n968), .Z(n976) );
  XNOR U1205 ( .A(n977), .B(sreg[157]), .Z(n971) );
  XNOR U1206 ( .A(n976), .B(n971), .Z(c[157]) );
  NAND U1207 ( .A(b[0]), .B(a[32]), .Z(n980) );
  AND U1208 ( .A(b[1]), .B(a[31]), .Z(n979) );
  XNOR U1209 ( .A(n981), .B(n979), .Z(n975) );
  XNOR U1210 ( .A(n980), .B(n975), .Z(n983) );
  XNOR U1211 ( .A(n984), .B(sreg[158]), .Z(n978) );
  XNOR U1212 ( .A(n983), .B(n978), .Z(c[158]) );
  NAND U1213 ( .A(b[0]), .B(a[33]), .Z(n987) );
  AND U1214 ( .A(b[1]), .B(a[32]), .Z(n986) );
  XNOR U1215 ( .A(n988), .B(n986), .Z(n982) );
  XNOR U1216 ( .A(n987), .B(n982), .Z(n990) );
  XNOR U1217 ( .A(n991), .B(sreg[159]), .Z(n985) );
  XNOR U1218 ( .A(n990), .B(n985), .Z(c[159]) );
  NAND U1219 ( .A(b[0]), .B(a[34]), .Z(n994) );
  AND U1220 ( .A(b[1]), .B(a[33]), .Z(n993) );
  XNOR U1221 ( .A(n995), .B(n993), .Z(n989) );
  XNOR U1222 ( .A(n994), .B(n989), .Z(n997) );
  XNOR U1223 ( .A(n998), .B(sreg[160]), .Z(n992) );
  XNOR U1224 ( .A(n997), .B(n992), .Z(c[160]) );
  NAND U1225 ( .A(b[0]), .B(a[35]), .Z(n1001) );
  AND U1226 ( .A(b[1]), .B(a[34]), .Z(n1000) );
  XNOR U1227 ( .A(n1002), .B(n1000), .Z(n996) );
  XNOR U1228 ( .A(n1001), .B(n996), .Z(n1004) );
  XNOR U1229 ( .A(n1005), .B(sreg[161]), .Z(n999) );
  XNOR U1230 ( .A(n1004), .B(n999), .Z(c[161]) );
  NAND U1231 ( .A(b[0]), .B(a[36]), .Z(n1008) );
  AND U1232 ( .A(b[1]), .B(a[35]), .Z(n1007) );
  XNOR U1233 ( .A(n1009), .B(n1007), .Z(n1003) );
  XNOR U1234 ( .A(n1008), .B(n1003), .Z(n1011) );
  XNOR U1235 ( .A(n1012), .B(sreg[162]), .Z(n1006) );
  XNOR U1236 ( .A(n1011), .B(n1006), .Z(c[162]) );
  NAND U1237 ( .A(b[0]), .B(a[37]), .Z(n1015) );
  AND U1238 ( .A(b[1]), .B(a[36]), .Z(n1014) );
  XNOR U1239 ( .A(n1016), .B(n1014), .Z(n1010) );
  XNOR U1240 ( .A(n1015), .B(n1010), .Z(n1018) );
  XNOR U1241 ( .A(n1019), .B(sreg[163]), .Z(n1013) );
  XNOR U1242 ( .A(n1018), .B(n1013), .Z(c[163]) );
  NAND U1243 ( .A(b[0]), .B(a[38]), .Z(n1022) );
  AND U1244 ( .A(b[1]), .B(a[37]), .Z(n1021) );
  XNOR U1245 ( .A(n1023), .B(n1021), .Z(n1017) );
  XNOR U1246 ( .A(n1022), .B(n1017), .Z(n1025) );
  XNOR U1247 ( .A(n1026), .B(sreg[164]), .Z(n1020) );
  XNOR U1248 ( .A(n1025), .B(n1020), .Z(c[164]) );
  NAND U1249 ( .A(b[0]), .B(a[39]), .Z(n1029) );
  AND U1250 ( .A(b[1]), .B(a[38]), .Z(n1028) );
  XNOR U1251 ( .A(n1030), .B(n1028), .Z(n1024) );
  XNOR U1252 ( .A(n1029), .B(n1024), .Z(n1032) );
  XNOR U1253 ( .A(n1033), .B(sreg[165]), .Z(n1027) );
  XNOR U1254 ( .A(n1032), .B(n1027), .Z(c[165]) );
  NAND U1255 ( .A(b[0]), .B(a[40]), .Z(n1036) );
  AND U1256 ( .A(b[1]), .B(a[39]), .Z(n1035) );
  XNOR U1257 ( .A(n1037), .B(n1035), .Z(n1031) );
  XNOR U1258 ( .A(n1036), .B(n1031), .Z(n1039) );
  XNOR U1259 ( .A(n1040), .B(sreg[166]), .Z(n1034) );
  XNOR U1260 ( .A(n1039), .B(n1034), .Z(c[166]) );
  NAND U1261 ( .A(b[0]), .B(a[41]), .Z(n1043) );
  AND U1262 ( .A(b[1]), .B(a[40]), .Z(n1042) );
  XNOR U1263 ( .A(n1044), .B(n1042), .Z(n1038) );
  XNOR U1264 ( .A(n1043), .B(n1038), .Z(n1046) );
  XNOR U1265 ( .A(n1047), .B(sreg[167]), .Z(n1041) );
  XNOR U1266 ( .A(n1046), .B(n1041), .Z(c[167]) );
  NAND U1267 ( .A(b[0]), .B(a[42]), .Z(n1050) );
  AND U1268 ( .A(b[1]), .B(a[41]), .Z(n1049) );
  XNOR U1269 ( .A(n1051), .B(n1049), .Z(n1045) );
  XNOR U1270 ( .A(n1050), .B(n1045), .Z(n1053) );
  XNOR U1271 ( .A(n1054), .B(sreg[168]), .Z(n1048) );
  XNOR U1272 ( .A(n1053), .B(n1048), .Z(c[168]) );
  NAND U1273 ( .A(b[0]), .B(a[43]), .Z(n1057) );
  AND U1274 ( .A(b[1]), .B(a[42]), .Z(n1056) );
  XNOR U1275 ( .A(n1058), .B(n1056), .Z(n1052) );
  XNOR U1276 ( .A(n1057), .B(n1052), .Z(n1060) );
  XNOR U1277 ( .A(n1061), .B(sreg[169]), .Z(n1055) );
  XNOR U1278 ( .A(n1060), .B(n1055), .Z(c[169]) );
  NAND U1279 ( .A(b[0]), .B(a[44]), .Z(n1064) );
  AND U1280 ( .A(b[1]), .B(a[43]), .Z(n1063) );
  XNOR U1281 ( .A(n1065), .B(n1063), .Z(n1059) );
  XNOR U1282 ( .A(n1064), .B(n1059), .Z(n1067) );
  XNOR U1283 ( .A(n1068), .B(sreg[170]), .Z(n1062) );
  XNOR U1284 ( .A(n1067), .B(n1062), .Z(c[170]) );
  NAND U1285 ( .A(b[0]), .B(a[45]), .Z(n1071) );
  AND U1286 ( .A(b[1]), .B(a[44]), .Z(n1070) );
  XNOR U1287 ( .A(n1072), .B(n1070), .Z(n1066) );
  XNOR U1288 ( .A(n1071), .B(n1066), .Z(n1074) );
  XNOR U1289 ( .A(n1075), .B(sreg[171]), .Z(n1069) );
  XNOR U1290 ( .A(n1074), .B(n1069), .Z(c[171]) );
  NAND U1291 ( .A(b[0]), .B(a[46]), .Z(n1078) );
  AND U1292 ( .A(b[1]), .B(a[45]), .Z(n1077) );
  XNOR U1293 ( .A(n1079), .B(n1077), .Z(n1073) );
  XNOR U1294 ( .A(n1078), .B(n1073), .Z(n1081) );
  XNOR U1295 ( .A(n1082), .B(sreg[172]), .Z(n1076) );
  XNOR U1296 ( .A(n1081), .B(n1076), .Z(c[172]) );
  NAND U1297 ( .A(b[0]), .B(a[47]), .Z(n1085) );
  AND U1298 ( .A(b[1]), .B(a[46]), .Z(n1084) );
  XNOR U1299 ( .A(n1086), .B(n1084), .Z(n1080) );
  XNOR U1300 ( .A(n1085), .B(n1080), .Z(n1088) );
  XNOR U1301 ( .A(n1089), .B(sreg[173]), .Z(n1083) );
  XNOR U1302 ( .A(n1088), .B(n1083), .Z(c[173]) );
  NAND U1303 ( .A(b[0]), .B(a[48]), .Z(n1092) );
  AND U1304 ( .A(b[1]), .B(a[47]), .Z(n1091) );
  XNOR U1305 ( .A(n1093), .B(n1091), .Z(n1087) );
  XNOR U1306 ( .A(n1092), .B(n1087), .Z(n1095) );
  XNOR U1307 ( .A(n1096), .B(sreg[174]), .Z(n1090) );
  XNOR U1308 ( .A(n1095), .B(n1090), .Z(c[174]) );
  NAND U1309 ( .A(b[0]), .B(a[49]), .Z(n1099) );
  AND U1310 ( .A(b[1]), .B(a[48]), .Z(n1098) );
  XNOR U1311 ( .A(n1100), .B(n1098), .Z(n1094) );
  XNOR U1312 ( .A(n1099), .B(n1094), .Z(n1102) );
  XNOR U1313 ( .A(n1103), .B(sreg[175]), .Z(n1097) );
  XNOR U1314 ( .A(n1102), .B(n1097), .Z(c[175]) );
  NAND U1315 ( .A(b[0]), .B(a[50]), .Z(n1106) );
  AND U1316 ( .A(b[1]), .B(a[49]), .Z(n1105) );
  XNOR U1317 ( .A(n1107), .B(n1105), .Z(n1101) );
  XNOR U1318 ( .A(n1106), .B(n1101), .Z(n1109) );
  XNOR U1319 ( .A(n1110), .B(sreg[176]), .Z(n1104) );
  XNOR U1320 ( .A(n1109), .B(n1104), .Z(c[176]) );
  NAND U1321 ( .A(b[0]), .B(a[51]), .Z(n1113) );
  AND U1322 ( .A(b[1]), .B(a[50]), .Z(n1112) );
  XNOR U1323 ( .A(n1114), .B(n1112), .Z(n1108) );
  XNOR U1324 ( .A(n1113), .B(n1108), .Z(n1116) );
  XNOR U1325 ( .A(n1117), .B(sreg[177]), .Z(n1111) );
  XNOR U1326 ( .A(n1116), .B(n1111), .Z(c[177]) );
  NAND U1327 ( .A(b[0]), .B(a[52]), .Z(n1120) );
  AND U1328 ( .A(b[1]), .B(a[51]), .Z(n1119) );
  XNOR U1329 ( .A(n1121), .B(n1119), .Z(n1115) );
  XNOR U1330 ( .A(n1120), .B(n1115), .Z(n1123) );
  XNOR U1331 ( .A(n1124), .B(sreg[178]), .Z(n1118) );
  XNOR U1332 ( .A(n1123), .B(n1118), .Z(c[178]) );
  NAND U1333 ( .A(b[0]), .B(a[53]), .Z(n1127) );
  AND U1334 ( .A(b[1]), .B(a[52]), .Z(n1126) );
  XNOR U1335 ( .A(n1128), .B(n1126), .Z(n1122) );
  XNOR U1336 ( .A(n1127), .B(n1122), .Z(n1130) );
  XNOR U1337 ( .A(n1131), .B(sreg[179]), .Z(n1125) );
  XNOR U1338 ( .A(n1130), .B(n1125), .Z(c[179]) );
  NAND U1339 ( .A(b[0]), .B(a[54]), .Z(n1134) );
  AND U1340 ( .A(b[1]), .B(a[53]), .Z(n1133) );
  XNOR U1341 ( .A(n1135), .B(n1133), .Z(n1129) );
  XNOR U1342 ( .A(n1134), .B(n1129), .Z(n1137) );
  XNOR U1343 ( .A(n1138), .B(sreg[180]), .Z(n1132) );
  XNOR U1344 ( .A(n1137), .B(n1132), .Z(c[180]) );
  NAND U1345 ( .A(b[0]), .B(a[55]), .Z(n1141) );
  AND U1346 ( .A(b[1]), .B(a[54]), .Z(n1140) );
  XNOR U1347 ( .A(n1142), .B(n1140), .Z(n1136) );
  XNOR U1348 ( .A(n1141), .B(n1136), .Z(n1144) );
  XNOR U1349 ( .A(n1145), .B(sreg[181]), .Z(n1139) );
  XNOR U1350 ( .A(n1144), .B(n1139), .Z(c[181]) );
  NAND U1351 ( .A(b[0]), .B(a[56]), .Z(n1148) );
  AND U1352 ( .A(b[1]), .B(a[55]), .Z(n1147) );
  XNOR U1353 ( .A(n1149), .B(n1147), .Z(n1143) );
  XNOR U1354 ( .A(n1148), .B(n1143), .Z(n1151) );
  XNOR U1355 ( .A(n1152), .B(sreg[182]), .Z(n1146) );
  XNOR U1356 ( .A(n1151), .B(n1146), .Z(c[182]) );
  NAND U1357 ( .A(b[0]), .B(a[57]), .Z(n1155) );
  AND U1358 ( .A(b[1]), .B(a[56]), .Z(n1154) );
  XNOR U1359 ( .A(n1156), .B(n1154), .Z(n1150) );
  XNOR U1360 ( .A(n1155), .B(n1150), .Z(n1158) );
  XNOR U1361 ( .A(n1159), .B(sreg[183]), .Z(n1153) );
  XNOR U1362 ( .A(n1158), .B(n1153), .Z(c[183]) );
  NAND U1363 ( .A(b[0]), .B(a[58]), .Z(n1162) );
  AND U1364 ( .A(b[1]), .B(a[57]), .Z(n1161) );
  XNOR U1365 ( .A(n1163), .B(n1161), .Z(n1157) );
  XNOR U1366 ( .A(n1162), .B(n1157), .Z(n1165) );
  XNOR U1367 ( .A(n1166), .B(sreg[184]), .Z(n1160) );
  XNOR U1368 ( .A(n1165), .B(n1160), .Z(c[184]) );
  NAND U1369 ( .A(b[0]), .B(a[59]), .Z(n1169) );
  AND U1370 ( .A(b[1]), .B(a[58]), .Z(n1168) );
  XNOR U1371 ( .A(n1170), .B(n1168), .Z(n1164) );
  XNOR U1372 ( .A(n1169), .B(n1164), .Z(n1172) );
  XNOR U1373 ( .A(n1173), .B(sreg[185]), .Z(n1167) );
  XNOR U1374 ( .A(n1172), .B(n1167), .Z(c[185]) );
  NAND U1375 ( .A(b[0]), .B(a[60]), .Z(n1176) );
  AND U1376 ( .A(b[1]), .B(a[59]), .Z(n1175) );
  XNOR U1377 ( .A(n1177), .B(n1175), .Z(n1171) );
  XNOR U1378 ( .A(n1176), .B(n1171), .Z(n1179) );
  XNOR U1379 ( .A(n1180), .B(sreg[186]), .Z(n1174) );
  XNOR U1380 ( .A(n1179), .B(n1174), .Z(c[186]) );
  NAND U1381 ( .A(b[0]), .B(a[61]), .Z(n1183) );
  AND U1382 ( .A(b[1]), .B(a[60]), .Z(n1182) );
  XNOR U1383 ( .A(n1184), .B(n1182), .Z(n1178) );
  XNOR U1384 ( .A(n1183), .B(n1178), .Z(n1186) );
  XNOR U1385 ( .A(n1187), .B(sreg[187]), .Z(n1181) );
  XNOR U1386 ( .A(n1186), .B(n1181), .Z(c[187]) );
  NAND U1387 ( .A(b[0]), .B(a[62]), .Z(n1190) );
  AND U1388 ( .A(b[1]), .B(a[61]), .Z(n1189) );
  XNOR U1389 ( .A(n1191), .B(n1189), .Z(n1185) );
  XNOR U1390 ( .A(n1190), .B(n1185), .Z(n1193) );
  XNOR U1391 ( .A(n1194), .B(sreg[188]), .Z(n1188) );
  XNOR U1392 ( .A(n1193), .B(n1188), .Z(c[188]) );
  NAND U1393 ( .A(b[0]), .B(a[63]), .Z(n1197) );
  AND U1394 ( .A(b[1]), .B(a[62]), .Z(n1196) );
  XNOR U1395 ( .A(n1198), .B(n1196), .Z(n1192) );
  XNOR U1396 ( .A(n1197), .B(n1192), .Z(n1200) );
  XNOR U1397 ( .A(n1201), .B(sreg[189]), .Z(n1195) );
  XNOR U1398 ( .A(n1200), .B(n1195), .Z(c[189]) );
  NAND U1399 ( .A(b[0]), .B(a[64]), .Z(n1204) );
  AND U1400 ( .A(b[1]), .B(a[63]), .Z(n1203) );
  XNOR U1401 ( .A(n1205), .B(n1203), .Z(n1199) );
  XNOR U1402 ( .A(n1204), .B(n1199), .Z(n1207) );
  XNOR U1403 ( .A(n1208), .B(sreg[190]), .Z(n1202) );
  XNOR U1404 ( .A(n1207), .B(n1202), .Z(c[190]) );
  NAND U1405 ( .A(b[0]), .B(a[65]), .Z(n1211) );
  AND U1406 ( .A(b[1]), .B(a[64]), .Z(n1210) );
  XNOR U1407 ( .A(n1212), .B(n1210), .Z(n1206) );
  XNOR U1408 ( .A(n1211), .B(n1206), .Z(n1214) );
  XNOR U1409 ( .A(n1215), .B(sreg[191]), .Z(n1209) );
  XNOR U1410 ( .A(n1214), .B(n1209), .Z(c[191]) );
  NAND U1411 ( .A(b[0]), .B(a[66]), .Z(n1218) );
  AND U1412 ( .A(b[1]), .B(a[65]), .Z(n1217) );
  XNOR U1413 ( .A(n1219), .B(n1217), .Z(n1213) );
  XNOR U1414 ( .A(n1218), .B(n1213), .Z(n1221) );
  XNOR U1415 ( .A(n1222), .B(sreg[192]), .Z(n1216) );
  XNOR U1416 ( .A(n1221), .B(n1216), .Z(c[192]) );
  NAND U1417 ( .A(b[0]), .B(a[67]), .Z(n1225) );
  AND U1418 ( .A(b[1]), .B(a[66]), .Z(n1224) );
  XNOR U1419 ( .A(n1226), .B(n1224), .Z(n1220) );
  XNOR U1420 ( .A(n1225), .B(n1220), .Z(n1228) );
  XNOR U1421 ( .A(n1229), .B(sreg[193]), .Z(n1223) );
  XNOR U1422 ( .A(n1228), .B(n1223), .Z(c[193]) );
  NAND U1423 ( .A(b[0]), .B(a[68]), .Z(n1232) );
  AND U1424 ( .A(b[1]), .B(a[67]), .Z(n1231) );
  XNOR U1425 ( .A(n1233), .B(n1231), .Z(n1227) );
  XNOR U1426 ( .A(n1232), .B(n1227), .Z(n1235) );
  XNOR U1427 ( .A(n1236), .B(sreg[194]), .Z(n1230) );
  XNOR U1428 ( .A(n1235), .B(n1230), .Z(c[194]) );
  NAND U1429 ( .A(b[0]), .B(a[69]), .Z(n1239) );
  AND U1430 ( .A(b[1]), .B(a[68]), .Z(n1238) );
  XNOR U1431 ( .A(n1240), .B(n1238), .Z(n1234) );
  XNOR U1432 ( .A(n1239), .B(n1234), .Z(n1242) );
  XNOR U1433 ( .A(n1243), .B(sreg[195]), .Z(n1237) );
  XNOR U1434 ( .A(n1242), .B(n1237), .Z(c[195]) );
  NAND U1435 ( .A(b[0]), .B(a[70]), .Z(n1246) );
  AND U1436 ( .A(b[1]), .B(a[69]), .Z(n1245) );
  XNOR U1437 ( .A(n1247), .B(n1245), .Z(n1241) );
  XNOR U1438 ( .A(n1246), .B(n1241), .Z(n1249) );
  XNOR U1439 ( .A(n1250), .B(sreg[196]), .Z(n1244) );
  XNOR U1440 ( .A(n1249), .B(n1244), .Z(c[196]) );
  NAND U1441 ( .A(b[0]), .B(a[71]), .Z(n1253) );
  AND U1442 ( .A(b[1]), .B(a[70]), .Z(n1252) );
  XNOR U1443 ( .A(n1254), .B(n1252), .Z(n1248) );
  XNOR U1444 ( .A(n1253), .B(n1248), .Z(n1256) );
  XNOR U1445 ( .A(n1257), .B(sreg[197]), .Z(n1251) );
  XNOR U1446 ( .A(n1256), .B(n1251), .Z(c[197]) );
  NAND U1447 ( .A(b[0]), .B(a[72]), .Z(n1260) );
  AND U1448 ( .A(b[1]), .B(a[71]), .Z(n1259) );
  XNOR U1449 ( .A(n1261), .B(n1259), .Z(n1255) );
  XNOR U1450 ( .A(n1260), .B(n1255), .Z(n1263) );
  XNOR U1451 ( .A(n1264), .B(sreg[198]), .Z(n1258) );
  XNOR U1452 ( .A(n1263), .B(n1258), .Z(c[198]) );
  NAND U1453 ( .A(b[0]), .B(a[73]), .Z(n1267) );
  AND U1454 ( .A(b[1]), .B(a[72]), .Z(n1266) );
  XNOR U1455 ( .A(n1268), .B(n1266), .Z(n1262) );
  XNOR U1456 ( .A(n1267), .B(n1262), .Z(n1270) );
  XNOR U1457 ( .A(n1271), .B(sreg[199]), .Z(n1265) );
  XNOR U1458 ( .A(n1270), .B(n1265), .Z(c[199]) );
  NAND U1459 ( .A(b[0]), .B(a[74]), .Z(n1274) );
  AND U1460 ( .A(b[1]), .B(a[73]), .Z(n1273) );
  XNOR U1461 ( .A(n1275), .B(n1273), .Z(n1269) );
  XNOR U1462 ( .A(n1274), .B(n1269), .Z(n1277) );
  XNOR U1463 ( .A(n1278), .B(sreg[200]), .Z(n1272) );
  XNOR U1464 ( .A(n1277), .B(n1272), .Z(c[200]) );
  NAND U1465 ( .A(b[0]), .B(a[75]), .Z(n1281) );
  AND U1466 ( .A(b[1]), .B(a[74]), .Z(n1280) );
  XNOR U1467 ( .A(n1282), .B(n1280), .Z(n1276) );
  XNOR U1468 ( .A(n1281), .B(n1276), .Z(n1284) );
  XNOR U1469 ( .A(n1285), .B(sreg[201]), .Z(n1279) );
  XNOR U1470 ( .A(n1284), .B(n1279), .Z(c[201]) );
  NAND U1471 ( .A(b[0]), .B(a[76]), .Z(n1288) );
  AND U1472 ( .A(b[1]), .B(a[75]), .Z(n1287) );
  XNOR U1473 ( .A(n1289), .B(n1287), .Z(n1283) );
  XNOR U1474 ( .A(n1288), .B(n1283), .Z(n1291) );
  XNOR U1475 ( .A(n1292), .B(sreg[202]), .Z(n1286) );
  XNOR U1476 ( .A(n1291), .B(n1286), .Z(c[202]) );
  NAND U1477 ( .A(b[0]), .B(a[77]), .Z(n1295) );
  AND U1478 ( .A(b[1]), .B(a[76]), .Z(n1294) );
  XNOR U1479 ( .A(n1296), .B(n1294), .Z(n1290) );
  XNOR U1480 ( .A(n1295), .B(n1290), .Z(n1298) );
  XNOR U1481 ( .A(n1299), .B(sreg[203]), .Z(n1293) );
  XNOR U1482 ( .A(n1298), .B(n1293), .Z(c[203]) );
  NAND U1483 ( .A(b[0]), .B(a[78]), .Z(n1302) );
  AND U1484 ( .A(b[1]), .B(a[77]), .Z(n1301) );
  XNOR U1485 ( .A(n1303), .B(n1301), .Z(n1297) );
  XNOR U1486 ( .A(n1302), .B(n1297), .Z(n1305) );
  XNOR U1487 ( .A(n1306), .B(sreg[204]), .Z(n1300) );
  XNOR U1488 ( .A(n1305), .B(n1300), .Z(c[204]) );
  NAND U1489 ( .A(b[0]), .B(a[79]), .Z(n1309) );
  AND U1490 ( .A(b[1]), .B(a[78]), .Z(n1308) );
  XNOR U1491 ( .A(n1310), .B(n1308), .Z(n1304) );
  XNOR U1492 ( .A(n1309), .B(n1304), .Z(n1312) );
  XNOR U1493 ( .A(n1313), .B(sreg[205]), .Z(n1307) );
  XNOR U1494 ( .A(n1312), .B(n1307), .Z(c[205]) );
  NAND U1495 ( .A(b[0]), .B(a[80]), .Z(n1316) );
  AND U1496 ( .A(b[1]), .B(a[79]), .Z(n1315) );
  XNOR U1497 ( .A(n1317), .B(n1315), .Z(n1311) );
  XNOR U1498 ( .A(n1316), .B(n1311), .Z(n1319) );
  XNOR U1499 ( .A(n1320), .B(sreg[206]), .Z(n1314) );
  XNOR U1500 ( .A(n1319), .B(n1314), .Z(c[206]) );
  NAND U1501 ( .A(b[0]), .B(a[81]), .Z(n1323) );
  AND U1502 ( .A(b[1]), .B(a[80]), .Z(n1322) );
  XNOR U1503 ( .A(n1324), .B(n1322), .Z(n1318) );
  XNOR U1504 ( .A(n1323), .B(n1318), .Z(n1326) );
  XNOR U1505 ( .A(n1327), .B(sreg[207]), .Z(n1321) );
  XNOR U1506 ( .A(n1326), .B(n1321), .Z(c[207]) );
  NAND U1507 ( .A(b[0]), .B(a[82]), .Z(n1330) );
  AND U1508 ( .A(b[1]), .B(a[81]), .Z(n1329) );
  XNOR U1509 ( .A(n1331), .B(n1329), .Z(n1325) );
  XNOR U1510 ( .A(n1330), .B(n1325), .Z(n1333) );
  XNOR U1511 ( .A(n1334), .B(sreg[208]), .Z(n1328) );
  XNOR U1512 ( .A(n1333), .B(n1328), .Z(c[208]) );
  NAND U1513 ( .A(b[0]), .B(a[83]), .Z(n1337) );
  AND U1514 ( .A(b[1]), .B(a[82]), .Z(n1336) );
  XNOR U1515 ( .A(n1338), .B(n1336), .Z(n1332) );
  XNOR U1516 ( .A(n1337), .B(n1332), .Z(n1340) );
  XNOR U1517 ( .A(n1341), .B(sreg[209]), .Z(n1335) );
  XNOR U1518 ( .A(n1340), .B(n1335), .Z(c[209]) );
  NAND U1519 ( .A(b[0]), .B(a[84]), .Z(n1344) );
  AND U1520 ( .A(b[1]), .B(a[83]), .Z(n1343) );
  XNOR U1521 ( .A(n1345), .B(n1343), .Z(n1339) );
  XNOR U1522 ( .A(n1344), .B(n1339), .Z(n1347) );
  XNOR U1523 ( .A(n1348), .B(sreg[210]), .Z(n1342) );
  XNOR U1524 ( .A(n1347), .B(n1342), .Z(c[210]) );
  NAND U1525 ( .A(b[0]), .B(a[85]), .Z(n1351) );
  AND U1526 ( .A(b[1]), .B(a[84]), .Z(n1350) );
  XNOR U1527 ( .A(n1352), .B(n1350), .Z(n1346) );
  XNOR U1528 ( .A(n1351), .B(n1346), .Z(n1354) );
  XNOR U1529 ( .A(n1355), .B(sreg[211]), .Z(n1349) );
  XNOR U1530 ( .A(n1354), .B(n1349), .Z(c[211]) );
  NAND U1531 ( .A(b[0]), .B(a[86]), .Z(n1358) );
  AND U1532 ( .A(b[1]), .B(a[85]), .Z(n1357) );
  XNOR U1533 ( .A(n1359), .B(n1357), .Z(n1353) );
  XNOR U1534 ( .A(n1358), .B(n1353), .Z(n1361) );
  XNOR U1535 ( .A(n1362), .B(sreg[212]), .Z(n1356) );
  XNOR U1536 ( .A(n1361), .B(n1356), .Z(c[212]) );
  NAND U1537 ( .A(b[0]), .B(a[87]), .Z(n1365) );
  AND U1538 ( .A(b[1]), .B(a[86]), .Z(n1364) );
  XNOR U1539 ( .A(n1366), .B(n1364), .Z(n1360) );
  XNOR U1540 ( .A(n1365), .B(n1360), .Z(n1368) );
  XNOR U1541 ( .A(n1369), .B(sreg[213]), .Z(n1363) );
  XNOR U1542 ( .A(n1368), .B(n1363), .Z(c[213]) );
  NAND U1543 ( .A(b[0]), .B(a[88]), .Z(n1372) );
  AND U1544 ( .A(b[1]), .B(a[87]), .Z(n1371) );
  XNOR U1545 ( .A(n1373), .B(n1371), .Z(n1367) );
  XNOR U1546 ( .A(n1372), .B(n1367), .Z(n1375) );
  XNOR U1547 ( .A(n1376), .B(sreg[214]), .Z(n1370) );
  XNOR U1548 ( .A(n1375), .B(n1370), .Z(c[214]) );
  NAND U1549 ( .A(b[0]), .B(a[89]), .Z(n1379) );
  AND U1550 ( .A(b[1]), .B(a[88]), .Z(n1378) );
  XNOR U1551 ( .A(n1380), .B(n1378), .Z(n1374) );
  XNOR U1552 ( .A(n1379), .B(n1374), .Z(n1382) );
  XNOR U1553 ( .A(n1383), .B(sreg[215]), .Z(n1377) );
  XNOR U1554 ( .A(n1382), .B(n1377), .Z(c[215]) );
  NAND U1555 ( .A(b[0]), .B(a[90]), .Z(n1386) );
  AND U1556 ( .A(b[1]), .B(a[89]), .Z(n1385) );
  XNOR U1557 ( .A(n1387), .B(n1385), .Z(n1381) );
  XNOR U1558 ( .A(n1386), .B(n1381), .Z(n1389) );
  XNOR U1559 ( .A(n1390), .B(sreg[216]), .Z(n1384) );
  XNOR U1560 ( .A(n1389), .B(n1384), .Z(c[216]) );
  NAND U1561 ( .A(b[0]), .B(a[91]), .Z(n1393) );
  AND U1562 ( .A(b[1]), .B(a[90]), .Z(n1392) );
  XNOR U1563 ( .A(n1394), .B(n1392), .Z(n1388) );
  XNOR U1564 ( .A(n1393), .B(n1388), .Z(n1396) );
  XNOR U1565 ( .A(n1397), .B(sreg[217]), .Z(n1391) );
  XNOR U1566 ( .A(n1396), .B(n1391), .Z(c[217]) );
  NAND U1567 ( .A(b[0]), .B(a[92]), .Z(n1400) );
  AND U1568 ( .A(b[1]), .B(a[91]), .Z(n1399) );
  XNOR U1569 ( .A(n1401), .B(n1399), .Z(n1395) );
  XNOR U1570 ( .A(n1400), .B(n1395), .Z(n1403) );
  XNOR U1571 ( .A(n1404), .B(sreg[218]), .Z(n1398) );
  XNOR U1572 ( .A(n1403), .B(n1398), .Z(c[218]) );
  NAND U1573 ( .A(b[0]), .B(a[93]), .Z(n1407) );
  AND U1574 ( .A(b[1]), .B(a[92]), .Z(n1406) );
  XNOR U1575 ( .A(n1408), .B(n1406), .Z(n1402) );
  XNOR U1576 ( .A(n1407), .B(n1402), .Z(n1410) );
  XNOR U1577 ( .A(n1411), .B(sreg[219]), .Z(n1405) );
  XNOR U1578 ( .A(n1410), .B(n1405), .Z(c[219]) );
  NAND U1579 ( .A(b[0]), .B(a[94]), .Z(n1414) );
  AND U1580 ( .A(b[1]), .B(a[93]), .Z(n1413) );
  XNOR U1581 ( .A(n1415), .B(n1413), .Z(n1409) );
  XNOR U1582 ( .A(n1414), .B(n1409), .Z(n1417) );
  XNOR U1583 ( .A(n1418), .B(sreg[220]), .Z(n1412) );
  XNOR U1584 ( .A(n1417), .B(n1412), .Z(c[220]) );
  NAND U1585 ( .A(b[0]), .B(a[95]), .Z(n1421) );
  AND U1586 ( .A(b[1]), .B(a[94]), .Z(n1420) );
  XNOR U1587 ( .A(n1422), .B(n1420), .Z(n1416) );
  XNOR U1588 ( .A(n1421), .B(n1416), .Z(n1424) );
  XNOR U1589 ( .A(n1425), .B(sreg[221]), .Z(n1419) );
  XNOR U1590 ( .A(n1424), .B(n1419), .Z(c[221]) );
  NAND U1591 ( .A(b[0]), .B(a[96]), .Z(n1428) );
  AND U1592 ( .A(b[1]), .B(a[95]), .Z(n1427) );
  XNOR U1593 ( .A(n1429), .B(n1427), .Z(n1423) );
  XNOR U1594 ( .A(n1428), .B(n1423), .Z(n1431) );
  XNOR U1595 ( .A(n1432), .B(sreg[222]), .Z(n1426) );
  XNOR U1596 ( .A(n1431), .B(n1426), .Z(c[222]) );
  NAND U1597 ( .A(b[0]), .B(a[97]), .Z(n1435) );
  AND U1598 ( .A(b[1]), .B(a[96]), .Z(n1434) );
  XNOR U1599 ( .A(n1436), .B(n1434), .Z(n1430) );
  XNOR U1600 ( .A(n1435), .B(n1430), .Z(n1438) );
  XNOR U1601 ( .A(n1439), .B(sreg[223]), .Z(n1433) );
  XNOR U1602 ( .A(n1438), .B(n1433), .Z(c[223]) );
  NAND U1603 ( .A(b[0]), .B(a[98]), .Z(n1442) );
  AND U1604 ( .A(b[1]), .B(a[97]), .Z(n1441) );
  XNOR U1605 ( .A(n1443), .B(n1441), .Z(n1437) );
  XNOR U1606 ( .A(n1442), .B(n1437), .Z(n1445) );
  XNOR U1607 ( .A(n1446), .B(sreg[224]), .Z(n1440) );
  XNOR U1608 ( .A(n1445), .B(n1440), .Z(c[224]) );
  NAND U1609 ( .A(b[0]), .B(a[99]), .Z(n1449) );
  AND U1610 ( .A(b[1]), .B(a[98]), .Z(n1448) );
  XNOR U1611 ( .A(n1450), .B(n1448), .Z(n1444) );
  XNOR U1612 ( .A(n1449), .B(n1444), .Z(n1452) );
  XNOR U1613 ( .A(n1453), .B(sreg[225]), .Z(n1447) );
  XNOR U1614 ( .A(n1452), .B(n1447), .Z(c[225]) );
  NAND U1615 ( .A(b[0]), .B(a[100]), .Z(n1456) );
  AND U1616 ( .A(b[1]), .B(a[99]), .Z(n1455) );
  XNOR U1617 ( .A(n1457), .B(n1455), .Z(n1451) );
  XNOR U1618 ( .A(n1456), .B(n1451), .Z(n1459) );
  XNOR U1619 ( .A(n1460), .B(sreg[226]), .Z(n1454) );
  XNOR U1620 ( .A(n1459), .B(n1454), .Z(c[226]) );
  NAND U1621 ( .A(b[0]), .B(a[101]), .Z(n1463) );
  AND U1622 ( .A(b[1]), .B(a[100]), .Z(n1462) );
  XNOR U1623 ( .A(n1464), .B(n1462), .Z(n1458) );
  XNOR U1624 ( .A(n1463), .B(n1458), .Z(n1466) );
  XNOR U1625 ( .A(n1467), .B(sreg[227]), .Z(n1461) );
  XNOR U1626 ( .A(n1466), .B(n1461), .Z(c[227]) );
  NAND U1627 ( .A(b[0]), .B(a[102]), .Z(n1470) );
  AND U1628 ( .A(b[1]), .B(a[101]), .Z(n1469) );
  XNOR U1629 ( .A(n1471), .B(n1469), .Z(n1465) );
  XNOR U1630 ( .A(n1470), .B(n1465), .Z(n1473) );
  XNOR U1631 ( .A(n1474), .B(sreg[228]), .Z(n1468) );
  XNOR U1632 ( .A(n1473), .B(n1468), .Z(c[228]) );
  NAND U1633 ( .A(b[0]), .B(a[103]), .Z(n1477) );
  AND U1634 ( .A(b[1]), .B(a[102]), .Z(n1476) );
  XNOR U1635 ( .A(n1478), .B(n1476), .Z(n1472) );
  XNOR U1636 ( .A(n1477), .B(n1472), .Z(n1480) );
  XNOR U1637 ( .A(n1481), .B(sreg[229]), .Z(n1475) );
  XNOR U1638 ( .A(n1480), .B(n1475), .Z(c[229]) );
  NAND U1639 ( .A(b[0]), .B(a[104]), .Z(n1484) );
  AND U1640 ( .A(b[1]), .B(a[103]), .Z(n1483) );
  XNOR U1641 ( .A(n1485), .B(n1483), .Z(n1479) );
  XNOR U1642 ( .A(n1484), .B(n1479), .Z(n1487) );
  XNOR U1643 ( .A(n1488), .B(sreg[230]), .Z(n1482) );
  XNOR U1644 ( .A(n1487), .B(n1482), .Z(c[230]) );
  NAND U1645 ( .A(b[0]), .B(a[105]), .Z(n1491) );
  AND U1646 ( .A(b[1]), .B(a[104]), .Z(n1490) );
  XNOR U1647 ( .A(n1492), .B(n1490), .Z(n1486) );
  XNOR U1648 ( .A(n1491), .B(n1486), .Z(n1494) );
  XNOR U1649 ( .A(n1495), .B(sreg[231]), .Z(n1489) );
  XNOR U1650 ( .A(n1494), .B(n1489), .Z(c[231]) );
  NAND U1651 ( .A(b[0]), .B(a[106]), .Z(n1498) );
  AND U1652 ( .A(b[1]), .B(a[105]), .Z(n1497) );
  XNOR U1653 ( .A(n1499), .B(n1497), .Z(n1493) );
  XNOR U1654 ( .A(n1498), .B(n1493), .Z(n1501) );
  XNOR U1655 ( .A(n1502), .B(sreg[232]), .Z(n1496) );
  XNOR U1656 ( .A(n1501), .B(n1496), .Z(c[232]) );
  NAND U1657 ( .A(b[0]), .B(a[107]), .Z(n1505) );
  AND U1658 ( .A(b[1]), .B(a[106]), .Z(n1504) );
  XNOR U1659 ( .A(n1506), .B(n1504), .Z(n1500) );
  XNOR U1660 ( .A(n1505), .B(n1500), .Z(n1508) );
  XNOR U1661 ( .A(n1509), .B(sreg[233]), .Z(n1503) );
  XNOR U1662 ( .A(n1508), .B(n1503), .Z(c[233]) );
  NAND U1663 ( .A(b[0]), .B(a[108]), .Z(n1512) );
  AND U1664 ( .A(b[1]), .B(a[107]), .Z(n1511) );
  XNOR U1665 ( .A(n1513), .B(n1511), .Z(n1507) );
  XNOR U1666 ( .A(n1512), .B(n1507), .Z(n1515) );
  XNOR U1667 ( .A(n1516), .B(sreg[234]), .Z(n1510) );
  XNOR U1668 ( .A(n1515), .B(n1510), .Z(c[234]) );
  NAND U1669 ( .A(b[0]), .B(a[109]), .Z(n1519) );
  AND U1670 ( .A(b[1]), .B(a[108]), .Z(n1518) );
  XNOR U1671 ( .A(n1520), .B(n1518), .Z(n1514) );
  XNOR U1672 ( .A(n1519), .B(n1514), .Z(n1522) );
  XNOR U1673 ( .A(n1523), .B(sreg[235]), .Z(n1517) );
  XNOR U1674 ( .A(n1522), .B(n1517), .Z(c[235]) );
  NAND U1675 ( .A(b[0]), .B(a[110]), .Z(n1526) );
  AND U1676 ( .A(b[1]), .B(a[109]), .Z(n1525) );
  XNOR U1677 ( .A(n1527), .B(n1525), .Z(n1521) );
  XNOR U1678 ( .A(n1526), .B(n1521), .Z(n1529) );
  XNOR U1679 ( .A(n1530), .B(sreg[236]), .Z(n1524) );
  XNOR U1680 ( .A(n1529), .B(n1524), .Z(c[236]) );
  NAND U1681 ( .A(b[0]), .B(a[111]), .Z(n1533) );
  AND U1682 ( .A(b[1]), .B(a[110]), .Z(n1532) );
  XNOR U1683 ( .A(n1534), .B(n1532), .Z(n1528) );
  XNOR U1684 ( .A(n1533), .B(n1528), .Z(n1536) );
  XNOR U1685 ( .A(n1537), .B(sreg[237]), .Z(n1531) );
  XNOR U1686 ( .A(n1536), .B(n1531), .Z(c[237]) );
  NAND U1687 ( .A(b[0]), .B(a[112]), .Z(n1540) );
  AND U1688 ( .A(b[1]), .B(a[111]), .Z(n1539) );
  XNOR U1689 ( .A(n1541), .B(n1539), .Z(n1535) );
  XNOR U1690 ( .A(n1540), .B(n1535), .Z(n1543) );
  XNOR U1691 ( .A(n1544), .B(sreg[238]), .Z(n1538) );
  XNOR U1692 ( .A(n1543), .B(n1538), .Z(c[238]) );
  NAND U1693 ( .A(b[0]), .B(a[113]), .Z(n1547) );
  AND U1694 ( .A(b[1]), .B(a[112]), .Z(n1546) );
  XNOR U1695 ( .A(n1548), .B(n1546), .Z(n1542) );
  XNOR U1696 ( .A(n1547), .B(n1542), .Z(n1550) );
  XNOR U1697 ( .A(n1551), .B(sreg[239]), .Z(n1545) );
  XNOR U1698 ( .A(n1550), .B(n1545), .Z(c[239]) );
  NAND U1699 ( .A(b[0]), .B(a[114]), .Z(n1554) );
  AND U1700 ( .A(b[1]), .B(a[113]), .Z(n1553) );
  XNOR U1701 ( .A(n1555), .B(n1553), .Z(n1549) );
  XNOR U1702 ( .A(n1554), .B(n1549), .Z(n1557) );
  XNOR U1703 ( .A(n1558), .B(sreg[240]), .Z(n1552) );
  XNOR U1704 ( .A(n1557), .B(n1552), .Z(c[240]) );
  NAND U1705 ( .A(b[0]), .B(a[115]), .Z(n1561) );
  AND U1706 ( .A(b[1]), .B(a[114]), .Z(n1560) );
  XNOR U1707 ( .A(n1562), .B(n1560), .Z(n1556) );
  XNOR U1708 ( .A(n1561), .B(n1556), .Z(n1564) );
  XNOR U1709 ( .A(n1565), .B(sreg[241]), .Z(n1559) );
  XNOR U1710 ( .A(n1564), .B(n1559), .Z(c[241]) );
  NAND U1711 ( .A(b[0]), .B(a[116]), .Z(n1568) );
  AND U1712 ( .A(b[1]), .B(a[115]), .Z(n1567) );
  XNOR U1713 ( .A(n1569), .B(n1567), .Z(n1563) );
  XNOR U1714 ( .A(n1568), .B(n1563), .Z(n1571) );
  XNOR U1715 ( .A(n1572), .B(sreg[242]), .Z(n1566) );
  XNOR U1716 ( .A(n1571), .B(n1566), .Z(c[242]) );
  NAND U1717 ( .A(b[0]), .B(a[117]), .Z(n1575) );
  AND U1718 ( .A(b[1]), .B(a[116]), .Z(n1574) );
  XNOR U1719 ( .A(n1576), .B(n1574), .Z(n1570) );
  XNOR U1720 ( .A(n1575), .B(n1570), .Z(n1578) );
  XNOR U1721 ( .A(n1579), .B(sreg[243]), .Z(n1573) );
  XNOR U1722 ( .A(n1578), .B(n1573), .Z(c[243]) );
  NAND U1723 ( .A(b[0]), .B(a[118]), .Z(n1582) );
  AND U1724 ( .A(b[1]), .B(a[117]), .Z(n1581) );
  XNOR U1725 ( .A(n1583), .B(n1581), .Z(n1577) );
  XNOR U1726 ( .A(n1582), .B(n1577), .Z(n1585) );
  XNOR U1727 ( .A(n1586), .B(sreg[244]), .Z(n1580) );
  XNOR U1728 ( .A(n1585), .B(n1580), .Z(c[244]) );
  NAND U1729 ( .A(b[0]), .B(a[119]), .Z(n1589) );
  AND U1730 ( .A(b[1]), .B(a[118]), .Z(n1588) );
  XNOR U1731 ( .A(n1590), .B(n1588), .Z(n1584) );
  XNOR U1732 ( .A(n1589), .B(n1584), .Z(n1592) );
  XNOR U1733 ( .A(n1593), .B(sreg[245]), .Z(n1587) );
  XNOR U1734 ( .A(n1592), .B(n1587), .Z(c[245]) );
  NAND U1735 ( .A(b[0]), .B(a[120]), .Z(n1596) );
  AND U1736 ( .A(b[1]), .B(a[119]), .Z(n1595) );
  XNOR U1737 ( .A(n1597), .B(n1595), .Z(n1591) );
  XNOR U1738 ( .A(n1596), .B(n1591), .Z(n1599) );
  XNOR U1739 ( .A(n1600), .B(sreg[246]), .Z(n1594) );
  XNOR U1740 ( .A(n1599), .B(n1594), .Z(c[246]) );
  NAND U1741 ( .A(b[0]), .B(a[121]), .Z(n1603) );
  AND U1742 ( .A(b[1]), .B(a[120]), .Z(n1602) );
  XNOR U1743 ( .A(n1604), .B(n1602), .Z(n1598) );
  XNOR U1744 ( .A(n1603), .B(n1598), .Z(n1606) );
  XNOR U1745 ( .A(n1607), .B(sreg[247]), .Z(n1601) );
  XNOR U1746 ( .A(n1606), .B(n1601), .Z(c[247]) );
  NAND U1747 ( .A(b[0]), .B(a[122]), .Z(n1610) );
  AND U1748 ( .A(b[1]), .B(a[121]), .Z(n1609) );
  XNOR U1749 ( .A(n1611), .B(n1609), .Z(n1605) );
  XNOR U1750 ( .A(n1610), .B(n1605), .Z(n1613) );
  XNOR U1751 ( .A(n1614), .B(sreg[248]), .Z(n1608) );
  XNOR U1752 ( .A(n1613), .B(n1608), .Z(c[248]) );
  NAND U1753 ( .A(b[0]), .B(a[123]), .Z(n1617) );
  AND U1754 ( .A(b[1]), .B(a[122]), .Z(n1616) );
  XNOR U1755 ( .A(n1618), .B(n1616), .Z(n1612) );
  XNOR U1756 ( .A(n1617), .B(n1612), .Z(n1620) );
  XNOR U1757 ( .A(n1621), .B(sreg[249]), .Z(n1615) );
  XNOR U1758 ( .A(n1620), .B(n1615), .Z(c[249]) );
  NAND U1759 ( .A(b[0]), .B(a[124]), .Z(n1624) );
  AND U1760 ( .A(b[1]), .B(a[123]), .Z(n1623) );
  XNOR U1761 ( .A(n1625), .B(n1623), .Z(n1619) );
  XNOR U1762 ( .A(n1624), .B(n1619), .Z(n1627) );
  XNOR U1763 ( .A(n1628), .B(sreg[250]), .Z(n1622) );
  XNOR U1764 ( .A(n1627), .B(n1622), .Z(c[250]) );
  NAND U1765 ( .A(b[0]), .B(a[125]), .Z(n1631) );
  AND U1766 ( .A(b[1]), .B(a[124]), .Z(n1630) );
  XNOR U1767 ( .A(n1632), .B(n1630), .Z(n1626) );
  XNOR U1768 ( .A(n1631), .B(n1626), .Z(n1634) );
  XNOR U1769 ( .A(n1635), .B(sreg[251]), .Z(n1629) );
  XNOR U1770 ( .A(n1634), .B(n1629), .Z(c[251]) );
  NAND U1771 ( .A(a[126]), .B(b[0]), .Z(n1638) );
  AND U1772 ( .A(b[1]), .B(a[125]), .Z(n1637) );
  XNOR U1773 ( .A(n1639), .B(n1637), .Z(n1633) );
  XNOR U1774 ( .A(n1638), .B(n1633), .Z(n1640) );
  XNOR U1775 ( .A(n1641), .B(sreg[252]), .Z(n1636) );
  XNOR U1776 ( .A(n1640), .B(n1636), .Z(c[252]) );
  AND U1777 ( .A(b[1]), .B(a[126]), .Z(n1645) );
  NAND U1778 ( .A(b[0]), .B(a[127]), .Z(n1646) );
  XNOR U1779 ( .A(n1645), .B(n1646), .Z(n1648) );
  XNOR U1780 ( .A(n1648), .B(n1647), .Z(n1643) );
  XNOR U1781 ( .A(n1644), .B(sreg[253]), .Z(n1642) );
  XNOR U1782 ( .A(n1643), .B(n1642), .Z(c[253]) );
  NANDN U1783 ( .A(n1646), .B(n1645), .Z(n1650) );
  NAND U1784 ( .A(n1648), .B(n1647), .Z(n1649) );
  AND U1785 ( .A(n1650), .B(n1649), .Z(n1654) );
  AND U1786 ( .A(b[1]), .B(a[127]), .Z(n1652) );
  XNOR U1787 ( .A(n1654), .B(n1652), .Z(n1651) );
  XNOR U1788 ( .A(n1653), .B(n1651), .Z(c[254]) );
endmodule

