
module mult_N256_CC128 ( clk, rst, a, b, c );
  input [255:0] a;
  input [1:0] b;
  output [511:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070;
  wire   [511:0] sreg;

  DFF \sreg_reg[509]  ( .D(c[511]), .CLK(clk), .RST(rst), .Q(sreg[509]) );
  DFF \sreg_reg[508]  ( .D(c[510]), .CLK(clk), .RST(rst), .Q(sreg[508]) );
  DFF \sreg_reg[507]  ( .D(c[509]), .CLK(clk), .RST(rst), .Q(sreg[507]) );
  DFF \sreg_reg[506]  ( .D(c[508]), .CLK(clk), .RST(rst), .Q(sreg[506]) );
  DFF \sreg_reg[505]  ( .D(c[507]), .CLK(clk), .RST(rst), .Q(sreg[505]) );
  DFF \sreg_reg[504]  ( .D(c[506]), .CLK(clk), .RST(rst), .Q(sreg[504]) );
  DFF \sreg_reg[503]  ( .D(c[505]), .CLK(clk), .RST(rst), .Q(sreg[503]) );
  DFF \sreg_reg[502]  ( .D(c[504]), .CLK(clk), .RST(rst), .Q(sreg[502]) );
  DFF \sreg_reg[501]  ( .D(c[503]), .CLK(clk), .RST(rst), .Q(sreg[501]) );
  DFF \sreg_reg[500]  ( .D(c[502]), .CLK(clk), .RST(rst), .Q(sreg[500]) );
  DFF \sreg_reg[499]  ( .D(c[501]), .CLK(clk), .RST(rst), .Q(sreg[499]) );
  DFF \sreg_reg[498]  ( .D(c[500]), .CLK(clk), .RST(rst), .Q(sreg[498]) );
  DFF \sreg_reg[497]  ( .D(c[499]), .CLK(clk), .RST(rst), .Q(sreg[497]) );
  DFF \sreg_reg[496]  ( .D(c[498]), .CLK(clk), .RST(rst), .Q(sreg[496]) );
  DFF \sreg_reg[495]  ( .D(c[497]), .CLK(clk), .RST(rst), .Q(sreg[495]) );
  DFF \sreg_reg[494]  ( .D(c[496]), .CLK(clk), .RST(rst), .Q(sreg[494]) );
  DFF \sreg_reg[493]  ( .D(c[495]), .CLK(clk), .RST(rst), .Q(sreg[493]) );
  DFF \sreg_reg[492]  ( .D(c[494]), .CLK(clk), .RST(rst), .Q(sreg[492]) );
  DFF \sreg_reg[491]  ( .D(c[493]), .CLK(clk), .RST(rst), .Q(sreg[491]) );
  DFF \sreg_reg[490]  ( .D(c[492]), .CLK(clk), .RST(rst), .Q(sreg[490]) );
  DFF \sreg_reg[489]  ( .D(c[491]), .CLK(clk), .RST(rst), .Q(sreg[489]) );
  DFF \sreg_reg[488]  ( .D(c[490]), .CLK(clk), .RST(rst), .Q(sreg[488]) );
  DFF \sreg_reg[487]  ( .D(c[489]), .CLK(clk), .RST(rst), .Q(sreg[487]) );
  DFF \sreg_reg[486]  ( .D(c[488]), .CLK(clk), .RST(rst), .Q(sreg[486]) );
  DFF \sreg_reg[485]  ( .D(c[487]), .CLK(clk), .RST(rst), .Q(sreg[485]) );
  DFF \sreg_reg[484]  ( .D(c[486]), .CLK(clk), .RST(rst), .Q(sreg[484]) );
  DFF \sreg_reg[483]  ( .D(c[485]), .CLK(clk), .RST(rst), .Q(sreg[483]) );
  DFF \sreg_reg[482]  ( .D(c[484]), .CLK(clk), .RST(rst), .Q(sreg[482]) );
  DFF \sreg_reg[481]  ( .D(c[483]), .CLK(clk), .RST(rst), .Q(sreg[481]) );
  DFF \sreg_reg[480]  ( .D(c[482]), .CLK(clk), .RST(rst), .Q(sreg[480]) );
  DFF \sreg_reg[479]  ( .D(c[481]), .CLK(clk), .RST(rst), .Q(sreg[479]) );
  DFF \sreg_reg[478]  ( .D(c[480]), .CLK(clk), .RST(rst), .Q(sreg[478]) );
  DFF \sreg_reg[477]  ( .D(c[479]), .CLK(clk), .RST(rst), .Q(sreg[477]) );
  DFF \sreg_reg[476]  ( .D(c[478]), .CLK(clk), .RST(rst), .Q(sreg[476]) );
  DFF \sreg_reg[475]  ( .D(c[477]), .CLK(clk), .RST(rst), .Q(sreg[475]) );
  DFF \sreg_reg[474]  ( .D(c[476]), .CLK(clk), .RST(rst), .Q(sreg[474]) );
  DFF \sreg_reg[473]  ( .D(c[475]), .CLK(clk), .RST(rst), .Q(sreg[473]) );
  DFF \sreg_reg[472]  ( .D(c[474]), .CLK(clk), .RST(rst), .Q(sreg[472]) );
  DFF \sreg_reg[471]  ( .D(c[473]), .CLK(clk), .RST(rst), .Q(sreg[471]) );
  DFF \sreg_reg[470]  ( .D(c[472]), .CLK(clk), .RST(rst), .Q(sreg[470]) );
  DFF \sreg_reg[469]  ( .D(c[471]), .CLK(clk), .RST(rst), .Q(sreg[469]) );
  DFF \sreg_reg[468]  ( .D(c[470]), .CLK(clk), .RST(rst), .Q(sreg[468]) );
  DFF \sreg_reg[467]  ( .D(c[469]), .CLK(clk), .RST(rst), .Q(sreg[467]) );
  DFF \sreg_reg[466]  ( .D(c[468]), .CLK(clk), .RST(rst), .Q(sreg[466]) );
  DFF \sreg_reg[465]  ( .D(c[467]), .CLK(clk), .RST(rst), .Q(sreg[465]) );
  DFF \sreg_reg[464]  ( .D(c[466]), .CLK(clk), .RST(rst), .Q(sreg[464]) );
  DFF \sreg_reg[463]  ( .D(c[465]), .CLK(clk), .RST(rst), .Q(sreg[463]) );
  DFF \sreg_reg[462]  ( .D(c[464]), .CLK(clk), .RST(rst), .Q(sreg[462]) );
  DFF \sreg_reg[461]  ( .D(c[463]), .CLK(clk), .RST(rst), .Q(sreg[461]) );
  DFF \sreg_reg[460]  ( .D(c[462]), .CLK(clk), .RST(rst), .Q(sreg[460]) );
  DFF \sreg_reg[459]  ( .D(c[461]), .CLK(clk), .RST(rst), .Q(sreg[459]) );
  DFF \sreg_reg[458]  ( .D(c[460]), .CLK(clk), .RST(rst), .Q(sreg[458]) );
  DFF \sreg_reg[457]  ( .D(c[459]), .CLK(clk), .RST(rst), .Q(sreg[457]) );
  DFF \sreg_reg[456]  ( .D(c[458]), .CLK(clk), .RST(rst), .Q(sreg[456]) );
  DFF \sreg_reg[455]  ( .D(c[457]), .CLK(clk), .RST(rst), .Q(sreg[455]) );
  DFF \sreg_reg[454]  ( .D(c[456]), .CLK(clk), .RST(rst), .Q(sreg[454]) );
  DFF \sreg_reg[453]  ( .D(c[455]), .CLK(clk), .RST(rst), .Q(sreg[453]) );
  DFF \sreg_reg[452]  ( .D(c[454]), .CLK(clk), .RST(rst), .Q(sreg[452]) );
  DFF \sreg_reg[451]  ( .D(c[453]), .CLK(clk), .RST(rst), .Q(sreg[451]) );
  DFF \sreg_reg[450]  ( .D(c[452]), .CLK(clk), .RST(rst), .Q(sreg[450]) );
  DFF \sreg_reg[449]  ( .D(c[451]), .CLK(clk), .RST(rst), .Q(sreg[449]) );
  DFF \sreg_reg[448]  ( .D(c[450]), .CLK(clk), .RST(rst), .Q(sreg[448]) );
  DFF \sreg_reg[447]  ( .D(c[449]), .CLK(clk), .RST(rst), .Q(sreg[447]) );
  DFF \sreg_reg[446]  ( .D(c[448]), .CLK(clk), .RST(rst), .Q(sreg[446]) );
  DFF \sreg_reg[445]  ( .D(c[447]), .CLK(clk), .RST(rst), .Q(sreg[445]) );
  DFF \sreg_reg[444]  ( .D(c[446]), .CLK(clk), .RST(rst), .Q(sreg[444]) );
  DFF \sreg_reg[443]  ( .D(c[445]), .CLK(clk), .RST(rst), .Q(sreg[443]) );
  DFF \sreg_reg[442]  ( .D(c[444]), .CLK(clk), .RST(rst), .Q(sreg[442]) );
  DFF \sreg_reg[441]  ( .D(c[443]), .CLK(clk), .RST(rst), .Q(sreg[441]) );
  DFF \sreg_reg[440]  ( .D(c[442]), .CLK(clk), .RST(rst), .Q(sreg[440]) );
  DFF \sreg_reg[439]  ( .D(c[441]), .CLK(clk), .RST(rst), .Q(sreg[439]) );
  DFF \sreg_reg[438]  ( .D(c[440]), .CLK(clk), .RST(rst), .Q(sreg[438]) );
  DFF \sreg_reg[437]  ( .D(c[439]), .CLK(clk), .RST(rst), .Q(sreg[437]) );
  DFF \sreg_reg[436]  ( .D(c[438]), .CLK(clk), .RST(rst), .Q(sreg[436]) );
  DFF \sreg_reg[435]  ( .D(c[437]), .CLK(clk), .RST(rst), .Q(sreg[435]) );
  DFF \sreg_reg[434]  ( .D(c[436]), .CLK(clk), .RST(rst), .Q(sreg[434]) );
  DFF \sreg_reg[433]  ( .D(c[435]), .CLK(clk), .RST(rst), .Q(sreg[433]) );
  DFF \sreg_reg[432]  ( .D(c[434]), .CLK(clk), .RST(rst), .Q(sreg[432]) );
  DFF \sreg_reg[431]  ( .D(c[433]), .CLK(clk), .RST(rst), .Q(sreg[431]) );
  DFF \sreg_reg[430]  ( .D(c[432]), .CLK(clk), .RST(rst), .Q(sreg[430]) );
  DFF \sreg_reg[429]  ( .D(c[431]), .CLK(clk), .RST(rst), .Q(sreg[429]) );
  DFF \sreg_reg[428]  ( .D(c[430]), .CLK(clk), .RST(rst), .Q(sreg[428]) );
  DFF \sreg_reg[427]  ( .D(c[429]), .CLK(clk), .RST(rst), .Q(sreg[427]) );
  DFF \sreg_reg[426]  ( .D(c[428]), .CLK(clk), .RST(rst), .Q(sreg[426]) );
  DFF \sreg_reg[425]  ( .D(c[427]), .CLK(clk), .RST(rst), .Q(sreg[425]) );
  DFF \sreg_reg[424]  ( .D(c[426]), .CLK(clk), .RST(rst), .Q(sreg[424]) );
  DFF \sreg_reg[423]  ( .D(c[425]), .CLK(clk), .RST(rst), .Q(sreg[423]) );
  DFF \sreg_reg[422]  ( .D(c[424]), .CLK(clk), .RST(rst), .Q(sreg[422]) );
  DFF \sreg_reg[421]  ( .D(c[423]), .CLK(clk), .RST(rst), .Q(sreg[421]) );
  DFF \sreg_reg[420]  ( .D(c[422]), .CLK(clk), .RST(rst), .Q(sreg[420]) );
  DFF \sreg_reg[419]  ( .D(c[421]), .CLK(clk), .RST(rst), .Q(sreg[419]) );
  DFF \sreg_reg[418]  ( .D(c[420]), .CLK(clk), .RST(rst), .Q(sreg[418]) );
  DFF \sreg_reg[417]  ( .D(c[419]), .CLK(clk), .RST(rst), .Q(sreg[417]) );
  DFF \sreg_reg[416]  ( .D(c[418]), .CLK(clk), .RST(rst), .Q(sreg[416]) );
  DFF \sreg_reg[415]  ( .D(c[417]), .CLK(clk), .RST(rst), .Q(sreg[415]) );
  DFF \sreg_reg[414]  ( .D(c[416]), .CLK(clk), .RST(rst), .Q(sreg[414]) );
  DFF \sreg_reg[413]  ( .D(c[415]), .CLK(clk), .RST(rst), .Q(sreg[413]) );
  DFF \sreg_reg[412]  ( .D(c[414]), .CLK(clk), .RST(rst), .Q(sreg[412]) );
  DFF \sreg_reg[411]  ( .D(c[413]), .CLK(clk), .RST(rst), .Q(sreg[411]) );
  DFF \sreg_reg[410]  ( .D(c[412]), .CLK(clk), .RST(rst), .Q(sreg[410]) );
  DFF \sreg_reg[409]  ( .D(c[411]), .CLK(clk), .RST(rst), .Q(sreg[409]) );
  DFF \sreg_reg[408]  ( .D(c[410]), .CLK(clk), .RST(rst), .Q(sreg[408]) );
  DFF \sreg_reg[407]  ( .D(c[409]), .CLK(clk), .RST(rst), .Q(sreg[407]) );
  DFF \sreg_reg[406]  ( .D(c[408]), .CLK(clk), .RST(rst), .Q(sreg[406]) );
  DFF \sreg_reg[405]  ( .D(c[407]), .CLK(clk), .RST(rst), .Q(sreg[405]) );
  DFF \sreg_reg[404]  ( .D(c[406]), .CLK(clk), .RST(rst), .Q(sreg[404]) );
  DFF \sreg_reg[403]  ( .D(c[405]), .CLK(clk), .RST(rst), .Q(sreg[403]) );
  DFF \sreg_reg[402]  ( .D(c[404]), .CLK(clk), .RST(rst), .Q(sreg[402]) );
  DFF \sreg_reg[401]  ( .D(c[403]), .CLK(clk), .RST(rst), .Q(sreg[401]) );
  DFF \sreg_reg[400]  ( .D(c[402]), .CLK(clk), .RST(rst), .Q(sreg[400]) );
  DFF \sreg_reg[399]  ( .D(c[401]), .CLK(clk), .RST(rst), .Q(sreg[399]) );
  DFF \sreg_reg[398]  ( .D(c[400]), .CLK(clk), .RST(rst), .Q(sreg[398]) );
  DFF \sreg_reg[397]  ( .D(c[399]), .CLK(clk), .RST(rst), .Q(sreg[397]) );
  DFF \sreg_reg[396]  ( .D(c[398]), .CLK(clk), .RST(rst), .Q(sreg[396]) );
  DFF \sreg_reg[395]  ( .D(c[397]), .CLK(clk), .RST(rst), .Q(sreg[395]) );
  DFF \sreg_reg[394]  ( .D(c[396]), .CLK(clk), .RST(rst), .Q(sreg[394]) );
  DFF \sreg_reg[393]  ( .D(c[395]), .CLK(clk), .RST(rst), .Q(sreg[393]) );
  DFF \sreg_reg[392]  ( .D(c[394]), .CLK(clk), .RST(rst), .Q(sreg[392]) );
  DFF \sreg_reg[391]  ( .D(c[393]), .CLK(clk), .RST(rst), .Q(sreg[391]) );
  DFF \sreg_reg[390]  ( .D(c[392]), .CLK(clk), .RST(rst), .Q(sreg[390]) );
  DFF \sreg_reg[389]  ( .D(c[391]), .CLK(clk), .RST(rst), .Q(sreg[389]) );
  DFF \sreg_reg[388]  ( .D(c[390]), .CLK(clk), .RST(rst), .Q(sreg[388]) );
  DFF \sreg_reg[387]  ( .D(c[389]), .CLK(clk), .RST(rst), .Q(sreg[387]) );
  DFF \sreg_reg[386]  ( .D(c[388]), .CLK(clk), .RST(rst), .Q(sreg[386]) );
  DFF \sreg_reg[385]  ( .D(c[387]), .CLK(clk), .RST(rst), .Q(sreg[385]) );
  DFF \sreg_reg[384]  ( .D(c[386]), .CLK(clk), .RST(rst), .Q(sreg[384]) );
  DFF \sreg_reg[383]  ( .D(c[385]), .CLK(clk), .RST(rst), .Q(sreg[383]) );
  DFF \sreg_reg[382]  ( .D(c[384]), .CLK(clk), .RST(rst), .Q(sreg[382]) );
  DFF \sreg_reg[381]  ( .D(c[383]), .CLK(clk), .RST(rst), .Q(sreg[381]) );
  DFF \sreg_reg[380]  ( .D(c[382]), .CLK(clk), .RST(rst), .Q(sreg[380]) );
  DFF \sreg_reg[379]  ( .D(c[381]), .CLK(clk), .RST(rst), .Q(sreg[379]) );
  DFF \sreg_reg[378]  ( .D(c[380]), .CLK(clk), .RST(rst), .Q(sreg[378]) );
  DFF \sreg_reg[377]  ( .D(c[379]), .CLK(clk), .RST(rst), .Q(sreg[377]) );
  DFF \sreg_reg[376]  ( .D(c[378]), .CLK(clk), .RST(rst), .Q(sreg[376]) );
  DFF \sreg_reg[375]  ( .D(c[377]), .CLK(clk), .RST(rst), .Q(sreg[375]) );
  DFF \sreg_reg[374]  ( .D(c[376]), .CLK(clk), .RST(rst), .Q(sreg[374]) );
  DFF \sreg_reg[373]  ( .D(c[375]), .CLK(clk), .RST(rst), .Q(sreg[373]) );
  DFF \sreg_reg[372]  ( .D(c[374]), .CLK(clk), .RST(rst), .Q(sreg[372]) );
  DFF \sreg_reg[371]  ( .D(c[373]), .CLK(clk), .RST(rst), .Q(sreg[371]) );
  DFF \sreg_reg[370]  ( .D(c[372]), .CLK(clk), .RST(rst), .Q(sreg[370]) );
  DFF \sreg_reg[369]  ( .D(c[371]), .CLK(clk), .RST(rst), .Q(sreg[369]) );
  DFF \sreg_reg[368]  ( .D(c[370]), .CLK(clk), .RST(rst), .Q(sreg[368]) );
  DFF \sreg_reg[367]  ( .D(c[369]), .CLK(clk), .RST(rst), .Q(sreg[367]) );
  DFF \sreg_reg[366]  ( .D(c[368]), .CLK(clk), .RST(rst), .Q(sreg[366]) );
  DFF \sreg_reg[365]  ( .D(c[367]), .CLK(clk), .RST(rst), .Q(sreg[365]) );
  DFF \sreg_reg[364]  ( .D(c[366]), .CLK(clk), .RST(rst), .Q(sreg[364]) );
  DFF \sreg_reg[363]  ( .D(c[365]), .CLK(clk), .RST(rst), .Q(sreg[363]) );
  DFF \sreg_reg[362]  ( .D(c[364]), .CLK(clk), .RST(rst), .Q(sreg[362]) );
  DFF \sreg_reg[361]  ( .D(c[363]), .CLK(clk), .RST(rst), .Q(sreg[361]) );
  DFF \sreg_reg[360]  ( .D(c[362]), .CLK(clk), .RST(rst), .Q(sreg[360]) );
  DFF \sreg_reg[359]  ( .D(c[361]), .CLK(clk), .RST(rst), .Q(sreg[359]) );
  DFF \sreg_reg[358]  ( .D(c[360]), .CLK(clk), .RST(rst), .Q(sreg[358]) );
  DFF \sreg_reg[357]  ( .D(c[359]), .CLK(clk), .RST(rst), .Q(sreg[357]) );
  DFF \sreg_reg[356]  ( .D(c[358]), .CLK(clk), .RST(rst), .Q(sreg[356]) );
  DFF \sreg_reg[355]  ( .D(c[357]), .CLK(clk), .RST(rst), .Q(sreg[355]) );
  DFF \sreg_reg[354]  ( .D(c[356]), .CLK(clk), .RST(rst), .Q(sreg[354]) );
  DFF \sreg_reg[353]  ( .D(c[355]), .CLK(clk), .RST(rst), .Q(sreg[353]) );
  DFF \sreg_reg[352]  ( .D(c[354]), .CLK(clk), .RST(rst), .Q(sreg[352]) );
  DFF \sreg_reg[351]  ( .D(c[353]), .CLK(clk), .RST(rst), .Q(sreg[351]) );
  DFF \sreg_reg[350]  ( .D(c[352]), .CLK(clk), .RST(rst), .Q(sreg[350]) );
  DFF \sreg_reg[349]  ( .D(c[351]), .CLK(clk), .RST(rst), .Q(sreg[349]) );
  DFF \sreg_reg[348]  ( .D(c[350]), .CLK(clk), .RST(rst), .Q(sreg[348]) );
  DFF \sreg_reg[347]  ( .D(c[349]), .CLK(clk), .RST(rst), .Q(sreg[347]) );
  DFF \sreg_reg[346]  ( .D(c[348]), .CLK(clk), .RST(rst), .Q(sreg[346]) );
  DFF \sreg_reg[345]  ( .D(c[347]), .CLK(clk), .RST(rst), .Q(sreg[345]) );
  DFF \sreg_reg[344]  ( .D(c[346]), .CLK(clk), .RST(rst), .Q(sreg[344]) );
  DFF \sreg_reg[343]  ( .D(c[345]), .CLK(clk), .RST(rst), .Q(sreg[343]) );
  DFF \sreg_reg[342]  ( .D(c[344]), .CLK(clk), .RST(rst), .Q(sreg[342]) );
  DFF \sreg_reg[341]  ( .D(c[343]), .CLK(clk), .RST(rst), .Q(sreg[341]) );
  DFF \sreg_reg[340]  ( .D(c[342]), .CLK(clk), .RST(rst), .Q(sreg[340]) );
  DFF \sreg_reg[339]  ( .D(c[341]), .CLK(clk), .RST(rst), .Q(sreg[339]) );
  DFF \sreg_reg[338]  ( .D(c[340]), .CLK(clk), .RST(rst), .Q(sreg[338]) );
  DFF \sreg_reg[337]  ( .D(c[339]), .CLK(clk), .RST(rst), .Q(sreg[337]) );
  DFF \sreg_reg[336]  ( .D(c[338]), .CLK(clk), .RST(rst), .Q(sreg[336]) );
  DFF \sreg_reg[335]  ( .D(c[337]), .CLK(clk), .RST(rst), .Q(sreg[335]) );
  DFF \sreg_reg[334]  ( .D(c[336]), .CLK(clk), .RST(rst), .Q(sreg[334]) );
  DFF \sreg_reg[333]  ( .D(c[335]), .CLK(clk), .RST(rst), .Q(sreg[333]) );
  DFF \sreg_reg[332]  ( .D(c[334]), .CLK(clk), .RST(rst), .Q(sreg[332]) );
  DFF \sreg_reg[331]  ( .D(c[333]), .CLK(clk), .RST(rst), .Q(sreg[331]) );
  DFF \sreg_reg[330]  ( .D(c[332]), .CLK(clk), .RST(rst), .Q(sreg[330]) );
  DFF \sreg_reg[329]  ( .D(c[331]), .CLK(clk), .RST(rst), .Q(sreg[329]) );
  DFF \sreg_reg[328]  ( .D(c[330]), .CLK(clk), .RST(rst), .Q(sreg[328]) );
  DFF \sreg_reg[327]  ( .D(c[329]), .CLK(clk), .RST(rst), .Q(sreg[327]) );
  DFF \sreg_reg[326]  ( .D(c[328]), .CLK(clk), .RST(rst), .Q(sreg[326]) );
  DFF \sreg_reg[325]  ( .D(c[327]), .CLK(clk), .RST(rst), .Q(sreg[325]) );
  DFF \sreg_reg[324]  ( .D(c[326]), .CLK(clk), .RST(rst), .Q(sreg[324]) );
  DFF \sreg_reg[323]  ( .D(c[325]), .CLK(clk), .RST(rst), .Q(sreg[323]) );
  DFF \sreg_reg[322]  ( .D(c[324]), .CLK(clk), .RST(rst), .Q(sreg[322]) );
  DFF \sreg_reg[321]  ( .D(c[323]), .CLK(clk), .RST(rst), .Q(sreg[321]) );
  DFF \sreg_reg[320]  ( .D(c[322]), .CLK(clk), .RST(rst), .Q(sreg[320]) );
  DFF \sreg_reg[319]  ( .D(c[321]), .CLK(clk), .RST(rst), .Q(sreg[319]) );
  DFF \sreg_reg[318]  ( .D(c[320]), .CLK(clk), .RST(rst), .Q(sreg[318]) );
  DFF \sreg_reg[317]  ( .D(c[319]), .CLK(clk), .RST(rst), .Q(sreg[317]) );
  DFF \sreg_reg[316]  ( .D(c[318]), .CLK(clk), .RST(rst), .Q(sreg[316]) );
  DFF \sreg_reg[315]  ( .D(c[317]), .CLK(clk), .RST(rst), .Q(sreg[315]) );
  DFF \sreg_reg[314]  ( .D(c[316]), .CLK(clk), .RST(rst), .Q(sreg[314]) );
  DFF \sreg_reg[313]  ( .D(c[315]), .CLK(clk), .RST(rst), .Q(sreg[313]) );
  DFF \sreg_reg[312]  ( .D(c[314]), .CLK(clk), .RST(rst), .Q(sreg[312]) );
  DFF \sreg_reg[311]  ( .D(c[313]), .CLK(clk), .RST(rst), .Q(sreg[311]) );
  DFF \sreg_reg[310]  ( .D(c[312]), .CLK(clk), .RST(rst), .Q(sreg[310]) );
  DFF \sreg_reg[309]  ( .D(c[311]), .CLK(clk), .RST(rst), .Q(sreg[309]) );
  DFF \sreg_reg[308]  ( .D(c[310]), .CLK(clk), .RST(rst), .Q(sreg[308]) );
  DFF \sreg_reg[307]  ( .D(c[309]), .CLK(clk), .RST(rst), .Q(sreg[307]) );
  DFF \sreg_reg[306]  ( .D(c[308]), .CLK(clk), .RST(rst), .Q(sreg[306]) );
  DFF \sreg_reg[305]  ( .D(c[307]), .CLK(clk), .RST(rst), .Q(sreg[305]) );
  DFF \sreg_reg[304]  ( .D(c[306]), .CLK(clk), .RST(rst), .Q(sreg[304]) );
  DFF \sreg_reg[303]  ( .D(c[305]), .CLK(clk), .RST(rst), .Q(sreg[303]) );
  DFF \sreg_reg[302]  ( .D(c[304]), .CLK(clk), .RST(rst), .Q(sreg[302]) );
  DFF \sreg_reg[301]  ( .D(c[303]), .CLK(clk), .RST(rst), .Q(sreg[301]) );
  DFF \sreg_reg[300]  ( .D(c[302]), .CLK(clk), .RST(rst), .Q(sreg[300]) );
  DFF \sreg_reg[299]  ( .D(c[301]), .CLK(clk), .RST(rst), .Q(sreg[299]) );
  DFF \sreg_reg[298]  ( .D(c[300]), .CLK(clk), .RST(rst), .Q(sreg[298]) );
  DFF \sreg_reg[297]  ( .D(c[299]), .CLK(clk), .RST(rst), .Q(sreg[297]) );
  DFF \sreg_reg[296]  ( .D(c[298]), .CLK(clk), .RST(rst), .Q(sreg[296]) );
  DFF \sreg_reg[295]  ( .D(c[297]), .CLK(clk), .RST(rst), .Q(sreg[295]) );
  DFF \sreg_reg[294]  ( .D(c[296]), .CLK(clk), .RST(rst), .Q(sreg[294]) );
  DFF \sreg_reg[293]  ( .D(c[295]), .CLK(clk), .RST(rst), .Q(sreg[293]) );
  DFF \sreg_reg[292]  ( .D(c[294]), .CLK(clk), .RST(rst), .Q(sreg[292]) );
  DFF \sreg_reg[291]  ( .D(c[293]), .CLK(clk), .RST(rst), .Q(sreg[291]) );
  DFF \sreg_reg[290]  ( .D(c[292]), .CLK(clk), .RST(rst), .Q(sreg[290]) );
  DFF \sreg_reg[289]  ( .D(c[291]), .CLK(clk), .RST(rst), .Q(sreg[289]) );
  DFF \sreg_reg[288]  ( .D(c[290]), .CLK(clk), .RST(rst), .Q(sreg[288]) );
  DFF \sreg_reg[287]  ( .D(c[289]), .CLK(clk), .RST(rst), .Q(sreg[287]) );
  DFF \sreg_reg[286]  ( .D(c[288]), .CLK(clk), .RST(rst), .Q(sreg[286]) );
  DFF \sreg_reg[285]  ( .D(c[287]), .CLK(clk), .RST(rst), .Q(sreg[285]) );
  DFF \sreg_reg[284]  ( .D(c[286]), .CLK(clk), .RST(rst), .Q(sreg[284]) );
  DFF \sreg_reg[283]  ( .D(c[285]), .CLK(clk), .RST(rst), .Q(sreg[283]) );
  DFF \sreg_reg[282]  ( .D(c[284]), .CLK(clk), .RST(rst), .Q(sreg[282]) );
  DFF \sreg_reg[281]  ( .D(c[283]), .CLK(clk), .RST(rst), .Q(sreg[281]) );
  DFF \sreg_reg[280]  ( .D(c[282]), .CLK(clk), .RST(rst), .Q(sreg[280]) );
  DFF \sreg_reg[279]  ( .D(c[281]), .CLK(clk), .RST(rst), .Q(sreg[279]) );
  DFF \sreg_reg[278]  ( .D(c[280]), .CLK(clk), .RST(rst), .Q(sreg[278]) );
  DFF \sreg_reg[277]  ( .D(c[279]), .CLK(clk), .RST(rst), .Q(sreg[277]) );
  DFF \sreg_reg[276]  ( .D(c[278]), .CLK(clk), .RST(rst), .Q(sreg[276]) );
  DFF \sreg_reg[275]  ( .D(c[277]), .CLK(clk), .RST(rst), .Q(sreg[275]) );
  DFF \sreg_reg[274]  ( .D(c[276]), .CLK(clk), .RST(rst), .Q(sreg[274]) );
  DFF \sreg_reg[273]  ( .D(c[275]), .CLK(clk), .RST(rst), .Q(sreg[273]) );
  DFF \sreg_reg[272]  ( .D(c[274]), .CLK(clk), .RST(rst), .Q(sreg[272]) );
  DFF \sreg_reg[271]  ( .D(c[273]), .CLK(clk), .RST(rst), .Q(sreg[271]) );
  DFF \sreg_reg[270]  ( .D(c[272]), .CLK(clk), .RST(rst), .Q(sreg[270]) );
  DFF \sreg_reg[269]  ( .D(c[271]), .CLK(clk), .RST(rst), .Q(sreg[269]) );
  DFF \sreg_reg[268]  ( .D(c[270]), .CLK(clk), .RST(rst), .Q(sreg[268]) );
  DFF \sreg_reg[267]  ( .D(c[269]), .CLK(clk), .RST(rst), .Q(sreg[267]) );
  DFF \sreg_reg[266]  ( .D(c[268]), .CLK(clk), .RST(rst), .Q(sreg[266]) );
  DFF \sreg_reg[265]  ( .D(c[267]), .CLK(clk), .RST(rst), .Q(sreg[265]) );
  DFF \sreg_reg[264]  ( .D(c[266]), .CLK(clk), .RST(rst), .Q(sreg[264]) );
  DFF \sreg_reg[263]  ( .D(c[265]), .CLK(clk), .RST(rst), .Q(sreg[263]) );
  DFF \sreg_reg[262]  ( .D(c[264]), .CLK(clk), .RST(rst), .Q(sreg[262]) );
  DFF \sreg_reg[261]  ( .D(c[263]), .CLK(clk), .RST(rst), .Q(sreg[261]) );
  DFF \sreg_reg[260]  ( .D(c[262]), .CLK(clk), .RST(rst), .Q(sreg[260]) );
  DFF \sreg_reg[259]  ( .D(c[261]), .CLK(clk), .RST(rst), .Q(sreg[259]) );
  DFF \sreg_reg[258]  ( .D(c[260]), .CLK(clk), .RST(rst), .Q(sreg[258]) );
  DFF \sreg_reg[257]  ( .D(c[259]), .CLK(clk), .RST(rst), .Q(sreg[257]) );
  DFF \sreg_reg[256]  ( .D(c[258]), .CLK(clk), .RST(rst), .Q(sreg[256]) );
  DFF \sreg_reg[255]  ( .D(c[257]), .CLK(clk), .RST(rst), .Q(sreg[255]) );
  DFF \sreg_reg[254]  ( .D(c[256]), .CLK(clk), .RST(rst), .Q(sreg[254]) );
  DFF \sreg_reg[253]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(c[253]) );
  DFF \sreg_reg[252]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(c[252]) );
  DFF \sreg_reg[251]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(c[251]) );
  DFF \sreg_reg[250]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(c[250]) );
  DFF \sreg_reg[249]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(c[249]) );
  DFF \sreg_reg[248]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(c[248]) );
  DFF \sreg_reg[247]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(c[247]) );
  DFF \sreg_reg[246]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(c[246]) );
  DFF \sreg_reg[245]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(c[245]) );
  DFF \sreg_reg[244]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(c[244]) );
  DFF \sreg_reg[243]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(c[243]) );
  DFF \sreg_reg[242]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(c[242]) );
  DFF \sreg_reg[241]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(c[241]) );
  DFF \sreg_reg[240]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(c[240]) );
  DFF \sreg_reg[239]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(c[239]) );
  DFF \sreg_reg[238]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(c[238]) );
  DFF \sreg_reg[237]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(c[237]) );
  DFF \sreg_reg[236]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(c[236]) );
  DFF \sreg_reg[235]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(c[235]) );
  DFF \sreg_reg[234]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(c[234]) );
  DFF \sreg_reg[233]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(c[233]) );
  DFF \sreg_reg[232]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(c[232]) );
  DFF \sreg_reg[231]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(c[231]) );
  DFF \sreg_reg[230]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(c[230]) );
  DFF \sreg_reg[229]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(c[229]) );
  DFF \sreg_reg[228]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(c[228]) );
  DFF \sreg_reg[227]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(c[227]) );
  DFF \sreg_reg[226]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(c[226]) );
  DFF \sreg_reg[225]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(c[225]) );
  DFF \sreg_reg[224]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(c[224]) );
  DFF \sreg_reg[223]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(c[223]) );
  DFF \sreg_reg[222]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(c[222]) );
  DFF \sreg_reg[221]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(c[221]) );
  DFF \sreg_reg[220]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(c[220]) );
  DFF \sreg_reg[219]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(c[219]) );
  DFF \sreg_reg[218]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(c[218]) );
  DFF \sreg_reg[217]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(c[217]) );
  DFF \sreg_reg[216]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(c[216]) );
  DFF \sreg_reg[215]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(c[215]) );
  DFF \sreg_reg[214]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(c[214]) );
  DFF \sreg_reg[213]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(c[213]) );
  DFF \sreg_reg[212]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(c[212]) );
  DFF \sreg_reg[211]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(c[211]) );
  DFF \sreg_reg[210]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(c[210]) );
  DFF \sreg_reg[209]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(c[209]) );
  DFF \sreg_reg[208]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(c[208]) );
  DFF \sreg_reg[207]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(c[207]) );
  DFF \sreg_reg[206]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(c[206]) );
  DFF \sreg_reg[205]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(c[205]) );
  DFF \sreg_reg[204]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(c[204]) );
  DFF \sreg_reg[203]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(c[203]) );
  DFF \sreg_reg[202]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(c[202]) );
  DFF \sreg_reg[201]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(c[201]) );
  DFF \sreg_reg[200]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(c[200]) );
  DFF \sreg_reg[199]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(c[199]) );
  DFF \sreg_reg[198]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(c[198]) );
  DFF \sreg_reg[197]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(c[197]) );
  DFF \sreg_reg[196]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(c[196]) );
  DFF \sreg_reg[195]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(c[195]) );
  DFF \sreg_reg[194]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(c[194]) );
  DFF \sreg_reg[193]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(c[193]) );
  DFF \sreg_reg[192]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(c[192]) );
  DFF \sreg_reg[191]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(c[191]) );
  DFF \sreg_reg[190]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(c[190]) );
  DFF \sreg_reg[189]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(c[189]) );
  DFF \sreg_reg[188]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(c[188]) );
  DFF \sreg_reg[187]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(c[187]) );
  DFF \sreg_reg[186]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(c[186]) );
  DFF \sreg_reg[185]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(c[185]) );
  DFF \sreg_reg[184]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(c[184]) );
  DFF \sreg_reg[183]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(c[183]) );
  DFF \sreg_reg[182]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(c[182]) );
  DFF \sreg_reg[181]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(c[181]) );
  DFF \sreg_reg[180]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(c[180]) );
  DFF \sreg_reg[179]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(c[179]) );
  DFF \sreg_reg[178]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(c[178]) );
  DFF \sreg_reg[177]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(c[177]) );
  DFF \sreg_reg[176]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(c[176]) );
  DFF \sreg_reg[175]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(c[175]) );
  DFF \sreg_reg[174]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(c[174]) );
  DFF \sreg_reg[173]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(c[173]) );
  DFF \sreg_reg[172]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(c[172]) );
  DFF \sreg_reg[171]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(c[171]) );
  DFF \sreg_reg[170]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(c[170]) );
  DFF \sreg_reg[169]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(c[169]) );
  DFF \sreg_reg[168]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(c[168]) );
  DFF \sreg_reg[167]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(c[167]) );
  DFF \sreg_reg[166]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(c[166]) );
  DFF \sreg_reg[165]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(c[165]) );
  DFF \sreg_reg[164]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(c[164]) );
  DFF \sreg_reg[163]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(c[163]) );
  DFF \sreg_reg[162]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(c[162]) );
  DFF \sreg_reg[161]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(c[161]) );
  DFF \sreg_reg[160]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(c[160]) );
  DFF \sreg_reg[159]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(c[159]) );
  DFF \sreg_reg[158]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(c[158]) );
  DFF \sreg_reg[157]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(c[157]) );
  DFF \sreg_reg[156]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(c[156]) );
  DFF \sreg_reg[155]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(c[155]) );
  DFF \sreg_reg[154]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(c[154]) );
  DFF \sreg_reg[153]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(c[153]) );
  DFF \sreg_reg[152]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(c[152]) );
  DFF \sreg_reg[151]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(c[151]) );
  DFF \sreg_reg[150]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(c[150]) );
  DFF \sreg_reg[149]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(c[149]) );
  DFF \sreg_reg[148]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(c[148]) );
  DFF \sreg_reg[147]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(c[147]) );
  DFF \sreg_reg[146]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(c[146]) );
  DFF \sreg_reg[145]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(c[145]) );
  DFF \sreg_reg[144]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(c[144]) );
  DFF \sreg_reg[143]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(c[143]) );
  DFF \sreg_reg[142]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(c[142]) );
  DFF \sreg_reg[141]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(c[141]) );
  DFF \sreg_reg[140]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(c[140]) );
  DFF \sreg_reg[139]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(c[139]) );
  DFF \sreg_reg[138]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(c[138]) );
  DFF \sreg_reg[137]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(c[137]) );
  DFF \sreg_reg[136]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(c[136]) );
  DFF \sreg_reg[135]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(c[135]) );
  DFF \sreg_reg[134]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(c[134]) );
  DFF \sreg_reg[133]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(c[133]) );
  DFF \sreg_reg[132]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(c[132]) );
  DFF \sreg_reg[131]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(c[131]) );
  DFF \sreg_reg[130]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(c[130]) );
  DFF \sreg_reg[129]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(c[129]) );
  DFF \sreg_reg[128]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(c[128]) );
  DFF \sreg_reg[127]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(c[127]) );
  DFF \sreg_reg[126]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(c[126]) );
  DFF \sreg_reg[125]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[125]) );
  DFF \sreg_reg[124]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[124]) );
  DFF \sreg_reg[123]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[123]) );
  DFF \sreg_reg[122]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[122]) );
  DFF \sreg_reg[121]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[121]) );
  DFF \sreg_reg[120]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[120]) );
  DFF \sreg_reg[119]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[118]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[117]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[116]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[115]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[114]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[113]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[112]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[111]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[110]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[109]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[108]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[107]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[106]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[105]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[104]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[103]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[102]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[101]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[100]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[99]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[98]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[97]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[96]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[95]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[94]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[93]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[92]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[91]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[90]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[89]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[88]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[87]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[86]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[85]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[84]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[83]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[82]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[81]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[80]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[79]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[78]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[77]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[76]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[75]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[74]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[73]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[72]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[71]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[70]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[69]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[68]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[67]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[66]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[65]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[64]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[63]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[62]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[3]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[2]), .CLK(clk), .RST(rst), .Q(c[0]) );
  OR U5 ( .A(n1042), .B(n1041), .Z(n1) );
  NAND U6 ( .A(n1044), .B(n1043), .Z(n2) );
  NAND U7 ( .A(n1), .B(n2), .Z(n1051) );
  OR U8 ( .A(n1065), .B(n1064), .Z(n3) );
  NAND U9 ( .A(n1067), .B(n1066), .Z(n4) );
  NAND U10 ( .A(n3), .B(n4), .Z(n1073) );
  OR U11 ( .A(n1097), .B(n1096), .Z(n5) );
  NAND U12 ( .A(n1099), .B(n1098), .Z(n6) );
  NAND U13 ( .A(n5), .B(n6), .Z(n1105) );
  OR U14 ( .A(n1129), .B(n1128), .Z(n7) );
  NAND U15 ( .A(n1131), .B(n1130), .Z(n8) );
  NAND U16 ( .A(n7), .B(n8), .Z(n1137) );
  OR U17 ( .A(n1215), .B(n1214), .Z(n9) );
  NAND U18 ( .A(n1217), .B(n1216), .Z(n10) );
  NAND U19 ( .A(n9), .B(n10), .Z(n1223) );
  OR U20 ( .A(n1247), .B(n1246), .Z(n11) );
  NAND U21 ( .A(n1249), .B(n1248), .Z(n12) );
  NAND U22 ( .A(n11), .B(n12), .Z(n1255) );
  OR U23 ( .A(n1279), .B(n1278), .Z(n13) );
  NAND U24 ( .A(n1281), .B(n1280), .Z(n14) );
  NAND U25 ( .A(n13), .B(n14), .Z(n1287) );
  OR U26 ( .A(n1311), .B(n1310), .Z(n15) );
  NAND U27 ( .A(n1313), .B(n1312), .Z(n16) );
  NAND U28 ( .A(n15), .B(n16), .Z(n1319) );
  OR U29 ( .A(n1343), .B(n1342), .Z(n17) );
  NAND U30 ( .A(n1345), .B(n1344), .Z(n18) );
  NAND U31 ( .A(n17), .B(n18), .Z(n1352) );
  OR U32 ( .A(n1391), .B(n1390), .Z(n19) );
  NAND U33 ( .A(n1393), .B(n1392), .Z(n20) );
  NAND U34 ( .A(n19), .B(n20), .Z(n1400) );
  OR U35 ( .A(n1439), .B(n1438), .Z(n21) );
  NAND U36 ( .A(n1441), .B(n1440), .Z(n22) );
  NAND U37 ( .A(n21), .B(n22), .Z(n1447) );
  OR U38 ( .A(n1471), .B(n1470), .Z(n23) );
  NAND U39 ( .A(n1473), .B(n1472), .Z(n24) );
  NAND U40 ( .A(n23), .B(n24), .Z(n1479) );
  OR U41 ( .A(n1521), .B(n1520), .Z(n25) );
  NAND U42 ( .A(n1523), .B(n1522), .Z(n26) );
  NAND U43 ( .A(n25), .B(n26), .Z(n1529) );
  OR U44 ( .A(n1589), .B(n1588), .Z(n27) );
  NAND U45 ( .A(n1591), .B(n1590), .Z(n28) );
  NAND U46 ( .A(n27), .B(n28), .Z(n1597) );
  OR U47 ( .A(n1621), .B(n1620), .Z(n29) );
  NAND U48 ( .A(n1623), .B(n1622), .Z(n30) );
  NAND U49 ( .A(n29), .B(n30), .Z(n1629) );
  OR U50 ( .A(n1653), .B(n1652), .Z(n31) );
  NAND U51 ( .A(n1655), .B(n1654), .Z(n32) );
  NAND U52 ( .A(n31), .B(n32), .Z(n1661) );
  OR U53 ( .A(n1823), .B(n1822), .Z(n33) );
  NAND U54 ( .A(n1825), .B(n1824), .Z(n34) );
  NAND U55 ( .A(n33), .B(n34), .Z(n1831) );
  OR U56 ( .A(n1855), .B(n1854), .Z(n35) );
  NAND U57 ( .A(n1857), .B(n1856), .Z(n36) );
  NAND U58 ( .A(n35), .B(n36), .Z(n1863) );
  OR U59 ( .A(n1905), .B(n1904), .Z(n37) );
  NAND U60 ( .A(n1907), .B(n1906), .Z(n38) );
  NAND U61 ( .A(n37), .B(n38), .Z(n1913) );
  OR U62 ( .A(n1937), .B(n1936), .Z(n39) );
  NAND U63 ( .A(n1939), .B(n1938), .Z(n40) );
  NAND U64 ( .A(n39), .B(n40), .Z(n1945) );
  OR U65 ( .A(n2003), .B(n2002), .Z(n41) );
  NAND U66 ( .A(n2005), .B(n2004), .Z(n42) );
  NAND U67 ( .A(n41), .B(n42), .Z(n2011) );
  OR U68 ( .A(n2104), .B(n2103), .Z(n43) );
  NAND U69 ( .A(n2106), .B(n2105), .Z(n44) );
  NAND U70 ( .A(n43), .B(n44), .Z(n2112) );
  OR U71 ( .A(n2136), .B(n2135), .Z(n45) );
  NAND U72 ( .A(n2138), .B(n2137), .Z(n46) );
  NAND U73 ( .A(n45), .B(n46), .Z(n2144) );
  OR U74 ( .A(n2204), .B(n2203), .Z(n47) );
  NAND U75 ( .A(n2206), .B(n2205), .Z(n48) );
  NAND U76 ( .A(n47), .B(n48), .Z(n2212) );
  OR U77 ( .A(n2236), .B(n2235), .Z(n49) );
  NAND U78 ( .A(n2238), .B(n2237), .Z(n50) );
  NAND U79 ( .A(n49), .B(n50), .Z(n2244) );
  OR U80 ( .A(n2312), .B(n2311), .Z(n51) );
  NAND U81 ( .A(n2314), .B(n2313), .Z(n52) );
  NAND U82 ( .A(n51), .B(n52), .Z(n2321) );
  OR U83 ( .A(n2335), .B(n2334), .Z(n53) );
  NAND U84 ( .A(n2337), .B(n2336), .Z(n54) );
  NAND U85 ( .A(n53), .B(n54), .Z(n2343) );
  OR U86 ( .A(n2367), .B(n2366), .Z(n55) );
  NAND U87 ( .A(n2369), .B(n2368), .Z(n56) );
  NAND U88 ( .A(n55), .B(n56), .Z(n2375) );
  OR U89 ( .A(n2399), .B(n2398), .Z(n57) );
  NAND U90 ( .A(n2401), .B(n2400), .Z(n58) );
  NAND U91 ( .A(n57), .B(n58), .Z(n2407) );
  OR U92 ( .A(n2449), .B(n2448), .Z(n59) );
  NAND U93 ( .A(n2451), .B(n2450), .Z(n60) );
  NAND U94 ( .A(n59), .B(n60), .Z(n2457) );
  OR U95 ( .A(n2481), .B(n2480), .Z(n61) );
  NAND U96 ( .A(n2483), .B(n2482), .Z(n62) );
  NAND U97 ( .A(n61), .B(n62), .Z(n2489) );
  OR U98 ( .A(n2513), .B(n2512), .Z(n63) );
  NAND U99 ( .A(n2515), .B(n2514), .Z(n64) );
  NAND U100 ( .A(n63), .B(n64), .Z(n2521) );
  OR U101 ( .A(n2545), .B(n2544), .Z(n65) );
  NAND U102 ( .A(n2547), .B(n2546), .Z(n66) );
  NAND U103 ( .A(n65), .B(n66), .Z(n2553) );
  OR U104 ( .A(n2577), .B(n2576), .Z(n67) );
  NAND U105 ( .A(n2579), .B(n2578), .Z(n68) );
  NAND U106 ( .A(n67), .B(n68), .Z(n2585) );
  OR U107 ( .A(n2609), .B(n2608), .Z(n69) );
  NAND U108 ( .A(n2611), .B(n2610), .Z(n70) );
  NAND U109 ( .A(n69), .B(n70), .Z(n2617) );
  OR U110 ( .A(n2641), .B(n2640), .Z(n71) );
  NAND U111 ( .A(n2643), .B(n2642), .Z(n72) );
  NAND U112 ( .A(n71), .B(n72), .Z(n2649) );
  OR U113 ( .A(n2691), .B(n2690), .Z(n73) );
  NAND U114 ( .A(n2693), .B(n2692), .Z(n74) );
  NAND U115 ( .A(n73), .B(n74), .Z(n2699) );
  OR U116 ( .A(n2723), .B(n2722), .Z(n75) );
  NAND U117 ( .A(n2725), .B(n2724), .Z(n76) );
  NAND U118 ( .A(n75), .B(n76), .Z(n2731) );
  OR U119 ( .A(n2755), .B(n2754), .Z(n77) );
  NAND U120 ( .A(n2757), .B(n2756), .Z(n78) );
  NAND U121 ( .A(n77), .B(n78), .Z(n2764) );
  OR U122 ( .A(n2787), .B(n2786), .Z(n79) );
  NAND U123 ( .A(n2789), .B(n2788), .Z(n80) );
  NAND U124 ( .A(n79), .B(n80), .Z(n2795) );
  OR U125 ( .A(n2819), .B(n2818), .Z(n81) );
  NAND U126 ( .A(n2821), .B(n2820), .Z(n82) );
  NAND U127 ( .A(n81), .B(n82), .Z(n2827) );
  OR U128 ( .A(n2851), .B(n2850), .Z(n83) );
  NAND U129 ( .A(n2853), .B(n2852), .Z(n84) );
  NAND U130 ( .A(n83), .B(n84), .Z(n2859) );
  OR U131 ( .A(n2883), .B(n2882), .Z(n85) );
  NAND U132 ( .A(n2885), .B(n2884), .Z(n86) );
  NAND U133 ( .A(n85), .B(n86), .Z(n2891) );
  OR U134 ( .A(n2925), .B(n2924), .Z(n87) );
  NAND U135 ( .A(n2927), .B(n2926), .Z(n88) );
  NAND U136 ( .A(n87), .B(n88), .Z(n2934) );
  OR U137 ( .A(n2982), .B(n2981), .Z(n89) );
  NAND U138 ( .A(n2984), .B(n2983), .Z(n90) );
  NAND U139 ( .A(n89), .B(n90), .Z(n2990) );
  OR U140 ( .A(n3024), .B(n3023), .Z(n91) );
  NAND U141 ( .A(n3026), .B(n3025), .Z(n92) );
  NAND U142 ( .A(n91), .B(n92), .Z(n3033) );
  OR U143 ( .A(n1049), .B(n1048), .Z(n93) );
  NAND U144 ( .A(n1051), .B(n1050), .Z(n94) );
  NAND U145 ( .A(n93), .B(n94), .Z(n1057) );
  OR U146 ( .A(n1081), .B(n1080), .Z(n95) );
  NAND U147 ( .A(n1083), .B(n1082), .Z(n96) );
  NAND U148 ( .A(n95), .B(n96), .Z(n1089) );
  OR U149 ( .A(n1113), .B(n1112), .Z(n97) );
  NAND U150 ( .A(n1115), .B(n1114), .Z(n98) );
  NAND U151 ( .A(n97), .B(n98), .Z(n1121) );
  OR U152 ( .A(n1145), .B(n1144), .Z(n99) );
  NAND U153 ( .A(n1147), .B(n1146), .Z(n100) );
  NAND U154 ( .A(n99), .B(n100), .Z(n1153) );
  OR U155 ( .A(n1181), .B(n1180), .Z(n101) );
  NAND U156 ( .A(n1183), .B(n1182), .Z(n102) );
  NAND U157 ( .A(n101), .B(n102), .Z(n1189) );
  OR U158 ( .A(n1231), .B(n1230), .Z(n103) );
  NAND U159 ( .A(n1233), .B(n1232), .Z(n104) );
  NAND U160 ( .A(n103), .B(n104), .Z(n1239) );
  OR U161 ( .A(n1263), .B(n1262), .Z(n105) );
  NAND U162 ( .A(n1265), .B(n1264), .Z(n106) );
  NAND U163 ( .A(n105), .B(n106), .Z(n1271) );
  OR U164 ( .A(n1295), .B(n1294), .Z(n107) );
  NAND U165 ( .A(n1297), .B(n1296), .Z(n108) );
  NAND U166 ( .A(n107), .B(n108), .Z(n1303) );
  OR U167 ( .A(n1327), .B(n1326), .Z(n109) );
  NAND U168 ( .A(n1329), .B(n1328), .Z(n110) );
  NAND U169 ( .A(n109), .B(n110), .Z(n1335) );
  OR U170 ( .A(n1350), .B(n1349), .Z(n111) );
  NAND U171 ( .A(n1352), .B(n1351), .Z(n112) );
  NAND U172 ( .A(n111), .B(n112), .Z(n1358) );
  OR U173 ( .A(n1375), .B(n1374), .Z(n113) );
  NAND U174 ( .A(n1377), .B(n1376), .Z(n114) );
  NAND U175 ( .A(n113), .B(n114), .Z(n1383) );
  OR U176 ( .A(n1398), .B(n1397), .Z(n115) );
  NAND U177 ( .A(n1400), .B(n1399), .Z(n116) );
  NAND U178 ( .A(n115), .B(n116), .Z(n1406) );
  OR U179 ( .A(n1423), .B(n1422), .Z(n117) );
  NAND U180 ( .A(n1425), .B(n1424), .Z(n118) );
  NAND U181 ( .A(n117), .B(n118), .Z(n1431) );
  OR U182 ( .A(n1455), .B(n1454), .Z(n119) );
  NAND U183 ( .A(n1457), .B(n1456), .Z(n120) );
  NAND U184 ( .A(n119), .B(n120), .Z(n1463) );
  OR U185 ( .A(n1487), .B(n1486), .Z(n121) );
  NAND U186 ( .A(n1489), .B(n1488), .Z(n122) );
  NAND U187 ( .A(n121), .B(n122), .Z(n1495) );
  OR U188 ( .A(n1537), .B(n1536), .Z(n123) );
  NAND U189 ( .A(n1539), .B(n1538), .Z(n124) );
  NAND U190 ( .A(n123), .B(n124), .Z(n1545) );
  OR U191 ( .A(n1605), .B(n1604), .Z(n125) );
  NAND U192 ( .A(n1607), .B(n1606), .Z(n126) );
  NAND U193 ( .A(n125), .B(n126), .Z(n1613) );
  OR U194 ( .A(n1637), .B(n1636), .Z(n127) );
  NAND U195 ( .A(n1639), .B(n1638), .Z(n128) );
  NAND U196 ( .A(n127), .B(n128), .Z(n1645) );
  OR U197 ( .A(n1669), .B(n1668), .Z(n129) );
  NAND U198 ( .A(n1671), .B(n1670), .Z(n130) );
  NAND U199 ( .A(n129), .B(n130), .Z(n1677) );
  OR U200 ( .A(n1703), .B(n1702), .Z(n131) );
  NAND U201 ( .A(n1705), .B(n1704), .Z(n132) );
  NAND U202 ( .A(n131), .B(n132), .Z(n1711) );
  OR U203 ( .A(n1737), .B(n1736), .Z(n133) );
  NAND U204 ( .A(n1739), .B(n1738), .Z(n134) );
  NAND U205 ( .A(n133), .B(n134), .Z(n1745) );
  OR U206 ( .A(n1807), .B(n1806), .Z(n135) );
  NAND U207 ( .A(n1809), .B(n1808), .Z(n136) );
  NAND U208 ( .A(n135), .B(n136), .Z(n1815) );
  OR U209 ( .A(n1839), .B(n1838), .Z(n137) );
  NAND U210 ( .A(n1841), .B(n1840), .Z(n138) );
  NAND U211 ( .A(n137), .B(n138), .Z(n1847) );
  OR U212 ( .A(n1871), .B(n1870), .Z(n139) );
  NAND U213 ( .A(n1873), .B(n1872), .Z(n140) );
  NAND U214 ( .A(n139), .B(n140), .Z(n1879) );
  OR U215 ( .A(n1921), .B(n1920), .Z(n141) );
  NAND U216 ( .A(n1923), .B(n1922), .Z(n142) );
  NAND U217 ( .A(n141), .B(n142), .Z(n1929) );
  OR U218 ( .A(n1953), .B(n1952), .Z(n143) );
  NAND U219 ( .A(n1955), .B(n1954), .Z(n144) );
  NAND U220 ( .A(n143), .B(n144), .Z(n1961) );
  OR U221 ( .A(n1987), .B(n1986), .Z(n145) );
  NAND U222 ( .A(n1989), .B(n1988), .Z(n146) );
  NAND U223 ( .A(n145), .B(n146), .Z(n1995) );
  OR U224 ( .A(n2019), .B(n2018), .Z(n147) );
  NAND U225 ( .A(n2021), .B(n2020), .Z(n148) );
  NAND U226 ( .A(n147), .B(n148), .Z(n2027) );
  OR U227 ( .A(n2053), .B(n2052), .Z(n149) );
  NAND U228 ( .A(n2055), .B(n2054), .Z(n150) );
  NAND U229 ( .A(n149), .B(n150), .Z(n2061) );
  OR U230 ( .A(n2097), .B(n2096), .Z(n151) );
  NAND U231 ( .A(n2099), .B(n2098), .Z(n152) );
  NAND U232 ( .A(n151), .B(n152), .Z(n2106) );
  OR U233 ( .A(n2120), .B(n2119), .Z(n153) );
  NAND U234 ( .A(n2122), .B(n2121), .Z(n154) );
  NAND U235 ( .A(n153), .B(n154), .Z(n2128) );
  OR U236 ( .A(n2152), .B(n2151), .Z(n155) );
  NAND U237 ( .A(n2154), .B(n2153), .Z(n156) );
  NAND U238 ( .A(n155), .B(n156), .Z(n2160) );
  OR U239 ( .A(n2220), .B(n2219), .Z(n157) );
  NAND U240 ( .A(n2222), .B(n2221), .Z(n158) );
  NAND U241 ( .A(n157), .B(n158), .Z(n2228) );
  OR U242 ( .A(n2252), .B(n2251), .Z(n159) );
  NAND U243 ( .A(n2254), .B(n2253), .Z(n160) );
  NAND U244 ( .A(n159), .B(n160), .Z(n2260) );
  OR U245 ( .A(n2286), .B(n2285), .Z(n161) );
  NAND U246 ( .A(n2288), .B(n2287), .Z(n162) );
  NAND U247 ( .A(n161), .B(n162), .Z(n2294) );
  OR U248 ( .A(n2319), .B(n2318), .Z(n163) );
  NAND U249 ( .A(n2321), .B(n2320), .Z(n164) );
  NAND U250 ( .A(n163), .B(n164), .Z(n2327) );
  OR U251 ( .A(n2351), .B(n2350), .Z(n165) );
  NAND U252 ( .A(n2353), .B(n2352), .Z(n166) );
  NAND U253 ( .A(n165), .B(n166), .Z(n2359) );
  OR U254 ( .A(n2383), .B(n2382), .Z(n167) );
  NAND U255 ( .A(n2385), .B(n2384), .Z(n168) );
  NAND U256 ( .A(n167), .B(n168), .Z(n2391) );
  OR U257 ( .A(n2415), .B(n2414), .Z(n169) );
  NAND U258 ( .A(n2417), .B(n2416), .Z(n170) );
  NAND U259 ( .A(n169), .B(n170), .Z(n2423) );
  OR U260 ( .A(n2465), .B(n2464), .Z(n171) );
  NAND U261 ( .A(n2467), .B(n2466), .Z(n172) );
  NAND U262 ( .A(n171), .B(n172), .Z(n2473) );
  OR U263 ( .A(n2497), .B(n2496), .Z(n173) );
  NAND U264 ( .A(n2499), .B(n2498), .Z(n174) );
  NAND U265 ( .A(n173), .B(n174), .Z(n2505) );
  OR U266 ( .A(n2529), .B(n2528), .Z(n175) );
  NAND U267 ( .A(n2531), .B(n2530), .Z(n176) );
  NAND U268 ( .A(n175), .B(n176), .Z(n2537) );
  OR U269 ( .A(n2561), .B(n2560), .Z(n177) );
  NAND U270 ( .A(n2563), .B(n2562), .Z(n178) );
  NAND U271 ( .A(n177), .B(n178), .Z(n2569) );
  OR U272 ( .A(n2593), .B(n2592), .Z(n179) );
  NAND U273 ( .A(n2595), .B(n2594), .Z(n180) );
  NAND U274 ( .A(n179), .B(n180), .Z(n2601) );
  OR U275 ( .A(n2625), .B(n2624), .Z(n181) );
  NAND U276 ( .A(n2627), .B(n2626), .Z(n182) );
  NAND U277 ( .A(n181), .B(n182), .Z(n2633) );
  OR U278 ( .A(n2657), .B(n2656), .Z(n183) );
  NAND U279 ( .A(n2659), .B(n2658), .Z(n184) );
  NAND U280 ( .A(n183), .B(n184), .Z(n2665) );
  OR U281 ( .A(n2707), .B(n2706), .Z(n185) );
  NAND U282 ( .A(n2709), .B(n2708), .Z(n186) );
  NAND U283 ( .A(n185), .B(n186), .Z(n2715) );
  OR U284 ( .A(n2739), .B(n2738), .Z(n187) );
  NAND U285 ( .A(n2741), .B(n2740), .Z(n188) );
  NAND U286 ( .A(n187), .B(n188), .Z(n2747) );
  OR U287 ( .A(n2762), .B(n2761), .Z(n189) );
  NAND U288 ( .A(n2764), .B(n2763), .Z(n190) );
  NAND U289 ( .A(n189), .B(n190), .Z(n2770) );
  OR U290 ( .A(n2803), .B(n2802), .Z(n191) );
  NAND U291 ( .A(n2805), .B(n2804), .Z(n192) );
  NAND U292 ( .A(n191), .B(n192), .Z(n2811) );
  OR U293 ( .A(n2835), .B(n2834), .Z(n193) );
  NAND U294 ( .A(n2837), .B(n2836), .Z(n194) );
  NAND U295 ( .A(n193), .B(n194), .Z(n2843) );
  OR U296 ( .A(n2867), .B(n2866), .Z(n195) );
  NAND U297 ( .A(n2869), .B(n2868), .Z(n196) );
  NAND U298 ( .A(n195), .B(n196), .Z(n2875) );
  OR U299 ( .A(n2899), .B(n2898), .Z(n197) );
  NAND U300 ( .A(n2901), .B(n2900), .Z(n198) );
  NAND U301 ( .A(n197), .B(n198), .Z(n2907) );
  OR U302 ( .A(n2932), .B(n2931), .Z(n199) );
  NAND U303 ( .A(n2934), .B(n2933), .Z(n200) );
  NAND U304 ( .A(n199), .B(n200), .Z(n2940) );
  OR U305 ( .A(n2966), .B(n2965), .Z(n201) );
  NAND U306 ( .A(n2968), .B(n2967), .Z(n202) );
  NAND U307 ( .A(n201), .B(n202), .Z(n2974) );
  OR U308 ( .A(n2998), .B(n2997), .Z(n203) );
  NAND U309 ( .A(n3000), .B(n2999), .Z(n204) );
  NAND U310 ( .A(n203), .B(n204), .Z(n3006) );
  OR U311 ( .A(n3031), .B(n3030), .Z(n205) );
  NAND U312 ( .A(n3033), .B(n3032), .Z(n206) );
  NAND U313 ( .A(n205), .B(n206), .Z(n3039) );
  NAND U314 ( .A(n1165), .B(sreg[278]), .Z(n207) );
  XOR U315 ( .A(sreg[278]), .B(n1165), .Z(n208) );
  NANDN U316 ( .A(n1164), .B(n208), .Z(n209) );
  NAND U317 ( .A(n207), .B(n209), .Z(n1174) );
  NAND U318 ( .A(n992), .B(sreg[257]), .Z(n210) );
  XOR U319 ( .A(sreg[257]), .B(n992), .Z(n211) );
  NANDN U320 ( .A(n991), .B(n211), .Z(n212) );
  NAND U321 ( .A(n210), .B(n212), .Z(n1000) );
  NAND U322 ( .A(n1022), .B(sreg[260]), .Z(n213) );
  XOR U323 ( .A(sreg[260]), .B(n1022), .Z(n214) );
  NANDN U324 ( .A(n1021), .B(n214), .Z(n215) );
  NAND U325 ( .A(n213), .B(n215), .Z(n1029) );
  NAND U326 ( .A(n1046), .B(sreg[263]), .Z(n216) );
  XOR U327 ( .A(sreg[263]), .B(n1046), .Z(n217) );
  NANDN U328 ( .A(n1045), .B(n217), .Z(n218) );
  NAND U329 ( .A(n216), .B(n218), .Z(n1052) );
  NAND U330 ( .A(n1069), .B(sreg[266]), .Z(n219) );
  XOR U331 ( .A(sreg[266]), .B(n1069), .Z(n220) );
  NANDN U332 ( .A(n1068), .B(n220), .Z(n221) );
  NAND U333 ( .A(n219), .B(n221), .Z(n1077) );
  XOR U334 ( .A(n1093), .B(sreg[269]), .Z(n222) );
  NANDN U335 ( .A(n1094), .B(n222), .Z(n223) );
  NAND U336 ( .A(n1093), .B(sreg[269]), .Z(n224) );
  AND U337 ( .A(n223), .B(n224), .Z(n1100) );
  NAND U338 ( .A(n1117), .B(sreg[272]), .Z(n225) );
  XOR U339 ( .A(sreg[272]), .B(n1117), .Z(n226) );
  NANDN U340 ( .A(n1116), .B(n226), .Z(n227) );
  NAND U341 ( .A(n225), .B(n227), .Z(n1125) );
  XOR U342 ( .A(n1141), .B(sreg[275]), .Z(n228) );
  NANDN U343 ( .A(n1142), .B(n228), .Z(n229) );
  NAND U344 ( .A(n1141), .B(sreg[275]), .Z(n230) );
  AND U345 ( .A(n229), .B(n230), .Z(n1148) );
  XOR U346 ( .A(n1202), .B(n1203), .Z(n231) );
  NANDN U347 ( .A(sreg[282]), .B(n231), .Z(n232) );
  NAND U348 ( .A(n1202), .B(n1203), .Z(n233) );
  AND U349 ( .A(n232), .B(n233), .Z(n1211) );
  XOR U350 ( .A(n1227), .B(sreg[285]), .Z(n234) );
  NANDN U351 ( .A(n1228), .B(n234), .Z(n235) );
  NAND U352 ( .A(n1227), .B(sreg[285]), .Z(n236) );
  AND U353 ( .A(n235), .B(n236), .Z(n1234) );
  NAND U354 ( .A(n1251), .B(sreg[288]), .Z(n237) );
  XOR U355 ( .A(sreg[288]), .B(n1251), .Z(n238) );
  NANDN U356 ( .A(n1250), .B(n238), .Z(n239) );
  NAND U357 ( .A(n237), .B(n239), .Z(n1259) );
  XOR U358 ( .A(n1275), .B(sreg[291]), .Z(n240) );
  NANDN U359 ( .A(n1276), .B(n240), .Z(n241) );
  NAND U360 ( .A(n1275), .B(sreg[291]), .Z(n242) );
  AND U361 ( .A(n241), .B(n242), .Z(n1282) );
  NAND U362 ( .A(n1299), .B(sreg[294]), .Z(n243) );
  XOR U363 ( .A(sreg[294]), .B(n1299), .Z(n244) );
  NANDN U364 ( .A(n1298), .B(n244), .Z(n245) );
  NAND U365 ( .A(n243), .B(n245), .Z(n1307) );
  XOR U366 ( .A(n1323), .B(sreg[297]), .Z(n246) );
  NANDN U367 ( .A(n1324), .B(n246), .Z(n247) );
  NAND U368 ( .A(n1323), .B(sreg[297]), .Z(n248) );
  AND U369 ( .A(n247), .B(n248), .Z(n1330) );
  NAND U370 ( .A(n1347), .B(sreg[300]), .Z(n249) );
  XOR U371 ( .A(sreg[300]), .B(n1347), .Z(n250) );
  NANDN U372 ( .A(n1346), .B(n250), .Z(n251) );
  NAND U373 ( .A(n249), .B(n251), .Z(n1353) );
  XOR U374 ( .A(n1371), .B(sreg[303]), .Z(n252) );
  NANDN U375 ( .A(n1372), .B(n252), .Z(n253) );
  NAND U376 ( .A(n1371), .B(sreg[303]), .Z(n254) );
  AND U377 ( .A(n253), .B(n254), .Z(n1378) );
  NAND U378 ( .A(n1395), .B(sreg[306]), .Z(n255) );
  XOR U379 ( .A(sreg[306]), .B(n1395), .Z(n256) );
  NANDN U380 ( .A(n1394), .B(n256), .Z(n257) );
  NAND U381 ( .A(n255), .B(n257), .Z(n1401) );
  XOR U382 ( .A(n1419), .B(sreg[309]), .Z(n258) );
  NANDN U383 ( .A(n1420), .B(n258), .Z(n259) );
  NAND U384 ( .A(n1419), .B(sreg[309]), .Z(n260) );
  AND U385 ( .A(n259), .B(n260), .Z(n1426) );
  NAND U386 ( .A(n1443), .B(sreg[312]), .Z(n261) );
  XOR U387 ( .A(sreg[312]), .B(n1443), .Z(n262) );
  NANDN U388 ( .A(n1442), .B(n262), .Z(n263) );
  NAND U389 ( .A(n261), .B(n263), .Z(n1451) );
  XOR U390 ( .A(n1467), .B(sreg[315]), .Z(n264) );
  NANDN U391 ( .A(n1468), .B(n264), .Z(n265) );
  NAND U392 ( .A(n1467), .B(sreg[315]), .Z(n266) );
  AND U393 ( .A(n265), .B(n266), .Z(n1474) );
  NAND U394 ( .A(n1491), .B(sreg[318]), .Z(n267) );
  XOR U395 ( .A(sreg[318]), .B(n1491), .Z(n268) );
  NANDN U396 ( .A(n1490), .B(n268), .Z(n269) );
  NAND U397 ( .A(n267), .B(n269), .Z(n1499) );
  XOR U398 ( .A(n1517), .B(sreg[321]), .Z(n270) );
  NANDN U399 ( .A(n1518), .B(n270), .Z(n271) );
  NAND U400 ( .A(n1517), .B(sreg[321]), .Z(n272) );
  AND U401 ( .A(n271), .B(n272), .Z(n1524) );
  NAND U402 ( .A(n1541), .B(sreg[324]), .Z(n273) );
  XOR U403 ( .A(sreg[324]), .B(n1541), .Z(n274) );
  NANDN U404 ( .A(n1540), .B(n274), .Z(n275) );
  NAND U405 ( .A(n273), .B(n275), .Z(n1549) );
  NAND U406 ( .A(n1567), .B(sreg[327]), .Z(n276) );
  XOR U407 ( .A(sreg[327]), .B(n1567), .Z(n277) );
  NANDN U408 ( .A(n1568), .B(n277), .Z(n278) );
  NAND U409 ( .A(n276), .B(n278), .Z(n1576) );
  NAND U410 ( .A(n1593), .B(sreg[330]), .Z(n279) );
  XOR U411 ( .A(sreg[330]), .B(n1593), .Z(n280) );
  NANDN U412 ( .A(n1592), .B(n280), .Z(n281) );
  NAND U413 ( .A(n279), .B(n281), .Z(n1601) );
  XOR U414 ( .A(n1617), .B(sreg[333]), .Z(n282) );
  NANDN U415 ( .A(n1618), .B(n282), .Z(n283) );
  NAND U416 ( .A(n1617), .B(sreg[333]), .Z(n284) );
  AND U417 ( .A(n283), .B(n284), .Z(n1624) );
  NAND U418 ( .A(n1641), .B(sreg[336]), .Z(n285) );
  XOR U419 ( .A(sreg[336]), .B(n1641), .Z(n286) );
  NANDN U420 ( .A(n1640), .B(n286), .Z(n287) );
  NAND U421 ( .A(n285), .B(n287), .Z(n1649) );
  XOR U422 ( .A(n1665), .B(sreg[339]), .Z(n288) );
  NANDN U423 ( .A(n1666), .B(n288), .Z(n289) );
  NAND U424 ( .A(n1665), .B(sreg[339]), .Z(n290) );
  AND U425 ( .A(n289), .B(n290), .Z(n1672) );
  NAND U426 ( .A(n1690), .B(sreg[342]), .Z(n291) );
  XOR U427 ( .A(sreg[342]), .B(n1690), .Z(n292) );
  NANDN U428 ( .A(n1691), .B(n292), .Z(n293) );
  NAND U429 ( .A(n291), .B(n293), .Z(n1699) );
  NAND U430 ( .A(n1715), .B(sreg[345]), .Z(n294) );
  XOR U431 ( .A(sreg[345]), .B(n1715), .Z(n295) );
  NANDN U432 ( .A(n1716), .B(n295), .Z(n296) );
  NAND U433 ( .A(n294), .B(n296), .Z(n1724) );
  NAND U434 ( .A(n1741), .B(sreg[348]), .Z(n297) );
  XOR U435 ( .A(sreg[348]), .B(n1741), .Z(n298) );
  NANDN U436 ( .A(n1740), .B(n298), .Z(n299) );
  NAND U437 ( .A(n297), .B(n299), .Z(n1749) );
  NAND U438 ( .A(n1767), .B(sreg[351]), .Z(n300) );
  XOR U439 ( .A(sreg[351]), .B(n1767), .Z(n301) );
  NANDN U440 ( .A(n1768), .B(n301), .Z(n302) );
  NAND U441 ( .A(n300), .B(n302), .Z(n1776) );
  NAND U442 ( .A(n1794), .B(sreg[354]), .Z(n303) );
  XOR U443 ( .A(sreg[354]), .B(n1794), .Z(n304) );
  NANDN U444 ( .A(n1795), .B(n304), .Z(n305) );
  NAND U445 ( .A(n303), .B(n305), .Z(n1803) );
  XOR U446 ( .A(n1819), .B(sreg[357]), .Z(n306) );
  NANDN U447 ( .A(n1820), .B(n306), .Z(n307) );
  NAND U448 ( .A(n1819), .B(sreg[357]), .Z(n308) );
  AND U449 ( .A(n307), .B(n308), .Z(n1826) );
  NAND U450 ( .A(n1843), .B(sreg[360]), .Z(n309) );
  XOR U451 ( .A(sreg[360]), .B(n1843), .Z(n310) );
  NANDN U452 ( .A(n1842), .B(n310), .Z(n311) );
  NAND U453 ( .A(n309), .B(n311), .Z(n1851) );
  XOR U454 ( .A(n1867), .B(sreg[363]), .Z(n312) );
  NANDN U455 ( .A(n1868), .B(n312), .Z(n313) );
  NAND U456 ( .A(n1867), .B(sreg[363]), .Z(n314) );
  AND U457 ( .A(n313), .B(n314), .Z(n1874) );
  NAND U458 ( .A(n1892), .B(sreg[366]), .Z(n315) );
  XOR U459 ( .A(sreg[366]), .B(n1892), .Z(n316) );
  NANDN U460 ( .A(n1893), .B(n316), .Z(n317) );
  NAND U461 ( .A(n315), .B(n317), .Z(n1901) );
  XOR U462 ( .A(n1917), .B(sreg[369]), .Z(n318) );
  NANDN U463 ( .A(n1918), .B(n318), .Z(n319) );
  NAND U464 ( .A(n1917), .B(sreg[369]), .Z(n320) );
  AND U465 ( .A(n319), .B(n320), .Z(n1924) );
  NAND U466 ( .A(n1941), .B(sreg[372]), .Z(n321) );
  XOR U467 ( .A(sreg[372]), .B(n1941), .Z(n322) );
  NANDN U468 ( .A(n1940), .B(n322), .Z(n323) );
  NAND U469 ( .A(n321), .B(n323), .Z(n1949) );
  NAND U470 ( .A(n1965), .B(sreg[375]), .Z(n324) );
  XOR U471 ( .A(sreg[375]), .B(n1965), .Z(n325) );
  NANDN U472 ( .A(n1966), .B(n325), .Z(n326) );
  NAND U473 ( .A(n324), .B(n326), .Z(n1974) );
  NAND U474 ( .A(n1991), .B(sreg[378]), .Z(n327) );
  XOR U475 ( .A(sreg[378]), .B(n1991), .Z(n328) );
  NANDN U476 ( .A(n1990), .B(n328), .Z(n329) );
  NAND U477 ( .A(n327), .B(n329), .Z(n1999) );
  XOR U478 ( .A(n2015), .B(sreg[381]), .Z(n330) );
  NANDN U479 ( .A(n2016), .B(n330), .Z(n331) );
  NAND U480 ( .A(n2015), .B(sreg[381]), .Z(n332) );
  AND U481 ( .A(n331), .B(n332), .Z(n2022) );
  NAND U482 ( .A(n2040), .B(sreg[384]), .Z(n333) );
  XOR U483 ( .A(sreg[384]), .B(n2040), .Z(n334) );
  NANDN U484 ( .A(n2041), .B(n334), .Z(n335) );
  NAND U485 ( .A(n333), .B(n335), .Z(n2049) );
  NAND U486 ( .A(n2065), .B(sreg[387]), .Z(n336) );
  XOR U487 ( .A(sreg[387]), .B(n2065), .Z(n337) );
  NANDN U488 ( .A(n2066), .B(n337), .Z(n338) );
  NAND U489 ( .A(n336), .B(n338), .Z(n2074) );
  NAND U490 ( .A(n2094), .B(sreg[390]), .Z(n339) );
  XOR U491 ( .A(sreg[390]), .B(n2094), .Z(n340) );
  NANDN U492 ( .A(n2093), .B(n340), .Z(n341) );
  NAND U493 ( .A(n339), .B(n341), .Z(n2100) );
  XOR U494 ( .A(n2116), .B(sreg[393]), .Z(n342) );
  NANDN U495 ( .A(n2117), .B(n342), .Z(n343) );
  NAND U496 ( .A(n2116), .B(sreg[393]), .Z(n344) );
  AND U497 ( .A(n343), .B(n344), .Z(n2123) );
  NAND U498 ( .A(n2140), .B(sreg[396]), .Z(n345) );
  XOR U499 ( .A(sreg[396]), .B(n2140), .Z(n346) );
  NANDN U500 ( .A(n2139), .B(n346), .Z(n347) );
  NAND U501 ( .A(n345), .B(n347), .Z(n2148) );
  NAND U502 ( .A(n2164), .B(sreg[399]), .Z(n348) );
  XOR U503 ( .A(sreg[399]), .B(n2164), .Z(n349) );
  NANDN U504 ( .A(n2165), .B(n349), .Z(n350) );
  NAND U505 ( .A(n348), .B(n350), .Z(n2173) );
  NAND U506 ( .A(n2191), .B(sreg[402]), .Z(n351) );
  XOR U507 ( .A(sreg[402]), .B(n2191), .Z(n352) );
  NANDN U508 ( .A(n2192), .B(n352), .Z(n353) );
  NAND U509 ( .A(n351), .B(n353), .Z(n2200) );
  XOR U510 ( .A(n2216), .B(sreg[405]), .Z(n354) );
  NANDN U511 ( .A(n2217), .B(n354), .Z(n355) );
  NAND U512 ( .A(n2216), .B(sreg[405]), .Z(n356) );
  AND U513 ( .A(n355), .B(n356), .Z(n2223) );
  NAND U514 ( .A(n2240), .B(sreg[408]), .Z(n357) );
  XOR U515 ( .A(sreg[408]), .B(n2240), .Z(n358) );
  NANDN U516 ( .A(n2239), .B(n358), .Z(n359) );
  NAND U517 ( .A(n357), .B(n359), .Z(n2248) );
  NAND U518 ( .A(n2264), .B(sreg[411]), .Z(n360) );
  XOR U519 ( .A(sreg[411]), .B(n2264), .Z(n361) );
  NANDN U520 ( .A(n2265), .B(n361), .Z(n362) );
  NAND U521 ( .A(n360), .B(n362), .Z(n2273) );
  NAND U522 ( .A(n2290), .B(sreg[414]), .Z(n363) );
  XOR U523 ( .A(sreg[414]), .B(n2290), .Z(n364) );
  NANDN U524 ( .A(n2289), .B(n364), .Z(n365) );
  NAND U525 ( .A(n363), .B(n365), .Z(n2298) );
  NAND U526 ( .A(n2316), .B(sreg[417]), .Z(n366) );
  XOR U527 ( .A(sreg[417]), .B(n2316), .Z(n367) );
  NAND U528 ( .A(n367), .B(n2315), .Z(n368) );
  NAND U529 ( .A(n366), .B(n368), .Z(n2322) );
  NAND U530 ( .A(n2339), .B(sreg[420]), .Z(n369) );
  XOR U531 ( .A(sreg[420]), .B(n2339), .Z(n370) );
  NANDN U532 ( .A(n2338), .B(n370), .Z(n371) );
  NAND U533 ( .A(n369), .B(n371), .Z(n2347) );
  XOR U534 ( .A(n2363), .B(sreg[423]), .Z(n372) );
  NANDN U535 ( .A(n2364), .B(n372), .Z(n373) );
  NAND U536 ( .A(n2363), .B(sreg[423]), .Z(n374) );
  AND U537 ( .A(n373), .B(n374), .Z(n2370) );
  NAND U538 ( .A(n2387), .B(sreg[426]), .Z(n375) );
  XOR U539 ( .A(sreg[426]), .B(n2387), .Z(n376) );
  NANDN U540 ( .A(n2386), .B(n376), .Z(n377) );
  NAND U541 ( .A(n375), .B(n377), .Z(n2395) );
  XOR U542 ( .A(n2411), .B(sreg[429]), .Z(n378) );
  NANDN U543 ( .A(n2412), .B(n378), .Z(n379) );
  NAND U544 ( .A(n2411), .B(sreg[429]), .Z(n380) );
  AND U545 ( .A(n379), .B(n380), .Z(n2418) );
  NAND U546 ( .A(n2436), .B(sreg[432]), .Z(n381) );
  XOR U547 ( .A(sreg[432]), .B(n2436), .Z(n382) );
  NANDN U548 ( .A(n2437), .B(n382), .Z(n383) );
  NAND U549 ( .A(n381), .B(n383), .Z(n2445) );
  XOR U550 ( .A(n2461), .B(sreg[435]), .Z(n384) );
  NANDN U551 ( .A(n2462), .B(n384), .Z(n385) );
  NAND U552 ( .A(n2461), .B(sreg[435]), .Z(n386) );
  AND U553 ( .A(n385), .B(n386), .Z(n2468) );
  NAND U554 ( .A(n2485), .B(sreg[438]), .Z(n387) );
  XOR U555 ( .A(sreg[438]), .B(n2485), .Z(n388) );
  NANDN U556 ( .A(n2484), .B(n388), .Z(n389) );
  NAND U557 ( .A(n387), .B(n389), .Z(n2493) );
  XOR U558 ( .A(n2509), .B(sreg[441]), .Z(n390) );
  NANDN U559 ( .A(n2510), .B(n390), .Z(n391) );
  NAND U560 ( .A(n2509), .B(sreg[441]), .Z(n392) );
  AND U561 ( .A(n391), .B(n392), .Z(n2516) );
  NAND U562 ( .A(n2533), .B(sreg[444]), .Z(n393) );
  XOR U563 ( .A(sreg[444]), .B(n2533), .Z(n394) );
  NANDN U564 ( .A(n2532), .B(n394), .Z(n395) );
  NAND U565 ( .A(n393), .B(n395), .Z(n2541) );
  XOR U566 ( .A(n2557), .B(sreg[447]), .Z(n396) );
  NANDN U567 ( .A(n2558), .B(n396), .Z(n397) );
  NAND U568 ( .A(n2557), .B(sreg[447]), .Z(n398) );
  AND U569 ( .A(n397), .B(n398), .Z(n2564) );
  NAND U570 ( .A(n2581), .B(sreg[450]), .Z(n399) );
  XOR U571 ( .A(sreg[450]), .B(n2581), .Z(n400) );
  NANDN U572 ( .A(n2580), .B(n400), .Z(n401) );
  NAND U573 ( .A(n399), .B(n401), .Z(n2589) );
  XOR U574 ( .A(n2605), .B(sreg[453]), .Z(n402) );
  NANDN U575 ( .A(n2606), .B(n402), .Z(n403) );
  NAND U576 ( .A(n2605), .B(sreg[453]), .Z(n404) );
  AND U577 ( .A(n403), .B(n404), .Z(n2612) );
  NAND U578 ( .A(n2629), .B(sreg[456]), .Z(n405) );
  XOR U579 ( .A(sreg[456]), .B(n2629), .Z(n406) );
  NANDN U580 ( .A(n2628), .B(n406), .Z(n407) );
  NAND U581 ( .A(n405), .B(n407), .Z(n2637) );
  XOR U582 ( .A(n2653), .B(sreg[459]), .Z(n408) );
  NANDN U583 ( .A(n2654), .B(n408), .Z(n409) );
  NAND U584 ( .A(n2653), .B(sreg[459]), .Z(n410) );
  AND U585 ( .A(n409), .B(n410), .Z(n2660) );
  NAND U586 ( .A(n2678), .B(sreg[462]), .Z(n411) );
  XOR U587 ( .A(sreg[462]), .B(n2678), .Z(n412) );
  NANDN U588 ( .A(n2679), .B(n412), .Z(n413) );
  NAND U589 ( .A(n411), .B(n413), .Z(n2687) );
  XOR U590 ( .A(n2703), .B(sreg[465]), .Z(n414) );
  NANDN U591 ( .A(n2704), .B(n414), .Z(n415) );
  NAND U592 ( .A(n2703), .B(sreg[465]), .Z(n416) );
  AND U593 ( .A(n415), .B(n416), .Z(n2710) );
  NAND U594 ( .A(n2727), .B(sreg[468]), .Z(n417) );
  XOR U595 ( .A(sreg[468]), .B(n2727), .Z(n418) );
  NANDN U596 ( .A(n2726), .B(n418), .Z(n419) );
  NAND U597 ( .A(n417), .B(n419), .Z(n2735) );
  XOR U598 ( .A(n2751), .B(sreg[471]), .Z(n420) );
  NANDN U599 ( .A(n2752), .B(n420), .Z(n421) );
  NAND U600 ( .A(n2751), .B(sreg[471]), .Z(n422) );
  AND U601 ( .A(n421), .B(n422), .Z(n2758) );
  NAND U602 ( .A(n2774), .B(sreg[474]), .Z(n423) );
  XOR U603 ( .A(sreg[474]), .B(n2774), .Z(n424) );
  NANDN U604 ( .A(n2775), .B(n424), .Z(n425) );
  NAND U605 ( .A(n423), .B(n425), .Z(n2783) );
  XOR U606 ( .A(n2799), .B(sreg[477]), .Z(n426) );
  NANDN U607 ( .A(n2800), .B(n426), .Z(n427) );
  NAND U608 ( .A(n2799), .B(sreg[477]), .Z(n428) );
  AND U609 ( .A(n427), .B(n428), .Z(n2806) );
  NAND U610 ( .A(n2823), .B(sreg[480]), .Z(n429) );
  XOR U611 ( .A(sreg[480]), .B(n2823), .Z(n430) );
  NANDN U612 ( .A(n2822), .B(n430), .Z(n431) );
  NAND U613 ( .A(n429), .B(n431), .Z(n2831) );
  XOR U614 ( .A(n2847), .B(sreg[483]), .Z(n432) );
  NANDN U615 ( .A(n2848), .B(n432), .Z(n433) );
  NAND U616 ( .A(n2847), .B(sreg[483]), .Z(n434) );
  AND U617 ( .A(n433), .B(n434), .Z(n2854) );
  NAND U618 ( .A(n2871), .B(sreg[486]), .Z(n435) );
  XOR U619 ( .A(sreg[486]), .B(n2871), .Z(n436) );
  NANDN U620 ( .A(n2870), .B(n436), .Z(n437) );
  NAND U621 ( .A(n435), .B(n437), .Z(n2879) );
  XOR U622 ( .A(n2895), .B(sreg[489]), .Z(n438) );
  NANDN U623 ( .A(n2896), .B(n438), .Z(n439) );
  NAND U624 ( .A(n2895), .B(sreg[489]), .Z(n440) );
  AND U625 ( .A(n439), .B(n440), .Z(n2902) );
  NAND U626 ( .A(n2922), .B(sreg[492]), .Z(n441) );
  XOR U627 ( .A(sreg[492]), .B(n2922), .Z(n442) );
  NANDN U628 ( .A(n2921), .B(n442), .Z(n443) );
  NAND U629 ( .A(n441), .B(n443), .Z(n2928) );
  NAND U630 ( .A(n2944), .B(sreg[495]), .Z(n444) );
  XOR U631 ( .A(sreg[495]), .B(n2944), .Z(n445) );
  NANDN U632 ( .A(n2945), .B(n445), .Z(n446) );
  NAND U633 ( .A(n444), .B(n446), .Z(n2953) );
  NAND U634 ( .A(n2970), .B(sreg[498]), .Z(n447) );
  XOR U635 ( .A(sreg[498]), .B(n2970), .Z(n448) );
  NANDN U636 ( .A(n2969), .B(n448), .Z(n449) );
  NAND U637 ( .A(n447), .B(n449), .Z(n2978) );
  XOR U638 ( .A(n2994), .B(sreg[501]), .Z(n450) );
  NANDN U639 ( .A(n2995), .B(n450), .Z(n451) );
  NAND U640 ( .A(n2994), .B(sreg[501]), .Z(n452) );
  AND U641 ( .A(n451), .B(n452), .Z(n3001) );
  NAND U642 ( .A(n3021), .B(sreg[504]), .Z(n453) );
  XOR U643 ( .A(sreg[504]), .B(n3021), .Z(n454) );
  NANDN U644 ( .A(n3020), .B(n454), .Z(n455) );
  NAND U645 ( .A(n453), .B(n455), .Z(n3027) );
  XOR U646 ( .A(n3043), .B(sreg[507]), .Z(n456) );
  NANDN U647 ( .A(n3044), .B(n456), .Z(n457) );
  NAND U648 ( .A(n3043), .B(sreg[507]), .Z(n458) );
  AND U649 ( .A(n457), .B(n458), .Z(n3054) );
  NAND U650 ( .A(n1000), .B(sreg[258]), .Z(n459) );
  XOR U651 ( .A(sreg[258]), .B(n1000), .Z(n460) );
  NANDN U652 ( .A(n1001), .B(n460), .Z(n461) );
  NAND U653 ( .A(n459), .B(n461), .Z(n1010) );
  NAND U654 ( .A(n1030), .B(sreg[261]), .Z(n462) );
  XOR U655 ( .A(sreg[261]), .B(n1030), .Z(n463) );
  NAND U656 ( .A(n463), .B(n1029), .Z(n464) );
  NAND U657 ( .A(n462), .B(n464), .Z(n1038) );
  NAND U658 ( .A(n1053), .B(sreg[264]), .Z(n465) );
  XOR U659 ( .A(sreg[264]), .B(n1053), .Z(n466) );
  NAND U660 ( .A(n466), .B(n1052), .Z(n467) );
  NAND U661 ( .A(n465), .B(n467), .Z(n1061) );
  XOR U662 ( .A(n1077), .B(sreg[267]), .Z(n468) );
  NANDN U663 ( .A(n1078), .B(n468), .Z(n469) );
  NAND U664 ( .A(n1077), .B(sreg[267]), .Z(n470) );
  AND U665 ( .A(n469), .B(n470), .Z(n1084) );
  NAND U666 ( .A(n1101), .B(sreg[270]), .Z(n471) );
  XOR U667 ( .A(sreg[270]), .B(n1101), .Z(n472) );
  NANDN U668 ( .A(n1100), .B(n472), .Z(n473) );
  NAND U669 ( .A(n471), .B(n473), .Z(n1109) );
  XOR U670 ( .A(n1125), .B(sreg[273]), .Z(n474) );
  NANDN U671 ( .A(n1126), .B(n474), .Z(n475) );
  NAND U672 ( .A(n1125), .B(sreg[273]), .Z(n476) );
  AND U673 ( .A(n475), .B(n476), .Z(n1132) );
  NAND U674 ( .A(n1149), .B(sreg[276]), .Z(n477) );
  XOR U675 ( .A(sreg[276]), .B(n1149), .Z(n478) );
  NANDN U676 ( .A(n1148), .B(n478), .Z(n479) );
  NAND U677 ( .A(n477), .B(n479), .Z(n1157) );
  NAND U678 ( .A(n1185), .B(sreg[280]), .Z(n480) );
  XOR U679 ( .A(sreg[280]), .B(n1185), .Z(n481) );
  NAND U680 ( .A(n481), .B(n1184), .Z(n482) );
  NAND U681 ( .A(n480), .B(n482), .Z(n1193) );
  XOR U682 ( .A(n1211), .B(sreg[283]), .Z(n483) );
  NANDN U683 ( .A(n1212), .B(n483), .Z(n484) );
  NAND U684 ( .A(n1211), .B(sreg[283]), .Z(n485) );
  AND U685 ( .A(n484), .B(n485), .Z(n1218) );
  NAND U686 ( .A(n1235), .B(sreg[286]), .Z(n486) );
  XOR U687 ( .A(sreg[286]), .B(n1235), .Z(n487) );
  NANDN U688 ( .A(n1234), .B(n487), .Z(n488) );
  NAND U689 ( .A(n486), .B(n488), .Z(n1243) );
  XOR U690 ( .A(n1259), .B(sreg[289]), .Z(n489) );
  NANDN U691 ( .A(n1260), .B(n489), .Z(n490) );
  NAND U692 ( .A(n1259), .B(sreg[289]), .Z(n491) );
  AND U693 ( .A(n490), .B(n491), .Z(n1266) );
  NAND U694 ( .A(n1283), .B(sreg[292]), .Z(n492) );
  XOR U695 ( .A(sreg[292]), .B(n1283), .Z(n493) );
  NANDN U696 ( .A(n1282), .B(n493), .Z(n494) );
  NAND U697 ( .A(n492), .B(n494), .Z(n1291) );
  XOR U698 ( .A(n1307), .B(sreg[295]), .Z(n495) );
  NANDN U699 ( .A(n1308), .B(n495), .Z(n496) );
  NAND U700 ( .A(n1307), .B(sreg[295]), .Z(n497) );
  AND U701 ( .A(n496), .B(n497), .Z(n1314) );
  NAND U702 ( .A(n1331), .B(sreg[298]), .Z(n498) );
  XOR U703 ( .A(sreg[298]), .B(n1331), .Z(n499) );
  NANDN U704 ( .A(n1330), .B(n499), .Z(n500) );
  NAND U705 ( .A(n498), .B(n500), .Z(n1339) );
  NAND U706 ( .A(n1354), .B(sreg[301]), .Z(n501) );
  XOR U707 ( .A(sreg[301]), .B(n1354), .Z(n502) );
  NAND U708 ( .A(n502), .B(n1353), .Z(n503) );
  NAND U709 ( .A(n501), .B(n503), .Z(n1362) );
  NAND U710 ( .A(n1379), .B(sreg[304]), .Z(n504) );
  XOR U711 ( .A(sreg[304]), .B(n1379), .Z(n505) );
  NANDN U712 ( .A(n1378), .B(n505), .Z(n506) );
  NAND U713 ( .A(n504), .B(n506), .Z(n1387) );
  NAND U714 ( .A(n1402), .B(sreg[307]), .Z(n507) );
  XOR U715 ( .A(sreg[307]), .B(n1402), .Z(n508) );
  NAND U716 ( .A(n508), .B(n1401), .Z(n509) );
  NAND U717 ( .A(n507), .B(n509), .Z(n1410) );
  NAND U718 ( .A(n1427), .B(sreg[310]), .Z(n510) );
  XOR U719 ( .A(sreg[310]), .B(n1427), .Z(n511) );
  NANDN U720 ( .A(n1426), .B(n511), .Z(n512) );
  NAND U721 ( .A(n510), .B(n512), .Z(n1435) );
  XOR U722 ( .A(n1451), .B(sreg[313]), .Z(n513) );
  NANDN U723 ( .A(n1452), .B(n513), .Z(n514) );
  NAND U724 ( .A(n1451), .B(sreg[313]), .Z(n515) );
  AND U725 ( .A(n514), .B(n515), .Z(n1458) );
  NAND U726 ( .A(n1475), .B(sreg[316]), .Z(n516) );
  XOR U727 ( .A(sreg[316]), .B(n1475), .Z(n517) );
  NANDN U728 ( .A(n1474), .B(n517), .Z(n518) );
  NAND U729 ( .A(n516), .B(n518), .Z(n1483) );
  NAND U730 ( .A(n1499), .B(sreg[319]), .Z(n519) );
  XOR U731 ( .A(sreg[319]), .B(n1499), .Z(n520) );
  NANDN U732 ( .A(n1500), .B(n520), .Z(n521) );
  NAND U733 ( .A(n519), .B(n521), .Z(n1508) );
  NAND U734 ( .A(n1525), .B(sreg[322]), .Z(n522) );
  XOR U735 ( .A(sreg[322]), .B(n1525), .Z(n523) );
  NANDN U736 ( .A(n1524), .B(n523), .Z(n524) );
  NAND U737 ( .A(n522), .B(n524), .Z(n1533) );
  NAND U738 ( .A(n1549), .B(sreg[325]), .Z(n525) );
  XOR U739 ( .A(sreg[325]), .B(n1549), .Z(n526) );
  NANDN U740 ( .A(n1550), .B(n526), .Z(n527) );
  NAND U741 ( .A(n525), .B(n527), .Z(n1558) );
  NAND U742 ( .A(n1576), .B(sreg[328]), .Z(n528) );
  XOR U743 ( .A(sreg[328]), .B(n1576), .Z(n529) );
  NANDN U744 ( .A(n1577), .B(n529), .Z(n530) );
  NAND U745 ( .A(n528), .B(n530), .Z(n1585) );
  XOR U746 ( .A(n1601), .B(sreg[331]), .Z(n531) );
  NANDN U747 ( .A(n1602), .B(n531), .Z(n532) );
  NAND U748 ( .A(n1601), .B(sreg[331]), .Z(n533) );
  AND U749 ( .A(n532), .B(n533), .Z(n1608) );
  NAND U750 ( .A(n1625), .B(sreg[334]), .Z(n534) );
  XOR U751 ( .A(sreg[334]), .B(n1625), .Z(n535) );
  NANDN U752 ( .A(n1624), .B(n535), .Z(n536) );
  NAND U753 ( .A(n534), .B(n536), .Z(n1633) );
  XOR U754 ( .A(n1649), .B(sreg[337]), .Z(n537) );
  NANDN U755 ( .A(n1650), .B(n537), .Z(n538) );
  NAND U756 ( .A(n1649), .B(sreg[337]), .Z(n539) );
  AND U757 ( .A(n538), .B(n539), .Z(n1656) );
  NAND U758 ( .A(n1673), .B(sreg[340]), .Z(n540) );
  XOR U759 ( .A(sreg[340]), .B(n1673), .Z(n541) );
  NANDN U760 ( .A(n1672), .B(n541), .Z(n542) );
  NAND U761 ( .A(n540), .B(n542), .Z(n1681) );
  XOR U762 ( .A(n1699), .B(sreg[343]), .Z(n543) );
  NANDN U763 ( .A(n1700), .B(n543), .Z(n544) );
  NAND U764 ( .A(n1699), .B(sreg[343]), .Z(n545) );
  AND U765 ( .A(n544), .B(n545), .Z(n1706) );
  NAND U766 ( .A(n1724), .B(sreg[346]), .Z(n546) );
  XOR U767 ( .A(sreg[346]), .B(n1724), .Z(n547) );
  NANDN U768 ( .A(n1725), .B(n547), .Z(n548) );
  NAND U769 ( .A(n546), .B(n548), .Z(n1733) );
  NAND U770 ( .A(n1749), .B(sreg[349]), .Z(n549) );
  XOR U771 ( .A(sreg[349]), .B(n1749), .Z(n550) );
  NANDN U772 ( .A(n1750), .B(n550), .Z(n551) );
  NAND U773 ( .A(n549), .B(n551), .Z(n1758) );
  NAND U774 ( .A(n1776), .B(sreg[352]), .Z(n552) );
  XOR U775 ( .A(sreg[352]), .B(n1776), .Z(n553) );
  NANDN U776 ( .A(n1777), .B(n553), .Z(n554) );
  NAND U777 ( .A(n552), .B(n554), .Z(n1785) );
  XOR U778 ( .A(n1803), .B(sreg[355]), .Z(n555) );
  NANDN U779 ( .A(n1804), .B(n555), .Z(n556) );
  NAND U780 ( .A(n1803), .B(sreg[355]), .Z(n557) );
  AND U781 ( .A(n556), .B(n557), .Z(n1810) );
  NAND U782 ( .A(n1827), .B(sreg[358]), .Z(n558) );
  XOR U783 ( .A(sreg[358]), .B(n1827), .Z(n559) );
  NANDN U784 ( .A(n1826), .B(n559), .Z(n560) );
  NAND U785 ( .A(n558), .B(n560), .Z(n1835) );
  XOR U786 ( .A(n1851), .B(sreg[361]), .Z(n561) );
  NANDN U787 ( .A(n1852), .B(n561), .Z(n562) );
  NAND U788 ( .A(n1851), .B(sreg[361]), .Z(n563) );
  AND U789 ( .A(n562), .B(n563), .Z(n1858) );
  NAND U790 ( .A(n1875), .B(sreg[364]), .Z(n564) );
  XOR U791 ( .A(sreg[364]), .B(n1875), .Z(n565) );
  NANDN U792 ( .A(n1874), .B(n565), .Z(n566) );
  NAND U793 ( .A(n564), .B(n566), .Z(n1883) );
  XOR U794 ( .A(n1901), .B(sreg[367]), .Z(n567) );
  NANDN U795 ( .A(n1902), .B(n567), .Z(n568) );
  NAND U796 ( .A(n1901), .B(sreg[367]), .Z(n569) );
  AND U797 ( .A(n568), .B(n569), .Z(n1908) );
  NAND U798 ( .A(n1925), .B(sreg[370]), .Z(n570) );
  XOR U799 ( .A(sreg[370]), .B(n1925), .Z(n571) );
  NANDN U800 ( .A(n1924), .B(n571), .Z(n572) );
  NAND U801 ( .A(n570), .B(n572), .Z(n1933) );
  XOR U802 ( .A(n1949), .B(sreg[373]), .Z(n573) );
  NANDN U803 ( .A(n1950), .B(n573), .Z(n574) );
  NAND U804 ( .A(n1949), .B(sreg[373]), .Z(n575) );
  AND U805 ( .A(n574), .B(n575), .Z(n1956) );
  NAND U806 ( .A(n1974), .B(sreg[376]), .Z(n576) );
  XOR U807 ( .A(sreg[376]), .B(n1974), .Z(n577) );
  NANDN U808 ( .A(n1975), .B(n577), .Z(n578) );
  NAND U809 ( .A(n576), .B(n578), .Z(n1983) );
  XOR U810 ( .A(n1999), .B(sreg[379]), .Z(n579) );
  NANDN U811 ( .A(n2000), .B(n579), .Z(n580) );
  NAND U812 ( .A(n1999), .B(sreg[379]), .Z(n581) );
  AND U813 ( .A(n580), .B(n581), .Z(n2006) );
  NAND U814 ( .A(n2023), .B(sreg[382]), .Z(n582) );
  XOR U815 ( .A(sreg[382]), .B(n2023), .Z(n583) );
  NANDN U816 ( .A(n2022), .B(n583), .Z(n584) );
  NAND U817 ( .A(n582), .B(n584), .Z(n2031) );
  XOR U818 ( .A(n2049), .B(sreg[385]), .Z(n585) );
  NANDN U819 ( .A(n2050), .B(n585), .Z(n586) );
  NAND U820 ( .A(n2049), .B(sreg[385]), .Z(n587) );
  AND U821 ( .A(n586), .B(n587), .Z(n2056) );
  NAND U822 ( .A(n2074), .B(sreg[388]), .Z(n588) );
  XOR U823 ( .A(sreg[388]), .B(n2074), .Z(n589) );
  NANDN U824 ( .A(n2075), .B(n589), .Z(n590) );
  NAND U825 ( .A(n588), .B(n590), .Z(n2083) );
  NAND U826 ( .A(n2101), .B(sreg[391]), .Z(n591) );
  XOR U827 ( .A(sreg[391]), .B(n2101), .Z(n592) );
  NAND U828 ( .A(n592), .B(n2100), .Z(n593) );
  NAND U829 ( .A(n591), .B(n593), .Z(n2107) );
  NAND U830 ( .A(n2124), .B(sreg[394]), .Z(n594) );
  XOR U831 ( .A(sreg[394]), .B(n2124), .Z(n595) );
  NANDN U832 ( .A(n2123), .B(n595), .Z(n596) );
  NAND U833 ( .A(n594), .B(n596), .Z(n2132) );
  XOR U834 ( .A(n2148), .B(sreg[397]), .Z(n597) );
  NANDN U835 ( .A(n2149), .B(n597), .Z(n598) );
  NAND U836 ( .A(n2148), .B(sreg[397]), .Z(n599) );
  AND U837 ( .A(n598), .B(n599), .Z(n2155) );
  NAND U838 ( .A(n2173), .B(sreg[400]), .Z(n600) );
  XOR U839 ( .A(sreg[400]), .B(n2173), .Z(n601) );
  NANDN U840 ( .A(n2174), .B(n601), .Z(n602) );
  NAND U841 ( .A(n600), .B(n602), .Z(n2182) );
  XOR U842 ( .A(n2200), .B(sreg[403]), .Z(n603) );
  NANDN U843 ( .A(n2201), .B(n603), .Z(n604) );
  NAND U844 ( .A(n2200), .B(sreg[403]), .Z(n605) );
  AND U845 ( .A(n604), .B(n605), .Z(n2207) );
  NAND U846 ( .A(n2224), .B(sreg[406]), .Z(n606) );
  XOR U847 ( .A(sreg[406]), .B(n2224), .Z(n607) );
  NANDN U848 ( .A(n2223), .B(n607), .Z(n608) );
  NAND U849 ( .A(n606), .B(n608), .Z(n2232) );
  XOR U850 ( .A(n2248), .B(sreg[409]), .Z(n609) );
  NANDN U851 ( .A(n2249), .B(n609), .Z(n610) );
  NAND U852 ( .A(n2248), .B(sreg[409]), .Z(n611) );
  AND U853 ( .A(n610), .B(n611), .Z(n2255) );
  NAND U854 ( .A(n2273), .B(sreg[412]), .Z(n612) );
  XOR U855 ( .A(sreg[412]), .B(n2273), .Z(n613) );
  NANDN U856 ( .A(n2274), .B(n613), .Z(n614) );
  NAND U857 ( .A(n612), .B(n614), .Z(n2282) );
  XOR U858 ( .A(n2298), .B(sreg[415]), .Z(n615) );
  NANDN U859 ( .A(n2299), .B(n615), .Z(n616) );
  NAND U860 ( .A(n2298), .B(sreg[415]), .Z(n617) );
  AND U861 ( .A(n616), .B(n617), .Z(n2308) );
  NAND U862 ( .A(n2323), .B(sreg[418]), .Z(n618) );
  XOR U863 ( .A(sreg[418]), .B(n2323), .Z(n619) );
  NAND U864 ( .A(n619), .B(n2322), .Z(n620) );
  NAND U865 ( .A(n618), .B(n620), .Z(n2331) );
  XOR U866 ( .A(n2347), .B(sreg[421]), .Z(n621) );
  NANDN U867 ( .A(n2348), .B(n621), .Z(n622) );
  NAND U868 ( .A(n2347), .B(sreg[421]), .Z(n623) );
  AND U869 ( .A(n622), .B(n623), .Z(n2354) );
  NAND U870 ( .A(n2371), .B(sreg[424]), .Z(n624) );
  XOR U871 ( .A(sreg[424]), .B(n2371), .Z(n625) );
  NANDN U872 ( .A(n2370), .B(n625), .Z(n626) );
  NAND U873 ( .A(n624), .B(n626), .Z(n2379) );
  XOR U874 ( .A(n2395), .B(sreg[427]), .Z(n627) );
  NANDN U875 ( .A(n2396), .B(n627), .Z(n628) );
  NAND U876 ( .A(n2395), .B(sreg[427]), .Z(n629) );
  AND U877 ( .A(n628), .B(n629), .Z(n2402) );
  NAND U878 ( .A(n2419), .B(sreg[430]), .Z(n630) );
  XOR U879 ( .A(sreg[430]), .B(n2419), .Z(n631) );
  NANDN U880 ( .A(n2418), .B(n631), .Z(n632) );
  NAND U881 ( .A(n630), .B(n632), .Z(n2427) );
  XOR U882 ( .A(n2445), .B(sreg[433]), .Z(n633) );
  NANDN U883 ( .A(n2446), .B(n633), .Z(n634) );
  NAND U884 ( .A(n2445), .B(sreg[433]), .Z(n635) );
  AND U885 ( .A(n634), .B(n635), .Z(n2452) );
  NAND U886 ( .A(n2469), .B(sreg[436]), .Z(n636) );
  XOR U887 ( .A(sreg[436]), .B(n2469), .Z(n637) );
  NANDN U888 ( .A(n2468), .B(n637), .Z(n638) );
  NAND U889 ( .A(n636), .B(n638), .Z(n2477) );
  XOR U890 ( .A(n2493), .B(sreg[439]), .Z(n639) );
  NANDN U891 ( .A(n2494), .B(n639), .Z(n640) );
  NAND U892 ( .A(n2493), .B(sreg[439]), .Z(n641) );
  AND U893 ( .A(n640), .B(n641), .Z(n2500) );
  NAND U894 ( .A(n2517), .B(sreg[442]), .Z(n642) );
  XOR U895 ( .A(sreg[442]), .B(n2517), .Z(n643) );
  NANDN U896 ( .A(n2516), .B(n643), .Z(n644) );
  NAND U897 ( .A(n642), .B(n644), .Z(n2525) );
  XOR U898 ( .A(n2541), .B(sreg[445]), .Z(n645) );
  NANDN U899 ( .A(n2542), .B(n645), .Z(n646) );
  NAND U900 ( .A(n2541), .B(sreg[445]), .Z(n647) );
  AND U901 ( .A(n646), .B(n647), .Z(n2548) );
  NAND U902 ( .A(n2565), .B(sreg[448]), .Z(n648) );
  XOR U903 ( .A(sreg[448]), .B(n2565), .Z(n649) );
  NANDN U904 ( .A(n2564), .B(n649), .Z(n650) );
  NAND U905 ( .A(n648), .B(n650), .Z(n2573) );
  XOR U906 ( .A(n2589), .B(sreg[451]), .Z(n651) );
  NANDN U907 ( .A(n2590), .B(n651), .Z(n652) );
  NAND U908 ( .A(n2589), .B(sreg[451]), .Z(n653) );
  AND U909 ( .A(n652), .B(n653), .Z(n2596) );
  NAND U910 ( .A(n2613), .B(sreg[454]), .Z(n654) );
  XOR U911 ( .A(sreg[454]), .B(n2613), .Z(n655) );
  NANDN U912 ( .A(n2612), .B(n655), .Z(n656) );
  NAND U913 ( .A(n654), .B(n656), .Z(n2621) );
  XOR U914 ( .A(n2637), .B(sreg[457]), .Z(n657) );
  NANDN U915 ( .A(n2638), .B(n657), .Z(n658) );
  NAND U916 ( .A(n2637), .B(sreg[457]), .Z(n659) );
  AND U917 ( .A(n658), .B(n659), .Z(n2644) );
  NAND U918 ( .A(n2661), .B(sreg[460]), .Z(n660) );
  XOR U919 ( .A(sreg[460]), .B(n2661), .Z(n661) );
  NANDN U920 ( .A(n2660), .B(n661), .Z(n662) );
  NAND U921 ( .A(n660), .B(n662), .Z(n2669) );
  XOR U922 ( .A(n2687), .B(sreg[463]), .Z(n663) );
  NANDN U923 ( .A(n2688), .B(n663), .Z(n664) );
  NAND U924 ( .A(n2687), .B(sreg[463]), .Z(n665) );
  AND U925 ( .A(n664), .B(n665), .Z(n2694) );
  NAND U926 ( .A(n2711), .B(sreg[466]), .Z(n666) );
  XOR U927 ( .A(sreg[466]), .B(n2711), .Z(n667) );
  NANDN U928 ( .A(n2710), .B(n667), .Z(n668) );
  NAND U929 ( .A(n666), .B(n668), .Z(n2719) );
  XOR U930 ( .A(n2735), .B(sreg[469]), .Z(n669) );
  NANDN U931 ( .A(n2736), .B(n669), .Z(n670) );
  NAND U932 ( .A(n2735), .B(sreg[469]), .Z(n671) );
  AND U933 ( .A(n670), .B(n671), .Z(n2742) );
  NAND U934 ( .A(n2759), .B(sreg[472]), .Z(n672) );
  XOR U935 ( .A(sreg[472]), .B(n2759), .Z(n673) );
  NANDN U936 ( .A(n2758), .B(n673), .Z(n674) );
  NAND U937 ( .A(n672), .B(n674), .Z(n2765) );
  XOR U938 ( .A(n2783), .B(sreg[475]), .Z(n675) );
  NANDN U939 ( .A(n2784), .B(n675), .Z(n676) );
  NAND U940 ( .A(n2783), .B(sreg[475]), .Z(n677) );
  AND U941 ( .A(n676), .B(n677), .Z(n2790) );
  NAND U942 ( .A(n2807), .B(sreg[478]), .Z(n678) );
  XOR U943 ( .A(sreg[478]), .B(n2807), .Z(n679) );
  NANDN U944 ( .A(n2806), .B(n679), .Z(n680) );
  NAND U945 ( .A(n678), .B(n680), .Z(n2815) );
  XOR U946 ( .A(n2831), .B(sreg[481]), .Z(n681) );
  NANDN U947 ( .A(n2832), .B(n681), .Z(n682) );
  NAND U948 ( .A(n2831), .B(sreg[481]), .Z(n683) );
  AND U949 ( .A(n682), .B(n683), .Z(n2838) );
  NAND U950 ( .A(n2855), .B(sreg[484]), .Z(n684) );
  XOR U951 ( .A(sreg[484]), .B(n2855), .Z(n685) );
  NANDN U952 ( .A(n2854), .B(n685), .Z(n686) );
  NAND U953 ( .A(n684), .B(n686), .Z(n2863) );
  XOR U954 ( .A(n2879), .B(sreg[487]), .Z(n687) );
  NANDN U955 ( .A(n2880), .B(n687), .Z(n688) );
  NAND U956 ( .A(n2879), .B(sreg[487]), .Z(n689) );
  AND U957 ( .A(n688), .B(n689), .Z(n2886) );
  NAND U958 ( .A(n2903), .B(sreg[490]), .Z(n690) );
  XOR U959 ( .A(sreg[490]), .B(n2903), .Z(n691) );
  NANDN U960 ( .A(n2902), .B(n691), .Z(n692) );
  NAND U961 ( .A(n690), .B(n692), .Z(n2911) );
  NAND U962 ( .A(n2929), .B(sreg[493]), .Z(n693) );
  XOR U963 ( .A(sreg[493]), .B(n2929), .Z(n694) );
  NAND U964 ( .A(n694), .B(n2928), .Z(n695) );
  NAND U965 ( .A(n693), .B(n695), .Z(n2935) );
  NAND U966 ( .A(n2953), .B(sreg[496]), .Z(n696) );
  XOR U967 ( .A(sreg[496]), .B(n2953), .Z(n697) );
  NANDN U968 ( .A(n2954), .B(n697), .Z(n698) );
  NAND U969 ( .A(n696), .B(n698), .Z(n2962) );
  XOR U970 ( .A(n2978), .B(sreg[499]), .Z(n699) );
  NANDN U971 ( .A(n2979), .B(n699), .Z(n700) );
  NAND U972 ( .A(n2978), .B(sreg[499]), .Z(n701) );
  AND U973 ( .A(n700), .B(n701), .Z(n2985) );
  NAND U974 ( .A(n3002), .B(sreg[502]), .Z(n702) );
  XOR U975 ( .A(sreg[502]), .B(n3002), .Z(n703) );
  NANDN U976 ( .A(n3001), .B(n703), .Z(n704) );
  NAND U977 ( .A(n702), .B(n704), .Z(n3010) );
  NAND U978 ( .A(n3028), .B(sreg[505]), .Z(n705) );
  XOR U979 ( .A(sreg[505]), .B(n3028), .Z(n706) );
  NAND U980 ( .A(n706), .B(n3027), .Z(n707) );
  NAND U981 ( .A(n705), .B(n707), .Z(n3034) );
  XOR U982 ( .A(n3055), .B(n3054), .Z(n708) );
  NANDN U983 ( .A(sreg[508]), .B(n708), .Z(n709) );
  NAND U984 ( .A(n3055), .B(n3054), .Z(n710) );
  AND U985 ( .A(n709), .B(n710), .Z(n3062) );
  OR U986 ( .A(n1161), .B(n1160), .Z(n711) );
  NAND U987 ( .A(n1163), .B(n1162), .Z(n712) );
  NAND U988 ( .A(n711), .B(n712), .Z(n1170) );
  XOR U989 ( .A(n1011), .B(n1010), .Z(n713) );
  NAND U990 ( .A(n713), .B(sreg[259]), .Z(n714) );
  NAND U991 ( .A(n1011), .B(n1010), .Z(n715) );
  AND U992 ( .A(n714), .B(n715), .Z(n1021) );
  XOR U993 ( .A(n1038), .B(sreg[262]), .Z(n716) );
  NANDN U994 ( .A(n1039), .B(n716), .Z(n717) );
  NAND U995 ( .A(n1038), .B(sreg[262]), .Z(n718) );
  AND U996 ( .A(n717), .B(n718), .Z(n1045) );
  XOR U997 ( .A(n1061), .B(sreg[265]), .Z(n719) );
  NANDN U998 ( .A(n1062), .B(n719), .Z(n720) );
  NAND U999 ( .A(n1061), .B(sreg[265]), .Z(n721) );
  AND U1000 ( .A(n720), .B(n721), .Z(n1068) );
  NAND U1001 ( .A(n1085), .B(sreg[268]), .Z(n722) );
  XOR U1002 ( .A(sreg[268]), .B(n1085), .Z(n723) );
  NANDN U1003 ( .A(n1084), .B(n723), .Z(n724) );
  NAND U1004 ( .A(n722), .B(n724), .Z(n1093) );
  XOR U1005 ( .A(n1109), .B(sreg[271]), .Z(n725) );
  NANDN U1006 ( .A(n1110), .B(n725), .Z(n726) );
  NAND U1007 ( .A(n1109), .B(sreg[271]), .Z(n727) );
  AND U1008 ( .A(n726), .B(n727), .Z(n1116) );
  NAND U1009 ( .A(n1133), .B(sreg[274]), .Z(n728) );
  XOR U1010 ( .A(sreg[274]), .B(n1133), .Z(n729) );
  NANDN U1011 ( .A(n1132), .B(n729), .Z(n730) );
  NAND U1012 ( .A(n728), .B(n730), .Z(n1141) );
  XOR U1013 ( .A(n1157), .B(sreg[277]), .Z(n731) );
  NANDN U1014 ( .A(n1158), .B(n731), .Z(n732) );
  NAND U1015 ( .A(n1157), .B(sreg[277]), .Z(n733) );
  AND U1016 ( .A(n732), .B(n733), .Z(n1164) );
  XOR U1017 ( .A(n1193), .B(sreg[281]), .Z(n734) );
  NANDN U1018 ( .A(n1194), .B(n734), .Z(n735) );
  NAND U1019 ( .A(n1193), .B(sreg[281]), .Z(n736) );
  AND U1020 ( .A(n735), .B(n736), .Z(n1202) );
  NAND U1021 ( .A(n1219), .B(sreg[284]), .Z(n737) );
  XOR U1022 ( .A(sreg[284]), .B(n1219), .Z(n738) );
  NANDN U1023 ( .A(n1218), .B(n738), .Z(n739) );
  NAND U1024 ( .A(n737), .B(n739), .Z(n1227) );
  XOR U1025 ( .A(n1243), .B(sreg[287]), .Z(n740) );
  NANDN U1026 ( .A(n1244), .B(n740), .Z(n741) );
  NAND U1027 ( .A(n1243), .B(sreg[287]), .Z(n742) );
  AND U1028 ( .A(n741), .B(n742), .Z(n1250) );
  NAND U1029 ( .A(n1267), .B(sreg[290]), .Z(n743) );
  XOR U1030 ( .A(sreg[290]), .B(n1267), .Z(n744) );
  NANDN U1031 ( .A(n1266), .B(n744), .Z(n745) );
  NAND U1032 ( .A(n743), .B(n745), .Z(n1275) );
  XOR U1033 ( .A(n1291), .B(sreg[293]), .Z(n746) );
  NANDN U1034 ( .A(n1292), .B(n746), .Z(n747) );
  NAND U1035 ( .A(n1291), .B(sreg[293]), .Z(n748) );
  AND U1036 ( .A(n747), .B(n748), .Z(n1298) );
  NAND U1037 ( .A(n1315), .B(sreg[296]), .Z(n749) );
  XOR U1038 ( .A(sreg[296]), .B(n1315), .Z(n750) );
  NANDN U1039 ( .A(n1314), .B(n750), .Z(n751) );
  NAND U1040 ( .A(n749), .B(n751), .Z(n1323) );
  XOR U1041 ( .A(n1339), .B(sreg[299]), .Z(n752) );
  NANDN U1042 ( .A(n1340), .B(n752), .Z(n753) );
  NAND U1043 ( .A(n1339), .B(sreg[299]), .Z(n754) );
  AND U1044 ( .A(n753), .B(n754), .Z(n1346) );
  NAND U1045 ( .A(n1362), .B(sreg[302]), .Z(n755) );
  XOR U1046 ( .A(sreg[302]), .B(n1362), .Z(n756) );
  NANDN U1047 ( .A(n1363), .B(n756), .Z(n757) );
  NAND U1048 ( .A(n755), .B(n757), .Z(n1371) );
  XOR U1049 ( .A(n1387), .B(sreg[305]), .Z(n758) );
  NANDN U1050 ( .A(n1388), .B(n758), .Z(n759) );
  NAND U1051 ( .A(n1387), .B(sreg[305]), .Z(n760) );
  AND U1052 ( .A(n759), .B(n760), .Z(n1394) );
  NAND U1053 ( .A(n1410), .B(sreg[308]), .Z(n761) );
  XOR U1054 ( .A(sreg[308]), .B(n1410), .Z(n762) );
  NANDN U1055 ( .A(n1411), .B(n762), .Z(n763) );
  NAND U1056 ( .A(n761), .B(n763), .Z(n1419) );
  XOR U1057 ( .A(n1435), .B(sreg[311]), .Z(n764) );
  NANDN U1058 ( .A(n1436), .B(n764), .Z(n765) );
  NAND U1059 ( .A(n1435), .B(sreg[311]), .Z(n766) );
  AND U1060 ( .A(n765), .B(n766), .Z(n1442) );
  NAND U1061 ( .A(n1459), .B(sreg[314]), .Z(n767) );
  XOR U1062 ( .A(sreg[314]), .B(n1459), .Z(n768) );
  NANDN U1063 ( .A(n1458), .B(n768), .Z(n769) );
  NAND U1064 ( .A(n767), .B(n769), .Z(n1467) );
  XOR U1065 ( .A(n1483), .B(sreg[317]), .Z(n770) );
  NANDN U1066 ( .A(n1484), .B(n770), .Z(n771) );
  NAND U1067 ( .A(n1483), .B(sreg[317]), .Z(n772) );
  AND U1068 ( .A(n771), .B(n772), .Z(n1490) );
  NAND U1069 ( .A(n1508), .B(sreg[320]), .Z(n773) );
  XOR U1070 ( .A(sreg[320]), .B(n1508), .Z(n774) );
  NANDN U1071 ( .A(n1509), .B(n774), .Z(n775) );
  NAND U1072 ( .A(n773), .B(n775), .Z(n1517) );
  XOR U1073 ( .A(n1533), .B(sreg[323]), .Z(n776) );
  NANDN U1074 ( .A(n1534), .B(n776), .Z(n777) );
  NAND U1075 ( .A(n1533), .B(sreg[323]), .Z(n778) );
  AND U1076 ( .A(n777), .B(n778), .Z(n1540) );
  NAND U1077 ( .A(n1558), .B(sreg[326]), .Z(n779) );
  XOR U1078 ( .A(sreg[326]), .B(n1558), .Z(n780) );
  NANDN U1079 ( .A(n1559), .B(n780), .Z(n781) );
  NAND U1080 ( .A(n779), .B(n781), .Z(n1567) );
  XOR U1081 ( .A(n1585), .B(sreg[329]), .Z(n782) );
  NANDN U1082 ( .A(n1586), .B(n782), .Z(n783) );
  NAND U1083 ( .A(n1585), .B(sreg[329]), .Z(n784) );
  AND U1084 ( .A(n783), .B(n784), .Z(n1592) );
  NAND U1085 ( .A(n1609), .B(sreg[332]), .Z(n785) );
  XOR U1086 ( .A(sreg[332]), .B(n1609), .Z(n786) );
  NANDN U1087 ( .A(n1608), .B(n786), .Z(n787) );
  NAND U1088 ( .A(n785), .B(n787), .Z(n1617) );
  XOR U1089 ( .A(n1633), .B(sreg[335]), .Z(n788) );
  NANDN U1090 ( .A(n1634), .B(n788), .Z(n789) );
  NAND U1091 ( .A(n1633), .B(sreg[335]), .Z(n790) );
  AND U1092 ( .A(n789), .B(n790), .Z(n1640) );
  NAND U1093 ( .A(n1657), .B(sreg[338]), .Z(n791) );
  XOR U1094 ( .A(sreg[338]), .B(n1657), .Z(n792) );
  NANDN U1095 ( .A(n1656), .B(n792), .Z(n793) );
  NAND U1096 ( .A(n791), .B(n793), .Z(n1665) );
  NAND U1097 ( .A(n1681), .B(sreg[341]), .Z(n794) );
  XOR U1098 ( .A(sreg[341]), .B(n1681), .Z(n795) );
  NANDN U1099 ( .A(n1682), .B(n795), .Z(n796) );
  NAND U1100 ( .A(n794), .B(n796), .Z(n1690) );
  NAND U1101 ( .A(n1707), .B(sreg[344]), .Z(n797) );
  XOR U1102 ( .A(sreg[344]), .B(n1707), .Z(n798) );
  NANDN U1103 ( .A(n1706), .B(n798), .Z(n799) );
  NAND U1104 ( .A(n797), .B(n799), .Z(n1715) );
  XOR U1105 ( .A(n1733), .B(sreg[347]), .Z(n800) );
  NANDN U1106 ( .A(n1734), .B(n800), .Z(n801) );
  NAND U1107 ( .A(n1733), .B(sreg[347]), .Z(n802) );
  AND U1108 ( .A(n801), .B(n802), .Z(n1740) );
  NAND U1109 ( .A(n1758), .B(sreg[350]), .Z(n803) );
  XOR U1110 ( .A(sreg[350]), .B(n1758), .Z(n804) );
  NANDN U1111 ( .A(n1759), .B(n804), .Z(n805) );
  NAND U1112 ( .A(n803), .B(n805), .Z(n1767) );
  NAND U1113 ( .A(n1785), .B(sreg[353]), .Z(n806) );
  XOR U1114 ( .A(sreg[353]), .B(n1785), .Z(n807) );
  NANDN U1115 ( .A(n1786), .B(n807), .Z(n808) );
  NAND U1116 ( .A(n806), .B(n808), .Z(n1794) );
  NAND U1117 ( .A(n1811), .B(sreg[356]), .Z(n809) );
  XOR U1118 ( .A(sreg[356]), .B(n1811), .Z(n810) );
  NANDN U1119 ( .A(n1810), .B(n810), .Z(n811) );
  NAND U1120 ( .A(n809), .B(n811), .Z(n1819) );
  XOR U1121 ( .A(n1835), .B(sreg[359]), .Z(n812) );
  NANDN U1122 ( .A(n1836), .B(n812), .Z(n813) );
  NAND U1123 ( .A(n1835), .B(sreg[359]), .Z(n814) );
  AND U1124 ( .A(n813), .B(n814), .Z(n1842) );
  NAND U1125 ( .A(n1859), .B(sreg[362]), .Z(n815) );
  XOR U1126 ( .A(sreg[362]), .B(n1859), .Z(n816) );
  NANDN U1127 ( .A(n1858), .B(n816), .Z(n817) );
  NAND U1128 ( .A(n815), .B(n817), .Z(n1867) );
  NAND U1129 ( .A(n1883), .B(sreg[365]), .Z(n818) );
  XOR U1130 ( .A(sreg[365]), .B(n1883), .Z(n819) );
  NANDN U1131 ( .A(n1884), .B(n819), .Z(n820) );
  NAND U1132 ( .A(n818), .B(n820), .Z(n1892) );
  NAND U1133 ( .A(n1909), .B(sreg[368]), .Z(n821) );
  XOR U1134 ( .A(sreg[368]), .B(n1909), .Z(n822) );
  NANDN U1135 ( .A(n1908), .B(n822), .Z(n823) );
  NAND U1136 ( .A(n821), .B(n823), .Z(n1917) );
  XOR U1137 ( .A(n1933), .B(sreg[371]), .Z(n824) );
  NANDN U1138 ( .A(n1934), .B(n824), .Z(n825) );
  NAND U1139 ( .A(n1933), .B(sreg[371]), .Z(n826) );
  AND U1140 ( .A(n825), .B(n826), .Z(n1940) );
  NAND U1141 ( .A(n1957), .B(sreg[374]), .Z(n827) );
  XOR U1142 ( .A(sreg[374]), .B(n1957), .Z(n828) );
  NANDN U1143 ( .A(n1956), .B(n828), .Z(n829) );
  NAND U1144 ( .A(n827), .B(n829), .Z(n1965) );
  XOR U1145 ( .A(n1983), .B(sreg[377]), .Z(n830) );
  NANDN U1146 ( .A(n1984), .B(n830), .Z(n831) );
  NAND U1147 ( .A(n1983), .B(sreg[377]), .Z(n832) );
  AND U1148 ( .A(n831), .B(n832), .Z(n1990) );
  NAND U1149 ( .A(n2007), .B(sreg[380]), .Z(n833) );
  XOR U1150 ( .A(sreg[380]), .B(n2007), .Z(n834) );
  NANDN U1151 ( .A(n2006), .B(n834), .Z(n835) );
  NAND U1152 ( .A(n833), .B(n835), .Z(n2015) );
  NAND U1153 ( .A(n2031), .B(sreg[383]), .Z(n836) );
  XOR U1154 ( .A(sreg[383]), .B(n2031), .Z(n837) );
  NANDN U1155 ( .A(n2032), .B(n837), .Z(n838) );
  NAND U1156 ( .A(n836), .B(n838), .Z(n2040) );
  NAND U1157 ( .A(n2057), .B(sreg[386]), .Z(n839) );
  XOR U1158 ( .A(sreg[386]), .B(n2057), .Z(n840) );
  NANDN U1159 ( .A(n2056), .B(n840), .Z(n841) );
  NAND U1160 ( .A(n839), .B(n841), .Z(n2065) );
  XOR U1161 ( .A(n2083), .B(sreg[389]), .Z(n842) );
  NANDN U1162 ( .A(n2084), .B(n842), .Z(n843) );
  NAND U1163 ( .A(n2083), .B(sreg[389]), .Z(n844) );
  AND U1164 ( .A(n843), .B(n844), .Z(n2093) );
  NAND U1165 ( .A(n2108), .B(sreg[392]), .Z(n845) );
  XOR U1166 ( .A(sreg[392]), .B(n2108), .Z(n846) );
  NAND U1167 ( .A(n846), .B(n2107), .Z(n847) );
  NAND U1168 ( .A(n845), .B(n847), .Z(n2116) );
  XOR U1169 ( .A(n2132), .B(sreg[395]), .Z(n848) );
  NANDN U1170 ( .A(n2133), .B(n848), .Z(n849) );
  NAND U1171 ( .A(n2132), .B(sreg[395]), .Z(n850) );
  AND U1172 ( .A(n849), .B(n850), .Z(n2139) );
  NAND U1173 ( .A(n2156), .B(sreg[398]), .Z(n851) );
  XOR U1174 ( .A(sreg[398]), .B(n2156), .Z(n852) );
  NANDN U1175 ( .A(n2155), .B(n852), .Z(n853) );
  NAND U1176 ( .A(n851), .B(n853), .Z(n2164) );
  NAND U1177 ( .A(n2182), .B(sreg[401]), .Z(n854) );
  XOR U1178 ( .A(sreg[401]), .B(n2182), .Z(n855) );
  NANDN U1179 ( .A(n2183), .B(n855), .Z(n856) );
  NAND U1180 ( .A(n854), .B(n856), .Z(n2191) );
  NAND U1181 ( .A(n2208), .B(sreg[404]), .Z(n857) );
  XOR U1182 ( .A(sreg[404]), .B(n2208), .Z(n858) );
  NANDN U1183 ( .A(n2207), .B(n858), .Z(n859) );
  NAND U1184 ( .A(n857), .B(n859), .Z(n2216) );
  XOR U1185 ( .A(n2232), .B(sreg[407]), .Z(n860) );
  NANDN U1186 ( .A(n2233), .B(n860), .Z(n861) );
  NAND U1187 ( .A(n2232), .B(sreg[407]), .Z(n862) );
  AND U1188 ( .A(n861), .B(n862), .Z(n2239) );
  NAND U1189 ( .A(n2256), .B(sreg[410]), .Z(n863) );
  XOR U1190 ( .A(sreg[410]), .B(n2256), .Z(n864) );
  NANDN U1191 ( .A(n2255), .B(n864), .Z(n865) );
  NAND U1192 ( .A(n863), .B(n865), .Z(n2264) );
  XOR U1193 ( .A(n2282), .B(sreg[413]), .Z(n866) );
  NANDN U1194 ( .A(n2283), .B(n866), .Z(n867) );
  NAND U1195 ( .A(n2282), .B(sreg[413]), .Z(n868) );
  AND U1196 ( .A(n867), .B(n868), .Z(n2289) );
  NAND U1197 ( .A(n2309), .B(sreg[416]), .Z(n869) );
  XOR U1198 ( .A(sreg[416]), .B(n2309), .Z(n870) );
  NANDN U1199 ( .A(n2308), .B(n870), .Z(n871) );
  NAND U1200 ( .A(n869), .B(n871), .Z(n2315) );
  XOR U1201 ( .A(n2331), .B(sreg[419]), .Z(n872) );
  NANDN U1202 ( .A(n2332), .B(n872), .Z(n873) );
  NAND U1203 ( .A(n2331), .B(sreg[419]), .Z(n874) );
  AND U1204 ( .A(n873), .B(n874), .Z(n2338) );
  NAND U1205 ( .A(n2355), .B(sreg[422]), .Z(n875) );
  XOR U1206 ( .A(sreg[422]), .B(n2355), .Z(n876) );
  NANDN U1207 ( .A(n2354), .B(n876), .Z(n877) );
  NAND U1208 ( .A(n875), .B(n877), .Z(n2363) );
  XOR U1209 ( .A(n2379), .B(sreg[425]), .Z(n878) );
  NANDN U1210 ( .A(n2380), .B(n878), .Z(n879) );
  NAND U1211 ( .A(n2379), .B(sreg[425]), .Z(n880) );
  AND U1212 ( .A(n879), .B(n880), .Z(n2386) );
  NAND U1213 ( .A(n2403), .B(sreg[428]), .Z(n881) );
  XOR U1214 ( .A(sreg[428]), .B(n2403), .Z(n882) );
  NANDN U1215 ( .A(n2402), .B(n882), .Z(n883) );
  NAND U1216 ( .A(n881), .B(n883), .Z(n2411) );
  NAND U1217 ( .A(n2427), .B(sreg[431]), .Z(n884) );
  XOR U1218 ( .A(sreg[431]), .B(n2427), .Z(n885) );
  NANDN U1219 ( .A(n2428), .B(n885), .Z(n886) );
  NAND U1220 ( .A(n884), .B(n886), .Z(n2436) );
  NAND U1221 ( .A(n2453), .B(sreg[434]), .Z(n887) );
  XOR U1222 ( .A(sreg[434]), .B(n2453), .Z(n888) );
  NANDN U1223 ( .A(n2452), .B(n888), .Z(n889) );
  NAND U1224 ( .A(n887), .B(n889), .Z(n2461) );
  XOR U1225 ( .A(n2477), .B(sreg[437]), .Z(n890) );
  NANDN U1226 ( .A(n2478), .B(n890), .Z(n891) );
  NAND U1227 ( .A(n2477), .B(sreg[437]), .Z(n892) );
  AND U1228 ( .A(n891), .B(n892), .Z(n2484) );
  NAND U1229 ( .A(n2501), .B(sreg[440]), .Z(n893) );
  XOR U1230 ( .A(sreg[440]), .B(n2501), .Z(n894) );
  NANDN U1231 ( .A(n2500), .B(n894), .Z(n895) );
  NAND U1232 ( .A(n893), .B(n895), .Z(n2509) );
  XOR U1233 ( .A(n2525), .B(sreg[443]), .Z(n896) );
  NANDN U1234 ( .A(n2526), .B(n896), .Z(n897) );
  NAND U1235 ( .A(n2525), .B(sreg[443]), .Z(n898) );
  AND U1236 ( .A(n897), .B(n898), .Z(n2532) );
  NAND U1237 ( .A(n2549), .B(sreg[446]), .Z(n899) );
  XOR U1238 ( .A(sreg[446]), .B(n2549), .Z(n900) );
  NANDN U1239 ( .A(n2548), .B(n900), .Z(n901) );
  NAND U1240 ( .A(n899), .B(n901), .Z(n2557) );
  XOR U1241 ( .A(n2573), .B(sreg[449]), .Z(n902) );
  NANDN U1242 ( .A(n2574), .B(n902), .Z(n903) );
  NAND U1243 ( .A(n2573), .B(sreg[449]), .Z(n904) );
  AND U1244 ( .A(n903), .B(n904), .Z(n2580) );
  NAND U1245 ( .A(n2597), .B(sreg[452]), .Z(n905) );
  XOR U1246 ( .A(sreg[452]), .B(n2597), .Z(n906) );
  NANDN U1247 ( .A(n2596), .B(n906), .Z(n907) );
  NAND U1248 ( .A(n905), .B(n907), .Z(n2605) );
  XOR U1249 ( .A(n2621), .B(sreg[455]), .Z(n908) );
  NANDN U1250 ( .A(n2622), .B(n908), .Z(n909) );
  NAND U1251 ( .A(n2621), .B(sreg[455]), .Z(n910) );
  AND U1252 ( .A(n909), .B(n910), .Z(n2628) );
  NAND U1253 ( .A(n2645), .B(sreg[458]), .Z(n911) );
  XOR U1254 ( .A(sreg[458]), .B(n2645), .Z(n912) );
  NANDN U1255 ( .A(n2644), .B(n912), .Z(n913) );
  NAND U1256 ( .A(n911), .B(n913), .Z(n2653) );
  NAND U1257 ( .A(n2669), .B(sreg[461]), .Z(n914) );
  XOR U1258 ( .A(sreg[461]), .B(n2669), .Z(n915) );
  NANDN U1259 ( .A(n2670), .B(n915), .Z(n916) );
  NAND U1260 ( .A(n914), .B(n916), .Z(n2678) );
  NAND U1261 ( .A(n2695), .B(sreg[464]), .Z(n917) );
  XOR U1262 ( .A(sreg[464]), .B(n2695), .Z(n918) );
  NANDN U1263 ( .A(n2694), .B(n918), .Z(n919) );
  NAND U1264 ( .A(n917), .B(n919), .Z(n2703) );
  XOR U1265 ( .A(n2719), .B(sreg[467]), .Z(n920) );
  NANDN U1266 ( .A(n2720), .B(n920), .Z(n921) );
  NAND U1267 ( .A(n2719), .B(sreg[467]), .Z(n922) );
  AND U1268 ( .A(n921), .B(n922), .Z(n2726) );
  NAND U1269 ( .A(n2743), .B(sreg[470]), .Z(n923) );
  XOR U1270 ( .A(sreg[470]), .B(n2743), .Z(n924) );
  NANDN U1271 ( .A(n2742), .B(n924), .Z(n925) );
  NAND U1272 ( .A(n923), .B(n925), .Z(n2751) );
  NAND U1273 ( .A(n2766), .B(sreg[473]), .Z(n926) );
  XOR U1274 ( .A(sreg[473]), .B(n2766), .Z(n927) );
  NAND U1275 ( .A(n927), .B(n2765), .Z(n928) );
  NAND U1276 ( .A(n926), .B(n928), .Z(n2774) );
  NAND U1277 ( .A(n2791), .B(sreg[476]), .Z(n929) );
  XOR U1278 ( .A(sreg[476]), .B(n2791), .Z(n930) );
  NANDN U1279 ( .A(n2790), .B(n930), .Z(n931) );
  NAND U1280 ( .A(n929), .B(n931), .Z(n2799) );
  XOR U1281 ( .A(n2815), .B(sreg[479]), .Z(n932) );
  NANDN U1282 ( .A(n2816), .B(n932), .Z(n933) );
  NAND U1283 ( .A(n2815), .B(sreg[479]), .Z(n934) );
  AND U1284 ( .A(n933), .B(n934), .Z(n2822) );
  NAND U1285 ( .A(n2839), .B(sreg[482]), .Z(n935) );
  XOR U1286 ( .A(sreg[482]), .B(n2839), .Z(n936) );
  NANDN U1287 ( .A(n2838), .B(n936), .Z(n937) );
  NAND U1288 ( .A(n935), .B(n937), .Z(n2847) );
  XOR U1289 ( .A(n2863), .B(sreg[485]), .Z(n938) );
  NANDN U1290 ( .A(n2864), .B(n938), .Z(n939) );
  NAND U1291 ( .A(n2863), .B(sreg[485]), .Z(n940) );
  AND U1292 ( .A(n939), .B(n940), .Z(n2870) );
  NAND U1293 ( .A(n2887), .B(sreg[488]), .Z(n941) );
  XOR U1294 ( .A(sreg[488]), .B(n2887), .Z(n942) );
  NANDN U1295 ( .A(n2886), .B(n942), .Z(n943) );
  NAND U1296 ( .A(n941), .B(n943), .Z(n2895) );
  XOR U1297 ( .A(n2911), .B(sreg[491]), .Z(n944) );
  NANDN U1298 ( .A(n2912), .B(n944), .Z(n945) );
  NAND U1299 ( .A(n2911), .B(sreg[491]), .Z(n946) );
  AND U1300 ( .A(n945), .B(n946), .Z(n2921) );
  NAND U1301 ( .A(n2936), .B(sreg[494]), .Z(n947) );
  XOR U1302 ( .A(sreg[494]), .B(n2936), .Z(n948) );
  NAND U1303 ( .A(n948), .B(n2935), .Z(n949) );
  NAND U1304 ( .A(n947), .B(n949), .Z(n2944) );
  XOR U1305 ( .A(n2962), .B(sreg[497]), .Z(n950) );
  NANDN U1306 ( .A(n2963), .B(n950), .Z(n951) );
  NAND U1307 ( .A(n2962), .B(sreg[497]), .Z(n952) );
  AND U1308 ( .A(n951), .B(n952), .Z(n2969) );
  NAND U1309 ( .A(n2986), .B(sreg[500]), .Z(n953) );
  XOR U1310 ( .A(sreg[500]), .B(n2986), .Z(n954) );
  NANDN U1311 ( .A(n2985), .B(n954), .Z(n955) );
  NAND U1312 ( .A(n953), .B(n955), .Z(n2994) );
  XOR U1313 ( .A(n3010), .B(sreg[503]), .Z(n956) );
  NANDN U1314 ( .A(n3011), .B(n956), .Z(n957) );
  NAND U1315 ( .A(n3010), .B(sreg[503]), .Z(n958) );
  AND U1316 ( .A(n957), .B(n958), .Z(n3020) );
  NAND U1317 ( .A(n3035), .B(sreg[506]), .Z(n959) );
  XOR U1318 ( .A(sreg[506]), .B(n3035), .Z(n960) );
  NAND U1319 ( .A(n960), .B(n3034), .Z(n961) );
  NAND U1320 ( .A(n959), .B(n961), .Z(n3043) );
  NAND U1321 ( .A(n3063), .B(n3062), .Z(n962) );
  XOR U1322 ( .A(n3062), .B(n3063), .Z(n963) );
  NAND U1323 ( .A(n963), .B(sreg[509]), .Z(n964) );
  NAND U1324 ( .A(n962), .B(n964), .Z(n3067) );
  IV U1325 ( .A(b[0]), .Z(n965) );
  IV U1326 ( .A(b[1]), .Z(n966) );
  ANDN U1327 ( .B(a[0]), .A(n965), .Z(n977) );
  XOR U1328 ( .A(n977), .B(sreg[254]), .Z(c[254]) );
  ANDN U1329 ( .B(a[1]), .A(n965), .Z(n968) );
  NANDN U1330 ( .A(n966), .B(a[0]), .Z(n967) );
  XNOR U1331 ( .A(n968), .B(n967), .Z(n970) );
  XNOR U1332 ( .A(sreg[255]), .B(n970), .Z(n972) );
  NAND U1333 ( .A(n977), .B(sreg[254]), .Z(n971) );
  XOR U1334 ( .A(n972), .B(n971), .Z(c[255]) );
  AND U1335 ( .A(a[2]), .B(b[0]), .Z(n986) );
  NANDN U1336 ( .A(n966), .B(a[1]), .Z(n979) );
  OR U1337 ( .A(n979), .B(n977), .Z(n969) );
  XNOR U1338 ( .A(n986), .B(n969), .Z(n980) );
  XNOR U1339 ( .A(sreg[256]), .B(n980), .Z(n982) );
  NAND U1340 ( .A(n970), .B(sreg[255]), .Z(n974) );
  OR U1341 ( .A(n972), .B(n971), .Z(n973) );
  AND U1342 ( .A(n974), .B(n973), .Z(n981) );
  XOR U1343 ( .A(n982), .B(n981), .Z(c[256]) );
  ANDN U1344 ( .B(a[3]), .A(n965), .Z(n976) );
  NANDN U1345 ( .A(n966), .B(a[2]), .Z(n975) );
  XOR U1346 ( .A(n976), .B(n975), .Z(n988) );
  OR U1347 ( .A(n986), .B(n977), .Z(n978) );
  NANDN U1348 ( .A(n979), .B(n978), .Z(n987) );
  XOR U1349 ( .A(n988), .B(n987), .Z(n992) );
  NAND U1350 ( .A(sreg[256]), .B(n980), .Z(n984) );
  OR U1351 ( .A(n982), .B(n981), .Z(n983) );
  AND U1352 ( .A(n984), .B(n983), .Z(n991) );
  XNOR U1353 ( .A(n991), .B(sreg[257]), .Z(n985) );
  XOR U1354 ( .A(n992), .B(n985), .Z(c[257]) );
  AND U1355 ( .A(a[3]), .B(b[1]), .Z(n995) );
  AND U1356 ( .A(a[4]), .B(b[0]), .Z(n1004) );
  NAND U1357 ( .A(n995), .B(n986), .Z(n990) );
  OR U1358 ( .A(n988), .B(n987), .Z(n989) );
  NAND U1359 ( .A(n990), .B(n989), .Z(n994) );
  XOR U1360 ( .A(n1004), .B(n994), .Z(n996) );
  XNOR U1361 ( .A(n995), .B(n996), .Z(n1001) );
  XOR U1362 ( .A(n1000), .B(sreg[258]), .Z(n993) );
  XNOR U1363 ( .A(n1001), .B(n993), .Z(c[258]) );
  NAND U1364 ( .A(n994), .B(n1004), .Z(n998) );
  NAND U1365 ( .A(n996), .B(n995), .Z(n997) );
  NAND U1366 ( .A(n998), .B(n997), .Z(n1006) );
  ANDN U1367 ( .B(a[5]), .A(n965), .Z(n1015) );
  NANDN U1368 ( .A(n966), .B(a[4]), .Z(n999) );
  XNOR U1369 ( .A(n1015), .B(n999), .Z(n1007) );
  XOR U1370 ( .A(n1006), .B(n1007), .Z(n1011) );
  XOR U1371 ( .A(n1010), .B(sreg[259]), .Z(n1002) );
  XOR U1372 ( .A(n1011), .B(n1002), .Z(c[259]) );
  ANDN U1373 ( .B(a[6]), .A(n965), .Z(n1024) );
  NANDN U1374 ( .A(n966), .B(a[5]), .Z(n1003) );
  XOR U1375 ( .A(n1024), .B(n1003), .Z(n1018) );
  ANDN U1376 ( .B(a[5]), .A(n966), .Z(n1005) );
  NAND U1377 ( .A(n1005), .B(n1004), .Z(n1009) );
  NAND U1378 ( .A(n1007), .B(n1006), .Z(n1008) );
  NAND U1379 ( .A(n1009), .B(n1008), .Z(n1017) );
  XNOR U1380 ( .A(n1018), .B(n1017), .Z(n1022) );
  XOR U1381 ( .A(sreg[260]), .B(n1021), .Z(n1012) );
  XNOR U1382 ( .A(n1022), .B(n1012), .Z(c[260]) );
  ANDN U1383 ( .B(a[7]), .A(n965), .Z(n1014) );
  NANDN U1384 ( .A(n966), .B(a[6]), .Z(n1013) );
  XOR U1385 ( .A(n1014), .B(n1013), .Z(n1026) );
  ANDN U1386 ( .B(a[6]), .A(n966), .Z(n1016) );
  NAND U1387 ( .A(n1016), .B(n1015), .Z(n1020) );
  NANDN U1388 ( .A(n1018), .B(n1017), .Z(n1019) );
  NAND U1389 ( .A(n1020), .B(n1019), .Z(n1025) );
  XNOR U1390 ( .A(n1026), .B(n1025), .Z(n1030) );
  XNOR U1391 ( .A(sreg[261]), .B(n1029), .Z(n1023) );
  XNOR U1392 ( .A(n1030), .B(n1023), .Z(c[261]) );
  ANDN U1393 ( .B(a[7]), .A(n966), .Z(n1033) );
  NAND U1394 ( .A(n1024), .B(n1033), .Z(n1028) );
  NANDN U1395 ( .A(n1026), .B(n1025), .Z(n1027) );
  NAND U1396 ( .A(n1028), .B(n1027), .Z(n1034) );
  ANDN U1397 ( .B(a[8]), .A(n965), .Z(n1032) );
  XNOR U1398 ( .A(n1033), .B(n1032), .Z(n1035) );
  XOR U1399 ( .A(n1034), .B(n1035), .Z(n1039) );
  XOR U1400 ( .A(n1038), .B(sreg[262]), .Z(n1031) );
  XNOR U1401 ( .A(n1039), .B(n1031), .Z(c[262]) );
  OR U1402 ( .A(n1033), .B(n1032), .Z(n1037) );
  OR U1403 ( .A(n1035), .B(n1034), .Z(n1036) );
  NAND U1404 ( .A(n1037), .B(n1036), .Z(n1044) );
  ANDN U1405 ( .B(a[9]), .A(n965), .Z(n1042) );
  ANDN U1406 ( .B(a[8]), .A(n966), .Z(n1041) );
  XOR U1407 ( .A(n1042), .B(n1041), .Z(n1043) );
  XNOR U1408 ( .A(n1044), .B(n1043), .Z(n1046) );
  XOR U1409 ( .A(sreg[263]), .B(n1045), .Z(n1040) );
  XNOR U1410 ( .A(n1046), .B(n1040), .Z(c[263]) );
  ANDN U1411 ( .B(a[10]), .A(n965), .Z(n1049) );
  ANDN U1412 ( .B(a[9]), .A(n966), .Z(n1048) );
  XOR U1413 ( .A(n1049), .B(n1048), .Z(n1050) );
  XNOR U1414 ( .A(n1051), .B(n1050), .Z(n1053) );
  XNOR U1415 ( .A(sreg[264]), .B(n1052), .Z(n1047) );
  XNOR U1416 ( .A(n1053), .B(n1047), .Z(c[264]) );
  NAND U1417 ( .A(b[0]), .B(a[11]), .Z(n1056) );
  NAND U1418 ( .A(b[1]), .B(a[10]), .Z(n1055) );
  XNOR U1419 ( .A(n1056), .B(n1055), .Z(n1058) );
  XNOR U1420 ( .A(n1057), .B(n1058), .Z(n1062) );
  XOR U1421 ( .A(n1061), .B(sreg[265]), .Z(n1054) );
  XNOR U1422 ( .A(n1062), .B(n1054), .Z(c[265]) );
  NAND U1423 ( .A(n1056), .B(n1055), .Z(n1060) );
  NANDN U1424 ( .A(n1058), .B(n1057), .Z(n1059) );
  NAND U1425 ( .A(n1060), .B(n1059), .Z(n1067) );
  ANDN U1426 ( .B(a[12]), .A(n965), .Z(n1065) );
  ANDN U1427 ( .B(a[11]), .A(n966), .Z(n1064) );
  XOR U1428 ( .A(n1065), .B(n1064), .Z(n1066) );
  XNOR U1429 ( .A(n1067), .B(n1066), .Z(n1069) );
  XOR U1430 ( .A(sreg[266]), .B(n1068), .Z(n1063) );
  XNOR U1431 ( .A(n1069), .B(n1063), .Z(c[266]) );
  NAND U1432 ( .A(b[0]), .B(a[13]), .Z(n1072) );
  NAND U1433 ( .A(b[1]), .B(a[12]), .Z(n1071) );
  XNOR U1434 ( .A(n1072), .B(n1071), .Z(n1074) );
  XNOR U1435 ( .A(n1073), .B(n1074), .Z(n1078) );
  XOR U1436 ( .A(n1077), .B(sreg[267]), .Z(n1070) );
  XNOR U1437 ( .A(n1078), .B(n1070), .Z(c[267]) );
  NAND U1438 ( .A(n1072), .B(n1071), .Z(n1076) );
  NANDN U1439 ( .A(n1074), .B(n1073), .Z(n1075) );
  NAND U1440 ( .A(n1076), .B(n1075), .Z(n1083) );
  ANDN U1441 ( .B(a[14]), .A(n965), .Z(n1081) );
  ANDN U1442 ( .B(a[13]), .A(n966), .Z(n1080) );
  XOR U1443 ( .A(n1081), .B(n1080), .Z(n1082) );
  XNOR U1444 ( .A(n1083), .B(n1082), .Z(n1085) );
  XOR U1445 ( .A(sreg[268]), .B(n1084), .Z(n1079) );
  XNOR U1446 ( .A(n1085), .B(n1079), .Z(c[268]) );
  NAND U1447 ( .A(b[0]), .B(a[15]), .Z(n1088) );
  NAND U1448 ( .A(b[1]), .B(a[14]), .Z(n1087) );
  XNOR U1449 ( .A(n1088), .B(n1087), .Z(n1090) );
  XNOR U1450 ( .A(n1089), .B(n1090), .Z(n1094) );
  XOR U1451 ( .A(n1093), .B(sreg[269]), .Z(n1086) );
  XNOR U1452 ( .A(n1094), .B(n1086), .Z(c[269]) );
  NAND U1453 ( .A(n1088), .B(n1087), .Z(n1092) );
  NANDN U1454 ( .A(n1090), .B(n1089), .Z(n1091) );
  NAND U1455 ( .A(n1092), .B(n1091), .Z(n1099) );
  ANDN U1456 ( .B(a[16]), .A(n965), .Z(n1097) );
  ANDN U1457 ( .B(a[15]), .A(n966), .Z(n1096) );
  XOR U1458 ( .A(n1097), .B(n1096), .Z(n1098) );
  XNOR U1459 ( .A(n1099), .B(n1098), .Z(n1101) );
  XOR U1460 ( .A(sreg[270]), .B(n1100), .Z(n1095) );
  XNOR U1461 ( .A(n1101), .B(n1095), .Z(c[270]) );
  NAND U1462 ( .A(b[0]), .B(a[17]), .Z(n1104) );
  NAND U1463 ( .A(b[1]), .B(a[16]), .Z(n1103) );
  XNOR U1464 ( .A(n1104), .B(n1103), .Z(n1106) );
  XNOR U1465 ( .A(n1105), .B(n1106), .Z(n1110) );
  XOR U1466 ( .A(n1109), .B(sreg[271]), .Z(n1102) );
  XNOR U1467 ( .A(n1110), .B(n1102), .Z(c[271]) );
  NAND U1468 ( .A(n1104), .B(n1103), .Z(n1108) );
  NANDN U1469 ( .A(n1106), .B(n1105), .Z(n1107) );
  NAND U1470 ( .A(n1108), .B(n1107), .Z(n1115) );
  ANDN U1471 ( .B(a[18]), .A(n965), .Z(n1113) );
  ANDN U1472 ( .B(a[17]), .A(n966), .Z(n1112) );
  XOR U1473 ( .A(n1113), .B(n1112), .Z(n1114) );
  XNOR U1474 ( .A(n1115), .B(n1114), .Z(n1117) );
  XOR U1475 ( .A(sreg[272]), .B(n1116), .Z(n1111) );
  XNOR U1476 ( .A(n1117), .B(n1111), .Z(c[272]) );
  NAND U1477 ( .A(b[0]), .B(a[19]), .Z(n1120) );
  NAND U1478 ( .A(b[1]), .B(a[18]), .Z(n1119) );
  XNOR U1479 ( .A(n1120), .B(n1119), .Z(n1122) );
  XNOR U1480 ( .A(n1121), .B(n1122), .Z(n1126) );
  XOR U1481 ( .A(n1125), .B(sreg[273]), .Z(n1118) );
  XNOR U1482 ( .A(n1126), .B(n1118), .Z(c[273]) );
  NAND U1483 ( .A(n1120), .B(n1119), .Z(n1124) );
  NANDN U1484 ( .A(n1122), .B(n1121), .Z(n1123) );
  NAND U1485 ( .A(n1124), .B(n1123), .Z(n1131) );
  ANDN U1486 ( .B(a[20]), .A(n965), .Z(n1129) );
  ANDN U1487 ( .B(a[19]), .A(n966), .Z(n1128) );
  XOR U1488 ( .A(n1129), .B(n1128), .Z(n1130) );
  XNOR U1489 ( .A(n1131), .B(n1130), .Z(n1133) );
  XOR U1490 ( .A(sreg[274]), .B(n1132), .Z(n1127) );
  XNOR U1491 ( .A(n1133), .B(n1127), .Z(c[274]) );
  NAND U1492 ( .A(b[0]), .B(a[21]), .Z(n1136) );
  NAND U1493 ( .A(b[1]), .B(a[20]), .Z(n1135) );
  XNOR U1494 ( .A(n1136), .B(n1135), .Z(n1138) );
  XNOR U1495 ( .A(n1137), .B(n1138), .Z(n1142) );
  XOR U1496 ( .A(n1141), .B(sreg[275]), .Z(n1134) );
  XNOR U1497 ( .A(n1142), .B(n1134), .Z(c[275]) );
  NAND U1498 ( .A(n1136), .B(n1135), .Z(n1140) );
  NANDN U1499 ( .A(n1138), .B(n1137), .Z(n1139) );
  NAND U1500 ( .A(n1140), .B(n1139), .Z(n1147) );
  ANDN U1501 ( .B(a[22]), .A(n965), .Z(n1145) );
  ANDN U1502 ( .B(a[21]), .A(n966), .Z(n1144) );
  XOR U1503 ( .A(n1145), .B(n1144), .Z(n1146) );
  XNOR U1504 ( .A(n1147), .B(n1146), .Z(n1149) );
  XOR U1505 ( .A(sreg[276]), .B(n1148), .Z(n1143) );
  XNOR U1506 ( .A(n1149), .B(n1143), .Z(c[276]) );
  NAND U1507 ( .A(b[0]), .B(a[23]), .Z(n1152) );
  NAND U1508 ( .A(b[1]), .B(a[22]), .Z(n1151) );
  XNOR U1509 ( .A(n1152), .B(n1151), .Z(n1154) );
  XNOR U1510 ( .A(n1153), .B(n1154), .Z(n1158) );
  XOR U1511 ( .A(n1157), .B(sreg[277]), .Z(n1150) );
  XNOR U1512 ( .A(n1158), .B(n1150), .Z(c[277]) );
  NAND U1513 ( .A(n1152), .B(n1151), .Z(n1156) );
  NANDN U1514 ( .A(n1154), .B(n1153), .Z(n1155) );
  NAND U1515 ( .A(n1156), .B(n1155), .Z(n1163) );
  ANDN U1516 ( .B(a[24]), .A(n965), .Z(n1161) );
  ANDN U1517 ( .B(a[23]), .A(n966), .Z(n1160) );
  XOR U1518 ( .A(n1161), .B(n1160), .Z(n1162) );
  XNOR U1519 ( .A(n1163), .B(n1162), .Z(n1165) );
  XOR U1520 ( .A(sreg[278]), .B(n1164), .Z(n1159) );
  XNOR U1521 ( .A(n1165), .B(n1159), .Z(c[278]) );
  ANDN U1522 ( .B(a[25]), .A(n965), .Z(n1168) );
  ANDN U1523 ( .B(a[24]), .A(n966), .Z(n1167) );
  XOR U1524 ( .A(n1168), .B(n1167), .Z(n1169) );
  XOR U1525 ( .A(n1170), .B(n1169), .Z(n1176) );
  IV U1526 ( .A(n1174), .Z(n1173) );
  XOR U1527 ( .A(n1173), .B(sreg[279]), .Z(n1166) );
  XOR U1528 ( .A(n1176), .B(n1166), .Z(c[279]) );
  OR U1529 ( .A(n1168), .B(n1167), .Z(n1172) );
  NAND U1530 ( .A(n1170), .B(n1169), .Z(n1171) );
  NAND U1531 ( .A(n1172), .B(n1171), .Z(n1183) );
  ANDN U1532 ( .B(a[26]), .A(n965), .Z(n1181) );
  ANDN U1533 ( .B(a[25]), .A(n966), .Z(n1180) );
  XOR U1534 ( .A(n1181), .B(n1180), .Z(n1182) );
  XNOR U1535 ( .A(n1183), .B(n1182), .Z(n1185) );
  NANDN U1536 ( .A(n1173), .B(sreg[279]), .Z(n1178) );
  OR U1537 ( .A(sreg[279]), .B(n1174), .Z(n1175) );
  NANDN U1538 ( .A(n1176), .B(n1175), .Z(n1177) );
  NAND U1539 ( .A(n1178), .B(n1177), .Z(n1184) );
  XNOR U1540 ( .A(sreg[280]), .B(n1184), .Z(n1179) );
  XNOR U1541 ( .A(n1185), .B(n1179), .Z(c[280]) );
  NAND U1542 ( .A(b[0]), .B(a[27]), .Z(n1188) );
  NAND U1543 ( .A(b[1]), .B(a[26]), .Z(n1187) );
  XNOR U1544 ( .A(n1188), .B(n1187), .Z(n1190) );
  XNOR U1545 ( .A(n1189), .B(n1190), .Z(n1194) );
  XOR U1546 ( .A(n1193), .B(sreg[281]), .Z(n1186) );
  XNOR U1547 ( .A(n1194), .B(n1186), .Z(c[281]) );
  NAND U1548 ( .A(n1188), .B(n1187), .Z(n1192) );
  NANDN U1549 ( .A(n1190), .B(n1189), .Z(n1191) );
  NAND U1550 ( .A(n1192), .B(n1191), .Z(n1198) );
  NAND U1551 ( .A(b[0]), .B(a[28]), .Z(n1197) );
  NAND U1552 ( .A(b[1]), .B(a[27]), .Z(n1196) );
  XNOR U1553 ( .A(n1197), .B(n1196), .Z(n1199) );
  XNOR U1554 ( .A(n1198), .B(n1199), .Z(n1203) );
  XNOR U1555 ( .A(n1202), .B(sreg[282]), .Z(n1195) );
  XNOR U1556 ( .A(n1203), .B(n1195), .Z(c[282]) );
  NAND U1557 ( .A(n1197), .B(n1196), .Z(n1201) );
  NANDN U1558 ( .A(n1199), .B(n1198), .Z(n1200) );
  NAND U1559 ( .A(n1201), .B(n1200), .Z(n1207) );
  NAND U1560 ( .A(b[0]), .B(a[29]), .Z(n1206) );
  NAND U1561 ( .A(b[1]), .B(a[28]), .Z(n1205) );
  XNOR U1562 ( .A(n1206), .B(n1205), .Z(n1208) );
  XNOR U1563 ( .A(n1207), .B(n1208), .Z(n1212) );
  XOR U1564 ( .A(n1211), .B(sreg[283]), .Z(n1204) );
  XNOR U1565 ( .A(n1212), .B(n1204), .Z(c[283]) );
  NAND U1566 ( .A(n1206), .B(n1205), .Z(n1210) );
  NANDN U1567 ( .A(n1208), .B(n1207), .Z(n1209) );
  NAND U1568 ( .A(n1210), .B(n1209), .Z(n1217) );
  ANDN U1569 ( .B(a[30]), .A(n965), .Z(n1215) );
  ANDN U1570 ( .B(a[29]), .A(n966), .Z(n1214) );
  XOR U1571 ( .A(n1215), .B(n1214), .Z(n1216) );
  XNOR U1572 ( .A(n1217), .B(n1216), .Z(n1219) );
  XOR U1573 ( .A(sreg[284]), .B(n1218), .Z(n1213) );
  XNOR U1574 ( .A(n1219), .B(n1213), .Z(c[284]) );
  NAND U1575 ( .A(b[0]), .B(a[31]), .Z(n1222) );
  NAND U1576 ( .A(b[1]), .B(a[30]), .Z(n1221) );
  XNOR U1577 ( .A(n1222), .B(n1221), .Z(n1224) );
  XNOR U1578 ( .A(n1223), .B(n1224), .Z(n1228) );
  XOR U1579 ( .A(n1227), .B(sreg[285]), .Z(n1220) );
  XNOR U1580 ( .A(n1228), .B(n1220), .Z(c[285]) );
  NAND U1581 ( .A(n1222), .B(n1221), .Z(n1226) );
  NANDN U1582 ( .A(n1224), .B(n1223), .Z(n1225) );
  NAND U1583 ( .A(n1226), .B(n1225), .Z(n1233) );
  ANDN U1584 ( .B(a[32]), .A(n965), .Z(n1231) );
  ANDN U1585 ( .B(a[31]), .A(n966), .Z(n1230) );
  XOR U1586 ( .A(n1231), .B(n1230), .Z(n1232) );
  XNOR U1587 ( .A(n1233), .B(n1232), .Z(n1235) );
  XOR U1588 ( .A(sreg[286]), .B(n1234), .Z(n1229) );
  XNOR U1589 ( .A(n1235), .B(n1229), .Z(c[286]) );
  NAND U1590 ( .A(b[0]), .B(a[33]), .Z(n1238) );
  NAND U1591 ( .A(b[1]), .B(a[32]), .Z(n1237) );
  XNOR U1592 ( .A(n1238), .B(n1237), .Z(n1240) );
  XNOR U1593 ( .A(n1239), .B(n1240), .Z(n1244) );
  XOR U1594 ( .A(n1243), .B(sreg[287]), .Z(n1236) );
  XNOR U1595 ( .A(n1244), .B(n1236), .Z(c[287]) );
  NAND U1596 ( .A(n1238), .B(n1237), .Z(n1242) );
  NANDN U1597 ( .A(n1240), .B(n1239), .Z(n1241) );
  NAND U1598 ( .A(n1242), .B(n1241), .Z(n1249) );
  ANDN U1599 ( .B(a[34]), .A(n965), .Z(n1247) );
  ANDN U1600 ( .B(a[33]), .A(n966), .Z(n1246) );
  XOR U1601 ( .A(n1247), .B(n1246), .Z(n1248) );
  XNOR U1602 ( .A(n1249), .B(n1248), .Z(n1251) );
  XOR U1603 ( .A(sreg[288]), .B(n1250), .Z(n1245) );
  XNOR U1604 ( .A(n1251), .B(n1245), .Z(c[288]) );
  NAND U1605 ( .A(b[0]), .B(a[35]), .Z(n1254) );
  NAND U1606 ( .A(b[1]), .B(a[34]), .Z(n1253) );
  XNOR U1607 ( .A(n1254), .B(n1253), .Z(n1256) );
  XNOR U1608 ( .A(n1255), .B(n1256), .Z(n1260) );
  XOR U1609 ( .A(n1259), .B(sreg[289]), .Z(n1252) );
  XNOR U1610 ( .A(n1260), .B(n1252), .Z(c[289]) );
  NAND U1611 ( .A(n1254), .B(n1253), .Z(n1258) );
  NANDN U1612 ( .A(n1256), .B(n1255), .Z(n1257) );
  NAND U1613 ( .A(n1258), .B(n1257), .Z(n1265) );
  ANDN U1614 ( .B(a[36]), .A(n965), .Z(n1263) );
  ANDN U1615 ( .B(a[35]), .A(n966), .Z(n1262) );
  XOR U1616 ( .A(n1263), .B(n1262), .Z(n1264) );
  XNOR U1617 ( .A(n1265), .B(n1264), .Z(n1267) );
  XOR U1618 ( .A(sreg[290]), .B(n1266), .Z(n1261) );
  XNOR U1619 ( .A(n1267), .B(n1261), .Z(c[290]) );
  NAND U1620 ( .A(b[0]), .B(a[37]), .Z(n1270) );
  NAND U1621 ( .A(b[1]), .B(a[36]), .Z(n1269) );
  XNOR U1622 ( .A(n1270), .B(n1269), .Z(n1272) );
  XNOR U1623 ( .A(n1271), .B(n1272), .Z(n1276) );
  XOR U1624 ( .A(n1275), .B(sreg[291]), .Z(n1268) );
  XNOR U1625 ( .A(n1276), .B(n1268), .Z(c[291]) );
  NAND U1626 ( .A(n1270), .B(n1269), .Z(n1274) );
  NANDN U1627 ( .A(n1272), .B(n1271), .Z(n1273) );
  NAND U1628 ( .A(n1274), .B(n1273), .Z(n1281) );
  ANDN U1629 ( .B(a[38]), .A(n965), .Z(n1279) );
  ANDN U1630 ( .B(a[37]), .A(n966), .Z(n1278) );
  XOR U1631 ( .A(n1279), .B(n1278), .Z(n1280) );
  XNOR U1632 ( .A(n1281), .B(n1280), .Z(n1283) );
  XOR U1633 ( .A(sreg[292]), .B(n1282), .Z(n1277) );
  XNOR U1634 ( .A(n1283), .B(n1277), .Z(c[292]) );
  NAND U1635 ( .A(b[0]), .B(a[39]), .Z(n1286) );
  NAND U1636 ( .A(b[1]), .B(a[38]), .Z(n1285) );
  XNOR U1637 ( .A(n1286), .B(n1285), .Z(n1288) );
  XNOR U1638 ( .A(n1287), .B(n1288), .Z(n1292) );
  XOR U1639 ( .A(n1291), .B(sreg[293]), .Z(n1284) );
  XNOR U1640 ( .A(n1292), .B(n1284), .Z(c[293]) );
  NAND U1641 ( .A(n1286), .B(n1285), .Z(n1290) );
  NANDN U1642 ( .A(n1288), .B(n1287), .Z(n1289) );
  NAND U1643 ( .A(n1290), .B(n1289), .Z(n1297) );
  ANDN U1644 ( .B(a[40]), .A(n965), .Z(n1295) );
  ANDN U1645 ( .B(a[39]), .A(n966), .Z(n1294) );
  XOR U1646 ( .A(n1295), .B(n1294), .Z(n1296) );
  XNOR U1647 ( .A(n1297), .B(n1296), .Z(n1299) );
  XOR U1648 ( .A(sreg[294]), .B(n1298), .Z(n1293) );
  XNOR U1649 ( .A(n1299), .B(n1293), .Z(c[294]) );
  NAND U1650 ( .A(b[0]), .B(a[41]), .Z(n1302) );
  NAND U1651 ( .A(b[1]), .B(a[40]), .Z(n1301) );
  XNOR U1652 ( .A(n1302), .B(n1301), .Z(n1304) );
  XNOR U1653 ( .A(n1303), .B(n1304), .Z(n1308) );
  XOR U1654 ( .A(n1307), .B(sreg[295]), .Z(n1300) );
  XNOR U1655 ( .A(n1308), .B(n1300), .Z(c[295]) );
  NAND U1656 ( .A(n1302), .B(n1301), .Z(n1306) );
  NANDN U1657 ( .A(n1304), .B(n1303), .Z(n1305) );
  NAND U1658 ( .A(n1306), .B(n1305), .Z(n1313) );
  ANDN U1659 ( .B(a[42]), .A(n965), .Z(n1311) );
  ANDN U1660 ( .B(a[41]), .A(n966), .Z(n1310) );
  XOR U1661 ( .A(n1311), .B(n1310), .Z(n1312) );
  XNOR U1662 ( .A(n1313), .B(n1312), .Z(n1315) );
  XOR U1663 ( .A(sreg[296]), .B(n1314), .Z(n1309) );
  XNOR U1664 ( .A(n1315), .B(n1309), .Z(c[296]) );
  NAND U1665 ( .A(b[0]), .B(a[43]), .Z(n1318) );
  NAND U1666 ( .A(b[1]), .B(a[42]), .Z(n1317) );
  XNOR U1667 ( .A(n1318), .B(n1317), .Z(n1320) );
  XNOR U1668 ( .A(n1319), .B(n1320), .Z(n1324) );
  XOR U1669 ( .A(n1323), .B(sreg[297]), .Z(n1316) );
  XNOR U1670 ( .A(n1324), .B(n1316), .Z(c[297]) );
  NAND U1671 ( .A(n1318), .B(n1317), .Z(n1322) );
  NANDN U1672 ( .A(n1320), .B(n1319), .Z(n1321) );
  NAND U1673 ( .A(n1322), .B(n1321), .Z(n1329) );
  ANDN U1674 ( .B(a[44]), .A(n965), .Z(n1327) );
  ANDN U1675 ( .B(a[43]), .A(n966), .Z(n1326) );
  XOR U1676 ( .A(n1327), .B(n1326), .Z(n1328) );
  XNOR U1677 ( .A(n1329), .B(n1328), .Z(n1331) );
  XOR U1678 ( .A(sreg[298]), .B(n1330), .Z(n1325) );
  XNOR U1679 ( .A(n1331), .B(n1325), .Z(c[298]) );
  NAND U1680 ( .A(b[0]), .B(a[45]), .Z(n1334) );
  NAND U1681 ( .A(b[1]), .B(a[44]), .Z(n1333) );
  XNOR U1682 ( .A(n1334), .B(n1333), .Z(n1336) );
  XNOR U1683 ( .A(n1335), .B(n1336), .Z(n1340) );
  XOR U1684 ( .A(n1339), .B(sreg[299]), .Z(n1332) );
  XNOR U1685 ( .A(n1340), .B(n1332), .Z(c[299]) );
  NAND U1686 ( .A(n1334), .B(n1333), .Z(n1338) );
  NANDN U1687 ( .A(n1336), .B(n1335), .Z(n1337) );
  NAND U1688 ( .A(n1338), .B(n1337), .Z(n1345) );
  ANDN U1689 ( .B(a[46]), .A(n965), .Z(n1343) );
  ANDN U1690 ( .B(a[45]), .A(n966), .Z(n1342) );
  XOR U1691 ( .A(n1343), .B(n1342), .Z(n1344) );
  XNOR U1692 ( .A(n1345), .B(n1344), .Z(n1347) );
  XOR U1693 ( .A(sreg[300]), .B(n1346), .Z(n1341) );
  XNOR U1694 ( .A(n1347), .B(n1341), .Z(c[300]) );
  ANDN U1695 ( .B(a[47]), .A(n965), .Z(n1350) );
  ANDN U1696 ( .B(a[46]), .A(n966), .Z(n1349) );
  XOR U1697 ( .A(n1350), .B(n1349), .Z(n1351) );
  XNOR U1698 ( .A(n1352), .B(n1351), .Z(n1354) );
  XNOR U1699 ( .A(sreg[301]), .B(n1353), .Z(n1348) );
  XNOR U1700 ( .A(n1354), .B(n1348), .Z(c[301]) );
  NAND U1701 ( .A(b[0]), .B(a[48]), .Z(n1357) );
  NAND U1702 ( .A(b[1]), .B(a[47]), .Z(n1356) );
  XNOR U1703 ( .A(n1357), .B(n1356), .Z(n1359) );
  XNOR U1704 ( .A(n1358), .B(n1359), .Z(n1363) );
  XOR U1705 ( .A(n1362), .B(sreg[302]), .Z(n1355) );
  XNOR U1706 ( .A(n1363), .B(n1355), .Z(c[302]) );
  NAND U1707 ( .A(n1357), .B(n1356), .Z(n1361) );
  NANDN U1708 ( .A(n1359), .B(n1358), .Z(n1360) );
  NAND U1709 ( .A(n1361), .B(n1360), .Z(n1367) );
  NAND U1710 ( .A(b[0]), .B(a[49]), .Z(n1366) );
  NAND U1711 ( .A(b[1]), .B(a[48]), .Z(n1365) );
  XNOR U1712 ( .A(n1366), .B(n1365), .Z(n1368) );
  XNOR U1713 ( .A(n1367), .B(n1368), .Z(n1372) );
  XOR U1714 ( .A(n1371), .B(sreg[303]), .Z(n1364) );
  XNOR U1715 ( .A(n1372), .B(n1364), .Z(c[303]) );
  NAND U1716 ( .A(n1366), .B(n1365), .Z(n1370) );
  NANDN U1717 ( .A(n1368), .B(n1367), .Z(n1369) );
  NAND U1718 ( .A(n1370), .B(n1369), .Z(n1377) );
  ANDN U1719 ( .B(a[50]), .A(n965), .Z(n1375) );
  ANDN U1720 ( .B(a[49]), .A(n966), .Z(n1374) );
  XOR U1721 ( .A(n1375), .B(n1374), .Z(n1376) );
  XNOR U1722 ( .A(n1377), .B(n1376), .Z(n1379) );
  XOR U1723 ( .A(sreg[304]), .B(n1378), .Z(n1373) );
  XNOR U1724 ( .A(n1379), .B(n1373), .Z(c[304]) );
  NAND U1725 ( .A(b[0]), .B(a[51]), .Z(n1382) );
  NAND U1726 ( .A(b[1]), .B(a[50]), .Z(n1381) );
  XNOR U1727 ( .A(n1382), .B(n1381), .Z(n1384) );
  XNOR U1728 ( .A(n1383), .B(n1384), .Z(n1388) );
  XOR U1729 ( .A(n1387), .B(sreg[305]), .Z(n1380) );
  XNOR U1730 ( .A(n1388), .B(n1380), .Z(c[305]) );
  NAND U1731 ( .A(n1382), .B(n1381), .Z(n1386) );
  NANDN U1732 ( .A(n1384), .B(n1383), .Z(n1385) );
  NAND U1733 ( .A(n1386), .B(n1385), .Z(n1393) );
  ANDN U1734 ( .B(a[52]), .A(n965), .Z(n1391) );
  ANDN U1735 ( .B(a[51]), .A(n966), .Z(n1390) );
  XOR U1736 ( .A(n1391), .B(n1390), .Z(n1392) );
  XNOR U1737 ( .A(n1393), .B(n1392), .Z(n1395) );
  XOR U1738 ( .A(sreg[306]), .B(n1394), .Z(n1389) );
  XNOR U1739 ( .A(n1395), .B(n1389), .Z(c[306]) );
  ANDN U1740 ( .B(a[53]), .A(n965), .Z(n1398) );
  ANDN U1741 ( .B(a[52]), .A(n966), .Z(n1397) );
  XOR U1742 ( .A(n1398), .B(n1397), .Z(n1399) );
  XNOR U1743 ( .A(n1400), .B(n1399), .Z(n1402) );
  XNOR U1744 ( .A(sreg[307]), .B(n1401), .Z(n1396) );
  XNOR U1745 ( .A(n1402), .B(n1396), .Z(c[307]) );
  NAND U1746 ( .A(b[0]), .B(a[54]), .Z(n1405) );
  NAND U1747 ( .A(b[1]), .B(a[53]), .Z(n1404) );
  XNOR U1748 ( .A(n1405), .B(n1404), .Z(n1407) );
  XNOR U1749 ( .A(n1406), .B(n1407), .Z(n1411) );
  XOR U1750 ( .A(n1410), .B(sreg[308]), .Z(n1403) );
  XNOR U1751 ( .A(n1411), .B(n1403), .Z(c[308]) );
  NAND U1752 ( .A(n1405), .B(n1404), .Z(n1409) );
  NANDN U1753 ( .A(n1407), .B(n1406), .Z(n1408) );
  NAND U1754 ( .A(n1409), .B(n1408), .Z(n1415) );
  NAND U1755 ( .A(b[0]), .B(a[55]), .Z(n1414) );
  NAND U1756 ( .A(b[1]), .B(a[54]), .Z(n1413) );
  XNOR U1757 ( .A(n1414), .B(n1413), .Z(n1416) );
  XNOR U1758 ( .A(n1415), .B(n1416), .Z(n1420) );
  XOR U1759 ( .A(n1419), .B(sreg[309]), .Z(n1412) );
  XNOR U1760 ( .A(n1420), .B(n1412), .Z(c[309]) );
  NAND U1761 ( .A(n1414), .B(n1413), .Z(n1418) );
  NANDN U1762 ( .A(n1416), .B(n1415), .Z(n1417) );
  NAND U1763 ( .A(n1418), .B(n1417), .Z(n1425) );
  ANDN U1764 ( .B(a[56]), .A(n965), .Z(n1423) );
  ANDN U1765 ( .B(a[55]), .A(n966), .Z(n1422) );
  XOR U1766 ( .A(n1423), .B(n1422), .Z(n1424) );
  XNOR U1767 ( .A(n1425), .B(n1424), .Z(n1427) );
  XOR U1768 ( .A(sreg[310]), .B(n1426), .Z(n1421) );
  XNOR U1769 ( .A(n1427), .B(n1421), .Z(c[310]) );
  NAND U1770 ( .A(b[0]), .B(a[57]), .Z(n1430) );
  NAND U1771 ( .A(b[1]), .B(a[56]), .Z(n1429) );
  XNOR U1772 ( .A(n1430), .B(n1429), .Z(n1432) );
  XNOR U1773 ( .A(n1431), .B(n1432), .Z(n1436) );
  XOR U1774 ( .A(n1435), .B(sreg[311]), .Z(n1428) );
  XNOR U1775 ( .A(n1436), .B(n1428), .Z(c[311]) );
  NAND U1776 ( .A(n1430), .B(n1429), .Z(n1434) );
  NANDN U1777 ( .A(n1432), .B(n1431), .Z(n1433) );
  NAND U1778 ( .A(n1434), .B(n1433), .Z(n1441) );
  ANDN U1779 ( .B(a[58]), .A(n965), .Z(n1439) );
  ANDN U1780 ( .B(a[57]), .A(n966), .Z(n1438) );
  XOR U1781 ( .A(n1439), .B(n1438), .Z(n1440) );
  XNOR U1782 ( .A(n1441), .B(n1440), .Z(n1443) );
  XOR U1783 ( .A(sreg[312]), .B(n1442), .Z(n1437) );
  XNOR U1784 ( .A(n1443), .B(n1437), .Z(c[312]) );
  NAND U1785 ( .A(b[0]), .B(a[59]), .Z(n1446) );
  NAND U1786 ( .A(b[1]), .B(a[58]), .Z(n1445) );
  XNOR U1787 ( .A(n1446), .B(n1445), .Z(n1448) );
  XNOR U1788 ( .A(n1447), .B(n1448), .Z(n1452) );
  XOR U1789 ( .A(n1451), .B(sreg[313]), .Z(n1444) );
  XNOR U1790 ( .A(n1452), .B(n1444), .Z(c[313]) );
  NAND U1791 ( .A(n1446), .B(n1445), .Z(n1450) );
  NANDN U1792 ( .A(n1448), .B(n1447), .Z(n1449) );
  NAND U1793 ( .A(n1450), .B(n1449), .Z(n1457) );
  ANDN U1794 ( .B(a[60]), .A(n965), .Z(n1455) );
  ANDN U1795 ( .B(a[59]), .A(n966), .Z(n1454) );
  XOR U1796 ( .A(n1455), .B(n1454), .Z(n1456) );
  XNOR U1797 ( .A(n1457), .B(n1456), .Z(n1459) );
  XOR U1798 ( .A(sreg[314]), .B(n1458), .Z(n1453) );
  XNOR U1799 ( .A(n1459), .B(n1453), .Z(c[314]) );
  NAND U1800 ( .A(b[0]), .B(a[61]), .Z(n1462) );
  NAND U1801 ( .A(b[1]), .B(a[60]), .Z(n1461) );
  XNOR U1802 ( .A(n1462), .B(n1461), .Z(n1464) );
  XNOR U1803 ( .A(n1463), .B(n1464), .Z(n1468) );
  XOR U1804 ( .A(n1467), .B(sreg[315]), .Z(n1460) );
  XNOR U1805 ( .A(n1468), .B(n1460), .Z(c[315]) );
  NAND U1806 ( .A(n1462), .B(n1461), .Z(n1466) );
  NANDN U1807 ( .A(n1464), .B(n1463), .Z(n1465) );
  NAND U1808 ( .A(n1466), .B(n1465), .Z(n1473) );
  ANDN U1809 ( .B(a[62]), .A(n965), .Z(n1471) );
  ANDN U1810 ( .B(a[61]), .A(n966), .Z(n1470) );
  XOR U1811 ( .A(n1471), .B(n1470), .Z(n1472) );
  XNOR U1812 ( .A(n1473), .B(n1472), .Z(n1475) );
  XOR U1813 ( .A(sreg[316]), .B(n1474), .Z(n1469) );
  XNOR U1814 ( .A(n1475), .B(n1469), .Z(c[316]) );
  NAND U1815 ( .A(b[0]), .B(a[63]), .Z(n1478) );
  NAND U1816 ( .A(b[1]), .B(a[62]), .Z(n1477) );
  XNOR U1817 ( .A(n1478), .B(n1477), .Z(n1480) );
  XNOR U1818 ( .A(n1479), .B(n1480), .Z(n1484) );
  XOR U1819 ( .A(n1483), .B(sreg[317]), .Z(n1476) );
  XNOR U1820 ( .A(n1484), .B(n1476), .Z(c[317]) );
  NAND U1821 ( .A(n1478), .B(n1477), .Z(n1482) );
  NANDN U1822 ( .A(n1480), .B(n1479), .Z(n1481) );
  NAND U1823 ( .A(n1482), .B(n1481), .Z(n1489) );
  ANDN U1824 ( .B(a[64]), .A(n965), .Z(n1487) );
  ANDN U1825 ( .B(a[63]), .A(n966), .Z(n1486) );
  XOR U1826 ( .A(n1487), .B(n1486), .Z(n1488) );
  XNOR U1827 ( .A(n1489), .B(n1488), .Z(n1491) );
  XOR U1828 ( .A(sreg[318]), .B(n1490), .Z(n1485) );
  XNOR U1829 ( .A(n1491), .B(n1485), .Z(c[318]) );
  NAND U1830 ( .A(b[0]), .B(a[65]), .Z(n1494) );
  NAND U1831 ( .A(b[1]), .B(a[64]), .Z(n1493) );
  XNOR U1832 ( .A(n1494), .B(n1493), .Z(n1496) );
  XNOR U1833 ( .A(n1495), .B(n1496), .Z(n1500) );
  XOR U1834 ( .A(n1499), .B(sreg[319]), .Z(n1492) );
  XNOR U1835 ( .A(n1500), .B(n1492), .Z(c[319]) );
  NAND U1836 ( .A(n1494), .B(n1493), .Z(n1498) );
  NANDN U1837 ( .A(n1496), .B(n1495), .Z(n1497) );
  NAND U1838 ( .A(n1498), .B(n1497), .Z(n1504) );
  NAND U1839 ( .A(b[0]), .B(a[66]), .Z(n1503) );
  NAND U1840 ( .A(b[1]), .B(a[65]), .Z(n1502) );
  XNOR U1841 ( .A(n1503), .B(n1502), .Z(n1505) );
  XNOR U1842 ( .A(n1504), .B(n1505), .Z(n1509) );
  XOR U1843 ( .A(n1508), .B(sreg[320]), .Z(n1501) );
  XNOR U1844 ( .A(n1509), .B(n1501), .Z(c[320]) );
  NAND U1845 ( .A(n1503), .B(n1502), .Z(n1507) );
  NANDN U1846 ( .A(n1505), .B(n1504), .Z(n1506) );
  NAND U1847 ( .A(n1507), .B(n1506), .Z(n1513) );
  NAND U1848 ( .A(b[0]), .B(a[67]), .Z(n1512) );
  NAND U1849 ( .A(b[1]), .B(a[66]), .Z(n1511) );
  XNOR U1850 ( .A(n1512), .B(n1511), .Z(n1514) );
  XNOR U1851 ( .A(n1513), .B(n1514), .Z(n1518) );
  XOR U1852 ( .A(n1517), .B(sreg[321]), .Z(n1510) );
  XNOR U1853 ( .A(n1518), .B(n1510), .Z(c[321]) );
  NAND U1854 ( .A(n1512), .B(n1511), .Z(n1516) );
  NANDN U1855 ( .A(n1514), .B(n1513), .Z(n1515) );
  NAND U1856 ( .A(n1516), .B(n1515), .Z(n1523) );
  ANDN U1857 ( .B(a[68]), .A(n965), .Z(n1521) );
  ANDN U1858 ( .B(a[67]), .A(n966), .Z(n1520) );
  XOR U1859 ( .A(n1521), .B(n1520), .Z(n1522) );
  XNOR U1860 ( .A(n1523), .B(n1522), .Z(n1525) );
  XOR U1861 ( .A(sreg[322]), .B(n1524), .Z(n1519) );
  XNOR U1862 ( .A(n1525), .B(n1519), .Z(c[322]) );
  NAND U1863 ( .A(b[0]), .B(a[69]), .Z(n1528) );
  NAND U1864 ( .A(b[1]), .B(a[68]), .Z(n1527) );
  XNOR U1865 ( .A(n1528), .B(n1527), .Z(n1530) );
  XNOR U1866 ( .A(n1529), .B(n1530), .Z(n1534) );
  XOR U1867 ( .A(n1533), .B(sreg[323]), .Z(n1526) );
  XNOR U1868 ( .A(n1534), .B(n1526), .Z(c[323]) );
  NAND U1869 ( .A(n1528), .B(n1527), .Z(n1532) );
  NANDN U1870 ( .A(n1530), .B(n1529), .Z(n1531) );
  NAND U1871 ( .A(n1532), .B(n1531), .Z(n1539) );
  ANDN U1872 ( .B(a[70]), .A(n965), .Z(n1537) );
  ANDN U1873 ( .B(a[69]), .A(n966), .Z(n1536) );
  XOR U1874 ( .A(n1537), .B(n1536), .Z(n1538) );
  XNOR U1875 ( .A(n1539), .B(n1538), .Z(n1541) );
  XOR U1876 ( .A(sreg[324]), .B(n1540), .Z(n1535) );
  XNOR U1877 ( .A(n1541), .B(n1535), .Z(c[324]) );
  NAND U1878 ( .A(b[0]), .B(a[71]), .Z(n1544) );
  NAND U1879 ( .A(b[1]), .B(a[70]), .Z(n1543) );
  XNOR U1880 ( .A(n1544), .B(n1543), .Z(n1546) );
  XNOR U1881 ( .A(n1545), .B(n1546), .Z(n1550) );
  XOR U1882 ( .A(n1549), .B(sreg[325]), .Z(n1542) );
  XNOR U1883 ( .A(n1550), .B(n1542), .Z(c[325]) );
  NAND U1884 ( .A(n1544), .B(n1543), .Z(n1548) );
  NANDN U1885 ( .A(n1546), .B(n1545), .Z(n1547) );
  NAND U1886 ( .A(n1548), .B(n1547), .Z(n1554) );
  NAND U1887 ( .A(b[0]), .B(a[72]), .Z(n1553) );
  NAND U1888 ( .A(b[1]), .B(a[71]), .Z(n1552) );
  XNOR U1889 ( .A(n1553), .B(n1552), .Z(n1555) );
  XNOR U1890 ( .A(n1554), .B(n1555), .Z(n1559) );
  XOR U1891 ( .A(n1558), .B(sreg[326]), .Z(n1551) );
  XNOR U1892 ( .A(n1559), .B(n1551), .Z(c[326]) );
  NAND U1893 ( .A(n1553), .B(n1552), .Z(n1557) );
  NANDN U1894 ( .A(n1555), .B(n1554), .Z(n1556) );
  NAND U1895 ( .A(n1557), .B(n1556), .Z(n1563) );
  NAND U1896 ( .A(b[0]), .B(a[73]), .Z(n1562) );
  NAND U1897 ( .A(b[1]), .B(a[72]), .Z(n1561) );
  XNOR U1898 ( .A(n1562), .B(n1561), .Z(n1564) );
  XNOR U1899 ( .A(n1563), .B(n1564), .Z(n1568) );
  XOR U1900 ( .A(n1567), .B(sreg[327]), .Z(n1560) );
  XNOR U1901 ( .A(n1568), .B(n1560), .Z(c[327]) );
  NAND U1902 ( .A(n1562), .B(n1561), .Z(n1566) );
  NANDN U1903 ( .A(n1564), .B(n1563), .Z(n1565) );
  NAND U1904 ( .A(n1566), .B(n1565), .Z(n1572) );
  NAND U1905 ( .A(b[0]), .B(a[74]), .Z(n1571) );
  NAND U1906 ( .A(b[1]), .B(a[73]), .Z(n1570) );
  XNOR U1907 ( .A(n1571), .B(n1570), .Z(n1573) );
  XNOR U1908 ( .A(n1572), .B(n1573), .Z(n1577) );
  XOR U1909 ( .A(n1576), .B(sreg[328]), .Z(n1569) );
  XNOR U1910 ( .A(n1577), .B(n1569), .Z(c[328]) );
  NAND U1911 ( .A(n1571), .B(n1570), .Z(n1575) );
  NANDN U1912 ( .A(n1573), .B(n1572), .Z(n1574) );
  NAND U1913 ( .A(n1575), .B(n1574), .Z(n1581) );
  NAND U1914 ( .A(b[0]), .B(a[75]), .Z(n1580) );
  NAND U1915 ( .A(b[1]), .B(a[74]), .Z(n1579) );
  XNOR U1916 ( .A(n1580), .B(n1579), .Z(n1582) );
  XNOR U1917 ( .A(n1581), .B(n1582), .Z(n1586) );
  XOR U1918 ( .A(n1585), .B(sreg[329]), .Z(n1578) );
  XNOR U1919 ( .A(n1586), .B(n1578), .Z(c[329]) );
  NAND U1920 ( .A(n1580), .B(n1579), .Z(n1584) );
  NANDN U1921 ( .A(n1582), .B(n1581), .Z(n1583) );
  NAND U1922 ( .A(n1584), .B(n1583), .Z(n1591) );
  ANDN U1923 ( .B(a[76]), .A(n965), .Z(n1589) );
  ANDN U1924 ( .B(a[75]), .A(n966), .Z(n1588) );
  XOR U1925 ( .A(n1589), .B(n1588), .Z(n1590) );
  XNOR U1926 ( .A(n1591), .B(n1590), .Z(n1593) );
  XOR U1927 ( .A(sreg[330]), .B(n1592), .Z(n1587) );
  XNOR U1928 ( .A(n1593), .B(n1587), .Z(c[330]) );
  NAND U1929 ( .A(b[0]), .B(a[77]), .Z(n1596) );
  NAND U1930 ( .A(b[1]), .B(a[76]), .Z(n1595) );
  XNOR U1931 ( .A(n1596), .B(n1595), .Z(n1598) );
  XNOR U1932 ( .A(n1597), .B(n1598), .Z(n1602) );
  XOR U1933 ( .A(n1601), .B(sreg[331]), .Z(n1594) );
  XNOR U1934 ( .A(n1602), .B(n1594), .Z(c[331]) );
  NAND U1935 ( .A(n1596), .B(n1595), .Z(n1600) );
  NANDN U1936 ( .A(n1598), .B(n1597), .Z(n1599) );
  NAND U1937 ( .A(n1600), .B(n1599), .Z(n1607) );
  ANDN U1938 ( .B(a[78]), .A(n965), .Z(n1605) );
  ANDN U1939 ( .B(a[77]), .A(n966), .Z(n1604) );
  XOR U1940 ( .A(n1605), .B(n1604), .Z(n1606) );
  XNOR U1941 ( .A(n1607), .B(n1606), .Z(n1609) );
  XOR U1942 ( .A(sreg[332]), .B(n1608), .Z(n1603) );
  XNOR U1943 ( .A(n1609), .B(n1603), .Z(c[332]) );
  NAND U1944 ( .A(b[0]), .B(a[79]), .Z(n1612) );
  NAND U1945 ( .A(b[1]), .B(a[78]), .Z(n1611) );
  XNOR U1946 ( .A(n1612), .B(n1611), .Z(n1614) );
  XNOR U1947 ( .A(n1613), .B(n1614), .Z(n1618) );
  XOR U1948 ( .A(n1617), .B(sreg[333]), .Z(n1610) );
  XNOR U1949 ( .A(n1618), .B(n1610), .Z(c[333]) );
  NAND U1950 ( .A(n1612), .B(n1611), .Z(n1616) );
  NANDN U1951 ( .A(n1614), .B(n1613), .Z(n1615) );
  NAND U1952 ( .A(n1616), .B(n1615), .Z(n1623) );
  ANDN U1953 ( .B(a[80]), .A(n965), .Z(n1621) );
  ANDN U1954 ( .B(a[79]), .A(n966), .Z(n1620) );
  XOR U1955 ( .A(n1621), .B(n1620), .Z(n1622) );
  XNOR U1956 ( .A(n1623), .B(n1622), .Z(n1625) );
  XOR U1957 ( .A(sreg[334]), .B(n1624), .Z(n1619) );
  XNOR U1958 ( .A(n1625), .B(n1619), .Z(c[334]) );
  NAND U1959 ( .A(b[0]), .B(a[81]), .Z(n1628) );
  NAND U1960 ( .A(b[1]), .B(a[80]), .Z(n1627) );
  XNOR U1961 ( .A(n1628), .B(n1627), .Z(n1630) );
  XNOR U1962 ( .A(n1629), .B(n1630), .Z(n1634) );
  XOR U1963 ( .A(n1633), .B(sreg[335]), .Z(n1626) );
  XNOR U1964 ( .A(n1634), .B(n1626), .Z(c[335]) );
  NAND U1965 ( .A(n1628), .B(n1627), .Z(n1632) );
  NANDN U1966 ( .A(n1630), .B(n1629), .Z(n1631) );
  NAND U1967 ( .A(n1632), .B(n1631), .Z(n1639) );
  ANDN U1968 ( .B(a[82]), .A(n965), .Z(n1637) );
  ANDN U1969 ( .B(a[81]), .A(n966), .Z(n1636) );
  XOR U1970 ( .A(n1637), .B(n1636), .Z(n1638) );
  XNOR U1971 ( .A(n1639), .B(n1638), .Z(n1641) );
  XOR U1972 ( .A(sreg[336]), .B(n1640), .Z(n1635) );
  XNOR U1973 ( .A(n1641), .B(n1635), .Z(c[336]) );
  NAND U1974 ( .A(b[0]), .B(a[83]), .Z(n1644) );
  NAND U1975 ( .A(b[1]), .B(a[82]), .Z(n1643) );
  XNOR U1976 ( .A(n1644), .B(n1643), .Z(n1646) );
  XNOR U1977 ( .A(n1645), .B(n1646), .Z(n1650) );
  XOR U1978 ( .A(n1649), .B(sreg[337]), .Z(n1642) );
  XNOR U1979 ( .A(n1650), .B(n1642), .Z(c[337]) );
  NAND U1980 ( .A(n1644), .B(n1643), .Z(n1648) );
  NANDN U1981 ( .A(n1646), .B(n1645), .Z(n1647) );
  NAND U1982 ( .A(n1648), .B(n1647), .Z(n1655) );
  ANDN U1983 ( .B(a[84]), .A(n965), .Z(n1653) );
  ANDN U1984 ( .B(a[83]), .A(n966), .Z(n1652) );
  XOR U1985 ( .A(n1653), .B(n1652), .Z(n1654) );
  XNOR U1986 ( .A(n1655), .B(n1654), .Z(n1657) );
  XOR U1987 ( .A(sreg[338]), .B(n1656), .Z(n1651) );
  XNOR U1988 ( .A(n1657), .B(n1651), .Z(c[338]) );
  NAND U1989 ( .A(b[0]), .B(a[85]), .Z(n1660) );
  NAND U1990 ( .A(b[1]), .B(a[84]), .Z(n1659) );
  XNOR U1991 ( .A(n1660), .B(n1659), .Z(n1662) );
  XNOR U1992 ( .A(n1661), .B(n1662), .Z(n1666) );
  XOR U1993 ( .A(n1665), .B(sreg[339]), .Z(n1658) );
  XNOR U1994 ( .A(n1666), .B(n1658), .Z(c[339]) );
  NAND U1995 ( .A(n1660), .B(n1659), .Z(n1664) );
  NANDN U1996 ( .A(n1662), .B(n1661), .Z(n1663) );
  NAND U1997 ( .A(n1664), .B(n1663), .Z(n1671) );
  ANDN U1998 ( .B(a[86]), .A(n965), .Z(n1669) );
  ANDN U1999 ( .B(a[85]), .A(n966), .Z(n1668) );
  XOR U2000 ( .A(n1669), .B(n1668), .Z(n1670) );
  XNOR U2001 ( .A(n1671), .B(n1670), .Z(n1673) );
  XOR U2002 ( .A(sreg[340]), .B(n1672), .Z(n1667) );
  XNOR U2003 ( .A(n1673), .B(n1667), .Z(c[340]) );
  NAND U2004 ( .A(b[0]), .B(a[87]), .Z(n1676) );
  NAND U2005 ( .A(b[1]), .B(a[86]), .Z(n1675) );
  XNOR U2006 ( .A(n1676), .B(n1675), .Z(n1678) );
  XNOR U2007 ( .A(n1677), .B(n1678), .Z(n1682) );
  XOR U2008 ( .A(n1681), .B(sreg[341]), .Z(n1674) );
  XNOR U2009 ( .A(n1682), .B(n1674), .Z(c[341]) );
  NAND U2010 ( .A(n1676), .B(n1675), .Z(n1680) );
  NANDN U2011 ( .A(n1678), .B(n1677), .Z(n1679) );
  NAND U2012 ( .A(n1680), .B(n1679), .Z(n1686) );
  NAND U2013 ( .A(b[0]), .B(a[88]), .Z(n1685) );
  NAND U2014 ( .A(b[1]), .B(a[87]), .Z(n1684) );
  XNOR U2015 ( .A(n1685), .B(n1684), .Z(n1687) );
  XNOR U2016 ( .A(n1686), .B(n1687), .Z(n1691) );
  XOR U2017 ( .A(n1690), .B(sreg[342]), .Z(n1683) );
  XNOR U2018 ( .A(n1691), .B(n1683), .Z(c[342]) );
  NAND U2019 ( .A(n1685), .B(n1684), .Z(n1689) );
  NANDN U2020 ( .A(n1687), .B(n1686), .Z(n1688) );
  NAND U2021 ( .A(n1689), .B(n1688), .Z(n1695) );
  NAND U2022 ( .A(b[0]), .B(a[89]), .Z(n1694) );
  NAND U2023 ( .A(b[1]), .B(a[88]), .Z(n1693) );
  XNOR U2024 ( .A(n1694), .B(n1693), .Z(n1696) );
  XNOR U2025 ( .A(n1695), .B(n1696), .Z(n1700) );
  XOR U2026 ( .A(n1699), .B(sreg[343]), .Z(n1692) );
  XNOR U2027 ( .A(n1700), .B(n1692), .Z(c[343]) );
  NAND U2028 ( .A(n1694), .B(n1693), .Z(n1698) );
  NANDN U2029 ( .A(n1696), .B(n1695), .Z(n1697) );
  NAND U2030 ( .A(n1698), .B(n1697), .Z(n1705) );
  ANDN U2031 ( .B(a[90]), .A(n965), .Z(n1703) );
  ANDN U2032 ( .B(a[89]), .A(n966), .Z(n1702) );
  XOR U2033 ( .A(n1703), .B(n1702), .Z(n1704) );
  XNOR U2034 ( .A(n1705), .B(n1704), .Z(n1707) );
  XOR U2035 ( .A(sreg[344]), .B(n1706), .Z(n1701) );
  XNOR U2036 ( .A(n1707), .B(n1701), .Z(c[344]) );
  NAND U2037 ( .A(b[0]), .B(a[91]), .Z(n1710) );
  NAND U2038 ( .A(b[1]), .B(a[90]), .Z(n1709) );
  XNOR U2039 ( .A(n1710), .B(n1709), .Z(n1712) );
  XNOR U2040 ( .A(n1711), .B(n1712), .Z(n1716) );
  XOR U2041 ( .A(n1715), .B(sreg[345]), .Z(n1708) );
  XNOR U2042 ( .A(n1716), .B(n1708), .Z(c[345]) );
  NAND U2043 ( .A(n1710), .B(n1709), .Z(n1714) );
  NANDN U2044 ( .A(n1712), .B(n1711), .Z(n1713) );
  NAND U2045 ( .A(n1714), .B(n1713), .Z(n1720) );
  NAND U2046 ( .A(b[0]), .B(a[92]), .Z(n1719) );
  NAND U2047 ( .A(b[1]), .B(a[91]), .Z(n1718) );
  XNOR U2048 ( .A(n1719), .B(n1718), .Z(n1721) );
  XNOR U2049 ( .A(n1720), .B(n1721), .Z(n1725) );
  XOR U2050 ( .A(n1724), .B(sreg[346]), .Z(n1717) );
  XNOR U2051 ( .A(n1725), .B(n1717), .Z(c[346]) );
  NAND U2052 ( .A(n1719), .B(n1718), .Z(n1723) );
  NANDN U2053 ( .A(n1721), .B(n1720), .Z(n1722) );
  NAND U2054 ( .A(n1723), .B(n1722), .Z(n1729) );
  NAND U2055 ( .A(b[0]), .B(a[93]), .Z(n1728) );
  NAND U2056 ( .A(b[1]), .B(a[92]), .Z(n1727) );
  XNOR U2057 ( .A(n1728), .B(n1727), .Z(n1730) );
  XNOR U2058 ( .A(n1729), .B(n1730), .Z(n1734) );
  XOR U2059 ( .A(n1733), .B(sreg[347]), .Z(n1726) );
  XNOR U2060 ( .A(n1734), .B(n1726), .Z(c[347]) );
  NAND U2061 ( .A(n1728), .B(n1727), .Z(n1732) );
  NANDN U2062 ( .A(n1730), .B(n1729), .Z(n1731) );
  NAND U2063 ( .A(n1732), .B(n1731), .Z(n1739) );
  ANDN U2064 ( .B(a[94]), .A(n965), .Z(n1737) );
  ANDN U2065 ( .B(a[93]), .A(n966), .Z(n1736) );
  XOR U2066 ( .A(n1737), .B(n1736), .Z(n1738) );
  XNOR U2067 ( .A(n1739), .B(n1738), .Z(n1741) );
  XOR U2068 ( .A(sreg[348]), .B(n1740), .Z(n1735) );
  XNOR U2069 ( .A(n1741), .B(n1735), .Z(c[348]) );
  NAND U2070 ( .A(b[0]), .B(a[95]), .Z(n1744) );
  NAND U2071 ( .A(b[1]), .B(a[94]), .Z(n1743) );
  XNOR U2072 ( .A(n1744), .B(n1743), .Z(n1746) );
  XNOR U2073 ( .A(n1745), .B(n1746), .Z(n1750) );
  XOR U2074 ( .A(n1749), .B(sreg[349]), .Z(n1742) );
  XNOR U2075 ( .A(n1750), .B(n1742), .Z(c[349]) );
  NAND U2076 ( .A(n1744), .B(n1743), .Z(n1748) );
  NANDN U2077 ( .A(n1746), .B(n1745), .Z(n1747) );
  NAND U2078 ( .A(n1748), .B(n1747), .Z(n1754) );
  NAND U2079 ( .A(b[0]), .B(a[96]), .Z(n1753) );
  NAND U2080 ( .A(b[1]), .B(a[95]), .Z(n1752) );
  XNOR U2081 ( .A(n1753), .B(n1752), .Z(n1755) );
  XNOR U2082 ( .A(n1754), .B(n1755), .Z(n1759) );
  XOR U2083 ( .A(n1758), .B(sreg[350]), .Z(n1751) );
  XNOR U2084 ( .A(n1759), .B(n1751), .Z(c[350]) );
  NAND U2085 ( .A(n1753), .B(n1752), .Z(n1757) );
  NANDN U2086 ( .A(n1755), .B(n1754), .Z(n1756) );
  NAND U2087 ( .A(n1757), .B(n1756), .Z(n1763) );
  NAND U2088 ( .A(b[0]), .B(a[97]), .Z(n1762) );
  NAND U2089 ( .A(b[1]), .B(a[96]), .Z(n1761) );
  XNOR U2090 ( .A(n1762), .B(n1761), .Z(n1764) );
  XNOR U2091 ( .A(n1763), .B(n1764), .Z(n1768) );
  XOR U2092 ( .A(n1767), .B(sreg[351]), .Z(n1760) );
  XNOR U2093 ( .A(n1768), .B(n1760), .Z(c[351]) );
  NAND U2094 ( .A(n1762), .B(n1761), .Z(n1766) );
  NANDN U2095 ( .A(n1764), .B(n1763), .Z(n1765) );
  NAND U2096 ( .A(n1766), .B(n1765), .Z(n1772) );
  NAND U2097 ( .A(b[0]), .B(a[98]), .Z(n1771) );
  NAND U2098 ( .A(b[1]), .B(a[97]), .Z(n1770) );
  XNOR U2099 ( .A(n1771), .B(n1770), .Z(n1773) );
  XNOR U2100 ( .A(n1772), .B(n1773), .Z(n1777) );
  XOR U2101 ( .A(n1776), .B(sreg[352]), .Z(n1769) );
  XNOR U2102 ( .A(n1777), .B(n1769), .Z(c[352]) );
  NAND U2103 ( .A(n1771), .B(n1770), .Z(n1775) );
  NANDN U2104 ( .A(n1773), .B(n1772), .Z(n1774) );
  NAND U2105 ( .A(n1775), .B(n1774), .Z(n1781) );
  NAND U2106 ( .A(b[0]), .B(a[99]), .Z(n1780) );
  NAND U2107 ( .A(b[1]), .B(a[98]), .Z(n1779) );
  XNOR U2108 ( .A(n1780), .B(n1779), .Z(n1782) );
  XNOR U2109 ( .A(n1781), .B(n1782), .Z(n1786) );
  XOR U2110 ( .A(n1785), .B(sreg[353]), .Z(n1778) );
  XNOR U2111 ( .A(n1786), .B(n1778), .Z(c[353]) );
  NAND U2112 ( .A(n1780), .B(n1779), .Z(n1784) );
  NANDN U2113 ( .A(n1782), .B(n1781), .Z(n1783) );
  NAND U2114 ( .A(n1784), .B(n1783), .Z(n1790) );
  NAND U2115 ( .A(b[0]), .B(a[100]), .Z(n1789) );
  NAND U2116 ( .A(b[1]), .B(a[99]), .Z(n1788) );
  XNOR U2117 ( .A(n1789), .B(n1788), .Z(n1791) );
  XNOR U2118 ( .A(n1790), .B(n1791), .Z(n1795) );
  XOR U2119 ( .A(n1794), .B(sreg[354]), .Z(n1787) );
  XNOR U2120 ( .A(n1795), .B(n1787), .Z(c[354]) );
  NAND U2121 ( .A(n1789), .B(n1788), .Z(n1793) );
  NANDN U2122 ( .A(n1791), .B(n1790), .Z(n1792) );
  NAND U2123 ( .A(n1793), .B(n1792), .Z(n1799) );
  NAND U2124 ( .A(b[0]), .B(a[101]), .Z(n1798) );
  NAND U2125 ( .A(b[1]), .B(a[100]), .Z(n1797) );
  XNOR U2126 ( .A(n1798), .B(n1797), .Z(n1800) );
  XNOR U2127 ( .A(n1799), .B(n1800), .Z(n1804) );
  XOR U2128 ( .A(n1803), .B(sreg[355]), .Z(n1796) );
  XNOR U2129 ( .A(n1804), .B(n1796), .Z(c[355]) );
  NAND U2130 ( .A(n1798), .B(n1797), .Z(n1802) );
  NANDN U2131 ( .A(n1800), .B(n1799), .Z(n1801) );
  NAND U2132 ( .A(n1802), .B(n1801), .Z(n1809) );
  ANDN U2133 ( .B(a[102]), .A(n965), .Z(n1807) );
  ANDN U2134 ( .B(a[101]), .A(n966), .Z(n1806) );
  XOR U2135 ( .A(n1807), .B(n1806), .Z(n1808) );
  XNOR U2136 ( .A(n1809), .B(n1808), .Z(n1811) );
  XOR U2137 ( .A(sreg[356]), .B(n1810), .Z(n1805) );
  XNOR U2138 ( .A(n1811), .B(n1805), .Z(c[356]) );
  NAND U2139 ( .A(b[0]), .B(a[103]), .Z(n1814) );
  NAND U2140 ( .A(b[1]), .B(a[102]), .Z(n1813) );
  XNOR U2141 ( .A(n1814), .B(n1813), .Z(n1816) );
  XNOR U2142 ( .A(n1815), .B(n1816), .Z(n1820) );
  XOR U2143 ( .A(n1819), .B(sreg[357]), .Z(n1812) );
  XNOR U2144 ( .A(n1820), .B(n1812), .Z(c[357]) );
  NAND U2145 ( .A(n1814), .B(n1813), .Z(n1818) );
  NANDN U2146 ( .A(n1816), .B(n1815), .Z(n1817) );
  NAND U2147 ( .A(n1818), .B(n1817), .Z(n1825) );
  ANDN U2148 ( .B(a[104]), .A(n965), .Z(n1823) );
  ANDN U2149 ( .B(a[103]), .A(n966), .Z(n1822) );
  XOR U2150 ( .A(n1823), .B(n1822), .Z(n1824) );
  XNOR U2151 ( .A(n1825), .B(n1824), .Z(n1827) );
  XOR U2152 ( .A(sreg[358]), .B(n1826), .Z(n1821) );
  XNOR U2153 ( .A(n1827), .B(n1821), .Z(c[358]) );
  NAND U2154 ( .A(b[0]), .B(a[105]), .Z(n1830) );
  NAND U2155 ( .A(b[1]), .B(a[104]), .Z(n1829) );
  XNOR U2156 ( .A(n1830), .B(n1829), .Z(n1832) );
  XNOR U2157 ( .A(n1831), .B(n1832), .Z(n1836) );
  XOR U2158 ( .A(n1835), .B(sreg[359]), .Z(n1828) );
  XNOR U2159 ( .A(n1836), .B(n1828), .Z(c[359]) );
  NAND U2160 ( .A(n1830), .B(n1829), .Z(n1834) );
  NANDN U2161 ( .A(n1832), .B(n1831), .Z(n1833) );
  NAND U2162 ( .A(n1834), .B(n1833), .Z(n1841) );
  ANDN U2163 ( .B(a[106]), .A(n965), .Z(n1839) );
  ANDN U2164 ( .B(a[105]), .A(n966), .Z(n1838) );
  XOR U2165 ( .A(n1839), .B(n1838), .Z(n1840) );
  XNOR U2166 ( .A(n1841), .B(n1840), .Z(n1843) );
  XOR U2167 ( .A(sreg[360]), .B(n1842), .Z(n1837) );
  XNOR U2168 ( .A(n1843), .B(n1837), .Z(c[360]) );
  NAND U2169 ( .A(b[0]), .B(a[107]), .Z(n1846) );
  NAND U2170 ( .A(b[1]), .B(a[106]), .Z(n1845) );
  XNOR U2171 ( .A(n1846), .B(n1845), .Z(n1848) );
  XNOR U2172 ( .A(n1847), .B(n1848), .Z(n1852) );
  XOR U2173 ( .A(n1851), .B(sreg[361]), .Z(n1844) );
  XNOR U2174 ( .A(n1852), .B(n1844), .Z(c[361]) );
  NAND U2175 ( .A(n1846), .B(n1845), .Z(n1850) );
  NANDN U2176 ( .A(n1848), .B(n1847), .Z(n1849) );
  NAND U2177 ( .A(n1850), .B(n1849), .Z(n1857) );
  ANDN U2178 ( .B(a[108]), .A(n965), .Z(n1855) );
  ANDN U2179 ( .B(a[107]), .A(n966), .Z(n1854) );
  XOR U2180 ( .A(n1855), .B(n1854), .Z(n1856) );
  XNOR U2181 ( .A(n1857), .B(n1856), .Z(n1859) );
  XOR U2182 ( .A(sreg[362]), .B(n1858), .Z(n1853) );
  XNOR U2183 ( .A(n1859), .B(n1853), .Z(c[362]) );
  NAND U2184 ( .A(b[0]), .B(a[109]), .Z(n1862) );
  NAND U2185 ( .A(b[1]), .B(a[108]), .Z(n1861) );
  XNOR U2186 ( .A(n1862), .B(n1861), .Z(n1864) );
  XNOR U2187 ( .A(n1863), .B(n1864), .Z(n1868) );
  XOR U2188 ( .A(n1867), .B(sreg[363]), .Z(n1860) );
  XNOR U2189 ( .A(n1868), .B(n1860), .Z(c[363]) );
  NAND U2190 ( .A(n1862), .B(n1861), .Z(n1866) );
  NANDN U2191 ( .A(n1864), .B(n1863), .Z(n1865) );
  NAND U2192 ( .A(n1866), .B(n1865), .Z(n1873) );
  ANDN U2193 ( .B(a[110]), .A(n965), .Z(n1871) );
  ANDN U2194 ( .B(a[109]), .A(n966), .Z(n1870) );
  XOR U2195 ( .A(n1871), .B(n1870), .Z(n1872) );
  XNOR U2196 ( .A(n1873), .B(n1872), .Z(n1875) );
  XOR U2197 ( .A(sreg[364]), .B(n1874), .Z(n1869) );
  XNOR U2198 ( .A(n1875), .B(n1869), .Z(c[364]) );
  NAND U2199 ( .A(b[0]), .B(a[111]), .Z(n1878) );
  NAND U2200 ( .A(b[1]), .B(a[110]), .Z(n1877) );
  XNOR U2201 ( .A(n1878), .B(n1877), .Z(n1880) );
  XNOR U2202 ( .A(n1879), .B(n1880), .Z(n1884) );
  XOR U2203 ( .A(n1883), .B(sreg[365]), .Z(n1876) );
  XNOR U2204 ( .A(n1884), .B(n1876), .Z(c[365]) );
  NAND U2205 ( .A(n1878), .B(n1877), .Z(n1882) );
  NANDN U2206 ( .A(n1880), .B(n1879), .Z(n1881) );
  NAND U2207 ( .A(n1882), .B(n1881), .Z(n1888) );
  NAND U2208 ( .A(b[0]), .B(a[112]), .Z(n1887) );
  NAND U2209 ( .A(b[1]), .B(a[111]), .Z(n1886) );
  XNOR U2210 ( .A(n1887), .B(n1886), .Z(n1889) );
  XNOR U2211 ( .A(n1888), .B(n1889), .Z(n1893) );
  XOR U2212 ( .A(n1892), .B(sreg[366]), .Z(n1885) );
  XNOR U2213 ( .A(n1893), .B(n1885), .Z(c[366]) );
  NAND U2214 ( .A(n1887), .B(n1886), .Z(n1891) );
  NANDN U2215 ( .A(n1889), .B(n1888), .Z(n1890) );
  NAND U2216 ( .A(n1891), .B(n1890), .Z(n1897) );
  NAND U2217 ( .A(b[0]), .B(a[113]), .Z(n1896) );
  NAND U2218 ( .A(b[1]), .B(a[112]), .Z(n1895) );
  XNOR U2219 ( .A(n1896), .B(n1895), .Z(n1898) );
  XNOR U2220 ( .A(n1897), .B(n1898), .Z(n1902) );
  XOR U2221 ( .A(n1901), .B(sreg[367]), .Z(n1894) );
  XNOR U2222 ( .A(n1902), .B(n1894), .Z(c[367]) );
  NAND U2223 ( .A(n1896), .B(n1895), .Z(n1900) );
  NANDN U2224 ( .A(n1898), .B(n1897), .Z(n1899) );
  NAND U2225 ( .A(n1900), .B(n1899), .Z(n1907) );
  ANDN U2226 ( .B(a[114]), .A(n965), .Z(n1905) );
  ANDN U2227 ( .B(a[113]), .A(n966), .Z(n1904) );
  XOR U2228 ( .A(n1905), .B(n1904), .Z(n1906) );
  XNOR U2229 ( .A(n1907), .B(n1906), .Z(n1909) );
  XOR U2230 ( .A(sreg[368]), .B(n1908), .Z(n1903) );
  XNOR U2231 ( .A(n1909), .B(n1903), .Z(c[368]) );
  NAND U2232 ( .A(b[0]), .B(a[115]), .Z(n1912) );
  NAND U2233 ( .A(b[1]), .B(a[114]), .Z(n1911) );
  XNOR U2234 ( .A(n1912), .B(n1911), .Z(n1914) );
  XNOR U2235 ( .A(n1913), .B(n1914), .Z(n1918) );
  XOR U2236 ( .A(n1917), .B(sreg[369]), .Z(n1910) );
  XNOR U2237 ( .A(n1918), .B(n1910), .Z(c[369]) );
  NAND U2238 ( .A(n1912), .B(n1911), .Z(n1916) );
  NANDN U2239 ( .A(n1914), .B(n1913), .Z(n1915) );
  NAND U2240 ( .A(n1916), .B(n1915), .Z(n1923) );
  ANDN U2241 ( .B(a[116]), .A(n965), .Z(n1921) );
  ANDN U2242 ( .B(a[115]), .A(n966), .Z(n1920) );
  XOR U2243 ( .A(n1921), .B(n1920), .Z(n1922) );
  XNOR U2244 ( .A(n1923), .B(n1922), .Z(n1925) );
  XOR U2245 ( .A(sreg[370]), .B(n1924), .Z(n1919) );
  XNOR U2246 ( .A(n1925), .B(n1919), .Z(c[370]) );
  NAND U2247 ( .A(b[0]), .B(a[117]), .Z(n1928) );
  NAND U2248 ( .A(b[1]), .B(a[116]), .Z(n1927) );
  XNOR U2249 ( .A(n1928), .B(n1927), .Z(n1930) );
  XNOR U2250 ( .A(n1929), .B(n1930), .Z(n1934) );
  XOR U2251 ( .A(n1933), .B(sreg[371]), .Z(n1926) );
  XNOR U2252 ( .A(n1934), .B(n1926), .Z(c[371]) );
  NAND U2253 ( .A(n1928), .B(n1927), .Z(n1932) );
  NANDN U2254 ( .A(n1930), .B(n1929), .Z(n1931) );
  NAND U2255 ( .A(n1932), .B(n1931), .Z(n1939) );
  ANDN U2256 ( .B(a[118]), .A(n965), .Z(n1937) );
  ANDN U2257 ( .B(a[117]), .A(n966), .Z(n1936) );
  XOR U2258 ( .A(n1937), .B(n1936), .Z(n1938) );
  XNOR U2259 ( .A(n1939), .B(n1938), .Z(n1941) );
  XOR U2260 ( .A(sreg[372]), .B(n1940), .Z(n1935) );
  XNOR U2261 ( .A(n1941), .B(n1935), .Z(c[372]) );
  NAND U2262 ( .A(b[0]), .B(a[119]), .Z(n1944) );
  NAND U2263 ( .A(b[1]), .B(a[118]), .Z(n1943) );
  XNOR U2264 ( .A(n1944), .B(n1943), .Z(n1946) );
  XNOR U2265 ( .A(n1945), .B(n1946), .Z(n1950) );
  XOR U2266 ( .A(n1949), .B(sreg[373]), .Z(n1942) );
  XNOR U2267 ( .A(n1950), .B(n1942), .Z(c[373]) );
  NAND U2268 ( .A(n1944), .B(n1943), .Z(n1948) );
  NANDN U2269 ( .A(n1946), .B(n1945), .Z(n1947) );
  NAND U2270 ( .A(n1948), .B(n1947), .Z(n1955) );
  ANDN U2271 ( .B(a[120]), .A(n965), .Z(n1953) );
  ANDN U2272 ( .B(a[119]), .A(n966), .Z(n1952) );
  XOR U2273 ( .A(n1953), .B(n1952), .Z(n1954) );
  XNOR U2274 ( .A(n1955), .B(n1954), .Z(n1957) );
  XOR U2275 ( .A(sreg[374]), .B(n1956), .Z(n1951) );
  XNOR U2276 ( .A(n1957), .B(n1951), .Z(c[374]) );
  NAND U2277 ( .A(b[0]), .B(a[121]), .Z(n1960) );
  NAND U2278 ( .A(b[1]), .B(a[120]), .Z(n1959) );
  XNOR U2279 ( .A(n1960), .B(n1959), .Z(n1962) );
  XNOR U2280 ( .A(n1961), .B(n1962), .Z(n1966) );
  XOR U2281 ( .A(n1965), .B(sreg[375]), .Z(n1958) );
  XNOR U2282 ( .A(n1966), .B(n1958), .Z(c[375]) );
  NAND U2283 ( .A(n1960), .B(n1959), .Z(n1964) );
  NANDN U2284 ( .A(n1962), .B(n1961), .Z(n1963) );
  NAND U2285 ( .A(n1964), .B(n1963), .Z(n1970) );
  NAND U2286 ( .A(b[0]), .B(a[122]), .Z(n1969) );
  NAND U2287 ( .A(b[1]), .B(a[121]), .Z(n1968) );
  XNOR U2288 ( .A(n1969), .B(n1968), .Z(n1971) );
  XNOR U2289 ( .A(n1970), .B(n1971), .Z(n1975) );
  XOR U2290 ( .A(n1974), .B(sreg[376]), .Z(n1967) );
  XNOR U2291 ( .A(n1975), .B(n1967), .Z(c[376]) );
  NAND U2292 ( .A(n1969), .B(n1968), .Z(n1973) );
  NANDN U2293 ( .A(n1971), .B(n1970), .Z(n1972) );
  NAND U2294 ( .A(n1973), .B(n1972), .Z(n1979) );
  NAND U2295 ( .A(b[0]), .B(a[123]), .Z(n1978) );
  NAND U2296 ( .A(b[1]), .B(a[122]), .Z(n1977) );
  XNOR U2297 ( .A(n1978), .B(n1977), .Z(n1980) );
  XNOR U2298 ( .A(n1979), .B(n1980), .Z(n1984) );
  XOR U2299 ( .A(n1983), .B(sreg[377]), .Z(n1976) );
  XNOR U2300 ( .A(n1984), .B(n1976), .Z(c[377]) );
  NAND U2301 ( .A(n1978), .B(n1977), .Z(n1982) );
  NANDN U2302 ( .A(n1980), .B(n1979), .Z(n1981) );
  NAND U2303 ( .A(n1982), .B(n1981), .Z(n1989) );
  ANDN U2304 ( .B(a[124]), .A(n965), .Z(n1987) );
  ANDN U2305 ( .B(a[123]), .A(n966), .Z(n1986) );
  XOR U2306 ( .A(n1987), .B(n1986), .Z(n1988) );
  XNOR U2307 ( .A(n1989), .B(n1988), .Z(n1991) );
  XOR U2308 ( .A(sreg[378]), .B(n1990), .Z(n1985) );
  XNOR U2309 ( .A(n1991), .B(n1985), .Z(c[378]) );
  NAND U2310 ( .A(b[0]), .B(a[125]), .Z(n1994) );
  NAND U2311 ( .A(b[1]), .B(a[124]), .Z(n1993) );
  XNOR U2312 ( .A(n1994), .B(n1993), .Z(n1996) );
  XNOR U2313 ( .A(n1995), .B(n1996), .Z(n2000) );
  XOR U2314 ( .A(n1999), .B(sreg[379]), .Z(n1992) );
  XNOR U2315 ( .A(n2000), .B(n1992), .Z(c[379]) );
  NAND U2316 ( .A(n1994), .B(n1993), .Z(n1998) );
  NANDN U2317 ( .A(n1996), .B(n1995), .Z(n1997) );
  NAND U2318 ( .A(n1998), .B(n1997), .Z(n2005) );
  ANDN U2319 ( .B(a[126]), .A(n965), .Z(n2003) );
  ANDN U2320 ( .B(a[125]), .A(n966), .Z(n2002) );
  XOR U2321 ( .A(n2003), .B(n2002), .Z(n2004) );
  XNOR U2322 ( .A(n2005), .B(n2004), .Z(n2007) );
  XOR U2323 ( .A(sreg[380]), .B(n2006), .Z(n2001) );
  XNOR U2324 ( .A(n2007), .B(n2001), .Z(c[380]) );
  NAND U2325 ( .A(b[0]), .B(a[127]), .Z(n2010) );
  NAND U2326 ( .A(b[1]), .B(a[126]), .Z(n2009) );
  XNOR U2327 ( .A(n2010), .B(n2009), .Z(n2012) );
  XNOR U2328 ( .A(n2011), .B(n2012), .Z(n2016) );
  XOR U2329 ( .A(n2015), .B(sreg[381]), .Z(n2008) );
  XNOR U2330 ( .A(n2016), .B(n2008), .Z(c[381]) );
  NAND U2331 ( .A(n2010), .B(n2009), .Z(n2014) );
  NANDN U2332 ( .A(n2012), .B(n2011), .Z(n2013) );
  NAND U2333 ( .A(n2014), .B(n2013), .Z(n2021) );
  ANDN U2334 ( .B(a[128]), .A(n965), .Z(n2019) );
  ANDN U2335 ( .B(a[127]), .A(n966), .Z(n2018) );
  XOR U2336 ( .A(n2019), .B(n2018), .Z(n2020) );
  XNOR U2337 ( .A(n2021), .B(n2020), .Z(n2023) );
  XOR U2338 ( .A(sreg[382]), .B(n2022), .Z(n2017) );
  XNOR U2339 ( .A(n2023), .B(n2017), .Z(c[382]) );
  NAND U2340 ( .A(b[0]), .B(a[129]), .Z(n2026) );
  NAND U2341 ( .A(b[1]), .B(a[128]), .Z(n2025) );
  XNOR U2342 ( .A(n2026), .B(n2025), .Z(n2028) );
  XNOR U2343 ( .A(n2027), .B(n2028), .Z(n2032) );
  XOR U2344 ( .A(n2031), .B(sreg[383]), .Z(n2024) );
  XNOR U2345 ( .A(n2032), .B(n2024), .Z(c[383]) );
  NAND U2346 ( .A(n2026), .B(n2025), .Z(n2030) );
  NANDN U2347 ( .A(n2028), .B(n2027), .Z(n2029) );
  NAND U2348 ( .A(n2030), .B(n2029), .Z(n2036) );
  NAND U2349 ( .A(b[0]), .B(a[130]), .Z(n2035) );
  NAND U2350 ( .A(b[1]), .B(a[129]), .Z(n2034) );
  XNOR U2351 ( .A(n2035), .B(n2034), .Z(n2037) );
  XNOR U2352 ( .A(n2036), .B(n2037), .Z(n2041) );
  XOR U2353 ( .A(n2040), .B(sreg[384]), .Z(n2033) );
  XNOR U2354 ( .A(n2041), .B(n2033), .Z(c[384]) );
  NAND U2355 ( .A(n2035), .B(n2034), .Z(n2039) );
  NANDN U2356 ( .A(n2037), .B(n2036), .Z(n2038) );
  NAND U2357 ( .A(n2039), .B(n2038), .Z(n2045) );
  NAND U2358 ( .A(b[0]), .B(a[131]), .Z(n2044) );
  NAND U2359 ( .A(b[1]), .B(a[130]), .Z(n2043) );
  XNOR U2360 ( .A(n2044), .B(n2043), .Z(n2046) );
  XNOR U2361 ( .A(n2045), .B(n2046), .Z(n2050) );
  XOR U2362 ( .A(n2049), .B(sreg[385]), .Z(n2042) );
  XNOR U2363 ( .A(n2050), .B(n2042), .Z(c[385]) );
  NAND U2364 ( .A(n2044), .B(n2043), .Z(n2048) );
  NANDN U2365 ( .A(n2046), .B(n2045), .Z(n2047) );
  NAND U2366 ( .A(n2048), .B(n2047), .Z(n2055) );
  ANDN U2367 ( .B(a[132]), .A(n965), .Z(n2053) );
  ANDN U2368 ( .B(a[131]), .A(n966), .Z(n2052) );
  XOR U2369 ( .A(n2053), .B(n2052), .Z(n2054) );
  XNOR U2370 ( .A(n2055), .B(n2054), .Z(n2057) );
  XOR U2371 ( .A(sreg[386]), .B(n2056), .Z(n2051) );
  XNOR U2372 ( .A(n2057), .B(n2051), .Z(c[386]) );
  NAND U2373 ( .A(b[0]), .B(a[133]), .Z(n2060) );
  NAND U2374 ( .A(b[1]), .B(a[132]), .Z(n2059) );
  XNOR U2375 ( .A(n2060), .B(n2059), .Z(n2062) );
  XNOR U2376 ( .A(n2061), .B(n2062), .Z(n2066) );
  XOR U2377 ( .A(n2065), .B(sreg[387]), .Z(n2058) );
  XNOR U2378 ( .A(n2066), .B(n2058), .Z(c[387]) );
  NAND U2379 ( .A(n2060), .B(n2059), .Z(n2064) );
  NANDN U2380 ( .A(n2062), .B(n2061), .Z(n2063) );
  NAND U2381 ( .A(n2064), .B(n2063), .Z(n2070) );
  NAND U2382 ( .A(b[0]), .B(a[134]), .Z(n2069) );
  NAND U2383 ( .A(b[1]), .B(a[133]), .Z(n2068) );
  XNOR U2384 ( .A(n2069), .B(n2068), .Z(n2071) );
  XNOR U2385 ( .A(n2070), .B(n2071), .Z(n2075) );
  XOR U2386 ( .A(n2074), .B(sreg[388]), .Z(n2067) );
  XNOR U2387 ( .A(n2075), .B(n2067), .Z(c[388]) );
  NAND U2388 ( .A(n2069), .B(n2068), .Z(n2073) );
  NANDN U2389 ( .A(n2071), .B(n2070), .Z(n2072) );
  NAND U2390 ( .A(n2073), .B(n2072), .Z(n2079) );
  NAND U2391 ( .A(b[0]), .B(a[135]), .Z(n2078) );
  NAND U2392 ( .A(b[1]), .B(a[134]), .Z(n2077) );
  XNOR U2393 ( .A(n2078), .B(n2077), .Z(n2080) );
  XNOR U2394 ( .A(n2079), .B(n2080), .Z(n2084) );
  XOR U2395 ( .A(n2083), .B(sreg[389]), .Z(n2076) );
  XNOR U2396 ( .A(n2084), .B(n2076), .Z(c[389]) );
  NAND U2397 ( .A(n2078), .B(n2077), .Z(n2082) );
  NANDN U2398 ( .A(n2080), .B(n2079), .Z(n2081) );
  NAND U2399 ( .A(n2082), .B(n2081), .Z(n2089) );
  ANDN U2400 ( .B(a[136]), .A(n965), .Z(n2087) );
  ANDN U2401 ( .B(a[135]), .A(n966), .Z(n2086) );
  XOR U2402 ( .A(n2087), .B(n2086), .Z(n2088) );
  XNOR U2403 ( .A(n2089), .B(n2088), .Z(n2094) );
  XOR U2404 ( .A(sreg[390]), .B(n2093), .Z(n2085) );
  XNOR U2405 ( .A(n2094), .B(n2085), .Z(c[390]) );
  OR U2406 ( .A(n2087), .B(n2086), .Z(n2092) );
  IV U2407 ( .A(n2088), .Z(n2090) );
  NANDN U2408 ( .A(n2090), .B(n2089), .Z(n2091) );
  NAND U2409 ( .A(n2092), .B(n2091), .Z(n2099) );
  ANDN U2410 ( .B(a[137]), .A(n965), .Z(n2097) );
  ANDN U2411 ( .B(a[136]), .A(n966), .Z(n2096) );
  XOR U2412 ( .A(n2097), .B(n2096), .Z(n2098) );
  XNOR U2413 ( .A(n2099), .B(n2098), .Z(n2101) );
  XNOR U2414 ( .A(sreg[391]), .B(n2100), .Z(n2095) );
  XNOR U2415 ( .A(n2101), .B(n2095), .Z(c[391]) );
  ANDN U2416 ( .B(a[138]), .A(n965), .Z(n2104) );
  ANDN U2417 ( .B(a[137]), .A(n966), .Z(n2103) );
  XOR U2418 ( .A(n2104), .B(n2103), .Z(n2105) );
  XNOR U2419 ( .A(n2106), .B(n2105), .Z(n2108) );
  XNOR U2420 ( .A(sreg[392]), .B(n2107), .Z(n2102) );
  XNOR U2421 ( .A(n2108), .B(n2102), .Z(c[392]) );
  NAND U2422 ( .A(b[0]), .B(a[139]), .Z(n2111) );
  NAND U2423 ( .A(b[1]), .B(a[138]), .Z(n2110) );
  XNOR U2424 ( .A(n2111), .B(n2110), .Z(n2113) );
  XNOR U2425 ( .A(n2112), .B(n2113), .Z(n2117) );
  XOR U2426 ( .A(n2116), .B(sreg[393]), .Z(n2109) );
  XNOR U2427 ( .A(n2117), .B(n2109), .Z(c[393]) );
  NAND U2428 ( .A(n2111), .B(n2110), .Z(n2115) );
  NANDN U2429 ( .A(n2113), .B(n2112), .Z(n2114) );
  NAND U2430 ( .A(n2115), .B(n2114), .Z(n2122) );
  ANDN U2431 ( .B(a[140]), .A(n965), .Z(n2120) );
  ANDN U2432 ( .B(a[139]), .A(n966), .Z(n2119) );
  XOR U2433 ( .A(n2120), .B(n2119), .Z(n2121) );
  XNOR U2434 ( .A(n2122), .B(n2121), .Z(n2124) );
  XOR U2435 ( .A(sreg[394]), .B(n2123), .Z(n2118) );
  XNOR U2436 ( .A(n2124), .B(n2118), .Z(c[394]) );
  NAND U2437 ( .A(b[0]), .B(a[141]), .Z(n2127) );
  NAND U2438 ( .A(b[1]), .B(a[140]), .Z(n2126) );
  XNOR U2439 ( .A(n2127), .B(n2126), .Z(n2129) );
  XNOR U2440 ( .A(n2128), .B(n2129), .Z(n2133) );
  XOR U2441 ( .A(n2132), .B(sreg[395]), .Z(n2125) );
  XNOR U2442 ( .A(n2133), .B(n2125), .Z(c[395]) );
  NAND U2443 ( .A(n2127), .B(n2126), .Z(n2131) );
  NANDN U2444 ( .A(n2129), .B(n2128), .Z(n2130) );
  NAND U2445 ( .A(n2131), .B(n2130), .Z(n2138) );
  ANDN U2446 ( .B(a[142]), .A(n965), .Z(n2136) );
  ANDN U2447 ( .B(a[141]), .A(n966), .Z(n2135) );
  XOR U2448 ( .A(n2136), .B(n2135), .Z(n2137) );
  XNOR U2449 ( .A(n2138), .B(n2137), .Z(n2140) );
  XOR U2450 ( .A(sreg[396]), .B(n2139), .Z(n2134) );
  XNOR U2451 ( .A(n2140), .B(n2134), .Z(c[396]) );
  NAND U2452 ( .A(b[0]), .B(a[143]), .Z(n2143) );
  NAND U2453 ( .A(b[1]), .B(a[142]), .Z(n2142) );
  XNOR U2454 ( .A(n2143), .B(n2142), .Z(n2145) );
  XNOR U2455 ( .A(n2144), .B(n2145), .Z(n2149) );
  XOR U2456 ( .A(n2148), .B(sreg[397]), .Z(n2141) );
  XNOR U2457 ( .A(n2149), .B(n2141), .Z(c[397]) );
  NAND U2458 ( .A(n2143), .B(n2142), .Z(n2147) );
  NANDN U2459 ( .A(n2145), .B(n2144), .Z(n2146) );
  NAND U2460 ( .A(n2147), .B(n2146), .Z(n2154) );
  ANDN U2461 ( .B(a[144]), .A(n965), .Z(n2152) );
  ANDN U2462 ( .B(a[143]), .A(n966), .Z(n2151) );
  XOR U2463 ( .A(n2152), .B(n2151), .Z(n2153) );
  XNOR U2464 ( .A(n2154), .B(n2153), .Z(n2156) );
  XOR U2465 ( .A(sreg[398]), .B(n2155), .Z(n2150) );
  XNOR U2466 ( .A(n2156), .B(n2150), .Z(c[398]) );
  NAND U2467 ( .A(b[0]), .B(a[145]), .Z(n2159) );
  NAND U2468 ( .A(b[1]), .B(a[144]), .Z(n2158) );
  XNOR U2469 ( .A(n2159), .B(n2158), .Z(n2161) );
  XNOR U2470 ( .A(n2160), .B(n2161), .Z(n2165) );
  XOR U2471 ( .A(n2164), .B(sreg[399]), .Z(n2157) );
  XNOR U2472 ( .A(n2165), .B(n2157), .Z(c[399]) );
  NAND U2473 ( .A(n2159), .B(n2158), .Z(n2163) );
  NANDN U2474 ( .A(n2161), .B(n2160), .Z(n2162) );
  NAND U2475 ( .A(n2163), .B(n2162), .Z(n2169) );
  NAND U2476 ( .A(b[0]), .B(a[146]), .Z(n2168) );
  NAND U2477 ( .A(b[1]), .B(a[145]), .Z(n2167) );
  XNOR U2478 ( .A(n2168), .B(n2167), .Z(n2170) );
  XNOR U2479 ( .A(n2169), .B(n2170), .Z(n2174) );
  XOR U2480 ( .A(n2173), .B(sreg[400]), .Z(n2166) );
  XNOR U2481 ( .A(n2174), .B(n2166), .Z(c[400]) );
  NAND U2482 ( .A(n2168), .B(n2167), .Z(n2172) );
  NANDN U2483 ( .A(n2170), .B(n2169), .Z(n2171) );
  NAND U2484 ( .A(n2172), .B(n2171), .Z(n2178) );
  NAND U2485 ( .A(b[0]), .B(a[147]), .Z(n2177) );
  NAND U2486 ( .A(b[1]), .B(a[146]), .Z(n2176) );
  XNOR U2487 ( .A(n2177), .B(n2176), .Z(n2179) );
  XNOR U2488 ( .A(n2178), .B(n2179), .Z(n2183) );
  XOR U2489 ( .A(n2182), .B(sreg[401]), .Z(n2175) );
  XNOR U2490 ( .A(n2183), .B(n2175), .Z(c[401]) );
  NAND U2491 ( .A(n2177), .B(n2176), .Z(n2181) );
  NANDN U2492 ( .A(n2179), .B(n2178), .Z(n2180) );
  NAND U2493 ( .A(n2181), .B(n2180), .Z(n2187) );
  NAND U2494 ( .A(b[0]), .B(a[148]), .Z(n2186) );
  NAND U2495 ( .A(b[1]), .B(a[147]), .Z(n2185) );
  XNOR U2496 ( .A(n2186), .B(n2185), .Z(n2188) );
  XNOR U2497 ( .A(n2187), .B(n2188), .Z(n2192) );
  XOR U2498 ( .A(n2191), .B(sreg[402]), .Z(n2184) );
  XNOR U2499 ( .A(n2192), .B(n2184), .Z(c[402]) );
  NAND U2500 ( .A(n2186), .B(n2185), .Z(n2190) );
  NANDN U2501 ( .A(n2188), .B(n2187), .Z(n2189) );
  NAND U2502 ( .A(n2190), .B(n2189), .Z(n2196) );
  NAND U2503 ( .A(b[0]), .B(a[149]), .Z(n2195) );
  NAND U2504 ( .A(b[1]), .B(a[148]), .Z(n2194) );
  XNOR U2505 ( .A(n2195), .B(n2194), .Z(n2197) );
  XNOR U2506 ( .A(n2196), .B(n2197), .Z(n2201) );
  XOR U2507 ( .A(n2200), .B(sreg[403]), .Z(n2193) );
  XNOR U2508 ( .A(n2201), .B(n2193), .Z(c[403]) );
  NAND U2509 ( .A(n2195), .B(n2194), .Z(n2199) );
  NANDN U2510 ( .A(n2197), .B(n2196), .Z(n2198) );
  NAND U2511 ( .A(n2199), .B(n2198), .Z(n2206) );
  ANDN U2512 ( .B(a[150]), .A(n965), .Z(n2204) );
  ANDN U2513 ( .B(a[149]), .A(n966), .Z(n2203) );
  XOR U2514 ( .A(n2204), .B(n2203), .Z(n2205) );
  XNOR U2515 ( .A(n2206), .B(n2205), .Z(n2208) );
  XOR U2516 ( .A(sreg[404]), .B(n2207), .Z(n2202) );
  XNOR U2517 ( .A(n2208), .B(n2202), .Z(c[404]) );
  NAND U2518 ( .A(b[0]), .B(a[151]), .Z(n2211) );
  NAND U2519 ( .A(b[1]), .B(a[150]), .Z(n2210) );
  XNOR U2520 ( .A(n2211), .B(n2210), .Z(n2213) );
  XNOR U2521 ( .A(n2212), .B(n2213), .Z(n2217) );
  XOR U2522 ( .A(n2216), .B(sreg[405]), .Z(n2209) );
  XNOR U2523 ( .A(n2217), .B(n2209), .Z(c[405]) );
  NAND U2524 ( .A(n2211), .B(n2210), .Z(n2215) );
  NANDN U2525 ( .A(n2213), .B(n2212), .Z(n2214) );
  NAND U2526 ( .A(n2215), .B(n2214), .Z(n2222) );
  ANDN U2527 ( .B(a[152]), .A(n965), .Z(n2220) );
  ANDN U2528 ( .B(a[151]), .A(n966), .Z(n2219) );
  XOR U2529 ( .A(n2220), .B(n2219), .Z(n2221) );
  XNOR U2530 ( .A(n2222), .B(n2221), .Z(n2224) );
  XOR U2531 ( .A(sreg[406]), .B(n2223), .Z(n2218) );
  XNOR U2532 ( .A(n2224), .B(n2218), .Z(c[406]) );
  NAND U2533 ( .A(b[0]), .B(a[153]), .Z(n2227) );
  NAND U2534 ( .A(b[1]), .B(a[152]), .Z(n2226) );
  XNOR U2535 ( .A(n2227), .B(n2226), .Z(n2229) );
  XNOR U2536 ( .A(n2228), .B(n2229), .Z(n2233) );
  XOR U2537 ( .A(n2232), .B(sreg[407]), .Z(n2225) );
  XNOR U2538 ( .A(n2233), .B(n2225), .Z(c[407]) );
  NAND U2539 ( .A(n2227), .B(n2226), .Z(n2231) );
  NANDN U2540 ( .A(n2229), .B(n2228), .Z(n2230) );
  NAND U2541 ( .A(n2231), .B(n2230), .Z(n2238) );
  ANDN U2542 ( .B(a[154]), .A(n965), .Z(n2236) );
  ANDN U2543 ( .B(a[153]), .A(n966), .Z(n2235) );
  XOR U2544 ( .A(n2236), .B(n2235), .Z(n2237) );
  XNOR U2545 ( .A(n2238), .B(n2237), .Z(n2240) );
  XOR U2546 ( .A(sreg[408]), .B(n2239), .Z(n2234) );
  XNOR U2547 ( .A(n2240), .B(n2234), .Z(c[408]) );
  NAND U2548 ( .A(b[0]), .B(a[155]), .Z(n2243) );
  NAND U2549 ( .A(b[1]), .B(a[154]), .Z(n2242) );
  XNOR U2550 ( .A(n2243), .B(n2242), .Z(n2245) );
  XNOR U2551 ( .A(n2244), .B(n2245), .Z(n2249) );
  XOR U2552 ( .A(n2248), .B(sreg[409]), .Z(n2241) );
  XNOR U2553 ( .A(n2249), .B(n2241), .Z(c[409]) );
  NAND U2554 ( .A(n2243), .B(n2242), .Z(n2247) );
  NANDN U2555 ( .A(n2245), .B(n2244), .Z(n2246) );
  NAND U2556 ( .A(n2247), .B(n2246), .Z(n2254) );
  ANDN U2557 ( .B(a[156]), .A(n965), .Z(n2252) );
  ANDN U2558 ( .B(a[155]), .A(n966), .Z(n2251) );
  XOR U2559 ( .A(n2252), .B(n2251), .Z(n2253) );
  XNOR U2560 ( .A(n2254), .B(n2253), .Z(n2256) );
  XOR U2561 ( .A(sreg[410]), .B(n2255), .Z(n2250) );
  XNOR U2562 ( .A(n2256), .B(n2250), .Z(c[410]) );
  NAND U2563 ( .A(b[0]), .B(a[157]), .Z(n2259) );
  NAND U2564 ( .A(b[1]), .B(a[156]), .Z(n2258) );
  XNOR U2565 ( .A(n2259), .B(n2258), .Z(n2261) );
  XNOR U2566 ( .A(n2260), .B(n2261), .Z(n2265) );
  XOR U2567 ( .A(n2264), .B(sreg[411]), .Z(n2257) );
  XNOR U2568 ( .A(n2265), .B(n2257), .Z(c[411]) );
  NAND U2569 ( .A(n2259), .B(n2258), .Z(n2263) );
  NANDN U2570 ( .A(n2261), .B(n2260), .Z(n2262) );
  NAND U2571 ( .A(n2263), .B(n2262), .Z(n2269) );
  NAND U2572 ( .A(b[0]), .B(a[158]), .Z(n2268) );
  NAND U2573 ( .A(b[1]), .B(a[157]), .Z(n2267) );
  XNOR U2574 ( .A(n2268), .B(n2267), .Z(n2270) );
  XNOR U2575 ( .A(n2269), .B(n2270), .Z(n2274) );
  XOR U2576 ( .A(n2273), .B(sreg[412]), .Z(n2266) );
  XNOR U2577 ( .A(n2274), .B(n2266), .Z(c[412]) );
  NAND U2578 ( .A(n2268), .B(n2267), .Z(n2272) );
  NANDN U2579 ( .A(n2270), .B(n2269), .Z(n2271) );
  NAND U2580 ( .A(n2272), .B(n2271), .Z(n2278) );
  NAND U2581 ( .A(b[0]), .B(a[159]), .Z(n2277) );
  NAND U2582 ( .A(b[1]), .B(a[158]), .Z(n2276) );
  XNOR U2583 ( .A(n2277), .B(n2276), .Z(n2279) );
  XNOR U2584 ( .A(n2278), .B(n2279), .Z(n2283) );
  XOR U2585 ( .A(n2282), .B(sreg[413]), .Z(n2275) );
  XNOR U2586 ( .A(n2283), .B(n2275), .Z(c[413]) );
  NAND U2587 ( .A(n2277), .B(n2276), .Z(n2281) );
  NANDN U2588 ( .A(n2279), .B(n2278), .Z(n2280) );
  NAND U2589 ( .A(n2281), .B(n2280), .Z(n2288) );
  ANDN U2590 ( .B(a[160]), .A(n965), .Z(n2286) );
  ANDN U2591 ( .B(a[159]), .A(n966), .Z(n2285) );
  XOR U2592 ( .A(n2286), .B(n2285), .Z(n2287) );
  XNOR U2593 ( .A(n2288), .B(n2287), .Z(n2290) );
  XOR U2594 ( .A(sreg[414]), .B(n2289), .Z(n2284) );
  XNOR U2595 ( .A(n2290), .B(n2284), .Z(c[414]) );
  NAND U2596 ( .A(b[0]), .B(a[161]), .Z(n2293) );
  NAND U2597 ( .A(b[1]), .B(a[160]), .Z(n2292) );
  XNOR U2598 ( .A(n2293), .B(n2292), .Z(n2295) );
  XNOR U2599 ( .A(n2294), .B(n2295), .Z(n2299) );
  XOR U2600 ( .A(n2298), .B(sreg[415]), .Z(n2291) );
  XNOR U2601 ( .A(n2299), .B(n2291), .Z(c[415]) );
  NAND U2602 ( .A(n2293), .B(n2292), .Z(n2297) );
  NANDN U2603 ( .A(n2295), .B(n2294), .Z(n2296) );
  NAND U2604 ( .A(n2297), .B(n2296), .Z(n2304) );
  ANDN U2605 ( .B(a[162]), .A(n965), .Z(n2302) );
  ANDN U2606 ( .B(a[161]), .A(n966), .Z(n2301) );
  XOR U2607 ( .A(n2302), .B(n2301), .Z(n2303) );
  XNOR U2608 ( .A(n2304), .B(n2303), .Z(n2309) );
  XOR U2609 ( .A(sreg[416]), .B(n2308), .Z(n2300) );
  XNOR U2610 ( .A(n2309), .B(n2300), .Z(c[416]) );
  OR U2611 ( .A(n2302), .B(n2301), .Z(n2307) );
  IV U2612 ( .A(n2303), .Z(n2305) );
  NANDN U2613 ( .A(n2305), .B(n2304), .Z(n2306) );
  NAND U2614 ( .A(n2307), .B(n2306), .Z(n2314) );
  ANDN U2615 ( .B(a[163]), .A(n965), .Z(n2312) );
  ANDN U2616 ( .B(a[162]), .A(n966), .Z(n2311) );
  XOR U2617 ( .A(n2312), .B(n2311), .Z(n2313) );
  XNOR U2618 ( .A(n2314), .B(n2313), .Z(n2316) );
  XNOR U2619 ( .A(sreg[417]), .B(n2315), .Z(n2310) );
  XNOR U2620 ( .A(n2316), .B(n2310), .Z(c[417]) );
  ANDN U2621 ( .B(a[164]), .A(n965), .Z(n2319) );
  ANDN U2622 ( .B(a[163]), .A(n966), .Z(n2318) );
  XOR U2623 ( .A(n2319), .B(n2318), .Z(n2320) );
  XNOR U2624 ( .A(n2321), .B(n2320), .Z(n2323) );
  XNOR U2625 ( .A(sreg[418]), .B(n2322), .Z(n2317) );
  XNOR U2626 ( .A(n2323), .B(n2317), .Z(c[418]) );
  NAND U2627 ( .A(b[0]), .B(a[165]), .Z(n2326) );
  NAND U2628 ( .A(b[1]), .B(a[164]), .Z(n2325) );
  XNOR U2629 ( .A(n2326), .B(n2325), .Z(n2328) );
  XNOR U2630 ( .A(n2327), .B(n2328), .Z(n2332) );
  XOR U2631 ( .A(n2331), .B(sreg[419]), .Z(n2324) );
  XNOR U2632 ( .A(n2332), .B(n2324), .Z(c[419]) );
  NAND U2633 ( .A(n2326), .B(n2325), .Z(n2330) );
  NANDN U2634 ( .A(n2328), .B(n2327), .Z(n2329) );
  NAND U2635 ( .A(n2330), .B(n2329), .Z(n2337) );
  ANDN U2636 ( .B(a[166]), .A(n965), .Z(n2335) );
  ANDN U2637 ( .B(a[165]), .A(n966), .Z(n2334) );
  XOR U2638 ( .A(n2335), .B(n2334), .Z(n2336) );
  XNOR U2639 ( .A(n2337), .B(n2336), .Z(n2339) );
  XOR U2640 ( .A(sreg[420]), .B(n2338), .Z(n2333) );
  XNOR U2641 ( .A(n2339), .B(n2333), .Z(c[420]) );
  NAND U2642 ( .A(b[0]), .B(a[167]), .Z(n2342) );
  NAND U2643 ( .A(b[1]), .B(a[166]), .Z(n2341) );
  XNOR U2644 ( .A(n2342), .B(n2341), .Z(n2344) );
  XNOR U2645 ( .A(n2343), .B(n2344), .Z(n2348) );
  XOR U2646 ( .A(n2347), .B(sreg[421]), .Z(n2340) );
  XNOR U2647 ( .A(n2348), .B(n2340), .Z(c[421]) );
  NAND U2648 ( .A(n2342), .B(n2341), .Z(n2346) );
  NANDN U2649 ( .A(n2344), .B(n2343), .Z(n2345) );
  NAND U2650 ( .A(n2346), .B(n2345), .Z(n2353) );
  ANDN U2651 ( .B(a[168]), .A(n965), .Z(n2351) );
  ANDN U2652 ( .B(a[167]), .A(n966), .Z(n2350) );
  XOR U2653 ( .A(n2351), .B(n2350), .Z(n2352) );
  XNOR U2654 ( .A(n2353), .B(n2352), .Z(n2355) );
  XOR U2655 ( .A(sreg[422]), .B(n2354), .Z(n2349) );
  XNOR U2656 ( .A(n2355), .B(n2349), .Z(c[422]) );
  NAND U2657 ( .A(b[0]), .B(a[169]), .Z(n2358) );
  NAND U2658 ( .A(b[1]), .B(a[168]), .Z(n2357) );
  XNOR U2659 ( .A(n2358), .B(n2357), .Z(n2360) );
  XNOR U2660 ( .A(n2359), .B(n2360), .Z(n2364) );
  XOR U2661 ( .A(n2363), .B(sreg[423]), .Z(n2356) );
  XNOR U2662 ( .A(n2364), .B(n2356), .Z(c[423]) );
  NAND U2663 ( .A(n2358), .B(n2357), .Z(n2362) );
  NANDN U2664 ( .A(n2360), .B(n2359), .Z(n2361) );
  NAND U2665 ( .A(n2362), .B(n2361), .Z(n2369) );
  ANDN U2666 ( .B(a[170]), .A(n965), .Z(n2367) );
  ANDN U2667 ( .B(a[169]), .A(n966), .Z(n2366) );
  XOR U2668 ( .A(n2367), .B(n2366), .Z(n2368) );
  XNOR U2669 ( .A(n2369), .B(n2368), .Z(n2371) );
  XOR U2670 ( .A(sreg[424]), .B(n2370), .Z(n2365) );
  XNOR U2671 ( .A(n2371), .B(n2365), .Z(c[424]) );
  NAND U2672 ( .A(b[0]), .B(a[171]), .Z(n2374) );
  NAND U2673 ( .A(b[1]), .B(a[170]), .Z(n2373) );
  XNOR U2674 ( .A(n2374), .B(n2373), .Z(n2376) );
  XNOR U2675 ( .A(n2375), .B(n2376), .Z(n2380) );
  XOR U2676 ( .A(n2379), .B(sreg[425]), .Z(n2372) );
  XNOR U2677 ( .A(n2380), .B(n2372), .Z(c[425]) );
  NAND U2678 ( .A(n2374), .B(n2373), .Z(n2378) );
  NANDN U2679 ( .A(n2376), .B(n2375), .Z(n2377) );
  NAND U2680 ( .A(n2378), .B(n2377), .Z(n2385) );
  ANDN U2681 ( .B(a[172]), .A(n965), .Z(n2383) );
  ANDN U2682 ( .B(a[171]), .A(n966), .Z(n2382) );
  XOR U2683 ( .A(n2383), .B(n2382), .Z(n2384) );
  XNOR U2684 ( .A(n2385), .B(n2384), .Z(n2387) );
  XOR U2685 ( .A(sreg[426]), .B(n2386), .Z(n2381) );
  XNOR U2686 ( .A(n2387), .B(n2381), .Z(c[426]) );
  NAND U2687 ( .A(b[0]), .B(a[173]), .Z(n2390) );
  NAND U2688 ( .A(b[1]), .B(a[172]), .Z(n2389) );
  XNOR U2689 ( .A(n2390), .B(n2389), .Z(n2392) );
  XNOR U2690 ( .A(n2391), .B(n2392), .Z(n2396) );
  XOR U2691 ( .A(n2395), .B(sreg[427]), .Z(n2388) );
  XNOR U2692 ( .A(n2396), .B(n2388), .Z(c[427]) );
  NAND U2693 ( .A(n2390), .B(n2389), .Z(n2394) );
  NANDN U2694 ( .A(n2392), .B(n2391), .Z(n2393) );
  NAND U2695 ( .A(n2394), .B(n2393), .Z(n2401) );
  ANDN U2696 ( .B(a[174]), .A(n965), .Z(n2399) );
  ANDN U2697 ( .B(a[173]), .A(n966), .Z(n2398) );
  XOR U2698 ( .A(n2399), .B(n2398), .Z(n2400) );
  XNOR U2699 ( .A(n2401), .B(n2400), .Z(n2403) );
  XOR U2700 ( .A(sreg[428]), .B(n2402), .Z(n2397) );
  XNOR U2701 ( .A(n2403), .B(n2397), .Z(c[428]) );
  NAND U2702 ( .A(b[0]), .B(a[175]), .Z(n2406) );
  NAND U2703 ( .A(b[1]), .B(a[174]), .Z(n2405) );
  XNOR U2704 ( .A(n2406), .B(n2405), .Z(n2408) );
  XNOR U2705 ( .A(n2407), .B(n2408), .Z(n2412) );
  XOR U2706 ( .A(n2411), .B(sreg[429]), .Z(n2404) );
  XNOR U2707 ( .A(n2412), .B(n2404), .Z(c[429]) );
  NAND U2708 ( .A(n2406), .B(n2405), .Z(n2410) );
  NANDN U2709 ( .A(n2408), .B(n2407), .Z(n2409) );
  NAND U2710 ( .A(n2410), .B(n2409), .Z(n2417) );
  ANDN U2711 ( .B(a[176]), .A(n965), .Z(n2415) );
  ANDN U2712 ( .B(a[175]), .A(n966), .Z(n2414) );
  XOR U2713 ( .A(n2415), .B(n2414), .Z(n2416) );
  XNOR U2714 ( .A(n2417), .B(n2416), .Z(n2419) );
  XOR U2715 ( .A(sreg[430]), .B(n2418), .Z(n2413) );
  XNOR U2716 ( .A(n2419), .B(n2413), .Z(c[430]) );
  NAND U2717 ( .A(b[0]), .B(a[177]), .Z(n2422) );
  NAND U2718 ( .A(b[1]), .B(a[176]), .Z(n2421) );
  XNOR U2719 ( .A(n2422), .B(n2421), .Z(n2424) );
  XNOR U2720 ( .A(n2423), .B(n2424), .Z(n2428) );
  XOR U2721 ( .A(n2427), .B(sreg[431]), .Z(n2420) );
  XNOR U2722 ( .A(n2428), .B(n2420), .Z(c[431]) );
  NAND U2723 ( .A(n2422), .B(n2421), .Z(n2426) );
  NANDN U2724 ( .A(n2424), .B(n2423), .Z(n2425) );
  NAND U2725 ( .A(n2426), .B(n2425), .Z(n2432) );
  NAND U2726 ( .A(b[0]), .B(a[178]), .Z(n2431) );
  NAND U2727 ( .A(b[1]), .B(a[177]), .Z(n2430) );
  XNOR U2728 ( .A(n2431), .B(n2430), .Z(n2433) );
  XNOR U2729 ( .A(n2432), .B(n2433), .Z(n2437) );
  XOR U2730 ( .A(n2436), .B(sreg[432]), .Z(n2429) );
  XNOR U2731 ( .A(n2437), .B(n2429), .Z(c[432]) );
  NAND U2732 ( .A(n2431), .B(n2430), .Z(n2435) );
  NANDN U2733 ( .A(n2433), .B(n2432), .Z(n2434) );
  NAND U2734 ( .A(n2435), .B(n2434), .Z(n2441) );
  NAND U2735 ( .A(b[0]), .B(a[179]), .Z(n2440) );
  NAND U2736 ( .A(b[1]), .B(a[178]), .Z(n2439) );
  XNOR U2737 ( .A(n2440), .B(n2439), .Z(n2442) );
  XNOR U2738 ( .A(n2441), .B(n2442), .Z(n2446) );
  XOR U2739 ( .A(n2445), .B(sreg[433]), .Z(n2438) );
  XNOR U2740 ( .A(n2446), .B(n2438), .Z(c[433]) );
  NAND U2741 ( .A(n2440), .B(n2439), .Z(n2444) );
  NANDN U2742 ( .A(n2442), .B(n2441), .Z(n2443) );
  NAND U2743 ( .A(n2444), .B(n2443), .Z(n2451) );
  ANDN U2744 ( .B(a[180]), .A(n965), .Z(n2449) );
  ANDN U2745 ( .B(a[179]), .A(n966), .Z(n2448) );
  XOR U2746 ( .A(n2449), .B(n2448), .Z(n2450) );
  XNOR U2747 ( .A(n2451), .B(n2450), .Z(n2453) );
  XOR U2748 ( .A(sreg[434]), .B(n2452), .Z(n2447) );
  XNOR U2749 ( .A(n2453), .B(n2447), .Z(c[434]) );
  NAND U2750 ( .A(b[0]), .B(a[181]), .Z(n2456) );
  NAND U2751 ( .A(b[1]), .B(a[180]), .Z(n2455) );
  XNOR U2752 ( .A(n2456), .B(n2455), .Z(n2458) );
  XNOR U2753 ( .A(n2457), .B(n2458), .Z(n2462) );
  XOR U2754 ( .A(n2461), .B(sreg[435]), .Z(n2454) );
  XNOR U2755 ( .A(n2462), .B(n2454), .Z(c[435]) );
  NAND U2756 ( .A(n2456), .B(n2455), .Z(n2460) );
  NANDN U2757 ( .A(n2458), .B(n2457), .Z(n2459) );
  NAND U2758 ( .A(n2460), .B(n2459), .Z(n2467) );
  ANDN U2759 ( .B(a[182]), .A(n965), .Z(n2465) );
  ANDN U2760 ( .B(a[181]), .A(n966), .Z(n2464) );
  XOR U2761 ( .A(n2465), .B(n2464), .Z(n2466) );
  XNOR U2762 ( .A(n2467), .B(n2466), .Z(n2469) );
  XOR U2763 ( .A(sreg[436]), .B(n2468), .Z(n2463) );
  XNOR U2764 ( .A(n2469), .B(n2463), .Z(c[436]) );
  NAND U2765 ( .A(b[0]), .B(a[183]), .Z(n2472) );
  NAND U2766 ( .A(b[1]), .B(a[182]), .Z(n2471) );
  XNOR U2767 ( .A(n2472), .B(n2471), .Z(n2474) );
  XNOR U2768 ( .A(n2473), .B(n2474), .Z(n2478) );
  XOR U2769 ( .A(n2477), .B(sreg[437]), .Z(n2470) );
  XNOR U2770 ( .A(n2478), .B(n2470), .Z(c[437]) );
  NAND U2771 ( .A(n2472), .B(n2471), .Z(n2476) );
  NANDN U2772 ( .A(n2474), .B(n2473), .Z(n2475) );
  NAND U2773 ( .A(n2476), .B(n2475), .Z(n2483) );
  ANDN U2774 ( .B(a[184]), .A(n965), .Z(n2481) );
  ANDN U2775 ( .B(a[183]), .A(n966), .Z(n2480) );
  XOR U2776 ( .A(n2481), .B(n2480), .Z(n2482) );
  XNOR U2777 ( .A(n2483), .B(n2482), .Z(n2485) );
  XOR U2778 ( .A(sreg[438]), .B(n2484), .Z(n2479) );
  XNOR U2779 ( .A(n2485), .B(n2479), .Z(c[438]) );
  NAND U2780 ( .A(b[0]), .B(a[185]), .Z(n2488) );
  NAND U2781 ( .A(b[1]), .B(a[184]), .Z(n2487) );
  XNOR U2782 ( .A(n2488), .B(n2487), .Z(n2490) );
  XNOR U2783 ( .A(n2489), .B(n2490), .Z(n2494) );
  XOR U2784 ( .A(n2493), .B(sreg[439]), .Z(n2486) );
  XNOR U2785 ( .A(n2494), .B(n2486), .Z(c[439]) );
  NAND U2786 ( .A(n2488), .B(n2487), .Z(n2492) );
  NANDN U2787 ( .A(n2490), .B(n2489), .Z(n2491) );
  NAND U2788 ( .A(n2492), .B(n2491), .Z(n2499) );
  ANDN U2789 ( .B(a[186]), .A(n965), .Z(n2497) );
  ANDN U2790 ( .B(a[185]), .A(n966), .Z(n2496) );
  XOR U2791 ( .A(n2497), .B(n2496), .Z(n2498) );
  XNOR U2792 ( .A(n2499), .B(n2498), .Z(n2501) );
  XOR U2793 ( .A(sreg[440]), .B(n2500), .Z(n2495) );
  XNOR U2794 ( .A(n2501), .B(n2495), .Z(c[440]) );
  NAND U2795 ( .A(b[0]), .B(a[187]), .Z(n2504) );
  NAND U2796 ( .A(b[1]), .B(a[186]), .Z(n2503) );
  XNOR U2797 ( .A(n2504), .B(n2503), .Z(n2506) );
  XNOR U2798 ( .A(n2505), .B(n2506), .Z(n2510) );
  XOR U2799 ( .A(n2509), .B(sreg[441]), .Z(n2502) );
  XNOR U2800 ( .A(n2510), .B(n2502), .Z(c[441]) );
  NAND U2801 ( .A(n2504), .B(n2503), .Z(n2508) );
  NANDN U2802 ( .A(n2506), .B(n2505), .Z(n2507) );
  NAND U2803 ( .A(n2508), .B(n2507), .Z(n2515) );
  ANDN U2804 ( .B(a[188]), .A(n965), .Z(n2513) );
  ANDN U2805 ( .B(a[187]), .A(n966), .Z(n2512) );
  XOR U2806 ( .A(n2513), .B(n2512), .Z(n2514) );
  XNOR U2807 ( .A(n2515), .B(n2514), .Z(n2517) );
  XOR U2808 ( .A(sreg[442]), .B(n2516), .Z(n2511) );
  XNOR U2809 ( .A(n2517), .B(n2511), .Z(c[442]) );
  NAND U2810 ( .A(b[0]), .B(a[189]), .Z(n2520) );
  NAND U2811 ( .A(b[1]), .B(a[188]), .Z(n2519) );
  XNOR U2812 ( .A(n2520), .B(n2519), .Z(n2522) );
  XNOR U2813 ( .A(n2521), .B(n2522), .Z(n2526) );
  XOR U2814 ( .A(n2525), .B(sreg[443]), .Z(n2518) );
  XNOR U2815 ( .A(n2526), .B(n2518), .Z(c[443]) );
  NAND U2816 ( .A(n2520), .B(n2519), .Z(n2524) );
  NANDN U2817 ( .A(n2522), .B(n2521), .Z(n2523) );
  NAND U2818 ( .A(n2524), .B(n2523), .Z(n2531) );
  ANDN U2819 ( .B(a[190]), .A(n965), .Z(n2529) );
  ANDN U2820 ( .B(a[189]), .A(n966), .Z(n2528) );
  XOR U2821 ( .A(n2529), .B(n2528), .Z(n2530) );
  XNOR U2822 ( .A(n2531), .B(n2530), .Z(n2533) );
  XOR U2823 ( .A(sreg[444]), .B(n2532), .Z(n2527) );
  XNOR U2824 ( .A(n2533), .B(n2527), .Z(c[444]) );
  NAND U2825 ( .A(b[0]), .B(a[191]), .Z(n2536) );
  NAND U2826 ( .A(b[1]), .B(a[190]), .Z(n2535) );
  XNOR U2827 ( .A(n2536), .B(n2535), .Z(n2538) );
  XNOR U2828 ( .A(n2537), .B(n2538), .Z(n2542) );
  XOR U2829 ( .A(n2541), .B(sreg[445]), .Z(n2534) );
  XNOR U2830 ( .A(n2542), .B(n2534), .Z(c[445]) );
  NAND U2831 ( .A(n2536), .B(n2535), .Z(n2540) );
  NANDN U2832 ( .A(n2538), .B(n2537), .Z(n2539) );
  NAND U2833 ( .A(n2540), .B(n2539), .Z(n2547) );
  ANDN U2834 ( .B(a[192]), .A(n965), .Z(n2545) );
  ANDN U2835 ( .B(a[191]), .A(n966), .Z(n2544) );
  XOR U2836 ( .A(n2545), .B(n2544), .Z(n2546) );
  XNOR U2837 ( .A(n2547), .B(n2546), .Z(n2549) );
  XOR U2838 ( .A(sreg[446]), .B(n2548), .Z(n2543) );
  XNOR U2839 ( .A(n2549), .B(n2543), .Z(c[446]) );
  NAND U2840 ( .A(b[0]), .B(a[193]), .Z(n2552) );
  NAND U2841 ( .A(b[1]), .B(a[192]), .Z(n2551) );
  XNOR U2842 ( .A(n2552), .B(n2551), .Z(n2554) );
  XNOR U2843 ( .A(n2553), .B(n2554), .Z(n2558) );
  XOR U2844 ( .A(n2557), .B(sreg[447]), .Z(n2550) );
  XNOR U2845 ( .A(n2558), .B(n2550), .Z(c[447]) );
  NAND U2846 ( .A(n2552), .B(n2551), .Z(n2556) );
  NANDN U2847 ( .A(n2554), .B(n2553), .Z(n2555) );
  NAND U2848 ( .A(n2556), .B(n2555), .Z(n2563) );
  ANDN U2849 ( .B(a[194]), .A(n965), .Z(n2561) );
  ANDN U2850 ( .B(a[193]), .A(n966), .Z(n2560) );
  XOR U2851 ( .A(n2561), .B(n2560), .Z(n2562) );
  XNOR U2852 ( .A(n2563), .B(n2562), .Z(n2565) );
  XOR U2853 ( .A(sreg[448]), .B(n2564), .Z(n2559) );
  XNOR U2854 ( .A(n2565), .B(n2559), .Z(c[448]) );
  NAND U2855 ( .A(b[0]), .B(a[195]), .Z(n2568) );
  NAND U2856 ( .A(b[1]), .B(a[194]), .Z(n2567) );
  XNOR U2857 ( .A(n2568), .B(n2567), .Z(n2570) );
  XNOR U2858 ( .A(n2569), .B(n2570), .Z(n2574) );
  XOR U2859 ( .A(n2573), .B(sreg[449]), .Z(n2566) );
  XNOR U2860 ( .A(n2574), .B(n2566), .Z(c[449]) );
  NAND U2861 ( .A(n2568), .B(n2567), .Z(n2572) );
  NANDN U2862 ( .A(n2570), .B(n2569), .Z(n2571) );
  NAND U2863 ( .A(n2572), .B(n2571), .Z(n2579) );
  ANDN U2864 ( .B(a[196]), .A(n965), .Z(n2577) );
  ANDN U2865 ( .B(a[195]), .A(n966), .Z(n2576) );
  XOR U2866 ( .A(n2577), .B(n2576), .Z(n2578) );
  XNOR U2867 ( .A(n2579), .B(n2578), .Z(n2581) );
  XOR U2868 ( .A(sreg[450]), .B(n2580), .Z(n2575) );
  XNOR U2869 ( .A(n2581), .B(n2575), .Z(c[450]) );
  NAND U2870 ( .A(b[0]), .B(a[197]), .Z(n2584) );
  NAND U2871 ( .A(b[1]), .B(a[196]), .Z(n2583) );
  XNOR U2872 ( .A(n2584), .B(n2583), .Z(n2586) );
  XNOR U2873 ( .A(n2585), .B(n2586), .Z(n2590) );
  XOR U2874 ( .A(n2589), .B(sreg[451]), .Z(n2582) );
  XNOR U2875 ( .A(n2590), .B(n2582), .Z(c[451]) );
  NAND U2876 ( .A(n2584), .B(n2583), .Z(n2588) );
  NANDN U2877 ( .A(n2586), .B(n2585), .Z(n2587) );
  NAND U2878 ( .A(n2588), .B(n2587), .Z(n2595) );
  ANDN U2879 ( .B(a[198]), .A(n965), .Z(n2593) );
  ANDN U2880 ( .B(a[197]), .A(n966), .Z(n2592) );
  XOR U2881 ( .A(n2593), .B(n2592), .Z(n2594) );
  XNOR U2882 ( .A(n2595), .B(n2594), .Z(n2597) );
  XOR U2883 ( .A(sreg[452]), .B(n2596), .Z(n2591) );
  XNOR U2884 ( .A(n2597), .B(n2591), .Z(c[452]) );
  NAND U2885 ( .A(b[0]), .B(a[199]), .Z(n2600) );
  NAND U2886 ( .A(b[1]), .B(a[198]), .Z(n2599) );
  XNOR U2887 ( .A(n2600), .B(n2599), .Z(n2602) );
  XNOR U2888 ( .A(n2601), .B(n2602), .Z(n2606) );
  XOR U2889 ( .A(n2605), .B(sreg[453]), .Z(n2598) );
  XNOR U2890 ( .A(n2606), .B(n2598), .Z(c[453]) );
  NAND U2891 ( .A(n2600), .B(n2599), .Z(n2604) );
  NANDN U2892 ( .A(n2602), .B(n2601), .Z(n2603) );
  NAND U2893 ( .A(n2604), .B(n2603), .Z(n2611) );
  ANDN U2894 ( .B(a[200]), .A(n965), .Z(n2609) );
  ANDN U2895 ( .B(a[199]), .A(n966), .Z(n2608) );
  XOR U2896 ( .A(n2609), .B(n2608), .Z(n2610) );
  XNOR U2897 ( .A(n2611), .B(n2610), .Z(n2613) );
  XOR U2898 ( .A(sreg[454]), .B(n2612), .Z(n2607) );
  XNOR U2899 ( .A(n2613), .B(n2607), .Z(c[454]) );
  NAND U2900 ( .A(b[0]), .B(a[201]), .Z(n2616) );
  NAND U2901 ( .A(b[1]), .B(a[200]), .Z(n2615) );
  XNOR U2902 ( .A(n2616), .B(n2615), .Z(n2618) );
  XNOR U2903 ( .A(n2617), .B(n2618), .Z(n2622) );
  XOR U2904 ( .A(n2621), .B(sreg[455]), .Z(n2614) );
  XNOR U2905 ( .A(n2622), .B(n2614), .Z(c[455]) );
  NAND U2906 ( .A(n2616), .B(n2615), .Z(n2620) );
  NANDN U2907 ( .A(n2618), .B(n2617), .Z(n2619) );
  NAND U2908 ( .A(n2620), .B(n2619), .Z(n2627) );
  ANDN U2909 ( .B(a[202]), .A(n965), .Z(n2625) );
  ANDN U2910 ( .B(a[201]), .A(n966), .Z(n2624) );
  XOR U2911 ( .A(n2625), .B(n2624), .Z(n2626) );
  XNOR U2912 ( .A(n2627), .B(n2626), .Z(n2629) );
  XOR U2913 ( .A(sreg[456]), .B(n2628), .Z(n2623) );
  XNOR U2914 ( .A(n2629), .B(n2623), .Z(c[456]) );
  NAND U2915 ( .A(b[0]), .B(a[203]), .Z(n2632) );
  NAND U2916 ( .A(b[1]), .B(a[202]), .Z(n2631) );
  XNOR U2917 ( .A(n2632), .B(n2631), .Z(n2634) );
  XNOR U2918 ( .A(n2633), .B(n2634), .Z(n2638) );
  XOR U2919 ( .A(n2637), .B(sreg[457]), .Z(n2630) );
  XNOR U2920 ( .A(n2638), .B(n2630), .Z(c[457]) );
  NAND U2921 ( .A(n2632), .B(n2631), .Z(n2636) );
  NANDN U2922 ( .A(n2634), .B(n2633), .Z(n2635) );
  NAND U2923 ( .A(n2636), .B(n2635), .Z(n2643) );
  ANDN U2924 ( .B(a[204]), .A(n965), .Z(n2641) );
  ANDN U2925 ( .B(a[203]), .A(n966), .Z(n2640) );
  XOR U2926 ( .A(n2641), .B(n2640), .Z(n2642) );
  XNOR U2927 ( .A(n2643), .B(n2642), .Z(n2645) );
  XOR U2928 ( .A(sreg[458]), .B(n2644), .Z(n2639) );
  XNOR U2929 ( .A(n2645), .B(n2639), .Z(c[458]) );
  NAND U2930 ( .A(b[0]), .B(a[205]), .Z(n2648) );
  NAND U2931 ( .A(b[1]), .B(a[204]), .Z(n2647) );
  XNOR U2932 ( .A(n2648), .B(n2647), .Z(n2650) );
  XNOR U2933 ( .A(n2649), .B(n2650), .Z(n2654) );
  XOR U2934 ( .A(n2653), .B(sreg[459]), .Z(n2646) );
  XNOR U2935 ( .A(n2654), .B(n2646), .Z(c[459]) );
  NAND U2936 ( .A(n2648), .B(n2647), .Z(n2652) );
  NANDN U2937 ( .A(n2650), .B(n2649), .Z(n2651) );
  NAND U2938 ( .A(n2652), .B(n2651), .Z(n2659) );
  ANDN U2939 ( .B(a[206]), .A(n965), .Z(n2657) );
  ANDN U2940 ( .B(a[205]), .A(n966), .Z(n2656) );
  XOR U2941 ( .A(n2657), .B(n2656), .Z(n2658) );
  XNOR U2942 ( .A(n2659), .B(n2658), .Z(n2661) );
  XOR U2943 ( .A(sreg[460]), .B(n2660), .Z(n2655) );
  XNOR U2944 ( .A(n2661), .B(n2655), .Z(c[460]) );
  NAND U2945 ( .A(b[0]), .B(a[207]), .Z(n2664) );
  NAND U2946 ( .A(b[1]), .B(a[206]), .Z(n2663) );
  XNOR U2947 ( .A(n2664), .B(n2663), .Z(n2666) );
  XNOR U2948 ( .A(n2665), .B(n2666), .Z(n2670) );
  XOR U2949 ( .A(n2669), .B(sreg[461]), .Z(n2662) );
  XNOR U2950 ( .A(n2670), .B(n2662), .Z(c[461]) );
  NAND U2951 ( .A(n2664), .B(n2663), .Z(n2668) );
  NANDN U2952 ( .A(n2666), .B(n2665), .Z(n2667) );
  NAND U2953 ( .A(n2668), .B(n2667), .Z(n2674) );
  NAND U2954 ( .A(b[0]), .B(a[208]), .Z(n2673) );
  NAND U2955 ( .A(b[1]), .B(a[207]), .Z(n2672) );
  XNOR U2956 ( .A(n2673), .B(n2672), .Z(n2675) );
  XNOR U2957 ( .A(n2674), .B(n2675), .Z(n2679) );
  XOR U2958 ( .A(n2678), .B(sreg[462]), .Z(n2671) );
  XNOR U2959 ( .A(n2679), .B(n2671), .Z(c[462]) );
  NAND U2960 ( .A(n2673), .B(n2672), .Z(n2677) );
  NANDN U2961 ( .A(n2675), .B(n2674), .Z(n2676) );
  NAND U2962 ( .A(n2677), .B(n2676), .Z(n2683) );
  NAND U2963 ( .A(b[0]), .B(a[209]), .Z(n2682) );
  NAND U2964 ( .A(b[1]), .B(a[208]), .Z(n2681) );
  XNOR U2965 ( .A(n2682), .B(n2681), .Z(n2684) );
  XNOR U2966 ( .A(n2683), .B(n2684), .Z(n2688) );
  XOR U2967 ( .A(n2687), .B(sreg[463]), .Z(n2680) );
  XNOR U2968 ( .A(n2688), .B(n2680), .Z(c[463]) );
  NAND U2969 ( .A(n2682), .B(n2681), .Z(n2686) );
  NANDN U2970 ( .A(n2684), .B(n2683), .Z(n2685) );
  NAND U2971 ( .A(n2686), .B(n2685), .Z(n2693) );
  ANDN U2972 ( .B(a[210]), .A(n965), .Z(n2691) );
  ANDN U2973 ( .B(a[209]), .A(n966), .Z(n2690) );
  XOR U2974 ( .A(n2691), .B(n2690), .Z(n2692) );
  XNOR U2975 ( .A(n2693), .B(n2692), .Z(n2695) );
  XOR U2976 ( .A(sreg[464]), .B(n2694), .Z(n2689) );
  XNOR U2977 ( .A(n2695), .B(n2689), .Z(c[464]) );
  NAND U2978 ( .A(b[0]), .B(a[211]), .Z(n2698) );
  NAND U2979 ( .A(b[1]), .B(a[210]), .Z(n2697) );
  XNOR U2980 ( .A(n2698), .B(n2697), .Z(n2700) );
  XNOR U2981 ( .A(n2699), .B(n2700), .Z(n2704) );
  XOR U2982 ( .A(n2703), .B(sreg[465]), .Z(n2696) );
  XNOR U2983 ( .A(n2704), .B(n2696), .Z(c[465]) );
  NAND U2984 ( .A(n2698), .B(n2697), .Z(n2702) );
  NANDN U2985 ( .A(n2700), .B(n2699), .Z(n2701) );
  NAND U2986 ( .A(n2702), .B(n2701), .Z(n2709) );
  ANDN U2987 ( .B(a[212]), .A(n965), .Z(n2707) );
  ANDN U2988 ( .B(a[211]), .A(n966), .Z(n2706) );
  XOR U2989 ( .A(n2707), .B(n2706), .Z(n2708) );
  XNOR U2990 ( .A(n2709), .B(n2708), .Z(n2711) );
  XOR U2991 ( .A(sreg[466]), .B(n2710), .Z(n2705) );
  XNOR U2992 ( .A(n2711), .B(n2705), .Z(c[466]) );
  NAND U2993 ( .A(b[0]), .B(a[213]), .Z(n2714) );
  NAND U2994 ( .A(b[1]), .B(a[212]), .Z(n2713) );
  XNOR U2995 ( .A(n2714), .B(n2713), .Z(n2716) );
  XNOR U2996 ( .A(n2715), .B(n2716), .Z(n2720) );
  XOR U2997 ( .A(n2719), .B(sreg[467]), .Z(n2712) );
  XNOR U2998 ( .A(n2720), .B(n2712), .Z(c[467]) );
  NAND U2999 ( .A(n2714), .B(n2713), .Z(n2718) );
  NANDN U3000 ( .A(n2716), .B(n2715), .Z(n2717) );
  NAND U3001 ( .A(n2718), .B(n2717), .Z(n2725) );
  ANDN U3002 ( .B(a[214]), .A(n965), .Z(n2723) );
  ANDN U3003 ( .B(a[213]), .A(n966), .Z(n2722) );
  XOR U3004 ( .A(n2723), .B(n2722), .Z(n2724) );
  XNOR U3005 ( .A(n2725), .B(n2724), .Z(n2727) );
  XOR U3006 ( .A(sreg[468]), .B(n2726), .Z(n2721) );
  XNOR U3007 ( .A(n2727), .B(n2721), .Z(c[468]) );
  NAND U3008 ( .A(b[0]), .B(a[215]), .Z(n2730) );
  NAND U3009 ( .A(b[1]), .B(a[214]), .Z(n2729) );
  XNOR U3010 ( .A(n2730), .B(n2729), .Z(n2732) );
  XNOR U3011 ( .A(n2731), .B(n2732), .Z(n2736) );
  XOR U3012 ( .A(n2735), .B(sreg[469]), .Z(n2728) );
  XNOR U3013 ( .A(n2736), .B(n2728), .Z(c[469]) );
  NAND U3014 ( .A(n2730), .B(n2729), .Z(n2734) );
  NANDN U3015 ( .A(n2732), .B(n2731), .Z(n2733) );
  NAND U3016 ( .A(n2734), .B(n2733), .Z(n2741) );
  ANDN U3017 ( .B(a[216]), .A(n965), .Z(n2739) );
  ANDN U3018 ( .B(a[215]), .A(n966), .Z(n2738) );
  XOR U3019 ( .A(n2739), .B(n2738), .Z(n2740) );
  XNOR U3020 ( .A(n2741), .B(n2740), .Z(n2743) );
  XOR U3021 ( .A(sreg[470]), .B(n2742), .Z(n2737) );
  XNOR U3022 ( .A(n2743), .B(n2737), .Z(c[470]) );
  NAND U3023 ( .A(b[0]), .B(a[217]), .Z(n2746) );
  NAND U3024 ( .A(b[1]), .B(a[216]), .Z(n2745) );
  XNOR U3025 ( .A(n2746), .B(n2745), .Z(n2748) );
  XNOR U3026 ( .A(n2747), .B(n2748), .Z(n2752) );
  XOR U3027 ( .A(n2751), .B(sreg[471]), .Z(n2744) );
  XNOR U3028 ( .A(n2752), .B(n2744), .Z(c[471]) );
  NAND U3029 ( .A(n2746), .B(n2745), .Z(n2750) );
  NANDN U3030 ( .A(n2748), .B(n2747), .Z(n2749) );
  NAND U3031 ( .A(n2750), .B(n2749), .Z(n2757) );
  ANDN U3032 ( .B(a[218]), .A(n965), .Z(n2755) );
  ANDN U3033 ( .B(a[217]), .A(n966), .Z(n2754) );
  XOR U3034 ( .A(n2755), .B(n2754), .Z(n2756) );
  XNOR U3035 ( .A(n2757), .B(n2756), .Z(n2759) );
  XOR U3036 ( .A(sreg[472]), .B(n2758), .Z(n2753) );
  XNOR U3037 ( .A(n2759), .B(n2753), .Z(c[472]) );
  ANDN U3038 ( .B(a[219]), .A(n965), .Z(n2762) );
  ANDN U3039 ( .B(a[218]), .A(n966), .Z(n2761) );
  XOR U3040 ( .A(n2762), .B(n2761), .Z(n2763) );
  XNOR U3041 ( .A(n2764), .B(n2763), .Z(n2766) );
  XNOR U3042 ( .A(sreg[473]), .B(n2765), .Z(n2760) );
  XNOR U3043 ( .A(n2766), .B(n2760), .Z(c[473]) );
  NAND U3044 ( .A(b[0]), .B(a[220]), .Z(n2769) );
  NAND U3045 ( .A(b[1]), .B(a[219]), .Z(n2768) );
  XNOR U3046 ( .A(n2769), .B(n2768), .Z(n2771) );
  XNOR U3047 ( .A(n2770), .B(n2771), .Z(n2775) );
  XOR U3048 ( .A(n2774), .B(sreg[474]), .Z(n2767) );
  XNOR U3049 ( .A(n2775), .B(n2767), .Z(c[474]) );
  NAND U3050 ( .A(n2769), .B(n2768), .Z(n2773) );
  NANDN U3051 ( .A(n2771), .B(n2770), .Z(n2772) );
  NAND U3052 ( .A(n2773), .B(n2772), .Z(n2779) );
  NAND U3053 ( .A(b[0]), .B(a[221]), .Z(n2778) );
  NAND U3054 ( .A(b[1]), .B(a[220]), .Z(n2777) );
  XNOR U3055 ( .A(n2778), .B(n2777), .Z(n2780) );
  XNOR U3056 ( .A(n2779), .B(n2780), .Z(n2784) );
  XOR U3057 ( .A(n2783), .B(sreg[475]), .Z(n2776) );
  XNOR U3058 ( .A(n2784), .B(n2776), .Z(c[475]) );
  NAND U3059 ( .A(n2778), .B(n2777), .Z(n2782) );
  NANDN U3060 ( .A(n2780), .B(n2779), .Z(n2781) );
  NAND U3061 ( .A(n2782), .B(n2781), .Z(n2789) );
  ANDN U3062 ( .B(a[222]), .A(n965), .Z(n2787) );
  ANDN U3063 ( .B(a[221]), .A(n966), .Z(n2786) );
  XOR U3064 ( .A(n2787), .B(n2786), .Z(n2788) );
  XNOR U3065 ( .A(n2789), .B(n2788), .Z(n2791) );
  XOR U3066 ( .A(sreg[476]), .B(n2790), .Z(n2785) );
  XNOR U3067 ( .A(n2791), .B(n2785), .Z(c[476]) );
  NAND U3068 ( .A(b[0]), .B(a[223]), .Z(n2794) );
  NAND U3069 ( .A(b[1]), .B(a[222]), .Z(n2793) );
  XNOR U3070 ( .A(n2794), .B(n2793), .Z(n2796) );
  XNOR U3071 ( .A(n2795), .B(n2796), .Z(n2800) );
  XOR U3072 ( .A(n2799), .B(sreg[477]), .Z(n2792) );
  XNOR U3073 ( .A(n2800), .B(n2792), .Z(c[477]) );
  NAND U3074 ( .A(n2794), .B(n2793), .Z(n2798) );
  NANDN U3075 ( .A(n2796), .B(n2795), .Z(n2797) );
  NAND U3076 ( .A(n2798), .B(n2797), .Z(n2805) );
  ANDN U3077 ( .B(a[224]), .A(n965), .Z(n2803) );
  ANDN U3078 ( .B(a[223]), .A(n966), .Z(n2802) );
  XOR U3079 ( .A(n2803), .B(n2802), .Z(n2804) );
  XNOR U3080 ( .A(n2805), .B(n2804), .Z(n2807) );
  XOR U3081 ( .A(sreg[478]), .B(n2806), .Z(n2801) );
  XNOR U3082 ( .A(n2807), .B(n2801), .Z(c[478]) );
  NAND U3083 ( .A(b[0]), .B(a[225]), .Z(n2810) );
  NAND U3084 ( .A(b[1]), .B(a[224]), .Z(n2809) );
  XNOR U3085 ( .A(n2810), .B(n2809), .Z(n2812) );
  XNOR U3086 ( .A(n2811), .B(n2812), .Z(n2816) );
  XOR U3087 ( .A(n2815), .B(sreg[479]), .Z(n2808) );
  XNOR U3088 ( .A(n2816), .B(n2808), .Z(c[479]) );
  NAND U3089 ( .A(n2810), .B(n2809), .Z(n2814) );
  NANDN U3090 ( .A(n2812), .B(n2811), .Z(n2813) );
  NAND U3091 ( .A(n2814), .B(n2813), .Z(n2821) );
  ANDN U3092 ( .B(a[226]), .A(n965), .Z(n2819) );
  ANDN U3093 ( .B(a[225]), .A(n966), .Z(n2818) );
  XOR U3094 ( .A(n2819), .B(n2818), .Z(n2820) );
  XNOR U3095 ( .A(n2821), .B(n2820), .Z(n2823) );
  XOR U3096 ( .A(sreg[480]), .B(n2822), .Z(n2817) );
  XNOR U3097 ( .A(n2823), .B(n2817), .Z(c[480]) );
  NAND U3098 ( .A(b[0]), .B(a[227]), .Z(n2826) );
  NAND U3099 ( .A(b[1]), .B(a[226]), .Z(n2825) );
  XNOR U3100 ( .A(n2826), .B(n2825), .Z(n2828) );
  XNOR U3101 ( .A(n2827), .B(n2828), .Z(n2832) );
  XOR U3102 ( .A(n2831), .B(sreg[481]), .Z(n2824) );
  XNOR U3103 ( .A(n2832), .B(n2824), .Z(c[481]) );
  NAND U3104 ( .A(n2826), .B(n2825), .Z(n2830) );
  NANDN U3105 ( .A(n2828), .B(n2827), .Z(n2829) );
  NAND U3106 ( .A(n2830), .B(n2829), .Z(n2837) );
  ANDN U3107 ( .B(a[228]), .A(n965), .Z(n2835) );
  ANDN U3108 ( .B(a[227]), .A(n966), .Z(n2834) );
  XOR U3109 ( .A(n2835), .B(n2834), .Z(n2836) );
  XNOR U3110 ( .A(n2837), .B(n2836), .Z(n2839) );
  XOR U3111 ( .A(sreg[482]), .B(n2838), .Z(n2833) );
  XNOR U3112 ( .A(n2839), .B(n2833), .Z(c[482]) );
  NAND U3113 ( .A(b[0]), .B(a[229]), .Z(n2842) );
  NAND U3114 ( .A(b[1]), .B(a[228]), .Z(n2841) );
  XNOR U3115 ( .A(n2842), .B(n2841), .Z(n2844) );
  XNOR U3116 ( .A(n2843), .B(n2844), .Z(n2848) );
  XOR U3117 ( .A(n2847), .B(sreg[483]), .Z(n2840) );
  XNOR U3118 ( .A(n2848), .B(n2840), .Z(c[483]) );
  NAND U3119 ( .A(n2842), .B(n2841), .Z(n2846) );
  NANDN U3120 ( .A(n2844), .B(n2843), .Z(n2845) );
  NAND U3121 ( .A(n2846), .B(n2845), .Z(n2853) );
  ANDN U3122 ( .B(a[230]), .A(n965), .Z(n2851) );
  ANDN U3123 ( .B(a[229]), .A(n966), .Z(n2850) );
  XOR U3124 ( .A(n2851), .B(n2850), .Z(n2852) );
  XNOR U3125 ( .A(n2853), .B(n2852), .Z(n2855) );
  XOR U3126 ( .A(sreg[484]), .B(n2854), .Z(n2849) );
  XNOR U3127 ( .A(n2855), .B(n2849), .Z(c[484]) );
  NAND U3128 ( .A(b[0]), .B(a[231]), .Z(n2858) );
  NAND U3129 ( .A(b[1]), .B(a[230]), .Z(n2857) );
  XNOR U3130 ( .A(n2858), .B(n2857), .Z(n2860) );
  XNOR U3131 ( .A(n2859), .B(n2860), .Z(n2864) );
  XOR U3132 ( .A(n2863), .B(sreg[485]), .Z(n2856) );
  XNOR U3133 ( .A(n2864), .B(n2856), .Z(c[485]) );
  NAND U3134 ( .A(n2858), .B(n2857), .Z(n2862) );
  NANDN U3135 ( .A(n2860), .B(n2859), .Z(n2861) );
  NAND U3136 ( .A(n2862), .B(n2861), .Z(n2869) );
  ANDN U3137 ( .B(a[232]), .A(n965), .Z(n2867) );
  ANDN U3138 ( .B(a[231]), .A(n966), .Z(n2866) );
  XOR U3139 ( .A(n2867), .B(n2866), .Z(n2868) );
  XNOR U3140 ( .A(n2869), .B(n2868), .Z(n2871) );
  XOR U3141 ( .A(sreg[486]), .B(n2870), .Z(n2865) );
  XNOR U3142 ( .A(n2871), .B(n2865), .Z(c[486]) );
  NAND U3143 ( .A(b[0]), .B(a[233]), .Z(n2874) );
  NAND U3144 ( .A(b[1]), .B(a[232]), .Z(n2873) );
  XNOR U3145 ( .A(n2874), .B(n2873), .Z(n2876) );
  XNOR U3146 ( .A(n2875), .B(n2876), .Z(n2880) );
  XOR U3147 ( .A(n2879), .B(sreg[487]), .Z(n2872) );
  XNOR U3148 ( .A(n2880), .B(n2872), .Z(c[487]) );
  NAND U3149 ( .A(n2874), .B(n2873), .Z(n2878) );
  NANDN U3150 ( .A(n2876), .B(n2875), .Z(n2877) );
  NAND U3151 ( .A(n2878), .B(n2877), .Z(n2885) );
  ANDN U3152 ( .B(a[234]), .A(n965), .Z(n2883) );
  ANDN U3153 ( .B(a[233]), .A(n966), .Z(n2882) );
  XOR U3154 ( .A(n2883), .B(n2882), .Z(n2884) );
  XNOR U3155 ( .A(n2885), .B(n2884), .Z(n2887) );
  XOR U3156 ( .A(sreg[488]), .B(n2886), .Z(n2881) );
  XNOR U3157 ( .A(n2887), .B(n2881), .Z(c[488]) );
  NAND U3158 ( .A(b[0]), .B(a[235]), .Z(n2890) );
  NAND U3159 ( .A(b[1]), .B(a[234]), .Z(n2889) );
  XNOR U3160 ( .A(n2890), .B(n2889), .Z(n2892) );
  XNOR U3161 ( .A(n2891), .B(n2892), .Z(n2896) );
  XOR U3162 ( .A(n2895), .B(sreg[489]), .Z(n2888) );
  XNOR U3163 ( .A(n2896), .B(n2888), .Z(c[489]) );
  NAND U3164 ( .A(n2890), .B(n2889), .Z(n2894) );
  NANDN U3165 ( .A(n2892), .B(n2891), .Z(n2893) );
  NAND U3166 ( .A(n2894), .B(n2893), .Z(n2901) );
  ANDN U3167 ( .B(a[236]), .A(n965), .Z(n2899) );
  ANDN U3168 ( .B(a[235]), .A(n966), .Z(n2898) );
  XOR U3169 ( .A(n2899), .B(n2898), .Z(n2900) );
  XNOR U3170 ( .A(n2901), .B(n2900), .Z(n2903) );
  XOR U3171 ( .A(sreg[490]), .B(n2902), .Z(n2897) );
  XNOR U3172 ( .A(n2903), .B(n2897), .Z(c[490]) );
  NAND U3173 ( .A(b[0]), .B(a[237]), .Z(n2906) );
  NAND U3174 ( .A(b[1]), .B(a[236]), .Z(n2905) );
  XNOR U3175 ( .A(n2906), .B(n2905), .Z(n2908) );
  XNOR U3176 ( .A(n2907), .B(n2908), .Z(n2912) );
  XOR U3177 ( .A(n2911), .B(sreg[491]), .Z(n2904) );
  XNOR U3178 ( .A(n2912), .B(n2904), .Z(c[491]) );
  NAND U3179 ( .A(n2906), .B(n2905), .Z(n2910) );
  NANDN U3180 ( .A(n2908), .B(n2907), .Z(n2909) );
  NAND U3181 ( .A(n2910), .B(n2909), .Z(n2917) );
  ANDN U3182 ( .B(a[238]), .A(n965), .Z(n2915) );
  ANDN U3183 ( .B(a[237]), .A(n966), .Z(n2914) );
  XOR U3184 ( .A(n2915), .B(n2914), .Z(n2916) );
  XNOR U3185 ( .A(n2917), .B(n2916), .Z(n2922) );
  XOR U3186 ( .A(sreg[492]), .B(n2921), .Z(n2913) );
  XNOR U3187 ( .A(n2922), .B(n2913), .Z(c[492]) );
  OR U3188 ( .A(n2915), .B(n2914), .Z(n2920) );
  IV U3189 ( .A(n2916), .Z(n2918) );
  NANDN U3190 ( .A(n2918), .B(n2917), .Z(n2919) );
  NAND U3191 ( .A(n2920), .B(n2919), .Z(n2927) );
  ANDN U3192 ( .B(a[239]), .A(n965), .Z(n2925) );
  ANDN U3193 ( .B(a[238]), .A(n966), .Z(n2924) );
  XOR U3194 ( .A(n2925), .B(n2924), .Z(n2926) );
  XNOR U3195 ( .A(n2927), .B(n2926), .Z(n2929) );
  XNOR U3196 ( .A(sreg[493]), .B(n2928), .Z(n2923) );
  XNOR U3197 ( .A(n2929), .B(n2923), .Z(c[493]) );
  ANDN U3198 ( .B(a[240]), .A(n965), .Z(n2932) );
  ANDN U3199 ( .B(a[239]), .A(n966), .Z(n2931) );
  XOR U3200 ( .A(n2932), .B(n2931), .Z(n2933) );
  XNOR U3201 ( .A(n2934), .B(n2933), .Z(n2936) );
  XNOR U3202 ( .A(sreg[494]), .B(n2935), .Z(n2930) );
  XNOR U3203 ( .A(n2936), .B(n2930), .Z(c[494]) );
  NAND U3204 ( .A(b[0]), .B(a[241]), .Z(n2939) );
  NAND U3205 ( .A(b[1]), .B(a[240]), .Z(n2938) );
  XNOR U3206 ( .A(n2939), .B(n2938), .Z(n2941) );
  XNOR U3207 ( .A(n2940), .B(n2941), .Z(n2945) );
  XOR U3208 ( .A(n2944), .B(sreg[495]), .Z(n2937) );
  XNOR U3209 ( .A(n2945), .B(n2937), .Z(c[495]) );
  NAND U3210 ( .A(n2939), .B(n2938), .Z(n2943) );
  NANDN U3211 ( .A(n2941), .B(n2940), .Z(n2942) );
  NAND U3212 ( .A(n2943), .B(n2942), .Z(n2949) );
  NAND U3213 ( .A(b[0]), .B(a[242]), .Z(n2948) );
  NAND U3214 ( .A(b[1]), .B(a[241]), .Z(n2947) );
  XNOR U3215 ( .A(n2948), .B(n2947), .Z(n2950) );
  XNOR U3216 ( .A(n2949), .B(n2950), .Z(n2954) );
  XOR U3217 ( .A(n2953), .B(sreg[496]), .Z(n2946) );
  XNOR U3218 ( .A(n2954), .B(n2946), .Z(c[496]) );
  NAND U3219 ( .A(n2948), .B(n2947), .Z(n2952) );
  NANDN U3220 ( .A(n2950), .B(n2949), .Z(n2951) );
  NAND U3221 ( .A(n2952), .B(n2951), .Z(n2958) );
  NAND U3222 ( .A(b[0]), .B(a[243]), .Z(n2957) );
  NAND U3223 ( .A(b[1]), .B(a[242]), .Z(n2956) );
  XNOR U3224 ( .A(n2957), .B(n2956), .Z(n2959) );
  XNOR U3225 ( .A(n2958), .B(n2959), .Z(n2963) );
  XOR U3226 ( .A(n2962), .B(sreg[497]), .Z(n2955) );
  XNOR U3227 ( .A(n2963), .B(n2955), .Z(c[497]) );
  NAND U3228 ( .A(n2957), .B(n2956), .Z(n2961) );
  NANDN U3229 ( .A(n2959), .B(n2958), .Z(n2960) );
  NAND U3230 ( .A(n2961), .B(n2960), .Z(n2968) );
  ANDN U3231 ( .B(a[244]), .A(n965), .Z(n2966) );
  ANDN U3232 ( .B(a[243]), .A(n966), .Z(n2965) );
  XOR U3233 ( .A(n2966), .B(n2965), .Z(n2967) );
  XNOR U3234 ( .A(n2968), .B(n2967), .Z(n2970) );
  XOR U3235 ( .A(sreg[498]), .B(n2969), .Z(n2964) );
  XNOR U3236 ( .A(n2970), .B(n2964), .Z(c[498]) );
  NAND U3237 ( .A(b[0]), .B(a[245]), .Z(n2973) );
  NAND U3238 ( .A(b[1]), .B(a[244]), .Z(n2972) );
  XNOR U3239 ( .A(n2973), .B(n2972), .Z(n2975) );
  XNOR U3240 ( .A(n2974), .B(n2975), .Z(n2979) );
  XOR U3241 ( .A(n2978), .B(sreg[499]), .Z(n2971) );
  XNOR U3242 ( .A(n2979), .B(n2971), .Z(c[499]) );
  NAND U3243 ( .A(n2973), .B(n2972), .Z(n2977) );
  NANDN U3244 ( .A(n2975), .B(n2974), .Z(n2976) );
  NAND U3245 ( .A(n2977), .B(n2976), .Z(n2984) );
  ANDN U3246 ( .B(a[246]), .A(n965), .Z(n2982) );
  ANDN U3247 ( .B(a[245]), .A(n966), .Z(n2981) );
  XOR U3248 ( .A(n2982), .B(n2981), .Z(n2983) );
  XNOR U3249 ( .A(n2984), .B(n2983), .Z(n2986) );
  XOR U3250 ( .A(sreg[500]), .B(n2985), .Z(n2980) );
  XNOR U3251 ( .A(n2986), .B(n2980), .Z(c[500]) );
  NAND U3252 ( .A(b[0]), .B(a[247]), .Z(n2989) );
  NAND U3253 ( .A(b[1]), .B(a[246]), .Z(n2988) );
  XNOR U3254 ( .A(n2989), .B(n2988), .Z(n2991) );
  XNOR U3255 ( .A(n2990), .B(n2991), .Z(n2995) );
  XOR U3256 ( .A(n2994), .B(sreg[501]), .Z(n2987) );
  XNOR U3257 ( .A(n2995), .B(n2987), .Z(c[501]) );
  NAND U3258 ( .A(n2989), .B(n2988), .Z(n2993) );
  NANDN U3259 ( .A(n2991), .B(n2990), .Z(n2992) );
  NAND U3260 ( .A(n2993), .B(n2992), .Z(n3000) );
  ANDN U3261 ( .B(a[248]), .A(n965), .Z(n2998) );
  ANDN U3262 ( .B(a[247]), .A(n966), .Z(n2997) );
  XOR U3263 ( .A(n2998), .B(n2997), .Z(n2999) );
  XNOR U3264 ( .A(n3000), .B(n2999), .Z(n3002) );
  XOR U3265 ( .A(sreg[502]), .B(n3001), .Z(n2996) );
  XNOR U3266 ( .A(n3002), .B(n2996), .Z(c[502]) );
  NAND U3267 ( .A(b[0]), .B(a[249]), .Z(n3005) );
  NAND U3268 ( .A(b[1]), .B(a[248]), .Z(n3004) );
  XNOR U3269 ( .A(n3005), .B(n3004), .Z(n3007) );
  XNOR U3270 ( .A(n3006), .B(n3007), .Z(n3011) );
  XOR U3271 ( .A(n3010), .B(sreg[503]), .Z(n3003) );
  XNOR U3272 ( .A(n3011), .B(n3003), .Z(c[503]) );
  NAND U3273 ( .A(n3005), .B(n3004), .Z(n3009) );
  NANDN U3274 ( .A(n3007), .B(n3006), .Z(n3008) );
  NAND U3275 ( .A(n3009), .B(n3008), .Z(n3016) );
  ANDN U3276 ( .B(a[250]), .A(n965), .Z(n3014) );
  ANDN U3277 ( .B(a[249]), .A(n966), .Z(n3013) );
  XOR U3278 ( .A(n3014), .B(n3013), .Z(n3015) );
  XNOR U3279 ( .A(n3016), .B(n3015), .Z(n3021) );
  XOR U3280 ( .A(sreg[504]), .B(n3020), .Z(n3012) );
  XNOR U3281 ( .A(n3021), .B(n3012), .Z(c[504]) );
  OR U3282 ( .A(n3014), .B(n3013), .Z(n3019) );
  IV U3283 ( .A(n3015), .Z(n3017) );
  NANDN U3284 ( .A(n3017), .B(n3016), .Z(n3018) );
  NAND U3285 ( .A(n3019), .B(n3018), .Z(n3026) );
  ANDN U3286 ( .B(a[251]), .A(n965), .Z(n3024) );
  ANDN U3287 ( .B(a[250]), .A(n966), .Z(n3023) );
  XOR U3288 ( .A(n3024), .B(n3023), .Z(n3025) );
  XNOR U3289 ( .A(n3026), .B(n3025), .Z(n3028) );
  XNOR U3290 ( .A(sreg[505]), .B(n3027), .Z(n3022) );
  XNOR U3291 ( .A(n3028), .B(n3022), .Z(c[505]) );
  ANDN U3292 ( .B(a[252]), .A(n965), .Z(n3031) );
  ANDN U3293 ( .B(a[251]), .A(n966), .Z(n3030) );
  XOR U3294 ( .A(n3031), .B(n3030), .Z(n3032) );
  XNOR U3295 ( .A(n3033), .B(n3032), .Z(n3035) );
  XNOR U3296 ( .A(sreg[506]), .B(n3034), .Z(n3029) );
  XNOR U3297 ( .A(n3035), .B(n3029), .Z(c[506]) );
  NAND U3298 ( .A(b[0]), .B(a[253]), .Z(n3038) );
  NAND U3299 ( .A(b[1]), .B(a[252]), .Z(n3037) );
  XNOR U3300 ( .A(n3038), .B(n3037), .Z(n3040) );
  XNOR U3301 ( .A(n3039), .B(n3040), .Z(n3044) );
  XOR U3302 ( .A(n3043), .B(sreg[507]), .Z(n3036) );
  XNOR U3303 ( .A(n3044), .B(n3036), .Z(c[507]) );
  NAND U3304 ( .A(n3038), .B(n3037), .Z(n3042) );
  NANDN U3305 ( .A(n3040), .B(n3039), .Z(n3041) );
  NAND U3306 ( .A(n3042), .B(n3041), .Z(n3049) );
  ANDN U3307 ( .B(a[254]), .A(n965), .Z(n3046) );
  IV U3308 ( .A(n3046), .Z(n3057) );
  AND U3309 ( .A(a[253]), .B(b[1]), .Z(n3047) );
  XNOR U3310 ( .A(n3057), .B(n3047), .Z(n3048) );
  XOR U3311 ( .A(n3049), .B(n3048), .Z(n3055) );
  XOR U3312 ( .A(sreg[508]), .B(n3054), .Z(n3045) );
  XOR U3313 ( .A(n3055), .B(n3045), .Z(c[508]) );
  OR U3314 ( .A(n3047), .B(n3046), .Z(n3051) );
  NAND U3315 ( .A(n3049), .B(n3048), .Z(n3050) );
  NAND U3316 ( .A(n3051), .B(n3050), .Z(n3059) );
  ANDN U3317 ( .B(a[255]), .A(n965), .Z(n3053) );
  NANDN U3318 ( .A(n966), .B(a[254]), .Z(n3052) );
  XOR U3319 ( .A(n3053), .B(n3052), .Z(n3058) );
  XOR U3320 ( .A(n3059), .B(n3058), .Z(n3063) );
  XOR U3321 ( .A(n3062), .B(sreg[509]), .Z(n3056) );
  XOR U3322 ( .A(n3063), .B(n3056), .Z(c[509]) );
  AND U3323 ( .A(a[255]), .B(b[1]), .Z(n3066) );
  NANDN U3324 ( .A(n3057), .B(n3066), .Z(n3061) );
  OR U3325 ( .A(n3059), .B(n3058), .Z(n3060) );
  NAND U3326 ( .A(n3061), .B(n3060), .Z(n3068) );
  XOR U3327 ( .A(n3066), .B(n3067), .Z(n3064) );
  XOR U3328 ( .A(n3068), .B(n3064), .Z(c[510]) );
  XOR U3329 ( .A(n3068), .B(n3067), .Z(n3065) );
  NANDN U3330 ( .A(n3066), .B(n3065), .Z(n3070) );
  OR U3331 ( .A(n3068), .B(n3067), .Z(n3069) );
  AND U3332 ( .A(n3070), .B(n3069), .Z(c[511]) );
endmodule

