
module mult_N64_CC8 ( clk, rst, a, b, c );
  input [63:0] a;
  input [7:0] b;
  output [127:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695;
  wire   [127:0] sreg;

  DFF \sreg_reg[119]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(sreg[119]) );
  DFF \sreg_reg[118]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(sreg[118]) );
  DFF \sreg_reg[117]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(sreg[117]) );
  DFF \sreg_reg[116]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(sreg[116]) );
  DFF \sreg_reg[115]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(sreg[115]) );
  DFF \sreg_reg[114]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(sreg[114]) );
  DFF \sreg_reg[113]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(sreg[113]) );
  DFF \sreg_reg[112]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(sreg[112]) );
  DFF \sreg_reg[111]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(sreg[111]) );
  DFF \sreg_reg[110]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(sreg[110]) );
  DFF \sreg_reg[109]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(sreg[109]) );
  DFF \sreg_reg[108]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(sreg[108]) );
  DFF \sreg_reg[107]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(sreg[107]) );
  DFF \sreg_reg[106]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(sreg[106]) );
  DFF \sreg_reg[105]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(sreg[105]) );
  DFF \sreg_reg[104]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(sreg[104]) );
  DFF \sreg_reg[103]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(sreg[103]) );
  DFF \sreg_reg[102]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(sreg[102]) );
  DFF \sreg_reg[101]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(sreg[101]) );
  DFF \sreg_reg[100]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(sreg[100]) );
  DFF \sreg_reg[99]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(sreg[99]) );
  DFF \sreg_reg[98]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(sreg[98]) );
  DFF \sreg_reg[97]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(sreg[97]) );
  DFF \sreg_reg[96]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(sreg[96]) );
  DFF \sreg_reg[95]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(sreg[95]) );
  DFF \sreg_reg[94]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(sreg[94]) );
  DFF \sreg_reg[93]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(sreg[93]) );
  DFF \sreg_reg[92]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(sreg[92]) );
  DFF \sreg_reg[91]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(sreg[91]) );
  DFF \sreg_reg[90]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(sreg[90]) );
  DFF \sreg_reg[89]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(sreg[89]) );
  DFF \sreg_reg[88]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(sreg[88]) );
  DFF \sreg_reg[87]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(sreg[87]) );
  DFF \sreg_reg[86]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(sreg[86]) );
  DFF \sreg_reg[85]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(sreg[85]) );
  DFF \sreg_reg[84]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(sreg[84]) );
  DFF \sreg_reg[83]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(sreg[83]) );
  DFF \sreg_reg[82]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(sreg[82]) );
  DFF \sreg_reg[81]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(sreg[81]) );
  DFF \sreg_reg[80]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(sreg[80]) );
  DFF \sreg_reg[79]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(sreg[79]) );
  DFF \sreg_reg[78]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(sreg[78]) );
  DFF \sreg_reg[77]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(sreg[77]) );
  DFF \sreg_reg[76]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(sreg[76]) );
  DFF \sreg_reg[75]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(sreg[75]) );
  DFF \sreg_reg[74]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(sreg[74]) );
  DFF \sreg_reg[73]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(sreg[73]) );
  DFF \sreg_reg[72]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(sreg[72]) );
  DFF \sreg_reg[71]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(sreg[71]) );
  DFF \sreg_reg[70]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(sreg[70]) );
  DFF \sreg_reg[69]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(sreg[69]) );
  DFF \sreg_reg[68]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(sreg[68]) );
  DFF \sreg_reg[67]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(sreg[67]) );
  DFF \sreg_reg[66]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(sreg[66]) );
  DFF \sreg_reg[65]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(sreg[65]) );
  DFF \sreg_reg[64]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(sreg[64]) );
  DFF \sreg_reg[63]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(sreg[63]) );
  DFF \sreg_reg[62]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(sreg[62]) );
  DFF \sreg_reg[61]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(sreg[61]) );
  DFF \sreg_reg[60]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(sreg[60]) );
  DFF \sreg_reg[59]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(sreg[59]) );
  DFF \sreg_reg[58]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(sreg[58]) );
  DFF \sreg_reg[57]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(sreg[57]) );
  DFF \sreg_reg[56]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(sreg[56]) );
  DFF \sreg_reg[55]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[0]) );
  NANDN U11 ( .A(b[0]), .B(a[63]), .Z(n1) );
  NAND U12 ( .A(b[1]), .B(n1), .Z(n2519) );
  XNOR U13 ( .A(n2497), .B(n2496), .Z(n2498) );
  XNOR U14 ( .A(n2517), .B(n2516), .Z(n2518) );
  NAND U15 ( .A(n2588), .B(n2633), .Z(n2) );
  NAND U16 ( .A(n2634), .B(n35), .Z(n3) );
  NAND U17 ( .A(n2), .B(n3), .Z(n2616) );
  NAND U18 ( .A(n88), .B(n87), .Z(n4) );
  NANDN U19 ( .A(n90), .B(n89), .Z(n5) );
  AND U20 ( .A(n4), .B(n5), .Z(n111) );
  XNOR U21 ( .A(n2532), .B(n2531), .Z(n2533) );
  XNOR U22 ( .A(n2551), .B(b[1]), .Z(n2553) );
  XNOR U23 ( .A(n2452), .B(n2451), .Z(n2453) );
  XNOR U24 ( .A(n2474), .B(n2473), .Z(n2475) );
  XNOR U25 ( .A(n2580), .B(n2579), .Z(n2581) );
  XNOR U26 ( .A(n2611), .B(n2610), .Z(n2612) );
  XNOR U27 ( .A(n2654), .B(n2653), .Z(n2645) );
  XOR U28 ( .A(n72), .B(n70), .Z(n6) );
  NANDN U29 ( .A(n71), .B(n6), .Z(n7) );
  NAND U30 ( .A(n72), .B(n70), .Z(n8) );
  AND U31 ( .A(n7), .B(n8), .Z(n90) );
  XNOR U32 ( .A(n2491), .B(n2490), .Z(n2492) );
  XNOR U33 ( .A(n2454), .B(n2453), .Z(n2421) );
  XOR U34 ( .A(n2534), .B(n2533), .Z(n2510) );
  XNOR U35 ( .A(n2617), .B(n2616), .Z(n2619) );
  XOR U36 ( .A(n2476), .B(n2475), .Z(n2468) );
  XNOR U37 ( .A(n2548), .B(n2547), .Z(n2539) );
  XNOR U38 ( .A(n2582), .B(n2581), .Z(n2573) );
  XNOR U39 ( .A(n2613), .B(n2612), .Z(n2604) );
  XNOR U40 ( .A(n2646), .B(n2645), .Z(n2647) );
  NAND U41 ( .A(sreg[59]), .B(n83), .Z(n9) );
  XOR U42 ( .A(sreg[59]), .B(n83), .Z(n10) );
  NANDN U43 ( .A(n82), .B(n10), .Z(n11) );
  NAND U44 ( .A(n9), .B(n11), .Z(n85) );
  XOR U45 ( .A(n138), .B(sreg[62]), .Z(n12) );
  NANDN U46 ( .A(n139), .B(n12), .Z(n13) );
  NAND U47 ( .A(n138), .B(sreg[62]), .Z(n14) );
  AND U48 ( .A(n13), .B(n14), .Z(n206) );
  XOR U49 ( .A(n2693), .B(n2694), .Z(n2689) );
  XNOR U50 ( .A(n2434), .B(n2433), .Z(n2435) );
  XNOR U51 ( .A(n2428), .B(n2427), .Z(n2430) );
  XNOR U52 ( .A(n2519), .B(n2518), .Z(n2531) );
  XOR U53 ( .A(n2568), .B(n2567), .Z(n2552) );
  XNOR U54 ( .A(n2597), .B(n2596), .Z(n2598) );
  XNOR U55 ( .A(n2499), .B(n2498), .Z(n2473) );
  XNOR U56 ( .A(n2513), .B(n2512), .Z(n2504) );
  XNOR U57 ( .A(n2470), .B(n2469), .Z(n2462) );
  XNOR U58 ( .A(n2540), .B(n2539), .Z(n2541) );
  XNOR U59 ( .A(n2574), .B(n2573), .Z(n2575) );
  XNOR U60 ( .A(n2605), .B(n2604), .Z(n2606) );
  XNOR U61 ( .A(n2640), .B(n2639), .Z(n2641) );
  XOR U62 ( .A(sreg[60]), .B(n85), .Z(n15) );
  NANDN U63 ( .A(n86), .B(n15), .Z(n16) );
  NAND U64 ( .A(sreg[60]), .B(n85), .Z(n17) );
  AND U65 ( .A(n16), .B(n17), .Z(n134) );
  XOR U66 ( .A(n210), .B(sreg[64]), .Z(n18) );
  NANDN U67 ( .A(n211), .B(n18), .Z(n19) );
  NAND U68 ( .A(n210), .B(sreg[64]), .Z(n20) );
  AND U69 ( .A(n19), .B(n20), .Z(n286) );
  XNOR U70 ( .A(n2688), .B(n2689), .Z(n21) );
  XNOR U71 ( .A(n2687), .B(n21), .Z(n22) );
  NAND U72 ( .A(n2690), .B(n22), .Z(n23) );
  NANDN U73 ( .A(n2688), .B(n2689), .Z(n24) );
  NAND U74 ( .A(n2687), .B(n21), .Z(n25) );
  NAND U75 ( .A(n24), .B(n25), .Z(n26) );
  NAND U76 ( .A(n23), .B(n26), .Z(n27) );
  NAND U77 ( .A(n2692), .B(n2691), .Z(n28) );
  NANDN U78 ( .A(n2693), .B(n2694), .Z(n29) );
  AND U79 ( .A(n28), .B(n29), .Z(n30) );
  XNOR U80 ( .A(a[63]), .B(a[62]), .Z(n31) );
  XNOR U81 ( .A(n2695), .B(n31), .Z(n32) );
  AND U82 ( .A(n32), .B(b[7]), .Z(n33) );
  XNOR U83 ( .A(n27), .B(n30), .Z(n34) );
  XNOR U84 ( .A(n33), .B(n34), .Z(c[127]) );
  XOR U85 ( .A(b[4]), .B(b[3]), .Z(n35) );
  IV U86 ( .A(n2484), .Z(n36) );
  IV U87 ( .A(n35), .Z(n37) );
  AND U88 ( .A(b[0]), .B(a[0]), .Z(n39) );
  XOR U89 ( .A(n39), .B(sreg[56]), .Z(c[56]) );
  AND U90 ( .A(b[0]), .B(a[1]), .Z(n46) );
  NAND U91 ( .A(a[0]), .B(b[1]), .Z(n38) );
  XOR U92 ( .A(n46), .B(n38), .Z(n40) );
  XNOR U93 ( .A(sreg[57]), .B(n40), .Z(n42) );
  AND U94 ( .A(n39), .B(sreg[56]), .Z(n41) );
  XOR U95 ( .A(n42), .B(n41), .Z(c[57]) );
  NANDN U96 ( .A(n40), .B(sreg[57]), .Z(n44) );
  NAND U97 ( .A(n42), .B(n41), .Z(n43) );
  AND U98 ( .A(n44), .B(n43), .Z(n52) );
  XNOR U99 ( .A(n52), .B(sreg[58]), .Z(n54) );
  NAND U100 ( .A(a[0]), .B(b[2]), .Z(n45) );
  XNOR U101 ( .A(b[1]), .B(n45), .Z(n48) );
  NANDN U102 ( .A(a[0]), .B(n46), .Z(n47) );
  NAND U103 ( .A(n48), .B(n47), .Z(n58) );
  NAND U104 ( .A(b[0]), .B(a[2]), .Z(n49) );
  XNOR U105 ( .A(b[1]), .B(n49), .Z(n51) );
  NANDN U106 ( .A(b[0]), .B(a[1]), .Z(n50) );
  NAND U107 ( .A(n51), .B(n50), .Z(n57) );
  XOR U108 ( .A(n58), .B(n57), .Z(n53) );
  XOR U109 ( .A(n54), .B(n53), .Z(c[58]) );
  NANDN U110 ( .A(n52), .B(sreg[58]), .Z(n56) );
  NAND U111 ( .A(n54), .B(n53), .Z(n55) );
  NAND U112 ( .A(n56), .B(n55), .Z(n83) );
  NOR U113 ( .A(n58), .B(n57), .Z(n72) );
  NAND U114 ( .A(b[0]), .B(a[3]), .Z(n59) );
  XNOR U115 ( .A(b[1]), .B(n59), .Z(n61) );
  NANDN U116 ( .A(b[0]), .B(a[2]), .Z(n60) );
  NAND U117 ( .A(n61), .B(n60), .Z(n80) );
  XOR U118 ( .A(b[3]), .B(b[2]), .Z(n73) );
  XOR U119 ( .A(b[3]), .B(a[0]), .Z(n62) );
  NAND U120 ( .A(n73), .B(n62), .Z(n63) );
  XNOR U121 ( .A(b[2]), .B(b[1]), .Z(n2484) );
  OR U122 ( .A(n63), .B(n36), .Z(n65) );
  XOR U123 ( .A(b[3]), .B(a[1]), .Z(n74) );
  NAND U124 ( .A(n36), .B(n74), .Z(n64) );
  AND U125 ( .A(n65), .B(n64), .Z(n81) );
  XNOR U126 ( .A(n80), .B(n81), .Z(n71) );
  NANDN U127 ( .A(n2484), .B(a[0]), .Z(n67) );
  NANDN U128 ( .A(b[2]), .B(b[3]), .Z(n66) );
  NANDN U129 ( .A(n2484), .B(b[3]), .Z(n2559) );
  NAND U130 ( .A(n66), .B(n2559), .Z(n2623) );
  IV U131 ( .A(n2623), .Z(n2589) );
  ANDN U132 ( .B(n67), .A(n2589), .Z(n70) );
  XOR U133 ( .A(n71), .B(n70), .Z(n68) );
  XOR U134 ( .A(n72), .B(n68), .Z(n82) );
  XOR U135 ( .A(sreg[59]), .B(n82), .Z(n69) );
  XNOR U136 ( .A(n83), .B(n69), .Z(c[59]) );
  ANDN U137 ( .B(n73), .A(n36), .Z(n2556) );
  IV U138 ( .A(n2556), .Z(n2483) );
  NANDN U139 ( .A(n2483), .B(n74), .Z(n76) );
  XOR U140 ( .A(b[3]), .B(a[2]), .Z(n91) );
  NANDN U141 ( .A(n2484), .B(n91), .Z(n75) );
  AND U142 ( .A(n76), .B(n75), .Z(n105) );
  ANDN U143 ( .B(a[0]), .A(n37), .Z(n102) );
  NAND U144 ( .A(b[0]), .B(a[4]), .Z(n77) );
  XNOR U145 ( .A(b[1]), .B(n77), .Z(n79) );
  NANDN U146 ( .A(b[0]), .B(a[3]), .Z(n78) );
  NAND U147 ( .A(n79), .B(n78), .Z(n103) );
  XNOR U148 ( .A(n102), .B(n103), .Z(n104) );
  XNOR U149 ( .A(n105), .B(n104), .Z(n88) );
  NOR U150 ( .A(n81), .B(n80), .Z(n87) );
  XOR U151 ( .A(n88), .B(n87), .Z(n89) );
  XOR U152 ( .A(n90), .B(n89), .Z(n86) );
  XOR U153 ( .A(n85), .B(sreg[60]), .Z(n84) );
  XNOR U154 ( .A(n86), .B(n84), .Z(c[60]) );
  NANDN U155 ( .A(n2483), .B(n91), .Z(n93) );
  XOR U156 ( .A(b[3]), .B(a[3]), .Z(n114) );
  NANDN U157 ( .A(n2484), .B(n114), .Z(n92) );
  AND U158 ( .A(n93), .B(n92), .Z(n127) );
  NANDN U159 ( .A(b[4]), .B(b[5]), .Z(n94) );
  NANDN U160 ( .A(n37), .B(b[5]), .Z(n2636) );
  NAND U161 ( .A(n94), .B(n2636), .Z(n2661) );
  ANDN U162 ( .B(n2661), .A(n102), .Z(n126) );
  XNOR U163 ( .A(n127), .B(n126), .Z(n129) );
  NAND U164 ( .A(b[0]), .B(a[5]), .Z(n95) );
  XNOR U165 ( .A(b[1]), .B(n95), .Z(n97) );
  NANDN U166 ( .A(b[0]), .B(a[4]), .Z(n96) );
  NAND U167 ( .A(n97), .B(n96), .Z(n124) );
  XOR U168 ( .A(b[5]), .B(b[4]), .Z(n120) );
  XOR U169 ( .A(b[5]), .B(a[0]), .Z(n98) );
  NAND U170 ( .A(n120), .B(n98), .Z(n99) );
  OR U171 ( .A(n99), .B(n35), .Z(n101) );
  XOR U172 ( .A(b[5]), .B(a[1]), .Z(n121) );
  NAND U173 ( .A(n35), .B(n121), .Z(n100) );
  NAND U174 ( .A(n101), .B(n100), .Z(n125) );
  XNOR U175 ( .A(n124), .B(n125), .Z(n128) );
  XOR U176 ( .A(n129), .B(n128), .Z(n109) );
  NANDN U177 ( .A(n103), .B(n102), .Z(n107) );
  NANDN U178 ( .A(n105), .B(n104), .Z(n106) );
  AND U179 ( .A(n107), .B(n106), .Z(n108) );
  XNOR U180 ( .A(n109), .B(n108), .Z(n110) );
  XOR U181 ( .A(n111), .B(n110), .Z(n132) );
  XNOR U182 ( .A(n132), .B(sreg[61]), .Z(n133) );
  XNOR U183 ( .A(n134), .B(n133), .Z(c[61]) );
  NANDN U184 ( .A(n109), .B(n108), .Z(n113) );
  NAND U185 ( .A(n111), .B(n110), .Z(n112) );
  AND U186 ( .A(n113), .B(n112), .Z(n143) );
  NANDN U187 ( .A(n2483), .B(n114), .Z(n116) );
  XOR U188 ( .A(b[3]), .B(a[4]), .Z(n157) );
  NANDN U189 ( .A(n2484), .B(n157), .Z(n115) );
  AND U190 ( .A(n116), .B(n115), .Z(n163) );
  XOR U191 ( .A(b[5]), .B(b[6]), .Z(n2666) );
  IV U192 ( .A(n2666), .Z(n2630) );
  ANDN U193 ( .B(a[0]), .A(n2630), .Z(n160) );
  NAND U194 ( .A(b[0]), .B(a[6]), .Z(n117) );
  XNOR U195 ( .A(b[1]), .B(n117), .Z(n119) );
  NANDN U196 ( .A(b[0]), .B(a[5]), .Z(n118) );
  NAND U197 ( .A(n119), .B(n118), .Z(n161) );
  XNOR U198 ( .A(n160), .B(n161), .Z(n162) );
  XNOR U199 ( .A(n163), .B(n162), .Z(n169) );
  ANDN U200 ( .B(n120), .A(n35), .Z(n2633) );
  NAND U201 ( .A(n2633), .B(n121), .Z(n123) );
  XOR U202 ( .A(b[5]), .B(a[2]), .Z(n146) );
  NANDN U203 ( .A(n37), .B(n146), .Z(n122) );
  AND U204 ( .A(n123), .B(n122), .Z(n167) );
  ANDN U205 ( .B(n125), .A(n124), .Z(n166) );
  XNOR U206 ( .A(n167), .B(n166), .Z(n168) );
  XOR U207 ( .A(n169), .B(n168), .Z(n141) );
  NANDN U208 ( .A(n127), .B(n126), .Z(n131) );
  NAND U209 ( .A(n129), .B(n128), .Z(n130) );
  AND U210 ( .A(n131), .B(n130), .Z(n140) );
  XNOR U211 ( .A(n141), .B(n140), .Z(n142) );
  XNOR U212 ( .A(n143), .B(n142), .Z(n139) );
  NANDN U213 ( .A(n132), .B(sreg[61]), .Z(n136) );
  NANDN U214 ( .A(n134), .B(n133), .Z(n135) );
  NAND U215 ( .A(n136), .B(n135), .Z(n138) );
  XOR U216 ( .A(n138), .B(sreg[62]), .Z(n137) );
  XNOR U217 ( .A(n139), .B(n137), .Z(c[62]) );
  NANDN U218 ( .A(n141), .B(n140), .Z(n145) );
  NANDN U219 ( .A(n143), .B(n142), .Z(n144) );
  AND U220 ( .A(n145), .B(n144), .Z(n174) );
  NAND U221 ( .A(n2633), .B(n146), .Z(n148) );
  XOR U222 ( .A(b[5]), .B(a[3]), .Z(n201) );
  NANDN U223 ( .A(n37), .B(n201), .Z(n147) );
  AND U224 ( .A(n148), .B(n147), .Z(n197) );
  XOR U225 ( .A(b[6]), .B(b[7]), .Z(n149) );
  ANDN U226 ( .B(n149), .A(n2666), .Z(n2667) );
  IV U227 ( .A(n2667), .Z(n2629) );
  XOR U228 ( .A(a[0]), .B(b[7]), .Z(n150) );
  NANDN U229 ( .A(n2629), .B(n150), .Z(n152) );
  XOR U230 ( .A(b[7]), .B(a[1]), .Z(n190) );
  ANDN U231 ( .B(n190), .A(n2630), .Z(n151) );
  ANDN U232 ( .B(n152), .A(n151), .Z(n196) );
  XOR U233 ( .A(n197), .B(n196), .Z(n187) );
  NAND U234 ( .A(b[5]), .B(b[6]), .Z(n2695) );
  AND U235 ( .A(b[7]), .B(n2695), .Z(n153) );
  ANDN U236 ( .B(n153), .A(n160), .Z(n185) );
  NAND U237 ( .A(b[0]), .B(a[7]), .Z(n154) );
  XNOR U238 ( .A(b[1]), .B(n154), .Z(n156) );
  NANDN U239 ( .A(b[0]), .B(a[6]), .Z(n155) );
  NAND U240 ( .A(n156), .B(n155), .Z(n184) );
  XNOR U241 ( .A(n185), .B(n184), .Z(n186) );
  XNOR U242 ( .A(n187), .B(n186), .Z(n178) );
  NAND U243 ( .A(n2556), .B(n157), .Z(n159) );
  XNOR U244 ( .A(b[3]), .B(a[5]), .Z(n193) );
  NANDN U245 ( .A(n193), .B(n36), .Z(n158) );
  NAND U246 ( .A(n159), .B(n158), .Z(n179) );
  XNOR U247 ( .A(n178), .B(n179), .Z(n180) );
  NANDN U248 ( .A(n161), .B(n160), .Z(n165) );
  NANDN U249 ( .A(n163), .B(n162), .Z(n164) );
  NAND U250 ( .A(n165), .B(n164), .Z(n181) );
  XNOR U251 ( .A(n180), .B(n181), .Z(n172) );
  NANDN U252 ( .A(n167), .B(n166), .Z(n171) );
  NAND U253 ( .A(n169), .B(n168), .Z(n170) );
  NAND U254 ( .A(n171), .B(n170), .Z(n173) );
  XOR U255 ( .A(n172), .B(n173), .Z(n175) );
  XOR U256 ( .A(n174), .B(n175), .Z(n204) );
  XNOR U257 ( .A(n204), .B(sreg[63]), .Z(n205) );
  XNOR U258 ( .A(n206), .B(n205), .Z(c[63]) );
  NANDN U259 ( .A(n173), .B(n172), .Z(n177) );
  OR U260 ( .A(n175), .B(n174), .Z(n176) );
  AND U261 ( .A(n177), .B(n176), .Z(n245) );
  NANDN U262 ( .A(n179), .B(n178), .Z(n183) );
  NANDN U263 ( .A(n181), .B(n180), .Z(n182) );
  AND U264 ( .A(n183), .B(n182), .Z(n243) );
  NANDN U265 ( .A(n185), .B(n184), .Z(n189) );
  NANDN U266 ( .A(n187), .B(n186), .Z(n188) );
  AND U267 ( .A(n189), .B(n188), .Z(n215) );
  NANDN U268 ( .A(n2629), .B(n190), .Z(n192) );
  XOR U269 ( .A(b[7]), .B(a[2]), .Z(n230) );
  NANDN U270 ( .A(n2630), .B(n230), .Z(n191) );
  AND U271 ( .A(n192), .B(n191), .Z(n219) );
  NANDN U272 ( .A(n193), .B(n2556), .Z(n195) );
  XOR U273 ( .A(b[3]), .B(a[6]), .Z(n233) );
  NANDN U274 ( .A(n2484), .B(n233), .Z(n194) );
  NAND U275 ( .A(n195), .B(n194), .Z(n218) );
  XNOR U276 ( .A(n219), .B(n218), .Z(n221) );
  NOR U277 ( .A(n197), .B(n196), .Z(n220) );
  XOR U278 ( .A(n221), .B(n220), .Z(n213) );
  NAND U279 ( .A(b[0]), .B(a[8]), .Z(n198) );
  XNOR U280 ( .A(b[1]), .B(n198), .Z(n200) );
  NANDN U281 ( .A(b[0]), .B(a[7]), .Z(n199) );
  NAND U282 ( .A(n200), .B(n199), .Z(n227) );
  NAND U283 ( .A(n2633), .B(n201), .Z(n203) );
  XOR U284 ( .A(b[5]), .B(a[4]), .Z(n236) );
  NANDN U285 ( .A(n37), .B(n236), .Z(n202) );
  AND U286 ( .A(n203), .B(n202), .Z(n225) );
  AND U287 ( .A(b[7]), .B(a[0]), .Z(n224) );
  XOR U288 ( .A(n225), .B(n224), .Z(n226) );
  XNOR U289 ( .A(n227), .B(n226), .Z(n212) );
  XNOR U290 ( .A(n213), .B(n212), .Z(n214) );
  XNOR U291 ( .A(n215), .B(n214), .Z(n242) );
  XNOR U292 ( .A(n243), .B(n242), .Z(n244) );
  XNOR U293 ( .A(n245), .B(n244), .Z(n211) );
  NANDN U294 ( .A(n204), .B(sreg[63]), .Z(n208) );
  NANDN U295 ( .A(n206), .B(n205), .Z(n207) );
  NAND U296 ( .A(n208), .B(n207), .Z(n210) );
  XOR U297 ( .A(n210), .B(sreg[64]), .Z(n209) );
  XNOR U298 ( .A(n211), .B(n209), .Z(c[64]) );
  NANDN U299 ( .A(n213), .B(n212), .Z(n217) );
  NANDN U300 ( .A(n215), .B(n214), .Z(n216) );
  AND U301 ( .A(n217), .B(n216), .Z(n248) );
  NANDN U302 ( .A(n219), .B(n218), .Z(n223) );
  NAND U303 ( .A(n221), .B(n220), .Z(n222) );
  AND U304 ( .A(n223), .B(n222), .Z(n281) );
  NANDN U305 ( .A(n225), .B(n224), .Z(n229) );
  OR U306 ( .A(n227), .B(n226), .Z(n228) );
  AND U307 ( .A(n229), .B(n228), .Z(n279) );
  NANDN U308 ( .A(n2629), .B(n230), .Z(n232) );
  XOR U309 ( .A(b[7]), .B(a[3]), .Z(n254) );
  NANDN U310 ( .A(n2630), .B(n254), .Z(n231) );
  AND U311 ( .A(n232), .B(n231), .Z(n273) );
  NANDN U312 ( .A(n2483), .B(n233), .Z(n235) );
  XOR U313 ( .A(b[3]), .B(a[7]), .Z(n257) );
  NANDN U314 ( .A(n2484), .B(n257), .Z(n234) );
  NAND U315 ( .A(n235), .B(n234), .Z(n272) );
  XNOR U316 ( .A(n273), .B(n272), .Z(n274) );
  NAND U317 ( .A(n2633), .B(n236), .Z(n238) );
  XOR U318 ( .A(b[5]), .B(a[5]), .Z(n263) );
  NANDN U319 ( .A(n37), .B(n263), .Z(n237) );
  AND U320 ( .A(n238), .B(n237), .Z(n267) );
  AND U321 ( .A(b[7]), .B(a[1]), .Z(n266) );
  XNOR U322 ( .A(n267), .B(n266), .Z(n268) );
  NAND U323 ( .A(b[0]), .B(a[9]), .Z(n239) );
  XNOR U324 ( .A(b[1]), .B(n239), .Z(n241) );
  NANDN U325 ( .A(b[0]), .B(a[8]), .Z(n240) );
  NAND U326 ( .A(n241), .B(n240), .Z(n269) );
  XOR U327 ( .A(n268), .B(n269), .Z(n275) );
  XNOR U328 ( .A(n274), .B(n275), .Z(n278) );
  XNOR U329 ( .A(n279), .B(n278), .Z(n280) );
  XOR U330 ( .A(n281), .B(n280), .Z(n249) );
  XNOR U331 ( .A(n248), .B(n249), .Z(n250) );
  NANDN U332 ( .A(n243), .B(n242), .Z(n247) );
  NANDN U333 ( .A(n245), .B(n244), .Z(n246) );
  NAND U334 ( .A(n247), .B(n246), .Z(n251) );
  XOR U335 ( .A(n250), .B(n251), .Z(n284) );
  XNOR U336 ( .A(sreg[65]), .B(n284), .Z(n285) );
  XNOR U337 ( .A(n286), .B(n285), .Z(c[65]) );
  NANDN U338 ( .A(n249), .B(n248), .Z(n253) );
  NANDN U339 ( .A(n251), .B(n250), .Z(n252) );
  AND U340 ( .A(n253), .B(n252), .Z(n297) );
  NANDN U341 ( .A(n2629), .B(n254), .Z(n256) );
  XOR U342 ( .A(b[7]), .B(a[4]), .Z(n306) );
  NANDN U343 ( .A(n2630), .B(n306), .Z(n255) );
  AND U344 ( .A(n256), .B(n255), .Z(n325) );
  NANDN U345 ( .A(n2483), .B(n257), .Z(n259) );
  XOR U346 ( .A(b[3]), .B(a[8]), .Z(n309) );
  NANDN U347 ( .A(n2484), .B(n309), .Z(n258) );
  NAND U348 ( .A(n259), .B(n258), .Z(n324) );
  XNOR U349 ( .A(n325), .B(n324), .Z(n327) );
  NAND U350 ( .A(b[0]), .B(a[10]), .Z(n260) );
  XNOR U351 ( .A(b[1]), .B(n260), .Z(n262) );
  NANDN U352 ( .A(b[0]), .B(a[9]), .Z(n261) );
  NAND U353 ( .A(n262), .B(n261), .Z(n321) );
  NAND U354 ( .A(n2633), .B(n263), .Z(n265) );
  XOR U355 ( .A(b[5]), .B(a[6]), .Z(n315) );
  NANDN U356 ( .A(n37), .B(n315), .Z(n264) );
  AND U357 ( .A(n265), .B(n264), .Z(n319) );
  AND U358 ( .A(b[7]), .B(a[2]), .Z(n318) );
  XNOR U359 ( .A(n319), .B(n318), .Z(n320) );
  XNOR U360 ( .A(n321), .B(n320), .Z(n326) );
  XOR U361 ( .A(n327), .B(n326), .Z(n301) );
  NANDN U362 ( .A(n267), .B(n266), .Z(n271) );
  NANDN U363 ( .A(n269), .B(n268), .Z(n270) );
  AND U364 ( .A(n271), .B(n270), .Z(n300) );
  XNOR U365 ( .A(n301), .B(n300), .Z(n302) );
  NANDN U366 ( .A(n273), .B(n272), .Z(n277) );
  NANDN U367 ( .A(n275), .B(n274), .Z(n276) );
  NAND U368 ( .A(n277), .B(n276), .Z(n303) );
  XNOR U369 ( .A(n302), .B(n303), .Z(n294) );
  NANDN U370 ( .A(n279), .B(n278), .Z(n283) );
  NANDN U371 ( .A(n281), .B(n280), .Z(n282) );
  NAND U372 ( .A(n283), .B(n282), .Z(n295) );
  XNOR U373 ( .A(n294), .B(n295), .Z(n296) );
  XOR U374 ( .A(n297), .B(n296), .Z(n289) );
  XNOR U375 ( .A(n289), .B(sreg[66]), .Z(n291) );
  NANDN U376 ( .A(n284), .B(sreg[65]), .Z(n288) );
  NANDN U377 ( .A(n286), .B(n285), .Z(n287) );
  NAND U378 ( .A(n288), .B(n287), .Z(n290) );
  XOR U379 ( .A(n291), .B(n290), .Z(c[66]) );
  NANDN U380 ( .A(n289), .B(sreg[66]), .Z(n293) );
  NAND U381 ( .A(n291), .B(n290), .Z(n292) );
  AND U382 ( .A(n293), .B(n292), .Z(n368) );
  NANDN U383 ( .A(n295), .B(n294), .Z(n299) );
  NAND U384 ( .A(n297), .B(n296), .Z(n298) );
  AND U385 ( .A(n299), .B(n298), .Z(n333) );
  NANDN U386 ( .A(n301), .B(n300), .Z(n305) );
  NANDN U387 ( .A(n303), .B(n302), .Z(n304) );
  AND U388 ( .A(n305), .B(n304), .Z(n331) );
  NANDN U389 ( .A(n2629), .B(n306), .Z(n308) );
  XOR U390 ( .A(b[7]), .B(a[5]), .Z(n342) );
  NANDN U391 ( .A(n2630), .B(n342), .Z(n307) );
  AND U392 ( .A(n308), .B(n307), .Z(n361) );
  NANDN U393 ( .A(n2483), .B(n309), .Z(n311) );
  XOR U394 ( .A(b[3]), .B(a[9]), .Z(n345) );
  NANDN U395 ( .A(n2484), .B(n345), .Z(n310) );
  NAND U396 ( .A(n311), .B(n310), .Z(n360) );
  XNOR U397 ( .A(n361), .B(n360), .Z(n363) );
  NAND U398 ( .A(b[0]), .B(a[11]), .Z(n312) );
  XNOR U399 ( .A(b[1]), .B(n312), .Z(n314) );
  NANDN U400 ( .A(b[0]), .B(a[10]), .Z(n313) );
  NAND U401 ( .A(n314), .B(n313), .Z(n357) );
  NAND U402 ( .A(n2633), .B(n315), .Z(n317) );
  XOR U403 ( .A(b[5]), .B(a[7]), .Z(n351) );
  NANDN U404 ( .A(n37), .B(n351), .Z(n316) );
  AND U405 ( .A(n317), .B(n316), .Z(n355) );
  AND U406 ( .A(b[7]), .B(a[3]), .Z(n354) );
  XNOR U407 ( .A(n355), .B(n354), .Z(n356) );
  XNOR U408 ( .A(n357), .B(n356), .Z(n362) );
  XOR U409 ( .A(n363), .B(n362), .Z(n337) );
  NANDN U410 ( .A(n319), .B(n318), .Z(n323) );
  NANDN U411 ( .A(n321), .B(n320), .Z(n322) );
  AND U412 ( .A(n323), .B(n322), .Z(n336) );
  XNOR U413 ( .A(n337), .B(n336), .Z(n338) );
  NANDN U414 ( .A(n325), .B(n324), .Z(n329) );
  NAND U415 ( .A(n327), .B(n326), .Z(n328) );
  NAND U416 ( .A(n329), .B(n328), .Z(n339) );
  XNOR U417 ( .A(n338), .B(n339), .Z(n330) );
  XNOR U418 ( .A(n331), .B(n330), .Z(n332) );
  XNOR U419 ( .A(n333), .B(n332), .Z(n366) );
  XNOR U420 ( .A(sreg[67]), .B(n366), .Z(n367) );
  XNOR U421 ( .A(n368), .B(n367), .Z(c[67]) );
  NANDN U422 ( .A(n331), .B(n330), .Z(n335) );
  NANDN U423 ( .A(n333), .B(n332), .Z(n334) );
  AND U424 ( .A(n335), .B(n334), .Z(n374) );
  NANDN U425 ( .A(n337), .B(n336), .Z(n341) );
  NANDN U426 ( .A(n339), .B(n338), .Z(n340) );
  AND U427 ( .A(n341), .B(n340), .Z(n372) );
  NANDN U428 ( .A(n2629), .B(n342), .Z(n344) );
  XOR U429 ( .A(b[7]), .B(a[6]), .Z(n383) );
  NANDN U430 ( .A(n2630), .B(n383), .Z(n343) );
  AND U431 ( .A(n344), .B(n343), .Z(n402) );
  NANDN U432 ( .A(n2483), .B(n345), .Z(n347) );
  XOR U433 ( .A(b[3]), .B(a[10]), .Z(n386) );
  NANDN U434 ( .A(n2484), .B(n386), .Z(n346) );
  NAND U435 ( .A(n347), .B(n346), .Z(n401) );
  XNOR U436 ( .A(n402), .B(n401), .Z(n404) );
  NAND U437 ( .A(b[0]), .B(a[12]), .Z(n348) );
  XNOR U438 ( .A(b[1]), .B(n348), .Z(n350) );
  NANDN U439 ( .A(b[0]), .B(a[11]), .Z(n349) );
  NAND U440 ( .A(n350), .B(n349), .Z(n398) );
  NAND U441 ( .A(n2633), .B(n351), .Z(n353) );
  XOR U442 ( .A(b[5]), .B(a[8]), .Z(n389) );
  NANDN U443 ( .A(n37), .B(n389), .Z(n352) );
  AND U444 ( .A(n353), .B(n352), .Z(n396) );
  AND U445 ( .A(b[7]), .B(a[4]), .Z(n395) );
  XNOR U446 ( .A(n396), .B(n395), .Z(n397) );
  XNOR U447 ( .A(n398), .B(n397), .Z(n403) );
  XOR U448 ( .A(n404), .B(n403), .Z(n378) );
  NANDN U449 ( .A(n355), .B(n354), .Z(n359) );
  NANDN U450 ( .A(n357), .B(n356), .Z(n358) );
  AND U451 ( .A(n359), .B(n358), .Z(n377) );
  XNOR U452 ( .A(n378), .B(n377), .Z(n379) );
  NANDN U453 ( .A(n361), .B(n360), .Z(n365) );
  NAND U454 ( .A(n363), .B(n362), .Z(n364) );
  NAND U455 ( .A(n365), .B(n364), .Z(n380) );
  XNOR U456 ( .A(n379), .B(n380), .Z(n371) );
  XNOR U457 ( .A(n372), .B(n371), .Z(n373) );
  XNOR U458 ( .A(n374), .B(n373), .Z(n407) );
  XNOR U459 ( .A(sreg[68]), .B(n407), .Z(n409) );
  NANDN U460 ( .A(sreg[67]), .B(n366), .Z(n370) );
  NAND U461 ( .A(n368), .B(n367), .Z(n369) );
  NAND U462 ( .A(n370), .B(n369), .Z(n408) );
  XNOR U463 ( .A(n409), .B(n408), .Z(c[68]) );
  NANDN U464 ( .A(n372), .B(n371), .Z(n376) );
  NANDN U465 ( .A(n374), .B(n373), .Z(n375) );
  AND U466 ( .A(n376), .B(n375), .Z(n419) );
  NANDN U467 ( .A(n378), .B(n377), .Z(n382) );
  NANDN U468 ( .A(n380), .B(n379), .Z(n381) );
  AND U469 ( .A(n382), .B(n381), .Z(n418) );
  NANDN U470 ( .A(n2629), .B(n383), .Z(n385) );
  XOR U471 ( .A(b[7]), .B(a[7]), .Z(n429) );
  NANDN U472 ( .A(n2630), .B(n429), .Z(n384) );
  AND U473 ( .A(n385), .B(n384), .Z(n448) );
  NANDN U474 ( .A(n2483), .B(n386), .Z(n388) );
  XOR U475 ( .A(b[3]), .B(a[11]), .Z(n432) );
  NANDN U476 ( .A(n2484), .B(n432), .Z(n387) );
  NAND U477 ( .A(n388), .B(n387), .Z(n447) );
  XNOR U478 ( .A(n448), .B(n447), .Z(n450) );
  NAND U479 ( .A(n2633), .B(n389), .Z(n391) );
  XOR U480 ( .A(b[5]), .B(a[9]), .Z(n438) );
  NANDN U481 ( .A(n37), .B(n438), .Z(n390) );
  AND U482 ( .A(n391), .B(n390), .Z(n442) );
  AND U483 ( .A(b[7]), .B(a[5]), .Z(n441) );
  XNOR U484 ( .A(n442), .B(n441), .Z(n443) );
  NAND U485 ( .A(b[0]), .B(a[13]), .Z(n392) );
  XNOR U486 ( .A(b[1]), .B(n392), .Z(n394) );
  NANDN U487 ( .A(b[0]), .B(a[12]), .Z(n393) );
  NAND U488 ( .A(n394), .B(n393), .Z(n444) );
  XNOR U489 ( .A(n443), .B(n444), .Z(n449) );
  XOR U490 ( .A(n450), .B(n449), .Z(n424) );
  NANDN U491 ( .A(n396), .B(n395), .Z(n400) );
  NANDN U492 ( .A(n398), .B(n397), .Z(n399) );
  AND U493 ( .A(n400), .B(n399), .Z(n423) );
  XNOR U494 ( .A(n424), .B(n423), .Z(n425) );
  NANDN U495 ( .A(n402), .B(n401), .Z(n406) );
  NAND U496 ( .A(n404), .B(n403), .Z(n405) );
  NAND U497 ( .A(n406), .B(n405), .Z(n426) );
  XNOR U498 ( .A(n425), .B(n426), .Z(n417) );
  XOR U499 ( .A(n418), .B(n417), .Z(n420) );
  XOR U500 ( .A(n419), .B(n420), .Z(n412) );
  XNOR U501 ( .A(n412), .B(sreg[69]), .Z(n414) );
  NANDN U502 ( .A(sreg[68]), .B(n407), .Z(n411) );
  NAND U503 ( .A(n409), .B(n408), .Z(n410) );
  AND U504 ( .A(n411), .B(n410), .Z(n413) );
  XOR U505 ( .A(n414), .B(n413), .Z(c[69]) );
  NANDN U506 ( .A(n412), .B(sreg[69]), .Z(n416) );
  NAND U507 ( .A(n414), .B(n413), .Z(n415) );
  AND U508 ( .A(n416), .B(n415), .Z(n491) );
  NANDN U509 ( .A(n418), .B(n417), .Z(n422) );
  OR U510 ( .A(n420), .B(n419), .Z(n421) );
  AND U511 ( .A(n422), .B(n421), .Z(n456) );
  NANDN U512 ( .A(n424), .B(n423), .Z(n428) );
  NANDN U513 ( .A(n426), .B(n425), .Z(n427) );
  AND U514 ( .A(n428), .B(n427), .Z(n454) );
  NANDN U515 ( .A(n2629), .B(n429), .Z(n431) );
  XOR U516 ( .A(b[7]), .B(a[8]), .Z(n465) );
  NANDN U517 ( .A(n2630), .B(n465), .Z(n430) );
  AND U518 ( .A(n431), .B(n430), .Z(n484) );
  NANDN U519 ( .A(n2483), .B(n432), .Z(n434) );
  XOR U520 ( .A(b[3]), .B(a[12]), .Z(n468) );
  NANDN U521 ( .A(n2484), .B(n468), .Z(n433) );
  NAND U522 ( .A(n434), .B(n433), .Z(n483) );
  XNOR U523 ( .A(n484), .B(n483), .Z(n486) );
  NAND U524 ( .A(b[0]), .B(a[14]), .Z(n435) );
  XNOR U525 ( .A(b[1]), .B(n435), .Z(n437) );
  NANDN U526 ( .A(b[0]), .B(a[13]), .Z(n436) );
  NAND U527 ( .A(n437), .B(n436), .Z(n480) );
  NAND U528 ( .A(n2633), .B(n438), .Z(n440) );
  XOR U529 ( .A(b[5]), .B(a[10]), .Z(n474) );
  NANDN U530 ( .A(n37), .B(n474), .Z(n439) );
  AND U531 ( .A(n440), .B(n439), .Z(n478) );
  AND U532 ( .A(b[7]), .B(a[6]), .Z(n477) );
  XNOR U533 ( .A(n478), .B(n477), .Z(n479) );
  XNOR U534 ( .A(n480), .B(n479), .Z(n485) );
  XOR U535 ( .A(n486), .B(n485), .Z(n460) );
  NANDN U536 ( .A(n442), .B(n441), .Z(n446) );
  NANDN U537 ( .A(n444), .B(n443), .Z(n445) );
  AND U538 ( .A(n446), .B(n445), .Z(n459) );
  XNOR U539 ( .A(n460), .B(n459), .Z(n461) );
  NANDN U540 ( .A(n448), .B(n447), .Z(n452) );
  NAND U541 ( .A(n450), .B(n449), .Z(n451) );
  NAND U542 ( .A(n452), .B(n451), .Z(n462) );
  XNOR U543 ( .A(n461), .B(n462), .Z(n453) );
  XNOR U544 ( .A(n454), .B(n453), .Z(n455) );
  XNOR U545 ( .A(n456), .B(n455), .Z(n489) );
  XNOR U546 ( .A(sreg[70]), .B(n489), .Z(n490) );
  XNOR U547 ( .A(n491), .B(n490), .Z(c[70]) );
  NANDN U548 ( .A(n454), .B(n453), .Z(n458) );
  NANDN U549 ( .A(n456), .B(n455), .Z(n457) );
  AND U550 ( .A(n458), .B(n457), .Z(n497) );
  NANDN U551 ( .A(n460), .B(n459), .Z(n464) );
  NANDN U552 ( .A(n462), .B(n461), .Z(n463) );
  AND U553 ( .A(n464), .B(n463), .Z(n495) );
  NANDN U554 ( .A(n2629), .B(n465), .Z(n467) );
  XOR U555 ( .A(b[7]), .B(a[9]), .Z(n506) );
  NANDN U556 ( .A(n2630), .B(n506), .Z(n466) );
  AND U557 ( .A(n467), .B(n466), .Z(n525) );
  NANDN U558 ( .A(n2483), .B(n468), .Z(n470) );
  XOR U559 ( .A(b[3]), .B(a[13]), .Z(n509) );
  NANDN U560 ( .A(n2484), .B(n509), .Z(n469) );
  NAND U561 ( .A(n470), .B(n469), .Z(n524) );
  XNOR U562 ( .A(n525), .B(n524), .Z(n527) );
  NAND U563 ( .A(b[0]), .B(a[15]), .Z(n471) );
  XNOR U564 ( .A(b[1]), .B(n471), .Z(n473) );
  NANDN U565 ( .A(b[0]), .B(a[14]), .Z(n472) );
  NAND U566 ( .A(n473), .B(n472), .Z(n521) );
  NAND U567 ( .A(n2633), .B(n474), .Z(n476) );
  XOR U568 ( .A(b[5]), .B(a[11]), .Z(n515) );
  NANDN U569 ( .A(n37), .B(n515), .Z(n475) );
  AND U570 ( .A(n476), .B(n475), .Z(n519) );
  AND U571 ( .A(b[7]), .B(a[7]), .Z(n518) );
  XNOR U572 ( .A(n519), .B(n518), .Z(n520) );
  XNOR U573 ( .A(n521), .B(n520), .Z(n526) );
  XOR U574 ( .A(n527), .B(n526), .Z(n501) );
  NANDN U575 ( .A(n478), .B(n477), .Z(n482) );
  NANDN U576 ( .A(n480), .B(n479), .Z(n481) );
  AND U577 ( .A(n482), .B(n481), .Z(n500) );
  XNOR U578 ( .A(n501), .B(n500), .Z(n502) );
  NANDN U579 ( .A(n484), .B(n483), .Z(n488) );
  NAND U580 ( .A(n486), .B(n485), .Z(n487) );
  NAND U581 ( .A(n488), .B(n487), .Z(n503) );
  XNOR U582 ( .A(n502), .B(n503), .Z(n494) );
  XNOR U583 ( .A(n495), .B(n494), .Z(n496) );
  XNOR U584 ( .A(n497), .B(n496), .Z(n530) );
  XNOR U585 ( .A(sreg[71]), .B(n530), .Z(n532) );
  NANDN U586 ( .A(sreg[70]), .B(n489), .Z(n493) );
  NAND U587 ( .A(n491), .B(n490), .Z(n492) );
  NAND U588 ( .A(n493), .B(n492), .Z(n531) );
  XNOR U589 ( .A(n532), .B(n531), .Z(c[71]) );
  NANDN U590 ( .A(n495), .B(n494), .Z(n499) );
  NANDN U591 ( .A(n497), .B(n496), .Z(n498) );
  AND U592 ( .A(n499), .B(n498), .Z(n538) );
  NANDN U593 ( .A(n501), .B(n500), .Z(n505) );
  NANDN U594 ( .A(n503), .B(n502), .Z(n504) );
  AND U595 ( .A(n505), .B(n504), .Z(n536) );
  NANDN U596 ( .A(n2629), .B(n506), .Z(n508) );
  XOR U597 ( .A(b[7]), .B(a[10]), .Z(n547) );
  NANDN U598 ( .A(n2630), .B(n547), .Z(n507) );
  AND U599 ( .A(n508), .B(n507), .Z(n566) );
  NANDN U600 ( .A(n2483), .B(n509), .Z(n511) );
  XOR U601 ( .A(b[3]), .B(a[14]), .Z(n550) );
  NANDN U602 ( .A(n2484), .B(n550), .Z(n510) );
  NAND U603 ( .A(n511), .B(n510), .Z(n565) );
  XNOR U604 ( .A(n566), .B(n565), .Z(n568) );
  NAND U605 ( .A(b[0]), .B(a[16]), .Z(n512) );
  XNOR U606 ( .A(b[1]), .B(n512), .Z(n514) );
  NANDN U607 ( .A(b[0]), .B(a[15]), .Z(n513) );
  NAND U608 ( .A(n514), .B(n513), .Z(n562) );
  NAND U609 ( .A(n2633), .B(n515), .Z(n517) );
  XOR U610 ( .A(b[5]), .B(a[12]), .Z(n553) );
  NANDN U611 ( .A(n37), .B(n553), .Z(n516) );
  AND U612 ( .A(n517), .B(n516), .Z(n560) );
  AND U613 ( .A(b[7]), .B(a[8]), .Z(n559) );
  XNOR U614 ( .A(n560), .B(n559), .Z(n561) );
  XNOR U615 ( .A(n562), .B(n561), .Z(n567) );
  XOR U616 ( .A(n568), .B(n567), .Z(n542) );
  NANDN U617 ( .A(n519), .B(n518), .Z(n523) );
  NANDN U618 ( .A(n521), .B(n520), .Z(n522) );
  AND U619 ( .A(n523), .B(n522), .Z(n541) );
  XNOR U620 ( .A(n542), .B(n541), .Z(n543) );
  NANDN U621 ( .A(n525), .B(n524), .Z(n529) );
  NAND U622 ( .A(n527), .B(n526), .Z(n528) );
  NAND U623 ( .A(n529), .B(n528), .Z(n544) );
  XNOR U624 ( .A(n543), .B(n544), .Z(n535) );
  XNOR U625 ( .A(n536), .B(n535), .Z(n537) );
  XNOR U626 ( .A(n538), .B(n537), .Z(n571) );
  XNOR U627 ( .A(sreg[72]), .B(n571), .Z(n573) );
  NANDN U628 ( .A(sreg[71]), .B(n530), .Z(n534) );
  NAND U629 ( .A(n532), .B(n531), .Z(n533) );
  NAND U630 ( .A(n534), .B(n533), .Z(n572) );
  XNOR U631 ( .A(n573), .B(n572), .Z(c[72]) );
  NANDN U632 ( .A(n536), .B(n535), .Z(n540) );
  NANDN U633 ( .A(n538), .B(n537), .Z(n539) );
  AND U634 ( .A(n540), .B(n539), .Z(n579) );
  NANDN U635 ( .A(n542), .B(n541), .Z(n546) );
  NANDN U636 ( .A(n544), .B(n543), .Z(n545) );
  AND U637 ( .A(n546), .B(n545), .Z(n577) );
  NANDN U638 ( .A(n2629), .B(n547), .Z(n549) );
  XOR U639 ( .A(b[7]), .B(a[11]), .Z(n588) );
  NANDN U640 ( .A(n2630), .B(n588), .Z(n548) );
  AND U641 ( .A(n549), .B(n548), .Z(n607) );
  NANDN U642 ( .A(n2483), .B(n550), .Z(n552) );
  XOR U643 ( .A(b[3]), .B(a[15]), .Z(n591) );
  NANDN U644 ( .A(n2484), .B(n591), .Z(n551) );
  NAND U645 ( .A(n552), .B(n551), .Z(n606) );
  XNOR U646 ( .A(n607), .B(n606), .Z(n609) );
  NAND U647 ( .A(n2633), .B(n553), .Z(n555) );
  XOR U648 ( .A(b[5]), .B(a[13]), .Z(n594) );
  NANDN U649 ( .A(n37), .B(n594), .Z(n554) );
  AND U650 ( .A(n555), .B(n554), .Z(n601) );
  AND U651 ( .A(b[7]), .B(a[9]), .Z(n600) );
  XNOR U652 ( .A(n601), .B(n600), .Z(n602) );
  NAND U653 ( .A(b[0]), .B(a[17]), .Z(n556) );
  XNOR U654 ( .A(b[1]), .B(n556), .Z(n558) );
  NANDN U655 ( .A(b[0]), .B(a[16]), .Z(n557) );
  NAND U656 ( .A(n558), .B(n557), .Z(n603) );
  XNOR U657 ( .A(n602), .B(n603), .Z(n608) );
  XOR U658 ( .A(n609), .B(n608), .Z(n583) );
  NANDN U659 ( .A(n560), .B(n559), .Z(n564) );
  NANDN U660 ( .A(n562), .B(n561), .Z(n563) );
  AND U661 ( .A(n564), .B(n563), .Z(n582) );
  XNOR U662 ( .A(n583), .B(n582), .Z(n584) );
  NANDN U663 ( .A(n566), .B(n565), .Z(n570) );
  NAND U664 ( .A(n568), .B(n567), .Z(n569) );
  NAND U665 ( .A(n570), .B(n569), .Z(n585) );
  XNOR U666 ( .A(n584), .B(n585), .Z(n576) );
  XNOR U667 ( .A(n577), .B(n576), .Z(n578) );
  XNOR U668 ( .A(n579), .B(n578), .Z(n612) );
  XNOR U669 ( .A(sreg[73]), .B(n612), .Z(n614) );
  NANDN U670 ( .A(sreg[72]), .B(n571), .Z(n575) );
  NAND U671 ( .A(n573), .B(n572), .Z(n574) );
  NAND U672 ( .A(n575), .B(n574), .Z(n613) );
  XNOR U673 ( .A(n614), .B(n613), .Z(c[73]) );
  NANDN U674 ( .A(n577), .B(n576), .Z(n581) );
  NANDN U675 ( .A(n579), .B(n578), .Z(n580) );
  AND U676 ( .A(n581), .B(n580), .Z(n620) );
  NANDN U677 ( .A(n583), .B(n582), .Z(n587) );
  NANDN U678 ( .A(n585), .B(n584), .Z(n586) );
  AND U679 ( .A(n587), .B(n586), .Z(n618) );
  NANDN U680 ( .A(n2629), .B(n588), .Z(n590) );
  XOR U681 ( .A(b[7]), .B(a[12]), .Z(n629) );
  NANDN U682 ( .A(n2630), .B(n629), .Z(n589) );
  AND U683 ( .A(n590), .B(n589), .Z(n648) );
  NANDN U684 ( .A(n2483), .B(n591), .Z(n593) );
  XOR U685 ( .A(b[3]), .B(a[16]), .Z(n632) );
  NANDN U686 ( .A(n2484), .B(n632), .Z(n592) );
  NAND U687 ( .A(n593), .B(n592), .Z(n647) );
  XNOR U688 ( .A(n648), .B(n647), .Z(n650) );
  NAND U689 ( .A(n2633), .B(n594), .Z(n596) );
  XOR U690 ( .A(b[5]), .B(a[14]), .Z(n638) );
  NANDN U691 ( .A(n37), .B(n638), .Z(n595) );
  AND U692 ( .A(n596), .B(n595), .Z(n642) );
  AND U693 ( .A(b[7]), .B(a[10]), .Z(n641) );
  XNOR U694 ( .A(n642), .B(n641), .Z(n643) );
  NAND U695 ( .A(b[0]), .B(a[18]), .Z(n597) );
  XNOR U696 ( .A(b[1]), .B(n597), .Z(n599) );
  NANDN U697 ( .A(b[0]), .B(a[17]), .Z(n598) );
  NAND U698 ( .A(n599), .B(n598), .Z(n644) );
  XNOR U699 ( .A(n643), .B(n644), .Z(n649) );
  XOR U700 ( .A(n650), .B(n649), .Z(n624) );
  NANDN U701 ( .A(n601), .B(n600), .Z(n605) );
  NANDN U702 ( .A(n603), .B(n602), .Z(n604) );
  AND U703 ( .A(n605), .B(n604), .Z(n623) );
  XNOR U704 ( .A(n624), .B(n623), .Z(n625) );
  NANDN U705 ( .A(n607), .B(n606), .Z(n611) );
  NAND U706 ( .A(n609), .B(n608), .Z(n610) );
  NAND U707 ( .A(n611), .B(n610), .Z(n626) );
  XNOR U708 ( .A(n625), .B(n626), .Z(n617) );
  XNOR U709 ( .A(n618), .B(n617), .Z(n619) );
  XNOR U710 ( .A(n620), .B(n619), .Z(n653) );
  XNOR U711 ( .A(sreg[74]), .B(n653), .Z(n655) );
  NANDN U712 ( .A(sreg[73]), .B(n612), .Z(n616) );
  NAND U713 ( .A(n614), .B(n613), .Z(n615) );
  NAND U714 ( .A(n616), .B(n615), .Z(n654) );
  XNOR U715 ( .A(n655), .B(n654), .Z(c[74]) );
  NANDN U716 ( .A(n618), .B(n617), .Z(n622) );
  NANDN U717 ( .A(n620), .B(n619), .Z(n621) );
  AND U718 ( .A(n622), .B(n621), .Z(n661) );
  NANDN U719 ( .A(n624), .B(n623), .Z(n628) );
  NANDN U720 ( .A(n626), .B(n625), .Z(n627) );
  AND U721 ( .A(n628), .B(n627), .Z(n659) );
  NANDN U722 ( .A(n2629), .B(n629), .Z(n631) );
  XOR U723 ( .A(b[7]), .B(a[13]), .Z(n670) );
  NANDN U724 ( .A(n2630), .B(n670), .Z(n630) );
  AND U725 ( .A(n631), .B(n630), .Z(n689) );
  NANDN U726 ( .A(n2483), .B(n632), .Z(n634) );
  XOR U727 ( .A(b[3]), .B(a[17]), .Z(n673) );
  NANDN U728 ( .A(n2484), .B(n673), .Z(n633) );
  NAND U729 ( .A(n634), .B(n633), .Z(n688) );
  XNOR U730 ( .A(n689), .B(n688), .Z(n691) );
  NAND U731 ( .A(b[0]), .B(a[19]), .Z(n635) );
  XNOR U732 ( .A(b[1]), .B(n635), .Z(n637) );
  NANDN U733 ( .A(b[0]), .B(a[18]), .Z(n636) );
  NAND U734 ( .A(n637), .B(n636), .Z(n685) );
  NAND U735 ( .A(n2633), .B(n638), .Z(n640) );
  XOR U736 ( .A(b[5]), .B(a[15]), .Z(n679) );
  NANDN U737 ( .A(n37), .B(n679), .Z(n639) );
  AND U738 ( .A(n640), .B(n639), .Z(n683) );
  AND U739 ( .A(b[7]), .B(a[11]), .Z(n682) );
  XNOR U740 ( .A(n683), .B(n682), .Z(n684) );
  XNOR U741 ( .A(n685), .B(n684), .Z(n690) );
  XOR U742 ( .A(n691), .B(n690), .Z(n665) );
  NANDN U743 ( .A(n642), .B(n641), .Z(n646) );
  NANDN U744 ( .A(n644), .B(n643), .Z(n645) );
  AND U745 ( .A(n646), .B(n645), .Z(n664) );
  XNOR U746 ( .A(n665), .B(n664), .Z(n666) );
  NANDN U747 ( .A(n648), .B(n647), .Z(n652) );
  NAND U748 ( .A(n650), .B(n649), .Z(n651) );
  NAND U749 ( .A(n652), .B(n651), .Z(n667) );
  XNOR U750 ( .A(n666), .B(n667), .Z(n658) );
  XNOR U751 ( .A(n659), .B(n658), .Z(n660) );
  XNOR U752 ( .A(n661), .B(n660), .Z(n694) );
  XNOR U753 ( .A(sreg[75]), .B(n694), .Z(n696) );
  NANDN U754 ( .A(sreg[74]), .B(n653), .Z(n657) );
  NAND U755 ( .A(n655), .B(n654), .Z(n656) );
  NAND U756 ( .A(n657), .B(n656), .Z(n695) );
  XNOR U757 ( .A(n696), .B(n695), .Z(c[75]) );
  NANDN U758 ( .A(n659), .B(n658), .Z(n663) );
  NANDN U759 ( .A(n661), .B(n660), .Z(n662) );
  AND U760 ( .A(n663), .B(n662), .Z(n702) );
  NANDN U761 ( .A(n665), .B(n664), .Z(n669) );
  NANDN U762 ( .A(n667), .B(n666), .Z(n668) );
  AND U763 ( .A(n669), .B(n668), .Z(n700) );
  NANDN U764 ( .A(n2629), .B(n670), .Z(n672) );
  XOR U765 ( .A(b[7]), .B(a[14]), .Z(n711) );
  NANDN U766 ( .A(n2630), .B(n711), .Z(n671) );
  AND U767 ( .A(n672), .B(n671), .Z(n730) );
  NANDN U768 ( .A(n2483), .B(n673), .Z(n675) );
  XOR U769 ( .A(b[3]), .B(a[18]), .Z(n714) );
  NANDN U770 ( .A(n2484), .B(n714), .Z(n674) );
  NAND U771 ( .A(n675), .B(n674), .Z(n729) );
  XNOR U772 ( .A(n730), .B(n729), .Z(n732) );
  NAND U773 ( .A(b[0]), .B(a[20]), .Z(n676) );
  XNOR U774 ( .A(b[1]), .B(n676), .Z(n678) );
  NANDN U775 ( .A(b[0]), .B(a[19]), .Z(n677) );
  NAND U776 ( .A(n678), .B(n677), .Z(n726) );
  NAND U777 ( .A(n2633), .B(n679), .Z(n681) );
  XOR U778 ( .A(b[5]), .B(a[16]), .Z(n717) );
  NANDN U779 ( .A(n37), .B(n717), .Z(n680) );
  AND U780 ( .A(n681), .B(n680), .Z(n724) );
  AND U781 ( .A(b[7]), .B(a[12]), .Z(n723) );
  XNOR U782 ( .A(n724), .B(n723), .Z(n725) );
  XNOR U783 ( .A(n726), .B(n725), .Z(n731) );
  XOR U784 ( .A(n732), .B(n731), .Z(n706) );
  NANDN U785 ( .A(n683), .B(n682), .Z(n687) );
  NANDN U786 ( .A(n685), .B(n684), .Z(n686) );
  AND U787 ( .A(n687), .B(n686), .Z(n705) );
  XNOR U788 ( .A(n706), .B(n705), .Z(n707) );
  NANDN U789 ( .A(n689), .B(n688), .Z(n693) );
  NAND U790 ( .A(n691), .B(n690), .Z(n692) );
  NAND U791 ( .A(n693), .B(n692), .Z(n708) );
  XNOR U792 ( .A(n707), .B(n708), .Z(n699) );
  XNOR U793 ( .A(n700), .B(n699), .Z(n701) );
  XNOR U794 ( .A(n702), .B(n701), .Z(n735) );
  XNOR U795 ( .A(sreg[76]), .B(n735), .Z(n737) );
  NANDN U796 ( .A(sreg[75]), .B(n694), .Z(n698) );
  NAND U797 ( .A(n696), .B(n695), .Z(n697) );
  NAND U798 ( .A(n698), .B(n697), .Z(n736) );
  XNOR U799 ( .A(n737), .B(n736), .Z(c[76]) );
  NANDN U800 ( .A(n700), .B(n699), .Z(n704) );
  NANDN U801 ( .A(n702), .B(n701), .Z(n703) );
  AND U802 ( .A(n704), .B(n703), .Z(n743) );
  NANDN U803 ( .A(n706), .B(n705), .Z(n710) );
  NANDN U804 ( .A(n708), .B(n707), .Z(n709) );
  AND U805 ( .A(n710), .B(n709), .Z(n741) );
  NANDN U806 ( .A(n2629), .B(n711), .Z(n713) );
  XOR U807 ( .A(b[7]), .B(a[15]), .Z(n752) );
  NANDN U808 ( .A(n2630), .B(n752), .Z(n712) );
  AND U809 ( .A(n713), .B(n712), .Z(n771) );
  NANDN U810 ( .A(n2483), .B(n714), .Z(n716) );
  XOR U811 ( .A(b[3]), .B(a[19]), .Z(n755) );
  NANDN U812 ( .A(n2484), .B(n755), .Z(n715) );
  NAND U813 ( .A(n716), .B(n715), .Z(n770) );
  XNOR U814 ( .A(n771), .B(n770), .Z(n773) );
  NAND U815 ( .A(n2633), .B(n717), .Z(n719) );
  XOR U816 ( .A(b[5]), .B(a[17]), .Z(n761) );
  NANDN U817 ( .A(n37), .B(n761), .Z(n718) );
  AND U818 ( .A(n719), .B(n718), .Z(n765) );
  AND U819 ( .A(b[7]), .B(a[13]), .Z(n764) );
  XNOR U820 ( .A(n765), .B(n764), .Z(n766) );
  NAND U821 ( .A(b[0]), .B(a[21]), .Z(n720) );
  XNOR U822 ( .A(b[1]), .B(n720), .Z(n722) );
  NANDN U823 ( .A(b[0]), .B(a[20]), .Z(n721) );
  NAND U824 ( .A(n722), .B(n721), .Z(n767) );
  XNOR U825 ( .A(n766), .B(n767), .Z(n772) );
  XOR U826 ( .A(n773), .B(n772), .Z(n747) );
  NANDN U827 ( .A(n724), .B(n723), .Z(n728) );
  NANDN U828 ( .A(n726), .B(n725), .Z(n727) );
  AND U829 ( .A(n728), .B(n727), .Z(n746) );
  XNOR U830 ( .A(n747), .B(n746), .Z(n748) );
  NANDN U831 ( .A(n730), .B(n729), .Z(n734) );
  NAND U832 ( .A(n732), .B(n731), .Z(n733) );
  NAND U833 ( .A(n734), .B(n733), .Z(n749) );
  XNOR U834 ( .A(n748), .B(n749), .Z(n740) );
  XNOR U835 ( .A(n741), .B(n740), .Z(n742) );
  XNOR U836 ( .A(n743), .B(n742), .Z(n776) );
  XNOR U837 ( .A(sreg[77]), .B(n776), .Z(n778) );
  NANDN U838 ( .A(sreg[76]), .B(n735), .Z(n739) );
  NAND U839 ( .A(n737), .B(n736), .Z(n738) );
  NAND U840 ( .A(n739), .B(n738), .Z(n777) );
  XNOR U841 ( .A(n778), .B(n777), .Z(c[77]) );
  NANDN U842 ( .A(n741), .B(n740), .Z(n745) );
  NANDN U843 ( .A(n743), .B(n742), .Z(n744) );
  AND U844 ( .A(n745), .B(n744), .Z(n784) );
  NANDN U845 ( .A(n747), .B(n746), .Z(n751) );
  NANDN U846 ( .A(n749), .B(n748), .Z(n750) );
  AND U847 ( .A(n751), .B(n750), .Z(n782) );
  NANDN U848 ( .A(n2629), .B(n752), .Z(n754) );
  XOR U849 ( .A(b[7]), .B(a[16]), .Z(n793) );
  NANDN U850 ( .A(n2630), .B(n793), .Z(n753) );
  AND U851 ( .A(n754), .B(n753), .Z(n812) );
  NANDN U852 ( .A(n2483), .B(n755), .Z(n757) );
  XOR U853 ( .A(b[3]), .B(a[20]), .Z(n796) );
  NANDN U854 ( .A(n2484), .B(n796), .Z(n756) );
  NAND U855 ( .A(n757), .B(n756), .Z(n811) );
  XNOR U856 ( .A(n812), .B(n811), .Z(n814) );
  AND U857 ( .A(b[0]), .B(a[22]), .Z(n758) );
  XOR U858 ( .A(b[1]), .B(n758), .Z(n760) );
  NANDN U859 ( .A(b[0]), .B(a[21]), .Z(n759) );
  AND U860 ( .A(n760), .B(n759), .Z(n807) );
  NAND U861 ( .A(n2633), .B(n761), .Z(n763) );
  XOR U862 ( .A(b[5]), .B(a[18]), .Z(n802) );
  NANDN U863 ( .A(n37), .B(n802), .Z(n762) );
  AND U864 ( .A(n763), .B(n762), .Z(n806) );
  AND U865 ( .A(b[7]), .B(a[14]), .Z(n805) );
  XOR U866 ( .A(n806), .B(n805), .Z(n808) );
  XNOR U867 ( .A(n807), .B(n808), .Z(n813) );
  XOR U868 ( .A(n814), .B(n813), .Z(n788) );
  NANDN U869 ( .A(n765), .B(n764), .Z(n769) );
  NANDN U870 ( .A(n767), .B(n766), .Z(n768) );
  AND U871 ( .A(n769), .B(n768), .Z(n787) );
  XNOR U872 ( .A(n788), .B(n787), .Z(n789) );
  NANDN U873 ( .A(n771), .B(n770), .Z(n775) );
  NAND U874 ( .A(n773), .B(n772), .Z(n774) );
  NAND U875 ( .A(n775), .B(n774), .Z(n790) );
  XNOR U876 ( .A(n789), .B(n790), .Z(n781) );
  XNOR U877 ( .A(n782), .B(n781), .Z(n783) );
  XNOR U878 ( .A(n784), .B(n783), .Z(n817) );
  XNOR U879 ( .A(sreg[78]), .B(n817), .Z(n819) );
  NANDN U880 ( .A(sreg[77]), .B(n776), .Z(n780) );
  NAND U881 ( .A(n778), .B(n777), .Z(n779) );
  NAND U882 ( .A(n780), .B(n779), .Z(n818) );
  XNOR U883 ( .A(n819), .B(n818), .Z(c[78]) );
  NANDN U884 ( .A(n782), .B(n781), .Z(n786) );
  NANDN U885 ( .A(n784), .B(n783), .Z(n785) );
  AND U886 ( .A(n786), .B(n785), .Z(n825) );
  NANDN U887 ( .A(n788), .B(n787), .Z(n792) );
  NANDN U888 ( .A(n790), .B(n789), .Z(n791) );
  AND U889 ( .A(n792), .B(n791), .Z(n823) );
  NANDN U890 ( .A(n2629), .B(n793), .Z(n795) );
  XOR U891 ( .A(b[7]), .B(a[17]), .Z(n834) );
  NANDN U892 ( .A(n2630), .B(n834), .Z(n794) );
  AND U893 ( .A(n795), .B(n794), .Z(n853) );
  NANDN U894 ( .A(n2483), .B(n796), .Z(n798) );
  XOR U895 ( .A(b[3]), .B(a[21]), .Z(n837) );
  NANDN U896 ( .A(n2484), .B(n837), .Z(n797) );
  NAND U897 ( .A(n798), .B(n797), .Z(n852) );
  XNOR U898 ( .A(n853), .B(n852), .Z(n855) );
  NAND U899 ( .A(b[0]), .B(a[23]), .Z(n799) );
  XNOR U900 ( .A(b[1]), .B(n799), .Z(n801) );
  NANDN U901 ( .A(b[0]), .B(a[22]), .Z(n800) );
  NAND U902 ( .A(n801), .B(n800), .Z(n849) );
  NAND U903 ( .A(n2633), .B(n802), .Z(n804) );
  XOR U904 ( .A(b[5]), .B(a[19]), .Z(n843) );
  NANDN U905 ( .A(n37), .B(n843), .Z(n803) );
  AND U906 ( .A(n804), .B(n803), .Z(n847) );
  AND U907 ( .A(b[7]), .B(a[15]), .Z(n846) );
  XNOR U908 ( .A(n847), .B(n846), .Z(n848) );
  XNOR U909 ( .A(n849), .B(n848), .Z(n854) );
  XOR U910 ( .A(n855), .B(n854), .Z(n829) );
  NANDN U911 ( .A(n806), .B(n805), .Z(n810) );
  NANDN U912 ( .A(n808), .B(n807), .Z(n809) );
  AND U913 ( .A(n810), .B(n809), .Z(n828) );
  XNOR U914 ( .A(n829), .B(n828), .Z(n830) );
  NANDN U915 ( .A(n812), .B(n811), .Z(n816) );
  NAND U916 ( .A(n814), .B(n813), .Z(n815) );
  NAND U917 ( .A(n816), .B(n815), .Z(n831) );
  XNOR U918 ( .A(n830), .B(n831), .Z(n822) );
  XNOR U919 ( .A(n823), .B(n822), .Z(n824) );
  XNOR U920 ( .A(n825), .B(n824), .Z(n858) );
  XNOR U921 ( .A(sreg[79]), .B(n858), .Z(n860) );
  NANDN U922 ( .A(sreg[78]), .B(n817), .Z(n821) );
  NAND U923 ( .A(n819), .B(n818), .Z(n820) );
  NAND U924 ( .A(n821), .B(n820), .Z(n859) );
  XNOR U925 ( .A(n860), .B(n859), .Z(c[79]) );
  NANDN U926 ( .A(n823), .B(n822), .Z(n827) );
  NANDN U927 ( .A(n825), .B(n824), .Z(n826) );
  AND U928 ( .A(n827), .B(n826), .Z(n866) );
  NANDN U929 ( .A(n829), .B(n828), .Z(n833) );
  NANDN U930 ( .A(n831), .B(n830), .Z(n832) );
  AND U931 ( .A(n833), .B(n832), .Z(n864) );
  NANDN U932 ( .A(n2629), .B(n834), .Z(n836) );
  XOR U933 ( .A(b[7]), .B(a[18]), .Z(n875) );
  NANDN U934 ( .A(n2630), .B(n875), .Z(n835) );
  AND U935 ( .A(n836), .B(n835), .Z(n894) );
  NANDN U936 ( .A(n2483), .B(n837), .Z(n839) );
  XOR U937 ( .A(b[3]), .B(a[22]), .Z(n878) );
  NANDN U938 ( .A(n2484), .B(n878), .Z(n838) );
  NAND U939 ( .A(n839), .B(n838), .Z(n893) );
  XNOR U940 ( .A(n894), .B(n893), .Z(n896) );
  NAND U941 ( .A(b[0]), .B(a[24]), .Z(n840) );
  XNOR U942 ( .A(b[1]), .B(n840), .Z(n842) );
  NANDN U943 ( .A(b[0]), .B(a[23]), .Z(n841) );
  NAND U944 ( .A(n842), .B(n841), .Z(n890) );
  NAND U945 ( .A(n2633), .B(n843), .Z(n845) );
  XOR U946 ( .A(b[5]), .B(a[20]), .Z(n884) );
  NANDN U947 ( .A(n37), .B(n884), .Z(n844) );
  AND U948 ( .A(n845), .B(n844), .Z(n888) );
  AND U949 ( .A(b[7]), .B(a[16]), .Z(n887) );
  XNOR U950 ( .A(n888), .B(n887), .Z(n889) );
  XNOR U951 ( .A(n890), .B(n889), .Z(n895) );
  XOR U952 ( .A(n896), .B(n895), .Z(n870) );
  NANDN U953 ( .A(n847), .B(n846), .Z(n851) );
  NANDN U954 ( .A(n849), .B(n848), .Z(n850) );
  AND U955 ( .A(n851), .B(n850), .Z(n869) );
  XNOR U956 ( .A(n870), .B(n869), .Z(n871) );
  NANDN U957 ( .A(n853), .B(n852), .Z(n857) );
  NAND U958 ( .A(n855), .B(n854), .Z(n856) );
  NAND U959 ( .A(n857), .B(n856), .Z(n872) );
  XNOR U960 ( .A(n871), .B(n872), .Z(n863) );
  XNOR U961 ( .A(n864), .B(n863), .Z(n865) );
  XNOR U962 ( .A(n866), .B(n865), .Z(n899) );
  XNOR U963 ( .A(sreg[80]), .B(n899), .Z(n901) );
  NANDN U964 ( .A(sreg[79]), .B(n858), .Z(n862) );
  NAND U965 ( .A(n860), .B(n859), .Z(n861) );
  NAND U966 ( .A(n862), .B(n861), .Z(n900) );
  XNOR U967 ( .A(n901), .B(n900), .Z(c[80]) );
  NANDN U968 ( .A(n864), .B(n863), .Z(n868) );
  NANDN U969 ( .A(n866), .B(n865), .Z(n867) );
  AND U970 ( .A(n868), .B(n867), .Z(n907) );
  NANDN U971 ( .A(n870), .B(n869), .Z(n874) );
  NANDN U972 ( .A(n872), .B(n871), .Z(n873) );
  AND U973 ( .A(n874), .B(n873), .Z(n905) );
  NANDN U974 ( .A(n2629), .B(n875), .Z(n877) );
  XOR U975 ( .A(b[7]), .B(a[19]), .Z(n916) );
  NANDN U976 ( .A(n2630), .B(n916), .Z(n876) );
  AND U977 ( .A(n877), .B(n876), .Z(n935) );
  NANDN U978 ( .A(n2483), .B(n878), .Z(n880) );
  XOR U979 ( .A(b[3]), .B(a[23]), .Z(n919) );
  NANDN U980 ( .A(n2484), .B(n919), .Z(n879) );
  NAND U981 ( .A(n880), .B(n879), .Z(n934) );
  XNOR U982 ( .A(n935), .B(n934), .Z(n937) );
  NAND U983 ( .A(b[0]), .B(a[25]), .Z(n881) );
  XNOR U984 ( .A(b[1]), .B(n881), .Z(n883) );
  NANDN U985 ( .A(b[0]), .B(a[24]), .Z(n882) );
  NAND U986 ( .A(n883), .B(n882), .Z(n931) );
  NAND U987 ( .A(n2633), .B(n884), .Z(n886) );
  XOR U988 ( .A(b[5]), .B(a[21]), .Z(n922) );
  NANDN U989 ( .A(n37), .B(n922), .Z(n885) );
  AND U990 ( .A(n886), .B(n885), .Z(n929) );
  AND U991 ( .A(b[7]), .B(a[17]), .Z(n928) );
  XNOR U992 ( .A(n929), .B(n928), .Z(n930) );
  XNOR U993 ( .A(n931), .B(n930), .Z(n936) );
  XOR U994 ( .A(n937), .B(n936), .Z(n911) );
  NANDN U995 ( .A(n888), .B(n887), .Z(n892) );
  NANDN U996 ( .A(n890), .B(n889), .Z(n891) );
  AND U997 ( .A(n892), .B(n891), .Z(n910) );
  XNOR U998 ( .A(n911), .B(n910), .Z(n912) );
  NANDN U999 ( .A(n894), .B(n893), .Z(n898) );
  NAND U1000 ( .A(n896), .B(n895), .Z(n897) );
  NAND U1001 ( .A(n898), .B(n897), .Z(n913) );
  XNOR U1002 ( .A(n912), .B(n913), .Z(n904) );
  XNOR U1003 ( .A(n905), .B(n904), .Z(n906) );
  XNOR U1004 ( .A(n907), .B(n906), .Z(n940) );
  XNOR U1005 ( .A(sreg[81]), .B(n940), .Z(n942) );
  NANDN U1006 ( .A(sreg[80]), .B(n899), .Z(n903) );
  NAND U1007 ( .A(n901), .B(n900), .Z(n902) );
  NAND U1008 ( .A(n903), .B(n902), .Z(n941) );
  XNOR U1009 ( .A(n942), .B(n941), .Z(c[81]) );
  NANDN U1010 ( .A(n905), .B(n904), .Z(n909) );
  NANDN U1011 ( .A(n907), .B(n906), .Z(n908) );
  AND U1012 ( .A(n909), .B(n908), .Z(n948) );
  NANDN U1013 ( .A(n911), .B(n910), .Z(n915) );
  NANDN U1014 ( .A(n913), .B(n912), .Z(n914) );
  AND U1015 ( .A(n915), .B(n914), .Z(n946) );
  NANDN U1016 ( .A(n2629), .B(n916), .Z(n918) );
  XOR U1017 ( .A(b[7]), .B(a[20]), .Z(n957) );
  NANDN U1018 ( .A(n2630), .B(n957), .Z(n917) );
  AND U1019 ( .A(n918), .B(n917), .Z(n976) );
  NANDN U1020 ( .A(n2483), .B(n919), .Z(n921) );
  XOR U1021 ( .A(b[3]), .B(a[24]), .Z(n960) );
  NANDN U1022 ( .A(n2484), .B(n960), .Z(n920) );
  NAND U1023 ( .A(n921), .B(n920), .Z(n975) );
  XNOR U1024 ( .A(n976), .B(n975), .Z(n978) );
  NAND U1025 ( .A(n2633), .B(n922), .Z(n924) );
  XOR U1026 ( .A(b[5]), .B(a[22]), .Z(n966) );
  NANDN U1027 ( .A(n37), .B(n966), .Z(n923) );
  AND U1028 ( .A(n924), .B(n923), .Z(n970) );
  AND U1029 ( .A(b[7]), .B(a[18]), .Z(n969) );
  XNOR U1030 ( .A(n970), .B(n969), .Z(n971) );
  NAND U1031 ( .A(b[0]), .B(a[26]), .Z(n925) );
  XNOR U1032 ( .A(b[1]), .B(n925), .Z(n927) );
  NANDN U1033 ( .A(b[0]), .B(a[25]), .Z(n926) );
  NAND U1034 ( .A(n927), .B(n926), .Z(n972) );
  XNOR U1035 ( .A(n971), .B(n972), .Z(n977) );
  XOR U1036 ( .A(n978), .B(n977), .Z(n952) );
  NANDN U1037 ( .A(n929), .B(n928), .Z(n933) );
  NANDN U1038 ( .A(n931), .B(n930), .Z(n932) );
  AND U1039 ( .A(n933), .B(n932), .Z(n951) );
  XNOR U1040 ( .A(n952), .B(n951), .Z(n953) );
  NANDN U1041 ( .A(n935), .B(n934), .Z(n939) );
  NAND U1042 ( .A(n937), .B(n936), .Z(n938) );
  NAND U1043 ( .A(n939), .B(n938), .Z(n954) );
  XNOR U1044 ( .A(n953), .B(n954), .Z(n945) );
  XNOR U1045 ( .A(n946), .B(n945), .Z(n947) );
  XNOR U1046 ( .A(n948), .B(n947), .Z(n981) );
  XNOR U1047 ( .A(sreg[82]), .B(n981), .Z(n983) );
  NANDN U1048 ( .A(sreg[81]), .B(n940), .Z(n944) );
  NAND U1049 ( .A(n942), .B(n941), .Z(n943) );
  NAND U1050 ( .A(n944), .B(n943), .Z(n982) );
  XNOR U1051 ( .A(n983), .B(n982), .Z(c[82]) );
  NANDN U1052 ( .A(n946), .B(n945), .Z(n950) );
  NANDN U1053 ( .A(n948), .B(n947), .Z(n949) );
  AND U1054 ( .A(n950), .B(n949), .Z(n989) );
  NANDN U1055 ( .A(n952), .B(n951), .Z(n956) );
  NANDN U1056 ( .A(n954), .B(n953), .Z(n955) );
  AND U1057 ( .A(n956), .B(n955), .Z(n987) );
  NANDN U1058 ( .A(n2629), .B(n957), .Z(n959) );
  XOR U1059 ( .A(b[7]), .B(a[21]), .Z(n998) );
  NANDN U1060 ( .A(n2630), .B(n998), .Z(n958) );
  AND U1061 ( .A(n959), .B(n958), .Z(n1017) );
  NANDN U1062 ( .A(n2483), .B(n960), .Z(n962) );
  XOR U1063 ( .A(b[3]), .B(a[25]), .Z(n1001) );
  NANDN U1064 ( .A(n2484), .B(n1001), .Z(n961) );
  NAND U1065 ( .A(n962), .B(n961), .Z(n1016) );
  XNOR U1066 ( .A(n1017), .B(n1016), .Z(n1019) );
  NAND U1067 ( .A(b[0]), .B(a[27]), .Z(n963) );
  XNOR U1068 ( .A(b[1]), .B(n963), .Z(n965) );
  NANDN U1069 ( .A(b[0]), .B(a[26]), .Z(n964) );
  NAND U1070 ( .A(n965), .B(n964), .Z(n1013) );
  NAND U1071 ( .A(n2633), .B(n966), .Z(n968) );
  XOR U1072 ( .A(b[5]), .B(a[23]), .Z(n1007) );
  NANDN U1073 ( .A(n37), .B(n1007), .Z(n967) );
  AND U1074 ( .A(n968), .B(n967), .Z(n1011) );
  AND U1075 ( .A(b[7]), .B(a[19]), .Z(n1010) );
  XNOR U1076 ( .A(n1011), .B(n1010), .Z(n1012) );
  XNOR U1077 ( .A(n1013), .B(n1012), .Z(n1018) );
  XOR U1078 ( .A(n1019), .B(n1018), .Z(n993) );
  NANDN U1079 ( .A(n970), .B(n969), .Z(n974) );
  NANDN U1080 ( .A(n972), .B(n971), .Z(n973) );
  AND U1081 ( .A(n974), .B(n973), .Z(n992) );
  XNOR U1082 ( .A(n993), .B(n992), .Z(n994) );
  NANDN U1083 ( .A(n976), .B(n975), .Z(n980) );
  NAND U1084 ( .A(n978), .B(n977), .Z(n979) );
  NAND U1085 ( .A(n980), .B(n979), .Z(n995) );
  XNOR U1086 ( .A(n994), .B(n995), .Z(n986) );
  XNOR U1087 ( .A(n987), .B(n986), .Z(n988) );
  XNOR U1088 ( .A(n989), .B(n988), .Z(n1022) );
  XNOR U1089 ( .A(sreg[83]), .B(n1022), .Z(n1024) );
  NANDN U1090 ( .A(sreg[82]), .B(n981), .Z(n985) );
  NAND U1091 ( .A(n983), .B(n982), .Z(n984) );
  NAND U1092 ( .A(n985), .B(n984), .Z(n1023) );
  XNOR U1093 ( .A(n1024), .B(n1023), .Z(c[83]) );
  NANDN U1094 ( .A(n987), .B(n986), .Z(n991) );
  NANDN U1095 ( .A(n989), .B(n988), .Z(n990) );
  AND U1096 ( .A(n991), .B(n990), .Z(n1030) );
  NANDN U1097 ( .A(n993), .B(n992), .Z(n997) );
  NANDN U1098 ( .A(n995), .B(n994), .Z(n996) );
  AND U1099 ( .A(n997), .B(n996), .Z(n1028) );
  NANDN U1100 ( .A(n2629), .B(n998), .Z(n1000) );
  XOR U1101 ( .A(b[7]), .B(a[22]), .Z(n1039) );
  NANDN U1102 ( .A(n2630), .B(n1039), .Z(n999) );
  AND U1103 ( .A(n1000), .B(n999), .Z(n1058) );
  NANDN U1104 ( .A(n2483), .B(n1001), .Z(n1003) );
  XOR U1105 ( .A(b[3]), .B(a[26]), .Z(n1042) );
  NANDN U1106 ( .A(n2484), .B(n1042), .Z(n1002) );
  NAND U1107 ( .A(n1003), .B(n1002), .Z(n1057) );
  XNOR U1108 ( .A(n1058), .B(n1057), .Z(n1060) );
  NAND U1109 ( .A(b[0]), .B(a[28]), .Z(n1004) );
  XNOR U1110 ( .A(b[1]), .B(n1004), .Z(n1006) );
  NANDN U1111 ( .A(b[0]), .B(a[27]), .Z(n1005) );
  NAND U1112 ( .A(n1006), .B(n1005), .Z(n1054) );
  NAND U1113 ( .A(n2633), .B(n1007), .Z(n1009) );
  XOR U1114 ( .A(b[5]), .B(a[24]), .Z(n1048) );
  NANDN U1115 ( .A(n37), .B(n1048), .Z(n1008) );
  AND U1116 ( .A(n1009), .B(n1008), .Z(n1052) );
  AND U1117 ( .A(b[7]), .B(a[20]), .Z(n1051) );
  XNOR U1118 ( .A(n1052), .B(n1051), .Z(n1053) );
  XNOR U1119 ( .A(n1054), .B(n1053), .Z(n1059) );
  XOR U1120 ( .A(n1060), .B(n1059), .Z(n1034) );
  NANDN U1121 ( .A(n1011), .B(n1010), .Z(n1015) );
  NANDN U1122 ( .A(n1013), .B(n1012), .Z(n1014) );
  AND U1123 ( .A(n1015), .B(n1014), .Z(n1033) );
  XNOR U1124 ( .A(n1034), .B(n1033), .Z(n1035) );
  NANDN U1125 ( .A(n1017), .B(n1016), .Z(n1021) );
  NAND U1126 ( .A(n1019), .B(n1018), .Z(n1020) );
  NAND U1127 ( .A(n1021), .B(n1020), .Z(n1036) );
  XNOR U1128 ( .A(n1035), .B(n1036), .Z(n1027) );
  XNOR U1129 ( .A(n1028), .B(n1027), .Z(n1029) );
  XNOR U1130 ( .A(n1030), .B(n1029), .Z(n1063) );
  XNOR U1131 ( .A(sreg[84]), .B(n1063), .Z(n1065) );
  NANDN U1132 ( .A(sreg[83]), .B(n1022), .Z(n1026) );
  NAND U1133 ( .A(n1024), .B(n1023), .Z(n1025) );
  NAND U1134 ( .A(n1026), .B(n1025), .Z(n1064) );
  XNOR U1135 ( .A(n1065), .B(n1064), .Z(c[84]) );
  NANDN U1136 ( .A(n1028), .B(n1027), .Z(n1032) );
  NANDN U1137 ( .A(n1030), .B(n1029), .Z(n1031) );
  AND U1138 ( .A(n1032), .B(n1031), .Z(n1071) );
  NANDN U1139 ( .A(n1034), .B(n1033), .Z(n1038) );
  NANDN U1140 ( .A(n1036), .B(n1035), .Z(n1037) );
  AND U1141 ( .A(n1038), .B(n1037), .Z(n1069) );
  NANDN U1142 ( .A(n2629), .B(n1039), .Z(n1041) );
  XOR U1143 ( .A(b[7]), .B(a[23]), .Z(n1080) );
  NANDN U1144 ( .A(n2630), .B(n1080), .Z(n1040) );
  AND U1145 ( .A(n1041), .B(n1040), .Z(n1099) );
  NANDN U1146 ( .A(n2483), .B(n1042), .Z(n1044) );
  XOR U1147 ( .A(b[3]), .B(a[27]), .Z(n1083) );
  NANDN U1148 ( .A(n2484), .B(n1083), .Z(n1043) );
  NAND U1149 ( .A(n1044), .B(n1043), .Z(n1098) );
  XNOR U1150 ( .A(n1099), .B(n1098), .Z(n1101) );
  NAND U1151 ( .A(b[0]), .B(a[29]), .Z(n1045) );
  XNOR U1152 ( .A(b[1]), .B(n1045), .Z(n1047) );
  NANDN U1153 ( .A(b[0]), .B(a[28]), .Z(n1046) );
  NAND U1154 ( .A(n1047), .B(n1046), .Z(n1095) );
  NAND U1155 ( .A(n2633), .B(n1048), .Z(n1050) );
  XOR U1156 ( .A(b[5]), .B(a[25]), .Z(n1086) );
  NANDN U1157 ( .A(n37), .B(n1086), .Z(n1049) );
  AND U1158 ( .A(n1050), .B(n1049), .Z(n1093) );
  AND U1159 ( .A(b[7]), .B(a[21]), .Z(n1092) );
  XNOR U1160 ( .A(n1093), .B(n1092), .Z(n1094) );
  XNOR U1161 ( .A(n1095), .B(n1094), .Z(n1100) );
  XOR U1162 ( .A(n1101), .B(n1100), .Z(n1075) );
  NANDN U1163 ( .A(n1052), .B(n1051), .Z(n1056) );
  NANDN U1164 ( .A(n1054), .B(n1053), .Z(n1055) );
  AND U1165 ( .A(n1056), .B(n1055), .Z(n1074) );
  XNOR U1166 ( .A(n1075), .B(n1074), .Z(n1076) );
  NANDN U1167 ( .A(n1058), .B(n1057), .Z(n1062) );
  NAND U1168 ( .A(n1060), .B(n1059), .Z(n1061) );
  NAND U1169 ( .A(n1062), .B(n1061), .Z(n1077) );
  XNOR U1170 ( .A(n1076), .B(n1077), .Z(n1068) );
  XNOR U1171 ( .A(n1069), .B(n1068), .Z(n1070) );
  XNOR U1172 ( .A(n1071), .B(n1070), .Z(n1104) );
  XNOR U1173 ( .A(sreg[85]), .B(n1104), .Z(n1106) );
  NANDN U1174 ( .A(sreg[84]), .B(n1063), .Z(n1067) );
  NAND U1175 ( .A(n1065), .B(n1064), .Z(n1066) );
  NAND U1176 ( .A(n1067), .B(n1066), .Z(n1105) );
  XNOR U1177 ( .A(n1106), .B(n1105), .Z(c[85]) );
  NANDN U1178 ( .A(n1069), .B(n1068), .Z(n1073) );
  NANDN U1179 ( .A(n1071), .B(n1070), .Z(n1072) );
  AND U1180 ( .A(n1073), .B(n1072), .Z(n1112) );
  NANDN U1181 ( .A(n1075), .B(n1074), .Z(n1079) );
  NANDN U1182 ( .A(n1077), .B(n1076), .Z(n1078) );
  AND U1183 ( .A(n1079), .B(n1078), .Z(n1110) );
  NANDN U1184 ( .A(n2629), .B(n1080), .Z(n1082) );
  XOR U1185 ( .A(b[7]), .B(a[24]), .Z(n1121) );
  NANDN U1186 ( .A(n2630), .B(n1121), .Z(n1081) );
  AND U1187 ( .A(n1082), .B(n1081), .Z(n1140) );
  NANDN U1188 ( .A(n2483), .B(n1083), .Z(n1085) );
  XOR U1189 ( .A(b[3]), .B(a[28]), .Z(n1124) );
  NANDN U1190 ( .A(n2484), .B(n1124), .Z(n1084) );
  NAND U1191 ( .A(n1085), .B(n1084), .Z(n1139) );
  XNOR U1192 ( .A(n1140), .B(n1139), .Z(n1142) );
  NAND U1193 ( .A(n2633), .B(n1086), .Z(n1088) );
  XOR U1194 ( .A(b[5]), .B(a[26]), .Z(n1130) );
  NANDN U1195 ( .A(n37), .B(n1130), .Z(n1087) );
  AND U1196 ( .A(n1088), .B(n1087), .Z(n1134) );
  AND U1197 ( .A(b[7]), .B(a[22]), .Z(n1133) );
  XNOR U1198 ( .A(n1134), .B(n1133), .Z(n1135) );
  NAND U1199 ( .A(b[0]), .B(a[30]), .Z(n1089) );
  XNOR U1200 ( .A(b[1]), .B(n1089), .Z(n1091) );
  NANDN U1201 ( .A(b[0]), .B(a[29]), .Z(n1090) );
  NAND U1202 ( .A(n1091), .B(n1090), .Z(n1136) );
  XNOR U1203 ( .A(n1135), .B(n1136), .Z(n1141) );
  XOR U1204 ( .A(n1142), .B(n1141), .Z(n1116) );
  NANDN U1205 ( .A(n1093), .B(n1092), .Z(n1097) );
  NANDN U1206 ( .A(n1095), .B(n1094), .Z(n1096) );
  AND U1207 ( .A(n1097), .B(n1096), .Z(n1115) );
  XNOR U1208 ( .A(n1116), .B(n1115), .Z(n1117) );
  NANDN U1209 ( .A(n1099), .B(n1098), .Z(n1103) );
  NAND U1210 ( .A(n1101), .B(n1100), .Z(n1102) );
  NAND U1211 ( .A(n1103), .B(n1102), .Z(n1118) );
  XNOR U1212 ( .A(n1117), .B(n1118), .Z(n1109) );
  XNOR U1213 ( .A(n1110), .B(n1109), .Z(n1111) );
  XNOR U1214 ( .A(n1112), .B(n1111), .Z(n1145) );
  XNOR U1215 ( .A(sreg[86]), .B(n1145), .Z(n1147) );
  NANDN U1216 ( .A(sreg[85]), .B(n1104), .Z(n1108) );
  NAND U1217 ( .A(n1106), .B(n1105), .Z(n1107) );
  NAND U1218 ( .A(n1108), .B(n1107), .Z(n1146) );
  XNOR U1219 ( .A(n1147), .B(n1146), .Z(c[86]) );
  NANDN U1220 ( .A(n1110), .B(n1109), .Z(n1114) );
  NANDN U1221 ( .A(n1112), .B(n1111), .Z(n1113) );
  AND U1222 ( .A(n1114), .B(n1113), .Z(n1153) );
  NANDN U1223 ( .A(n1116), .B(n1115), .Z(n1120) );
  NANDN U1224 ( .A(n1118), .B(n1117), .Z(n1119) );
  AND U1225 ( .A(n1120), .B(n1119), .Z(n1151) );
  NANDN U1226 ( .A(n2629), .B(n1121), .Z(n1123) );
  XOR U1227 ( .A(b[7]), .B(a[25]), .Z(n1162) );
  NANDN U1228 ( .A(n2630), .B(n1162), .Z(n1122) );
  AND U1229 ( .A(n1123), .B(n1122), .Z(n1181) );
  NANDN U1230 ( .A(n2483), .B(n1124), .Z(n1126) );
  XOR U1231 ( .A(b[3]), .B(a[29]), .Z(n1165) );
  NANDN U1232 ( .A(n2484), .B(n1165), .Z(n1125) );
  NAND U1233 ( .A(n1126), .B(n1125), .Z(n1180) );
  XNOR U1234 ( .A(n1181), .B(n1180), .Z(n1183) );
  NAND U1235 ( .A(b[0]), .B(a[31]), .Z(n1127) );
  XNOR U1236 ( .A(b[1]), .B(n1127), .Z(n1129) );
  NANDN U1237 ( .A(b[0]), .B(a[30]), .Z(n1128) );
  NAND U1238 ( .A(n1129), .B(n1128), .Z(n1177) );
  NAND U1239 ( .A(n2633), .B(n1130), .Z(n1132) );
  XOR U1240 ( .A(b[5]), .B(a[27]), .Z(n1168) );
  NANDN U1241 ( .A(n37), .B(n1168), .Z(n1131) );
  AND U1242 ( .A(n1132), .B(n1131), .Z(n1175) );
  AND U1243 ( .A(b[7]), .B(a[23]), .Z(n1174) );
  XNOR U1244 ( .A(n1175), .B(n1174), .Z(n1176) );
  XNOR U1245 ( .A(n1177), .B(n1176), .Z(n1182) );
  XOR U1246 ( .A(n1183), .B(n1182), .Z(n1157) );
  NANDN U1247 ( .A(n1134), .B(n1133), .Z(n1138) );
  NANDN U1248 ( .A(n1136), .B(n1135), .Z(n1137) );
  AND U1249 ( .A(n1138), .B(n1137), .Z(n1156) );
  XNOR U1250 ( .A(n1157), .B(n1156), .Z(n1158) );
  NANDN U1251 ( .A(n1140), .B(n1139), .Z(n1144) );
  NAND U1252 ( .A(n1142), .B(n1141), .Z(n1143) );
  NAND U1253 ( .A(n1144), .B(n1143), .Z(n1159) );
  XNOR U1254 ( .A(n1158), .B(n1159), .Z(n1150) );
  XNOR U1255 ( .A(n1151), .B(n1150), .Z(n1152) );
  XNOR U1256 ( .A(n1153), .B(n1152), .Z(n1186) );
  XNOR U1257 ( .A(sreg[87]), .B(n1186), .Z(n1188) );
  NANDN U1258 ( .A(sreg[86]), .B(n1145), .Z(n1149) );
  NAND U1259 ( .A(n1147), .B(n1146), .Z(n1148) );
  NAND U1260 ( .A(n1149), .B(n1148), .Z(n1187) );
  XNOR U1261 ( .A(n1188), .B(n1187), .Z(c[87]) );
  NANDN U1262 ( .A(n1151), .B(n1150), .Z(n1155) );
  NANDN U1263 ( .A(n1153), .B(n1152), .Z(n1154) );
  AND U1264 ( .A(n1155), .B(n1154), .Z(n1194) );
  NANDN U1265 ( .A(n1157), .B(n1156), .Z(n1161) );
  NANDN U1266 ( .A(n1159), .B(n1158), .Z(n1160) );
  AND U1267 ( .A(n1161), .B(n1160), .Z(n1192) );
  NANDN U1268 ( .A(n2629), .B(n1162), .Z(n1164) );
  XOR U1269 ( .A(b[7]), .B(a[26]), .Z(n1203) );
  NANDN U1270 ( .A(n2630), .B(n1203), .Z(n1163) );
  AND U1271 ( .A(n1164), .B(n1163), .Z(n1222) );
  NANDN U1272 ( .A(n2483), .B(n1165), .Z(n1167) );
  XOR U1273 ( .A(b[3]), .B(a[30]), .Z(n1206) );
  NANDN U1274 ( .A(n2484), .B(n1206), .Z(n1166) );
  NAND U1275 ( .A(n1167), .B(n1166), .Z(n1221) );
  XNOR U1276 ( .A(n1222), .B(n1221), .Z(n1224) );
  NAND U1277 ( .A(n2633), .B(n1168), .Z(n1170) );
  XOR U1278 ( .A(b[5]), .B(a[28]), .Z(n1212) );
  NANDN U1279 ( .A(n37), .B(n1212), .Z(n1169) );
  AND U1280 ( .A(n1170), .B(n1169), .Z(n1216) );
  AND U1281 ( .A(b[7]), .B(a[24]), .Z(n1215) );
  XNOR U1282 ( .A(n1216), .B(n1215), .Z(n1217) );
  NAND U1283 ( .A(b[0]), .B(a[32]), .Z(n1171) );
  XNOR U1284 ( .A(b[1]), .B(n1171), .Z(n1173) );
  NANDN U1285 ( .A(b[0]), .B(a[31]), .Z(n1172) );
  NAND U1286 ( .A(n1173), .B(n1172), .Z(n1218) );
  XNOR U1287 ( .A(n1217), .B(n1218), .Z(n1223) );
  XOR U1288 ( .A(n1224), .B(n1223), .Z(n1198) );
  NANDN U1289 ( .A(n1175), .B(n1174), .Z(n1179) );
  NANDN U1290 ( .A(n1177), .B(n1176), .Z(n1178) );
  AND U1291 ( .A(n1179), .B(n1178), .Z(n1197) );
  XNOR U1292 ( .A(n1198), .B(n1197), .Z(n1199) );
  NANDN U1293 ( .A(n1181), .B(n1180), .Z(n1185) );
  NAND U1294 ( .A(n1183), .B(n1182), .Z(n1184) );
  NAND U1295 ( .A(n1185), .B(n1184), .Z(n1200) );
  XNOR U1296 ( .A(n1199), .B(n1200), .Z(n1191) );
  XNOR U1297 ( .A(n1192), .B(n1191), .Z(n1193) );
  XNOR U1298 ( .A(n1194), .B(n1193), .Z(n1227) );
  XNOR U1299 ( .A(sreg[88]), .B(n1227), .Z(n1229) );
  NANDN U1300 ( .A(sreg[87]), .B(n1186), .Z(n1190) );
  NAND U1301 ( .A(n1188), .B(n1187), .Z(n1189) );
  NAND U1302 ( .A(n1190), .B(n1189), .Z(n1228) );
  XNOR U1303 ( .A(n1229), .B(n1228), .Z(c[88]) );
  NANDN U1304 ( .A(n1192), .B(n1191), .Z(n1196) );
  NANDN U1305 ( .A(n1194), .B(n1193), .Z(n1195) );
  AND U1306 ( .A(n1196), .B(n1195), .Z(n1235) );
  NANDN U1307 ( .A(n1198), .B(n1197), .Z(n1202) );
  NANDN U1308 ( .A(n1200), .B(n1199), .Z(n1201) );
  AND U1309 ( .A(n1202), .B(n1201), .Z(n1233) );
  NANDN U1310 ( .A(n2629), .B(n1203), .Z(n1205) );
  XOR U1311 ( .A(b[7]), .B(a[27]), .Z(n1244) );
  NANDN U1312 ( .A(n2630), .B(n1244), .Z(n1204) );
  AND U1313 ( .A(n1205), .B(n1204), .Z(n1263) );
  NANDN U1314 ( .A(n2483), .B(n1206), .Z(n1208) );
  XOR U1315 ( .A(b[3]), .B(a[31]), .Z(n1247) );
  NANDN U1316 ( .A(n2484), .B(n1247), .Z(n1207) );
  NAND U1317 ( .A(n1208), .B(n1207), .Z(n1262) );
  XNOR U1318 ( .A(n1263), .B(n1262), .Z(n1265) );
  NAND U1319 ( .A(b[0]), .B(a[33]), .Z(n1209) );
  XNOR U1320 ( .A(b[1]), .B(n1209), .Z(n1211) );
  NANDN U1321 ( .A(b[0]), .B(a[32]), .Z(n1210) );
  NAND U1322 ( .A(n1211), .B(n1210), .Z(n1259) );
  NAND U1323 ( .A(n2633), .B(n1212), .Z(n1214) );
  XOR U1324 ( .A(b[5]), .B(a[29]), .Z(n1253) );
  NANDN U1325 ( .A(n37), .B(n1253), .Z(n1213) );
  AND U1326 ( .A(n1214), .B(n1213), .Z(n1257) );
  AND U1327 ( .A(b[7]), .B(a[25]), .Z(n1256) );
  XNOR U1328 ( .A(n1257), .B(n1256), .Z(n1258) );
  XNOR U1329 ( .A(n1259), .B(n1258), .Z(n1264) );
  XOR U1330 ( .A(n1265), .B(n1264), .Z(n1239) );
  NANDN U1331 ( .A(n1216), .B(n1215), .Z(n1220) );
  NANDN U1332 ( .A(n1218), .B(n1217), .Z(n1219) );
  AND U1333 ( .A(n1220), .B(n1219), .Z(n1238) );
  XNOR U1334 ( .A(n1239), .B(n1238), .Z(n1240) );
  NANDN U1335 ( .A(n1222), .B(n1221), .Z(n1226) );
  NAND U1336 ( .A(n1224), .B(n1223), .Z(n1225) );
  NAND U1337 ( .A(n1226), .B(n1225), .Z(n1241) );
  XNOR U1338 ( .A(n1240), .B(n1241), .Z(n1232) );
  XNOR U1339 ( .A(n1233), .B(n1232), .Z(n1234) );
  XNOR U1340 ( .A(n1235), .B(n1234), .Z(n1268) );
  XNOR U1341 ( .A(sreg[89]), .B(n1268), .Z(n1270) );
  NANDN U1342 ( .A(sreg[88]), .B(n1227), .Z(n1231) );
  NAND U1343 ( .A(n1229), .B(n1228), .Z(n1230) );
  NAND U1344 ( .A(n1231), .B(n1230), .Z(n1269) );
  XNOR U1345 ( .A(n1270), .B(n1269), .Z(c[89]) );
  NANDN U1346 ( .A(n1233), .B(n1232), .Z(n1237) );
  NANDN U1347 ( .A(n1235), .B(n1234), .Z(n1236) );
  AND U1348 ( .A(n1237), .B(n1236), .Z(n1276) );
  NANDN U1349 ( .A(n1239), .B(n1238), .Z(n1243) );
  NANDN U1350 ( .A(n1241), .B(n1240), .Z(n1242) );
  AND U1351 ( .A(n1243), .B(n1242), .Z(n1274) );
  NANDN U1352 ( .A(n2629), .B(n1244), .Z(n1246) );
  XOR U1353 ( .A(b[7]), .B(a[28]), .Z(n1285) );
  NANDN U1354 ( .A(n2630), .B(n1285), .Z(n1245) );
  AND U1355 ( .A(n1246), .B(n1245), .Z(n1304) );
  NANDN U1356 ( .A(n2483), .B(n1247), .Z(n1249) );
  XOR U1357 ( .A(b[3]), .B(a[32]), .Z(n1288) );
  NANDN U1358 ( .A(n2484), .B(n1288), .Z(n1248) );
  NAND U1359 ( .A(n1249), .B(n1248), .Z(n1303) );
  XNOR U1360 ( .A(n1304), .B(n1303), .Z(n1306) );
  NAND U1361 ( .A(b[0]), .B(a[34]), .Z(n1250) );
  XNOR U1362 ( .A(b[1]), .B(n1250), .Z(n1252) );
  NANDN U1363 ( .A(b[0]), .B(a[33]), .Z(n1251) );
  NAND U1364 ( .A(n1252), .B(n1251), .Z(n1300) );
  NAND U1365 ( .A(n2633), .B(n1253), .Z(n1255) );
  XOR U1366 ( .A(b[5]), .B(a[30]), .Z(n1294) );
  NANDN U1367 ( .A(n37), .B(n1294), .Z(n1254) );
  AND U1368 ( .A(n1255), .B(n1254), .Z(n1298) );
  AND U1369 ( .A(b[7]), .B(a[26]), .Z(n1297) );
  XNOR U1370 ( .A(n1298), .B(n1297), .Z(n1299) );
  XNOR U1371 ( .A(n1300), .B(n1299), .Z(n1305) );
  XOR U1372 ( .A(n1306), .B(n1305), .Z(n1280) );
  NANDN U1373 ( .A(n1257), .B(n1256), .Z(n1261) );
  NANDN U1374 ( .A(n1259), .B(n1258), .Z(n1260) );
  AND U1375 ( .A(n1261), .B(n1260), .Z(n1279) );
  XNOR U1376 ( .A(n1280), .B(n1279), .Z(n1281) );
  NANDN U1377 ( .A(n1263), .B(n1262), .Z(n1267) );
  NAND U1378 ( .A(n1265), .B(n1264), .Z(n1266) );
  NAND U1379 ( .A(n1267), .B(n1266), .Z(n1282) );
  XNOR U1380 ( .A(n1281), .B(n1282), .Z(n1273) );
  XNOR U1381 ( .A(n1274), .B(n1273), .Z(n1275) );
  XNOR U1382 ( .A(n1276), .B(n1275), .Z(n1309) );
  XNOR U1383 ( .A(sreg[90]), .B(n1309), .Z(n1311) );
  NANDN U1384 ( .A(sreg[89]), .B(n1268), .Z(n1272) );
  NAND U1385 ( .A(n1270), .B(n1269), .Z(n1271) );
  NAND U1386 ( .A(n1272), .B(n1271), .Z(n1310) );
  XNOR U1387 ( .A(n1311), .B(n1310), .Z(c[90]) );
  NANDN U1388 ( .A(n1274), .B(n1273), .Z(n1278) );
  NANDN U1389 ( .A(n1276), .B(n1275), .Z(n1277) );
  AND U1390 ( .A(n1278), .B(n1277), .Z(n1317) );
  NANDN U1391 ( .A(n1280), .B(n1279), .Z(n1284) );
  NANDN U1392 ( .A(n1282), .B(n1281), .Z(n1283) );
  AND U1393 ( .A(n1284), .B(n1283), .Z(n1315) );
  NANDN U1394 ( .A(n2629), .B(n1285), .Z(n1287) );
  XOR U1395 ( .A(b[7]), .B(a[29]), .Z(n1326) );
  NANDN U1396 ( .A(n2630), .B(n1326), .Z(n1286) );
  AND U1397 ( .A(n1287), .B(n1286), .Z(n1345) );
  NANDN U1398 ( .A(n2483), .B(n1288), .Z(n1290) );
  XOR U1399 ( .A(b[3]), .B(a[33]), .Z(n1329) );
  NANDN U1400 ( .A(n2484), .B(n1329), .Z(n1289) );
  NAND U1401 ( .A(n1290), .B(n1289), .Z(n1344) );
  XNOR U1402 ( .A(n1345), .B(n1344), .Z(n1347) );
  NAND U1403 ( .A(b[0]), .B(a[35]), .Z(n1291) );
  XNOR U1404 ( .A(b[1]), .B(n1291), .Z(n1293) );
  NANDN U1405 ( .A(b[0]), .B(a[34]), .Z(n1292) );
  NAND U1406 ( .A(n1293), .B(n1292), .Z(n1341) );
  NAND U1407 ( .A(n2633), .B(n1294), .Z(n1296) );
  XOR U1408 ( .A(b[5]), .B(a[31]), .Z(n1335) );
  NANDN U1409 ( .A(n37), .B(n1335), .Z(n1295) );
  AND U1410 ( .A(n1296), .B(n1295), .Z(n1339) );
  AND U1411 ( .A(b[7]), .B(a[27]), .Z(n1338) );
  XNOR U1412 ( .A(n1339), .B(n1338), .Z(n1340) );
  XNOR U1413 ( .A(n1341), .B(n1340), .Z(n1346) );
  XOR U1414 ( .A(n1347), .B(n1346), .Z(n1321) );
  NANDN U1415 ( .A(n1298), .B(n1297), .Z(n1302) );
  NANDN U1416 ( .A(n1300), .B(n1299), .Z(n1301) );
  AND U1417 ( .A(n1302), .B(n1301), .Z(n1320) );
  XNOR U1418 ( .A(n1321), .B(n1320), .Z(n1322) );
  NANDN U1419 ( .A(n1304), .B(n1303), .Z(n1308) );
  NAND U1420 ( .A(n1306), .B(n1305), .Z(n1307) );
  NAND U1421 ( .A(n1308), .B(n1307), .Z(n1323) );
  XNOR U1422 ( .A(n1322), .B(n1323), .Z(n1314) );
  XNOR U1423 ( .A(n1315), .B(n1314), .Z(n1316) );
  XNOR U1424 ( .A(n1317), .B(n1316), .Z(n1350) );
  XNOR U1425 ( .A(sreg[91]), .B(n1350), .Z(n1352) );
  NANDN U1426 ( .A(sreg[90]), .B(n1309), .Z(n1313) );
  NAND U1427 ( .A(n1311), .B(n1310), .Z(n1312) );
  NAND U1428 ( .A(n1313), .B(n1312), .Z(n1351) );
  XNOR U1429 ( .A(n1352), .B(n1351), .Z(c[91]) );
  NANDN U1430 ( .A(n1315), .B(n1314), .Z(n1319) );
  NANDN U1431 ( .A(n1317), .B(n1316), .Z(n1318) );
  AND U1432 ( .A(n1319), .B(n1318), .Z(n1358) );
  NANDN U1433 ( .A(n1321), .B(n1320), .Z(n1325) );
  NANDN U1434 ( .A(n1323), .B(n1322), .Z(n1324) );
  AND U1435 ( .A(n1325), .B(n1324), .Z(n1356) );
  NANDN U1436 ( .A(n2629), .B(n1326), .Z(n1328) );
  XOR U1437 ( .A(b[7]), .B(a[30]), .Z(n1367) );
  NANDN U1438 ( .A(n2630), .B(n1367), .Z(n1327) );
  AND U1439 ( .A(n1328), .B(n1327), .Z(n1386) );
  NANDN U1440 ( .A(n2483), .B(n1329), .Z(n1331) );
  XOR U1441 ( .A(b[3]), .B(a[34]), .Z(n1370) );
  NANDN U1442 ( .A(n2484), .B(n1370), .Z(n1330) );
  NAND U1443 ( .A(n1331), .B(n1330), .Z(n1385) );
  XNOR U1444 ( .A(n1386), .B(n1385), .Z(n1388) );
  NAND U1445 ( .A(b[0]), .B(a[36]), .Z(n1332) );
  XNOR U1446 ( .A(b[1]), .B(n1332), .Z(n1334) );
  NANDN U1447 ( .A(b[0]), .B(a[35]), .Z(n1333) );
  NAND U1448 ( .A(n1334), .B(n1333), .Z(n1382) );
  NAND U1449 ( .A(n2633), .B(n1335), .Z(n1337) );
  XOR U1450 ( .A(b[5]), .B(a[32]), .Z(n1376) );
  NANDN U1451 ( .A(n37), .B(n1376), .Z(n1336) );
  AND U1452 ( .A(n1337), .B(n1336), .Z(n1380) );
  AND U1453 ( .A(b[7]), .B(a[28]), .Z(n1379) );
  XNOR U1454 ( .A(n1380), .B(n1379), .Z(n1381) );
  XNOR U1455 ( .A(n1382), .B(n1381), .Z(n1387) );
  XOR U1456 ( .A(n1388), .B(n1387), .Z(n1362) );
  NANDN U1457 ( .A(n1339), .B(n1338), .Z(n1343) );
  NANDN U1458 ( .A(n1341), .B(n1340), .Z(n1342) );
  AND U1459 ( .A(n1343), .B(n1342), .Z(n1361) );
  XNOR U1460 ( .A(n1362), .B(n1361), .Z(n1363) );
  NANDN U1461 ( .A(n1345), .B(n1344), .Z(n1349) );
  NAND U1462 ( .A(n1347), .B(n1346), .Z(n1348) );
  NAND U1463 ( .A(n1349), .B(n1348), .Z(n1364) );
  XNOR U1464 ( .A(n1363), .B(n1364), .Z(n1355) );
  XNOR U1465 ( .A(n1356), .B(n1355), .Z(n1357) );
  XNOR U1466 ( .A(n1358), .B(n1357), .Z(n1391) );
  XNOR U1467 ( .A(sreg[92]), .B(n1391), .Z(n1393) );
  NANDN U1468 ( .A(sreg[91]), .B(n1350), .Z(n1354) );
  NAND U1469 ( .A(n1352), .B(n1351), .Z(n1353) );
  NAND U1470 ( .A(n1354), .B(n1353), .Z(n1392) );
  XNOR U1471 ( .A(n1393), .B(n1392), .Z(c[92]) );
  NANDN U1472 ( .A(n1356), .B(n1355), .Z(n1360) );
  NANDN U1473 ( .A(n1358), .B(n1357), .Z(n1359) );
  AND U1474 ( .A(n1360), .B(n1359), .Z(n1399) );
  NANDN U1475 ( .A(n1362), .B(n1361), .Z(n1366) );
  NANDN U1476 ( .A(n1364), .B(n1363), .Z(n1365) );
  AND U1477 ( .A(n1366), .B(n1365), .Z(n1397) );
  NANDN U1478 ( .A(n2629), .B(n1367), .Z(n1369) );
  XOR U1479 ( .A(b[7]), .B(a[31]), .Z(n1408) );
  NANDN U1480 ( .A(n2630), .B(n1408), .Z(n1368) );
  AND U1481 ( .A(n1369), .B(n1368), .Z(n1427) );
  NANDN U1482 ( .A(n2483), .B(n1370), .Z(n1372) );
  XOR U1483 ( .A(b[3]), .B(a[35]), .Z(n1411) );
  NANDN U1484 ( .A(n2484), .B(n1411), .Z(n1371) );
  NAND U1485 ( .A(n1372), .B(n1371), .Z(n1426) );
  XNOR U1486 ( .A(n1427), .B(n1426), .Z(n1429) );
  NAND U1487 ( .A(b[0]), .B(a[37]), .Z(n1373) );
  XNOR U1488 ( .A(b[1]), .B(n1373), .Z(n1375) );
  NANDN U1489 ( .A(b[0]), .B(a[36]), .Z(n1374) );
  NAND U1490 ( .A(n1375), .B(n1374), .Z(n1423) );
  NAND U1491 ( .A(n2633), .B(n1376), .Z(n1378) );
  XOR U1492 ( .A(b[5]), .B(a[33]), .Z(n1417) );
  NANDN U1493 ( .A(n37), .B(n1417), .Z(n1377) );
  AND U1494 ( .A(n1378), .B(n1377), .Z(n1421) );
  AND U1495 ( .A(b[7]), .B(a[29]), .Z(n1420) );
  XNOR U1496 ( .A(n1421), .B(n1420), .Z(n1422) );
  XNOR U1497 ( .A(n1423), .B(n1422), .Z(n1428) );
  XOR U1498 ( .A(n1429), .B(n1428), .Z(n1403) );
  NANDN U1499 ( .A(n1380), .B(n1379), .Z(n1384) );
  NANDN U1500 ( .A(n1382), .B(n1381), .Z(n1383) );
  AND U1501 ( .A(n1384), .B(n1383), .Z(n1402) );
  XNOR U1502 ( .A(n1403), .B(n1402), .Z(n1404) );
  NANDN U1503 ( .A(n1386), .B(n1385), .Z(n1390) );
  NAND U1504 ( .A(n1388), .B(n1387), .Z(n1389) );
  NAND U1505 ( .A(n1390), .B(n1389), .Z(n1405) );
  XNOR U1506 ( .A(n1404), .B(n1405), .Z(n1396) );
  XNOR U1507 ( .A(n1397), .B(n1396), .Z(n1398) );
  XNOR U1508 ( .A(n1399), .B(n1398), .Z(n1432) );
  XNOR U1509 ( .A(sreg[93]), .B(n1432), .Z(n1434) );
  NANDN U1510 ( .A(sreg[92]), .B(n1391), .Z(n1395) );
  NAND U1511 ( .A(n1393), .B(n1392), .Z(n1394) );
  NAND U1512 ( .A(n1395), .B(n1394), .Z(n1433) );
  XNOR U1513 ( .A(n1434), .B(n1433), .Z(c[93]) );
  NANDN U1514 ( .A(n1397), .B(n1396), .Z(n1401) );
  NANDN U1515 ( .A(n1399), .B(n1398), .Z(n1400) );
  AND U1516 ( .A(n1401), .B(n1400), .Z(n1440) );
  NANDN U1517 ( .A(n1403), .B(n1402), .Z(n1407) );
  NANDN U1518 ( .A(n1405), .B(n1404), .Z(n1406) );
  AND U1519 ( .A(n1407), .B(n1406), .Z(n1438) );
  NANDN U1520 ( .A(n2629), .B(n1408), .Z(n1410) );
  XOR U1521 ( .A(b[7]), .B(a[32]), .Z(n1449) );
  NANDN U1522 ( .A(n2630), .B(n1449), .Z(n1409) );
  AND U1523 ( .A(n1410), .B(n1409), .Z(n1468) );
  NANDN U1524 ( .A(n2483), .B(n1411), .Z(n1413) );
  XOR U1525 ( .A(b[3]), .B(a[36]), .Z(n1452) );
  NANDN U1526 ( .A(n2484), .B(n1452), .Z(n1412) );
  NAND U1527 ( .A(n1413), .B(n1412), .Z(n1467) );
  XNOR U1528 ( .A(n1468), .B(n1467), .Z(n1470) );
  NAND U1529 ( .A(b[0]), .B(a[38]), .Z(n1414) );
  XNOR U1530 ( .A(b[1]), .B(n1414), .Z(n1416) );
  NANDN U1531 ( .A(b[0]), .B(a[37]), .Z(n1415) );
  NAND U1532 ( .A(n1416), .B(n1415), .Z(n1464) );
  NAND U1533 ( .A(n2633), .B(n1417), .Z(n1419) );
  XOR U1534 ( .A(b[5]), .B(a[34]), .Z(n1458) );
  NANDN U1535 ( .A(n37), .B(n1458), .Z(n1418) );
  AND U1536 ( .A(n1419), .B(n1418), .Z(n1462) );
  AND U1537 ( .A(b[7]), .B(a[30]), .Z(n1461) );
  XNOR U1538 ( .A(n1462), .B(n1461), .Z(n1463) );
  XNOR U1539 ( .A(n1464), .B(n1463), .Z(n1469) );
  XOR U1540 ( .A(n1470), .B(n1469), .Z(n1444) );
  NANDN U1541 ( .A(n1421), .B(n1420), .Z(n1425) );
  NANDN U1542 ( .A(n1423), .B(n1422), .Z(n1424) );
  AND U1543 ( .A(n1425), .B(n1424), .Z(n1443) );
  XNOR U1544 ( .A(n1444), .B(n1443), .Z(n1445) );
  NANDN U1545 ( .A(n1427), .B(n1426), .Z(n1431) );
  NAND U1546 ( .A(n1429), .B(n1428), .Z(n1430) );
  NAND U1547 ( .A(n1431), .B(n1430), .Z(n1446) );
  XNOR U1548 ( .A(n1445), .B(n1446), .Z(n1437) );
  XNOR U1549 ( .A(n1438), .B(n1437), .Z(n1439) );
  XNOR U1550 ( .A(n1440), .B(n1439), .Z(n1473) );
  XNOR U1551 ( .A(sreg[94]), .B(n1473), .Z(n1475) );
  NANDN U1552 ( .A(sreg[93]), .B(n1432), .Z(n1436) );
  NAND U1553 ( .A(n1434), .B(n1433), .Z(n1435) );
  NAND U1554 ( .A(n1436), .B(n1435), .Z(n1474) );
  XNOR U1555 ( .A(n1475), .B(n1474), .Z(c[94]) );
  NANDN U1556 ( .A(n1438), .B(n1437), .Z(n1442) );
  NANDN U1557 ( .A(n1440), .B(n1439), .Z(n1441) );
  AND U1558 ( .A(n1442), .B(n1441), .Z(n1481) );
  NANDN U1559 ( .A(n1444), .B(n1443), .Z(n1448) );
  NANDN U1560 ( .A(n1446), .B(n1445), .Z(n1447) );
  AND U1561 ( .A(n1448), .B(n1447), .Z(n1479) );
  NANDN U1562 ( .A(n2629), .B(n1449), .Z(n1451) );
  XOR U1563 ( .A(b[7]), .B(a[33]), .Z(n1490) );
  NANDN U1564 ( .A(n2630), .B(n1490), .Z(n1450) );
  AND U1565 ( .A(n1451), .B(n1450), .Z(n1509) );
  NANDN U1566 ( .A(n2483), .B(n1452), .Z(n1454) );
  XOR U1567 ( .A(b[3]), .B(a[37]), .Z(n1493) );
  NANDN U1568 ( .A(n2484), .B(n1493), .Z(n1453) );
  NAND U1569 ( .A(n1454), .B(n1453), .Z(n1508) );
  XNOR U1570 ( .A(n1509), .B(n1508), .Z(n1511) );
  NAND U1571 ( .A(b[0]), .B(a[39]), .Z(n1455) );
  XNOR U1572 ( .A(b[1]), .B(n1455), .Z(n1457) );
  NANDN U1573 ( .A(b[0]), .B(a[38]), .Z(n1456) );
  NAND U1574 ( .A(n1457), .B(n1456), .Z(n1505) );
  NAND U1575 ( .A(n2633), .B(n1458), .Z(n1460) );
  XOR U1576 ( .A(b[5]), .B(a[35]), .Z(n1496) );
  NANDN U1577 ( .A(n37), .B(n1496), .Z(n1459) );
  AND U1578 ( .A(n1460), .B(n1459), .Z(n1503) );
  AND U1579 ( .A(b[7]), .B(a[31]), .Z(n1502) );
  XNOR U1580 ( .A(n1503), .B(n1502), .Z(n1504) );
  XNOR U1581 ( .A(n1505), .B(n1504), .Z(n1510) );
  XOR U1582 ( .A(n1511), .B(n1510), .Z(n1485) );
  NANDN U1583 ( .A(n1462), .B(n1461), .Z(n1466) );
  NANDN U1584 ( .A(n1464), .B(n1463), .Z(n1465) );
  AND U1585 ( .A(n1466), .B(n1465), .Z(n1484) );
  XNOR U1586 ( .A(n1485), .B(n1484), .Z(n1486) );
  NANDN U1587 ( .A(n1468), .B(n1467), .Z(n1472) );
  NAND U1588 ( .A(n1470), .B(n1469), .Z(n1471) );
  NAND U1589 ( .A(n1472), .B(n1471), .Z(n1487) );
  XNOR U1590 ( .A(n1486), .B(n1487), .Z(n1478) );
  XNOR U1591 ( .A(n1479), .B(n1478), .Z(n1480) );
  XNOR U1592 ( .A(n1481), .B(n1480), .Z(n1514) );
  XNOR U1593 ( .A(sreg[95]), .B(n1514), .Z(n1516) );
  NANDN U1594 ( .A(sreg[94]), .B(n1473), .Z(n1477) );
  NAND U1595 ( .A(n1475), .B(n1474), .Z(n1476) );
  NAND U1596 ( .A(n1477), .B(n1476), .Z(n1515) );
  XNOR U1597 ( .A(n1516), .B(n1515), .Z(c[95]) );
  NANDN U1598 ( .A(n1479), .B(n1478), .Z(n1483) );
  NANDN U1599 ( .A(n1481), .B(n1480), .Z(n1482) );
  AND U1600 ( .A(n1483), .B(n1482), .Z(n1522) );
  NANDN U1601 ( .A(n1485), .B(n1484), .Z(n1489) );
  NANDN U1602 ( .A(n1487), .B(n1486), .Z(n1488) );
  AND U1603 ( .A(n1489), .B(n1488), .Z(n1520) );
  NANDN U1604 ( .A(n2629), .B(n1490), .Z(n1492) );
  XOR U1605 ( .A(b[7]), .B(a[34]), .Z(n1531) );
  NANDN U1606 ( .A(n2630), .B(n1531), .Z(n1491) );
  AND U1607 ( .A(n1492), .B(n1491), .Z(n1550) );
  NANDN U1608 ( .A(n2483), .B(n1493), .Z(n1495) );
  XOR U1609 ( .A(b[3]), .B(a[38]), .Z(n1534) );
  NANDN U1610 ( .A(n2484), .B(n1534), .Z(n1494) );
  NAND U1611 ( .A(n1495), .B(n1494), .Z(n1549) );
  XNOR U1612 ( .A(n1550), .B(n1549), .Z(n1552) );
  NAND U1613 ( .A(n2633), .B(n1496), .Z(n1498) );
  XOR U1614 ( .A(b[5]), .B(a[36]), .Z(n1540) );
  NANDN U1615 ( .A(n37), .B(n1540), .Z(n1497) );
  AND U1616 ( .A(n1498), .B(n1497), .Z(n1544) );
  AND U1617 ( .A(b[7]), .B(a[32]), .Z(n1543) );
  XNOR U1618 ( .A(n1544), .B(n1543), .Z(n1545) );
  NAND U1619 ( .A(b[0]), .B(a[40]), .Z(n1499) );
  XNOR U1620 ( .A(b[1]), .B(n1499), .Z(n1501) );
  NANDN U1621 ( .A(b[0]), .B(a[39]), .Z(n1500) );
  NAND U1622 ( .A(n1501), .B(n1500), .Z(n1546) );
  XNOR U1623 ( .A(n1545), .B(n1546), .Z(n1551) );
  XOR U1624 ( .A(n1552), .B(n1551), .Z(n1526) );
  NANDN U1625 ( .A(n1503), .B(n1502), .Z(n1507) );
  NANDN U1626 ( .A(n1505), .B(n1504), .Z(n1506) );
  AND U1627 ( .A(n1507), .B(n1506), .Z(n1525) );
  XNOR U1628 ( .A(n1526), .B(n1525), .Z(n1527) );
  NANDN U1629 ( .A(n1509), .B(n1508), .Z(n1513) );
  NAND U1630 ( .A(n1511), .B(n1510), .Z(n1512) );
  NAND U1631 ( .A(n1513), .B(n1512), .Z(n1528) );
  XNOR U1632 ( .A(n1527), .B(n1528), .Z(n1519) );
  XNOR U1633 ( .A(n1520), .B(n1519), .Z(n1521) );
  XNOR U1634 ( .A(n1522), .B(n1521), .Z(n1555) );
  XNOR U1635 ( .A(sreg[96]), .B(n1555), .Z(n1557) );
  NANDN U1636 ( .A(sreg[95]), .B(n1514), .Z(n1518) );
  NAND U1637 ( .A(n1516), .B(n1515), .Z(n1517) );
  NAND U1638 ( .A(n1518), .B(n1517), .Z(n1556) );
  XNOR U1639 ( .A(n1557), .B(n1556), .Z(c[96]) );
  NANDN U1640 ( .A(n1520), .B(n1519), .Z(n1524) );
  NANDN U1641 ( .A(n1522), .B(n1521), .Z(n1523) );
  AND U1642 ( .A(n1524), .B(n1523), .Z(n1563) );
  NANDN U1643 ( .A(n1526), .B(n1525), .Z(n1530) );
  NANDN U1644 ( .A(n1528), .B(n1527), .Z(n1529) );
  AND U1645 ( .A(n1530), .B(n1529), .Z(n1561) );
  NANDN U1646 ( .A(n2629), .B(n1531), .Z(n1533) );
  XOR U1647 ( .A(b[7]), .B(a[35]), .Z(n1572) );
  NANDN U1648 ( .A(n2630), .B(n1572), .Z(n1532) );
  AND U1649 ( .A(n1533), .B(n1532), .Z(n1591) );
  NANDN U1650 ( .A(n2483), .B(n1534), .Z(n1536) );
  XOR U1651 ( .A(b[3]), .B(a[39]), .Z(n1575) );
  NANDN U1652 ( .A(n2484), .B(n1575), .Z(n1535) );
  NAND U1653 ( .A(n1536), .B(n1535), .Z(n1590) );
  XNOR U1654 ( .A(n1591), .B(n1590), .Z(n1593) );
  NAND U1655 ( .A(b[0]), .B(a[41]), .Z(n1537) );
  XNOR U1656 ( .A(b[1]), .B(n1537), .Z(n1539) );
  NANDN U1657 ( .A(b[0]), .B(a[40]), .Z(n1538) );
  NAND U1658 ( .A(n1539), .B(n1538), .Z(n1587) );
  NAND U1659 ( .A(n2633), .B(n1540), .Z(n1542) );
  XOR U1660 ( .A(b[5]), .B(a[37]), .Z(n1581) );
  NANDN U1661 ( .A(n37), .B(n1581), .Z(n1541) );
  AND U1662 ( .A(n1542), .B(n1541), .Z(n1585) );
  AND U1663 ( .A(b[7]), .B(a[33]), .Z(n1584) );
  XNOR U1664 ( .A(n1585), .B(n1584), .Z(n1586) );
  XNOR U1665 ( .A(n1587), .B(n1586), .Z(n1592) );
  XOR U1666 ( .A(n1593), .B(n1592), .Z(n1567) );
  NANDN U1667 ( .A(n1544), .B(n1543), .Z(n1548) );
  NANDN U1668 ( .A(n1546), .B(n1545), .Z(n1547) );
  AND U1669 ( .A(n1548), .B(n1547), .Z(n1566) );
  XNOR U1670 ( .A(n1567), .B(n1566), .Z(n1568) );
  NANDN U1671 ( .A(n1550), .B(n1549), .Z(n1554) );
  NAND U1672 ( .A(n1552), .B(n1551), .Z(n1553) );
  NAND U1673 ( .A(n1554), .B(n1553), .Z(n1569) );
  XNOR U1674 ( .A(n1568), .B(n1569), .Z(n1560) );
  XNOR U1675 ( .A(n1561), .B(n1560), .Z(n1562) );
  XNOR U1676 ( .A(n1563), .B(n1562), .Z(n1596) );
  XNOR U1677 ( .A(sreg[97]), .B(n1596), .Z(n1598) );
  NANDN U1678 ( .A(sreg[96]), .B(n1555), .Z(n1559) );
  NAND U1679 ( .A(n1557), .B(n1556), .Z(n1558) );
  NAND U1680 ( .A(n1559), .B(n1558), .Z(n1597) );
  XNOR U1681 ( .A(n1598), .B(n1597), .Z(c[97]) );
  NANDN U1682 ( .A(n1561), .B(n1560), .Z(n1565) );
  NANDN U1683 ( .A(n1563), .B(n1562), .Z(n1564) );
  AND U1684 ( .A(n1565), .B(n1564), .Z(n1604) );
  NANDN U1685 ( .A(n1567), .B(n1566), .Z(n1571) );
  NANDN U1686 ( .A(n1569), .B(n1568), .Z(n1570) );
  AND U1687 ( .A(n1571), .B(n1570), .Z(n1602) );
  NANDN U1688 ( .A(n2629), .B(n1572), .Z(n1574) );
  XOR U1689 ( .A(b[7]), .B(a[36]), .Z(n1613) );
  NANDN U1690 ( .A(n2630), .B(n1613), .Z(n1573) );
  AND U1691 ( .A(n1574), .B(n1573), .Z(n1632) );
  NANDN U1692 ( .A(n2483), .B(n1575), .Z(n1577) );
  XOR U1693 ( .A(b[3]), .B(a[40]), .Z(n1616) );
  NANDN U1694 ( .A(n2484), .B(n1616), .Z(n1576) );
  NAND U1695 ( .A(n1577), .B(n1576), .Z(n1631) );
  XNOR U1696 ( .A(n1632), .B(n1631), .Z(n1634) );
  NAND U1697 ( .A(b[0]), .B(a[42]), .Z(n1578) );
  XNOR U1698 ( .A(b[1]), .B(n1578), .Z(n1580) );
  NANDN U1699 ( .A(b[0]), .B(a[41]), .Z(n1579) );
  NAND U1700 ( .A(n1580), .B(n1579), .Z(n1628) );
  NAND U1701 ( .A(n2633), .B(n1581), .Z(n1583) );
  XOR U1702 ( .A(b[5]), .B(a[38]), .Z(n1619) );
  NANDN U1703 ( .A(n37), .B(n1619), .Z(n1582) );
  AND U1704 ( .A(n1583), .B(n1582), .Z(n1626) );
  AND U1705 ( .A(b[7]), .B(a[34]), .Z(n1625) );
  XNOR U1706 ( .A(n1626), .B(n1625), .Z(n1627) );
  XNOR U1707 ( .A(n1628), .B(n1627), .Z(n1633) );
  XOR U1708 ( .A(n1634), .B(n1633), .Z(n1608) );
  NANDN U1709 ( .A(n1585), .B(n1584), .Z(n1589) );
  NANDN U1710 ( .A(n1587), .B(n1586), .Z(n1588) );
  AND U1711 ( .A(n1589), .B(n1588), .Z(n1607) );
  XNOR U1712 ( .A(n1608), .B(n1607), .Z(n1609) );
  NANDN U1713 ( .A(n1591), .B(n1590), .Z(n1595) );
  NAND U1714 ( .A(n1593), .B(n1592), .Z(n1594) );
  NAND U1715 ( .A(n1595), .B(n1594), .Z(n1610) );
  XNOR U1716 ( .A(n1609), .B(n1610), .Z(n1601) );
  XNOR U1717 ( .A(n1602), .B(n1601), .Z(n1603) );
  XNOR U1718 ( .A(n1604), .B(n1603), .Z(n1637) );
  XNOR U1719 ( .A(sreg[98]), .B(n1637), .Z(n1639) );
  NANDN U1720 ( .A(sreg[97]), .B(n1596), .Z(n1600) );
  NAND U1721 ( .A(n1598), .B(n1597), .Z(n1599) );
  NAND U1722 ( .A(n1600), .B(n1599), .Z(n1638) );
  XNOR U1723 ( .A(n1639), .B(n1638), .Z(c[98]) );
  NANDN U1724 ( .A(n1602), .B(n1601), .Z(n1606) );
  NANDN U1725 ( .A(n1604), .B(n1603), .Z(n1605) );
  AND U1726 ( .A(n1606), .B(n1605), .Z(n1645) );
  NANDN U1727 ( .A(n1608), .B(n1607), .Z(n1612) );
  NANDN U1728 ( .A(n1610), .B(n1609), .Z(n1611) );
  AND U1729 ( .A(n1612), .B(n1611), .Z(n1643) );
  NANDN U1730 ( .A(n2629), .B(n1613), .Z(n1615) );
  XOR U1731 ( .A(b[7]), .B(a[37]), .Z(n1654) );
  NANDN U1732 ( .A(n2630), .B(n1654), .Z(n1614) );
  AND U1733 ( .A(n1615), .B(n1614), .Z(n1673) );
  NANDN U1734 ( .A(n2483), .B(n1616), .Z(n1618) );
  XOR U1735 ( .A(b[3]), .B(a[41]), .Z(n1657) );
  NANDN U1736 ( .A(n2484), .B(n1657), .Z(n1617) );
  NAND U1737 ( .A(n1618), .B(n1617), .Z(n1672) );
  XNOR U1738 ( .A(n1673), .B(n1672), .Z(n1675) );
  NAND U1739 ( .A(n2633), .B(n1619), .Z(n1621) );
  XOR U1740 ( .A(b[5]), .B(a[39]), .Z(n1660) );
  NANDN U1741 ( .A(n37), .B(n1660), .Z(n1620) );
  AND U1742 ( .A(n1621), .B(n1620), .Z(n1667) );
  AND U1743 ( .A(b[7]), .B(a[35]), .Z(n1666) );
  XNOR U1744 ( .A(n1667), .B(n1666), .Z(n1668) );
  NAND U1745 ( .A(b[0]), .B(a[43]), .Z(n1622) );
  XNOR U1746 ( .A(b[1]), .B(n1622), .Z(n1624) );
  NANDN U1747 ( .A(b[0]), .B(a[42]), .Z(n1623) );
  NAND U1748 ( .A(n1624), .B(n1623), .Z(n1669) );
  XNOR U1749 ( .A(n1668), .B(n1669), .Z(n1674) );
  XOR U1750 ( .A(n1675), .B(n1674), .Z(n1649) );
  NANDN U1751 ( .A(n1626), .B(n1625), .Z(n1630) );
  NANDN U1752 ( .A(n1628), .B(n1627), .Z(n1629) );
  AND U1753 ( .A(n1630), .B(n1629), .Z(n1648) );
  XNOR U1754 ( .A(n1649), .B(n1648), .Z(n1650) );
  NANDN U1755 ( .A(n1632), .B(n1631), .Z(n1636) );
  NAND U1756 ( .A(n1634), .B(n1633), .Z(n1635) );
  NAND U1757 ( .A(n1636), .B(n1635), .Z(n1651) );
  XNOR U1758 ( .A(n1650), .B(n1651), .Z(n1642) );
  XNOR U1759 ( .A(n1643), .B(n1642), .Z(n1644) );
  XNOR U1760 ( .A(n1645), .B(n1644), .Z(n1678) );
  XNOR U1761 ( .A(sreg[99]), .B(n1678), .Z(n1680) );
  NANDN U1762 ( .A(sreg[98]), .B(n1637), .Z(n1641) );
  NAND U1763 ( .A(n1639), .B(n1638), .Z(n1640) );
  NAND U1764 ( .A(n1641), .B(n1640), .Z(n1679) );
  XNOR U1765 ( .A(n1680), .B(n1679), .Z(c[99]) );
  NANDN U1766 ( .A(n1643), .B(n1642), .Z(n1647) );
  NANDN U1767 ( .A(n1645), .B(n1644), .Z(n1646) );
  AND U1768 ( .A(n1647), .B(n1646), .Z(n1686) );
  NANDN U1769 ( .A(n1649), .B(n1648), .Z(n1653) );
  NANDN U1770 ( .A(n1651), .B(n1650), .Z(n1652) );
  AND U1771 ( .A(n1653), .B(n1652), .Z(n1684) );
  NANDN U1772 ( .A(n2629), .B(n1654), .Z(n1656) );
  XOR U1773 ( .A(b[7]), .B(a[38]), .Z(n1695) );
  NANDN U1774 ( .A(n2630), .B(n1695), .Z(n1655) );
  AND U1775 ( .A(n1656), .B(n1655), .Z(n1714) );
  NANDN U1776 ( .A(n2483), .B(n1657), .Z(n1659) );
  XOR U1777 ( .A(b[3]), .B(a[42]), .Z(n1698) );
  NANDN U1778 ( .A(n2484), .B(n1698), .Z(n1658) );
  NAND U1779 ( .A(n1659), .B(n1658), .Z(n1713) );
  XNOR U1780 ( .A(n1714), .B(n1713), .Z(n1716) );
  NAND U1781 ( .A(n2633), .B(n1660), .Z(n1662) );
  XOR U1782 ( .A(b[5]), .B(a[40]), .Z(n1704) );
  NANDN U1783 ( .A(n37), .B(n1704), .Z(n1661) );
  AND U1784 ( .A(n1662), .B(n1661), .Z(n1708) );
  AND U1785 ( .A(b[7]), .B(a[36]), .Z(n1707) );
  XNOR U1786 ( .A(n1708), .B(n1707), .Z(n1709) );
  NAND U1787 ( .A(b[0]), .B(a[44]), .Z(n1663) );
  XNOR U1788 ( .A(b[1]), .B(n1663), .Z(n1665) );
  NANDN U1789 ( .A(b[0]), .B(a[43]), .Z(n1664) );
  NAND U1790 ( .A(n1665), .B(n1664), .Z(n1710) );
  XNOR U1791 ( .A(n1709), .B(n1710), .Z(n1715) );
  XOR U1792 ( .A(n1716), .B(n1715), .Z(n1690) );
  NANDN U1793 ( .A(n1667), .B(n1666), .Z(n1671) );
  NANDN U1794 ( .A(n1669), .B(n1668), .Z(n1670) );
  AND U1795 ( .A(n1671), .B(n1670), .Z(n1689) );
  XNOR U1796 ( .A(n1690), .B(n1689), .Z(n1691) );
  NANDN U1797 ( .A(n1673), .B(n1672), .Z(n1677) );
  NAND U1798 ( .A(n1675), .B(n1674), .Z(n1676) );
  NAND U1799 ( .A(n1677), .B(n1676), .Z(n1692) );
  XNOR U1800 ( .A(n1691), .B(n1692), .Z(n1683) );
  XNOR U1801 ( .A(n1684), .B(n1683), .Z(n1685) );
  XNOR U1802 ( .A(n1686), .B(n1685), .Z(n1719) );
  XNOR U1803 ( .A(sreg[100]), .B(n1719), .Z(n1721) );
  NANDN U1804 ( .A(sreg[99]), .B(n1678), .Z(n1682) );
  NAND U1805 ( .A(n1680), .B(n1679), .Z(n1681) );
  NAND U1806 ( .A(n1682), .B(n1681), .Z(n1720) );
  XNOR U1807 ( .A(n1721), .B(n1720), .Z(c[100]) );
  NANDN U1808 ( .A(n1684), .B(n1683), .Z(n1688) );
  NANDN U1809 ( .A(n1686), .B(n1685), .Z(n1687) );
  AND U1810 ( .A(n1688), .B(n1687), .Z(n1727) );
  NANDN U1811 ( .A(n1690), .B(n1689), .Z(n1694) );
  NANDN U1812 ( .A(n1692), .B(n1691), .Z(n1693) );
  AND U1813 ( .A(n1694), .B(n1693), .Z(n1725) );
  NANDN U1814 ( .A(n2629), .B(n1695), .Z(n1697) );
  XOR U1815 ( .A(b[7]), .B(a[39]), .Z(n1736) );
  NANDN U1816 ( .A(n2630), .B(n1736), .Z(n1696) );
  AND U1817 ( .A(n1697), .B(n1696), .Z(n1755) );
  NANDN U1818 ( .A(n2483), .B(n1698), .Z(n1700) );
  XOR U1819 ( .A(b[3]), .B(a[43]), .Z(n1739) );
  NANDN U1820 ( .A(n2484), .B(n1739), .Z(n1699) );
  NAND U1821 ( .A(n1700), .B(n1699), .Z(n1754) );
  XNOR U1822 ( .A(n1755), .B(n1754), .Z(n1757) );
  NAND U1823 ( .A(b[0]), .B(a[45]), .Z(n1701) );
  XNOR U1824 ( .A(b[1]), .B(n1701), .Z(n1703) );
  NANDN U1825 ( .A(b[0]), .B(a[44]), .Z(n1702) );
  NAND U1826 ( .A(n1703), .B(n1702), .Z(n1751) );
  NAND U1827 ( .A(n2633), .B(n1704), .Z(n1706) );
  XOR U1828 ( .A(b[5]), .B(a[41]), .Z(n1745) );
  NANDN U1829 ( .A(n37), .B(n1745), .Z(n1705) );
  AND U1830 ( .A(n1706), .B(n1705), .Z(n1749) );
  AND U1831 ( .A(b[7]), .B(a[37]), .Z(n1748) );
  XNOR U1832 ( .A(n1749), .B(n1748), .Z(n1750) );
  XNOR U1833 ( .A(n1751), .B(n1750), .Z(n1756) );
  XOR U1834 ( .A(n1757), .B(n1756), .Z(n1731) );
  NANDN U1835 ( .A(n1708), .B(n1707), .Z(n1712) );
  NANDN U1836 ( .A(n1710), .B(n1709), .Z(n1711) );
  AND U1837 ( .A(n1712), .B(n1711), .Z(n1730) );
  XNOR U1838 ( .A(n1731), .B(n1730), .Z(n1732) );
  NANDN U1839 ( .A(n1714), .B(n1713), .Z(n1718) );
  NAND U1840 ( .A(n1716), .B(n1715), .Z(n1717) );
  NAND U1841 ( .A(n1718), .B(n1717), .Z(n1733) );
  XNOR U1842 ( .A(n1732), .B(n1733), .Z(n1724) );
  XNOR U1843 ( .A(n1725), .B(n1724), .Z(n1726) );
  XNOR U1844 ( .A(n1727), .B(n1726), .Z(n1760) );
  XNOR U1845 ( .A(sreg[101]), .B(n1760), .Z(n1762) );
  NANDN U1846 ( .A(sreg[100]), .B(n1719), .Z(n1723) );
  NAND U1847 ( .A(n1721), .B(n1720), .Z(n1722) );
  NAND U1848 ( .A(n1723), .B(n1722), .Z(n1761) );
  XNOR U1849 ( .A(n1762), .B(n1761), .Z(c[101]) );
  NANDN U1850 ( .A(n1725), .B(n1724), .Z(n1729) );
  NANDN U1851 ( .A(n1727), .B(n1726), .Z(n1728) );
  AND U1852 ( .A(n1729), .B(n1728), .Z(n1768) );
  NANDN U1853 ( .A(n1731), .B(n1730), .Z(n1735) );
  NANDN U1854 ( .A(n1733), .B(n1732), .Z(n1734) );
  AND U1855 ( .A(n1735), .B(n1734), .Z(n1766) );
  NANDN U1856 ( .A(n2629), .B(n1736), .Z(n1738) );
  XOR U1857 ( .A(b[7]), .B(a[40]), .Z(n1777) );
  NANDN U1858 ( .A(n2630), .B(n1777), .Z(n1737) );
  AND U1859 ( .A(n1738), .B(n1737), .Z(n1796) );
  NANDN U1860 ( .A(n2483), .B(n1739), .Z(n1741) );
  XOR U1861 ( .A(b[3]), .B(a[44]), .Z(n1780) );
  NANDN U1862 ( .A(n2484), .B(n1780), .Z(n1740) );
  NAND U1863 ( .A(n1741), .B(n1740), .Z(n1795) );
  XNOR U1864 ( .A(n1796), .B(n1795), .Z(n1798) );
  NAND U1865 ( .A(b[0]), .B(a[46]), .Z(n1742) );
  XNOR U1866 ( .A(b[1]), .B(n1742), .Z(n1744) );
  NANDN U1867 ( .A(b[0]), .B(a[45]), .Z(n1743) );
  NAND U1868 ( .A(n1744), .B(n1743), .Z(n1792) );
  NAND U1869 ( .A(n2633), .B(n1745), .Z(n1747) );
  XOR U1870 ( .A(b[5]), .B(a[42]), .Z(n1786) );
  NANDN U1871 ( .A(n37), .B(n1786), .Z(n1746) );
  AND U1872 ( .A(n1747), .B(n1746), .Z(n1790) );
  AND U1873 ( .A(b[7]), .B(a[38]), .Z(n1789) );
  XNOR U1874 ( .A(n1790), .B(n1789), .Z(n1791) );
  XNOR U1875 ( .A(n1792), .B(n1791), .Z(n1797) );
  XOR U1876 ( .A(n1798), .B(n1797), .Z(n1772) );
  NANDN U1877 ( .A(n1749), .B(n1748), .Z(n1753) );
  NANDN U1878 ( .A(n1751), .B(n1750), .Z(n1752) );
  AND U1879 ( .A(n1753), .B(n1752), .Z(n1771) );
  XNOR U1880 ( .A(n1772), .B(n1771), .Z(n1773) );
  NANDN U1881 ( .A(n1755), .B(n1754), .Z(n1759) );
  NAND U1882 ( .A(n1757), .B(n1756), .Z(n1758) );
  NAND U1883 ( .A(n1759), .B(n1758), .Z(n1774) );
  XNOR U1884 ( .A(n1773), .B(n1774), .Z(n1765) );
  XNOR U1885 ( .A(n1766), .B(n1765), .Z(n1767) );
  XNOR U1886 ( .A(n1768), .B(n1767), .Z(n1801) );
  XNOR U1887 ( .A(sreg[102]), .B(n1801), .Z(n1803) );
  NANDN U1888 ( .A(sreg[101]), .B(n1760), .Z(n1764) );
  NAND U1889 ( .A(n1762), .B(n1761), .Z(n1763) );
  NAND U1890 ( .A(n1764), .B(n1763), .Z(n1802) );
  XNOR U1891 ( .A(n1803), .B(n1802), .Z(c[102]) );
  NANDN U1892 ( .A(n1766), .B(n1765), .Z(n1770) );
  NANDN U1893 ( .A(n1768), .B(n1767), .Z(n1769) );
  AND U1894 ( .A(n1770), .B(n1769), .Z(n1809) );
  NANDN U1895 ( .A(n1772), .B(n1771), .Z(n1776) );
  NANDN U1896 ( .A(n1774), .B(n1773), .Z(n1775) );
  AND U1897 ( .A(n1776), .B(n1775), .Z(n1807) );
  NANDN U1898 ( .A(n2629), .B(n1777), .Z(n1779) );
  XOR U1899 ( .A(b[7]), .B(a[41]), .Z(n1818) );
  NANDN U1900 ( .A(n2630), .B(n1818), .Z(n1778) );
  AND U1901 ( .A(n1779), .B(n1778), .Z(n1837) );
  NANDN U1902 ( .A(n2483), .B(n1780), .Z(n1782) );
  XOR U1903 ( .A(b[3]), .B(a[45]), .Z(n1821) );
  NANDN U1904 ( .A(n2484), .B(n1821), .Z(n1781) );
  NAND U1905 ( .A(n1782), .B(n1781), .Z(n1836) );
  XNOR U1906 ( .A(n1837), .B(n1836), .Z(n1839) );
  NAND U1907 ( .A(b[0]), .B(a[47]), .Z(n1783) );
  XNOR U1908 ( .A(b[1]), .B(n1783), .Z(n1785) );
  NANDN U1909 ( .A(b[0]), .B(a[46]), .Z(n1784) );
  NAND U1910 ( .A(n1785), .B(n1784), .Z(n1833) );
  NAND U1911 ( .A(n2633), .B(n1786), .Z(n1788) );
  XOR U1912 ( .A(b[5]), .B(a[43]), .Z(n1827) );
  NANDN U1913 ( .A(n37), .B(n1827), .Z(n1787) );
  AND U1914 ( .A(n1788), .B(n1787), .Z(n1831) );
  AND U1915 ( .A(b[7]), .B(a[39]), .Z(n1830) );
  XNOR U1916 ( .A(n1831), .B(n1830), .Z(n1832) );
  XNOR U1917 ( .A(n1833), .B(n1832), .Z(n1838) );
  XOR U1918 ( .A(n1839), .B(n1838), .Z(n1813) );
  NANDN U1919 ( .A(n1790), .B(n1789), .Z(n1794) );
  NANDN U1920 ( .A(n1792), .B(n1791), .Z(n1793) );
  AND U1921 ( .A(n1794), .B(n1793), .Z(n1812) );
  XNOR U1922 ( .A(n1813), .B(n1812), .Z(n1814) );
  NANDN U1923 ( .A(n1796), .B(n1795), .Z(n1800) );
  NAND U1924 ( .A(n1798), .B(n1797), .Z(n1799) );
  NAND U1925 ( .A(n1800), .B(n1799), .Z(n1815) );
  XNOR U1926 ( .A(n1814), .B(n1815), .Z(n1806) );
  XNOR U1927 ( .A(n1807), .B(n1806), .Z(n1808) );
  XNOR U1928 ( .A(n1809), .B(n1808), .Z(n1842) );
  XNOR U1929 ( .A(sreg[103]), .B(n1842), .Z(n1844) );
  NANDN U1930 ( .A(sreg[102]), .B(n1801), .Z(n1805) );
  NAND U1931 ( .A(n1803), .B(n1802), .Z(n1804) );
  NAND U1932 ( .A(n1805), .B(n1804), .Z(n1843) );
  XNOR U1933 ( .A(n1844), .B(n1843), .Z(c[103]) );
  NANDN U1934 ( .A(n1807), .B(n1806), .Z(n1811) );
  NANDN U1935 ( .A(n1809), .B(n1808), .Z(n1810) );
  AND U1936 ( .A(n1811), .B(n1810), .Z(n1850) );
  NANDN U1937 ( .A(n1813), .B(n1812), .Z(n1817) );
  NANDN U1938 ( .A(n1815), .B(n1814), .Z(n1816) );
  AND U1939 ( .A(n1817), .B(n1816), .Z(n1848) );
  NANDN U1940 ( .A(n2629), .B(n1818), .Z(n1820) );
  XOR U1941 ( .A(b[7]), .B(a[42]), .Z(n1859) );
  NANDN U1942 ( .A(n2630), .B(n1859), .Z(n1819) );
  AND U1943 ( .A(n1820), .B(n1819), .Z(n1878) );
  NANDN U1944 ( .A(n2483), .B(n1821), .Z(n1823) );
  XOR U1945 ( .A(b[3]), .B(a[46]), .Z(n1862) );
  NANDN U1946 ( .A(n2484), .B(n1862), .Z(n1822) );
  NAND U1947 ( .A(n1823), .B(n1822), .Z(n1877) );
  XNOR U1948 ( .A(n1878), .B(n1877), .Z(n1880) );
  NAND U1949 ( .A(b[0]), .B(a[48]), .Z(n1824) );
  XNOR U1950 ( .A(b[1]), .B(n1824), .Z(n1826) );
  NANDN U1951 ( .A(b[0]), .B(a[47]), .Z(n1825) );
  NAND U1952 ( .A(n1826), .B(n1825), .Z(n1874) );
  NAND U1953 ( .A(n2633), .B(n1827), .Z(n1829) );
  XOR U1954 ( .A(b[5]), .B(a[44]), .Z(n1868) );
  NANDN U1955 ( .A(n37), .B(n1868), .Z(n1828) );
  AND U1956 ( .A(n1829), .B(n1828), .Z(n1872) );
  AND U1957 ( .A(b[7]), .B(a[40]), .Z(n1871) );
  XNOR U1958 ( .A(n1872), .B(n1871), .Z(n1873) );
  XNOR U1959 ( .A(n1874), .B(n1873), .Z(n1879) );
  XOR U1960 ( .A(n1880), .B(n1879), .Z(n1854) );
  NANDN U1961 ( .A(n1831), .B(n1830), .Z(n1835) );
  NANDN U1962 ( .A(n1833), .B(n1832), .Z(n1834) );
  AND U1963 ( .A(n1835), .B(n1834), .Z(n1853) );
  XNOR U1964 ( .A(n1854), .B(n1853), .Z(n1855) );
  NANDN U1965 ( .A(n1837), .B(n1836), .Z(n1841) );
  NAND U1966 ( .A(n1839), .B(n1838), .Z(n1840) );
  NAND U1967 ( .A(n1841), .B(n1840), .Z(n1856) );
  XNOR U1968 ( .A(n1855), .B(n1856), .Z(n1847) );
  XNOR U1969 ( .A(n1848), .B(n1847), .Z(n1849) );
  XNOR U1970 ( .A(n1850), .B(n1849), .Z(n1883) );
  XNOR U1971 ( .A(sreg[104]), .B(n1883), .Z(n1885) );
  NANDN U1972 ( .A(sreg[103]), .B(n1842), .Z(n1846) );
  NAND U1973 ( .A(n1844), .B(n1843), .Z(n1845) );
  NAND U1974 ( .A(n1846), .B(n1845), .Z(n1884) );
  XNOR U1975 ( .A(n1885), .B(n1884), .Z(c[104]) );
  NANDN U1976 ( .A(n1848), .B(n1847), .Z(n1852) );
  NANDN U1977 ( .A(n1850), .B(n1849), .Z(n1851) );
  AND U1978 ( .A(n1852), .B(n1851), .Z(n1891) );
  NANDN U1979 ( .A(n1854), .B(n1853), .Z(n1858) );
  NANDN U1980 ( .A(n1856), .B(n1855), .Z(n1857) );
  AND U1981 ( .A(n1858), .B(n1857), .Z(n1889) );
  NANDN U1982 ( .A(n2629), .B(n1859), .Z(n1861) );
  XOR U1983 ( .A(b[7]), .B(a[43]), .Z(n1900) );
  NANDN U1984 ( .A(n2630), .B(n1900), .Z(n1860) );
  AND U1985 ( .A(n1861), .B(n1860), .Z(n1919) );
  NANDN U1986 ( .A(n2483), .B(n1862), .Z(n1864) );
  XOR U1987 ( .A(b[3]), .B(a[47]), .Z(n1903) );
  NANDN U1988 ( .A(n2484), .B(n1903), .Z(n1863) );
  NAND U1989 ( .A(n1864), .B(n1863), .Z(n1918) );
  XNOR U1990 ( .A(n1919), .B(n1918), .Z(n1921) );
  NAND U1991 ( .A(b[0]), .B(a[49]), .Z(n1865) );
  XNOR U1992 ( .A(b[1]), .B(n1865), .Z(n1867) );
  NANDN U1993 ( .A(b[0]), .B(a[48]), .Z(n1866) );
  NAND U1994 ( .A(n1867), .B(n1866), .Z(n1915) );
  NAND U1995 ( .A(n2633), .B(n1868), .Z(n1870) );
  XOR U1996 ( .A(b[5]), .B(a[45]), .Z(n1906) );
  NANDN U1997 ( .A(n37), .B(n1906), .Z(n1869) );
  AND U1998 ( .A(n1870), .B(n1869), .Z(n1913) );
  AND U1999 ( .A(b[7]), .B(a[41]), .Z(n1912) );
  XNOR U2000 ( .A(n1913), .B(n1912), .Z(n1914) );
  XNOR U2001 ( .A(n1915), .B(n1914), .Z(n1920) );
  XOR U2002 ( .A(n1921), .B(n1920), .Z(n1895) );
  NANDN U2003 ( .A(n1872), .B(n1871), .Z(n1876) );
  NANDN U2004 ( .A(n1874), .B(n1873), .Z(n1875) );
  AND U2005 ( .A(n1876), .B(n1875), .Z(n1894) );
  XNOR U2006 ( .A(n1895), .B(n1894), .Z(n1896) );
  NANDN U2007 ( .A(n1878), .B(n1877), .Z(n1882) );
  NAND U2008 ( .A(n1880), .B(n1879), .Z(n1881) );
  NAND U2009 ( .A(n1882), .B(n1881), .Z(n1897) );
  XNOR U2010 ( .A(n1896), .B(n1897), .Z(n1888) );
  XNOR U2011 ( .A(n1889), .B(n1888), .Z(n1890) );
  XNOR U2012 ( .A(n1891), .B(n1890), .Z(n1924) );
  XNOR U2013 ( .A(sreg[105]), .B(n1924), .Z(n1926) );
  NANDN U2014 ( .A(sreg[104]), .B(n1883), .Z(n1887) );
  NAND U2015 ( .A(n1885), .B(n1884), .Z(n1886) );
  NAND U2016 ( .A(n1887), .B(n1886), .Z(n1925) );
  XNOR U2017 ( .A(n1926), .B(n1925), .Z(c[105]) );
  NANDN U2018 ( .A(n1889), .B(n1888), .Z(n1893) );
  NANDN U2019 ( .A(n1891), .B(n1890), .Z(n1892) );
  AND U2020 ( .A(n1893), .B(n1892), .Z(n1932) );
  NANDN U2021 ( .A(n1895), .B(n1894), .Z(n1899) );
  NANDN U2022 ( .A(n1897), .B(n1896), .Z(n1898) );
  AND U2023 ( .A(n1899), .B(n1898), .Z(n1930) );
  NANDN U2024 ( .A(n2629), .B(n1900), .Z(n1902) );
  XOR U2025 ( .A(b[7]), .B(a[44]), .Z(n1941) );
  NANDN U2026 ( .A(n2630), .B(n1941), .Z(n1901) );
  AND U2027 ( .A(n1902), .B(n1901), .Z(n1960) );
  NANDN U2028 ( .A(n2483), .B(n1903), .Z(n1905) );
  XOR U2029 ( .A(b[3]), .B(a[48]), .Z(n1944) );
  NANDN U2030 ( .A(n2484), .B(n1944), .Z(n1904) );
  NAND U2031 ( .A(n1905), .B(n1904), .Z(n1959) );
  XNOR U2032 ( .A(n1960), .B(n1959), .Z(n1962) );
  NAND U2033 ( .A(n2633), .B(n1906), .Z(n1908) );
  XOR U2034 ( .A(b[5]), .B(a[46]), .Z(n1950) );
  NANDN U2035 ( .A(n37), .B(n1950), .Z(n1907) );
  AND U2036 ( .A(n1908), .B(n1907), .Z(n1954) );
  AND U2037 ( .A(b[7]), .B(a[42]), .Z(n1953) );
  XNOR U2038 ( .A(n1954), .B(n1953), .Z(n1955) );
  NAND U2039 ( .A(b[0]), .B(a[50]), .Z(n1909) );
  XNOR U2040 ( .A(b[1]), .B(n1909), .Z(n1911) );
  NANDN U2041 ( .A(b[0]), .B(a[49]), .Z(n1910) );
  NAND U2042 ( .A(n1911), .B(n1910), .Z(n1956) );
  XNOR U2043 ( .A(n1955), .B(n1956), .Z(n1961) );
  XOR U2044 ( .A(n1962), .B(n1961), .Z(n1936) );
  NANDN U2045 ( .A(n1913), .B(n1912), .Z(n1917) );
  NANDN U2046 ( .A(n1915), .B(n1914), .Z(n1916) );
  AND U2047 ( .A(n1917), .B(n1916), .Z(n1935) );
  XNOR U2048 ( .A(n1936), .B(n1935), .Z(n1937) );
  NANDN U2049 ( .A(n1919), .B(n1918), .Z(n1923) );
  NAND U2050 ( .A(n1921), .B(n1920), .Z(n1922) );
  NAND U2051 ( .A(n1923), .B(n1922), .Z(n1938) );
  XNOR U2052 ( .A(n1937), .B(n1938), .Z(n1929) );
  XNOR U2053 ( .A(n1930), .B(n1929), .Z(n1931) );
  XNOR U2054 ( .A(n1932), .B(n1931), .Z(n1965) );
  XNOR U2055 ( .A(sreg[106]), .B(n1965), .Z(n1967) );
  NANDN U2056 ( .A(sreg[105]), .B(n1924), .Z(n1928) );
  NAND U2057 ( .A(n1926), .B(n1925), .Z(n1927) );
  NAND U2058 ( .A(n1928), .B(n1927), .Z(n1966) );
  XNOR U2059 ( .A(n1967), .B(n1966), .Z(c[106]) );
  NANDN U2060 ( .A(n1930), .B(n1929), .Z(n1934) );
  NANDN U2061 ( .A(n1932), .B(n1931), .Z(n1933) );
  AND U2062 ( .A(n1934), .B(n1933), .Z(n1973) );
  NANDN U2063 ( .A(n1936), .B(n1935), .Z(n1940) );
  NANDN U2064 ( .A(n1938), .B(n1937), .Z(n1939) );
  AND U2065 ( .A(n1940), .B(n1939), .Z(n1971) );
  NANDN U2066 ( .A(n2629), .B(n1941), .Z(n1943) );
  XOR U2067 ( .A(b[7]), .B(a[45]), .Z(n1982) );
  NANDN U2068 ( .A(n2630), .B(n1982), .Z(n1942) );
  AND U2069 ( .A(n1943), .B(n1942), .Z(n2001) );
  NANDN U2070 ( .A(n2483), .B(n1944), .Z(n1946) );
  XOR U2071 ( .A(b[3]), .B(a[49]), .Z(n1985) );
  NANDN U2072 ( .A(n2484), .B(n1985), .Z(n1945) );
  NAND U2073 ( .A(n1946), .B(n1945), .Z(n2000) );
  XNOR U2074 ( .A(n2001), .B(n2000), .Z(n2003) );
  NAND U2075 ( .A(b[0]), .B(a[51]), .Z(n1947) );
  XNOR U2076 ( .A(b[1]), .B(n1947), .Z(n1949) );
  NANDN U2077 ( .A(b[0]), .B(a[50]), .Z(n1948) );
  NAND U2078 ( .A(n1949), .B(n1948), .Z(n1997) );
  NAND U2079 ( .A(n2633), .B(n1950), .Z(n1952) );
  XOR U2080 ( .A(b[5]), .B(a[47]), .Z(n1991) );
  NANDN U2081 ( .A(n37), .B(n1991), .Z(n1951) );
  AND U2082 ( .A(n1952), .B(n1951), .Z(n1995) );
  AND U2083 ( .A(b[7]), .B(a[43]), .Z(n1994) );
  XNOR U2084 ( .A(n1995), .B(n1994), .Z(n1996) );
  XNOR U2085 ( .A(n1997), .B(n1996), .Z(n2002) );
  XOR U2086 ( .A(n2003), .B(n2002), .Z(n1977) );
  NANDN U2087 ( .A(n1954), .B(n1953), .Z(n1958) );
  NANDN U2088 ( .A(n1956), .B(n1955), .Z(n1957) );
  AND U2089 ( .A(n1958), .B(n1957), .Z(n1976) );
  XNOR U2090 ( .A(n1977), .B(n1976), .Z(n1978) );
  NANDN U2091 ( .A(n1960), .B(n1959), .Z(n1964) );
  NAND U2092 ( .A(n1962), .B(n1961), .Z(n1963) );
  NAND U2093 ( .A(n1964), .B(n1963), .Z(n1979) );
  XNOR U2094 ( .A(n1978), .B(n1979), .Z(n1970) );
  XNOR U2095 ( .A(n1971), .B(n1970), .Z(n1972) );
  XNOR U2096 ( .A(n1973), .B(n1972), .Z(n2006) );
  XNOR U2097 ( .A(sreg[107]), .B(n2006), .Z(n2008) );
  NANDN U2098 ( .A(sreg[106]), .B(n1965), .Z(n1969) );
  NAND U2099 ( .A(n1967), .B(n1966), .Z(n1968) );
  NAND U2100 ( .A(n1969), .B(n1968), .Z(n2007) );
  XNOR U2101 ( .A(n2008), .B(n2007), .Z(c[107]) );
  NANDN U2102 ( .A(n1971), .B(n1970), .Z(n1975) );
  NANDN U2103 ( .A(n1973), .B(n1972), .Z(n1974) );
  AND U2104 ( .A(n1975), .B(n1974), .Z(n2014) );
  NANDN U2105 ( .A(n1977), .B(n1976), .Z(n1981) );
  NANDN U2106 ( .A(n1979), .B(n1978), .Z(n1980) );
  AND U2107 ( .A(n1981), .B(n1980), .Z(n2012) );
  NANDN U2108 ( .A(n2629), .B(n1982), .Z(n1984) );
  XOR U2109 ( .A(b[7]), .B(a[46]), .Z(n2023) );
  NANDN U2110 ( .A(n2630), .B(n2023), .Z(n1983) );
  AND U2111 ( .A(n1984), .B(n1983), .Z(n2042) );
  NANDN U2112 ( .A(n2483), .B(n1985), .Z(n1987) );
  XOR U2113 ( .A(b[3]), .B(a[50]), .Z(n2026) );
  NANDN U2114 ( .A(n2484), .B(n2026), .Z(n1986) );
  NAND U2115 ( .A(n1987), .B(n1986), .Z(n2041) );
  XNOR U2116 ( .A(n2042), .B(n2041), .Z(n2044) );
  NAND U2117 ( .A(b[0]), .B(a[52]), .Z(n1988) );
  XNOR U2118 ( .A(b[1]), .B(n1988), .Z(n1990) );
  NANDN U2119 ( .A(b[0]), .B(a[51]), .Z(n1989) );
  NAND U2120 ( .A(n1990), .B(n1989), .Z(n2038) );
  NAND U2121 ( .A(n2633), .B(n1991), .Z(n1993) );
  XOR U2122 ( .A(b[5]), .B(a[48]), .Z(n2032) );
  NANDN U2123 ( .A(n37), .B(n2032), .Z(n1992) );
  AND U2124 ( .A(n1993), .B(n1992), .Z(n2036) );
  AND U2125 ( .A(b[7]), .B(a[44]), .Z(n2035) );
  XNOR U2126 ( .A(n2036), .B(n2035), .Z(n2037) );
  XNOR U2127 ( .A(n2038), .B(n2037), .Z(n2043) );
  XOR U2128 ( .A(n2044), .B(n2043), .Z(n2018) );
  NANDN U2129 ( .A(n1995), .B(n1994), .Z(n1999) );
  NANDN U2130 ( .A(n1997), .B(n1996), .Z(n1998) );
  AND U2131 ( .A(n1999), .B(n1998), .Z(n2017) );
  XNOR U2132 ( .A(n2018), .B(n2017), .Z(n2019) );
  NANDN U2133 ( .A(n2001), .B(n2000), .Z(n2005) );
  NAND U2134 ( .A(n2003), .B(n2002), .Z(n2004) );
  NAND U2135 ( .A(n2005), .B(n2004), .Z(n2020) );
  XNOR U2136 ( .A(n2019), .B(n2020), .Z(n2011) );
  XNOR U2137 ( .A(n2012), .B(n2011), .Z(n2013) );
  XNOR U2138 ( .A(n2014), .B(n2013), .Z(n2047) );
  XNOR U2139 ( .A(sreg[108]), .B(n2047), .Z(n2049) );
  NANDN U2140 ( .A(sreg[107]), .B(n2006), .Z(n2010) );
  NAND U2141 ( .A(n2008), .B(n2007), .Z(n2009) );
  NAND U2142 ( .A(n2010), .B(n2009), .Z(n2048) );
  XNOR U2143 ( .A(n2049), .B(n2048), .Z(c[108]) );
  NANDN U2144 ( .A(n2012), .B(n2011), .Z(n2016) );
  NANDN U2145 ( .A(n2014), .B(n2013), .Z(n2015) );
  AND U2146 ( .A(n2016), .B(n2015), .Z(n2055) );
  NANDN U2147 ( .A(n2018), .B(n2017), .Z(n2022) );
  NANDN U2148 ( .A(n2020), .B(n2019), .Z(n2021) );
  AND U2149 ( .A(n2022), .B(n2021), .Z(n2053) );
  NANDN U2150 ( .A(n2629), .B(n2023), .Z(n2025) );
  XOR U2151 ( .A(b[7]), .B(a[47]), .Z(n2064) );
  NANDN U2152 ( .A(n2630), .B(n2064), .Z(n2024) );
  AND U2153 ( .A(n2025), .B(n2024), .Z(n2083) );
  NANDN U2154 ( .A(n2483), .B(n2026), .Z(n2028) );
  XOR U2155 ( .A(b[3]), .B(a[51]), .Z(n2067) );
  NANDN U2156 ( .A(n2484), .B(n2067), .Z(n2027) );
  NAND U2157 ( .A(n2028), .B(n2027), .Z(n2082) );
  XNOR U2158 ( .A(n2083), .B(n2082), .Z(n2085) );
  NAND U2159 ( .A(b[0]), .B(a[53]), .Z(n2029) );
  XNOR U2160 ( .A(b[1]), .B(n2029), .Z(n2031) );
  NANDN U2161 ( .A(b[0]), .B(a[52]), .Z(n2030) );
  NAND U2162 ( .A(n2031), .B(n2030), .Z(n2079) );
  NAND U2163 ( .A(n2633), .B(n2032), .Z(n2034) );
  XOR U2164 ( .A(b[5]), .B(a[49]), .Z(n2073) );
  NANDN U2165 ( .A(n37), .B(n2073), .Z(n2033) );
  AND U2166 ( .A(n2034), .B(n2033), .Z(n2077) );
  AND U2167 ( .A(b[7]), .B(a[45]), .Z(n2076) );
  XNOR U2168 ( .A(n2077), .B(n2076), .Z(n2078) );
  XNOR U2169 ( .A(n2079), .B(n2078), .Z(n2084) );
  XOR U2170 ( .A(n2085), .B(n2084), .Z(n2059) );
  NANDN U2171 ( .A(n2036), .B(n2035), .Z(n2040) );
  NANDN U2172 ( .A(n2038), .B(n2037), .Z(n2039) );
  AND U2173 ( .A(n2040), .B(n2039), .Z(n2058) );
  XNOR U2174 ( .A(n2059), .B(n2058), .Z(n2060) );
  NANDN U2175 ( .A(n2042), .B(n2041), .Z(n2046) );
  NAND U2176 ( .A(n2044), .B(n2043), .Z(n2045) );
  NAND U2177 ( .A(n2046), .B(n2045), .Z(n2061) );
  XNOR U2178 ( .A(n2060), .B(n2061), .Z(n2052) );
  XNOR U2179 ( .A(n2053), .B(n2052), .Z(n2054) );
  XNOR U2180 ( .A(n2055), .B(n2054), .Z(n2088) );
  XNOR U2181 ( .A(sreg[109]), .B(n2088), .Z(n2090) );
  NANDN U2182 ( .A(sreg[108]), .B(n2047), .Z(n2051) );
  NAND U2183 ( .A(n2049), .B(n2048), .Z(n2050) );
  NAND U2184 ( .A(n2051), .B(n2050), .Z(n2089) );
  XNOR U2185 ( .A(n2090), .B(n2089), .Z(c[109]) );
  NANDN U2186 ( .A(n2053), .B(n2052), .Z(n2057) );
  NANDN U2187 ( .A(n2055), .B(n2054), .Z(n2056) );
  AND U2188 ( .A(n2057), .B(n2056), .Z(n2096) );
  NANDN U2189 ( .A(n2059), .B(n2058), .Z(n2063) );
  NANDN U2190 ( .A(n2061), .B(n2060), .Z(n2062) );
  AND U2191 ( .A(n2063), .B(n2062), .Z(n2094) );
  NANDN U2192 ( .A(n2629), .B(n2064), .Z(n2066) );
  XOR U2193 ( .A(b[7]), .B(a[48]), .Z(n2105) );
  NANDN U2194 ( .A(n2630), .B(n2105), .Z(n2065) );
  AND U2195 ( .A(n2066), .B(n2065), .Z(n2124) );
  NANDN U2196 ( .A(n2483), .B(n2067), .Z(n2069) );
  XOR U2197 ( .A(b[3]), .B(a[52]), .Z(n2108) );
  NANDN U2198 ( .A(n2484), .B(n2108), .Z(n2068) );
  NAND U2199 ( .A(n2069), .B(n2068), .Z(n2123) );
  XNOR U2200 ( .A(n2124), .B(n2123), .Z(n2126) );
  NAND U2201 ( .A(b[0]), .B(a[54]), .Z(n2070) );
  XNOR U2202 ( .A(b[1]), .B(n2070), .Z(n2072) );
  NANDN U2203 ( .A(b[0]), .B(a[53]), .Z(n2071) );
  NAND U2204 ( .A(n2072), .B(n2071), .Z(n2120) );
  NAND U2205 ( .A(n2633), .B(n2073), .Z(n2075) );
  XOR U2206 ( .A(b[5]), .B(a[50]), .Z(n2114) );
  NANDN U2207 ( .A(n37), .B(n2114), .Z(n2074) );
  AND U2208 ( .A(n2075), .B(n2074), .Z(n2118) );
  AND U2209 ( .A(b[7]), .B(a[46]), .Z(n2117) );
  XNOR U2210 ( .A(n2118), .B(n2117), .Z(n2119) );
  XNOR U2211 ( .A(n2120), .B(n2119), .Z(n2125) );
  XOR U2212 ( .A(n2126), .B(n2125), .Z(n2100) );
  NANDN U2213 ( .A(n2077), .B(n2076), .Z(n2081) );
  NANDN U2214 ( .A(n2079), .B(n2078), .Z(n2080) );
  AND U2215 ( .A(n2081), .B(n2080), .Z(n2099) );
  XNOR U2216 ( .A(n2100), .B(n2099), .Z(n2101) );
  NANDN U2217 ( .A(n2083), .B(n2082), .Z(n2087) );
  NAND U2218 ( .A(n2085), .B(n2084), .Z(n2086) );
  NAND U2219 ( .A(n2087), .B(n2086), .Z(n2102) );
  XNOR U2220 ( .A(n2101), .B(n2102), .Z(n2093) );
  XNOR U2221 ( .A(n2094), .B(n2093), .Z(n2095) );
  XNOR U2222 ( .A(n2096), .B(n2095), .Z(n2129) );
  XNOR U2223 ( .A(sreg[110]), .B(n2129), .Z(n2131) );
  NANDN U2224 ( .A(sreg[109]), .B(n2088), .Z(n2092) );
  NAND U2225 ( .A(n2090), .B(n2089), .Z(n2091) );
  NAND U2226 ( .A(n2092), .B(n2091), .Z(n2130) );
  XNOR U2227 ( .A(n2131), .B(n2130), .Z(c[110]) );
  NANDN U2228 ( .A(n2094), .B(n2093), .Z(n2098) );
  NANDN U2229 ( .A(n2096), .B(n2095), .Z(n2097) );
  AND U2230 ( .A(n2098), .B(n2097), .Z(n2137) );
  NANDN U2231 ( .A(n2100), .B(n2099), .Z(n2104) );
  NANDN U2232 ( .A(n2102), .B(n2101), .Z(n2103) );
  AND U2233 ( .A(n2104), .B(n2103), .Z(n2135) );
  NANDN U2234 ( .A(n2629), .B(n2105), .Z(n2107) );
  XOR U2235 ( .A(b[7]), .B(a[49]), .Z(n2146) );
  NANDN U2236 ( .A(n2630), .B(n2146), .Z(n2106) );
  AND U2237 ( .A(n2107), .B(n2106), .Z(n2165) );
  NANDN U2238 ( .A(n2483), .B(n2108), .Z(n2110) );
  XOR U2239 ( .A(b[3]), .B(a[53]), .Z(n2149) );
  NANDN U2240 ( .A(n2484), .B(n2149), .Z(n2109) );
  NAND U2241 ( .A(n2110), .B(n2109), .Z(n2164) );
  XNOR U2242 ( .A(n2165), .B(n2164), .Z(n2167) );
  NAND U2243 ( .A(b[0]), .B(a[55]), .Z(n2111) );
  XNOR U2244 ( .A(b[1]), .B(n2111), .Z(n2113) );
  NANDN U2245 ( .A(b[0]), .B(a[54]), .Z(n2112) );
  NAND U2246 ( .A(n2113), .B(n2112), .Z(n2161) );
  NAND U2247 ( .A(n2633), .B(n2114), .Z(n2116) );
  XOR U2248 ( .A(b[5]), .B(a[51]), .Z(n2155) );
  NANDN U2249 ( .A(n37), .B(n2155), .Z(n2115) );
  AND U2250 ( .A(n2116), .B(n2115), .Z(n2159) );
  AND U2251 ( .A(b[7]), .B(a[47]), .Z(n2158) );
  XNOR U2252 ( .A(n2159), .B(n2158), .Z(n2160) );
  XNOR U2253 ( .A(n2161), .B(n2160), .Z(n2166) );
  XOR U2254 ( .A(n2167), .B(n2166), .Z(n2141) );
  NANDN U2255 ( .A(n2118), .B(n2117), .Z(n2122) );
  NANDN U2256 ( .A(n2120), .B(n2119), .Z(n2121) );
  AND U2257 ( .A(n2122), .B(n2121), .Z(n2140) );
  XNOR U2258 ( .A(n2141), .B(n2140), .Z(n2142) );
  NANDN U2259 ( .A(n2124), .B(n2123), .Z(n2128) );
  NAND U2260 ( .A(n2126), .B(n2125), .Z(n2127) );
  NAND U2261 ( .A(n2128), .B(n2127), .Z(n2143) );
  XNOR U2262 ( .A(n2142), .B(n2143), .Z(n2134) );
  XNOR U2263 ( .A(n2135), .B(n2134), .Z(n2136) );
  XNOR U2264 ( .A(n2137), .B(n2136), .Z(n2170) );
  XNOR U2265 ( .A(sreg[111]), .B(n2170), .Z(n2172) );
  NANDN U2266 ( .A(sreg[110]), .B(n2129), .Z(n2133) );
  NAND U2267 ( .A(n2131), .B(n2130), .Z(n2132) );
  NAND U2268 ( .A(n2133), .B(n2132), .Z(n2171) );
  XNOR U2269 ( .A(n2172), .B(n2171), .Z(c[111]) );
  NANDN U2270 ( .A(n2135), .B(n2134), .Z(n2139) );
  NANDN U2271 ( .A(n2137), .B(n2136), .Z(n2138) );
  AND U2272 ( .A(n2139), .B(n2138), .Z(n2178) );
  NANDN U2273 ( .A(n2141), .B(n2140), .Z(n2145) );
  NANDN U2274 ( .A(n2143), .B(n2142), .Z(n2144) );
  AND U2275 ( .A(n2145), .B(n2144), .Z(n2176) );
  NANDN U2276 ( .A(n2629), .B(n2146), .Z(n2148) );
  XOR U2277 ( .A(b[7]), .B(a[50]), .Z(n2187) );
  NANDN U2278 ( .A(n2630), .B(n2187), .Z(n2147) );
  AND U2279 ( .A(n2148), .B(n2147), .Z(n2206) );
  NANDN U2280 ( .A(n2483), .B(n2149), .Z(n2151) );
  XOR U2281 ( .A(b[3]), .B(a[54]), .Z(n2190) );
  NANDN U2282 ( .A(n2484), .B(n2190), .Z(n2150) );
  NAND U2283 ( .A(n2151), .B(n2150), .Z(n2205) );
  XNOR U2284 ( .A(n2206), .B(n2205), .Z(n2208) );
  NAND U2285 ( .A(b[0]), .B(a[56]), .Z(n2152) );
  XNOR U2286 ( .A(b[1]), .B(n2152), .Z(n2154) );
  NANDN U2287 ( .A(b[0]), .B(a[55]), .Z(n2153) );
  NAND U2288 ( .A(n2154), .B(n2153), .Z(n2202) );
  NAND U2289 ( .A(n2633), .B(n2155), .Z(n2157) );
  XOR U2290 ( .A(b[5]), .B(a[52]), .Z(n2196) );
  NANDN U2291 ( .A(n37), .B(n2196), .Z(n2156) );
  AND U2292 ( .A(n2157), .B(n2156), .Z(n2200) );
  AND U2293 ( .A(b[7]), .B(a[48]), .Z(n2199) );
  XNOR U2294 ( .A(n2200), .B(n2199), .Z(n2201) );
  XNOR U2295 ( .A(n2202), .B(n2201), .Z(n2207) );
  XOR U2296 ( .A(n2208), .B(n2207), .Z(n2182) );
  NANDN U2297 ( .A(n2159), .B(n2158), .Z(n2163) );
  NANDN U2298 ( .A(n2161), .B(n2160), .Z(n2162) );
  AND U2299 ( .A(n2163), .B(n2162), .Z(n2181) );
  XNOR U2300 ( .A(n2182), .B(n2181), .Z(n2183) );
  NANDN U2301 ( .A(n2165), .B(n2164), .Z(n2169) );
  NAND U2302 ( .A(n2167), .B(n2166), .Z(n2168) );
  NAND U2303 ( .A(n2169), .B(n2168), .Z(n2184) );
  XNOR U2304 ( .A(n2183), .B(n2184), .Z(n2175) );
  XNOR U2305 ( .A(n2176), .B(n2175), .Z(n2177) );
  XNOR U2306 ( .A(n2178), .B(n2177), .Z(n2211) );
  XNOR U2307 ( .A(sreg[112]), .B(n2211), .Z(n2213) );
  NANDN U2308 ( .A(sreg[111]), .B(n2170), .Z(n2174) );
  NAND U2309 ( .A(n2172), .B(n2171), .Z(n2173) );
  NAND U2310 ( .A(n2174), .B(n2173), .Z(n2212) );
  XNOR U2311 ( .A(n2213), .B(n2212), .Z(c[112]) );
  NANDN U2312 ( .A(n2176), .B(n2175), .Z(n2180) );
  NANDN U2313 ( .A(n2178), .B(n2177), .Z(n2179) );
  AND U2314 ( .A(n2180), .B(n2179), .Z(n2219) );
  NANDN U2315 ( .A(n2182), .B(n2181), .Z(n2186) );
  NANDN U2316 ( .A(n2184), .B(n2183), .Z(n2185) );
  AND U2317 ( .A(n2186), .B(n2185), .Z(n2217) );
  NANDN U2318 ( .A(n2629), .B(n2187), .Z(n2189) );
  XOR U2319 ( .A(b[7]), .B(a[51]), .Z(n2228) );
  NANDN U2320 ( .A(n2630), .B(n2228), .Z(n2188) );
  AND U2321 ( .A(n2189), .B(n2188), .Z(n2247) );
  NANDN U2322 ( .A(n2483), .B(n2190), .Z(n2192) );
  XOR U2323 ( .A(b[3]), .B(a[55]), .Z(n2231) );
  NANDN U2324 ( .A(n2484), .B(n2231), .Z(n2191) );
  NAND U2325 ( .A(n2192), .B(n2191), .Z(n2246) );
  XNOR U2326 ( .A(n2247), .B(n2246), .Z(n2249) );
  NAND U2327 ( .A(b[0]), .B(a[57]), .Z(n2193) );
  XNOR U2328 ( .A(b[1]), .B(n2193), .Z(n2195) );
  NANDN U2329 ( .A(b[0]), .B(a[56]), .Z(n2194) );
  NAND U2330 ( .A(n2195), .B(n2194), .Z(n2243) );
  NAND U2331 ( .A(n2633), .B(n2196), .Z(n2198) );
  XOR U2332 ( .A(b[5]), .B(a[53]), .Z(n2237) );
  NANDN U2333 ( .A(n37), .B(n2237), .Z(n2197) );
  AND U2334 ( .A(n2198), .B(n2197), .Z(n2241) );
  AND U2335 ( .A(b[7]), .B(a[49]), .Z(n2240) );
  XNOR U2336 ( .A(n2241), .B(n2240), .Z(n2242) );
  XNOR U2337 ( .A(n2243), .B(n2242), .Z(n2248) );
  XOR U2338 ( .A(n2249), .B(n2248), .Z(n2223) );
  NANDN U2339 ( .A(n2200), .B(n2199), .Z(n2204) );
  NANDN U2340 ( .A(n2202), .B(n2201), .Z(n2203) );
  AND U2341 ( .A(n2204), .B(n2203), .Z(n2222) );
  XNOR U2342 ( .A(n2223), .B(n2222), .Z(n2224) );
  NANDN U2343 ( .A(n2206), .B(n2205), .Z(n2210) );
  NAND U2344 ( .A(n2208), .B(n2207), .Z(n2209) );
  NAND U2345 ( .A(n2210), .B(n2209), .Z(n2225) );
  XNOR U2346 ( .A(n2224), .B(n2225), .Z(n2216) );
  XNOR U2347 ( .A(n2217), .B(n2216), .Z(n2218) );
  XNOR U2348 ( .A(n2219), .B(n2218), .Z(n2252) );
  XNOR U2349 ( .A(sreg[113]), .B(n2252), .Z(n2254) );
  NANDN U2350 ( .A(sreg[112]), .B(n2211), .Z(n2215) );
  NAND U2351 ( .A(n2213), .B(n2212), .Z(n2214) );
  NAND U2352 ( .A(n2215), .B(n2214), .Z(n2253) );
  XNOR U2353 ( .A(n2254), .B(n2253), .Z(c[113]) );
  NANDN U2354 ( .A(n2217), .B(n2216), .Z(n2221) );
  NANDN U2355 ( .A(n2219), .B(n2218), .Z(n2220) );
  AND U2356 ( .A(n2221), .B(n2220), .Z(n2260) );
  NANDN U2357 ( .A(n2223), .B(n2222), .Z(n2227) );
  NANDN U2358 ( .A(n2225), .B(n2224), .Z(n2226) );
  AND U2359 ( .A(n2227), .B(n2226), .Z(n2258) );
  NANDN U2360 ( .A(n2629), .B(n2228), .Z(n2230) );
  XOR U2361 ( .A(b[7]), .B(a[52]), .Z(n2269) );
  NANDN U2362 ( .A(n2630), .B(n2269), .Z(n2229) );
  AND U2363 ( .A(n2230), .B(n2229), .Z(n2288) );
  NANDN U2364 ( .A(n2483), .B(n2231), .Z(n2233) );
  XOR U2365 ( .A(b[3]), .B(a[56]), .Z(n2272) );
  NANDN U2366 ( .A(n2484), .B(n2272), .Z(n2232) );
  NAND U2367 ( .A(n2233), .B(n2232), .Z(n2287) );
  XNOR U2368 ( .A(n2288), .B(n2287), .Z(n2290) );
  NAND U2369 ( .A(b[0]), .B(a[58]), .Z(n2234) );
  XNOR U2370 ( .A(b[1]), .B(n2234), .Z(n2236) );
  NANDN U2371 ( .A(b[0]), .B(a[57]), .Z(n2235) );
  NAND U2372 ( .A(n2236), .B(n2235), .Z(n2284) );
  NAND U2373 ( .A(n2633), .B(n2237), .Z(n2239) );
  XOR U2374 ( .A(b[5]), .B(a[54]), .Z(n2275) );
  NANDN U2375 ( .A(n37), .B(n2275), .Z(n2238) );
  AND U2376 ( .A(n2239), .B(n2238), .Z(n2282) );
  AND U2377 ( .A(b[7]), .B(a[50]), .Z(n2281) );
  XNOR U2378 ( .A(n2282), .B(n2281), .Z(n2283) );
  XNOR U2379 ( .A(n2284), .B(n2283), .Z(n2289) );
  XOR U2380 ( .A(n2290), .B(n2289), .Z(n2264) );
  NANDN U2381 ( .A(n2241), .B(n2240), .Z(n2245) );
  NANDN U2382 ( .A(n2243), .B(n2242), .Z(n2244) );
  AND U2383 ( .A(n2245), .B(n2244), .Z(n2263) );
  XNOR U2384 ( .A(n2264), .B(n2263), .Z(n2265) );
  NANDN U2385 ( .A(n2247), .B(n2246), .Z(n2251) );
  NAND U2386 ( .A(n2249), .B(n2248), .Z(n2250) );
  NAND U2387 ( .A(n2251), .B(n2250), .Z(n2266) );
  XNOR U2388 ( .A(n2265), .B(n2266), .Z(n2257) );
  XNOR U2389 ( .A(n2258), .B(n2257), .Z(n2259) );
  XNOR U2390 ( .A(n2260), .B(n2259), .Z(n2293) );
  XNOR U2391 ( .A(sreg[114]), .B(n2293), .Z(n2295) );
  NANDN U2392 ( .A(sreg[113]), .B(n2252), .Z(n2256) );
  NAND U2393 ( .A(n2254), .B(n2253), .Z(n2255) );
  NAND U2394 ( .A(n2256), .B(n2255), .Z(n2294) );
  XNOR U2395 ( .A(n2295), .B(n2294), .Z(c[114]) );
  NANDN U2396 ( .A(n2258), .B(n2257), .Z(n2262) );
  NANDN U2397 ( .A(n2260), .B(n2259), .Z(n2261) );
  AND U2398 ( .A(n2262), .B(n2261), .Z(n2301) );
  NANDN U2399 ( .A(n2264), .B(n2263), .Z(n2268) );
  NANDN U2400 ( .A(n2266), .B(n2265), .Z(n2267) );
  AND U2401 ( .A(n2268), .B(n2267), .Z(n2299) );
  NANDN U2402 ( .A(n2629), .B(n2269), .Z(n2271) );
  XOR U2403 ( .A(b[7]), .B(a[53]), .Z(n2310) );
  NANDN U2404 ( .A(n2630), .B(n2310), .Z(n2270) );
  AND U2405 ( .A(n2271), .B(n2270), .Z(n2329) );
  NANDN U2406 ( .A(n2483), .B(n2272), .Z(n2274) );
  XOR U2407 ( .A(b[3]), .B(a[57]), .Z(n2313) );
  NANDN U2408 ( .A(n2484), .B(n2313), .Z(n2273) );
  NAND U2409 ( .A(n2274), .B(n2273), .Z(n2328) );
  XNOR U2410 ( .A(n2329), .B(n2328), .Z(n2331) );
  NAND U2411 ( .A(n2633), .B(n2275), .Z(n2277) );
  XOR U2412 ( .A(b[5]), .B(a[55]), .Z(n2319) );
  NANDN U2413 ( .A(n37), .B(n2319), .Z(n2276) );
  AND U2414 ( .A(n2277), .B(n2276), .Z(n2323) );
  AND U2415 ( .A(b[7]), .B(a[51]), .Z(n2322) );
  XNOR U2416 ( .A(n2323), .B(n2322), .Z(n2324) );
  NAND U2417 ( .A(b[0]), .B(a[59]), .Z(n2278) );
  XNOR U2418 ( .A(b[1]), .B(n2278), .Z(n2280) );
  NANDN U2419 ( .A(b[0]), .B(a[58]), .Z(n2279) );
  NAND U2420 ( .A(n2280), .B(n2279), .Z(n2325) );
  XNOR U2421 ( .A(n2324), .B(n2325), .Z(n2330) );
  XOR U2422 ( .A(n2331), .B(n2330), .Z(n2305) );
  NANDN U2423 ( .A(n2282), .B(n2281), .Z(n2286) );
  NANDN U2424 ( .A(n2284), .B(n2283), .Z(n2285) );
  AND U2425 ( .A(n2286), .B(n2285), .Z(n2304) );
  XNOR U2426 ( .A(n2305), .B(n2304), .Z(n2306) );
  NANDN U2427 ( .A(n2288), .B(n2287), .Z(n2292) );
  NAND U2428 ( .A(n2290), .B(n2289), .Z(n2291) );
  NAND U2429 ( .A(n2292), .B(n2291), .Z(n2307) );
  XNOR U2430 ( .A(n2306), .B(n2307), .Z(n2298) );
  XNOR U2431 ( .A(n2299), .B(n2298), .Z(n2300) );
  XNOR U2432 ( .A(n2301), .B(n2300), .Z(n2334) );
  XNOR U2433 ( .A(sreg[115]), .B(n2334), .Z(n2336) );
  NANDN U2434 ( .A(sreg[114]), .B(n2293), .Z(n2297) );
  NAND U2435 ( .A(n2295), .B(n2294), .Z(n2296) );
  NAND U2436 ( .A(n2297), .B(n2296), .Z(n2335) );
  XNOR U2437 ( .A(n2336), .B(n2335), .Z(c[115]) );
  NANDN U2438 ( .A(n2299), .B(n2298), .Z(n2303) );
  NANDN U2439 ( .A(n2301), .B(n2300), .Z(n2302) );
  AND U2440 ( .A(n2303), .B(n2302), .Z(n2342) );
  NANDN U2441 ( .A(n2305), .B(n2304), .Z(n2309) );
  NANDN U2442 ( .A(n2307), .B(n2306), .Z(n2308) );
  AND U2443 ( .A(n2309), .B(n2308), .Z(n2340) );
  NANDN U2444 ( .A(n2629), .B(n2310), .Z(n2312) );
  XOR U2445 ( .A(b[7]), .B(a[54]), .Z(n2351) );
  NANDN U2446 ( .A(n2630), .B(n2351), .Z(n2311) );
  AND U2447 ( .A(n2312), .B(n2311), .Z(n2370) );
  NANDN U2448 ( .A(n2483), .B(n2313), .Z(n2315) );
  XOR U2449 ( .A(b[3]), .B(a[58]), .Z(n2354) );
  NANDN U2450 ( .A(n2484), .B(n2354), .Z(n2314) );
  NAND U2451 ( .A(n2315), .B(n2314), .Z(n2369) );
  XNOR U2452 ( .A(n2370), .B(n2369), .Z(n2372) );
  NAND U2453 ( .A(b[0]), .B(a[60]), .Z(n2316) );
  XNOR U2454 ( .A(b[1]), .B(n2316), .Z(n2318) );
  NANDN U2455 ( .A(b[0]), .B(a[59]), .Z(n2317) );
  NAND U2456 ( .A(n2318), .B(n2317), .Z(n2366) );
  NAND U2457 ( .A(n2633), .B(n2319), .Z(n2321) );
  XOR U2458 ( .A(b[5]), .B(a[56]), .Z(n2357) );
  NANDN U2459 ( .A(n37), .B(n2357), .Z(n2320) );
  AND U2460 ( .A(n2321), .B(n2320), .Z(n2364) );
  AND U2461 ( .A(b[7]), .B(a[52]), .Z(n2363) );
  XNOR U2462 ( .A(n2364), .B(n2363), .Z(n2365) );
  XNOR U2463 ( .A(n2366), .B(n2365), .Z(n2371) );
  XOR U2464 ( .A(n2372), .B(n2371), .Z(n2346) );
  NANDN U2465 ( .A(n2323), .B(n2322), .Z(n2327) );
  NANDN U2466 ( .A(n2325), .B(n2324), .Z(n2326) );
  AND U2467 ( .A(n2327), .B(n2326), .Z(n2345) );
  XNOR U2468 ( .A(n2346), .B(n2345), .Z(n2347) );
  NANDN U2469 ( .A(n2329), .B(n2328), .Z(n2333) );
  NAND U2470 ( .A(n2331), .B(n2330), .Z(n2332) );
  NAND U2471 ( .A(n2333), .B(n2332), .Z(n2348) );
  XNOR U2472 ( .A(n2347), .B(n2348), .Z(n2339) );
  XNOR U2473 ( .A(n2340), .B(n2339), .Z(n2341) );
  XNOR U2474 ( .A(n2342), .B(n2341), .Z(n2375) );
  XNOR U2475 ( .A(sreg[116]), .B(n2375), .Z(n2377) );
  NANDN U2476 ( .A(sreg[115]), .B(n2334), .Z(n2338) );
  NAND U2477 ( .A(n2336), .B(n2335), .Z(n2337) );
  NAND U2478 ( .A(n2338), .B(n2337), .Z(n2376) );
  XNOR U2479 ( .A(n2377), .B(n2376), .Z(c[116]) );
  NANDN U2480 ( .A(n2340), .B(n2339), .Z(n2344) );
  NANDN U2481 ( .A(n2342), .B(n2341), .Z(n2343) );
  AND U2482 ( .A(n2344), .B(n2343), .Z(n2383) );
  NANDN U2483 ( .A(n2346), .B(n2345), .Z(n2350) );
  NANDN U2484 ( .A(n2348), .B(n2347), .Z(n2349) );
  AND U2485 ( .A(n2350), .B(n2349), .Z(n2381) );
  NANDN U2486 ( .A(n2629), .B(n2351), .Z(n2353) );
  XOR U2487 ( .A(b[7]), .B(a[55]), .Z(n2392) );
  NANDN U2488 ( .A(n2630), .B(n2392), .Z(n2352) );
  AND U2489 ( .A(n2353), .B(n2352), .Z(n2411) );
  NANDN U2490 ( .A(n2483), .B(n2354), .Z(n2356) );
  XOR U2491 ( .A(b[3]), .B(a[59]), .Z(n2395) );
  NANDN U2492 ( .A(n2484), .B(n2395), .Z(n2355) );
  NAND U2493 ( .A(n2356), .B(n2355), .Z(n2410) );
  XNOR U2494 ( .A(n2411), .B(n2410), .Z(n2413) );
  NAND U2495 ( .A(n2633), .B(n2357), .Z(n2359) );
  XOR U2496 ( .A(b[5]), .B(a[57]), .Z(n2398) );
  NANDN U2497 ( .A(n37), .B(n2398), .Z(n2358) );
  AND U2498 ( .A(n2359), .B(n2358), .Z(n2405) );
  AND U2499 ( .A(b[7]), .B(a[53]), .Z(n2404) );
  XNOR U2500 ( .A(n2405), .B(n2404), .Z(n2406) );
  NAND U2501 ( .A(b[0]), .B(a[61]), .Z(n2360) );
  XNOR U2502 ( .A(b[1]), .B(n2360), .Z(n2362) );
  NANDN U2503 ( .A(b[0]), .B(a[60]), .Z(n2361) );
  NAND U2504 ( .A(n2362), .B(n2361), .Z(n2407) );
  XNOR U2505 ( .A(n2406), .B(n2407), .Z(n2412) );
  XOR U2506 ( .A(n2413), .B(n2412), .Z(n2387) );
  NANDN U2507 ( .A(n2364), .B(n2363), .Z(n2368) );
  NANDN U2508 ( .A(n2366), .B(n2365), .Z(n2367) );
  AND U2509 ( .A(n2368), .B(n2367), .Z(n2386) );
  XNOR U2510 ( .A(n2387), .B(n2386), .Z(n2388) );
  NANDN U2511 ( .A(n2370), .B(n2369), .Z(n2374) );
  NAND U2512 ( .A(n2372), .B(n2371), .Z(n2373) );
  NAND U2513 ( .A(n2374), .B(n2373), .Z(n2389) );
  XNOR U2514 ( .A(n2388), .B(n2389), .Z(n2380) );
  XNOR U2515 ( .A(n2381), .B(n2380), .Z(n2382) );
  XNOR U2516 ( .A(n2383), .B(n2382), .Z(n2416) );
  XNOR U2517 ( .A(sreg[117]), .B(n2416), .Z(n2418) );
  NANDN U2518 ( .A(sreg[116]), .B(n2375), .Z(n2379) );
  NAND U2519 ( .A(n2377), .B(n2376), .Z(n2378) );
  NAND U2520 ( .A(n2379), .B(n2378), .Z(n2417) );
  XNOR U2521 ( .A(n2418), .B(n2417), .Z(c[117]) );
  NANDN U2522 ( .A(n2381), .B(n2380), .Z(n2385) );
  NANDN U2523 ( .A(n2383), .B(n2382), .Z(n2384) );
  AND U2524 ( .A(n2385), .B(n2384), .Z(n2424) );
  NANDN U2525 ( .A(n2387), .B(n2386), .Z(n2391) );
  NANDN U2526 ( .A(n2389), .B(n2388), .Z(n2390) );
  AND U2527 ( .A(n2391), .B(n2390), .Z(n2422) );
  NANDN U2528 ( .A(n2629), .B(n2392), .Z(n2394) );
  XOR U2529 ( .A(b[7]), .B(a[56]), .Z(n2439) );
  NANDN U2530 ( .A(n2630), .B(n2439), .Z(n2393) );
  AND U2531 ( .A(n2394), .B(n2393), .Z(n2428) );
  NANDN U2532 ( .A(n2483), .B(n2395), .Z(n2397) );
  XOR U2533 ( .A(b[3]), .B(a[60]), .Z(n2442) );
  NANDN U2534 ( .A(n2484), .B(n2442), .Z(n2396) );
  NAND U2535 ( .A(n2397), .B(n2396), .Z(n2427) );
  NAND U2536 ( .A(n2633), .B(n2398), .Z(n2400) );
  XOR U2537 ( .A(b[5]), .B(a[58]), .Z(n2445) );
  NANDN U2538 ( .A(n37), .B(n2445), .Z(n2399) );
  AND U2539 ( .A(n2400), .B(n2399), .Z(n2434) );
  AND U2540 ( .A(b[7]), .B(a[54]), .Z(n2433) );
  NAND U2541 ( .A(b[0]), .B(a[62]), .Z(n2401) );
  XNOR U2542 ( .A(b[1]), .B(n2401), .Z(n2403) );
  NANDN U2543 ( .A(b[0]), .B(a[61]), .Z(n2402) );
  NAND U2544 ( .A(n2403), .B(n2402), .Z(n2436) );
  XNOR U2545 ( .A(n2435), .B(n2436), .Z(n2429) );
  XOR U2546 ( .A(n2430), .B(n2429), .Z(n2452) );
  NANDN U2547 ( .A(n2405), .B(n2404), .Z(n2409) );
  NANDN U2548 ( .A(n2407), .B(n2406), .Z(n2408) );
  AND U2549 ( .A(n2409), .B(n2408), .Z(n2451) );
  NANDN U2550 ( .A(n2411), .B(n2410), .Z(n2415) );
  NAND U2551 ( .A(n2413), .B(n2412), .Z(n2414) );
  NAND U2552 ( .A(n2415), .B(n2414), .Z(n2454) );
  XNOR U2553 ( .A(n2422), .B(n2421), .Z(n2423) );
  XNOR U2554 ( .A(n2424), .B(n2423), .Z(n2457) );
  XNOR U2555 ( .A(sreg[118]), .B(n2457), .Z(n2459) );
  NANDN U2556 ( .A(sreg[117]), .B(n2416), .Z(n2420) );
  NAND U2557 ( .A(n2418), .B(n2417), .Z(n2419) );
  NAND U2558 ( .A(n2420), .B(n2419), .Z(n2458) );
  XNOR U2559 ( .A(n2459), .B(n2458), .Z(c[118]) );
  NANDN U2560 ( .A(n2422), .B(n2421), .Z(n2426) );
  NANDN U2561 ( .A(n2424), .B(n2423), .Z(n2425) );
  AND U2562 ( .A(n2426), .B(n2425), .Z(n2470) );
  NANDN U2563 ( .A(n2428), .B(n2427), .Z(n2432) );
  NAND U2564 ( .A(n2430), .B(n2429), .Z(n2431) );
  AND U2565 ( .A(n2432), .B(n2431), .Z(n2476) );
  NANDN U2566 ( .A(n2434), .B(n2433), .Z(n2438) );
  NANDN U2567 ( .A(n2436), .B(n2435), .Z(n2437) );
  AND U2568 ( .A(n2438), .B(n2437), .Z(n2474) );
  NANDN U2569 ( .A(n2629), .B(n2439), .Z(n2441) );
  XOR U2570 ( .A(b[7]), .B(a[57]), .Z(n2479) );
  NANDN U2571 ( .A(n2630), .B(n2479), .Z(n2440) );
  AND U2572 ( .A(n2441), .B(n2440), .Z(n2499) );
  NANDN U2573 ( .A(n2483), .B(n2442), .Z(n2444) );
  XOR U2574 ( .A(b[3]), .B(a[61]), .Z(n2482) );
  NANDN U2575 ( .A(n2484), .B(n2482), .Z(n2443) );
  AND U2576 ( .A(n2444), .B(n2443), .Z(n2497) );
  NAND U2577 ( .A(n2633), .B(n2445), .Z(n2447) );
  XOR U2578 ( .A(b[5]), .B(a[59]), .Z(n2487) );
  NANDN U2579 ( .A(n37), .B(n2487), .Z(n2446) );
  AND U2580 ( .A(n2447), .B(n2446), .Z(n2491) );
  AND U2581 ( .A(b[7]), .B(a[55]), .Z(n2490) );
  NAND U2582 ( .A(b[0]), .B(a[63]), .Z(n2448) );
  XNOR U2583 ( .A(b[1]), .B(n2448), .Z(n2450) );
  NANDN U2584 ( .A(b[0]), .B(a[62]), .Z(n2449) );
  NAND U2585 ( .A(n2450), .B(n2449), .Z(n2493) );
  XNOR U2586 ( .A(n2492), .B(n2493), .Z(n2496) );
  NANDN U2587 ( .A(n2452), .B(n2451), .Z(n2456) );
  NANDN U2588 ( .A(n2454), .B(n2453), .Z(n2455) );
  NAND U2589 ( .A(n2456), .B(n2455), .Z(n2467) );
  XOR U2590 ( .A(n2468), .B(n2467), .Z(n2469) );
  XNOR U2591 ( .A(sreg[119]), .B(n2462), .Z(n2464) );
  NANDN U2592 ( .A(sreg[118]), .B(n2457), .Z(n2461) );
  NAND U2593 ( .A(n2459), .B(n2458), .Z(n2460) );
  NAND U2594 ( .A(n2461), .B(n2460), .Z(n2463) );
  XNOR U2595 ( .A(n2464), .B(n2463), .Z(c[119]) );
  NANDN U2596 ( .A(sreg[119]), .B(n2462), .Z(n2466) );
  NAND U2597 ( .A(n2464), .B(n2463), .Z(n2465) );
  AND U2598 ( .A(n2466), .B(n2465), .Z(n2503) );
  NAND U2599 ( .A(n2468), .B(n2467), .Z(n2472) );
  NANDN U2600 ( .A(n2470), .B(n2469), .Z(n2471) );
  AND U2601 ( .A(n2472), .B(n2471), .Z(n2507) );
  NANDN U2602 ( .A(n2474), .B(n2473), .Z(n2478) );
  NANDN U2603 ( .A(n2476), .B(n2475), .Z(n2477) );
  AND U2604 ( .A(n2478), .B(n2477), .Z(n2505) );
  NANDN U2605 ( .A(n2629), .B(n2479), .Z(n2481) );
  XOR U2606 ( .A(b[7]), .B(a[58]), .Z(n2522) );
  NANDN U2607 ( .A(n2630), .B(n2522), .Z(n2480) );
  AND U2608 ( .A(n2481), .B(n2480), .Z(n2534) );
  NANDN U2609 ( .A(n2483), .B(n2482), .Z(n2486) );
  XOR U2610 ( .A(b[3]), .B(a[62]), .Z(n2528) );
  NANDN U2611 ( .A(n2484), .B(n2528), .Z(n2485) );
  AND U2612 ( .A(n2486), .B(n2485), .Z(n2532) );
  NAND U2613 ( .A(n2633), .B(n2487), .Z(n2489) );
  XOR U2614 ( .A(b[5]), .B(a[60]), .Z(n2525) );
  NANDN U2615 ( .A(n37), .B(n2525), .Z(n2488) );
  AND U2616 ( .A(n2489), .B(n2488), .Z(n2517) );
  AND U2617 ( .A(b[7]), .B(a[56]), .Z(n2516) );
  NANDN U2618 ( .A(n2491), .B(n2490), .Z(n2495) );
  NANDN U2619 ( .A(n2493), .B(n2492), .Z(n2494) );
  AND U2620 ( .A(n2495), .B(n2494), .Z(n2511) );
  XOR U2621 ( .A(n2510), .B(n2511), .Z(n2512) );
  NANDN U2622 ( .A(n2497), .B(n2496), .Z(n2501) );
  NANDN U2623 ( .A(n2499), .B(n2498), .Z(n2500) );
  NAND U2624 ( .A(n2501), .B(n2500), .Z(n2513) );
  XOR U2625 ( .A(n2505), .B(n2504), .Z(n2506) );
  XOR U2626 ( .A(n2507), .B(n2506), .Z(n2502) );
  XOR U2627 ( .A(n2503), .B(n2502), .Z(c[120]) );
  AND U2628 ( .A(n2503), .B(n2502), .Z(n2538) );
  NAND U2629 ( .A(n2505), .B(n2504), .Z(n2509) );
  NANDN U2630 ( .A(n2507), .B(n2506), .Z(n2508) );
  AND U2631 ( .A(n2509), .B(n2508), .Z(n2542) );
  NAND U2632 ( .A(n2511), .B(n2510), .Z(n2515) );
  NANDN U2633 ( .A(n2513), .B(n2512), .Z(n2514) );
  AND U2634 ( .A(n2515), .B(n2514), .Z(n2540) );
  NANDN U2635 ( .A(n2517), .B(n2516), .Z(n2521) );
  NANDN U2636 ( .A(n2519), .B(n2518), .Z(n2520) );
  AND U2637 ( .A(n2521), .B(n2520), .Z(n2546) );
  NANDN U2638 ( .A(n2629), .B(n2522), .Z(n2524) );
  XOR U2639 ( .A(b[7]), .B(a[59]), .Z(n2560) );
  NANDN U2640 ( .A(n2630), .B(n2560), .Z(n2523) );
  AND U2641 ( .A(n2524), .B(n2523), .Z(n2568) );
  NAND U2642 ( .A(b[7]), .B(a[57]), .Z(n2625) );
  NAND U2643 ( .A(n2633), .B(n2525), .Z(n2527) );
  XOR U2644 ( .A(b[5]), .B(a[61]), .Z(n2563) );
  NANDN U2645 ( .A(n37), .B(n2563), .Z(n2526) );
  NAND U2646 ( .A(n2527), .B(n2526), .Z(n2566) );
  XOR U2647 ( .A(n2625), .B(n2566), .Z(n2567) );
  NAND U2648 ( .A(n2556), .B(n2528), .Z(n2530) );
  XNOR U2649 ( .A(b[3]), .B(a[63]), .Z(n2557) );
  NANDN U2650 ( .A(n2557), .B(n36), .Z(n2529) );
  NAND U2651 ( .A(n2530), .B(n2529), .Z(n2551) );
  XOR U2652 ( .A(n2552), .B(n2553), .Z(n2545) );
  XOR U2653 ( .A(n2546), .B(n2545), .Z(n2547) );
  NANDN U2654 ( .A(n2532), .B(n2531), .Z(n2536) );
  NANDN U2655 ( .A(n2534), .B(n2533), .Z(n2535) );
  NAND U2656 ( .A(n2536), .B(n2535), .Z(n2548) );
  XOR U2657 ( .A(n2542), .B(n2541), .Z(n2537) );
  XOR U2658 ( .A(n2538), .B(n2537), .Z(c[121]) );
  AND U2659 ( .A(n2538), .B(n2537), .Z(n2572) );
  NANDN U2660 ( .A(n2540), .B(n2539), .Z(n2544) );
  NANDN U2661 ( .A(n2542), .B(n2541), .Z(n2543) );
  AND U2662 ( .A(n2544), .B(n2543), .Z(n2576) );
  NAND U2663 ( .A(n2546), .B(n2545), .Z(n2550) );
  NANDN U2664 ( .A(n2548), .B(n2547), .Z(n2549) );
  AND U2665 ( .A(n2550), .B(n2549), .Z(n2574) );
  NANDN U2666 ( .A(n2551), .B(b[1]), .Z(n2555) );
  NAND U2667 ( .A(n2553), .B(n2552), .Z(n2554) );
  AND U2668 ( .A(n2555), .B(n2554), .Z(n2582) );
  NANDN U2669 ( .A(n2557), .B(n2556), .Z(n2558) );
  AND U2670 ( .A(n2559), .B(n2558), .Z(n2591) );
  AND U2671 ( .A(b[7]), .B(a[58]), .Z(n2590) );
  XNOR U2672 ( .A(n2591), .B(n2590), .Z(n2592) );
  XOR U2673 ( .A(n2625), .B(n2592), .Z(n2599) );
  NANDN U2674 ( .A(n2629), .B(n2560), .Z(n2562) );
  XOR U2675 ( .A(b[7]), .B(a[60]), .Z(n2585) );
  NANDN U2676 ( .A(n2630), .B(n2585), .Z(n2561) );
  AND U2677 ( .A(n2562), .B(n2561), .Z(n2597) );
  NAND U2678 ( .A(n2633), .B(n2563), .Z(n2565) );
  XOR U2679 ( .A(b[5]), .B(a[62]), .Z(n2588) );
  NANDN U2680 ( .A(n37), .B(n2588), .Z(n2564) );
  NAND U2681 ( .A(n2565), .B(n2564), .Z(n2596) );
  XOR U2682 ( .A(n2599), .B(n2598), .Z(n2580) );
  IV U2683 ( .A(n2625), .Z(n2593) );
  NANDN U2684 ( .A(n2593), .B(n2566), .Z(n2570) );
  NANDN U2685 ( .A(n2568), .B(n2567), .Z(n2569) );
  AND U2686 ( .A(n2570), .B(n2569), .Z(n2579) );
  XOR U2687 ( .A(n2576), .B(n2575), .Z(n2571) );
  XOR U2688 ( .A(n2572), .B(n2571), .Z(c[122]) );
  AND U2689 ( .A(n2572), .B(n2571), .Z(n2603) );
  NANDN U2690 ( .A(n2574), .B(n2573), .Z(n2578) );
  NANDN U2691 ( .A(n2576), .B(n2575), .Z(n2577) );
  AND U2692 ( .A(n2578), .B(n2577), .Z(n2607) );
  NANDN U2693 ( .A(n2580), .B(n2579), .Z(n2584) );
  NANDN U2694 ( .A(n2582), .B(n2581), .Z(n2583) );
  AND U2695 ( .A(n2584), .B(n2583), .Z(n2605) );
  NANDN U2696 ( .A(n2629), .B(n2585), .Z(n2587) );
  XOR U2697 ( .A(b[7]), .B(a[61]), .Z(n2628) );
  NANDN U2698 ( .A(n2630), .B(n2628), .Z(n2586) );
  AND U2699 ( .A(n2587), .B(n2586), .Z(n2617) );
  XOR U2700 ( .A(b[5]), .B(a[63]), .Z(n2634) );
  AND U2701 ( .A(b[7]), .B(a[59]), .Z(n2622) );
  XOR U2702 ( .A(n2622), .B(n2589), .Z(n2624) );
  XOR U2703 ( .A(n2593), .B(n2624), .Z(n2618) );
  XOR U2704 ( .A(n2619), .B(n2618), .Z(n2611) );
  NANDN U2705 ( .A(n2591), .B(n2590), .Z(n2595) );
  NANDN U2706 ( .A(n2593), .B(n2592), .Z(n2594) );
  AND U2707 ( .A(n2595), .B(n2594), .Z(n2610) );
  NANDN U2708 ( .A(n2597), .B(n2596), .Z(n2601) );
  NAND U2709 ( .A(n2599), .B(n2598), .Z(n2600) );
  NAND U2710 ( .A(n2601), .B(n2600), .Z(n2613) );
  XOR U2711 ( .A(n2607), .B(n2606), .Z(n2602) );
  XOR U2712 ( .A(n2603), .B(n2602), .Z(c[123]) );
  AND U2713 ( .A(n2603), .B(n2602), .Z(n2638) );
  NANDN U2714 ( .A(n2605), .B(n2604), .Z(n2609) );
  NANDN U2715 ( .A(n2607), .B(n2606), .Z(n2608) );
  AND U2716 ( .A(n2609), .B(n2608), .Z(n2642) );
  NANDN U2717 ( .A(n2611), .B(n2610), .Z(n2615) );
  NANDN U2718 ( .A(n2613), .B(n2612), .Z(n2614) );
  AND U2719 ( .A(n2615), .B(n2614), .Z(n2640) );
  NANDN U2720 ( .A(n2617), .B(n2616), .Z(n2621) );
  NAND U2721 ( .A(n2619), .B(n2618), .Z(n2620) );
  AND U2722 ( .A(n2621), .B(n2620), .Z(n2648) );
  NANDN U2723 ( .A(n2623), .B(n2622), .Z(n2627) );
  NANDN U2724 ( .A(n2625), .B(n2624), .Z(n2626) );
  AND U2725 ( .A(n2627), .B(n2626), .Z(n2646) );
  NANDN U2726 ( .A(n2629), .B(n2628), .Z(n2632) );
  XOR U2727 ( .A(b[7]), .B(a[62]), .Z(n2657) );
  NANDN U2728 ( .A(n2630), .B(n2657), .Z(n2631) );
  AND U2729 ( .A(n2632), .B(n2631), .Z(n2654) );
  NAND U2730 ( .A(n2634), .B(n2633), .Z(n2635) );
  AND U2731 ( .A(n2636), .B(n2635), .Z(n2652) );
  NAND U2732 ( .A(b[7]), .B(a[60]), .Z(n2663) );
  IV U2733 ( .A(n2663), .Z(n2651) );
  XOR U2734 ( .A(n2652), .B(n2651), .Z(n2653) );
  XOR U2735 ( .A(n2648), .B(n2647), .Z(n2639) );
  XOR U2736 ( .A(n2642), .B(n2641), .Z(n2637) );
  XOR U2737 ( .A(n2638), .B(n2637), .Z(c[124]) );
  AND U2738 ( .A(n2638), .B(n2637), .Z(n2672) );
  NANDN U2739 ( .A(n2640), .B(n2639), .Z(n2644) );
  NANDN U2740 ( .A(n2642), .B(n2641), .Z(n2643) );
  AND U2741 ( .A(n2644), .B(n2643), .Z(n2682) );
  NANDN U2742 ( .A(n2646), .B(n2645), .Z(n2650) );
  NANDN U2743 ( .A(n2648), .B(n2647), .Z(n2649) );
  AND U2744 ( .A(n2650), .B(n2649), .Z(n2680) );
  OR U2745 ( .A(n2652), .B(n2651), .Z(n2656) );
  NANDN U2746 ( .A(n2654), .B(n2653), .Z(n2655) );
  AND U2747 ( .A(n2656), .B(n2655), .Z(n2676) );
  AND U2748 ( .A(b[7]), .B(a[61]), .Z(n2660) );
  XNOR U2749 ( .A(n2661), .B(n2660), .Z(n2662) );
  XOR U2750 ( .A(n2662), .B(n2663), .Z(n2673) );
  NAND U2751 ( .A(n2667), .B(n2657), .Z(n2659) );
  XNOR U2752 ( .A(b[7]), .B(a[63]), .Z(n2668) );
  NANDN U2753 ( .A(n2668), .B(n2666), .Z(n2658) );
  AND U2754 ( .A(n2659), .B(n2658), .Z(n2674) );
  XOR U2755 ( .A(n2673), .B(n2674), .Z(n2675) );
  XOR U2756 ( .A(n2676), .B(n2675), .Z(n2679) );
  XOR U2757 ( .A(n2680), .B(n2679), .Z(n2681) );
  XOR U2758 ( .A(n2682), .B(n2681), .Z(n2671) );
  XOR U2759 ( .A(n2672), .B(n2671), .Z(c[125]) );
  NANDN U2760 ( .A(n2661), .B(n2660), .Z(n2665) );
  NANDN U2761 ( .A(n2663), .B(n2662), .Z(n2664) );
  NAND U2762 ( .A(n2665), .B(n2664), .Z(n2694) );
  NAND U2763 ( .A(b[7]), .B(a[62]), .Z(n2692) );
  NAND U2764 ( .A(b[7]), .B(n2666), .Z(n2670) );
  NANDN U2765 ( .A(n2668), .B(n2667), .Z(n2669) );
  NAND U2766 ( .A(n2670), .B(n2669), .Z(n2691) );
  XNOR U2767 ( .A(n2692), .B(n2691), .Z(n2693) );
  AND U2768 ( .A(n2672), .B(n2671), .Z(n2690) );
  XNOR U2769 ( .A(n2689), .B(n2690), .Z(n2686) );
  NAND U2770 ( .A(n2674), .B(n2673), .Z(n2678) );
  NAND U2771 ( .A(n2676), .B(n2675), .Z(n2677) );
  AND U2772 ( .A(n2678), .B(n2677), .Z(n2688) );
  NAND U2773 ( .A(n2680), .B(n2679), .Z(n2684) );
  NANDN U2774 ( .A(n2682), .B(n2681), .Z(n2683) );
  NAND U2775 ( .A(n2684), .B(n2683), .Z(n2687) );
  XOR U2776 ( .A(n2688), .B(n2687), .Z(n2685) );
  XNOR U2777 ( .A(n2686), .B(n2685), .Z(c[126]) );
endmodule

