
module mult_N64_CC16 ( clk, rst, a, b, c );
  input [63:0] a;
  input [3:0] b;
  output [63:0] c;
  input clk, rst;
  wire   \mult_44/PROD1[3] , \mult_44/SUMB[1][1] , \mult_44/SUMB[1][2] ,
         \mult_44/SUMB[2][1] , \mult_44/SUMB[2][2] , \mult_44/SUMB[3][1] ,
         \mult_44/SUMB[3][2] , \mult_44/SUMB[4][1] , \mult_44/SUMB[4][2] ,
         \mult_44/SUMB[5][1] , \mult_44/SUMB[5][2] , \mult_44/SUMB[6][1] ,
         \mult_44/SUMB[6][2] , \mult_44/SUMB[7][1] , \mult_44/SUMB[7][2] ,
         \mult_44/SUMB[8][1] , \mult_44/SUMB[8][2] , \mult_44/SUMB[9][1] ,
         \mult_44/SUMB[9][2] , \mult_44/SUMB[10][1] , \mult_44/SUMB[10][2] ,
         \mult_44/SUMB[11][1] , \mult_44/SUMB[11][2] , \mult_44/SUMB[12][1] ,
         \mult_44/SUMB[12][2] , \mult_44/SUMB[13][1] , \mult_44/SUMB[13][2] ,
         \mult_44/SUMB[14][1] , \mult_44/SUMB[14][2] , \mult_44/SUMB[15][1] ,
         \mult_44/SUMB[15][2] , \mult_44/SUMB[16][1] , \mult_44/SUMB[16][2] ,
         \mult_44/SUMB[17][1] , \mult_44/SUMB[17][2] , \mult_44/SUMB[18][1] ,
         \mult_44/SUMB[18][2] , \mult_44/SUMB[19][1] , \mult_44/SUMB[19][2] ,
         \mult_44/SUMB[20][1] , \mult_44/SUMB[20][2] , \mult_44/SUMB[21][1] ,
         \mult_44/SUMB[21][2] , \mult_44/SUMB[22][1] , \mult_44/SUMB[22][2] ,
         \mult_44/SUMB[23][1] , \mult_44/SUMB[23][2] , \mult_44/SUMB[24][1] ,
         \mult_44/SUMB[24][2] , \mult_44/SUMB[25][1] , \mult_44/SUMB[25][2] ,
         \mult_44/SUMB[26][1] , \mult_44/SUMB[26][2] , \mult_44/SUMB[27][1] ,
         \mult_44/SUMB[27][2] , \mult_44/SUMB[28][1] , \mult_44/SUMB[28][2] ,
         \mult_44/SUMB[29][1] , \mult_44/SUMB[29][2] , \mult_44/SUMB[30][1] ,
         \mult_44/SUMB[30][2] , \mult_44/SUMB[31][1] , \mult_44/SUMB[31][2] ,
         \mult_44/SUMB[32][1] , \mult_44/SUMB[32][2] , \mult_44/SUMB[33][1] ,
         \mult_44/SUMB[33][2] , \mult_44/SUMB[34][1] , \mult_44/SUMB[34][2] ,
         \mult_44/SUMB[35][1] , \mult_44/SUMB[35][2] , \mult_44/SUMB[36][1] ,
         \mult_44/SUMB[36][2] , \mult_44/SUMB[37][1] , \mult_44/SUMB[37][2] ,
         \mult_44/SUMB[38][1] , \mult_44/SUMB[38][2] , \mult_44/SUMB[39][1] ,
         \mult_44/SUMB[39][2] , \mult_44/SUMB[40][1] , \mult_44/SUMB[40][2] ,
         \mult_44/SUMB[41][1] , \mult_44/SUMB[41][2] , \mult_44/SUMB[42][1] ,
         \mult_44/SUMB[42][2] , \mult_44/SUMB[43][1] , \mult_44/SUMB[43][2] ,
         \mult_44/SUMB[44][1] , \mult_44/SUMB[44][2] , \mult_44/SUMB[45][1] ,
         \mult_44/SUMB[45][2] , \mult_44/SUMB[46][1] , \mult_44/SUMB[46][2] ,
         \mult_44/SUMB[47][1] , \mult_44/SUMB[47][2] , \mult_44/SUMB[48][1] ,
         \mult_44/SUMB[48][2] , \mult_44/SUMB[49][1] , \mult_44/SUMB[49][2] ,
         \mult_44/SUMB[50][1] , \mult_44/SUMB[50][2] , \mult_44/SUMB[51][1] ,
         \mult_44/SUMB[51][2] , \mult_44/SUMB[52][1] , \mult_44/SUMB[52][2] ,
         \mult_44/SUMB[53][1] , \mult_44/SUMB[53][2] , \mult_44/SUMB[54][1] ,
         \mult_44/SUMB[54][2] , \mult_44/SUMB[55][1] , \mult_44/SUMB[55][2] ,
         \mult_44/SUMB[56][1] , \mult_44/SUMB[56][2] , \mult_44/SUMB[57][1] ,
         \mult_44/SUMB[57][2] , \mult_44/SUMB[58][1] , \mult_44/SUMB[58][2] ,
         \mult_44/SUMB[59][1] , \mult_44/SUMB[59][2] , \mult_44/SUMB[60][1] ,
         \mult_44/SUMB[60][2] , \mult_44/SUMB[61][1] , \mult_44/SUMB[61][2] ,
         \mult_44/SUMB[62][1] , \mult_44/SUMB[63][0] , \mult_44/CARRYB[1][0] ,
         \mult_44/CARRYB[1][1] , \mult_44/CARRYB[1][2] ,
         \mult_44/CARRYB[2][0] , \mult_44/CARRYB[2][1] ,
         \mult_44/CARRYB[2][2] , \mult_44/CARRYB[3][0] ,
         \mult_44/CARRYB[3][1] , \mult_44/CARRYB[3][2] ,
         \mult_44/CARRYB[4][0] , \mult_44/CARRYB[4][1] ,
         \mult_44/CARRYB[4][2] , \mult_44/CARRYB[5][0] ,
         \mult_44/CARRYB[5][1] , \mult_44/CARRYB[5][2] ,
         \mult_44/CARRYB[6][0] , \mult_44/CARRYB[6][1] ,
         \mult_44/CARRYB[6][2] , \mult_44/CARRYB[7][0] ,
         \mult_44/CARRYB[7][1] , \mult_44/CARRYB[7][2] ,
         \mult_44/CARRYB[8][0] , \mult_44/CARRYB[8][1] ,
         \mult_44/CARRYB[8][2] , \mult_44/CARRYB[9][0] ,
         \mult_44/CARRYB[9][1] , \mult_44/CARRYB[9][2] ,
         \mult_44/CARRYB[10][0] , \mult_44/CARRYB[10][1] ,
         \mult_44/CARRYB[10][2] , \mult_44/CARRYB[11][0] ,
         \mult_44/CARRYB[11][1] , \mult_44/CARRYB[11][2] ,
         \mult_44/CARRYB[12][0] , \mult_44/CARRYB[12][1] ,
         \mult_44/CARRYB[12][2] , \mult_44/CARRYB[13][0] ,
         \mult_44/CARRYB[13][1] , \mult_44/CARRYB[13][2] ,
         \mult_44/CARRYB[14][0] , \mult_44/CARRYB[14][1] ,
         \mult_44/CARRYB[14][2] , \mult_44/CARRYB[15][0] ,
         \mult_44/CARRYB[15][1] , \mult_44/CARRYB[15][2] ,
         \mult_44/CARRYB[16][0] , \mult_44/CARRYB[16][1] ,
         \mult_44/CARRYB[16][2] , \mult_44/CARRYB[17][0] ,
         \mult_44/CARRYB[17][1] , \mult_44/CARRYB[17][2] ,
         \mult_44/CARRYB[18][0] , \mult_44/CARRYB[18][1] ,
         \mult_44/CARRYB[18][2] , \mult_44/CARRYB[19][0] ,
         \mult_44/CARRYB[19][1] , \mult_44/CARRYB[19][2] ,
         \mult_44/CARRYB[20][0] , \mult_44/CARRYB[20][1] ,
         \mult_44/CARRYB[20][2] , \mult_44/CARRYB[21][0] ,
         \mult_44/CARRYB[21][1] , \mult_44/CARRYB[21][2] ,
         \mult_44/CARRYB[22][0] , \mult_44/CARRYB[22][1] ,
         \mult_44/CARRYB[22][2] , \mult_44/CARRYB[23][0] ,
         \mult_44/CARRYB[23][1] , \mult_44/CARRYB[23][2] ,
         \mult_44/CARRYB[24][0] , \mult_44/CARRYB[24][1] ,
         \mult_44/CARRYB[24][2] , \mult_44/CARRYB[25][0] ,
         \mult_44/CARRYB[25][1] , \mult_44/CARRYB[25][2] ,
         \mult_44/CARRYB[26][0] , \mult_44/CARRYB[26][1] ,
         \mult_44/CARRYB[26][2] , \mult_44/CARRYB[27][0] ,
         \mult_44/CARRYB[27][1] , \mult_44/CARRYB[27][2] ,
         \mult_44/CARRYB[28][0] , \mult_44/CARRYB[28][1] ,
         \mult_44/CARRYB[28][2] , \mult_44/CARRYB[29][0] ,
         \mult_44/CARRYB[29][1] , \mult_44/CARRYB[29][2] ,
         \mult_44/CARRYB[30][0] , \mult_44/CARRYB[30][1] ,
         \mult_44/CARRYB[30][2] , \mult_44/CARRYB[31][0] ,
         \mult_44/CARRYB[31][1] , \mult_44/CARRYB[31][2] ,
         \mult_44/CARRYB[32][0] , \mult_44/CARRYB[32][1] ,
         \mult_44/CARRYB[32][2] , \mult_44/CARRYB[33][0] ,
         \mult_44/CARRYB[33][1] , \mult_44/CARRYB[33][2] ,
         \mult_44/CARRYB[34][0] , \mult_44/CARRYB[34][1] ,
         \mult_44/CARRYB[34][2] , \mult_44/CARRYB[35][0] ,
         \mult_44/CARRYB[35][1] , \mult_44/CARRYB[35][2] ,
         \mult_44/CARRYB[36][0] , \mult_44/CARRYB[36][1] ,
         \mult_44/CARRYB[36][2] , \mult_44/CARRYB[37][0] ,
         \mult_44/CARRYB[37][1] , \mult_44/CARRYB[37][2] ,
         \mult_44/CARRYB[38][0] , \mult_44/CARRYB[38][1] ,
         \mult_44/CARRYB[38][2] , \mult_44/CARRYB[39][0] ,
         \mult_44/CARRYB[39][1] , \mult_44/CARRYB[39][2] ,
         \mult_44/CARRYB[40][0] , \mult_44/CARRYB[40][1] ,
         \mult_44/CARRYB[40][2] , \mult_44/CARRYB[41][0] ,
         \mult_44/CARRYB[41][1] , \mult_44/CARRYB[41][2] ,
         \mult_44/CARRYB[42][0] , \mult_44/CARRYB[42][1] ,
         \mult_44/CARRYB[42][2] , \mult_44/CARRYB[43][0] ,
         \mult_44/CARRYB[43][1] , \mult_44/CARRYB[43][2] ,
         \mult_44/CARRYB[44][0] , \mult_44/CARRYB[44][1] ,
         \mult_44/CARRYB[44][2] , \mult_44/CARRYB[45][0] ,
         \mult_44/CARRYB[45][1] , \mult_44/CARRYB[45][2] ,
         \mult_44/CARRYB[46][0] , \mult_44/CARRYB[46][1] ,
         \mult_44/CARRYB[46][2] , \mult_44/CARRYB[47][0] ,
         \mult_44/CARRYB[47][1] , \mult_44/CARRYB[47][2] ,
         \mult_44/CARRYB[48][0] , \mult_44/CARRYB[48][1] ,
         \mult_44/CARRYB[48][2] , \mult_44/CARRYB[49][0] ,
         \mult_44/CARRYB[49][1] , \mult_44/CARRYB[49][2] ,
         \mult_44/CARRYB[50][0] , \mult_44/CARRYB[50][1] ,
         \mult_44/CARRYB[50][2] , \mult_44/CARRYB[51][0] ,
         \mult_44/CARRYB[51][1] , \mult_44/CARRYB[51][2] ,
         \mult_44/CARRYB[52][0] , \mult_44/CARRYB[52][1] ,
         \mult_44/CARRYB[52][2] , \mult_44/CARRYB[53][0] ,
         \mult_44/CARRYB[53][1] , \mult_44/CARRYB[53][2] ,
         \mult_44/CARRYB[54][0] , \mult_44/CARRYB[54][1] ,
         \mult_44/CARRYB[54][2] , \mult_44/CARRYB[55][0] ,
         \mult_44/CARRYB[55][1] , \mult_44/CARRYB[55][2] ,
         \mult_44/CARRYB[56][0] , \mult_44/CARRYB[56][1] ,
         \mult_44/CARRYB[56][2] , \mult_44/CARRYB[57][0] ,
         \mult_44/CARRYB[57][1] , \mult_44/CARRYB[57][2] ,
         \mult_44/CARRYB[58][0] , \mult_44/CARRYB[58][1] ,
         \mult_44/CARRYB[58][2] , \mult_44/CARRYB[59][0] ,
         \mult_44/CARRYB[59][1] , \mult_44/CARRYB[59][2] ,
         \mult_44/CARRYB[60][0] , \mult_44/CARRYB[60][1] ,
         \mult_44/CARRYB[60][2] , \mult_44/CARRYB[61][0] ,
         \mult_44/CARRYB[61][1] , \mult_44/CARRYB[62][0] , \mult_44/ab[0][1] ,
         \mult_44/ab[0][2] , \mult_44/ab[0][3] , \mult_44/ab[1][0] ,
         \mult_44/ab[1][1] , \mult_44/ab[1][2] , \mult_44/ab[1][3] ,
         \mult_44/ab[2][0] , \mult_44/ab[2][1] , \mult_44/ab[2][2] ,
         \mult_44/ab[2][3] , \mult_44/ab[3][0] , \mult_44/ab[3][1] ,
         \mult_44/ab[3][2] , \mult_44/ab[3][3] , \mult_44/ab[4][0] ,
         \mult_44/ab[4][1] , \mult_44/ab[4][2] , \mult_44/ab[4][3] ,
         \mult_44/ab[5][0] , \mult_44/ab[5][1] , \mult_44/ab[5][2] ,
         \mult_44/ab[5][3] , \mult_44/ab[6][0] , \mult_44/ab[6][1] ,
         \mult_44/ab[6][2] , \mult_44/ab[6][3] , \mult_44/ab[7][0] ,
         \mult_44/ab[7][1] , \mult_44/ab[7][2] , \mult_44/ab[7][3] ,
         \mult_44/ab[8][0] , \mult_44/ab[8][1] , \mult_44/ab[8][2] ,
         \mult_44/ab[8][3] , \mult_44/ab[9][0] , \mult_44/ab[9][1] ,
         \mult_44/ab[9][2] , \mult_44/ab[9][3] , \mult_44/ab[10][0] ,
         \mult_44/ab[10][1] , \mult_44/ab[10][2] , \mult_44/ab[10][3] ,
         \mult_44/ab[11][0] , \mult_44/ab[11][1] , \mult_44/ab[11][2] ,
         \mult_44/ab[11][3] , \mult_44/ab[12][0] , \mult_44/ab[12][1] ,
         \mult_44/ab[12][2] , \mult_44/ab[12][3] , \mult_44/ab[13][0] ,
         \mult_44/ab[13][1] , \mult_44/ab[13][2] , \mult_44/ab[13][3] ,
         \mult_44/ab[14][0] , \mult_44/ab[14][1] , \mult_44/ab[14][2] ,
         \mult_44/ab[14][3] , \mult_44/ab[15][0] , \mult_44/ab[15][1] ,
         \mult_44/ab[15][2] , \mult_44/ab[15][3] , \mult_44/ab[16][0] ,
         \mult_44/ab[16][1] , \mult_44/ab[16][2] , \mult_44/ab[16][3] ,
         \mult_44/ab[17][0] , \mult_44/ab[17][1] , \mult_44/ab[17][2] ,
         \mult_44/ab[17][3] , \mult_44/ab[18][0] , \mult_44/ab[18][1] ,
         \mult_44/ab[18][2] , \mult_44/ab[18][3] , \mult_44/ab[19][0] ,
         \mult_44/ab[19][1] , \mult_44/ab[19][2] , \mult_44/ab[19][3] ,
         \mult_44/ab[20][0] , \mult_44/ab[20][1] , \mult_44/ab[20][2] ,
         \mult_44/ab[20][3] , \mult_44/ab[21][0] , \mult_44/ab[21][1] ,
         \mult_44/ab[21][2] , \mult_44/ab[21][3] , \mult_44/ab[22][0] ,
         \mult_44/ab[22][1] , \mult_44/ab[22][2] , \mult_44/ab[22][3] ,
         \mult_44/ab[23][0] , \mult_44/ab[23][1] , \mult_44/ab[23][2] ,
         \mult_44/ab[23][3] , \mult_44/ab[24][0] , \mult_44/ab[24][1] ,
         \mult_44/ab[24][2] , \mult_44/ab[24][3] , \mult_44/ab[25][0] ,
         \mult_44/ab[25][1] , \mult_44/ab[25][2] , \mult_44/ab[25][3] ,
         \mult_44/ab[26][0] , \mult_44/ab[26][1] , \mult_44/ab[26][2] ,
         \mult_44/ab[26][3] , \mult_44/ab[27][0] , \mult_44/ab[27][1] ,
         \mult_44/ab[27][2] , \mult_44/ab[27][3] , \mult_44/ab[28][0] ,
         \mult_44/ab[28][1] , \mult_44/ab[28][2] , \mult_44/ab[28][3] ,
         \mult_44/ab[29][0] , \mult_44/ab[29][1] , \mult_44/ab[29][2] ,
         \mult_44/ab[29][3] , \mult_44/ab[30][0] , \mult_44/ab[30][1] ,
         \mult_44/ab[30][2] , \mult_44/ab[30][3] , \mult_44/ab[31][0] ,
         \mult_44/ab[31][1] , \mult_44/ab[31][2] , \mult_44/ab[31][3] ,
         \mult_44/ab[32][0] , \mult_44/ab[32][1] , \mult_44/ab[32][2] ,
         \mult_44/ab[32][3] , \mult_44/ab[33][0] , \mult_44/ab[33][1] ,
         \mult_44/ab[33][2] , \mult_44/ab[33][3] , \mult_44/ab[34][0] ,
         \mult_44/ab[34][1] , \mult_44/ab[34][2] , \mult_44/ab[34][3] ,
         \mult_44/ab[35][0] , \mult_44/ab[35][1] , \mult_44/ab[35][2] ,
         \mult_44/ab[35][3] , \mult_44/ab[36][0] , \mult_44/ab[36][1] ,
         \mult_44/ab[36][2] , \mult_44/ab[36][3] , \mult_44/ab[37][0] ,
         \mult_44/ab[37][1] , \mult_44/ab[37][2] , \mult_44/ab[37][3] ,
         \mult_44/ab[38][0] , \mult_44/ab[38][1] , \mult_44/ab[38][2] ,
         \mult_44/ab[38][3] , \mult_44/ab[39][0] , \mult_44/ab[39][1] ,
         \mult_44/ab[39][2] , \mult_44/ab[39][3] , \mult_44/ab[40][0] ,
         \mult_44/ab[40][1] , \mult_44/ab[40][2] , \mult_44/ab[40][3] ,
         \mult_44/ab[41][0] , \mult_44/ab[41][1] , \mult_44/ab[41][2] ,
         \mult_44/ab[41][3] , \mult_44/ab[42][0] , \mult_44/ab[42][1] ,
         \mult_44/ab[42][2] , \mult_44/ab[42][3] , \mult_44/ab[43][0] ,
         \mult_44/ab[43][1] , \mult_44/ab[43][2] , \mult_44/ab[43][3] ,
         \mult_44/ab[44][0] , \mult_44/ab[44][1] , \mult_44/ab[44][2] ,
         \mult_44/ab[44][3] , \mult_44/ab[45][0] , \mult_44/ab[45][1] ,
         \mult_44/ab[45][2] , \mult_44/ab[45][3] , \mult_44/ab[46][0] ,
         \mult_44/ab[46][1] , \mult_44/ab[46][2] , \mult_44/ab[46][3] ,
         \mult_44/ab[47][0] , \mult_44/ab[47][1] , \mult_44/ab[47][2] ,
         \mult_44/ab[47][3] , \mult_44/ab[48][0] , \mult_44/ab[48][1] ,
         \mult_44/ab[48][2] , \mult_44/ab[48][3] , \mult_44/ab[49][0] ,
         \mult_44/ab[49][1] , \mult_44/ab[49][2] , \mult_44/ab[49][3] ,
         \mult_44/ab[50][0] , \mult_44/ab[50][1] , \mult_44/ab[50][2] ,
         \mult_44/ab[50][3] , \mult_44/ab[51][0] , \mult_44/ab[51][1] ,
         \mult_44/ab[51][2] , \mult_44/ab[51][3] , \mult_44/ab[52][0] ,
         \mult_44/ab[52][1] , \mult_44/ab[52][2] , \mult_44/ab[52][3] ,
         \mult_44/ab[53][0] , \mult_44/ab[53][1] , \mult_44/ab[53][2] ,
         \mult_44/ab[53][3] , \mult_44/ab[54][0] , \mult_44/ab[54][1] ,
         \mult_44/ab[54][2] , \mult_44/ab[54][3] , \mult_44/ab[55][0] ,
         \mult_44/ab[55][1] , \mult_44/ab[55][2] , \mult_44/ab[55][3] ,
         \mult_44/ab[56][0] , \mult_44/ab[56][1] , \mult_44/ab[56][2] ,
         \mult_44/ab[56][3] , \mult_44/ab[57][0] , \mult_44/ab[57][1] ,
         \mult_44/ab[57][2] , \mult_44/ab[57][3] , \mult_44/ab[58][0] ,
         \mult_44/ab[58][1] , \mult_44/ab[58][2] , \mult_44/ab[58][3] ,
         \mult_44/ab[59][0] , \mult_44/ab[59][1] , \mult_44/ab[59][2] ,
         \mult_44/ab[59][3] , \mult_44/ab[60][0] , \mult_44/ab[60][1] ,
         \mult_44/ab[60][2] , \mult_44/ab[60][3] , \mult_44/ab[61][0] ,
         \mult_44/ab[61][1] , \mult_44/ab[61][2] , \mult_44/ab[62][0] ,
         \mult_44/ab[62][1] , \mult_44/ab[63][0] , n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305;
  wire   [63:4] swire;
  wire   [127:64] sreg;
  wire   [63:0] clocal;

  DFF \sreg_reg[64]  ( .D(swire[4]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[64]) );
  DFF \sreg_reg[65]  ( .D(swire[5]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[65]) );
  DFF \sreg_reg[66]  ( .D(swire[6]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[66]) );
  DFF \sreg_reg[67]  ( .D(swire[7]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[67]) );
  DFF \sreg_reg[68]  ( .D(swire[8]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[68]) );
  DFF \sreg_reg[69]  ( .D(swire[9]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[69]) );
  DFF \sreg_reg[70]  ( .D(swire[10]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[70]) );
  DFF \sreg_reg[71]  ( .D(swire[11]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[71]) );
  DFF \sreg_reg[72]  ( .D(swire[12]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[72]) );
  DFF \sreg_reg[73]  ( .D(swire[13]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[73]) );
  DFF \sreg_reg[74]  ( .D(swire[14]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[74]) );
  DFF \sreg_reg[75]  ( .D(swire[15]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[75]) );
  DFF \sreg_reg[76]  ( .D(swire[16]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[76]) );
  DFF \sreg_reg[77]  ( .D(swire[17]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[77]) );
  DFF \sreg_reg[78]  ( .D(swire[18]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[78]) );
  DFF \sreg_reg[79]  ( .D(swire[19]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[79]) );
  DFF \sreg_reg[80]  ( .D(swire[20]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[80]) );
  DFF \sreg_reg[81]  ( .D(swire[21]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[81]) );
  DFF \sreg_reg[82]  ( .D(swire[22]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[82]) );
  DFF \sreg_reg[83]  ( .D(swire[23]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[83]) );
  DFF \sreg_reg[84]  ( .D(swire[24]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[84]) );
  DFF \sreg_reg[85]  ( .D(swire[25]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[85]) );
  DFF \sreg_reg[86]  ( .D(swire[26]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[86]) );
  DFF \sreg_reg[87]  ( .D(swire[27]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[87]) );
  DFF \sreg_reg[88]  ( .D(swire[28]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[88]) );
  DFF \sreg_reg[89]  ( .D(swire[29]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[89]) );
  DFF \sreg_reg[90]  ( .D(swire[30]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[90]) );
  DFF \sreg_reg[91]  ( .D(swire[31]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[91]) );
  DFF \sreg_reg[92]  ( .D(swire[32]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[92]) );
  DFF \sreg_reg[93]  ( .D(swire[33]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[93]) );
  DFF \sreg_reg[94]  ( .D(swire[34]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[94]) );
  DFF \sreg_reg[95]  ( .D(swire[35]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[95]) );
  DFF \sreg_reg[96]  ( .D(swire[36]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[96]) );
  DFF \sreg_reg[97]  ( .D(swire[37]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[97]) );
  DFF \sreg_reg[98]  ( .D(swire[38]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[98]) );
  DFF \sreg_reg[99]  ( .D(swire[39]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[99]) );
  DFF \sreg_reg[100]  ( .D(swire[40]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[100]) );
  DFF \sreg_reg[101]  ( .D(swire[41]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[101]) );
  DFF \sreg_reg[102]  ( .D(swire[42]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[102]) );
  DFF \sreg_reg[103]  ( .D(swire[43]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[103]) );
  DFF \sreg_reg[104]  ( .D(swire[44]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[104]) );
  DFF \sreg_reg[105]  ( .D(swire[45]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[105]) );
  DFF \sreg_reg[106]  ( .D(swire[46]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[106]) );
  DFF \sreg_reg[107]  ( .D(swire[47]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[107]) );
  DFF \sreg_reg[108]  ( .D(swire[48]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[108]) );
  DFF \sreg_reg[109]  ( .D(swire[49]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[109]) );
  DFF \sreg_reg[110]  ( .D(swire[50]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[110]) );
  DFF \sreg_reg[111]  ( .D(swire[51]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[111]) );
  DFF \sreg_reg[112]  ( .D(swire[52]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[112]) );
  DFF \sreg_reg[113]  ( .D(swire[53]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[113]) );
  DFF \sreg_reg[114]  ( .D(swire[54]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[114]) );
  DFF \sreg_reg[115]  ( .D(swire[55]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[115]) );
  DFF \sreg_reg[116]  ( .D(swire[56]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[116]) );
  DFF \sreg_reg[117]  ( .D(swire[57]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[117]) );
  DFF \sreg_reg[118]  ( .D(swire[58]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[118]) );
  DFF \sreg_reg[119]  ( .D(swire[59]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[119]) );
  DFF \sreg_reg[120]  ( .D(swire[60]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[120]) );
  DFF \sreg_reg[121]  ( .D(swire[61]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[121]) );
  DFF \sreg_reg[122]  ( .D(swire[62]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[122]) );
  DFF \sreg_reg[123]  ( .D(swire[63]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[123]) );
  DFF \sreg_reg[63]  ( .D(c[63]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[59]) );
  DFF \sreg_reg[62]  ( .D(c[62]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[58]) );
  DFF \sreg_reg[61]  ( .D(c[61]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[57]) );
  DFF \sreg_reg[60]  ( .D(c[60]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[56]) );
  DFF \sreg_reg[59]  ( .D(c[59]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[55]) );
  DFF \sreg_reg[58]  ( .D(c[58]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[54]) );
  DFF \sreg_reg[57]  ( .D(c[57]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[53]) );
  DFF \sreg_reg[56]  ( .D(c[56]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[52]) );
  DFF \sreg_reg[55]  ( .D(c[55]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[51]) );
  DFF \sreg_reg[54]  ( .D(c[54]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[50]) );
  DFF \sreg_reg[53]  ( .D(c[53]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[49]) );
  DFF \sreg_reg[52]  ( .D(c[52]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[48]) );
  DFF \sreg_reg[51]  ( .D(c[51]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[47]) );
  DFF \sreg_reg[50]  ( .D(c[50]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[46]) );
  DFF \sreg_reg[49]  ( .D(c[49]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[45]) );
  DFF \sreg_reg[48]  ( .D(c[48]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[44]) );
  DFF \sreg_reg[47]  ( .D(c[47]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[43]) );
  DFF \sreg_reg[46]  ( .D(c[46]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[42]) );
  DFF \sreg_reg[45]  ( .D(c[45]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[41]) );
  DFF \sreg_reg[44]  ( .D(c[44]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[40]) );
  DFF \sreg_reg[43]  ( .D(c[43]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[39]) );
  DFF \sreg_reg[42]  ( .D(c[42]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[38]) );
  DFF \sreg_reg[41]  ( .D(c[41]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[37]) );
  DFF \sreg_reg[40]  ( .D(c[40]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[36]) );
  DFF \sreg_reg[39]  ( .D(c[39]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[35]) );
  DFF \sreg_reg[38]  ( .D(c[38]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[34]) );
  DFF \sreg_reg[37]  ( .D(c[37]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[33]) );
  DFF \sreg_reg[36]  ( .D(c[36]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[32]) );
  DFF \sreg_reg[35]  ( .D(c[35]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[31]) );
  DFF \sreg_reg[34]  ( .D(c[34]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[30]) );
  DFF \sreg_reg[33]  ( .D(c[33]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[29]) );
  DFF \sreg_reg[32]  ( .D(c[32]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[28]) );
  DFF \sreg_reg[31]  ( .D(c[31]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[27]) );
  DFF \sreg_reg[30]  ( .D(c[30]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[26]) );
  DFF \sreg_reg[29]  ( .D(c[29]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[25]) );
  DFF \sreg_reg[28]  ( .D(c[28]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[24]) );
  DFF \sreg_reg[27]  ( .D(c[27]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[23]) );
  DFF \sreg_reg[26]  ( .D(c[26]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[22]) );
  DFF \sreg_reg[25]  ( .D(c[25]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[21]) );
  DFF \sreg_reg[24]  ( .D(c[24]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[20]) );
  DFF \sreg_reg[23]  ( .D(c[23]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[19]) );
  DFF \sreg_reg[22]  ( .D(c[22]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[18]) );
  DFF \sreg_reg[21]  ( .D(c[21]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[17]) );
  DFF \sreg_reg[20]  ( .D(c[20]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[16]) );
  DFF \sreg_reg[19]  ( .D(c[19]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[15]) );
  DFF \sreg_reg[18]  ( .D(c[18]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[14]) );
  DFF \sreg_reg[17]  ( .D(c[17]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[13]) );
  DFF \sreg_reg[16]  ( .D(c[16]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[12]) );
  DFF \sreg_reg[15]  ( .D(c[15]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[11]) );
  DFF \sreg_reg[14]  ( .D(c[14]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[10]) );
  DFF \sreg_reg[13]  ( .D(c[13]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[9]) );
  DFF \sreg_reg[12]  ( .D(c[12]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[8]) );
  DFF \sreg_reg[11]  ( .D(c[11]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[7]) );
  DFF \sreg_reg[10]  ( .D(c[10]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[6]) );
  DFF \sreg_reg[9]  ( .D(c[9]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[5]) );
  DFF \sreg_reg[8]  ( .D(c[8]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[4]) );
  DFF \sreg_reg[7]  ( .D(c[7]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[3]) );
  DFF \sreg_reg[6]  ( .D(c[6]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[2]) );
  DFF \sreg_reg[5]  ( .D(c[5]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[1]) );
  DFF \sreg_reg[4]  ( .D(c[4]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[0]) );
  FADDER \mult_44/S3_2_2  ( .CIN(\mult_44/ab[2][2] ), .IN0(
        \mult_44/CARRYB[1][2] ), .IN1(\mult_44/ab[1][3] ), .COUT(
        \mult_44/CARRYB[2][2] ), .SUM(\mult_44/SUMB[2][2] ) );
  FADDER \mult_44/S2_2_1  ( .CIN(\mult_44/ab[2][1] ), .IN0(
        \mult_44/CARRYB[1][1] ), .IN1(\mult_44/SUMB[1][2] ), .COUT(
        \mult_44/CARRYB[2][1] ), .SUM(\mult_44/SUMB[2][1] ) );
  FADDER \mult_44/S1_2_0  ( .CIN(\mult_44/ab[2][0] ), .IN0(
        \mult_44/CARRYB[1][0] ), .IN1(\mult_44/SUMB[1][1] ), .COUT(
        \mult_44/CARRYB[2][0] ), .SUM(clocal[2]) );
  FADDER \mult_44/S3_3_2  ( .CIN(\mult_44/ab[3][2] ), .IN0(
        \mult_44/CARRYB[2][2] ), .IN1(\mult_44/ab[2][3] ), .COUT(
        \mult_44/CARRYB[3][2] ), .SUM(\mult_44/SUMB[3][2] ) );
  FADDER \mult_44/S2_3_1  ( .CIN(\mult_44/ab[3][1] ), .IN0(
        \mult_44/CARRYB[2][1] ), .IN1(\mult_44/SUMB[2][2] ), .COUT(
        \mult_44/CARRYB[3][1] ), .SUM(\mult_44/SUMB[3][1] ) );
  FADDER \mult_44/S1_3_0  ( .CIN(\mult_44/ab[3][0] ), .IN0(
        \mult_44/CARRYB[2][0] ), .IN1(\mult_44/SUMB[2][1] ), .COUT(
        \mult_44/CARRYB[3][0] ), .SUM(\mult_44/PROD1[3] ) );
  FADDER \mult_44/S3_4_2  ( .CIN(\mult_44/ab[4][2] ), .IN0(
        \mult_44/CARRYB[3][2] ), .IN1(\mult_44/ab[3][3] ), .COUT(
        \mult_44/CARRYB[4][2] ), .SUM(\mult_44/SUMB[4][2] ) );
  FADDER \mult_44/S2_4_1  ( .CIN(\mult_44/ab[4][1] ), .IN0(
        \mult_44/CARRYB[3][1] ), .IN1(\mult_44/SUMB[3][2] ), .COUT(
        \mult_44/CARRYB[4][1] ), .SUM(\mult_44/SUMB[4][1] ) );
  FADDER \mult_44/S1_4_0  ( .CIN(\mult_44/ab[4][0] ), .IN0(
        \mult_44/CARRYB[3][0] ), .IN1(\mult_44/SUMB[3][1] ), .COUT(
        \mult_44/CARRYB[4][0] ), .SUM(clocal[4]) );
  FADDER \mult_44/S3_5_2  ( .CIN(\mult_44/ab[5][2] ), .IN0(
        \mult_44/CARRYB[4][2] ), .IN1(\mult_44/ab[4][3] ), .COUT(
        \mult_44/CARRYB[5][2] ), .SUM(\mult_44/SUMB[5][2] ) );
  FADDER \mult_44/S2_5_1  ( .CIN(\mult_44/ab[5][1] ), .IN0(
        \mult_44/CARRYB[4][1] ), .IN1(\mult_44/SUMB[4][2] ), .COUT(
        \mult_44/CARRYB[5][1] ), .SUM(\mult_44/SUMB[5][1] ) );
  FADDER \mult_44/S1_5_0  ( .CIN(\mult_44/ab[5][0] ), .IN0(
        \mult_44/CARRYB[4][0] ), .IN1(\mult_44/SUMB[4][1] ), .COUT(
        \mult_44/CARRYB[5][0] ), .SUM(clocal[5]) );
  FADDER \mult_44/S3_6_2  ( .CIN(\mult_44/ab[6][2] ), .IN0(
        \mult_44/CARRYB[5][2] ), .IN1(\mult_44/ab[5][3] ), .COUT(
        \mult_44/CARRYB[6][2] ), .SUM(\mult_44/SUMB[6][2] ) );
  FADDER \mult_44/S2_6_1  ( .CIN(\mult_44/ab[6][1] ), .IN0(
        \mult_44/CARRYB[5][1] ), .IN1(\mult_44/SUMB[5][2] ), .COUT(
        \mult_44/CARRYB[6][1] ), .SUM(\mult_44/SUMB[6][1] ) );
  FADDER \mult_44/S1_6_0  ( .CIN(\mult_44/ab[6][0] ), .IN0(
        \mult_44/CARRYB[5][0] ), .IN1(\mult_44/SUMB[5][1] ), .COUT(
        \mult_44/CARRYB[6][0] ), .SUM(clocal[6]) );
  FADDER \mult_44/S3_7_2  ( .CIN(\mult_44/ab[7][2] ), .IN0(
        \mult_44/CARRYB[6][2] ), .IN1(\mult_44/ab[6][3] ), .COUT(
        \mult_44/CARRYB[7][2] ), .SUM(\mult_44/SUMB[7][2] ) );
  FADDER \mult_44/S2_7_1  ( .CIN(\mult_44/ab[7][1] ), .IN0(
        \mult_44/CARRYB[6][1] ), .IN1(\mult_44/SUMB[6][2] ), .COUT(
        \mult_44/CARRYB[7][1] ), .SUM(\mult_44/SUMB[7][1] ) );
  FADDER \mult_44/S1_7_0  ( .CIN(\mult_44/ab[7][0] ), .IN0(
        \mult_44/CARRYB[6][0] ), .IN1(\mult_44/SUMB[6][1] ), .COUT(
        \mult_44/CARRYB[7][0] ), .SUM(clocal[7]) );
  FADDER \mult_44/S3_8_2  ( .CIN(\mult_44/ab[8][2] ), .IN0(
        \mult_44/CARRYB[7][2] ), .IN1(\mult_44/ab[7][3] ), .COUT(
        \mult_44/CARRYB[8][2] ), .SUM(\mult_44/SUMB[8][2] ) );
  FADDER \mult_44/S2_8_1  ( .CIN(\mult_44/ab[8][1] ), .IN0(
        \mult_44/CARRYB[7][1] ), .IN1(\mult_44/SUMB[7][2] ), .COUT(
        \mult_44/CARRYB[8][1] ), .SUM(\mult_44/SUMB[8][1] ) );
  FADDER \mult_44/S1_8_0  ( .CIN(\mult_44/ab[8][0] ), .IN0(
        \mult_44/CARRYB[7][0] ), .IN1(\mult_44/SUMB[7][1] ), .COUT(
        \mult_44/CARRYB[8][0] ), .SUM(clocal[8]) );
  FADDER \mult_44/S3_9_2  ( .CIN(\mult_44/ab[9][2] ), .IN0(
        \mult_44/CARRYB[8][2] ), .IN1(\mult_44/ab[8][3] ), .COUT(
        \mult_44/CARRYB[9][2] ), .SUM(\mult_44/SUMB[9][2] ) );
  FADDER \mult_44/S2_9_1  ( .CIN(\mult_44/ab[9][1] ), .IN0(
        \mult_44/CARRYB[8][1] ), .IN1(\mult_44/SUMB[8][2] ), .COUT(
        \mult_44/CARRYB[9][1] ), .SUM(\mult_44/SUMB[9][1] ) );
  FADDER \mult_44/S1_9_0  ( .CIN(\mult_44/ab[9][0] ), .IN0(
        \mult_44/CARRYB[8][0] ), .IN1(\mult_44/SUMB[8][1] ), .COUT(
        \mult_44/CARRYB[9][0] ), .SUM(clocal[9]) );
  FADDER \mult_44/S3_10_2  ( .CIN(\mult_44/ab[10][2] ), .IN0(
        \mult_44/CARRYB[9][2] ), .IN1(\mult_44/ab[9][3] ), .COUT(
        \mult_44/CARRYB[10][2] ), .SUM(\mult_44/SUMB[10][2] ) );
  FADDER \mult_44/S2_10_1  ( .CIN(\mult_44/ab[10][1] ), .IN0(
        \mult_44/CARRYB[9][1] ), .IN1(\mult_44/SUMB[9][2] ), .COUT(
        \mult_44/CARRYB[10][1] ), .SUM(\mult_44/SUMB[10][1] ) );
  FADDER \mult_44/S1_10_0  ( .CIN(\mult_44/ab[10][0] ), .IN0(
        \mult_44/CARRYB[9][0] ), .IN1(\mult_44/SUMB[9][1] ), .COUT(
        \mult_44/CARRYB[10][0] ), .SUM(clocal[10]) );
  FADDER \mult_44/S3_11_2  ( .CIN(\mult_44/ab[11][2] ), .IN0(
        \mult_44/CARRYB[10][2] ), .IN1(\mult_44/ab[10][3] ), .COUT(
        \mult_44/CARRYB[11][2] ), .SUM(\mult_44/SUMB[11][2] ) );
  FADDER \mult_44/S2_11_1  ( .CIN(\mult_44/ab[11][1] ), .IN0(
        \mult_44/CARRYB[10][1] ), .IN1(\mult_44/SUMB[10][2] ), .COUT(
        \mult_44/CARRYB[11][1] ), .SUM(\mult_44/SUMB[11][1] ) );
  FADDER \mult_44/S1_11_0  ( .CIN(\mult_44/ab[11][0] ), .IN0(
        \mult_44/CARRYB[10][0] ), .IN1(\mult_44/SUMB[10][1] ), .COUT(
        \mult_44/CARRYB[11][0] ), .SUM(clocal[11]) );
  FADDER \mult_44/S3_12_2  ( .CIN(\mult_44/ab[12][2] ), .IN0(
        \mult_44/CARRYB[11][2] ), .IN1(\mult_44/ab[11][3] ), .COUT(
        \mult_44/CARRYB[12][2] ), .SUM(\mult_44/SUMB[12][2] ) );
  FADDER \mult_44/S2_12_1  ( .CIN(\mult_44/ab[12][1] ), .IN0(
        \mult_44/CARRYB[11][1] ), .IN1(\mult_44/SUMB[11][2] ), .COUT(
        \mult_44/CARRYB[12][1] ), .SUM(\mult_44/SUMB[12][1] ) );
  FADDER \mult_44/S1_12_0  ( .CIN(\mult_44/ab[12][0] ), .IN0(
        \mult_44/CARRYB[11][0] ), .IN1(\mult_44/SUMB[11][1] ), .COUT(
        \mult_44/CARRYB[12][0] ), .SUM(clocal[12]) );
  FADDER \mult_44/S3_13_2  ( .CIN(\mult_44/ab[13][2] ), .IN0(
        \mult_44/CARRYB[12][2] ), .IN1(\mult_44/ab[12][3] ), .COUT(
        \mult_44/CARRYB[13][2] ), .SUM(\mult_44/SUMB[13][2] ) );
  FADDER \mult_44/S2_13_1  ( .CIN(\mult_44/ab[13][1] ), .IN0(
        \mult_44/CARRYB[12][1] ), .IN1(\mult_44/SUMB[12][2] ), .COUT(
        \mult_44/CARRYB[13][1] ), .SUM(\mult_44/SUMB[13][1] ) );
  FADDER \mult_44/S1_13_0  ( .CIN(\mult_44/ab[13][0] ), .IN0(
        \mult_44/CARRYB[12][0] ), .IN1(\mult_44/SUMB[12][1] ), .COUT(
        \mult_44/CARRYB[13][0] ), .SUM(clocal[13]) );
  FADDER \mult_44/S3_14_2  ( .CIN(\mult_44/ab[14][2] ), .IN0(
        \mult_44/CARRYB[13][2] ), .IN1(\mult_44/ab[13][3] ), .COUT(
        \mult_44/CARRYB[14][2] ), .SUM(\mult_44/SUMB[14][2] ) );
  FADDER \mult_44/S2_14_1  ( .CIN(\mult_44/ab[14][1] ), .IN0(
        \mult_44/CARRYB[13][1] ), .IN1(\mult_44/SUMB[13][2] ), .COUT(
        \mult_44/CARRYB[14][1] ), .SUM(\mult_44/SUMB[14][1] ) );
  FADDER \mult_44/S1_14_0  ( .CIN(\mult_44/ab[14][0] ), .IN0(
        \mult_44/CARRYB[13][0] ), .IN1(\mult_44/SUMB[13][1] ), .COUT(
        \mult_44/CARRYB[14][0] ), .SUM(clocal[14]) );
  FADDER \mult_44/S3_15_2  ( .CIN(\mult_44/ab[15][2] ), .IN0(
        \mult_44/CARRYB[14][2] ), .IN1(\mult_44/ab[14][3] ), .COUT(
        \mult_44/CARRYB[15][2] ), .SUM(\mult_44/SUMB[15][2] ) );
  FADDER \mult_44/S2_15_1  ( .CIN(\mult_44/ab[15][1] ), .IN0(
        \mult_44/CARRYB[14][1] ), .IN1(\mult_44/SUMB[14][2] ), .COUT(
        \mult_44/CARRYB[15][1] ), .SUM(\mult_44/SUMB[15][1] ) );
  FADDER \mult_44/S1_15_0  ( .CIN(\mult_44/ab[15][0] ), .IN0(
        \mult_44/CARRYB[14][0] ), .IN1(\mult_44/SUMB[14][1] ), .COUT(
        \mult_44/CARRYB[15][0] ), .SUM(clocal[15]) );
  FADDER \mult_44/S3_16_2  ( .CIN(\mult_44/ab[16][2] ), .IN0(
        \mult_44/CARRYB[15][2] ), .IN1(\mult_44/ab[15][3] ), .COUT(
        \mult_44/CARRYB[16][2] ), .SUM(\mult_44/SUMB[16][2] ) );
  FADDER \mult_44/S2_16_1  ( .CIN(\mult_44/ab[16][1] ), .IN0(
        \mult_44/CARRYB[15][1] ), .IN1(\mult_44/SUMB[15][2] ), .COUT(
        \mult_44/CARRYB[16][1] ), .SUM(\mult_44/SUMB[16][1] ) );
  FADDER \mult_44/S1_16_0  ( .CIN(\mult_44/ab[16][0] ), .IN0(
        \mult_44/CARRYB[15][0] ), .IN1(\mult_44/SUMB[15][1] ), .COUT(
        \mult_44/CARRYB[16][0] ), .SUM(clocal[16]) );
  FADDER \mult_44/S3_17_2  ( .CIN(\mult_44/ab[17][2] ), .IN0(
        \mult_44/CARRYB[16][2] ), .IN1(\mult_44/ab[16][3] ), .COUT(
        \mult_44/CARRYB[17][2] ), .SUM(\mult_44/SUMB[17][2] ) );
  FADDER \mult_44/S2_17_1  ( .CIN(\mult_44/ab[17][1] ), .IN0(
        \mult_44/CARRYB[16][1] ), .IN1(\mult_44/SUMB[16][2] ), .COUT(
        \mult_44/CARRYB[17][1] ), .SUM(\mult_44/SUMB[17][1] ) );
  FADDER \mult_44/S1_17_0  ( .CIN(\mult_44/ab[17][0] ), .IN0(
        \mult_44/CARRYB[16][0] ), .IN1(\mult_44/SUMB[16][1] ), .COUT(
        \mult_44/CARRYB[17][0] ), .SUM(clocal[17]) );
  FADDER \mult_44/S3_18_2  ( .CIN(\mult_44/ab[18][2] ), .IN0(
        \mult_44/CARRYB[17][2] ), .IN1(\mult_44/ab[17][3] ), .COUT(
        \mult_44/CARRYB[18][2] ), .SUM(\mult_44/SUMB[18][2] ) );
  FADDER \mult_44/S2_18_1  ( .CIN(\mult_44/ab[18][1] ), .IN0(
        \mult_44/CARRYB[17][1] ), .IN1(\mult_44/SUMB[17][2] ), .COUT(
        \mult_44/CARRYB[18][1] ), .SUM(\mult_44/SUMB[18][1] ) );
  FADDER \mult_44/S1_18_0  ( .CIN(\mult_44/ab[18][0] ), .IN0(
        \mult_44/CARRYB[17][0] ), .IN1(\mult_44/SUMB[17][1] ), .COUT(
        \mult_44/CARRYB[18][0] ), .SUM(clocal[18]) );
  FADDER \mult_44/S3_19_2  ( .CIN(\mult_44/ab[19][2] ), .IN0(
        \mult_44/CARRYB[18][2] ), .IN1(\mult_44/ab[18][3] ), .COUT(
        \mult_44/CARRYB[19][2] ), .SUM(\mult_44/SUMB[19][2] ) );
  FADDER \mult_44/S2_19_1  ( .CIN(\mult_44/ab[19][1] ), .IN0(
        \mult_44/CARRYB[18][1] ), .IN1(\mult_44/SUMB[18][2] ), .COUT(
        \mult_44/CARRYB[19][1] ), .SUM(\mult_44/SUMB[19][1] ) );
  FADDER \mult_44/S1_19_0  ( .CIN(\mult_44/ab[19][0] ), .IN0(
        \mult_44/CARRYB[18][0] ), .IN1(\mult_44/SUMB[18][1] ), .COUT(
        \mult_44/CARRYB[19][0] ), .SUM(clocal[19]) );
  FADDER \mult_44/S3_20_2  ( .CIN(\mult_44/ab[20][2] ), .IN0(
        \mult_44/CARRYB[19][2] ), .IN1(\mult_44/ab[19][3] ), .COUT(
        \mult_44/CARRYB[20][2] ), .SUM(\mult_44/SUMB[20][2] ) );
  FADDER \mult_44/S2_20_1  ( .CIN(\mult_44/ab[20][1] ), .IN0(
        \mult_44/CARRYB[19][1] ), .IN1(\mult_44/SUMB[19][2] ), .COUT(
        \mult_44/CARRYB[20][1] ), .SUM(\mult_44/SUMB[20][1] ) );
  FADDER \mult_44/S1_20_0  ( .CIN(\mult_44/ab[20][0] ), .IN0(
        \mult_44/CARRYB[19][0] ), .IN1(\mult_44/SUMB[19][1] ), .COUT(
        \mult_44/CARRYB[20][0] ), .SUM(clocal[20]) );
  FADDER \mult_44/S3_21_2  ( .CIN(\mult_44/ab[21][2] ), .IN0(
        \mult_44/CARRYB[20][2] ), .IN1(\mult_44/ab[20][3] ), .COUT(
        \mult_44/CARRYB[21][2] ), .SUM(\mult_44/SUMB[21][2] ) );
  FADDER \mult_44/S2_21_1  ( .CIN(\mult_44/ab[21][1] ), .IN0(
        \mult_44/CARRYB[20][1] ), .IN1(\mult_44/SUMB[20][2] ), .COUT(
        \mult_44/CARRYB[21][1] ), .SUM(\mult_44/SUMB[21][1] ) );
  FADDER \mult_44/S1_21_0  ( .CIN(\mult_44/ab[21][0] ), .IN0(
        \mult_44/CARRYB[20][0] ), .IN1(\mult_44/SUMB[20][1] ), .COUT(
        \mult_44/CARRYB[21][0] ), .SUM(clocal[21]) );
  FADDER \mult_44/S3_22_2  ( .CIN(\mult_44/ab[22][2] ), .IN0(
        \mult_44/CARRYB[21][2] ), .IN1(\mult_44/ab[21][3] ), .COUT(
        \mult_44/CARRYB[22][2] ), .SUM(\mult_44/SUMB[22][2] ) );
  FADDER \mult_44/S2_22_1  ( .CIN(\mult_44/ab[22][1] ), .IN0(
        \mult_44/CARRYB[21][1] ), .IN1(\mult_44/SUMB[21][2] ), .COUT(
        \mult_44/CARRYB[22][1] ), .SUM(\mult_44/SUMB[22][1] ) );
  FADDER \mult_44/S1_22_0  ( .CIN(\mult_44/ab[22][0] ), .IN0(
        \mult_44/CARRYB[21][0] ), .IN1(\mult_44/SUMB[21][1] ), .COUT(
        \mult_44/CARRYB[22][0] ), .SUM(clocal[22]) );
  FADDER \mult_44/S3_23_2  ( .CIN(\mult_44/ab[23][2] ), .IN0(
        \mult_44/CARRYB[22][2] ), .IN1(\mult_44/ab[22][3] ), .COUT(
        \mult_44/CARRYB[23][2] ), .SUM(\mult_44/SUMB[23][2] ) );
  FADDER \mult_44/S2_23_1  ( .CIN(\mult_44/ab[23][1] ), .IN0(
        \mult_44/CARRYB[22][1] ), .IN1(\mult_44/SUMB[22][2] ), .COUT(
        \mult_44/CARRYB[23][1] ), .SUM(\mult_44/SUMB[23][1] ) );
  FADDER \mult_44/S1_23_0  ( .CIN(\mult_44/ab[23][0] ), .IN0(
        \mult_44/CARRYB[22][0] ), .IN1(\mult_44/SUMB[22][1] ), .COUT(
        \mult_44/CARRYB[23][0] ), .SUM(clocal[23]) );
  FADDER \mult_44/S3_24_2  ( .CIN(\mult_44/ab[24][2] ), .IN0(
        \mult_44/CARRYB[23][2] ), .IN1(\mult_44/ab[23][3] ), .COUT(
        \mult_44/CARRYB[24][2] ), .SUM(\mult_44/SUMB[24][2] ) );
  FADDER \mult_44/S2_24_1  ( .CIN(\mult_44/ab[24][1] ), .IN0(
        \mult_44/CARRYB[23][1] ), .IN1(\mult_44/SUMB[23][2] ), .COUT(
        \mult_44/CARRYB[24][1] ), .SUM(\mult_44/SUMB[24][1] ) );
  FADDER \mult_44/S1_24_0  ( .CIN(\mult_44/ab[24][0] ), .IN0(
        \mult_44/CARRYB[23][0] ), .IN1(\mult_44/SUMB[23][1] ), .COUT(
        \mult_44/CARRYB[24][0] ), .SUM(clocal[24]) );
  FADDER \mult_44/S3_25_2  ( .CIN(\mult_44/ab[25][2] ), .IN0(
        \mult_44/CARRYB[24][2] ), .IN1(\mult_44/ab[24][3] ), .COUT(
        \mult_44/CARRYB[25][2] ), .SUM(\mult_44/SUMB[25][2] ) );
  FADDER \mult_44/S2_25_1  ( .CIN(\mult_44/ab[25][1] ), .IN0(
        \mult_44/CARRYB[24][1] ), .IN1(\mult_44/SUMB[24][2] ), .COUT(
        \mult_44/CARRYB[25][1] ), .SUM(\mult_44/SUMB[25][1] ) );
  FADDER \mult_44/S1_25_0  ( .CIN(\mult_44/ab[25][0] ), .IN0(
        \mult_44/CARRYB[24][0] ), .IN1(\mult_44/SUMB[24][1] ), .COUT(
        \mult_44/CARRYB[25][0] ), .SUM(clocal[25]) );
  FADDER \mult_44/S3_26_2  ( .CIN(\mult_44/ab[26][2] ), .IN0(
        \mult_44/CARRYB[25][2] ), .IN1(\mult_44/ab[25][3] ), .COUT(
        \mult_44/CARRYB[26][2] ), .SUM(\mult_44/SUMB[26][2] ) );
  FADDER \mult_44/S2_26_1  ( .CIN(\mult_44/ab[26][1] ), .IN0(
        \mult_44/CARRYB[25][1] ), .IN1(\mult_44/SUMB[25][2] ), .COUT(
        \mult_44/CARRYB[26][1] ), .SUM(\mult_44/SUMB[26][1] ) );
  FADDER \mult_44/S1_26_0  ( .CIN(\mult_44/ab[26][0] ), .IN0(
        \mult_44/CARRYB[25][0] ), .IN1(\mult_44/SUMB[25][1] ), .COUT(
        \mult_44/CARRYB[26][0] ), .SUM(clocal[26]) );
  FADDER \mult_44/S3_27_2  ( .CIN(\mult_44/ab[27][2] ), .IN0(
        \mult_44/CARRYB[26][2] ), .IN1(\mult_44/ab[26][3] ), .COUT(
        \mult_44/CARRYB[27][2] ), .SUM(\mult_44/SUMB[27][2] ) );
  FADDER \mult_44/S2_27_1  ( .CIN(\mult_44/ab[27][1] ), .IN0(
        \mult_44/CARRYB[26][1] ), .IN1(\mult_44/SUMB[26][2] ), .COUT(
        \mult_44/CARRYB[27][1] ), .SUM(\mult_44/SUMB[27][1] ) );
  FADDER \mult_44/S1_27_0  ( .CIN(\mult_44/ab[27][0] ), .IN0(
        \mult_44/CARRYB[26][0] ), .IN1(\mult_44/SUMB[26][1] ), .COUT(
        \mult_44/CARRYB[27][0] ), .SUM(clocal[27]) );
  FADDER \mult_44/S3_28_2  ( .CIN(\mult_44/ab[28][2] ), .IN0(
        \mult_44/CARRYB[27][2] ), .IN1(\mult_44/ab[27][3] ), .COUT(
        \mult_44/CARRYB[28][2] ), .SUM(\mult_44/SUMB[28][2] ) );
  FADDER \mult_44/S2_28_1  ( .CIN(\mult_44/ab[28][1] ), .IN0(
        \mult_44/CARRYB[27][1] ), .IN1(\mult_44/SUMB[27][2] ), .COUT(
        \mult_44/CARRYB[28][1] ), .SUM(\mult_44/SUMB[28][1] ) );
  FADDER \mult_44/S1_28_0  ( .CIN(\mult_44/ab[28][0] ), .IN0(
        \mult_44/CARRYB[27][0] ), .IN1(\mult_44/SUMB[27][1] ), .COUT(
        \mult_44/CARRYB[28][0] ), .SUM(clocal[28]) );
  FADDER \mult_44/S3_29_2  ( .CIN(\mult_44/ab[29][2] ), .IN0(
        \mult_44/CARRYB[28][2] ), .IN1(\mult_44/ab[28][3] ), .COUT(
        \mult_44/CARRYB[29][2] ), .SUM(\mult_44/SUMB[29][2] ) );
  FADDER \mult_44/S2_29_1  ( .CIN(\mult_44/ab[29][1] ), .IN0(
        \mult_44/CARRYB[28][1] ), .IN1(\mult_44/SUMB[28][2] ), .COUT(
        \mult_44/CARRYB[29][1] ), .SUM(\mult_44/SUMB[29][1] ) );
  FADDER \mult_44/S1_29_0  ( .CIN(\mult_44/ab[29][0] ), .IN0(
        \mult_44/CARRYB[28][0] ), .IN1(\mult_44/SUMB[28][1] ), .COUT(
        \mult_44/CARRYB[29][0] ), .SUM(clocal[29]) );
  FADDER \mult_44/S3_30_2  ( .CIN(\mult_44/ab[30][2] ), .IN0(
        \mult_44/CARRYB[29][2] ), .IN1(\mult_44/ab[29][3] ), .COUT(
        \mult_44/CARRYB[30][2] ), .SUM(\mult_44/SUMB[30][2] ) );
  FADDER \mult_44/S2_30_1  ( .CIN(\mult_44/ab[30][1] ), .IN0(
        \mult_44/CARRYB[29][1] ), .IN1(\mult_44/SUMB[29][2] ), .COUT(
        \mult_44/CARRYB[30][1] ), .SUM(\mult_44/SUMB[30][1] ) );
  FADDER \mult_44/S1_30_0  ( .CIN(\mult_44/ab[30][0] ), .IN0(
        \mult_44/CARRYB[29][0] ), .IN1(\mult_44/SUMB[29][1] ), .COUT(
        \mult_44/CARRYB[30][0] ), .SUM(clocal[30]) );
  FADDER \mult_44/S3_31_2  ( .CIN(\mult_44/ab[31][2] ), .IN0(
        \mult_44/CARRYB[30][2] ), .IN1(\mult_44/ab[30][3] ), .COUT(
        \mult_44/CARRYB[31][2] ), .SUM(\mult_44/SUMB[31][2] ) );
  FADDER \mult_44/S2_31_1  ( .CIN(\mult_44/ab[31][1] ), .IN0(
        \mult_44/CARRYB[30][1] ), .IN1(\mult_44/SUMB[30][2] ), .COUT(
        \mult_44/CARRYB[31][1] ), .SUM(\mult_44/SUMB[31][1] ) );
  FADDER \mult_44/S1_31_0  ( .CIN(\mult_44/ab[31][0] ), .IN0(
        \mult_44/CARRYB[30][0] ), .IN1(\mult_44/SUMB[30][1] ), .COUT(
        \mult_44/CARRYB[31][0] ), .SUM(clocal[31]) );
  FADDER \mult_44/S3_32_2  ( .CIN(\mult_44/ab[32][2] ), .IN0(
        \mult_44/CARRYB[31][2] ), .IN1(\mult_44/ab[31][3] ), .COUT(
        \mult_44/CARRYB[32][2] ), .SUM(\mult_44/SUMB[32][2] ) );
  FADDER \mult_44/S2_32_1  ( .CIN(\mult_44/ab[32][1] ), .IN0(
        \mult_44/CARRYB[31][1] ), .IN1(\mult_44/SUMB[31][2] ), .COUT(
        \mult_44/CARRYB[32][1] ), .SUM(\mult_44/SUMB[32][1] ) );
  FADDER \mult_44/S1_32_0  ( .CIN(\mult_44/ab[32][0] ), .IN0(
        \mult_44/CARRYB[31][0] ), .IN1(\mult_44/SUMB[31][1] ), .COUT(
        \mult_44/CARRYB[32][0] ), .SUM(clocal[32]) );
  FADDER \mult_44/S3_33_2  ( .CIN(\mult_44/ab[33][2] ), .IN0(
        \mult_44/CARRYB[32][2] ), .IN1(\mult_44/ab[32][3] ), .COUT(
        \mult_44/CARRYB[33][2] ), .SUM(\mult_44/SUMB[33][2] ) );
  FADDER \mult_44/S2_33_1  ( .CIN(\mult_44/ab[33][1] ), .IN0(
        \mult_44/CARRYB[32][1] ), .IN1(\mult_44/SUMB[32][2] ), .COUT(
        \mult_44/CARRYB[33][1] ), .SUM(\mult_44/SUMB[33][1] ) );
  FADDER \mult_44/S1_33_0  ( .CIN(\mult_44/ab[33][0] ), .IN0(
        \mult_44/CARRYB[32][0] ), .IN1(\mult_44/SUMB[32][1] ), .COUT(
        \mult_44/CARRYB[33][0] ), .SUM(clocal[33]) );
  FADDER \mult_44/S3_34_2  ( .CIN(\mult_44/ab[34][2] ), .IN0(
        \mult_44/CARRYB[33][2] ), .IN1(\mult_44/ab[33][3] ), .COUT(
        \mult_44/CARRYB[34][2] ), .SUM(\mult_44/SUMB[34][2] ) );
  FADDER \mult_44/S2_34_1  ( .CIN(\mult_44/ab[34][1] ), .IN0(
        \mult_44/CARRYB[33][1] ), .IN1(\mult_44/SUMB[33][2] ), .COUT(
        \mult_44/CARRYB[34][1] ), .SUM(\mult_44/SUMB[34][1] ) );
  FADDER \mult_44/S1_34_0  ( .CIN(\mult_44/ab[34][0] ), .IN0(
        \mult_44/CARRYB[33][0] ), .IN1(\mult_44/SUMB[33][1] ), .COUT(
        \mult_44/CARRYB[34][0] ), .SUM(clocal[34]) );
  FADDER \mult_44/S3_35_2  ( .CIN(\mult_44/ab[35][2] ), .IN0(
        \mult_44/CARRYB[34][2] ), .IN1(\mult_44/ab[34][3] ), .COUT(
        \mult_44/CARRYB[35][2] ), .SUM(\mult_44/SUMB[35][2] ) );
  FADDER \mult_44/S2_35_1  ( .CIN(\mult_44/ab[35][1] ), .IN0(
        \mult_44/CARRYB[34][1] ), .IN1(\mult_44/SUMB[34][2] ), .COUT(
        \mult_44/CARRYB[35][1] ), .SUM(\mult_44/SUMB[35][1] ) );
  FADDER \mult_44/S1_35_0  ( .CIN(\mult_44/ab[35][0] ), .IN0(
        \mult_44/CARRYB[34][0] ), .IN1(\mult_44/SUMB[34][1] ), .COUT(
        \mult_44/CARRYB[35][0] ), .SUM(clocal[35]) );
  FADDER \mult_44/S3_36_2  ( .CIN(\mult_44/ab[36][2] ), .IN0(
        \mult_44/CARRYB[35][2] ), .IN1(\mult_44/ab[35][3] ), .COUT(
        \mult_44/CARRYB[36][2] ), .SUM(\mult_44/SUMB[36][2] ) );
  FADDER \mult_44/S2_36_1  ( .CIN(\mult_44/ab[36][1] ), .IN0(
        \mult_44/CARRYB[35][1] ), .IN1(\mult_44/SUMB[35][2] ), .COUT(
        \mult_44/CARRYB[36][1] ), .SUM(\mult_44/SUMB[36][1] ) );
  FADDER \mult_44/S1_36_0  ( .CIN(\mult_44/ab[36][0] ), .IN0(
        \mult_44/CARRYB[35][0] ), .IN1(\mult_44/SUMB[35][1] ), .COUT(
        \mult_44/CARRYB[36][0] ), .SUM(clocal[36]) );
  FADDER \mult_44/S3_37_2  ( .CIN(\mult_44/ab[37][2] ), .IN0(
        \mult_44/CARRYB[36][2] ), .IN1(\mult_44/ab[36][3] ), .COUT(
        \mult_44/CARRYB[37][2] ), .SUM(\mult_44/SUMB[37][2] ) );
  FADDER \mult_44/S2_37_1  ( .CIN(\mult_44/ab[37][1] ), .IN0(
        \mult_44/CARRYB[36][1] ), .IN1(\mult_44/SUMB[36][2] ), .COUT(
        \mult_44/CARRYB[37][1] ), .SUM(\mult_44/SUMB[37][1] ) );
  FADDER \mult_44/S1_37_0  ( .CIN(\mult_44/ab[37][0] ), .IN0(
        \mult_44/CARRYB[36][0] ), .IN1(\mult_44/SUMB[36][1] ), .COUT(
        \mult_44/CARRYB[37][0] ), .SUM(clocal[37]) );
  FADDER \mult_44/S3_38_2  ( .CIN(\mult_44/ab[38][2] ), .IN0(
        \mult_44/CARRYB[37][2] ), .IN1(\mult_44/ab[37][3] ), .COUT(
        \mult_44/CARRYB[38][2] ), .SUM(\mult_44/SUMB[38][2] ) );
  FADDER \mult_44/S2_38_1  ( .CIN(\mult_44/ab[38][1] ), .IN0(
        \mult_44/CARRYB[37][1] ), .IN1(\mult_44/SUMB[37][2] ), .COUT(
        \mult_44/CARRYB[38][1] ), .SUM(\mult_44/SUMB[38][1] ) );
  FADDER \mult_44/S1_38_0  ( .CIN(\mult_44/ab[38][0] ), .IN0(
        \mult_44/CARRYB[37][0] ), .IN1(\mult_44/SUMB[37][1] ), .COUT(
        \mult_44/CARRYB[38][0] ), .SUM(clocal[38]) );
  FADDER \mult_44/S3_39_2  ( .CIN(\mult_44/ab[39][2] ), .IN0(
        \mult_44/CARRYB[38][2] ), .IN1(\mult_44/ab[38][3] ), .COUT(
        \mult_44/CARRYB[39][2] ), .SUM(\mult_44/SUMB[39][2] ) );
  FADDER \mult_44/S2_39_1  ( .CIN(\mult_44/ab[39][1] ), .IN0(
        \mult_44/CARRYB[38][1] ), .IN1(\mult_44/SUMB[38][2] ), .COUT(
        \mult_44/CARRYB[39][1] ), .SUM(\mult_44/SUMB[39][1] ) );
  FADDER \mult_44/S1_39_0  ( .CIN(\mult_44/ab[39][0] ), .IN0(
        \mult_44/CARRYB[38][0] ), .IN1(\mult_44/SUMB[38][1] ), .COUT(
        \mult_44/CARRYB[39][0] ), .SUM(clocal[39]) );
  FADDER \mult_44/S3_40_2  ( .CIN(\mult_44/ab[40][2] ), .IN0(
        \mult_44/CARRYB[39][2] ), .IN1(\mult_44/ab[39][3] ), .COUT(
        \mult_44/CARRYB[40][2] ), .SUM(\mult_44/SUMB[40][2] ) );
  FADDER \mult_44/S2_40_1  ( .CIN(\mult_44/ab[40][1] ), .IN0(
        \mult_44/CARRYB[39][1] ), .IN1(\mult_44/SUMB[39][2] ), .COUT(
        \mult_44/CARRYB[40][1] ), .SUM(\mult_44/SUMB[40][1] ) );
  FADDER \mult_44/S1_40_0  ( .CIN(\mult_44/ab[40][0] ), .IN0(
        \mult_44/CARRYB[39][0] ), .IN1(\mult_44/SUMB[39][1] ), .COUT(
        \mult_44/CARRYB[40][0] ), .SUM(clocal[40]) );
  FADDER \mult_44/S3_41_2  ( .CIN(\mult_44/ab[41][2] ), .IN0(
        \mult_44/CARRYB[40][2] ), .IN1(\mult_44/ab[40][3] ), .COUT(
        \mult_44/CARRYB[41][2] ), .SUM(\mult_44/SUMB[41][2] ) );
  FADDER \mult_44/S2_41_1  ( .CIN(\mult_44/ab[41][1] ), .IN0(
        \mult_44/CARRYB[40][1] ), .IN1(\mult_44/SUMB[40][2] ), .COUT(
        \mult_44/CARRYB[41][1] ), .SUM(\mult_44/SUMB[41][1] ) );
  FADDER \mult_44/S1_41_0  ( .CIN(\mult_44/ab[41][0] ), .IN0(
        \mult_44/CARRYB[40][0] ), .IN1(\mult_44/SUMB[40][1] ), .COUT(
        \mult_44/CARRYB[41][0] ), .SUM(clocal[41]) );
  FADDER \mult_44/S3_42_2  ( .CIN(\mult_44/ab[42][2] ), .IN0(
        \mult_44/CARRYB[41][2] ), .IN1(\mult_44/ab[41][3] ), .COUT(
        \mult_44/CARRYB[42][2] ), .SUM(\mult_44/SUMB[42][2] ) );
  FADDER \mult_44/S2_42_1  ( .CIN(\mult_44/ab[42][1] ), .IN0(
        \mult_44/CARRYB[41][1] ), .IN1(\mult_44/SUMB[41][2] ), .COUT(
        \mult_44/CARRYB[42][1] ), .SUM(\mult_44/SUMB[42][1] ) );
  FADDER \mult_44/S1_42_0  ( .CIN(\mult_44/ab[42][0] ), .IN0(
        \mult_44/CARRYB[41][0] ), .IN1(\mult_44/SUMB[41][1] ), .COUT(
        \mult_44/CARRYB[42][0] ), .SUM(clocal[42]) );
  FADDER \mult_44/S3_43_2  ( .CIN(\mult_44/ab[43][2] ), .IN0(
        \mult_44/CARRYB[42][2] ), .IN1(\mult_44/ab[42][3] ), .COUT(
        \mult_44/CARRYB[43][2] ), .SUM(\mult_44/SUMB[43][2] ) );
  FADDER \mult_44/S2_43_1  ( .CIN(\mult_44/ab[43][1] ), .IN0(
        \mult_44/CARRYB[42][1] ), .IN1(\mult_44/SUMB[42][2] ), .COUT(
        \mult_44/CARRYB[43][1] ), .SUM(\mult_44/SUMB[43][1] ) );
  FADDER \mult_44/S1_43_0  ( .CIN(\mult_44/ab[43][0] ), .IN0(
        \mult_44/CARRYB[42][0] ), .IN1(\mult_44/SUMB[42][1] ), .COUT(
        \mult_44/CARRYB[43][0] ), .SUM(clocal[43]) );
  FADDER \mult_44/S3_44_2  ( .CIN(\mult_44/ab[44][2] ), .IN0(
        \mult_44/CARRYB[43][2] ), .IN1(\mult_44/ab[43][3] ), .COUT(
        \mult_44/CARRYB[44][2] ), .SUM(\mult_44/SUMB[44][2] ) );
  FADDER \mult_44/S2_44_1  ( .CIN(\mult_44/ab[44][1] ), .IN0(
        \mult_44/CARRYB[43][1] ), .IN1(\mult_44/SUMB[43][2] ), .COUT(
        \mult_44/CARRYB[44][1] ), .SUM(\mult_44/SUMB[44][1] ) );
  FADDER \mult_44/S1_44_0  ( .CIN(\mult_44/ab[44][0] ), .IN0(
        \mult_44/CARRYB[43][0] ), .IN1(\mult_44/SUMB[43][1] ), .COUT(
        \mult_44/CARRYB[44][0] ), .SUM(clocal[44]) );
  FADDER \mult_44/S3_45_2  ( .CIN(\mult_44/ab[45][2] ), .IN0(
        \mult_44/CARRYB[44][2] ), .IN1(\mult_44/ab[44][3] ), .COUT(
        \mult_44/CARRYB[45][2] ), .SUM(\mult_44/SUMB[45][2] ) );
  FADDER \mult_44/S2_45_1  ( .CIN(\mult_44/ab[45][1] ), .IN0(
        \mult_44/CARRYB[44][1] ), .IN1(\mult_44/SUMB[44][2] ), .COUT(
        \mult_44/CARRYB[45][1] ), .SUM(\mult_44/SUMB[45][1] ) );
  FADDER \mult_44/S1_45_0  ( .CIN(\mult_44/ab[45][0] ), .IN0(
        \mult_44/CARRYB[44][0] ), .IN1(\mult_44/SUMB[44][1] ), .COUT(
        \mult_44/CARRYB[45][0] ), .SUM(clocal[45]) );
  FADDER \mult_44/S3_46_2  ( .CIN(\mult_44/ab[46][2] ), .IN0(
        \mult_44/CARRYB[45][2] ), .IN1(\mult_44/ab[45][3] ), .COUT(
        \mult_44/CARRYB[46][2] ), .SUM(\mult_44/SUMB[46][2] ) );
  FADDER \mult_44/S2_46_1  ( .CIN(\mult_44/ab[46][1] ), .IN0(
        \mult_44/CARRYB[45][1] ), .IN1(\mult_44/SUMB[45][2] ), .COUT(
        \mult_44/CARRYB[46][1] ), .SUM(\mult_44/SUMB[46][1] ) );
  FADDER \mult_44/S1_46_0  ( .CIN(\mult_44/ab[46][0] ), .IN0(
        \mult_44/CARRYB[45][0] ), .IN1(\mult_44/SUMB[45][1] ), .COUT(
        \mult_44/CARRYB[46][0] ), .SUM(clocal[46]) );
  FADDER \mult_44/S3_47_2  ( .CIN(\mult_44/ab[47][2] ), .IN0(
        \mult_44/CARRYB[46][2] ), .IN1(\mult_44/ab[46][3] ), .COUT(
        \mult_44/CARRYB[47][2] ), .SUM(\mult_44/SUMB[47][2] ) );
  FADDER \mult_44/S2_47_1  ( .CIN(\mult_44/ab[47][1] ), .IN0(
        \mult_44/CARRYB[46][1] ), .IN1(\mult_44/SUMB[46][2] ), .COUT(
        \mult_44/CARRYB[47][1] ), .SUM(\mult_44/SUMB[47][1] ) );
  FADDER \mult_44/S1_47_0  ( .CIN(\mult_44/ab[47][0] ), .IN0(
        \mult_44/CARRYB[46][0] ), .IN1(\mult_44/SUMB[46][1] ), .COUT(
        \mult_44/CARRYB[47][0] ), .SUM(clocal[47]) );
  FADDER \mult_44/S3_48_2  ( .CIN(\mult_44/ab[48][2] ), .IN0(
        \mult_44/CARRYB[47][2] ), .IN1(\mult_44/ab[47][3] ), .COUT(
        \mult_44/CARRYB[48][2] ), .SUM(\mult_44/SUMB[48][2] ) );
  FADDER \mult_44/S2_48_1  ( .CIN(\mult_44/ab[48][1] ), .IN0(
        \mult_44/CARRYB[47][1] ), .IN1(\mult_44/SUMB[47][2] ), .COUT(
        \mult_44/CARRYB[48][1] ), .SUM(\mult_44/SUMB[48][1] ) );
  FADDER \mult_44/S1_48_0  ( .CIN(\mult_44/ab[48][0] ), .IN0(
        \mult_44/CARRYB[47][0] ), .IN1(\mult_44/SUMB[47][1] ), .COUT(
        \mult_44/CARRYB[48][0] ), .SUM(clocal[48]) );
  FADDER \mult_44/S3_49_2  ( .CIN(\mult_44/ab[49][2] ), .IN0(
        \mult_44/CARRYB[48][2] ), .IN1(\mult_44/ab[48][3] ), .COUT(
        \mult_44/CARRYB[49][2] ), .SUM(\mult_44/SUMB[49][2] ) );
  FADDER \mult_44/S2_49_1  ( .CIN(\mult_44/ab[49][1] ), .IN0(
        \mult_44/CARRYB[48][1] ), .IN1(\mult_44/SUMB[48][2] ), .COUT(
        \mult_44/CARRYB[49][1] ), .SUM(\mult_44/SUMB[49][1] ) );
  FADDER \mult_44/S1_49_0  ( .CIN(\mult_44/ab[49][0] ), .IN0(
        \mult_44/CARRYB[48][0] ), .IN1(\mult_44/SUMB[48][1] ), .COUT(
        \mult_44/CARRYB[49][0] ), .SUM(clocal[49]) );
  FADDER \mult_44/S3_50_2  ( .CIN(\mult_44/ab[50][2] ), .IN0(
        \mult_44/CARRYB[49][2] ), .IN1(\mult_44/ab[49][3] ), .COUT(
        \mult_44/CARRYB[50][2] ), .SUM(\mult_44/SUMB[50][2] ) );
  FADDER \mult_44/S2_50_1  ( .CIN(\mult_44/ab[50][1] ), .IN0(
        \mult_44/CARRYB[49][1] ), .IN1(\mult_44/SUMB[49][2] ), .COUT(
        \mult_44/CARRYB[50][1] ), .SUM(\mult_44/SUMB[50][1] ) );
  FADDER \mult_44/S1_50_0  ( .CIN(\mult_44/ab[50][0] ), .IN0(
        \mult_44/CARRYB[49][0] ), .IN1(\mult_44/SUMB[49][1] ), .COUT(
        \mult_44/CARRYB[50][0] ), .SUM(clocal[50]) );
  FADDER \mult_44/S3_51_2  ( .CIN(\mult_44/ab[51][2] ), .IN0(
        \mult_44/CARRYB[50][2] ), .IN1(\mult_44/ab[50][3] ), .COUT(
        \mult_44/CARRYB[51][2] ), .SUM(\mult_44/SUMB[51][2] ) );
  FADDER \mult_44/S2_51_1  ( .CIN(\mult_44/ab[51][1] ), .IN0(
        \mult_44/CARRYB[50][1] ), .IN1(\mult_44/SUMB[50][2] ), .COUT(
        \mult_44/CARRYB[51][1] ), .SUM(\mult_44/SUMB[51][1] ) );
  FADDER \mult_44/S1_51_0  ( .CIN(\mult_44/ab[51][0] ), .IN0(
        \mult_44/CARRYB[50][0] ), .IN1(\mult_44/SUMB[50][1] ), .COUT(
        \mult_44/CARRYB[51][0] ), .SUM(clocal[51]) );
  FADDER \mult_44/S3_52_2  ( .CIN(\mult_44/ab[52][2] ), .IN0(
        \mult_44/CARRYB[51][2] ), .IN1(\mult_44/ab[51][3] ), .COUT(
        \mult_44/CARRYB[52][2] ), .SUM(\mult_44/SUMB[52][2] ) );
  FADDER \mult_44/S2_52_1  ( .CIN(\mult_44/ab[52][1] ), .IN0(
        \mult_44/CARRYB[51][1] ), .IN1(\mult_44/SUMB[51][2] ), .COUT(
        \mult_44/CARRYB[52][1] ), .SUM(\mult_44/SUMB[52][1] ) );
  FADDER \mult_44/S1_52_0  ( .CIN(\mult_44/ab[52][0] ), .IN0(
        \mult_44/CARRYB[51][0] ), .IN1(\mult_44/SUMB[51][1] ), .COUT(
        \mult_44/CARRYB[52][0] ), .SUM(clocal[52]) );
  FADDER \mult_44/S3_53_2  ( .CIN(\mult_44/ab[53][2] ), .IN0(
        \mult_44/CARRYB[52][2] ), .IN1(\mult_44/ab[52][3] ), .COUT(
        \mult_44/CARRYB[53][2] ), .SUM(\mult_44/SUMB[53][2] ) );
  FADDER \mult_44/S2_53_1  ( .CIN(\mult_44/ab[53][1] ), .IN0(
        \mult_44/CARRYB[52][1] ), .IN1(\mult_44/SUMB[52][2] ), .COUT(
        \mult_44/CARRYB[53][1] ), .SUM(\mult_44/SUMB[53][1] ) );
  FADDER \mult_44/S1_53_0  ( .CIN(\mult_44/ab[53][0] ), .IN0(
        \mult_44/CARRYB[52][0] ), .IN1(\mult_44/SUMB[52][1] ), .COUT(
        \mult_44/CARRYB[53][0] ), .SUM(clocal[53]) );
  FADDER \mult_44/S3_54_2  ( .CIN(\mult_44/ab[54][2] ), .IN0(
        \mult_44/CARRYB[53][2] ), .IN1(\mult_44/ab[53][3] ), .COUT(
        \mult_44/CARRYB[54][2] ), .SUM(\mult_44/SUMB[54][2] ) );
  FADDER \mult_44/S2_54_1  ( .CIN(\mult_44/ab[54][1] ), .IN0(
        \mult_44/CARRYB[53][1] ), .IN1(\mult_44/SUMB[53][2] ), .COUT(
        \mult_44/CARRYB[54][1] ), .SUM(\mult_44/SUMB[54][1] ) );
  FADDER \mult_44/S1_54_0  ( .CIN(\mult_44/ab[54][0] ), .IN0(
        \mult_44/CARRYB[53][0] ), .IN1(\mult_44/SUMB[53][1] ), .COUT(
        \mult_44/CARRYB[54][0] ), .SUM(clocal[54]) );
  FADDER \mult_44/S3_55_2  ( .CIN(\mult_44/ab[55][2] ), .IN0(
        \mult_44/CARRYB[54][2] ), .IN1(\mult_44/ab[54][3] ), .COUT(
        \mult_44/CARRYB[55][2] ), .SUM(\mult_44/SUMB[55][2] ) );
  FADDER \mult_44/S2_55_1  ( .CIN(\mult_44/ab[55][1] ), .IN0(
        \mult_44/CARRYB[54][1] ), .IN1(\mult_44/SUMB[54][2] ), .COUT(
        \mult_44/CARRYB[55][1] ), .SUM(\mult_44/SUMB[55][1] ) );
  FADDER \mult_44/S1_55_0  ( .CIN(\mult_44/ab[55][0] ), .IN0(
        \mult_44/CARRYB[54][0] ), .IN1(\mult_44/SUMB[54][1] ), .COUT(
        \mult_44/CARRYB[55][0] ), .SUM(clocal[55]) );
  FADDER \mult_44/S3_56_2  ( .CIN(\mult_44/ab[56][2] ), .IN0(
        \mult_44/CARRYB[55][2] ), .IN1(\mult_44/ab[55][3] ), .COUT(
        \mult_44/CARRYB[56][2] ), .SUM(\mult_44/SUMB[56][2] ) );
  FADDER \mult_44/S2_56_1  ( .CIN(\mult_44/ab[56][1] ), .IN0(
        \mult_44/CARRYB[55][1] ), .IN1(\mult_44/SUMB[55][2] ), .COUT(
        \mult_44/CARRYB[56][1] ), .SUM(\mult_44/SUMB[56][1] ) );
  FADDER \mult_44/S1_56_0  ( .CIN(\mult_44/ab[56][0] ), .IN0(
        \mult_44/CARRYB[55][0] ), .IN1(\mult_44/SUMB[55][1] ), .COUT(
        \mult_44/CARRYB[56][0] ), .SUM(clocal[56]) );
  FADDER \mult_44/S3_57_2  ( .CIN(\mult_44/ab[57][2] ), .IN0(
        \mult_44/CARRYB[56][2] ), .IN1(\mult_44/ab[56][3] ), .COUT(
        \mult_44/CARRYB[57][2] ), .SUM(\mult_44/SUMB[57][2] ) );
  FADDER \mult_44/S2_57_1  ( .CIN(\mult_44/ab[57][1] ), .IN0(
        \mult_44/CARRYB[56][1] ), .IN1(\mult_44/SUMB[56][2] ), .COUT(
        \mult_44/CARRYB[57][1] ), .SUM(\mult_44/SUMB[57][1] ) );
  FADDER \mult_44/S1_57_0  ( .CIN(\mult_44/ab[57][0] ), .IN0(
        \mult_44/CARRYB[56][0] ), .IN1(\mult_44/SUMB[56][1] ), .COUT(
        \mult_44/CARRYB[57][0] ), .SUM(clocal[57]) );
  FADDER \mult_44/S3_58_2  ( .CIN(\mult_44/ab[58][2] ), .IN0(
        \mult_44/CARRYB[57][2] ), .IN1(\mult_44/ab[57][3] ), .COUT(
        \mult_44/CARRYB[58][2] ), .SUM(\mult_44/SUMB[58][2] ) );
  FADDER \mult_44/S2_58_1  ( .CIN(\mult_44/ab[58][1] ), .IN0(
        \mult_44/CARRYB[57][1] ), .IN1(\mult_44/SUMB[57][2] ), .COUT(
        \mult_44/CARRYB[58][1] ), .SUM(\mult_44/SUMB[58][1] ) );
  FADDER \mult_44/S1_58_0  ( .CIN(\mult_44/ab[58][0] ), .IN0(
        \mult_44/CARRYB[57][0] ), .IN1(\mult_44/SUMB[57][1] ), .COUT(
        \mult_44/CARRYB[58][0] ), .SUM(clocal[58]) );
  FADDER \mult_44/S3_59_2  ( .CIN(\mult_44/ab[59][2] ), .IN0(
        \mult_44/CARRYB[58][2] ), .IN1(\mult_44/ab[58][3] ), .COUT(
        \mult_44/CARRYB[59][2] ), .SUM(\mult_44/SUMB[59][2] ) );
  FADDER \mult_44/S2_59_1  ( .CIN(\mult_44/ab[59][1] ), .IN0(
        \mult_44/CARRYB[58][1] ), .IN1(\mult_44/SUMB[58][2] ), .COUT(
        \mult_44/CARRYB[59][1] ), .SUM(\mult_44/SUMB[59][1] ) );
  FADDER \mult_44/S1_59_0  ( .CIN(\mult_44/ab[59][0] ), .IN0(
        \mult_44/CARRYB[58][0] ), .IN1(\mult_44/SUMB[58][1] ), .COUT(
        \mult_44/CARRYB[59][0] ), .SUM(clocal[59]) );
  FADDER \mult_44/S3_60_2  ( .CIN(\mult_44/ab[60][2] ), .IN0(
        \mult_44/CARRYB[59][2] ), .IN1(\mult_44/ab[59][3] ), .COUT(
        \mult_44/CARRYB[60][2] ), .SUM(\mult_44/SUMB[60][2] ) );
  FADDER \mult_44/S2_60_1  ( .CIN(\mult_44/ab[60][1] ), .IN0(
        \mult_44/CARRYB[59][1] ), .IN1(\mult_44/SUMB[59][2] ), .COUT(
        \mult_44/CARRYB[60][1] ), .SUM(\mult_44/SUMB[60][1] ) );
  FADDER \mult_44/S1_60_0  ( .CIN(\mult_44/ab[60][0] ), .IN0(
        \mult_44/CARRYB[59][0] ), .IN1(\mult_44/SUMB[59][1] ), .COUT(
        \mult_44/CARRYB[60][0] ), .SUM(clocal[60]) );
  FADDER \mult_44/S3_61_2  ( .CIN(\mult_44/ab[61][2] ), .IN0(
        \mult_44/CARRYB[60][2] ), .IN1(\mult_44/ab[60][3] ), .SUM(
        \mult_44/SUMB[61][2] ) );
  FADDER \mult_44/S2_61_1  ( .CIN(\mult_44/ab[61][1] ), .IN0(
        \mult_44/CARRYB[60][1] ), .IN1(\mult_44/SUMB[60][2] ), .COUT(
        \mult_44/CARRYB[61][1] ), .SUM(\mult_44/SUMB[61][1] ) );
  FADDER \mult_44/S1_61_0  ( .CIN(\mult_44/ab[61][0] ), .IN0(
        \mult_44/CARRYB[60][0] ), .IN1(\mult_44/SUMB[60][1] ), .COUT(
        \mult_44/CARRYB[61][0] ), .SUM(clocal[61]) );
  FADDER \mult_44/S2_62_1  ( .CIN(\mult_44/ab[62][1] ), .IN0(
        \mult_44/CARRYB[61][1] ), .IN1(\mult_44/SUMB[61][2] ), .SUM(
        \mult_44/SUMB[62][1] ) );
  FADDER \mult_44/S1_62_0  ( .CIN(\mult_44/ab[62][0] ), .IN0(
        \mult_44/CARRYB[61][0] ), .IN1(\mult_44/SUMB[61][1] ), .COUT(
        \mult_44/CARRYB[62][0] ), .SUM(clocal[62]) );
  FADDER \mult_44/S4_0  ( .CIN(\mult_44/ab[63][0] ), .IN0(
        \mult_44/CARRYB[62][0] ), .IN1(\mult_44/SUMB[62][1] ), .SUM(
        \mult_44/SUMB[63][0] ) );
  MUX U128 ( .IN0(clocal[56]), .IN1(n142), .SEL(n143), .F(n138) );
  MUX U129 ( .IN0(clocal[52]), .IN1(n154), .SEL(n155), .F(n150) );
  MUX U130 ( .IN0(clocal[48]), .IN1(n167), .SEL(n168), .F(n162) );
  MUX U131 ( .IN0(clocal[44]), .IN1(n179), .SEL(n180), .F(n175) );
  MUX U132 ( .IN0(clocal[40]), .IN1(n191), .SEL(n192), .F(n187) );
  MUX U133 ( .IN0(clocal[36]), .IN1(n203), .SEL(n204), .F(n199) );
  MUX U134 ( .IN0(clocal[32]), .IN1(n215), .SEL(n216), .F(n211) );
  MUX U135 ( .IN0(clocal[28]), .IN1(n227), .SEL(n228), .F(n223) );
  MUX U136 ( .IN0(clocal[24]), .IN1(n239), .SEL(n240), .F(n235) );
  MUX U137 ( .IN0(clocal[20]), .IN1(n251), .SEL(n252), .F(n247) );
  MUX U138 ( .IN0(clocal[16]), .IN1(n263), .SEL(n264), .F(n259) );
  MUX U139 ( .IN0(clocal[12]), .IN1(n275), .SEL(n276), .F(n271) );
  MUX U140 ( .IN0(clocal[8]), .IN1(n286), .SEL(n123), .F(n283) );
  MUX U141 ( .IN0(clocal[4]), .IN1(n294), .SEL(n166), .F(n291) );
  MUX U142 ( .IN0(clocal[55]), .IN1(n144), .SEL(n145), .F(n142) );
  MUX U143 ( .IN0(clocal[51]), .IN1(n156), .SEL(n157), .F(n154) );
  MUX U144 ( .IN0(clocal[47]), .IN1(n169), .SEL(n170), .F(n167) );
  MUX U145 ( .IN0(clocal[43]), .IN1(n181), .SEL(n182), .F(n179) );
  MUX U146 ( .IN0(clocal[39]), .IN1(n193), .SEL(n194), .F(n191) );
  MUX U147 ( .IN0(clocal[35]), .IN1(n205), .SEL(n206), .F(n203) );
  MUX U148 ( .IN0(clocal[31]), .IN1(n217), .SEL(n218), .F(n215) );
  MUX U149 ( .IN0(clocal[27]), .IN1(n229), .SEL(n230), .F(n227) );
  MUX U150 ( .IN0(clocal[23]), .IN1(n241), .SEL(n242), .F(n239) );
  MUX U151 ( .IN0(clocal[19]), .IN1(n253), .SEL(n254), .F(n251) );
  MUX U152 ( .IN0(clocal[15]), .IN1(n265), .SEL(n266), .F(n263) );
  MUX U153 ( .IN0(clocal[11]), .IN1(n277), .SEL(n278), .F(n275) );
  MUX U154 ( .IN0(clocal[7]), .IN1(n287), .SEL(n124), .F(n286) );
  MUX U155 ( .IN0(\mult_44/PROD1[3] ), .IN1(n295), .SEL(n296), .F(n294) );
  MUX U156 ( .IN0(clocal[59]), .IN1(n131), .SEL(n132), .F(n130) );
  XNOR U157 ( .A(n295), .B(sreg[67]), .Z(n296) );
  XNOR U158 ( .A(n138), .B(sreg[121]), .Z(n141) );
  XNOR U159 ( .A(n146), .B(sreg[118]), .Z(n149) );
  XNOR U160 ( .A(n156), .B(sreg[115]), .Z(n157) );
  XNOR U161 ( .A(n167), .B(sreg[112]), .Z(n168) );
  XNOR U162 ( .A(n175), .B(sreg[109]), .Z(n178) );
  XNOR U163 ( .A(n183), .B(sreg[106]), .Z(n186) );
  XNOR U164 ( .A(n193), .B(sreg[103]), .Z(n194) );
  XNOR U165 ( .A(n203), .B(sreg[100]), .Z(n204) );
  XNOR U166 ( .A(n211), .B(sreg[97]), .Z(n214) );
  XNOR U167 ( .A(n219), .B(sreg[94]), .Z(n222) );
  XNOR U168 ( .A(n229), .B(sreg[91]), .Z(n230) );
  XNOR U169 ( .A(n239), .B(sreg[88]), .Z(n240) );
  XNOR U170 ( .A(n247), .B(sreg[85]), .Z(n250) );
  XNOR U171 ( .A(n255), .B(sreg[82]), .Z(n258) );
  XNOR U172 ( .A(n265), .B(sreg[79]), .Z(n266) );
  XNOR U173 ( .A(n275), .B(sreg[76]), .Z(n276) );
  XNOR U174 ( .A(n283), .B(sreg[73]), .Z(n122) );
  XNOR U175 ( .A(n288), .B(sreg[70]), .Z(n125) );
  XNOR U176 ( .A(n297), .B(sreg[66]), .Z(n300) );
  XNOR U177 ( .A(n131), .B(sreg[123]), .Z(n132) );
  XNOR U178 ( .A(n142), .B(sreg[120]), .Z(n143) );
  XNOR U179 ( .A(n150), .B(sreg[117]), .Z(n153) );
  XNOR U180 ( .A(n158), .B(sreg[114]), .Z(n161) );
  XNOR U181 ( .A(n169), .B(sreg[111]), .Z(n170) );
  XNOR U182 ( .A(n179), .B(sreg[108]), .Z(n180) );
  XNOR U183 ( .A(n187), .B(sreg[105]), .Z(n190) );
  XNOR U184 ( .A(n195), .B(sreg[102]), .Z(n198) );
  XNOR U185 ( .A(n205), .B(sreg[99]), .Z(n206) );
  XNOR U186 ( .A(n215), .B(sreg[96]), .Z(n216) );
  XNOR U187 ( .A(n223), .B(sreg[93]), .Z(n226) );
  XNOR U188 ( .A(n231), .B(sreg[90]), .Z(n234) );
  XNOR U189 ( .A(n241), .B(sreg[87]), .Z(n242) );
  XNOR U190 ( .A(n251), .B(sreg[84]), .Z(n252) );
  XNOR U191 ( .A(n259), .B(sreg[81]), .Z(n262) );
  XNOR U192 ( .A(n267), .B(sreg[78]), .Z(n270) );
  XNOR U193 ( .A(n277), .B(sreg[75]), .Z(n278) );
  XNOR U194 ( .A(n286), .B(sreg[72]), .Z(n123) );
  XNOR U195 ( .A(n291), .B(sreg[69]), .Z(n133) );
  XNOR U196 ( .A(n134), .B(sreg[122]), .Z(n137) );
  XNOR U197 ( .A(n144), .B(sreg[119]), .Z(n145) );
  XNOR U198 ( .A(n154), .B(sreg[116]), .Z(n155) );
  XNOR U199 ( .A(n162), .B(sreg[113]), .Z(n165) );
  XNOR U200 ( .A(n171), .B(sreg[110]), .Z(n174) );
  XNOR U201 ( .A(n181), .B(sreg[107]), .Z(n182) );
  XNOR U202 ( .A(n191), .B(sreg[104]), .Z(n192) );
  XNOR U203 ( .A(n199), .B(sreg[101]), .Z(n202) );
  XNOR U204 ( .A(n207), .B(sreg[98]), .Z(n210) );
  XNOR U205 ( .A(n217), .B(sreg[95]), .Z(n218) );
  XNOR U206 ( .A(n227), .B(sreg[92]), .Z(n228) );
  XNOR U207 ( .A(n235), .B(sreg[89]), .Z(n238) );
  XNOR U208 ( .A(n243), .B(sreg[86]), .Z(n246) );
  XNOR U209 ( .A(n253), .B(sreg[83]), .Z(n254) );
  XNOR U210 ( .A(n263), .B(sreg[80]), .Z(n264) );
  XNOR U211 ( .A(n271), .B(sreg[77]), .Z(n274) );
  XNOR U212 ( .A(n279), .B(sreg[74]), .Z(n282) );
  XNOR U213 ( .A(n287), .B(sreg[71]), .Z(n124) );
  XNOR U214 ( .A(n294), .B(sreg[68]), .Z(n166) );
  AND U215 ( .A(\mult_44/ab[0][1] ), .B(\mult_44/ab[1][0] ), .Z(
        \mult_44/CARRYB[1][0] ) );
  XOR U216 ( .A(\mult_44/ab[0][1] ), .B(\mult_44/ab[1][0] ), .Z(clocal[1]) );
  AND U217 ( .A(\mult_44/ab[1][1] ), .B(\mult_44/ab[0][2] ), .Z(
        \mult_44/CARRYB[1][1] ) );
  XOR U218 ( .A(\mult_44/ab[0][2] ), .B(\mult_44/ab[1][1] ), .Z(
        \mult_44/SUMB[1][1] ) );
  AND U219 ( .A(\mult_44/ab[1][2] ), .B(\mult_44/ab[0][3] ), .Z(
        \mult_44/CARRYB[1][2] ) );
  XOR U220 ( .A(\mult_44/ab[0][3] ), .B(\mult_44/ab[1][2] ), .Z(
        \mult_44/SUMB[1][2] ) );
  XNOR U221 ( .A(clocal[9]), .B(n122), .Z(swire[9]) );
  XNOR U222 ( .A(clocal[8]), .B(n123), .Z(swire[8]) );
  XNOR U223 ( .A(clocal[7]), .B(n124), .Z(swire[7]) );
  XNOR U224 ( .A(clocal[6]), .B(n125), .Z(swire[6]) );
  XOR U225 ( .A(n126), .B(n127), .Z(swire[63]) );
  XOR U226 ( .A(\mult_44/SUMB[63][0] ), .B(n128), .Z(n127) );
  ANDN U227 ( .B(n126), .A(clocal[62]), .Z(n128) );
  XOR U228 ( .A(clocal[62]), .B(n126), .Z(swire[62]) );
  ANDN U229 ( .B(clocal[61]), .A(n129), .Z(n126) );
  XNOR U230 ( .A(clocal[61]), .B(n129), .Z(swire[61]) );
  NAND U231 ( .A(n130), .B(clocal[60]), .Z(n129) );
  XOR U232 ( .A(clocal[60]), .B(n130), .Z(swire[60]) );
  XNOR U233 ( .A(clocal[5]), .B(n133), .Z(swire[5]) );
  XNOR U234 ( .A(clocal[59]), .B(n132), .Z(swire[59]) );
  XOR U235 ( .A(n134), .B(n135), .Z(n131) );
  ANDN U236 ( .B(n136), .A(n137), .Z(n135) );
  XOR U237 ( .A(clocal[58]), .B(n134), .Z(n136) );
  XNOR U238 ( .A(clocal[58]), .B(n137), .Z(swire[58]) );
  XOR U239 ( .A(n138), .B(n139), .Z(n134) );
  ANDN U240 ( .B(n140), .A(n141), .Z(n139) );
  XOR U241 ( .A(clocal[57]), .B(n138), .Z(n140) );
  XNOR U242 ( .A(clocal[57]), .B(n141), .Z(swire[57]) );
  XNOR U243 ( .A(clocal[56]), .B(n143), .Z(swire[56]) );
  XNOR U244 ( .A(clocal[55]), .B(n145), .Z(swire[55]) );
  XOR U245 ( .A(n146), .B(n147), .Z(n144) );
  ANDN U246 ( .B(n148), .A(n149), .Z(n147) );
  XOR U247 ( .A(clocal[54]), .B(n146), .Z(n148) );
  XNOR U248 ( .A(clocal[54]), .B(n149), .Z(swire[54]) );
  XOR U249 ( .A(n150), .B(n151), .Z(n146) );
  ANDN U250 ( .B(n152), .A(n153), .Z(n151) );
  XOR U251 ( .A(clocal[53]), .B(n150), .Z(n152) );
  XNOR U252 ( .A(clocal[53]), .B(n153), .Z(swire[53]) );
  XNOR U253 ( .A(clocal[52]), .B(n155), .Z(swire[52]) );
  XNOR U254 ( .A(clocal[51]), .B(n157), .Z(swire[51]) );
  XOR U255 ( .A(n158), .B(n159), .Z(n156) );
  ANDN U256 ( .B(n160), .A(n161), .Z(n159) );
  XOR U257 ( .A(clocal[50]), .B(n158), .Z(n160) );
  XNOR U258 ( .A(clocal[50]), .B(n161), .Z(swire[50]) );
  XOR U259 ( .A(n162), .B(n163), .Z(n158) );
  ANDN U260 ( .B(n164), .A(n165), .Z(n163) );
  XOR U261 ( .A(clocal[49]), .B(n162), .Z(n164) );
  XNOR U262 ( .A(clocal[4]), .B(n166), .Z(swire[4]) );
  XNOR U263 ( .A(clocal[49]), .B(n165), .Z(swire[49]) );
  XNOR U264 ( .A(clocal[48]), .B(n168), .Z(swire[48]) );
  XNOR U265 ( .A(clocal[47]), .B(n170), .Z(swire[47]) );
  XOR U266 ( .A(n171), .B(n172), .Z(n169) );
  ANDN U267 ( .B(n173), .A(n174), .Z(n172) );
  XOR U268 ( .A(clocal[46]), .B(n171), .Z(n173) );
  XNOR U269 ( .A(clocal[46]), .B(n174), .Z(swire[46]) );
  XOR U270 ( .A(n175), .B(n176), .Z(n171) );
  ANDN U271 ( .B(n177), .A(n178), .Z(n176) );
  XOR U272 ( .A(clocal[45]), .B(n175), .Z(n177) );
  XNOR U273 ( .A(clocal[45]), .B(n178), .Z(swire[45]) );
  XNOR U274 ( .A(clocal[44]), .B(n180), .Z(swire[44]) );
  XNOR U275 ( .A(clocal[43]), .B(n182), .Z(swire[43]) );
  XOR U276 ( .A(n183), .B(n184), .Z(n181) );
  ANDN U277 ( .B(n185), .A(n186), .Z(n184) );
  XOR U278 ( .A(clocal[42]), .B(n183), .Z(n185) );
  XNOR U279 ( .A(clocal[42]), .B(n186), .Z(swire[42]) );
  XOR U280 ( .A(n187), .B(n188), .Z(n183) );
  ANDN U281 ( .B(n189), .A(n190), .Z(n188) );
  XOR U282 ( .A(clocal[41]), .B(n187), .Z(n189) );
  XNOR U283 ( .A(clocal[41]), .B(n190), .Z(swire[41]) );
  XNOR U284 ( .A(clocal[40]), .B(n192), .Z(swire[40]) );
  XNOR U285 ( .A(clocal[39]), .B(n194), .Z(swire[39]) );
  XOR U286 ( .A(n195), .B(n196), .Z(n193) );
  ANDN U287 ( .B(n197), .A(n198), .Z(n196) );
  XOR U288 ( .A(clocal[38]), .B(n195), .Z(n197) );
  XNOR U289 ( .A(clocal[38]), .B(n198), .Z(swire[38]) );
  XOR U290 ( .A(n199), .B(n200), .Z(n195) );
  ANDN U291 ( .B(n201), .A(n202), .Z(n200) );
  XOR U292 ( .A(clocal[37]), .B(n199), .Z(n201) );
  XNOR U293 ( .A(clocal[37]), .B(n202), .Z(swire[37]) );
  XNOR U294 ( .A(clocal[36]), .B(n204), .Z(swire[36]) );
  XNOR U295 ( .A(clocal[35]), .B(n206), .Z(swire[35]) );
  XOR U296 ( .A(n207), .B(n208), .Z(n205) );
  ANDN U297 ( .B(n209), .A(n210), .Z(n208) );
  XOR U298 ( .A(clocal[34]), .B(n207), .Z(n209) );
  XNOR U299 ( .A(clocal[34]), .B(n210), .Z(swire[34]) );
  XOR U300 ( .A(n211), .B(n212), .Z(n207) );
  ANDN U301 ( .B(n213), .A(n214), .Z(n212) );
  XOR U302 ( .A(clocal[33]), .B(n211), .Z(n213) );
  XNOR U303 ( .A(clocal[33]), .B(n214), .Z(swire[33]) );
  XNOR U304 ( .A(clocal[32]), .B(n216), .Z(swire[32]) );
  XNOR U305 ( .A(clocal[31]), .B(n218), .Z(swire[31]) );
  XOR U306 ( .A(n219), .B(n220), .Z(n217) );
  ANDN U307 ( .B(n221), .A(n222), .Z(n220) );
  XOR U308 ( .A(clocal[30]), .B(n219), .Z(n221) );
  XNOR U309 ( .A(clocal[30]), .B(n222), .Z(swire[30]) );
  XOR U310 ( .A(n223), .B(n224), .Z(n219) );
  ANDN U311 ( .B(n225), .A(n226), .Z(n224) );
  XOR U312 ( .A(clocal[29]), .B(n223), .Z(n225) );
  XNOR U313 ( .A(clocal[29]), .B(n226), .Z(swire[29]) );
  XNOR U314 ( .A(clocal[28]), .B(n228), .Z(swire[28]) );
  XNOR U315 ( .A(clocal[27]), .B(n230), .Z(swire[27]) );
  XOR U316 ( .A(n231), .B(n232), .Z(n229) );
  ANDN U317 ( .B(n233), .A(n234), .Z(n232) );
  XOR U318 ( .A(clocal[26]), .B(n231), .Z(n233) );
  XNOR U319 ( .A(clocal[26]), .B(n234), .Z(swire[26]) );
  XOR U320 ( .A(n235), .B(n236), .Z(n231) );
  ANDN U321 ( .B(n237), .A(n238), .Z(n236) );
  XOR U322 ( .A(clocal[25]), .B(n235), .Z(n237) );
  XNOR U323 ( .A(clocal[25]), .B(n238), .Z(swire[25]) );
  XNOR U324 ( .A(clocal[24]), .B(n240), .Z(swire[24]) );
  XNOR U325 ( .A(clocal[23]), .B(n242), .Z(swire[23]) );
  XOR U326 ( .A(n243), .B(n244), .Z(n241) );
  ANDN U327 ( .B(n245), .A(n246), .Z(n244) );
  XOR U328 ( .A(clocal[22]), .B(n243), .Z(n245) );
  XNOR U329 ( .A(clocal[22]), .B(n246), .Z(swire[22]) );
  XOR U330 ( .A(n247), .B(n248), .Z(n243) );
  ANDN U331 ( .B(n249), .A(n250), .Z(n248) );
  XOR U332 ( .A(clocal[21]), .B(n247), .Z(n249) );
  XNOR U333 ( .A(clocal[21]), .B(n250), .Z(swire[21]) );
  XNOR U334 ( .A(clocal[20]), .B(n252), .Z(swire[20]) );
  XNOR U335 ( .A(clocal[19]), .B(n254), .Z(swire[19]) );
  XOR U336 ( .A(n255), .B(n256), .Z(n253) );
  ANDN U337 ( .B(n257), .A(n258), .Z(n256) );
  XOR U338 ( .A(clocal[18]), .B(n255), .Z(n257) );
  XNOR U339 ( .A(clocal[18]), .B(n258), .Z(swire[18]) );
  XOR U340 ( .A(n259), .B(n260), .Z(n255) );
  ANDN U341 ( .B(n261), .A(n262), .Z(n260) );
  XOR U342 ( .A(clocal[17]), .B(n259), .Z(n261) );
  XNOR U343 ( .A(clocal[17]), .B(n262), .Z(swire[17]) );
  XNOR U344 ( .A(clocal[16]), .B(n264), .Z(swire[16]) );
  XNOR U345 ( .A(clocal[15]), .B(n266), .Z(swire[15]) );
  XOR U346 ( .A(n267), .B(n268), .Z(n265) );
  ANDN U347 ( .B(n269), .A(n270), .Z(n268) );
  XOR U348 ( .A(clocal[14]), .B(n267), .Z(n269) );
  XNOR U349 ( .A(clocal[14]), .B(n270), .Z(swire[14]) );
  XOR U350 ( .A(n271), .B(n272), .Z(n267) );
  ANDN U351 ( .B(n273), .A(n274), .Z(n272) );
  XOR U352 ( .A(clocal[13]), .B(n271), .Z(n273) );
  XNOR U353 ( .A(clocal[13]), .B(n274), .Z(swire[13]) );
  XNOR U354 ( .A(clocal[12]), .B(n276), .Z(swire[12]) );
  XNOR U355 ( .A(clocal[11]), .B(n278), .Z(swire[11]) );
  XOR U356 ( .A(n279), .B(n280), .Z(n277) );
  ANDN U357 ( .B(n281), .A(n282), .Z(n280) );
  XOR U358 ( .A(clocal[10]), .B(n279), .Z(n281) );
  XNOR U359 ( .A(clocal[10]), .B(n282), .Z(swire[10]) );
  XOR U360 ( .A(n283), .B(n284), .Z(n279) );
  ANDN U361 ( .B(n285), .A(n122), .Z(n284) );
  XOR U362 ( .A(clocal[9]), .B(n283), .Z(n285) );
  XOR U363 ( .A(n288), .B(n289), .Z(n287) );
  ANDN U364 ( .B(n290), .A(n125), .Z(n289) );
  XOR U365 ( .A(clocal[6]), .B(n288), .Z(n290) );
  XOR U366 ( .A(n291), .B(n292), .Z(n288) );
  ANDN U367 ( .B(n293), .A(n133), .Z(n292) );
  XOR U368 ( .A(clocal[5]), .B(n291), .Z(n293) );
  AND U369 ( .A(a[9]), .B(b[3]), .Z(\mult_44/ab[9][3] ) );
  AND U370 ( .A(a[9]), .B(b[2]), .Z(\mult_44/ab[9][2] ) );
  AND U371 ( .A(a[9]), .B(b[1]), .Z(\mult_44/ab[9][1] ) );
  AND U372 ( .A(b[0]), .B(a[9]), .Z(\mult_44/ab[9][0] ) );
  AND U373 ( .A(b[3]), .B(a[8]), .Z(\mult_44/ab[8][3] ) );
  AND U374 ( .A(b[2]), .B(a[8]), .Z(\mult_44/ab[8][2] ) );
  AND U375 ( .A(b[1]), .B(a[8]), .Z(\mult_44/ab[8][1] ) );
  AND U376 ( .A(a[8]), .B(b[0]), .Z(\mult_44/ab[8][0] ) );
  AND U377 ( .A(b[3]), .B(a[7]), .Z(\mult_44/ab[7][3] ) );
  AND U378 ( .A(b[2]), .B(a[7]), .Z(\mult_44/ab[7][2] ) );
  AND U379 ( .A(b[1]), .B(a[7]), .Z(\mult_44/ab[7][1] ) );
  AND U380 ( .A(a[7]), .B(b[0]), .Z(\mult_44/ab[7][0] ) );
  AND U381 ( .A(b[3]), .B(a[6]), .Z(\mult_44/ab[6][3] ) );
  AND U382 ( .A(b[2]), .B(a[6]), .Z(\mult_44/ab[6][2] ) );
  AND U383 ( .A(b[1]), .B(a[6]), .Z(\mult_44/ab[6][1] ) );
  AND U384 ( .A(a[6]), .B(b[0]), .Z(\mult_44/ab[6][0] ) );
  AND U385 ( .A(a[63]), .B(b[0]), .Z(\mult_44/ab[63][0] ) );
  AND U386 ( .A(b[1]), .B(a[62]), .Z(\mult_44/ab[62][1] ) );
  AND U387 ( .A(a[62]), .B(b[0]), .Z(\mult_44/ab[62][0] ) );
  AND U388 ( .A(b[2]), .B(a[61]), .Z(\mult_44/ab[61][2] ) );
  AND U389 ( .A(b[1]), .B(a[61]), .Z(\mult_44/ab[61][1] ) );
  AND U390 ( .A(a[61]), .B(b[0]), .Z(\mult_44/ab[61][0] ) );
  AND U391 ( .A(b[3]), .B(a[60]), .Z(\mult_44/ab[60][3] ) );
  AND U392 ( .A(b[2]), .B(a[60]), .Z(\mult_44/ab[60][2] ) );
  AND U393 ( .A(b[1]), .B(a[60]), .Z(\mult_44/ab[60][1] ) );
  AND U394 ( .A(a[60]), .B(b[0]), .Z(\mult_44/ab[60][0] ) );
  AND U395 ( .A(b[3]), .B(a[5]), .Z(\mult_44/ab[5][3] ) );
  AND U396 ( .A(b[2]), .B(a[5]), .Z(\mult_44/ab[5][2] ) );
  AND U397 ( .A(b[1]), .B(a[5]), .Z(\mult_44/ab[5][1] ) );
  AND U398 ( .A(a[5]), .B(b[0]), .Z(\mult_44/ab[5][0] ) );
  AND U399 ( .A(b[3]), .B(a[59]), .Z(\mult_44/ab[59][3] ) );
  AND U400 ( .A(b[2]), .B(a[59]), .Z(\mult_44/ab[59][2] ) );
  AND U401 ( .A(b[1]), .B(a[59]), .Z(\mult_44/ab[59][1] ) );
  AND U402 ( .A(a[59]), .B(b[0]), .Z(\mult_44/ab[59][0] ) );
  AND U403 ( .A(b[3]), .B(a[58]), .Z(\mult_44/ab[58][3] ) );
  AND U404 ( .A(b[2]), .B(a[58]), .Z(\mult_44/ab[58][2] ) );
  AND U405 ( .A(b[1]), .B(a[58]), .Z(\mult_44/ab[58][1] ) );
  AND U406 ( .A(a[58]), .B(b[0]), .Z(\mult_44/ab[58][0] ) );
  AND U407 ( .A(b[3]), .B(a[57]), .Z(\mult_44/ab[57][3] ) );
  AND U408 ( .A(b[2]), .B(a[57]), .Z(\mult_44/ab[57][2] ) );
  AND U409 ( .A(b[1]), .B(a[57]), .Z(\mult_44/ab[57][1] ) );
  AND U410 ( .A(a[57]), .B(b[0]), .Z(\mult_44/ab[57][0] ) );
  AND U411 ( .A(b[3]), .B(a[56]), .Z(\mult_44/ab[56][3] ) );
  AND U412 ( .A(b[2]), .B(a[56]), .Z(\mult_44/ab[56][2] ) );
  AND U413 ( .A(b[1]), .B(a[56]), .Z(\mult_44/ab[56][1] ) );
  AND U414 ( .A(a[56]), .B(b[0]), .Z(\mult_44/ab[56][0] ) );
  AND U415 ( .A(b[3]), .B(a[55]), .Z(\mult_44/ab[55][3] ) );
  AND U416 ( .A(b[2]), .B(a[55]), .Z(\mult_44/ab[55][2] ) );
  AND U417 ( .A(b[1]), .B(a[55]), .Z(\mult_44/ab[55][1] ) );
  AND U418 ( .A(a[55]), .B(b[0]), .Z(\mult_44/ab[55][0] ) );
  AND U419 ( .A(b[3]), .B(a[54]), .Z(\mult_44/ab[54][3] ) );
  AND U420 ( .A(b[2]), .B(a[54]), .Z(\mult_44/ab[54][2] ) );
  AND U421 ( .A(b[1]), .B(a[54]), .Z(\mult_44/ab[54][1] ) );
  AND U422 ( .A(a[54]), .B(b[0]), .Z(\mult_44/ab[54][0] ) );
  AND U423 ( .A(b[3]), .B(a[53]), .Z(\mult_44/ab[53][3] ) );
  AND U424 ( .A(b[2]), .B(a[53]), .Z(\mult_44/ab[53][2] ) );
  AND U425 ( .A(b[1]), .B(a[53]), .Z(\mult_44/ab[53][1] ) );
  AND U426 ( .A(a[53]), .B(b[0]), .Z(\mult_44/ab[53][0] ) );
  AND U427 ( .A(b[3]), .B(a[52]), .Z(\mult_44/ab[52][3] ) );
  AND U428 ( .A(b[2]), .B(a[52]), .Z(\mult_44/ab[52][2] ) );
  AND U429 ( .A(b[1]), .B(a[52]), .Z(\mult_44/ab[52][1] ) );
  AND U430 ( .A(a[52]), .B(b[0]), .Z(\mult_44/ab[52][0] ) );
  AND U431 ( .A(b[3]), .B(a[51]), .Z(\mult_44/ab[51][3] ) );
  AND U432 ( .A(b[2]), .B(a[51]), .Z(\mult_44/ab[51][2] ) );
  AND U433 ( .A(b[1]), .B(a[51]), .Z(\mult_44/ab[51][1] ) );
  AND U434 ( .A(a[51]), .B(b[0]), .Z(\mult_44/ab[51][0] ) );
  AND U435 ( .A(b[3]), .B(a[50]), .Z(\mult_44/ab[50][3] ) );
  AND U436 ( .A(b[2]), .B(a[50]), .Z(\mult_44/ab[50][2] ) );
  AND U437 ( .A(b[1]), .B(a[50]), .Z(\mult_44/ab[50][1] ) );
  AND U438 ( .A(a[50]), .B(b[0]), .Z(\mult_44/ab[50][0] ) );
  AND U439 ( .A(b[3]), .B(a[4]), .Z(\mult_44/ab[4][3] ) );
  AND U440 ( .A(b[2]), .B(a[4]), .Z(\mult_44/ab[4][2] ) );
  AND U441 ( .A(b[1]), .B(a[4]), .Z(\mult_44/ab[4][1] ) );
  AND U442 ( .A(a[4]), .B(b[0]), .Z(\mult_44/ab[4][0] ) );
  AND U443 ( .A(b[3]), .B(a[49]), .Z(\mult_44/ab[49][3] ) );
  AND U444 ( .A(b[2]), .B(a[49]), .Z(\mult_44/ab[49][2] ) );
  AND U445 ( .A(b[1]), .B(a[49]), .Z(\mult_44/ab[49][1] ) );
  AND U446 ( .A(a[49]), .B(b[0]), .Z(\mult_44/ab[49][0] ) );
  AND U447 ( .A(b[3]), .B(a[48]), .Z(\mult_44/ab[48][3] ) );
  AND U448 ( .A(b[2]), .B(a[48]), .Z(\mult_44/ab[48][2] ) );
  AND U449 ( .A(b[1]), .B(a[48]), .Z(\mult_44/ab[48][1] ) );
  AND U450 ( .A(a[48]), .B(b[0]), .Z(\mult_44/ab[48][0] ) );
  AND U451 ( .A(b[3]), .B(a[47]), .Z(\mult_44/ab[47][3] ) );
  AND U452 ( .A(b[2]), .B(a[47]), .Z(\mult_44/ab[47][2] ) );
  AND U453 ( .A(b[1]), .B(a[47]), .Z(\mult_44/ab[47][1] ) );
  AND U454 ( .A(a[47]), .B(b[0]), .Z(\mult_44/ab[47][0] ) );
  AND U455 ( .A(b[3]), .B(a[46]), .Z(\mult_44/ab[46][3] ) );
  AND U456 ( .A(b[2]), .B(a[46]), .Z(\mult_44/ab[46][2] ) );
  AND U457 ( .A(b[1]), .B(a[46]), .Z(\mult_44/ab[46][1] ) );
  AND U458 ( .A(a[46]), .B(b[0]), .Z(\mult_44/ab[46][0] ) );
  AND U459 ( .A(b[3]), .B(a[45]), .Z(\mult_44/ab[45][3] ) );
  AND U460 ( .A(b[2]), .B(a[45]), .Z(\mult_44/ab[45][2] ) );
  AND U461 ( .A(b[1]), .B(a[45]), .Z(\mult_44/ab[45][1] ) );
  AND U462 ( .A(a[45]), .B(b[0]), .Z(\mult_44/ab[45][0] ) );
  AND U463 ( .A(b[3]), .B(a[44]), .Z(\mult_44/ab[44][3] ) );
  AND U464 ( .A(b[2]), .B(a[44]), .Z(\mult_44/ab[44][2] ) );
  AND U465 ( .A(b[1]), .B(a[44]), .Z(\mult_44/ab[44][1] ) );
  AND U466 ( .A(a[44]), .B(b[0]), .Z(\mult_44/ab[44][0] ) );
  AND U467 ( .A(b[3]), .B(a[43]), .Z(\mult_44/ab[43][3] ) );
  AND U468 ( .A(b[2]), .B(a[43]), .Z(\mult_44/ab[43][2] ) );
  AND U469 ( .A(b[1]), .B(a[43]), .Z(\mult_44/ab[43][1] ) );
  AND U470 ( .A(a[43]), .B(b[0]), .Z(\mult_44/ab[43][0] ) );
  AND U471 ( .A(b[3]), .B(a[42]), .Z(\mult_44/ab[42][3] ) );
  AND U472 ( .A(b[2]), .B(a[42]), .Z(\mult_44/ab[42][2] ) );
  AND U473 ( .A(b[1]), .B(a[42]), .Z(\mult_44/ab[42][1] ) );
  AND U474 ( .A(a[42]), .B(b[0]), .Z(\mult_44/ab[42][0] ) );
  AND U475 ( .A(b[3]), .B(a[41]), .Z(\mult_44/ab[41][3] ) );
  AND U476 ( .A(b[2]), .B(a[41]), .Z(\mult_44/ab[41][2] ) );
  AND U477 ( .A(b[1]), .B(a[41]), .Z(\mult_44/ab[41][1] ) );
  AND U478 ( .A(a[41]), .B(b[0]), .Z(\mult_44/ab[41][0] ) );
  AND U479 ( .A(b[3]), .B(a[40]), .Z(\mult_44/ab[40][3] ) );
  AND U480 ( .A(b[2]), .B(a[40]), .Z(\mult_44/ab[40][2] ) );
  AND U481 ( .A(b[1]), .B(a[40]), .Z(\mult_44/ab[40][1] ) );
  AND U482 ( .A(a[40]), .B(b[0]), .Z(\mult_44/ab[40][0] ) );
  AND U483 ( .A(b[3]), .B(a[3]), .Z(\mult_44/ab[3][3] ) );
  AND U484 ( .A(b[2]), .B(a[3]), .Z(\mult_44/ab[3][2] ) );
  AND U485 ( .A(b[1]), .B(a[3]), .Z(\mult_44/ab[3][1] ) );
  AND U486 ( .A(a[3]), .B(b[0]), .Z(\mult_44/ab[3][0] ) );
  AND U487 ( .A(b[3]), .B(a[39]), .Z(\mult_44/ab[39][3] ) );
  AND U488 ( .A(b[2]), .B(a[39]), .Z(\mult_44/ab[39][2] ) );
  AND U489 ( .A(b[1]), .B(a[39]), .Z(\mult_44/ab[39][1] ) );
  AND U490 ( .A(a[39]), .B(b[0]), .Z(\mult_44/ab[39][0] ) );
  AND U491 ( .A(b[3]), .B(a[38]), .Z(\mult_44/ab[38][3] ) );
  AND U492 ( .A(b[2]), .B(a[38]), .Z(\mult_44/ab[38][2] ) );
  AND U493 ( .A(b[1]), .B(a[38]), .Z(\mult_44/ab[38][1] ) );
  AND U494 ( .A(a[38]), .B(b[0]), .Z(\mult_44/ab[38][0] ) );
  AND U495 ( .A(b[3]), .B(a[37]), .Z(\mult_44/ab[37][3] ) );
  AND U496 ( .A(b[2]), .B(a[37]), .Z(\mult_44/ab[37][2] ) );
  AND U497 ( .A(b[1]), .B(a[37]), .Z(\mult_44/ab[37][1] ) );
  AND U498 ( .A(a[37]), .B(b[0]), .Z(\mult_44/ab[37][0] ) );
  AND U499 ( .A(b[3]), .B(a[36]), .Z(\mult_44/ab[36][3] ) );
  AND U500 ( .A(b[2]), .B(a[36]), .Z(\mult_44/ab[36][2] ) );
  AND U501 ( .A(b[1]), .B(a[36]), .Z(\mult_44/ab[36][1] ) );
  AND U502 ( .A(a[36]), .B(b[0]), .Z(\mult_44/ab[36][0] ) );
  AND U503 ( .A(b[3]), .B(a[35]), .Z(\mult_44/ab[35][3] ) );
  AND U504 ( .A(b[2]), .B(a[35]), .Z(\mult_44/ab[35][2] ) );
  AND U505 ( .A(b[1]), .B(a[35]), .Z(\mult_44/ab[35][1] ) );
  AND U506 ( .A(a[35]), .B(b[0]), .Z(\mult_44/ab[35][0] ) );
  AND U507 ( .A(b[3]), .B(a[34]), .Z(\mult_44/ab[34][3] ) );
  AND U508 ( .A(b[2]), .B(a[34]), .Z(\mult_44/ab[34][2] ) );
  AND U509 ( .A(b[1]), .B(a[34]), .Z(\mult_44/ab[34][1] ) );
  AND U510 ( .A(a[34]), .B(b[0]), .Z(\mult_44/ab[34][0] ) );
  AND U511 ( .A(b[3]), .B(a[33]), .Z(\mult_44/ab[33][3] ) );
  AND U512 ( .A(b[2]), .B(a[33]), .Z(\mult_44/ab[33][2] ) );
  AND U513 ( .A(b[1]), .B(a[33]), .Z(\mult_44/ab[33][1] ) );
  AND U514 ( .A(a[33]), .B(b[0]), .Z(\mult_44/ab[33][0] ) );
  AND U515 ( .A(b[3]), .B(a[32]), .Z(\mult_44/ab[32][3] ) );
  AND U516 ( .A(b[2]), .B(a[32]), .Z(\mult_44/ab[32][2] ) );
  AND U517 ( .A(b[1]), .B(a[32]), .Z(\mult_44/ab[32][1] ) );
  AND U518 ( .A(a[32]), .B(b[0]), .Z(\mult_44/ab[32][0] ) );
  AND U519 ( .A(b[3]), .B(a[31]), .Z(\mult_44/ab[31][3] ) );
  AND U520 ( .A(b[2]), .B(a[31]), .Z(\mult_44/ab[31][2] ) );
  AND U521 ( .A(b[1]), .B(a[31]), .Z(\mult_44/ab[31][1] ) );
  AND U522 ( .A(a[31]), .B(b[0]), .Z(\mult_44/ab[31][0] ) );
  AND U523 ( .A(b[3]), .B(a[30]), .Z(\mult_44/ab[30][3] ) );
  AND U524 ( .A(b[2]), .B(a[30]), .Z(\mult_44/ab[30][2] ) );
  AND U525 ( .A(b[1]), .B(a[30]), .Z(\mult_44/ab[30][1] ) );
  AND U526 ( .A(a[30]), .B(b[0]), .Z(\mult_44/ab[30][0] ) );
  AND U527 ( .A(b[3]), .B(a[2]), .Z(\mult_44/ab[2][3] ) );
  AND U528 ( .A(b[2]), .B(a[2]), .Z(\mult_44/ab[2][2] ) );
  AND U529 ( .A(b[1]), .B(a[2]), .Z(\mult_44/ab[2][1] ) );
  AND U530 ( .A(a[2]), .B(b[0]), .Z(\mult_44/ab[2][0] ) );
  AND U531 ( .A(b[3]), .B(a[29]), .Z(\mult_44/ab[29][3] ) );
  AND U532 ( .A(b[2]), .B(a[29]), .Z(\mult_44/ab[29][2] ) );
  AND U533 ( .A(b[1]), .B(a[29]), .Z(\mult_44/ab[29][1] ) );
  AND U534 ( .A(a[29]), .B(b[0]), .Z(\mult_44/ab[29][0] ) );
  AND U535 ( .A(b[3]), .B(a[28]), .Z(\mult_44/ab[28][3] ) );
  AND U536 ( .A(b[2]), .B(a[28]), .Z(\mult_44/ab[28][2] ) );
  AND U537 ( .A(b[1]), .B(a[28]), .Z(\mult_44/ab[28][1] ) );
  AND U538 ( .A(a[28]), .B(b[0]), .Z(\mult_44/ab[28][0] ) );
  AND U539 ( .A(b[3]), .B(a[27]), .Z(\mult_44/ab[27][3] ) );
  AND U540 ( .A(b[2]), .B(a[27]), .Z(\mult_44/ab[27][2] ) );
  AND U541 ( .A(b[1]), .B(a[27]), .Z(\mult_44/ab[27][1] ) );
  AND U542 ( .A(a[27]), .B(b[0]), .Z(\mult_44/ab[27][0] ) );
  AND U543 ( .A(b[3]), .B(a[26]), .Z(\mult_44/ab[26][3] ) );
  AND U544 ( .A(b[2]), .B(a[26]), .Z(\mult_44/ab[26][2] ) );
  AND U545 ( .A(b[1]), .B(a[26]), .Z(\mult_44/ab[26][1] ) );
  AND U546 ( .A(a[26]), .B(b[0]), .Z(\mult_44/ab[26][0] ) );
  AND U547 ( .A(b[3]), .B(a[25]), .Z(\mult_44/ab[25][3] ) );
  AND U548 ( .A(b[2]), .B(a[25]), .Z(\mult_44/ab[25][2] ) );
  AND U549 ( .A(b[1]), .B(a[25]), .Z(\mult_44/ab[25][1] ) );
  AND U550 ( .A(a[25]), .B(b[0]), .Z(\mult_44/ab[25][0] ) );
  AND U551 ( .A(b[3]), .B(a[24]), .Z(\mult_44/ab[24][3] ) );
  AND U552 ( .A(b[2]), .B(a[24]), .Z(\mult_44/ab[24][2] ) );
  AND U553 ( .A(b[1]), .B(a[24]), .Z(\mult_44/ab[24][1] ) );
  AND U554 ( .A(a[24]), .B(b[0]), .Z(\mult_44/ab[24][0] ) );
  AND U555 ( .A(b[3]), .B(a[23]), .Z(\mult_44/ab[23][3] ) );
  AND U556 ( .A(b[2]), .B(a[23]), .Z(\mult_44/ab[23][2] ) );
  AND U557 ( .A(b[1]), .B(a[23]), .Z(\mult_44/ab[23][1] ) );
  AND U558 ( .A(a[23]), .B(b[0]), .Z(\mult_44/ab[23][0] ) );
  AND U559 ( .A(b[3]), .B(a[22]), .Z(\mult_44/ab[22][3] ) );
  AND U560 ( .A(b[2]), .B(a[22]), .Z(\mult_44/ab[22][2] ) );
  AND U561 ( .A(b[1]), .B(a[22]), .Z(\mult_44/ab[22][1] ) );
  AND U562 ( .A(a[22]), .B(b[0]), .Z(\mult_44/ab[22][0] ) );
  AND U563 ( .A(b[3]), .B(a[21]), .Z(\mult_44/ab[21][3] ) );
  AND U564 ( .A(b[2]), .B(a[21]), .Z(\mult_44/ab[21][2] ) );
  AND U565 ( .A(b[1]), .B(a[21]), .Z(\mult_44/ab[21][1] ) );
  AND U566 ( .A(a[21]), .B(b[0]), .Z(\mult_44/ab[21][0] ) );
  AND U567 ( .A(b[3]), .B(a[20]), .Z(\mult_44/ab[20][3] ) );
  AND U568 ( .A(b[2]), .B(a[20]), .Z(\mult_44/ab[20][2] ) );
  AND U569 ( .A(b[1]), .B(a[20]), .Z(\mult_44/ab[20][1] ) );
  AND U570 ( .A(a[20]), .B(b[0]), .Z(\mult_44/ab[20][0] ) );
  AND U571 ( .A(b[3]), .B(a[1]), .Z(\mult_44/ab[1][3] ) );
  AND U572 ( .A(b[2]), .B(a[1]), .Z(\mult_44/ab[1][2] ) );
  AND U573 ( .A(b[1]), .B(a[1]), .Z(\mult_44/ab[1][1] ) );
  AND U574 ( .A(a[1]), .B(b[0]), .Z(\mult_44/ab[1][0] ) );
  AND U575 ( .A(b[3]), .B(a[19]), .Z(\mult_44/ab[19][3] ) );
  AND U576 ( .A(b[2]), .B(a[19]), .Z(\mult_44/ab[19][2] ) );
  AND U577 ( .A(b[1]), .B(a[19]), .Z(\mult_44/ab[19][1] ) );
  AND U578 ( .A(a[19]), .B(b[0]), .Z(\mult_44/ab[19][0] ) );
  AND U579 ( .A(b[3]), .B(a[18]), .Z(\mult_44/ab[18][3] ) );
  AND U580 ( .A(b[2]), .B(a[18]), .Z(\mult_44/ab[18][2] ) );
  AND U581 ( .A(b[1]), .B(a[18]), .Z(\mult_44/ab[18][1] ) );
  AND U582 ( .A(a[18]), .B(b[0]), .Z(\mult_44/ab[18][0] ) );
  AND U583 ( .A(b[3]), .B(a[17]), .Z(\mult_44/ab[17][3] ) );
  AND U584 ( .A(b[2]), .B(a[17]), .Z(\mult_44/ab[17][2] ) );
  AND U585 ( .A(b[1]), .B(a[17]), .Z(\mult_44/ab[17][1] ) );
  AND U586 ( .A(a[17]), .B(b[0]), .Z(\mult_44/ab[17][0] ) );
  AND U587 ( .A(b[3]), .B(a[16]), .Z(\mult_44/ab[16][3] ) );
  AND U588 ( .A(b[2]), .B(a[16]), .Z(\mult_44/ab[16][2] ) );
  AND U589 ( .A(b[1]), .B(a[16]), .Z(\mult_44/ab[16][1] ) );
  AND U590 ( .A(a[16]), .B(b[0]), .Z(\mult_44/ab[16][0] ) );
  AND U591 ( .A(b[3]), .B(a[15]), .Z(\mult_44/ab[15][3] ) );
  AND U592 ( .A(b[2]), .B(a[15]), .Z(\mult_44/ab[15][2] ) );
  AND U593 ( .A(b[1]), .B(a[15]), .Z(\mult_44/ab[15][1] ) );
  AND U594 ( .A(a[15]), .B(b[0]), .Z(\mult_44/ab[15][0] ) );
  AND U595 ( .A(b[3]), .B(a[14]), .Z(\mult_44/ab[14][3] ) );
  AND U596 ( .A(b[2]), .B(a[14]), .Z(\mult_44/ab[14][2] ) );
  AND U597 ( .A(b[1]), .B(a[14]), .Z(\mult_44/ab[14][1] ) );
  AND U598 ( .A(a[14]), .B(b[0]), .Z(\mult_44/ab[14][0] ) );
  AND U599 ( .A(b[3]), .B(a[13]), .Z(\mult_44/ab[13][3] ) );
  AND U600 ( .A(b[2]), .B(a[13]), .Z(\mult_44/ab[13][2] ) );
  AND U601 ( .A(b[1]), .B(a[13]), .Z(\mult_44/ab[13][1] ) );
  AND U602 ( .A(a[13]), .B(b[0]), .Z(\mult_44/ab[13][0] ) );
  AND U603 ( .A(b[3]), .B(a[12]), .Z(\mult_44/ab[12][3] ) );
  AND U604 ( .A(b[2]), .B(a[12]), .Z(\mult_44/ab[12][2] ) );
  AND U605 ( .A(b[1]), .B(a[12]), .Z(\mult_44/ab[12][1] ) );
  AND U606 ( .A(a[12]), .B(b[0]), .Z(\mult_44/ab[12][0] ) );
  AND U607 ( .A(b[3]), .B(a[11]), .Z(\mult_44/ab[11][3] ) );
  AND U608 ( .A(b[2]), .B(a[11]), .Z(\mult_44/ab[11][2] ) );
  AND U609 ( .A(b[1]), .B(a[11]), .Z(\mult_44/ab[11][1] ) );
  AND U610 ( .A(a[11]), .B(b[0]), .Z(\mult_44/ab[11][0] ) );
  AND U611 ( .A(b[3]), .B(a[10]), .Z(\mult_44/ab[10][3] ) );
  AND U612 ( .A(b[2]), .B(a[10]), .Z(\mult_44/ab[10][2] ) );
  AND U613 ( .A(b[1]), .B(a[10]), .Z(\mult_44/ab[10][1] ) );
  AND U614 ( .A(a[10]), .B(b[0]), .Z(\mult_44/ab[10][0] ) );
  AND U615 ( .A(a[0]), .B(b[3]), .Z(\mult_44/ab[0][3] ) );
  AND U616 ( .A(a[0]), .B(b[2]), .Z(\mult_44/ab[0][2] ) );
  AND U617 ( .A(a[0]), .B(b[1]), .Z(\mult_44/ab[0][1] ) );
  XNOR U618 ( .A(\mult_44/PROD1[3] ), .B(n296), .Z(c[63]) );
  XOR U619 ( .A(n297), .B(n298), .Z(n295) );
  ANDN U620 ( .B(n299), .A(n300), .Z(n298) );
  XOR U621 ( .A(clocal[2]), .B(n297), .Z(n299) );
  XNOR U622 ( .A(clocal[2]), .B(n300), .Z(c[62]) );
  XNOR U623 ( .A(n301), .B(n302), .Z(n297) );
  NANDN U624 ( .A(n303), .B(n304), .Z(n301) );
  XOR U625 ( .A(clocal[1]), .B(n302), .Z(n304) );
  XNOR U626 ( .A(clocal[1]), .B(n303), .Z(c[61]) );
  XNOR U627 ( .A(n302), .B(sreg[65]), .Z(n303) );
  ANDN U628 ( .B(sreg[64]), .A(n305), .Z(n302) );
  XNOR U629 ( .A(sreg[64]), .B(n305), .Z(c[60]) );
  NAND U630 ( .A(b[0]), .B(a[0]), .Z(n305) );
endmodule

