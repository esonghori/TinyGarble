
module modexp_1_N_N4_CC4 ( clk, rst, m, e, n, c );
  input [3:0] m;
  input [3:0] e;
  input [3:0] n;
  output [3:0] c;
  input clk, rst;
  wire   \cin[0][2] , \cin[0][1] , init, \keep_1[0] , N8, N9, N10, N11,
         \MODMULT1[0].modmult_1/MODMULT_STEP[0].modmult_step_/z2[3] ,
         \MODMULT1[0].modmult_1/MODMULT_STEP[1].modmult_step_/N4 ,
         \MODMULT2[0].modmult_2/MODMULT_STEP[1].modmult_step_/N4 , n3, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912;
  wire   [3:0] ein;
  wire   [3:0] ereg;
  assign \MODMULT2[0].modmult_2/MODMULT_STEP[1].modmult_step_/N4  = m[0];

  DFF init_reg ( .D(1'b1), .CLK(clk), .RST(rst), .Q(init) );
  DFF \ereg_reg[1]  ( .D(ein[0]), .CLK(clk), .RST(rst), .Q(ereg[1]) );
  DFF \ereg_reg[2]  ( .D(ein[1]), .CLK(clk), .RST(rst), .Q(ereg[2]) );
  DFF \ereg_reg[3]  ( .D(ein[2]), .CLK(clk), .RST(rst), .Q(ereg[3]) );
  DFF \creg_reg[1]  ( .D(N9), .CLK(clk), .RST(rst), .Q(\cin[0][1] ) );
  DFF \creg_reg[0]  ( .D(N8), .CLK(clk), .RST(rst), .Q(
        \MODMULT1[0].modmult_1/MODMULT_STEP[1].modmult_step_/N4 ) );
  DFF \creg_reg[3]  ( .D(N11), .CLK(clk), .RST(rst), .Q(
        \MODMULT1[0].modmult_1/MODMULT_STEP[0].modmult_step_/z2[3] ) );
  DFF \creg_reg[2]  ( .D(N10), .CLK(clk), .RST(rst), .Q(\cin[0][2] ) );
  DFF first_one_reg ( .D(n3), .CLK(clk), .RST(rst), .Q(\keep_1[0] ) );
  XOR U289 ( .A(n636), .B(n633), .Z(n185) );
  NANDN U290 ( .A(n[1]), .B(n185), .Z(n186) );
  NAND U291 ( .A(n636), .B(n633), .Z(n187) );
  AND U292 ( .A(n186), .B(n187), .Z(n639) );
  NOR U293 ( .A(n[0]), .B(n631), .Z(n188) );
  NAND U294 ( .A(n188), .B(n636), .Z(n189) );
  XOR U295 ( .A(n188), .B(n636), .Z(n190) );
  NANDN U296 ( .A(n[1]), .B(n190), .Z(n191) );
  NAND U297 ( .A(n189), .B(n191), .Z(n192) );
  XOR U298 ( .A(n866), .B(n638), .Z(n193) );
  NAND U299 ( .A(n193), .B(n192), .Z(n194) );
  NAND U300 ( .A(n866), .B(n638), .Z(n195) );
  AND U301 ( .A(n194), .B(n195), .Z(n646) );
  ANDN U302 ( .B(n511), .A(n[1]), .Z(n503) );
  NANDN U303 ( .A(n832), .B(m[3]), .Z(n196) );
  XOR U304 ( .A(m[3]), .B(n819), .Z(n197) );
  NAND U305 ( .A(n829), .B(n197), .Z(n198) );
  NAND U306 ( .A(n196), .B(n198), .Z(n199) );
  ANDN U307 ( .B(n199), .A(n890), .Z(n841) );
  XOR U308 ( .A(n853), .B(n850), .Z(n200) );
  NANDN U309 ( .A(n[1]), .B(n200), .Z(n201) );
  NAND U310 ( .A(n853), .B(n850), .Z(n202) );
  AND U311 ( .A(n201), .B(n202), .Z(n855) );
  NOR U312 ( .A(n[0]), .B(n359), .Z(n203) );
  NAND U313 ( .A(n203), .B(n377), .Z(n204) );
  XOR U314 ( .A(n203), .B(n377), .Z(n205) );
  NANDN U315 ( .A(n[1]), .B(n205), .Z(n206) );
  NAND U316 ( .A(n204), .B(n206), .Z(n207) );
  XNOR U317 ( .A(n866), .B(n372), .Z(n208) );
  AND U318 ( .A(n207), .B(n208), .Z(n209) );
  NOR U319 ( .A(n209), .B(n880), .Z(n210) );
  OR U320 ( .A(n[2]), .B(n372), .Z(n211) );
  NAND U321 ( .A(n210), .B(n211), .Z(n212) );
  AND U322 ( .A(\MODMULT1[0].modmult_1/MODMULT_STEP[0].modmult_step_/z2[3] ), 
        .B(n212), .Z(n375) );
  NAND U323 ( .A(n[0]), .B(n649), .Z(n213) );
  NANDN U324 ( .A(n[1]), .B(n652), .Z(n214) );
  XNOR U325 ( .A(n[1]), .B(n652), .Z(n215) );
  NAND U326 ( .A(n215), .B(n213), .Z(n216) );
  NAND U327 ( .A(n214), .B(n216), .Z(n217) );
  XOR U328 ( .A(n866), .B(n664), .Z(n218) );
  NAND U329 ( .A(n218), .B(n217), .Z(n219) );
  NAND U330 ( .A(n866), .B(n664), .Z(n220) );
  AND U331 ( .A(n219), .B(n220), .Z(n221) );
  NANDN U332 ( .A(n646), .B(n[3]), .Z(n222) );
  NANDN U333 ( .A(n880), .B(n645), .Z(n223) );
  NANDN U334 ( .A(n645), .B(n222), .Z(n224) );
  AND U335 ( .A(n223), .B(n224), .Z(n225) );
  NAND U336 ( .A(n647), .B(n225), .Z(n226) );
  OR U337 ( .A(n880), .B(n679), .Z(n227) );
  NANDN U338 ( .A(n221), .B(n227), .Z(n228) );
  AND U339 ( .A(n226), .B(n228), .Z(n677) );
  XNOR U340 ( .A(m[3]), .B(n672), .Z(n229) );
  AND U341 ( .A(n688), .B(n229), .Z(n230) );
  XNOR U342 ( .A(n670), .B(n230), .Z(n725) );
  AND U343 ( .A(n[0]), .B(n529), .Z(n231) );
  XOR U344 ( .A(n[1]), .B(n535), .Z(n232) );
  NAND U345 ( .A(n232), .B(n231), .Z(n233) );
  NAND U346 ( .A(n[1]), .B(n535), .Z(n234) );
  AND U347 ( .A(n233), .B(n234), .Z(n235) );
  XNOR U348 ( .A(n[2]), .B(n548), .Z(n236) );
  NAND U349 ( .A(n236), .B(n235), .Z(n237) );
  NANDN U350 ( .A(n[2]), .B(n548), .Z(n238) );
  NAND U351 ( .A(n237), .B(n238), .Z(n239) );
  OR U352 ( .A(n564), .B(n522), .Z(n240) );
  NANDN U353 ( .A(n[3]), .B(n239), .Z(n241) );
  ANDN U354 ( .B(n241), .A(n240), .Z(n242) );
  XNOR U355 ( .A(n[3]), .B(n239), .Z(n243) );
  NAND U356 ( .A(n243), .B(n557), .Z(n244) );
  NAND U357 ( .A(n242), .B(n244), .Z(n554) );
  NAND U358 ( .A(n[1]), .B(n801), .Z(n245) );
  XOR U359 ( .A(n[1]), .B(n801), .Z(n246) );
  NANDN U360 ( .A(n797), .B(n246), .Z(n247) );
  NAND U361 ( .A(n245), .B(n247), .Z(n793) );
  NANDN U362 ( .A(n[1]), .B(n853), .Z(n248) );
  NANDN U363 ( .A(n854), .B(n866), .Z(n249) );
  AND U364 ( .A(n248), .B(n249), .Z(n250) );
  NANDN U365 ( .A(n854), .B(n865), .Z(n251) );
  NAND U366 ( .A(n833), .B(n251), .Z(n252) );
  NANDN U367 ( .A(n250), .B(n252), .Z(n253) );
  ANDN U368 ( .B(n253), .A(n860), .Z(n254) );
  NAND U369 ( .A(n880), .B(n865), .Z(n255) );
  AND U370 ( .A(n254), .B(n255), .Z(n256) );
  NANDN U371 ( .A(n859), .B(n256), .Z(n863) );
  XNOR U372 ( .A(n653), .B(n652), .Z(n654) );
  AND U373 ( .A(n[0]), .B(n380), .Z(n257) );
  NAND U374 ( .A(n257), .B(n[1]), .Z(n258) );
  XOR U375 ( .A(n257), .B(n[1]), .Z(n259) );
  NANDN U376 ( .A(n383), .B(n259), .Z(n260) );
  NAND U377 ( .A(n258), .B(n260), .Z(n261) );
  NANDN U378 ( .A(n880), .B(n407), .Z(n262) );
  NANDN U379 ( .A(n407), .B(n866), .Z(n263) );
  NANDN U380 ( .A(n410), .B(n263), .Z(n264) );
  NAND U381 ( .A(n262), .B(n264), .Z(n265) );
  NAND U382 ( .A(n866), .B(n410), .Z(n266) );
  NAND U383 ( .A(n261), .B(n266), .Z(n267) );
  NANDN U384 ( .A(n265), .B(n267), .Z(n406) );
  ANDN U385 ( .B(n427), .A(n[1]), .Z(n419) );
  NANDN U386 ( .A(n537), .B(n536), .Z(n268) );
  NANDN U387 ( .A(n535), .B(n534), .Z(n269) );
  NAND U388 ( .A(n268), .B(n269), .Z(n550) );
  XNOR U389 ( .A(n755), .B(n756), .Z(n786) );
  AND U390 ( .A(n[0]), .B(n805), .Z(n270) );
  XOR U391 ( .A(n[1]), .B(n814), .Z(n271) );
  NAND U392 ( .A(n271), .B(n270), .Z(n272) );
  NAND U393 ( .A(n[1]), .B(n814), .Z(n273) );
  AND U394 ( .A(n272), .B(n273), .Z(n274) );
  XNOR U395 ( .A(n866), .B(n810), .Z(n275) );
  NANDN U396 ( .A(n274), .B(n275), .Z(n276) );
  AND U397 ( .A(n808), .B(n276), .Z(n277) );
  OR U398 ( .A(n880), .B(n836), .Z(n278) );
  NAND U399 ( .A(n277), .B(n278), .Z(n279) );
  NAND U400 ( .A(n809), .B(n279), .Z(n826) );
  NAND U401 ( .A(n[0]), .B(n803), .Z(n280) );
  NANDN U402 ( .A(n[1]), .B(n613), .Z(n281) );
  XNOR U403 ( .A(n[1]), .B(n613), .Z(n282) );
  NAND U404 ( .A(n282), .B(n280), .Z(n283) );
  NAND U405 ( .A(n281), .B(n283), .Z(n284) );
  XNOR U406 ( .A(n617), .B(n866), .Z(n285) );
  NANDN U407 ( .A(n284), .B(n285), .Z(n286) );
  NANDN U408 ( .A(n866), .B(n617), .Z(n287) );
  AND U409 ( .A(n286), .B(n287), .Z(n288) );
  ANDN U410 ( .B(n597), .A(n880), .Z(n289) );
  NANDN U411 ( .A(n605), .B(n609), .Z(n290) );
  AND U412 ( .A(n289), .B(n290), .Z(n291) );
  XNOR U413 ( .A(n291), .B(n603), .Z(n292) );
  NANDN U414 ( .A(n604), .B(n292), .Z(n293) );
  NANDN U415 ( .A(n[3]), .B(n288), .Z(n294) );
  ANDN U416 ( .B(n294), .A(n293), .Z(n295) );
  XNOR U417 ( .A(n288), .B(n[3]), .Z(n296) );
  NAND U418 ( .A(n296), .B(n626), .Z(n297) );
  NAND U419 ( .A(n295), .B(n297), .Z(n622) );
  AND U420 ( .A(n[0]), .B(n892), .Z(n298) );
  XOR U421 ( .A(n[1]), .B(n902), .Z(n299) );
  NAND U422 ( .A(n299), .B(n298), .Z(n300) );
  NAND U423 ( .A(n[1]), .B(n902), .Z(n301) );
  AND U424 ( .A(n300), .B(n301), .Z(n302) );
  XNOR U425 ( .A(n875), .B(n866), .Z(n303) );
  NANDN U426 ( .A(n302), .B(n303), .Z(n304) );
  NANDN U427 ( .A(n866), .B(n875), .Z(n305) );
  AND U428 ( .A(n304), .B(n305), .Z(n306) );
  ANDN U429 ( .B(n863), .A(n880), .Z(n307) );
  NANDN U430 ( .A(n861), .B(n865), .Z(n308) );
  AND U431 ( .A(n307), .B(n308), .Z(n309) );
  XNOR U432 ( .A(n309), .B(n859), .Z(n310) );
  NANDN U433 ( .A(n860), .B(n310), .Z(n311) );
  NANDN U434 ( .A(n[3]), .B(n306), .Z(n312) );
  ANDN U435 ( .B(n312), .A(n311), .Z(n313) );
  XNOR U436 ( .A(n306), .B(n[3]), .Z(n314) );
  NAND U437 ( .A(n314), .B(n883), .Z(n315) );
  NAND U438 ( .A(n313), .B(n315), .Z(n879) );
  XNOR U439 ( .A(n655), .B(n654), .Z(n659) );
  ANDN U440 ( .B(n[0]), .A(n449), .Z(n316) );
  XOR U441 ( .A(n[1]), .B(n453), .Z(n317) );
  NAND U442 ( .A(n317), .B(n316), .Z(n318) );
  NAND U443 ( .A(n[1]), .B(n453), .Z(n319) );
  AND U444 ( .A(n318), .B(n319), .Z(n320) );
  XNOR U445 ( .A(n[2]), .B(n478), .Z(n321) );
  NAND U446 ( .A(n321), .B(n320), .Z(n322) );
  NANDN U447 ( .A(n[2]), .B(n478), .Z(n323) );
  NAND U448 ( .A(n322), .B(n323), .Z(n324) );
  NAND U449 ( .A(n442), .B(n441), .Z(n325) );
  NANDN U450 ( .A(n494), .B(n325), .Z(n326) );
  NANDN U451 ( .A(n[3]), .B(n324), .Z(n327) );
  ANDN U452 ( .B(n327), .A(n326), .Z(n328) );
  XNOR U453 ( .A(n[3]), .B(n324), .Z(n329) );
  NAND U454 ( .A(n329), .B(n488), .Z(n330) );
  NAND U455 ( .A(n328), .B(n330), .Z(n484) );
  ANDN U456 ( .B(n[0]), .A(n734), .Z(n331) );
  XOR U457 ( .A(n[1]), .B(n727), .Z(n332) );
  NAND U458 ( .A(n332), .B(n331), .Z(n333) );
  NAND U459 ( .A(n[1]), .B(n727), .Z(n334) );
  AND U460 ( .A(n333), .B(n334), .Z(n335) );
  XNOR U461 ( .A(n[2]), .B(n742), .Z(n336) );
  NAND U462 ( .A(n336), .B(n335), .Z(n337) );
  NANDN U463 ( .A(n[2]), .B(n742), .Z(n338) );
  NAND U464 ( .A(n337), .B(n338), .Z(n339) );
  NANDN U465 ( .A(n758), .B(n720), .Z(n340) );
  NANDN U466 ( .A(n[3]), .B(n339), .Z(n341) );
  ANDN U467 ( .B(n341), .A(n340), .Z(n342) );
  XNOR U468 ( .A(n[3]), .B(n339), .Z(n343) );
  NAND U469 ( .A(n343), .B(n752), .Z(n344) );
  NAND U470 ( .A(n342), .B(n344), .Z(n748) );
  XNOR U471 ( .A(n491), .B(n492), .Z(n521) );
  XNOR U472 ( .A(n556), .B(n555), .Z(n561) );
  NAND U473 ( .A(n820), .B(m[2]), .Z(n345) );
  XOR U474 ( .A(n820), .B(m[2]), .Z(n346) );
  NAND U475 ( .A(n346), .B(n821), .Z(n347) );
  NAND U476 ( .A(n345), .B(n347), .Z(n829) );
  NANDN U477 ( .A(n[3]), .B(n785), .Z(n348) );
  ANDN U478 ( .B(n348), .A(n799), .Z(n349) );
  NAND U479 ( .A(n788), .B(n790), .Z(n350) );
  NAND U480 ( .A(n349), .B(n350), .Z(n351) );
  XNOR U481 ( .A(n786), .B(n351), .Z(n843) );
  NAND U482 ( .A(n612), .B(n613), .Z(n352) );
  XOR U483 ( .A(n612), .B(n613), .Z(n353) );
  NANDN U484 ( .A(n615), .B(n353), .Z(n354) );
  NAND U485 ( .A(n352), .B(n354), .Z(n616) );
  XOR U486 ( .A(n902), .B(n900), .Z(n355) );
  NAND U487 ( .A(n355), .B(n899), .Z(n356) );
  NAND U488 ( .A(n902), .B(n900), .Z(n357) );
  AND U489 ( .A(n356), .B(n357), .Z(n876) );
  NAND U490 ( .A(\MODMULT1[0].modmult_1/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(\cin[0][1] ), .Z(n585) );
  IV U491 ( .A(n585), .Z(n501) );
  NAND U492 ( .A(\MODMULT1[0].modmult_1/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(\MODMULT1[0].modmult_1/MODMULT_STEP[0].modmult_step_/z2[3] ), .Z(
        n359) );
  NAND U493 ( .A(\MODMULT1[0].modmult_1/MODMULT_STEP[0].modmult_step_/z2[3] ), 
        .B(\cin[0][2] ), .Z(n372) );
  IV U494 ( .A(n[3]), .Z(n880) );
  AND U495 ( .A(\MODMULT1[0].modmult_1/MODMULT_STEP[0].modmult_step_/z2[3] ), 
        .B(\cin[0][1] ), .Z(n377) );
  IV U496 ( .A(n[2]), .Z(n866) );
  NAND U497 ( .A(n375), .B(n[0]), .Z(n358) );
  XNOR U498 ( .A(n359), .B(n358), .Z(n380) );
  AND U499 ( .A(n[0]), .B(n359), .Z(n361) );
  IV U500 ( .A(n361), .Z(n373) );
  ANDN U501 ( .B(n[1]), .A(n373), .Z(n360) );
  NANDN U502 ( .A(n360), .B(n377), .Z(n363) );
  NOR U503 ( .A(n361), .B(n[1]), .Z(n362) );
  ANDN U504 ( .B(n363), .A(n362), .Z(n364) );
  NANDN U505 ( .A(n866), .B(n364), .Z(n366) );
  XNOR U506 ( .A(n866), .B(n364), .Z(n370) );
  NAND U507 ( .A(n372), .B(n370), .Z(n365) );
  NAND U508 ( .A(n366), .B(n365), .Z(n367) );
  NANDN U509 ( .A(n367), .B(n880), .Z(n368) );
  NAND U510 ( .A(n375), .B(n368), .Z(n369) );
  NAND U511 ( .A(\MODMULT1[0].modmult_1/MODMULT_STEP[0].modmult_step_/z2[3] ), 
        .B(n369), .Z(n407) );
  NAND U512 ( .A(n375), .B(n370), .Z(n371) );
  XOR U513 ( .A(n372), .B(n371), .Z(n410) );
  XNOR U514 ( .A(n[1]), .B(n373), .Z(n374) );
  NAND U515 ( .A(n375), .B(n374), .Z(n376) );
  XNOR U516 ( .A(n377), .B(n376), .Z(n383) );
  NANDN U517 ( .A(n407), .B(n880), .Z(n378) );
  AND U518 ( .A(n406), .B(n378), .Z(n382) );
  ANDN U519 ( .B(n[0]), .A(n382), .Z(n379) );
  AND U520 ( .A(n380), .B(n379), .Z(n386) );
  ANDN U521 ( .B(n[1]), .A(n382), .Z(n384) );
  XNOR U522 ( .A(n383), .B(n384), .Z(n385) );
  XNOR U523 ( .A(n386), .B(n385), .Z(n389) );
  XOR U524 ( .A(n380), .B(n379), .Z(n396) );
  NANDN U525 ( .A(n396), .B(\cin[0][1] ), .Z(n390) );
  NAND U526 ( .A(n390), .B(\cin[0][2] ), .Z(n381) );
  XOR U527 ( .A(n389), .B(n381), .Z(n432) );
  NOR U528 ( .A(n866), .B(n382), .Z(n409) );
  XNOR U529 ( .A(n410), .B(n409), .Z(n412) );
  NANDN U530 ( .A(n384), .B(n383), .Z(n388) );
  NANDN U531 ( .A(n386), .B(n385), .Z(n387) );
  NAND U532 ( .A(n388), .B(n387), .Z(n411) );
  XOR U533 ( .A(n412), .B(n411), .Z(n404) );
  OR U534 ( .A(n404), .B(\cin[0][2] ), .Z(n394) );
  ANDN U535 ( .B(n390), .A(n389), .Z(n403) );
  NANDN U536 ( .A(n404), .B(
        \MODMULT1[0].modmult_1/MODMULT_STEP[0].modmult_step_/z2[3] ), .Z(n391)
         );
  XNOR U537 ( .A(n403), .B(n391), .Z(n392) );
  NAND U538 ( .A(\cin[0][2] ), .B(n392), .Z(n393) );
  NAND U539 ( .A(n394), .B(n393), .Z(n447) );
  NANDN U540 ( .A(n880), .B(n447), .Z(n435) );
  NAND U541 ( .A(\cin[0][2] ), .B(\cin[0][1] ), .Z(n395) );
  XOR U542 ( .A(n396), .B(n395), .Z(n427) );
  NANDN U543 ( .A(n427), .B(n[1]), .Z(n421) );
  NAND U544 ( .A(\MODMULT1[0].modmult_1/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(\cin[0][2] ), .Z(n429) );
  NOR U545 ( .A(n429), .B(n[0]), .Z(n397) );
  NAND U546 ( .A(n421), .B(n397), .Z(n398) );
  NANDN U547 ( .A(n419), .B(n398), .Z(n399) );
  OR U548 ( .A(n399), .B(n866), .Z(n400) );
  AND U549 ( .A(n435), .B(n400), .Z(n401) );
  NANDN U550 ( .A(n432), .B(n401), .Z(n402) );
  ANDN U551 ( .B(n880), .A(n447), .Z(n438) );
  ANDN U552 ( .B(n402), .A(n438), .Z(n418) );
  NANDN U553 ( .A(n404), .B(n403), .Z(n405) );
  AND U554 ( .A(\cin[0][2] ), .B(n405), .Z(n442) );
  OR U555 ( .A(n406), .B(n880), .Z(n408) );
  ANDN U556 ( .B(n408), .A(n407), .Z(n416) );
  ANDN U557 ( .B(n410), .A(n409), .Z(n414) );
  AND U558 ( .A(n412), .B(n411), .Z(n413) );
  NOR U559 ( .A(n414), .B(n413), .Z(n415) );
  XOR U560 ( .A(n416), .B(n415), .Z(n441) );
  OR U561 ( .A(n442), .B(n441), .Z(n417) );
  ANDN U562 ( .B(n418), .A(n417), .Z(n444) );
  AND U563 ( .A(n[0]), .B(n429), .Z(n424) );
  NANDN U564 ( .A(n419), .B(n424), .Z(n420) );
  NAND U565 ( .A(n421), .B(n420), .Z(n430) );
  XOR U566 ( .A(n[2]), .B(n430), .Z(n422) );
  NANDN U567 ( .A(n444), .B(n422), .Z(n423) );
  XOR U568 ( .A(n432), .B(n423), .Z(n478) );
  XOR U569 ( .A(n[1]), .B(n424), .Z(n425) );
  NANDN U570 ( .A(n444), .B(n425), .Z(n426) );
  XOR U571 ( .A(n427), .B(n426), .Z(n453) );
  NANDN U572 ( .A(n444), .B(n[0]), .Z(n428) );
  XOR U573 ( .A(n429), .B(n428), .Z(n449) );
  XNOR U574 ( .A(n866), .B(n432), .Z(n431) );
  NAND U575 ( .A(n431), .B(n430), .Z(n434) );
  NANDN U576 ( .A(n866), .B(n432), .Z(n433) );
  AND U577 ( .A(n434), .B(n433), .Z(n443) );
  NAND U578 ( .A(n443), .B(n435), .Z(n436) );
  ANDN U579 ( .B(n436), .A(n444), .Z(n437) );
  NANDN U580 ( .A(n438), .B(n437), .Z(n440) );
  XNOR U581 ( .A(n442), .B(n441), .Z(n439) );
  XOR U582 ( .A(n440), .B(n439), .Z(n494) );
  XOR U583 ( .A(n443), .B(n880), .Z(n445) );
  ANDN U584 ( .B(n445), .A(n444), .Z(n446) );
  XNOR U585 ( .A(n447), .B(n446), .Z(n488) );
  AND U586 ( .A(n[0]), .B(n484), .Z(n448) );
  ANDN U587 ( .B(n448), .A(n449), .Z(n455) );
  NAND U588 ( .A(n[1]), .B(n484), .Z(n452) );
  XNOR U589 ( .A(n453), .B(n452), .Z(n454) );
  XNOR U590 ( .A(n455), .B(n454), .Z(n459) );
  IV U591 ( .A(n459), .Z(n458) );
  XOR U592 ( .A(n449), .B(n448), .Z(n465) );
  XOR U593 ( .A(\cin[0][2] ), .B(n465), .Z(n450) );
  NAND U594 ( .A(\cin[0][1] ), .B(n450), .Z(n451) );
  XOR U595 ( .A(n458), .B(n451), .Z(n507) );
  OR U596 ( .A(n507), .B(n866), .Z(n516) );
  ANDN U597 ( .B(n484), .A(n866), .Z(n479) );
  XNOR U598 ( .A(n478), .B(n479), .Z(n481) );
  NANDN U599 ( .A(n453), .B(n452), .Z(n457) );
  NANDN U600 ( .A(n455), .B(n454), .Z(n456) );
  NAND U601 ( .A(n457), .B(n456), .Z(n480) );
  XOR U602 ( .A(n481), .B(n480), .Z(n472) );
  IV U603 ( .A(n472), .Z(n471) );
  NANDN U604 ( .A(n458), .B(\cin[0][2] ), .Z(n462) );
  XOR U605 ( .A(\cin[0][2] ), .B(n459), .Z(n460) );
  NAND U606 ( .A(n460), .B(n465), .Z(n461) );
  NAND U607 ( .A(n462), .B(n461), .Z(n473) );
  XOR U608 ( .A(\MODMULT1[0].modmult_1/MODMULT_STEP[0].modmult_step_/z2[3] ), 
        .B(n473), .Z(n463) );
  NAND U609 ( .A(\cin[0][1] ), .B(n463), .Z(n464) );
  XOR U610 ( .A(n471), .B(n464), .Z(n527) );
  NOR U611 ( .A(n880), .B(n527), .Z(n517) );
  ANDN U612 ( .B(n516), .A(n517), .Z(n470) );
  XOR U613 ( .A(\cin[0][1] ), .B(n465), .Z(n511) );
  ANDN U614 ( .B(n[1]), .A(n511), .Z(n502) );
  NOR U615 ( .A(n585), .B(n[0]), .Z(n466) );
  NANDN U616 ( .A(n502), .B(n466), .Z(n467) );
  NANDN U617 ( .A(n503), .B(n467), .Z(n468) );
  AND U618 ( .A(n507), .B(n866), .Z(n514) );
  OR U619 ( .A(n468), .B(n514), .Z(n469) );
  AND U620 ( .A(n470), .B(n469), .Z(n499) );
  AND U621 ( .A(n527), .B(n880), .Z(n512) );
  ANDN U622 ( .B(\MODMULT1[0].modmult_1/MODMULT_STEP[0].modmult_step_/z2[3] ), 
        .A(n471), .Z(n476) );
  XOR U623 ( .A(\MODMULT1[0].modmult_1/MODMULT_STEP[0].modmult_step_/z2[3] ), 
        .B(n472), .Z(n474) );
  AND U624 ( .A(n474), .B(n473), .Z(n475) );
  OR U625 ( .A(n476), .B(n475), .Z(n477) );
  AND U626 ( .A(\cin[0][1] ), .B(n477), .Z(n492) );
  NANDN U627 ( .A(n479), .B(n478), .Z(n483) );
  NAND U628 ( .A(n481), .B(n480), .Z(n482) );
  NAND U629 ( .A(n483), .B(n482), .Z(n485) );
  NANDN U630 ( .A(n880), .B(n484), .Z(n487) );
  XOR U631 ( .A(n488), .B(n487), .Z(n486) );
  XNOR U632 ( .A(n485), .B(n486), .Z(n491) );
  NOR U633 ( .A(n512), .B(n521), .Z(n497) );
  NAND U634 ( .A(n486), .B(n485), .Z(n490) );
  NAND U635 ( .A(n488), .B(n487), .Z(n489) );
  AND U636 ( .A(n490), .B(n489), .Z(n496) );
  ANDN U637 ( .B(n492), .A(n491), .Z(n493) );
  XNOR U638 ( .A(n494), .B(n493), .Z(n495) );
  XNOR U639 ( .A(n496), .B(n495), .Z(n522) );
  ANDN U640 ( .B(n497), .A(n522), .Z(n498) );
  NANDN U641 ( .A(n499), .B(n498), .Z(n525) );
  NAND U642 ( .A(n525), .B(n[0]), .Z(n500) );
  XOR U643 ( .A(n501), .B(n500), .Z(n529) );
  ANDN U644 ( .B(n[0]), .A(n501), .Z(n508) );
  OR U645 ( .A(n502), .B(n508), .Z(n504) );
  ANDN U646 ( .B(n504), .A(n503), .Z(n513) );
  XNOR U647 ( .A(n866), .B(n513), .Z(n505) );
  NAND U648 ( .A(n525), .B(n505), .Z(n506) );
  XNOR U649 ( .A(n507), .B(n506), .Z(n548) );
  XOR U650 ( .A(n[1]), .B(n508), .Z(n509) );
  NAND U651 ( .A(n525), .B(n509), .Z(n510) );
  XOR U652 ( .A(n511), .B(n510), .Z(n535) );
  ANDN U653 ( .B(n525), .A(n512), .Z(n519) );
  NANDN U654 ( .A(n514), .B(n513), .Z(n515) );
  AND U655 ( .A(n516), .B(n515), .Z(n523) );
  NANDN U656 ( .A(n517), .B(n523), .Z(n518) );
  AND U657 ( .A(n519), .B(n518), .Z(n520) );
  XOR U658 ( .A(n521), .B(n520), .Z(n564) );
  XOR U659 ( .A(n880), .B(n523), .Z(n524) );
  NAND U660 ( .A(n525), .B(n524), .Z(n526) );
  XNOR U661 ( .A(n527), .B(n526), .Z(n557) );
  AND U662 ( .A(n[0]), .B(n554), .Z(n528) );
  NAND U663 ( .A(n529), .B(n528), .Z(n536) );
  NAND U664 ( .A(n[1]), .B(n554), .Z(n534) );
  XOR U665 ( .A(n535), .B(n534), .Z(n537) );
  XOR U666 ( .A(n536), .B(n537), .Z(n539) );
  XOR U667 ( .A(\cin[0][2] ), .B(n539), .Z(n540) );
  XOR U668 ( .A(n529), .B(n528), .Z(n586) );
  ANDN U669 ( .B(\cin[0][1] ), .A(n586), .Z(n530) );
  XNOR U670 ( .A(n540), .B(n530), .Z(n531) );
  NAND U671 ( .A(\MODMULT1[0].modmult_1/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(n531), .Z(n533) );
  OR U672 ( .A(\MODMULT1[0].modmult_1/MODMULT_STEP[1].modmult_step_/N4 ), .B(
        n539), .Z(n532) );
  AND U673 ( .A(n533), .B(n532), .Z(n598) );
  ANDN U674 ( .B(n554), .A(n866), .Z(n549) );
  XNOR U675 ( .A(n548), .B(n549), .Z(n551) );
  XOR U676 ( .A(n551), .B(n550), .Z(n538) );
  IV U677 ( .A(n538), .Z(n570) );
  ANDN U678 ( .B(\MODMULT1[0].modmult_1/MODMULT_STEP[0].modmult_step_/z2[3] ), 
        .A(n570), .Z(n546) );
  XOR U679 ( .A(\MODMULT1[0].modmult_1/MODMULT_STEP[0].modmult_step_/z2[3] ), 
        .B(n538), .Z(n544) );
  NANDN U680 ( .A(n539), .B(\cin[0][2] ), .Z(n543) );
  NANDN U681 ( .A(n586), .B(\cin[0][1] ), .Z(n541) );
  OR U682 ( .A(n541), .B(n540), .Z(n542) );
  AND U683 ( .A(n543), .B(n542), .Z(n567) );
  ANDN U684 ( .B(n544), .A(n567), .Z(n545) );
  OR U685 ( .A(n546), .B(n545), .Z(n547) );
  AND U686 ( .A(\MODMULT1[0].modmult_1/MODMULT_STEP[1].modmult_step_/N4 ), .B(
        n547), .Z(n562) );
  NANDN U687 ( .A(n549), .B(n548), .Z(n553) );
  NAND U688 ( .A(n551), .B(n550), .Z(n552) );
  AND U689 ( .A(n553), .B(n552), .Z(n556) );
  ANDN U690 ( .B(n554), .A(n880), .Z(n558) );
  XNOR U691 ( .A(n557), .B(n558), .Z(n555) );
  XOR U692 ( .A(n562), .B(n561), .Z(n603) );
  NANDN U693 ( .A(n556), .B(n555), .Z(n560) );
  NANDN U694 ( .A(n558), .B(n557), .Z(n559) );
  AND U695 ( .A(n560), .B(n559), .Z(n566) );
  AND U696 ( .A(n562), .B(n561), .Z(n563) );
  XNOR U697 ( .A(n564), .B(n563), .Z(n565) );
  XNOR U698 ( .A(n566), .B(n565), .Z(n604) );
  XNOR U699 ( .A(\MODMULT1[0].modmult_1/MODMULT_STEP[0].modmult_step_/z2[3] ), 
        .B(n567), .Z(n568) );
  NAND U700 ( .A(\MODMULT1[0].modmult_1/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(n568), .Z(n569) );
  XOR U701 ( .A(n570), .B(n569), .Z(n609) );
  NAND U702 ( .A(n866), .B(n609), .Z(n573) );
  OR U703 ( .A(n609), .B(n880), .Z(n571) );
  NANDN U704 ( .A(n598), .B(n571), .Z(n572) );
  NAND U705 ( .A(n573), .B(n572), .Z(n579) );
  XOR U706 ( .A(n585), .B(n586), .Z(n596) );
  NANDN U707 ( .A(n[0]), .B(
        \MODMULT1[0].modmult_1/MODMULT_STEP[1].modmult_step_/N4 ), .Z(n574) );
  NANDN U708 ( .A(n596), .B(n574), .Z(n575) );
  ANDN U709 ( .B(n575), .A(n[1]), .Z(n577) );
  ANDN U710 ( .B(n866), .A(n598), .Z(n576) );
  OR U711 ( .A(n577), .B(n576), .Z(n578) );
  NAND U712 ( .A(n579), .B(n578), .Z(n580) );
  NANDN U713 ( .A(n604), .B(n580), .Z(n581) );
  NOR U714 ( .A(n603), .B(n581), .Z(n583) );
  NAND U715 ( .A(n880), .B(n609), .Z(n582) );
  AND U716 ( .A(n583), .B(n582), .Z(n607) );
  ANDN U717 ( .B(n[0]), .A(
        \MODMULT1[0].modmult_1/MODMULT_STEP[1].modmult_step_/N4 ), .Z(n593) );
  OR U718 ( .A(n586), .B(n[1]), .Z(n584) );
  NAND U719 ( .A(n593), .B(n584), .Z(n589) );
  XNOR U720 ( .A(n586), .B(n585), .Z(n587) );
  NAND U721 ( .A(n[1]), .B(n587), .Z(n588) );
  AND U722 ( .A(n589), .B(n588), .Z(n600) );
  XOR U723 ( .A(n866), .B(n600), .Z(n590) );
  NANDN U724 ( .A(n607), .B(n590), .Z(n591) );
  XNOR U725 ( .A(n598), .B(n591), .Z(n617) );
  IV U726 ( .A(n607), .Z(n597) );
  AND U727 ( .A(n[0]), .B(n597), .Z(n592) );
  XNOR U728 ( .A(\MODMULT1[0].modmult_1/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(n592), .Z(n803) );
  XOR U729 ( .A(n[1]), .B(n593), .Z(n594) );
  ANDN U730 ( .B(n594), .A(n607), .Z(n595) );
  XOR U731 ( .A(n596), .B(n595), .Z(n613) );
  NANDN U732 ( .A(n866), .B(n598), .Z(n602) );
  XNOR U733 ( .A(n866), .B(n598), .Z(n599) );
  NANDN U734 ( .A(n600), .B(n599), .Z(n601) );
  NAND U735 ( .A(n602), .B(n601), .Z(n605) );
  XNOR U736 ( .A(n880), .B(n605), .Z(n606) );
  NANDN U737 ( .A(n607), .B(n606), .Z(n608) );
  XNOR U738 ( .A(n609), .B(n608), .Z(n626) );
  AND U739 ( .A(n[0]), .B(n622), .Z(n802) );
  NAND U740 ( .A(n803), .B(n802), .Z(n612) );
  AND U741 ( .A(n[1]), .B(n622), .Z(n615) );
  XNOR U742 ( .A(n617), .B(n616), .Z(n619) );
  ANDN U743 ( .B(n622), .A(n866), .Z(n618) );
  XNOR U744 ( .A(n619), .B(n618), .Z(n688) );
  NANDN U745 ( .A(ereg[3]), .B(init), .Z(n611) );
  OR U746 ( .A(init), .B(e[3]), .Z(n610) );
  NAND U747 ( .A(n611), .B(n610), .Z(n912) );
  NAND U748 ( .A(n688), .B(n912), .Z(n869) );
  XOR U749 ( .A(n613), .B(n612), .Z(n614) );
  XNOR U750 ( .A(n615), .B(n614), .Z(n898) );
  NAND U751 ( .A(n898), .B(
        \MODMULT2[0].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), .Z(n781) );
  ANDN U752 ( .B(n617), .A(n616), .Z(n621) );
  AND U753 ( .A(n619), .B(n618), .Z(n620) );
  NOR U754 ( .A(n621), .B(n620), .Z(n624) );
  ANDN U755 ( .B(n622), .A(n880), .Z(n623) );
  XNOR U756 ( .A(n624), .B(n623), .Z(n625) );
  XOR U757 ( .A(n626), .B(n625), .Z(n872) );
  NAND U758 ( .A(\MODMULT2[0].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(n872), .Z(n631) );
  AND U759 ( .A(m[3]), .B(n872), .Z(n647) );
  AND U760 ( .A(m[1]), .B(n872), .Z(n636) );
  AND U761 ( .A(m[2]), .B(n872), .Z(n638) );
  XNOR U762 ( .A(n880), .B(n646), .Z(n627) );
  NANDN U763 ( .A(n647), .B(n627), .Z(n629) );
  NANDN U764 ( .A(n880), .B(n646), .Z(n628) );
  NAND U765 ( .A(n629), .B(n628), .Z(n643) );
  NANDN U766 ( .A(n643), .B(n[0]), .Z(n630) );
  XNOR U767 ( .A(n631), .B(n630), .Z(n649) );
  NAND U768 ( .A(n[0]), .B(n631), .Z(n633) );
  XNOR U769 ( .A(n866), .B(n639), .Z(n637) );
  ANDN U770 ( .B(n637), .A(n643), .Z(n632) );
  XOR U771 ( .A(n638), .B(n632), .Z(n664) );
  XNOR U772 ( .A(n[1]), .B(n633), .Z(n634) );
  NANDN U773 ( .A(n643), .B(n634), .Z(n635) );
  XNOR U774 ( .A(n636), .B(n635), .Z(n652) );
  NANDN U775 ( .A(n638), .B(n637), .Z(n641) );
  NANDN U776 ( .A(n866), .B(n639), .Z(n640) );
  AND U777 ( .A(n641), .B(n640), .Z(n645) );
  XOR U778 ( .A(n880), .B(n645), .Z(n642) );
  NANDN U779 ( .A(n643), .B(n642), .Z(n644) );
  AND U780 ( .A(n647), .B(n644), .Z(n679) );
  ANDN U781 ( .B(n[0]), .A(n677), .Z(n648) );
  AND U782 ( .A(n649), .B(n648), .Z(n655) );
  ANDN U783 ( .B(n[1]), .A(n677), .Z(n653) );
  IV U784 ( .A(n659), .Z(n658) );
  XNOR U785 ( .A(n649), .B(n648), .Z(n687) );
  AND U786 ( .A(m[1]), .B(n687), .Z(n661) );
  XOR U787 ( .A(m[2]), .B(n661), .Z(n650) );
  NAND U788 ( .A(n688), .B(n650), .Z(n651) );
  XOR U789 ( .A(n658), .B(n651), .Z(n703) );
  NOR U790 ( .A(n866), .B(n677), .Z(n665) );
  XNOR U791 ( .A(n664), .B(n665), .Z(n667) );
  NANDN U792 ( .A(n653), .B(n652), .Z(n657) );
  NANDN U793 ( .A(n655), .B(n654), .Z(n656) );
  NAND U794 ( .A(n657), .B(n656), .Z(n666) );
  XOR U795 ( .A(n667), .B(n666), .Z(n671) );
  IV U796 ( .A(n671), .Z(n670) );
  NANDN U797 ( .A(n658), .B(m[2]), .Z(n663) );
  XOR U798 ( .A(m[2]), .B(n659), .Z(n660) );
  NAND U799 ( .A(n661), .B(n660), .Z(n662) );
  AND U800 ( .A(n663), .B(n662), .Z(n672) );
  AND U801 ( .A(n725), .B(n880), .Z(n710) );
  NANDN U802 ( .A(n665), .B(n664), .Z(n669) );
  NAND U803 ( .A(n667), .B(n666), .Z(n668) );
  AND U804 ( .A(n669), .B(n668), .Z(n683) );
  ANDN U805 ( .B(m[3]), .A(n670), .Z(n675) );
  XOR U806 ( .A(m[3]), .B(n671), .Z(n673) );
  ANDN U807 ( .B(n673), .A(n672), .Z(n674) );
  OR U808 ( .A(n675), .B(n674), .Z(n676) );
  AND U809 ( .A(n688), .B(n676), .Z(n685) );
  XOR U810 ( .A(n683), .B(n685), .Z(n681) );
  OR U811 ( .A(n677), .B(n880), .Z(n678) );
  AND U812 ( .A(n679), .B(n678), .Z(n682) );
  XNOR U813 ( .A(n685), .B(n682), .Z(n680) );
  NAND U814 ( .A(n681), .B(n680), .Z(n720) );
  XNOR U815 ( .A(n683), .B(n682), .Z(n684) );
  XNOR U816 ( .A(n685), .B(n684), .Z(n719) );
  ANDN U817 ( .B(n720), .A(n719), .Z(n695) );
  OR U818 ( .A(n703), .B(n866), .Z(n714) );
  NOR U819 ( .A(n880), .B(n725), .Z(n715) );
  ANDN U820 ( .B(n714), .A(n715), .Z(n693) );
  NAND U821 ( .A(n688), .B(m[1]), .Z(n686) );
  XOR U822 ( .A(n687), .B(n686), .Z(n707) );
  NOR U823 ( .A(n707), .B(n[1]), .Z(n698) );
  NAND U824 ( .A(n[1]), .B(n707), .Z(n700) );
  AND U825 ( .A(\MODMULT2[0].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), .B(
        n688), .Z(n697) );
  IV U826 ( .A(n697), .Z(n709) );
  NOR U827 ( .A(n709), .B(n[0]), .Z(n689) );
  NAND U828 ( .A(n700), .B(n689), .Z(n690) );
  NANDN U829 ( .A(n698), .B(n690), .Z(n691) );
  AND U830 ( .A(n703), .B(n866), .Z(n712) );
  OR U831 ( .A(n691), .B(n712), .Z(n692) );
  AND U832 ( .A(n693), .B(n692), .Z(n694) );
  ANDN U833 ( .B(n695), .A(n694), .Z(n696) );
  NANDN U834 ( .A(n710), .B(n696), .Z(n723) );
  ANDN U835 ( .B(n[0]), .A(n697), .Z(n704) );
  NANDN U836 ( .A(n698), .B(n704), .Z(n699) );
  AND U837 ( .A(n700), .B(n699), .Z(n711) );
  XOR U838 ( .A(n866), .B(n711), .Z(n701) );
  NAND U839 ( .A(n723), .B(n701), .Z(n702) );
  XNOR U840 ( .A(n703), .B(n702), .Z(n742) );
  XOR U841 ( .A(n[1]), .B(n704), .Z(n705) );
  NAND U842 ( .A(n723), .B(n705), .Z(n706) );
  XNOR U843 ( .A(n707), .B(n706), .Z(n727) );
  NAND U844 ( .A(n723), .B(n[0]), .Z(n708) );
  XOR U845 ( .A(n709), .B(n708), .Z(n734) );
  ANDN U846 ( .B(n723), .A(n710), .Z(n717) );
  OR U847 ( .A(n712), .B(n711), .Z(n713) );
  AND U848 ( .A(n714), .B(n713), .Z(n721) );
  NANDN U849 ( .A(n715), .B(n721), .Z(n716) );
  AND U850 ( .A(n717), .B(n716), .Z(n718) );
  XOR U851 ( .A(n719), .B(n718), .Z(n758) );
  XOR U852 ( .A(n880), .B(n721), .Z(n722) );
  NAND U853 ( .A(n723), .B(n722), .Z(n724) );
  XNOR U854 ( .A(n725), .B(n724), .Z(n752) );
  ANDN U855 ( .B(n748), .A(n866), .Z(n743) );
  XNOR U856 ( .A(n742), .B(n743), .Z(n745) );
  NAND U857 ( .A(n[1]), .B(n748), .Z(n726) );
  NANDN U858 ( .A(n727), .B(n726), .Z(n729) );
  AND U859 ( .A(n[0]), .B(n748), .Z(n733) );
  ANDN U860 ( .B(n733), .A(n734), .Z(n732) );
  XNOR U861 ( .A(n727), .B(n726), .Z(n731) );
  NANDN U862 ( .A(n732), .B(n731), .Z(n728) );
  NAND U863 ( .A(n729), .B(n728), .Z(n744) );
  XOR U864 ( .A(n745), .B(n744), .Z(n730) );
  IV U865 ( .A(n730), .Z(n772) );
  ANDN U866 ( .B(m[3]), .A(n772), .Z(n740) );
  XOR U867 ( .A(m[3]), .B(n730), .Z(n738) );
  XOR U868 ( .A(n732), .B(n731), .Z(n764) );
  NANDN U869 ( .A(n764), .B(m[2]), .Z(n737) );
  XNOR U870 ( .A(m[2]), .B(n764), .Z(n735) );
  XOR U871 ( .A(n734), .B(n733), .Z(n766) );
  AND U872 ( .A(m[1]), .B(n766), .Z(n761) );
  NAND U873 ( .A(n735), .B(n761), .Z(n736) );
  NAND U874 ( .A(n737), .B(n736), .Z(n769) );
  AND U875 ( .A(n738), .B(n769), .Z(n739) );
  OR U876 ( .A(n740), .B(n739), .Z(n741) );
  AND U877 ( .A(n898), .B(n741), .Z(n756) );
  NANDN U878 ( .A(n743), .B(n742), .Z(n747) );
  NAND U879 ( .A(n745), .B(n744), .Z(n746) );
  NAND U880 ( .A(n747), .B(n746), .Z(n749) );
  NANDN U881 ( .A(n880), .B(n748), .Z(n751) );
  XOR U882 ( .A(n752), .B(n751), .Z(n750) );
  XNOR U883 ( .A(n749), .B(n750), .Z(n755) );
  NAND U884 ( .A(n750), .B(n749), .Z(n754) );
  NAND U885 ( .A(n752), .B(n751), .Z(n753) );
  AND U886 ( .A(n754), .B(n753), .Z(n760) );
  ANDN U887 ( .B(n756), .A(n755), .Z(n757) );
  XNOR U888 ( .A(n758), .B(n757), .Z(n759) );
  XNOR U889 ( .A(n760), .B(n759), .Z(n787) );
  NOR U890 ( .A(n786), .B(n787), .Z(n777) );
  XOR U891 ( .A(n761), .B(m[2]), .Z(n762) );
  NAND U892 ( .A(n898), .B(n762), .Z(n763) );
  XNOR U893 ( .A(n764), .B(n763), .Z(n796) );
  ANDN U894 ( .B(n866), .A(n796), .Z(n768) );
  NAND U895 ( .A(m[1]), .B(n898), .Z(n765) );
  XOR U896 ( .A(n766), .B(n765), .Z(n801) );
  OR U897 ( .A(n[1]), .B(n801), .Z(n767) );
  NANDN U898 ( .A(n768), .B(n767), .Z(n775) );
  NAND U899 ( .A(n880), .B(n866), .Z(n833) );
  XOR U900 ( .A(m[3]), .B(n769), .Z(n770) );
  NAND U901 ( .A(n898), .B(n770), .Z(n771) );
  XOR U902 ( .A(n772), .B(n771), .Z(n790) );
  NANDN U903 ( .A(n796), .B(n790), .Z(n773) );
  AND U904 ( .A(n833), .B(n773), .Z(n774) );
  ANDN U905 ( .B(n775), .A(n774), .Z(n776) );
  ANDN U906 ( .B(n777), .A(n776), .Z(n779) );
  AND U907 ( .A(n790), .B(n880), .Z(n778) );
  ANDN U908 ( .B(n779), .A(n778), .Z(n799) );
  NANDN U909 ( .A(n799), .B(n[0]), .Z(n780) );
  XNOR U910 ( .A(n781), .B(n780), .Z(n805) );
  NANDN U911 ( .A(n866), .B(n796), .Z(n784) );
  XNOR U912 ( .A(n796), .B(n866), .Z(n782) );
  NAND U913 ( .A(n[0]), .B(n781), .Z(n797) );
  NAND U914 ( .A(n782), .B(n793), .Z(n783) );
  AND U915 ( .A(n784), .B(n783), .Z(n785) );
  XNOR U916 ( .A(n[3]), .B(n785), .Z(n788) );
  NOR U917 ( .A(n843), .B(n787), .Z(n792) );
  NANDN U918 ( .A(n799), .B(n788), .Z(n789) );
  XNOR U919 ( .A(n790), .B(n789), .Z(n836) );
  NAND U920 ( .A(n880), .B(n836), .Z(n791) );
  AND U921 ( .A(n792), .B(n791), .Z(n809) );
  XNOR U922 ( .A(n866), .B(n793), .Z(n794) );
  NANDN U923 ( .A(n799), .B(n794), .Z(n795) );
  XNOR U924 ( .A(n796), .B(n795), .Z(n810) );
  XNOR U925 ( .A(n[1]), .B(n797), .Z(n798) );
  NANDN U926 ( .A(n799), .B(n798), .Z(n800) );
  XNOR U927 ( .A(n801), .B(n800), .Z(n814) );
  NANDN U928 ( .A(n866), .B(n810), .Z(n808) );
  AND U929 ( .A(n[0]), .B(n826), .Z(n804) );
  AND U930 ( .A(n805), .B(n804), .Z(n816) );
  NAND U931 ( .A(n826), .B(n[1]), .Z(n813) );
  XNOR U932 ( .A(n814), .B(n813), .Z(n815) );
  XNOR U933 ( .A(n816), .B(n815), .Z(n820) );
  XOR U934 ( .A(n803), .B(n802), .Z(n890) );
  XOR U935 ( .A(n805), .B(n804), .Z(n828) );
  ANDN U936 ( .B(m[1]), .A(n828), .Z(n821) );
  XOR U937 ( .A(n821), .B(m[2]), .Z(n806) );
  NANDN U938 ( .A(n890), .B(n806), .Z(n807) );
  XOR U939 ( .A(n820), .B(n807), .Z(n854) );
  OR U940 ( .A(n809), .B(n808), .Z(n812) );
  NAND U941 ( .A(n[2]), .B(n826), .Z(n811) );
  ANDN U942 ( .B(n811), .A(n810), .Z(n824) );
  ANDN U943 ( .B(n812), .A(n824), .Z(n823) );
  NANDN U944 ( .A(n814), .B(n813), .Z(n818) );
  NANDN U945 ( .A(n816), .B(n815), .Z(n817) );
  NAND U946 ( .A(n818), .B(n817), .Z(n822) );
  XOR U947 ( .A(n823), .B(n822), .Z(n819) );
  IV U948 ( .A(n819), .Z(n832) );
  NAND U949 ( .A(n823), .B(n822), .Z(n825) );
  ANDN U950 ( .B(n825), .A(n824), .Z(n835) );
  AND U951 ( .A(n826), .B(n[3]), .Z(n837) );
  XNOR U952 ( .A(n836), .B(n837), .Z(n834) );
  XNOR U953 ( .A(n835), .B(n834), .Z(n840) );
  XOR U954 ( .A(n841), .B(n840), .Z(n859) );
  NANDN U955 ( .A(n890), .B(m[1]), .Z(n827) );
  XOR U956 ( .A(n828), .B(n827), .Z(n853) );
  XOR U957 ( .A(m[3]), .B(n829), .Z(n830) );
  NANDN U958 ( .A(n890), .B(n830), .Z(n831) );
  XOR U959 ( .A(n832), .B(n831), .Z(n865) );
  NANDN U960 ( .A(n835), .B(n834), .Z(n839) );
  NANDN U961 ( .A(n837), .B(n836), .Z(n838) );
  AND U962 ( .A(n839), .B(n838), .Z(n845) );
  AND U963 ( .A(n841), .B(n840), .Z(n842) );
  XNOR U964 ( .A(n843), .B(n842), .Z(n844) );
  XNOR U965 ( .A(n845), .B(n844), .Z(n860) );
  NANDN U966 ( .A(n890), .B(
        \MODMULT2[0].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), .Z(n849) );
  NAND U967 ( .A(n[0]), .B(n849), .Z(n850) );
  XNOR U968 ( .A(n866), .B(n855), .Z(n846) );
  NAND U969 ( .A(n863), .B(n846), .Z(n847) );
  XNOR U970 ( .A(n854), .B(n847), .Z(n875) );
  NAND U971 ( .A(n863), .B(n[0]), .Z(n848) );
  XNOR U972 ( .A(n849), .B(n848), .Z(n892) );
  XNOR U973 ( .A(n[1]), .B(n850), .Z(n851) );
  NAND U974 ( .A(n863), .B(n851), .Z(n852) );
  XOR U975 ( .A(n853), .B(n852), .Z(n902) );
  NANDN U976 ( .A(n866), .B(n854), .Z(n858) );
  XNOR U977 ( .A(n854), .B(n866), .Z(n856) );
  NAND U978 ( .A(n856), .B(n855), .Z(n857) );
  NAND U979 ( .A(n858), .B(n857), .Z(n861) );
  XNOR U980 ( .A(n880), .B(n861), .Z(n862) );
  NAND U981 ( .A(n863), .B(n862), .Z(n864) );
  XNOR U982 ( .A(n865), .B(n864), .Z(n883) );
  AND U983 ( .A(n[0]), .B(n879), .Z(n891) );
  AND U984 ( .A(n892), .B(n891), .Z(n900) );
  AND U985 ( .A(n[1]), .B(n879), .Z(n899) );
  XNOR U986 ( .A(n875), .B(n876), .Z(n874) );
  ANDN U987 ( .B(n879), .A(n866), .Z(n873) );
  XNOR U988 ( .A(n874), .B(n873), .Z(n867) );
  NANDN U989 ( .A(n912), .B(n867), .Z(n868) );
  NAND U990 ( .A(n869), .B(n868), .Z(c[2]) );
  NAND U991 ( .A(c[2]), .B(\keep_1[0] ), .Z(n871) );
  NANDN U992 ( .A(\keep_1[0] ), .B(m[2]), .Z(n870) );
  NAND U993 ( .A(n871), .B(n870), .Z(N10) );
  NAND U994 ( .A(n872), .B(n912), .Z(n887) );
  NAND U995 ( .A(n874), .B(n873), .Z(n878) );
  NANDN U996 ( .A(n876), .B(n875), .Z(n877) );
  AND U997 ( .A(n878), .B(n877), .Z(n882) );
  NANDN U998 ( .A(n880), .B(n879), .Z(n881) );
  XNOR U999 ( .A(n882), .B(n881), .Z(n884) );
  XNOR U1000 ( .A(n884), .B(n883), .Z(n885) );
  NANDN U1001 ( .A(n912), .B(n885), .Z(n886) );
  NAND U1002 ( .A(n887), .B(n886), .Z(c[3]) );
  NAND U1003 ( .A(c[3]), .B(\keep_1[0] ), .Z(n889) );
  NANDN U1004 ( .A(\keep_1[0] ), .B(m[3]), .Z(n888) );
  NAND U1005 ( .A(n889), .B(n888), .Z(N11) );
  NANDN U1006 ( .A(n890), .B(n912), .Z(n895) );
  XNOR U1007 ( .A(n892), .B(n891), .Z(n893) );
  NANDN U1008 ( .A(n912), .B(n893), .Z(n894) );
  NAND U1009 ( .A(n895), .B(n894), .Z(c[0]) );
  NAND U1010 ( .A(c[0]), .B(\keep_1[0] ), .Z(n897) );
  NANDN U1011 ( .A(\keep_1[0] ), .B(
        \MODMULT2[0].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), .Z(n896) );
  NAND U1012 ( .A(n897), .B(n896), .Z(N8) );
  NAND U1013 ( .A(n898), .B(n912), .Z(n905) );
  XOR U1014 ( .A(n900), .B(n899), .Z(n901) );
  XNOR U1015 ( .A(n902), .B(n901), .Z(n903) );
  NANDN U1016 ( .A(n912), .B(n903), .Z(n904) );
  NAND U1017 ( .A(n905), .B(n904), .Z(c[1]) );
  NAND U1018 ( .A(c[1]), .B(\keep_1[0] ), .Z(n907) );
  NANDN U1019 ( .A(\keep_1[0] ), .B(m[1]), .Z(n906) );
  NAND U1020 ( .A(n907), .B(n906), .Z(N9) );
  ANDN U1021 ( .B(e[0]), .A(init), .Z(ein[0]) );
  NAND U1022 ( .A(ereg[1]), .B(init), .Z(n909) );
  NANDN U1023 ( .A(init), .B(e[1]), .Z(n908) );
  NAND U1024 ( .A(n909), .B(n908), .Z(ein[1]) );
  NAND U1025 ( .A(ereg[2]), .B(init), .Z(n911) );
  NANDN U1026 ( .A(init), .B(e[2]), .Z(n910) );
  NAND U1027 ( .A(n911), .B(n910), .Z(ein[2]) );
  NANDN U1028 ( .A(\keep_1[0] ), .B(n912), .Z(n3) );
endmodule

